module basic_5000_50000_5000_50_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
and U0 (N_0,In_1744,In_4781);
xnor U1 (N_1,In_427,In_4953);
nor U2 (N_2,In_1399,In_2769);
xor U3 (N_3,In_3861,In_3145);
and U4 (N_4,In_688,In_2601);
xor U5 (N_5,In_3760,In_4984);
xnor U6 (N_6,In_1803,In_1383);
xnor U7 (N_7,In_1545,In_3479);
or U8 (N_8,In_682,In_4976);
and U9 (N_9,In_2980,In_2628);
or U10 (N_10,In_4146,In_170);
nand U11 (N_11,In_557,In_2495);
or U12 (N_12,In_2213,In_1449);
or U13 (N_13,In_4552,In_4968);
nor U14 (N_14,In_2819,In_3697);
nor U15 (N_15,In_2293,In_1662);
nor U16 (N_16,In_3296,In_1024);
or U17 (N_17,In_1579,In_966);
xnor U18 (N_18,In_232,In_3657);
or U19 (N_19,In_286,In_344);
and U20 (N_20,In_2817,In_2622);
nand U21 (N_21,In_1310,In_1092);
nor U22 (N_22,In_2123,In_1936);
and U23 (N_23,In_2,In_985);
and U24 (N_24,In_4259,In_4003);
xor U25 (N_25,In_2913,In_1126);
nand U26 (N_26,In_3355,In_3088);
and U27 (N_27,In_4002,In_1627);
nand U28 (N_28,In_3465,In_536);
nor U29 (N_29,In_840,In_774);
nand U30 (N_30,In_541,In_1316);
nor U31 (N_31,In_3186,In_2954);
nor U32 (N_32,In_3124,In_289);
nor U33 (N_33,In_3680,In_3816);
xnor U34 (N_34,In_1299,In_1355);
or U35 (N_35,In_2818,In_680);
and U36 (N_36,In_4596,In_4969);
xnor U37 (N_37,In_1655,In_1526);
nand U38 (N_38,In_2221,In_4831);
xnor U39 (N_39,In_2800,In_2245);
and U40 (N_40,In_2858,In_2244);
xnor U41 (N_41,In_2488,In_1736);
or U42 (N_42,In_3298,In_3159);
xnor U43 (N_43,In_3445,In_4550);
xnor U44 (N_44,In_1287,In_821);
nand U45 (N_45,In_3315,In_1318);
nor U46 (N_46,In_1821,In_3341);
or U47 (N_47,In_3530,In_1056);
xnor U48 (N_48,In_3721,In_3609);
or U49 (N_49,In_2681,In_2162);
or U50 (N_50,In_9,In_4206);
or U51 (N_51,In_3288,In_188);
nor U52 (N_52,In_4279,In_2182);
nand U53 (N_53,In_752,In_2361);
or U54 (N_54,In_3228,In_4386);
xor U55 (N_55,In_940,In_4646);
and U56 (N_56,In_1765,In_909);
nand U57 (N_57,In_2694,In_4869);
xnor U58 (N_58,In_2515,In_19);
xor U59 (N_59,In_1238,In_2201);
and U60 (N_60,In_2815,In_4276);
or U61 (N_61,In_2352,In_1439);
xor U62 (N_62,In_2549,In_1186);
xnor U63 (N_63,In_4027,In_3417);
xor U64 (N_64,In_3224,In_1790);
nor U65 (N_65,In_1952,In_3703);
nor U66 (N_66,In_594,In_2422);
or U67 (N_67,In_2340,In_1575);
and U68 (N_68,In_3090,In_2327);
nor U69 (N_69,In_4157,In_4114);
nand U70 (N_70,In_3297,In_1137);
xor U71 (N_71,In_3193,In_1217);
or U72 (N_72,In_4963,In_1386);
and U73 (N_73,In_920,In_4494);
xor U74 (N_74,In_2696,In_3085);
nand U75 (N_75,In_3739,In_3622);
and U76 (N_76,In_2442,In_1367);
and U77 (N_77,In_746,In_2982);
and U78 (N_78,In_3049,In_1325);
xnor U79 (N_79,In_2969,In_2375);
xor U80 (N_80,In_550,In_3958);
nand U81 (N_81,In_2968,In_4632);
nor U82 (N_82,In_51,In_3755);
nand U83 (N_83,In_3521,In_4359);
nor U84 (N_84,In_2270,In_2540);
and U85 (N_85,In_851,In_2770);
nand U86 (N_86,In_3026,In_2015);
nand U87 (N_87,In_2714,In_1062);
xnor U88 (N_88,In_4294,In_4760);
or U89 (N_89,In_4881,In_4077);
xnor U90 (N_90,In_1590,In_3108);
or U91 (N_91,In_613,In_653);
or U92 (N_92,In_1068,In_3318);
nand U93 (N_93,In_3854,In_4904);
and U94 (N_94,In_4022,In_3937);
and U95 (N_95,In_2315,In_1876);
and U96 (N_96,In_1739,In_590);
nand U97 (N_97,In_4529,In_772);
and U98 (N_98,In_1650,In_3008);
nor U99 (N_99,In_4052,In_15);
and U100 (N_100,In_1670,In_110);
and U101 (N_101,In_947,In_1456);
or U102 (N_102,In_4515,In_4221);
nand U103 (N_103,In_3592,In_642);
nand U104 (N_104,In_4802,In_4830);
or U105 (N_105,In_1073,In_4698);
xor U106 (N_106,In_4567,In_1505);
or U107 (N_107,In_3178,In_2779);
nand U108 (N_108,In_3157,In_2029);
xor U109 (N_109,In_4610,In_2481);
nor U110 (N_110,In_3659,In_1695);
xor U111 (N_111,In_3652,In_506);
and U112 (N_112,In_2059,In_1281);
nand U113 (N_113,In_1511,In_1551);
or U114 (N_114,In_2144,In_4587);
nor U115 (N_115,In_74,In_2736);
nand U116 (N_116,In_914,In_2590);
nor U117 (N_117,In_4970,In_1189);
nor U118 (N_118,In_3520,In_1199);
and U119 (N_119,In_757,In_1103);
nor U120 (N_120,In_2838,In_277);
nand U121 (N_121,In_2639,In_410);
or U122 (N_122,In_4162,In_723);
nor U123 (N_123,In_3851,In_4240);
and U124 (N_124,In_4629,In_2135);
xnor U125 (N_125,In_3208,In_4798);
nand U126 (N_126,In_4859,In_860);
or U127 (N_127,In_788,In_3243);
nand U128 (N_128,In_2084,In_342);
or U129 (N_129,In_196,In_78);
and U130 (N_130,In_260,In_3316);
nand U131 (N_131,In_4109,In_1136);
nor U132 (N_132,In_2204,In_679);
nor U133 (N_133,In_3859,In_2874);
nand U134 (N_134,In_4440,In_1866);
and U135 (N_135,In_711,In_3122);
xor U136 (N_136,In_4019,In_2305);
or U137 (N_137,In_200,In_957);
xor U138 (N_138,In_1605,In_3782);
and U139 (N_139,In_3735,In_370);
nor U140 (N_140,In_4617,In_3640);
nor U141 (N_141,In_422,In_3849);
nor U142 (N_142,In_3545,In_4058);
xor U143 (N_143,In_4161,In_4991);
nor U144 (N_144,In_1753,In_625);
nand U145 (N_145,In_3738,In_4250);
nor U146 (N_146,In_3292,In_4996);
nor U147 (N_147,In_2768,In_2808);
and U148 (N_148,In_4813,In_535);
nand U149 (N_149,In_2928,In_1586);
or U150 (N_150,In_1324,In_2598);
xor U151 (N_151,In_2740,In_935);
xnor U152 (N_152,In_34,In_831);
nand U153 (N_153,In_160,In_810);
xor U154 (N_154,In_3671,In_522);
xor U155 (N_155,In_3528,In_1442);
nor U156 (N_156,In_82,In_1606);
nand U157 (N_157,In_3940,In_1672);
nand U158 (N_158,In_234,In_1100);
nand U159 (N_159,In_2259,In_2518);
and U160 (N_160,In_1241,In_2406);
and U161 (N_161,In_4224,In_2618);
nand U162 (N_162,In_2919,In_1413);
and U163 (N_163,In_4305,In_3718);
nor U164 (N_164,In_1444,In_2658);
and U165 (N_165,In_1969,In_3063);
or U166 (N_166,In_2712,In_2003);
xor U167 (N_167,In_849,In_3836);
nor U168 (N_168,In_2955,In_4731);
xnor U169 (N_169,In_3134,In_990);
xnor U170 (N_170,In_3955,In_1888);
nand U171 (N_171,In_1289,In_458);
xor U172 (N_172,In_1539,In_2137);
nor U173 (N_173,In_2234,In_2828);
xor U174 (N_174,In_2594,In_166);
and U175 (N_175,In_4643,In_566);
xnor U176 (N_176,In_1990,In_3077);
or U177 (N_177,In_4964,In_1194);
and U178 (N_178,In_1038,In_1081);
nand U179 (N_179,In_4193,In_3792);
or U180 (N_180,In_3757,In_1378);
nor U181 (N_181,In_4809,In_306);
nor U182 (N_182,In_3919,In_464);
xnor U183 (N_183,In_1019,In_2847);
or U184 (N_184,In_4310,In_777);
xor U185 (N_185,In_1686,In_1981);
xor U186 (N_186,In_3686,In_2755);
or U187 (N_187,In_2957,In_2239);
nor U188 (N_188,In_367,In_1554);
and U189 (N_189,In_4764,In_2931);
nor U190 (N_190,In_2366,In_4761);
xor U191 (N_191,In_3751,In_3429);
or U192 (N_192,In_2429,In_4825);
or U193 (N_193,In_433,In_162);
or U194 (N_194,In_205,In_2306);
nand U195 (N_195,In_319,In_2855);
xor U196 (N_196,In_339,In_4481);
and U197 (N_197,In_4675,In_2039);
nand U198 (N_198,In_4907,In_4269);
or U199 (N_199,In_2412,In_3843);
or U200 (N_200,In_1577,In_3889);
xnor U201 (N_201,In_2972,In_3804);
nor U202 (N_202,In_4464,In_4076);
nor U203 (N_203,In_1302,In_3013);
and U204 (N_204,In_3881,In_3428);
xnor U205 (N_205,In_4799,In_3991);
nor U206 (N_206,In_2932,In_3375);
nor U207 (N_207,In_2258,In_925);
and U208 (N_208,In_3020,In_2216);
nor U209 (N_209,In_2977,In_197);
and U210 (N_210,In_3709,In_3299);
xnor U211 (N_211,In_4362,In_1935);
nand U212 (N_212,In_948,In_4068);
nor U213 (N_213,In_2192,In_2876);
and U214 (N_214,In_4364,In_2583);
xor U215 (N_215,In_2981,In_2921);
nor U216 (N_216,In_3708,In_95);
or U217 (N_217,In_4080,In_1967);
or U218 (N_218,In_4028,In_2906);
and U219 (N_219,In_2537,In_4349);
xor U220 (N_220,In_4167,In_989);
or U221 (N_221,In_1342,In_304);
and U222 (N_222,In_3486,In_4606);
and U223 (N_223,In_537,In_1770);
nor U224 (N_224,In_4278,In_3207);
nor U225 (N_225,In_4605,In_2675);
nand U226 (N_226,In_3339,In_1298);
or U227 (N_227,In_3372,In_4918);
and U228 (N_228,In_4820,In_4067);
or U229 (N_229,In_3019,In_3311);
nand U230 (N_230,In_1761,In_800);
or U231 (N_231,In_4381,In_146);
nor U232 (N_232,In_2298,In_2302);
and U233 (N_233,In_4674,In_2099);
or U234 (N_234,In_2215,In_766);
or U235 (N_235,In_1400,In_73);
nor U236 (N_236,In_3052,In_1360);
nand U237 (N_237,In_2742,In_3456);
nand U238 (N_238,In_55,In_2734);
and U239 (N_239,In_136,In_1313);
nor U240 (N_240,In_2942,In_8);
or U241 (N_241,In_4709,In_2431);
nand U242 (N_242,In_2196,In_3745);
nor U243 (N_243,In_2979,In_1003);
nand U244 (N_244,In_3396,In_4916);
or U245 (N_245,In_2348,In_296);
and U246 (N_246,In_3129,In_3506);
nand U247 (N_247,In_1276,In_4630);
and U248 (N_248,In_4326,In_3332);
nor U249 (N_249,In_4782,In_1645);
and U250 (N_250,In_111,In_1564);
nand U251 (N_251,In_4480,In_4465);
nor U252 (N_252,In_4062,In_3131);
nor U253 (N_253,In_4443,In_2297);
and U254 (N_254,In_237,In_4817);
and U255 (N_255,In_4286,In_3409);
nor U256 (N_256,In_1283,In_2606);
nand U257 (N_257,In_1164,In_4090);
or U258 (N_258,In_4424,In_3571);
nand U259 (N_259,In_4780,In_1948);
and U260 (N_260,In_1393,In_1291);
nor U261 (N_261,In_316,In_3631);
nand U262 (N_262,In_2507,In_262);
and U263 (N_263,In_3998,In_1249);
nor U264 (N_264,In_4733,In_4473);
nor U265 (N_265,In_4974,In_2023);
xnor U266 (N_266,In_2459,In_4860);
nor U267 (N_267,In_2061,In_66);
xnor U268 (N_268,In_2745,In_4582);
and U269 (N_269,In_2242,In_2220);
nor U270 (N_270,In_953,In_4336);
and U271 (N_271,In_4982,In_1934);
nor U272 (N_272,In_3661,In_693);
or U273 (N_273,In_2255,In_2994);
nand U274 (N_274,In_4599,In_3083);
xnor U275 (N_275,In_3407,In_2247);
or U276 (N_276,In_159,In_3365);
nor U277 (N_277,In_3149,In_1565);
xor U278 (N_278,In_2308,In_4422);
nand U279 (N_279,In_2822,In_1885);
or U280 (N_280,In_4046,In_823);
and U281 (N_281,In_3608,In_2797);
or U282 (N_282,In_4367,In_3139);
or U283 (N_283,In_3029,In_1788);
or U284 (N_284,In_3320,In_1580);
xor U285 (N_285,In_4382,In_3256);
nand U286 (N_286,In_1917,In_184);
or U287 (N_287,In_3076,In_448);
nor U288 (N_288,In_2299,In_3408);
and U289 (N_289,In_259,In_890);
or U290 (N_290,In_3378,In_3534);
or U291 (N_291,In_2591,In_3754);
or U292 (N_292,In_2288,In_4639);
and U293 (N_293,In_23,In_2365);
xnor U294 (N_294,In_2186,In_3691);
and U295 (N_295,In_819,In_4086);
nor U296 (N_296,In_4118,In_2376);
nand U297 (N_297,In_2542,In_1746);
nand U298 (N_298,In_127,In_1905);
nand U299 (N_299,In_2564,In_1729);
or U300 (N_300,In_2814,In_1951);
and U301 (N_301,In_4670,In_1516);
and U302 (N_302,In_629,In_2859);
xnor U303 (N_303,In_4999,In_1576);
and U304 (N_304,In_4393,In_2014);
and U305 (N_305,In_3404,In_507);
or U306 (N_306,In_3823,In_3100);
or U307 (N_307,In_4958,In_2063);
nand U308 (N_308,In_968,In_689);
nand U309 (N_309,In_218,In_123);
and U310 (N_310,In_3471,In_1849);
xnor U311 (N_311,In_4031,In_3639);
xnor U312 (N_312,In_2320,In_266);
nand U313 (N_313,In_3477,In_1110);
nor U314 (N_314,In_931,In_3112);
xnor U315 (N_315,In_3130,In_3566);
or U316 (N_316,In_2571,In_1151);
and U317 (N_317,In_2790,In_632);
nor U318 (N_318,In_3061,In_4654);
or U319 (N_319,In_1895,In_1085);
and U320 (N_320,In_326,In_3786);
nand U321 (N_321,In_1608,In_2539);
xnor U322 (N_322,In_3656,In_203);
and U323 (N_323,In_1070,In_1013);
nor U324 (N_324,In_4477,In_1387);
nand U325 (N_325,In_426,In_3234);
nand U326 (N_326,In_2316,In_2881);
nor U327 (N_327,In_1230,In_3384);
nand U328 (N_328,In_4729,In_4705);
nand U329 (N_329,In_855,In_912);
nor U330 (N_330,In_3988,In_133);
and U331 (N_331,In_3437,In_4322);
and U332 (N_332,In_3969,In_939);
nor U333 (N_333,In_4363,In_1420);
xnor U334 (N_334,In_1163,In_1180);
nand U335 (N_335,In_279,In_1688);
or U336 (N_336,In_2716,In_4213);
nor U337 (N_337,In_1540,In_532);
nor U338 (N_338,In_3478,In_3964);
nor U339 (N_339,In_2663,In_3865);
or U340 (N_340,In_1370,In_3719);
xor U341 (N_341,In_3853,In_2816);
or U342 (N_342,In_1010,In_871);
nand U343 (N_343,In_4434,In_3189);
and U344 (N_344,In_798,In_4516);
xnor U345 (N_345,In_239,In_4502);
xor U346 (N_346,In_1896,In_2230);
or U347 (N_347,In_2036,In_4898);
nand U348 (N_348,In_3303,In_2494);
xnor U349 (N_349,In_4750,In_1220);
or U350 (N_350,In_3993,In_4343);
nor U351 (N_351,In_431,In_3831);
and U352 (N_352,In_4255,In_4472);
nor U353 (N_353,In_3504,In_2056);
nor U354 (N_354,In_57,In_1705);
or U355 (N_355,In_1837,In_1634);
nor U356 (N_356,In_4660,In_4191);
nor U357 (N_357,In_2492,In_2538);
nand U358 (N_358,In_984,In_3539);
and U359 (N_359,In_2866,In_2053);
or U360 (N_360,In_3573,In_4132);
and U361 (N_361,In_1156,In_4330);
xor U362 (N_362,In_1963,In_44);
nand U363 (N_363,In_4693,In_3280);
nand U364 (N_364,In_4720,In_4956);
and U365 (N_365,In_4688,In_2108);
nor U366 (N_366,In_4864,In_898);
and U367 (N_367,In_2393,In_2892);
or U368 (N_368,In_119,In_404);
xnor U369 (N_369,In_1904,In_157);
nor U370 (N_370,In_3595,In_3440);
nand U371 (N_371,In_4694,In_71);
and U372 (N_372,In_4774,In_1247);
and U373 (N_373,In_395,In_1315);
and U374 (N_374,In_4112,In_4198);
nor U375 (N_375,In_2565,In_3283);
nor U376 (N_376,In_4843,In_1831);
xor U377 (N_377,In_2392,In_3784);
nand U378 (N_378,In_1450,In_2134);
or U379 (N_379,In_3644,In_84);
and U380 (N_380,In_3434,In_2952);
or U381 (N_381,In_1512,In_895);
and U382 (N_382,In_908,In_4274);
or U383 (N_383,In_2498,In_503);
or U384 (N_384,In_1914,In_2737);
nand U385 (N_385,In_1433,In_4572);
or U386 (N_386,In_3514,In_1219);
nand U387 (N_387,In_3097,In_3069);
and U388 (N_388,In_4656,In_4789);
xnor U389 (N_389,In_2075,In_1543);
or U390 (N_390,In_4538,In_893);
xor U391 (N_391,In_4983,In_280);
and U392 (N_392,In_1028,In_4337);
or U393 (N_393,In_2852,In_4862);
or U394 (N_394,In_4350,In_2472);
nor U395 (N_395,In_2350,In_4758);
xor U396 (N_396,In_4426,In_1784);
and U397 (N_397,In_3240,In_2555);
and U398 (N_398,In_3126,In_2080);
or U399 (N_399,In_3327,In_3676);
or U400 (N_400,In_420,In_222);
nor U401 (N_401,In_3229,In_4297);
and U402 (N_402,In_785,In_121);
nand U403 (N_403,In_3003,In_2501);
nand U404 (N_404,In_685,In_4923);
xnor U405 (N_405,In_2129,In_94);
nand U406 (N_406,In_2959,In_4535);
or U407 (N_407,In_2657,In_1776);
or U408 (N_408,In_1020,In_523);
nand U409 (N_409,In_3802,In_1411);
nor U410 (N_410,In_4779,In_4770);
and U411 (N_411,In_1679,In_1593);
nor U412 (N_412,In_951,In_2926);
xnor U413 (N_413,In_716,In_2068);
xor U414 (N_414,In_3577,In_1232);
nor U415 (N_415,In_4395,In_4264);
nand U416 (N_416,In_3930,In_4586);
nor U417 (N_417,In_4275,In_274);
or U418 (N_418,In_4858,In_3681);
nor U419 (N_419,In_3732,In_804);
or U420 (N_420,In_884,In_1932);
nor U421 (N_421,In_4827,In_3574);
or U422 (N_422,In_11,In_667);
or U423 (N_423,In_718,In_1827);
nor U424 (N_424,In_906,In_4773);
nand U425 (N_425,In_1716,In_4555);
nand U426 (N_426,In_1804,In_1359);
or U427 (N_427,In_60,In_3634);
or U428 (N_428,In_1350,In_4889);
or U429 (N_429,In_3326,In_915);
nand U430 (N_430,In_4836,In_4174);
or U431 (N_431,In_1692,In_421);
or U432 (N_432,In_3450,In_4111);
nor U433 (N_433,In_2741,In_325);
and U434 (N_434,In_4549,In_2190);
nor U435 (N_435,In_3822,In_4501);
nor U436 (N_436,In_4792,In_4253);
or U437 (N_437,In_567,In_3394);
and U438 (N_438,In_1084,In_1527);
and U439 (N_439,In_2329,In_608);
nand U440 (N_440,In_1182,In_206);
xor U441 (N_441,In_1996,In_3887);
and U442 (N_442,In_2575,In_3977);
xor U443 (N_443,In_2191,In_4919);
xnor U444 (N_444,In_4875,In_4565);
nor U445 (N_445,In_240,In_3057);
nand U446 (N_446,In_3864,In_551);
nor U447 (N_447,In_1780,In_3314);
nand U448 (N_448,In_2567,In_1703);
nand U449 (N_449,In_4876,In_930);
and U450 (N_450,In_1382,In_1177);
nand U451 (N_451,In_712,In_4292);
and U452 (N_452,In_1883,In_2281);
xnor U453 (N_453,In_2856,In_41);
xor U454 (N_454,In_243,In_3120);
nor U455 (N_455,In_2304,In_322);
and U456 (N_456,In_5,In_4060);
or U457 (N_457,In_4436,In_1920);
or U458 (N_458,In_4676,In_1025);
nor U459 (N_459,In_2698,In_1001);
or U460 (N_460,In_3218,In_2976);
or U461 (N_461,In_3105,In_3074);
or U462 (N_462,In_1998,In_1596);
and U463 (N_463,In_379,In_134);
nor U464 (N_464,In_543,In_2707);
nand U465 (N_465,In_2222,In_4070);
and U466 (N_466,In_651,In_4690);
nand U467 (N_467,In_3679,In_4220);
and U468 (N_468,In_854,In_3089);
nand U469 (N_469,In_4728,In_2967);
xor U470 (N_470,In_3908,In_3948);
nor U471 (N_471,In_868,In_635);
nand U472 (N_472,In_3589,In_1353);
nand U473 (N_473,In_2608,In_1436);
nand U474 (N_474,In_4208,In_378);
or U475 (N_475,In_1203,In_684);
or U476 (N_476,In_1262,In_3321);
xor U477 (N_477,In_4469,In_181);
or U478 (N_478,In_2659,In_2451);
and U479 (N_479,In_338,In_3337);
or U480 (N_480,In_2898,In_1144);
and U481 (N_481,In_3322,In_1079);
xnor U482 (N_482,In_903,In_2197);
or U483 (N_483,In_666,In_68);
or U484 (N_484,In_1987,In_2795);
nor U485 (N_485,In_1314,In_1758);
nor U486 (N_486,In_2851,In_2971);
nand U487 (N_487,In_2027,In_3929);
nand U488 (N_488,In_3230,In_3611);
nand U489 (N_489,In_2593,In_1838);
and U490 (N_490,In_2343,In_250);
and U491 (N_491,In_2307,In_3250);
or U492 (N_492,In_3770,In_315);
nor U493 (N_493,In_3737,In_4929);
nand U494 (N_494,In_4245,In_1653);
xor U495 (N_495,In_2098,In_2699);
or U496 (N_496,In_3340,In_1042);
or U497 (N_497,In_750,In_2223);
nand U498 (N_498,In_369,In_4937);
nand U499 (N_499,In_4828,In_2342);
xnor U500 (N_500,In_4768,In_209);
nor U501 (N_501,In_3890,In_570);
nor U502 (N_502,In_4569,In_1534);
and U503 (N_503,In_4287,In_3127);
nor U504 (N_504,In_681,In_1466);
xnor U505 (N_505,In_2689,In_958);
or U506 (N_506,In_476,In_591);
nand U507 (N_507,In_1850,In_1021);
nand U508 (N_508,In_1226,In_4551);
nor U509 (N_509,In_2560,In_1982);
and U510 (N_510,In_1926,In_1529);
xor U511 (N_511,In_690,In_4176);
xor U512 (N_512,In_4725,In_1810);
and U513 (N_513,In_4797,In_2878);
nand U514 (N_514,In_1423,In_1616);
xor U515 (N_515,In_36,In_4204);
nand U516 (N_516,In_29,In_1799);
nor U517 (N_517,In_4769,In_1395);
or U518 (N_518,In_4329,In_3841);
and U519 (N_519,In_1162,In_3674);
nand U520 (N_520,In_2332,In_4749);
and U521 (N_521,In_4513,In_4236);
or U522 (N_522,In_2408,In_4718);
nand U523 (N_523,In_1970,In_658);
or U524 (N_524,In_3349,In_2579);
nand U525 (N_525,In_3564,In_4965);
nor U526 (N_526,In_3979,In_3377);
xor U527 (N_527,In_118,In_1334);
nand U528 (N_528,In_2566,In_2106);
or U529 (N_529,In_4029,In_1246);
nand U530 (N_530,In_3030,In_732);
or U531 (N_531,In_1778,In_727);
xnor U532 (N_532,In_4104,In_4971);
nand U533 (N_533,In_1928,In_2941);
or U534 (N_534,In_1652,In_471);
and U535 (N_535,In_3148,In_2469);
nor U536 (N_536,In_4576,In_2026);
or U537 (N_537,In_4906,In_70);
nand U538 (N_538,In_3848,In_455);
nand U539 (N_539,In_3232,In_381);
xnor U540 (N_540,In_1421,In_413);
and U541 (N_541,In_26,In_1547);
and U542 (N_542,In_2863,In_2367);
xnor U543 (N_543,In_3420,In_4812);
xnor U544 (N_544,In_3548,In_2394);
nor U545 (N_545,In_238,In_2973);
or U546 (N_546,In_2044,In_3418);
nor U547 (N_547,In_3594,In_1721);
xor U548 (N_548,In_425,In_284);
or U549 (N_549,In_140,In_1394);
or U550 (N_550,In_2224,In_4214);
or U551 (N_551,In_4554,In_4416);
nor U552 (N_552,In_3916,In_2368);
and U553 (N_553,In_3258,In_2541);
nor U554 (N_554,In_2377,In_3800);
nand U555 (N_555,In_79,In_115);
nand U556 (N_556,In_4891,In_1694);
nand U557 (N_557,In_4852,In_3812);
nor U558 (N_558,In_1069,In_2651);
and U559 (N_559,In_4883,In_3794);
nand U560 (N_560,In_4272,In_2490);
nor U561 (N_561,In_3414,In_714);
nand U562 (N_562,In_3362,In_4324);
and U563 (N_563,In_65,In_796);
and U564 (N_564,In_2918,In_4835);
nor U565 (N_565,In_944,In_2465);
or U566 (N_566,In_3987,In_3704);
nand U567 (N_567,In_3617,In_4189);
and U568 (N_568,In_2263,In_3162);
nand U569 (N_569,In_526,In_3559);
and U570 (N_570,In_2167,In_2067);
nor U571 (N_571,In_457,In_1889);
nor U572 (N_572,In_3426,In_1735);
or U573 (N_573,In_2140,In_1133);
xor U574 (N_574,In_3809,In_1641);
and U575 (N_575,In_4517,In_1253);
xnor U576 (N_576,In_4137,In_2319);
or U577 (N_577,In_1875,In_3878);
nand U578 (N_578,In_3798,In_1724);
nor U579 (N_579,In_4173,In_4702);
nand U580 (N_580,In_1345,In_2206);
nor U581 (N_581,In_2912,In_2474);
nand U582 (N_582,In_4861,In_3926);
and U583 (N_583,In_4180,In_3210);
nand U584 (N_584,In_4377,In_2253);
nor U585 (N_585,In_4402,In_867);
nor U586 (N_586,In_923,In_4893);
nor U587 (N_587,In_4897,In_2886);
xor U588 (N_588,In_2232,In_4701);
nand U589 (N_589,In_69,In_3845);
or U590 (N_590,In_1012,In_1971);
or U591 (N_591,In_2616,In_2387);
or U592 (N_592,In_2599,In_4231);
nor U593 (N_593,In_1451,In_2425);
nand U594 (N_594,In_1897,In_2916);
xor U595 (N_595,In_4839,In_2662);
nand U596 (N_596,In_4475,In_3984);
xor U597 (N_597,In_3204,In_1496);
nand U598 (N_598,In_4973,In_4360);
xor U599 (N_599,In_2849,In_2523);
and U600 (N_600,In_139,In_17);
and U601 (N_601,In_3764,In_678);
nor U602 (N_602,In_3275,In_2750);
and U603 (N_603,In_4662,In_3923);
xor U604 (N_604,In_2677,In_4564);
nor U605 (N_605,In_962,In_4354);
and U606 (N_606,In_4047,In_2043);
xnor U607 (N_607,In_671,In_644);
or U608 (N_608,In_1720,In_3423);
or U609 (N_609,In_3892,In_4966);
and U610 (N_610,In_683,In_3761);
xor U611 (N_611,In_4412,In_538);
nand U612 (N_612,In_2497,In_1504);
nand U613 (N_613,In_4369,In_1515);
nor U614 (N_614,In_88,In_1484);
nand U615 (N_615,In_875,In_1448);
nand U616 (N_616,In_1054,In_1294);
nor U617 (N_617,In_1809,In_3808);
or U618 (N_618,In_1159,In_3701);
or U619 (N_619,In_934,In_372);
nor U620 (N_620,In_847,In_1854);
nor U621 (N_621,In_4410,In_938);
nand U622 (N_622,In_4810,In_1552);
and U623 (N_623,In_3035,In_3181);
xnor U624 (N_624,In_332,In_1045);
or U625 (N_625,In_1664,In_520);
nor U626 (N_626,In_3785,In_2766);
and U627 (N_627,In_3358,In_2500);
and U628 (N_628,In_288,In_4506);
or U629 (N_629,In_2019,In_4800);
or U630 (N_630,In_1431,In_2935);
nand U631 (N_631,In_3082,In_972);
and U632 (N_632,In_3529,In_217);
or U633 (N_633,In_892,In_853);
or U634 (N_634,In_1106,In_3222);
nand U635 (N_635,In_3614,In_1535);
nand U636 (N_636,In_3796,In_3813);
nor U637 (N_637,In_956,In_2672);
and U638 (N_638,In_2034,In_438);
nand U639 (N_639,In_2121,In_813);
nor U640 (N_640,In_3788,In_3301);
nor U641 (N_641,In_2759,In_3006);
and U642 (N_642,In_517,In_3253);
xnor U643 (N_643,In_362,In_1901);
nor U644 (N_644,In_3510,In_129);
nand U645 (N_645,In_2482,In_470);
nor U646 (N_646,In_3966,In_4653);
xor U647 (N_647,In_4263,In_3155);
or U648 (N_648,In_4219,In_2811);
and U649 (N_649,In_1869,In_1048);
and U650 (N_650,In_3689,In_3868);
or U651 (N_651,In_2841,In_835);
or U652 (N_652,In_2054,In_2165);
nand U653 (N_653,In_1902,In_3675);
or U654 (N_654,In_1710,In_3982);
nor U655 (N_655,In_4061,In_576);
or U656 (N_656,In_3163,In_4442);
or U657 (N_657,In_2194,In_564);
nand U658 (N_658,In_4571,In_4722);
nand U659 (N_659,In_3501,In_2411);
nor U660 (N_660,In_2827,In_3169);
xor U661 (N_661,In_3424,In_3620);
and U662 (N_662,In_3435,In_1786);
xor U663 (N_663,In_4331,In_54);
and U664 (N_664,In_2509,In_2691);
nor U665 (N_665,In_169,In_3206);
and U666 (N_666,In_2141,In_4697);
or U667 (N_667,In_1624,In_148);
xnor U668 (N_668,In_619,In_607);
and U669 (N_669,In_444,In_3427);
and U670 (N_670,In_4099,In_2173);
nand U671 (N_671,In_1819,In_3055);
or U672 (N_672,In_4030,In_1629);
xnor U673 (N_673,In_1884,In_2910);
or U674 (N_674,In_2520,In_2205);
xor U675 (N_675,In_2163,In_4452);
and U676 (N_676,In_3343,In_707);
and U677 (N_677,In_3586,In_3072);
nand U678 (N_678,In_1043,In_2286);
or U679 (N_679,In_2939,In_67);
or U680 (N_680,In_3464,In_4265);
nor U681 (N_681,In_2810,In_3905);
nand U682 (N_682,In_1430,In_3654);
xnor U683 (N_683,In_1254,In_124);
and U684 (N_684,In_147,In_351);
and U685 (N_685,In_1782,In_4703);
and U686 (N_686,In_1822,In_1317);
xor U687 (N_687,In_3482,In_1007);
nor U688 (N_688,In_2452,In_2953);
nor U689 (N_689,In_3176,In_449);
nand U690 (N_690,In_2788,In_3266);
nor U691 (N_691,In_4225,In_320);
nor U692 (N_692,In_278,In_2004);
and U693 (N_693,In_1832,In_3273);
or U694 (N_694,In_3313,In_4009);
nand U695 (N_695,In_2728,In_1726);
nor U696 (N_696,In_2240,In_3983);
nand U697 (N_697,In_3160,In_4372);
nand U698 (N_698,In_1892,In_1417);
xnor U699 (N_699,In_827,In_4691);
nand U700 (N_700,In_4902,In_528);
nor U701 (N_701,In_937,In_4500);
and U702 (N_702,In_4420,In_3819);
nand U703 (N_703,In_4730,In_3835);
nor U704 (N_704,In_435,In_3436);
xor U705 (N_705,In_3852,In_1792);
nor U706 (N_706,In_1145,In_3128);
nor U707 (N_707,In_263,In_933);
and U708 (N_708,In_2517,In_3663);
and U709 (N_709,In_2966,In_3491);
xnor U710 (N_710,In_1916,In_4612);
and U711 (N_711,In_329,In_3306);
xor U712 (N_712,In_4144,In_806);
nor U713 (N_713,In_866,In_4977);
xnor U714 (N_714,In_2374,In_4578);
or U715 (N_715,In_4147,In_4742);
or U716 (N_716,In_2479,In_3259);
nor U717 (N_717,In_2420,In_973);
nor U718 (N_718,In_1853,In_2391);
xnor U719 (N_719,In_1609,In_3877);
and U720 (N_720,In_2680,In_829);
nor U721 (N_721,In_1057,In_2218);
nor U722 (N_722,In_548,In_2762);
nand U723 (N_723,In_611,In_2552);
and U724 (N_724,In_2199,In_360);
and U725 (N_725,In_397,In_3950);
or U726 (N_726,In_2546,In_561);
nor U727 (N_727,In_2568,In_4379);
and U728 (N_728,In_373,In_3197);
and U729 (N_729,In_225,In_1894);
nor U730 (N_730,In_3746,In_531);
xor U731 (N_731,In_4095,In_4153);
or U732 (N_732,In_3125,In_1635);
nand U733 (N_733,In_3469,In_4280);
or U734 (N_734,In_1063,In_4358);
nor U735 (N_735,In_1994,In_4498);
and U736 (N_736,In_2867,In_4462);
nor U737 (N_737,In_461,In_1728);
nand U738 (N_738,In_3274,In_2217);
and U739 (N_739,In_2437,In_406);
nand U740 (N_740,In_4975,In_27);
nand U741 (N_741,In_3276,In_1312);
nand U742 (N_742,In_1800,In_4986);
or U743 (N_743,In_1229,In_4863);
and U744 (N_744,In_4928,In_822);
xor U745 (N_745,In_24,In_2399);
nor U746 (N_746,In_490,In_1260);
nand U747 (N_747,In_3619,In_4115);
nand U748 (N_748,In_1548,In_4524);
and U749 (N_749,In_1129,In_2850);
nor U750 (N_750,In_4409,In_285);
nor U751 (N_751,In_3121,In_2547);
nor U752 (N_752,In_4739,In_1371);
or U753 (N_753,In_3585,In_1755);
nand U754 (N_754,In_1587,In_64);
nor U755 (N_755,In_3220,In_1975);
nand U756 (N_756,In_4271,In_3387);
nor U757 (N_757,In_1893,In_2081);
nor U758 (N_758,In_2559,In_3934);
nand U759 (N_759,In_3810,In_1519);
nor U760 (N_760,In_3227,In_2002);
or U761 (N_761,In_2073,In_2100);
and U762 (N_762,In_4327,In_2773);
nor U763 (N_763,In_4595,In_1508);
xor U764 (N_764,In_3269,In_2661);
or U765 (N_765,In_1076,In_3214);
or U766 (N_766,In_3507,In_1111);
and U767 (N_767,In_4015,In_3123);
or U768 (N_768,In_3028,In_2301);
and U769 (N_769,In_4542,In_1737);
or U770 (N_770,In_2296,In_3711);
and U771 (N_771,In_2620,In_4788);
nand U772 (N_772,In_2991,In_4133);
and U773 (N_773,In_1006,In_1960);
and U774 (N_774,In_4121,In_4447);
nor U775 (N_775,In_3138,In_3281);
nor U776 (N_776,In_1094,In_983);
or U777 (N_777,In_3772,In_2285);
nand U778 (N_778,In_4021,In_2256);
or U779 (N_779,In_2122,In_1956);
or U780 (N_780,In_1676,In_877);
xor U781 (N_781,In_2709,In_4757);
nand U782 (N_782,In_3896,In_477);
xor U783 (N_783,In_4915,In_4601);
nand U784 (N_784,In_459,In_3135);
or U785 (N_785,In_163,In_1175);
xor U786 (N_786,In_2962,In_4527);
nand U787 (N_787,In_4140,In_737);
nand U788 (N_788,In_334,In_1107);
and U789 (N_789,In_1067,In_1120);
nand U790 (N_790,In_4400,In_3565);
xor U791 (N_791,In_3295,In_1480);
and U792 (N_792,In_1210,In_636);
or U793 (N_793,In_4190,In_778);
xor U794 (N_794,In_857,In_2754);
nand U795 (N_795,In_1255,In_988);
xnor U796 (N_796,In_1528,In_4135);
nand U797 (N_797,In_4608,In_1460);
nand U798 (N_798,In_33,In_3187);
or U799 (N_799,In_356,In_483);
or U800 (N_800,In_2102,In_2776);
nor U801 (N_801,In_4487,In_56);
or U802 (N_802,In_1647,In_1447);
nand U803 (N_803,In_1797,In_3094);
xor U804 (N_804,In_709,In_2702);
and U805 (N_805,In_630,In_1698);
and U806 (N_806,In_2619,In_45);
and U807 (N_807,In_4390,In_4223);
or U808 (N_808,In_2600,In_809);
or U809 (N_809,In_2048,In_4281);
xor U810 (N_810,In_4952,In_2064);
nor U811 (N_811,In_400,In_1581);
xor U812 (N_812,In_826,In_2664);
or U813 (N_813,In_3168,In_2085);
nand U814 (N_814,In_4584,In_4508);
and U815 (N_815,In_1116,In_4621);
and U816 (N_816,In_1125,In_950);
and U817 (N_817,In_3492,In_1392);
or U818 (N_818,In_4183,In_3673);
xor U819 (N_819,In_2556,In_2860);
or U820 (N_820,In_1099,In_574);
xnor U821 (N_821,In_1979,In_4634);
xor U822 (N_822,In_584,In_276);
nor U823 (N_823,In_2115,In_3699);
or U824 (N_824,In_3357,In_3004);
nand U825 (N_825,In_2901,In_3544);
nor U826 (N_826,In_575,In_2321);
and U827 (N_827,In_3402,In_1514);
nor U828 (N_828,In_224,In_1993);
nor U829 (N_829,In_2103,In_2292);
xnor U830 (N_830,In_3669,In_572);
nand U831 (N_831,In_643,In_4560);
nor U832 (N_832,In_323,In_1168);
nand U833 (N_833,In_1510,In_641);
nand U834 (N_834,In_2569,In_1135);
nor U835 (N_835,In_3883,In_4865);
or U836 (N_836,In_2782,In_4719);
nand U837 (N_837,In_1617,In_3194);
and U838 (N_838,In_3971,In_1864);
nand U839 (N_839,In_542,In_2380);
xnor U840 (N_840,In_2865,In_3448);
xor U841 (N_841,In_1090,In_1071);
or U842 (N_842,In_2584,In_4439);
and U843 (N_843,In_2386,In_1890);
xor U844 (N_844,In_4394,In_3744);
or U845 (N_845,In_2829,In_2409);
nor U846 (N_846,In_1621,In_30);
xor U847 (N_847,In_3215,In_4127);
nor U848 (N_848,In_2927,In_1366);
or U849 (N_849,In_1829,In_4683);
or U850 (N_850,In_1491,In_3512);
xor U851 (N_851,In_177,In_4783);
or U852 (N_852,In_53,In_1487);
nand U853 (N_853,In_3524,In_1083);
xnor U854 (N_854,In_1187,In_301);
nand U855 (N_855,In_2096,In_2463);
xor U856 (N_856,In_830,In_248);
and U857 (N_857,In_2438,In_227);
nor U858 (N_858,In_3540,In_2627);
and U859 (N_859,In_946,In_4428);
nor U860 (N_860,In_1681,In_3068);
and U861 (N_861,In_4514,In_1331);
nand U862 (N_862,In_3364,In_272);
xnor U863 (N_863,In_37,In_3683);
xnor U864 (N_864,In_1416,In_4832);
or U865 (N_865,In_1455,In_1265);
or U866 (N_866,In_4961,In_3570);
xnor U867 (N_867,In_4192,In_3925);
nor U868 (N_868,In_495,In_1174);
nor U869 (N_869,In_2534,In_2630);
nor U870 (N_870,In_1016,In_588);
and U871 (N_871,In_1861,In_2330);
nor U872 (N_872,In_1477,In_861);
or U873 (N_873,In_4681,In_4237);
and U874 (N_874,In_3990,In_592);
and U875 (N_875,In_1858,In_4154);
or U876 (N_876,In_2870,In_949);
nor U877 (N_877,In_3547,In_4035);
and U878 (N_878,In_4609,In_3141);
or U879 (N_879,In_1055,In_3444);
xor U880 (N_880,In_489,In_770);
xnor U881 (N_881,In_1155,In_467);
or U882 (N_882,In_2249,In_2832);
nand U883 (N_883,In_1404,In_4563);
nand U884 (N_884,In_109,In_4631);
and U885 (N_885,In_4945,In_3118);
xor U886 (N_886,In_4593,In_4597);
nor U887 (N_887,In_1005,In_350);
nand U888 (N_888,In_4922,In_154);
or U889 (N_889,In_1855,In_2903);
nor U890 (N_890,In_878,In_3264);
nand U891 (N_891,In_2890,In_3027);
nor U892 (N_892,In_1874,In_1127);
and U893 (N_893,In_1984,In_1147);
xnor U894 (N_894,In_1305,In_4184);
and U895 (N_895,In_452,In_4557);
nand U896 (N_896,In_2456,In_4665);
or U897 (N_897,In_3047,In_3490);
or U898 (N_898,In_3533,In_4700);
or U899 (N_899,In_2235,In_4950);
and U900 (N_900,In_767,In_705);
nor U901 (N_901,In_1040,In_965);
or U902 (N_902,In_742,In_547);
or U903 (N_903,In_1852,In_2640);
and U904 (N_904,In_293,In_2676);
xor U905 (N_905,In_779,In_3817);
and U906 (N_906,In_1429,In_3484);
nor U907 (N_907,In_3101,In_2405);
nor U908 (N_908,In_595,In_3348);
nand U909 (N_909,In_3342,In_4581);
nand U910 (N_910,In_391,In_1173);
xor U911 (N_911,In_986,In_2489);
or U912 (N_912,In_2880,In_1983);
nor U913 (N_913,In_3073,In_460);
xnor U914 (N_914,In_2227,In_4210);
or U915 (N_915,In_3353,In_945);
and U916 (N_916,In_1805,In_1095);
nand U917 (N_917,In_4940,In_1690);
nand U918 (N_918,In_3576,In_1467);
or U919 (N_919,In_4087,In_2355);
nand U920 (N_920,In_1381,In_3556);
xor U921 (N_921,In_2652,In_3084);
or U922 (N_922,In_4784,In_4229);
nor U923 (N_923,In_1170,In_631);
and U924 (N_924,In_3568,In_3912);
or U925 (N_925,In_430,In_4441);
or U926 (N_926,In_3730,In_4633);
nand U927 (N_927,In_2944,In_1270);
xor U928 (N_928,In_3985,In_475);
xor U929 (N_929,In_3637,In_1036);
or U930 (N_930,In_3960,In_1405);
nand U931 (N_931,In_558,In_4497);
xor U932 (N_932,In_975,In_2763);
nor U933 (N_933,In_424,In_4490);
and U934 (N_934,In_1950,In_1424);
nand U935 (N_935,In_4438,In_3827);
nor U936 (N_936,In_2149,In_3741);
nand U937 (N_937,In_2700,In_89);
or U938 (N_938,In_62,In_1221);
or U939 (N_939,In_1656,In_2883);
or U940 (N_940,In_4944,In_1131);
or U941 (N_941,In_4680,In_1171);
nor U942 (N_942,In_1122,In_245);
nand U943 (N_943,In_4094,In_4635);
xor U944 (N_944,In_4339,In_4583);
nor U945 (N_945,In_4946,In_2756);
xor U946 (N_946,In_1354,In_2553);
or U947 (N_947,In_3371,In_3382);
xor U948 (N_948,In_516,In_3750);
nor U949 (N_949,In_4078,In_3549);
or U950 (N_950,In_720,In_3583);
or U951 (N_951,In_3351,In_199);
nor U952 (N_952,In_2964,In_1292);
and U953 (N_953,In_1344,In_4342);
and U954 (N_954,In_2226,In_4814);
nor U955 (N_955,In_4707,In_4704);
nand U956 (N_956,In_1925,In_3336);
or U957 (N_957,In_4743,In_212);
xnor U958 (N_958,In_3062,In_1053);
nand U959 (N_959,In_3376,In_412);
nor U960 (N_960,In_4598,In_704);
and U961 (N_961,In_2708,In_3904);
nor U962 (N_962,In_1955,In_3662);
nor U963 (N_963,In_1732,In_1909);
nor U964 (N_964,In_3307,In_1201);
and U965 (N_965,In_1198,In_2248);
nor U966 (N_966,In_1088,In_1113);
nor U967 (N_967,In_1205,In_4476);
or U968 (N_968,In_1665,In_4525);
and U969 (N_969,In_1795,In_488);
xor U970 (N_970,In_1346,In_4391);
nor U971 (N_971,In_4126,In_998);
nand U972 (N_972,In_3282,In_3152);
nor U973 (N_973,In_4616,In_2156);
or U974 (N_974,In_2629,In_1913);
or U975 (N_975,In_4589,In_768);
xor U976 (N_976,In_879,In_4216);
xor U977 (N_977,In_954,In_3665);
or U978 (N_978,In_3651,In_4816);
nand U979 (N_979,In_3179,In_59);
nand U980 (N_980,In_4491,In_2638);
xor U981 (N_981,In_4880,In_2440);
or U982 (N_982,In_863,In_3888);
xnor U983 (N_983,In_144,In_4577);
nor U984 (N_984,In_3066,In_4244);
and U985 (N_985,In_2532,In_3106);
nand U986 (N_986,In_673,In_1300);
or U987 (N_987,In_2956,In_3602);
and U988 (N_988,In_573,In_2780);
or U989 (N_989,In_1051,In_1432);
xor U990 (N_990,In_1807,In_3499);
or U991 (N_991,In_1102,In_2379);
and U992 (N_992,In_3438,In_4107);
nand U993 (N_993,In_2785,In_4960);
nor U994 (N_994,In_2834,In_524);
nand U995 (N_995,In_715,In_2088);
nor U996 (N_996,In_1,In_816);
xor U997 (N_997,In_207,In_2493);
and U998 (N_998,In_4254,In_3773);
nand U999 (N_999,In_1929,In_77);
nor U1000 (N_1000,In_3759,In_3495);
nand U1001 (N_1001,In_581,In_4566);
and U1002 (N_1002,In_1252,In_2519);
nand U1003 (N_1003,In_726,In_761);
or U1004 (N_1004,In_2545,In_3200);
nor U1005 (N_1005,In_1096,In_4171);
nor U1006 (N_1006,In_4695,N_766);
or U1007 (N_1007,In_3762,In_1372);
xor U1008 (N_1008,In_2272,In_4466);
or U1009 (N_1009,In_4580,In_3454);
and U1010 (N_1010,In_1488,In_4613);
or U1011 (N_1011,N_225,In_2146);
xor U1012 (N_1012,In_2076,N_973);
or U1013 (N_1013,N_538,N_364);
or U1014 (N_1014,In_2153,In_2624);
xnor U1015 (N_1015,In_1522,In_4962);
and U1016 (N_1016,In_4526,N_997);
xnor U1017 (N_1017,N_882,In_518);
nor U1018 (N_1018,In_533,N_305);
nor U1019 (N_1019,N_159,In_1598);
and U1020 (N_1020,N_927,In_2444);
nor U1021 (N_1021,In_2873,N_943);
nand U1022 (N_1022,N_961,In_0);
nor U1023 (N_1023,N_265,In_3184);
nor U1024 (N_1024,N_842,In_242);
nor U1025 (N_1025,In_2840,N_565);
xnor U1026 (N_1026,N_475,In_3954);
and U1027 (N_1027,In_993,In_733);
xor U1028 (N_1028,In_3879,In_185);
or U1029 (N_1029,N_680,In_1274);
nand U1030 (N_1030,In_4425,In_3221);
nand U1031 (N_1031,In_1693,In_2426);
xor U1032 (N_1032,N_107,In_3058);
or U1033 (N_1033,In_1957,In_2645);
and U1034 (N_1034,In_247,N_430);
nand U1035 (N_1035,In_3635,N_970);
or U1036 (N_1036,In_3370,In_2450);
nand U1037 (N_1037,In_2731,In_1835);
nor U1038 (N_1038,In_1454,In_2264);
or U1039 (N_1039,In_3632,N_467);
and U1040 (N_1040,In_4668,In_3613);
xnor U1041 (N_1041,In_2576,In_2794);
nor U1042 (N_1042,In_2347,N_223);
and U1043 (N_1043,In_2077,N_40);
nor U1044 (N_1044,In_3485,In_3715);
or U1045 (N_1045,In_2842,In_3857);
nor U1046 (N_1046,N_748,N_283);
or U1047 (N_1047,In_3333,In_4136);
xnor U1048 (N_1048,In_107,In_3781);
nor U1049 (N_1049,In_943,N_414);
nor U1050 (N_1050,In_2751,In_375);
xnor U1051 (N_1051,N_70,In_4775);
nor U1052 (N_1052,N_67,In_1412);
and U1053 (N_1053,In_4874,N_620);
nor U1054 (N_1054,N_907,N_647);
or U1055 (N_1055,In_355,N_511);
or U1056 (N_1056,N_694,In_1714);
nor U1057 (N_1057,In_559,N_755);
and U1058 (N_1058,N_412,In_3328);
or U1059 (N_1059,In_1707,N_626);
xor U1060 (N_1060,In_3795,In_1725);
and U1061 (N_1061,In_2950,In_4684);
nor U1062 (N_1062,N_561,In_4288);
xnor U1063 (N_1063,In_1369,In_4892);
xor U1064 (N_1064,In_1419,In_3278);
nand U1065 (N_1065,N_247,In_3310);
and U1066 (N_1066,In_3192,In_1351);
nor U1067 (N_1067,In_4931,In_1183);
and U1068 (N_1068,In_2656,In_4065);
nand U1069 (N_1069,In_3956,In_2726);
nand U1070 (N_1070,N_632,N_378);
xnor U1071 (N_1071,In_4912,In_4539);
nor U1072 (N_1072,N_457,In_86);
nor U1073 (N_1073,In_3705,In_4556);
and U1074 (N_1074,In_4007,In_254);
or U1075 (N_1075,N_901,In_3974);
and U1076 (N_1076,In_3516,In_610);
or U1077 (N_1077,In_1027,In_4446);
xnor U1078 (N_1078,N_258,N_570);
nand U1079 (N_1079,In_1337,In_2710);
nand U1080 (N_1080,N_42,In_3140);
xor U1081 (N_1081,N_298,In_1644);
nand U1082 (N_1082,In_2138,N_497);
and U1083 (N_1083,In_2464,In_3367);
or U1084 (N_1084,In_3968,In_2282);
xnor U1085 (N_1085,In_1607,In_4913);
and U1086 (N_1086,In_3399,In_2682);
or U1087 (N_1087,In_2853,In_1767);
nand U1088 (N_1088,N_77,In_1937);
nand U1089 (N_1089,N_541,N_614);
xnor U1090 (N_1090,In_4546,N_873);
or U1091 (N_1091,In_3251,In_2211);
or U1092 (N_1092,N_783,N_628);
xnor U1093 (N_1093,In_880,In_3756);
nor U1094 (N_1094,N_373,In_3626);
xnor U1095 (N_1095,In_1375,N_665);
nor U1096 (N_1096,In_1682,In_710);
nor U1097 (N_1097,N_267,In_2116);
and U1098 (N_1098,In_4600,In_2533);
nand U1099 (N_1099,In_173,N_161);
or U1100 (N_1100,In_2767,In_2857);
and U1101 (N_1101,In_728,In_4492);
or U1102 (N_1102,In_4791,In_3317);
nand U1103 (N_1103,N_420,In_2655);
nand U1104 (N_1104,In_50,N_636);
nor U1105 (N_1105,In_665,In_3392);
and U1106 (N_1106,In_4201,In_1989);
and U1107 (N_1107,N_205,In_2909);
nand U1108 (N_1108,In_2017,In_4686);
xnor U1109 (N_1109,In_214,In_2558);
nand U1110 (N_1110,N_635,In_628);
nand U1111 (N_1111,In_2725,In_1743);
xnor U1112 (N_1112,In_4306,N_958);
or U1113 (N_1113,N_94,In_1503);
nand U1114 (N_1114,In_3561,In_4366);
or U1115 (N_1115,In_1215,In_3461);
nand U1116 (N_1116,N_175,In_241);
xnor U1117 (N_1117,In_2187,In_4141);
and U1118 (N_1118,In_4437,In_2310);
nor U1119 (N_1119,In_3552,In_4079);
nor U1120 (N_1120,N_323,N_607);
nor U1121 (N_1121,N_763,In_4134);
and U1122 (N_1122,In_3334,In_4398);
or U1123 (N_1123,In_2139,In_4622);
and U1124 (N_1124,In_2899,In_2268);
nand U1125 (N_1125,In_3385,In_1910);
nor U1126 (N_1126,In_2686,In_2423);
and U1127 (N_1127,N_508,N_466);
or U1128 (N_1128,In_2683,In_2389);
nand U1129 (N_1129,In_1434,In_1766);
nor U1130 (N_1130,N_336,In_2783);
nand U1131 (N_1131,In_1518,N_764);
or U1132 (N_1132,N_252,In_3257);
and U1133 (N_1133,In_3670,N_193);
or U1134 (N_1134,In_4628,In_415);
or U1135 (N_1135,N_594,In_3748);
nor U1136 (N_1136,In_2772,In_781);
xor U1137 (N_1137,In_2813,In_652);
nor U1138 (N_1138,In_1323,In_80);
or U1139 (N_1139,In_762,In_1244);
nand U1140 (N_1140,N_521,In_4014);
nor U1141 (N_1141,N_355,In_1032);
and U1142 (N_1142,In_2920,N_633);
xor U1143 (N_1143,In_310,N_80);
nand U1144 (N_1144,In_530,N_254);
nand U1145 (N_1145,In_3913,N_933);
nand U1146 (N_1146,In_3706,In_1762);
nand U1147 (N_1147,In_1273,In_4175);
nor U1148 (N_1148,N_921,In_4340);
or U1149 (N_1149,In_2949,In_1825);
and U1150 (N_1150,N_965,N_512);
xnor U1151 (N_1151,In_4233,In_4972);
or U1152 (N_1152,N_658,N_84);
nor U1153 (N_1153,In_627,In_3858);
and U1154 (N_1154,In_1571,N_232);
nor U1155 (N_1155,In_2012,In_1878);
and U1156 (N_1156,In_4682,In_4499);
xnor U1157 (N_1157,In_3335,In_1379);
nor U1158 (N_1158,In_614,In_2424);
nand U1159 (N_1159,In_1207,In_253);
xor U1160 (N_1160,In_2531,In_4049);
or U1161 (N_1161,In_3369,In_4834);
xor U1162 (N_1162,N_64,In_192);
nor U1163 (N_1163,N_772,In_3015);
or U1164 (N_1164,In_1407,In_2445);
nand U1165 (N_1165,In_2632,In_4445);
nor U1166 (N_1166,In_856,N_855);
and U1167 (N_1167,In_674,N_509);
or U1168 (N_1168,In_4222,In_2335);
and U1169 (N_1169,In_1277,In_1973);
nand U1170 (N_1170,In_2037,In_405);
or U1171 (N_1171,In_4938,In_2435);
nand U1172 (N_1172,In_1498,In_1868);
nor U1173 (N_1173,In_168,In_4752);
xnor U1174 (N_1174,N_822,N_945);
nor U1175 (N_1175,N_662,N_912);
xnor U1176 (N_1176,In_546,In_2266);
and U1177 (N_1177,N_656,In_3921);
and U1178 (N_1178,In_1697,In_4921);
nand U1179 (N_1179,In_1601,In_1942);
nor U1180 (N_1180,In_1015,In_3226);
xnor U1181 (N_1181,In_4650,N_868);
or U1182 (N_1182,In_3531,N_833);
xnor U1183 (N_1183,In_1793,N_953);
or U1184 (N_1184,In_1844,In_1348);
and U1185 (N_1185,N_66,In_4226);
xnor U1186 (N_1186,In_189,In_2824);
nor U1187 (N_1187,N_435,In_4247);
and U1188 (N_1188,In_1773,In_3600);
nor U1189 (N_1189,In_150,In_502);
nand U1190 (N_1190,N_580,In_740);
nor U1191 (N_1191,In_3086,N_82);
xnor U1192 (N_1192,In_743,In_622);
nor U1193 (N_1193,In_1806,In_3844);
or U1194 (N_1194,In_4097,In_98);
nor U1195 (N_1195,In_2127,In_2446);
or U1196 (N_1196,N_381,In_4249);
nand U1197 (N_1197,In_2013,In_2902);
or U1198 (N_1198,N_645,In_3398);
and U1199 (N_1199,In_555,In_215);
or U1200 (N_1200,In_1557,N_61);
nand U1201 (N_1201,In_4032,In_3870);
and U1202 (N_1202,In_3601,In_1919);
nand U1203 (N_1203,N_208,In_1402);
or U1204 (N_1204,In_4389,In_3467);
nand U1205 (N_1205,In_2203,In_2209);
nand U1206 (N_1206,In_2649,In_1206);
or U1207 (N_1207,In_213,In_4611);
nand U1208 (N_1208,In_2524,In_1209);
nor U1209 (N_1209,In_2033,N_870);
xor U1210 (N_1210,In_3915,In_2551);
xnor U1211 (N_1211,N_393,In_3021);
xnor U1212 (N_1212,N_885,In_3899);
or U1213 (N_1213,N_331,In_4038);
xor U1214 (N_1214,N_689,N_666);
xnor U1215 (N_1215,N_309,In_3986);
xor U1216 (N_1216,In_3957,In_1098);
nand U1217 (N_1217,In_3000,In_105);
nand U1218 (N_1218,N_785,In_4242);
or U1219 (N_1219,In_4642,In_597);
or U1220 (N_1220,N_100,In_4745);
nor U1221 (N_1221,In_2721,In_2550);
nand U1222 (N_1222,In_4075,In_1741);
or U1223 (N_1223,In_4403,In_4301);
or U1224 (N_1224,In_3826,In_1329);
and U1225 (N_1225,N_423,In_1643);
xnor U1226 (N_1226,In_2091,In_2007);
and U1227 (N_1227,N_667,In_553);
and U1228 (N_1228,In_138,In_1228);
nor U1229 (N_1229,N_552,In_1760);
and U1230 (N_1230,In_2178,N_306);
and U1231 (N_1231,N_856,In_3455);
xor U1232 (N_1232,In_4110,In_4888);
nor U1233 (N_1233,In_4540,In_3188);
nor U1234 (N_1234,N_173,N_354);
nand U1235 (N_1235,In_2732,In_4579);
nand U1236 (N_1236,In_1339,In_3605);
xnor U1237 (N_1237,In_2311,In_1101);
nand U1238 (N_1238,N_967,N_276);
or U1239 (N_1239,In_3196,In_12);
xor U1240 (N_1240,In_4651,In_1972);
nand U1241 (N_1241,N_403,In_1408);
nand U1242 (N_1242,In_702,In_3707);
nand U1243 (N_1243,In_910,N_101);
xor U1244 (N_1244,In_314,In_3406);
xor U1245 (N_1245,In_579,In_1978);
nor U1246 (N_1246,In_416,N_453);
and U1247 (N_1247,In_2261,In_4010);
xnor U1248 (N_1248,N_455,In_3638);
xnor U1249 (N_1249,N_180,In_4267);
nor U1250 (N_1250,In_3087,N_5);
xnor U1251 (N_1251,In_2373,In_4328);
and U1252 (N_1252,In_164,N_153);
and U1253 (N_1253,In_324,N_793);
or U1254 (N_1254,In_4341,In_2729);
or U1255 (N_1255,In_1352,In_3245);
and U1256 (N_1256,In_3832,N_824);
and U1257 (N_1257,In_308,In_1087);
nor U1258 (N_1258,N_639,In_3005);
nand U1259 (N_1259,N_296,In_4872);
nor U1260 (N_1260,In_4365,In_1414);
nand U1261 (N_1261,In_2038,N_81);
or U1262 (N_1262,N_391,N_473);
xnor U1263 (N_1263,In_3900,N_281);
nor U1264 (N_1264,In_2612,In_1242);
and U1265 (N_1265,In_3623,In_2748);
xor U1266 (N_1266,In_3951,In_2521);
and U1267 (N_1267,In_514,In_1008);
or U1268 (N_1268,N_606,N_974);
xor U1269 (N_1269,In_1772,In_1867);
nand U1270 (N_1270,In_2611,In_3714);
nor U1271 (N_1271,In_1977,In_3195);
or U1272 (N_1272,In_521,In_4954);
nand U1273 (N_1273,N_21,In_4925);
nand U1274 (N_1274,N_390,In_2328);
nor U1275 (N_1275,In_4048,In_2830);
nand U1276 (N_1276,In_824,In_353);
nand U1277 (N_1277,In_442,In_179);
nor U1278 (N_1278,N_471,In_2279);
and U1279 (N_1279,N_179,N_280);
nand U1280 (N_1280,In_3692,In_1525);
and U1281 (N_1281,N_458,In_3381);
or U1282 (N_1282,In_3572,In_2453);
nand U1283 (N_1283,In_4648,In_2904);
or U1284 (N_1284,In_1435,In_354);
and U1285 (N_1285,In_1560,In_725);
nor U1286 (N_1286,N_279,In_3862);
xor U1287 (N_1287,N_827,N_367);
xor U1288 (N_1288,In_2032,In_1931);
or U1289 (N_1289,N_648,In_4948);
xor U1290 (N_1290,In_1523,N_798);
or U1291 (N_1291,N_820,In_1271);
nor U1292 (N_1292,In_1178,In_2548);
nor U1293 (N_1293,In_4096,In_1777);
nor U1294 (N_1294,In_4116,In_1536);
and U1295 (N_1295,In_271,In_2246);
or U1296 (N_1296,N_91,In_2607);
or U1297 (N_1297,N_747,In_4033);
nor U1298 (N_1298,In_3596,In_1530);
or U1299 (N_1299,In_4017,N_73);
and U1300 (N_1300,In_1468,In_2688);
xnor U1301 (N_1301,In_4811,In_2243);
or U1302 (N_1302,In_2862,In_4163);
nor U1303 (N_1303,In_2833,N_337);
or U1304 (N_1304,In_4311,In_2900);
or U1305 (N_1305,N_522,In_889);
nor U1306 (N_1306,N_922,In_389);
nor U1307 (N_1307,In_2642,In_2170);
nand U1308 (N_1308,In_2747,In_2046);
xnor U1309 (N_1309,In_4935,In_3603);
or U1310 (N_1310,In_1443,In_4939);
nand U1311 (N_1311,In_4870,In_3976);
xor U1312 (N_1312,N_424,In_802);
xnor U1313 (N_1313,In_1166,N_568);
and U1314 (N_1314,In_4855,In_838);
xnor U1315 (N_1315,N_637,In_2095);
or U1316 (N_1316,In_450,In_4266);
xnor U1317 (N_1317,N_794,In_469);
and U1318 (N_1318,N_698,In_2617);
xor U1319 (N_1319,N_745,N_31);
xor U1320 (N_1320,In_3244,In_4185);
nand U1321 (N_1321,In_1358,In_1768);
nor U1322 (N_1322,N_796,In_4383);
xnor U1323 (N_1323,In_3033,In_4504);
nor U1324 (N_1324,N_110,N_760);
and U1325 (N_1325,In_4252,In_3147);
or U1326 (N_1326,In_411,In_4706);
or U1327 (N_1327,N_869,In_3650);
nor U1328 (N_1328,N_761,In_4588);
xor U1329 (N_1329,In_3277,In_4429);
and U1330 (N_1330,N_41,In_3405);
xor U1331 (N_1331,In_3038,In_3219);
or U1332 (N_1332,In_1752,In_2390);
nor U1333 (N_1333,In_3776,In_2784);
or U1334 (N_1334,In_2812,N_11);
and U1335 (N_1335,In_1426,N_872);
and U1336 (N_1336,In_2062,N_671);
nand U1337 (N_1337,N_87,In_4818);
nand U1338 (N_1338,In_2284,In_4);
or U1339 (N_1339,In_3048,N_562);
and U1340 (N_1340,In_2502,In_1715);
xor U1341 (N_1341,In_3992,N_203);
xnor U1342 (N_1342,In_899,In_2359);
or U1343 (N_1343,In_1296,In_3352);
and U1344 (N_1344,In_695,N_460);
and U1345 (N_1345,In_4871,In_3443);
nand U1346 (N_1346,N_454,N_691);
or U1347 (N_1347,In_4460,N_95);
nor U1348 (N_1348,In_190,In_2356);
xnor U1349 (N_1349,In_2936,N_998);
or U1350 (N_1350,In_2018,In_3142);
xnor U1351 (N_1351,In_4505,In_4734);
nand U1352 (N_1352,In_3309,In_3347);
nor U1353 (N_1353,In_3717,N_384);
xor U1354 (N_1354,In_3522,N_44);
and U1355 (N_1355,In_2181,In_3562);
and U1356 (N_1356,In_1308,N_705);
and U1357 (N_1357,In_4323,In_1709);
and U1358 (N_1358,In_1463,N_732);
nand U1359 (N_1359,In_2483,In_480);
nand U1360 (N_1360,In_987,In_341);
xnor U1361 (N_1361,N_476,In_2529);
and U1362 (N_1362,N_625,In_336);
or U1363 (N_1363,In_4967,N_776);
xnor U1364 (N_1364,In_932,In_4351);
and U1365 (N_1365,In_1817,In_2433);
and U1366 (N_1366,In_2049,N_60);
and U1367 (N_1367,N_621,In_443);
xnor U1368 (N_1368,In_3927,In_1326);
nor U1369 (N_1369,In_4661,N_816);
or U1370 (N_1370,In_2896,In_4767);
or U1371 (N_1371,N_896,In_1427);
and U1372 (N_1372,In_4819,In_2371);
nand U1373 (N_1373,In_4655,In_3373);
or U1374 (N_1374,N_165,In_2885);
nand U1375 (N_1375,In_198,In_2183);
xor U1376 (N_1376,In_843,In_1796);
or U1377 (N_1377,In_1357,N_241);
nand U1378 (N_1378,N_934,In_3354);
nor U1379 (N_1379,In_2128,In_616);
nand U1380 (N_1380,In_487,In_440);
or U1381 (N_1381,In_1915,In_4138);
or U1382 (N_1382,In_3973,In_122);
xnor U1383 (N_1383,In_2943,In_1626);
nor U1384 (N_1384,In_1469,In_4335);
and U1385 (N_1385,In_16,In_4794);
and U1386 (N_1386,N_358,In_887);
and U1387 (N_1387,In_2999,In_1620);
and U1388 (N_1388,In_2030,N_494);
nor U1389 (N_1389,N_195,In_2388);
nand U1390 (N_1390,In_432,N_994);
and U1391 (N_1391,N_212,In_3509);
and U1392 (N_1392,In_1839,N_589);
nor U1393 (N_1393,In_1464,In_3113);
and U1394 (N_1394,In_2861,In_4293);
or U1395 (N_1395,In_1513,In_1481);
xor U1396 (N_1396,N_861,In_4663);
or U1397 (N_1397,In_2086,In_3834);
xnor U1398 (N_1398,In_4421,In_936);
and U1399 (N_1399,In_1471,N_24);
or U1400 (N_1400,In_3962,In_1834);
nor U1401 (N_1401,In_3161,In_2176);
nor U1402 (N_1402,In_3833,In_2528);
or U1403 (N_1403,In_4806,In_2970);
xnor U1404 (N_1404,In_741,In_4371);
xor U1405 (N_1405,In_3493,In_1037);
or U1406 (N_1406,In_3263,In_2713);
or U1407 (N_1407,In_911,In_221);
and U1408 (N_1408,In_4234,N_495);
nand U1409 (N_1409,In_942,In_1237);
nand U1410 (N_1410,In_1333,In_780);
and U1411 (N_1411,N_275,In_3053);
nand U1412 (N_1412,In_4166,In_392);
nand U1413 (N_1413,N_320,In_3515);
nand U1414 (N_1414,In_182,In_4156);
nand U1415 (N_1415,In_4829,N_389);
and U1416 (N_1416,In_4637,In_4528);
nand U1417 (N_1417,In_492,In_3933);
and U1418 (N_1418,In_3803,In_617);
xor U1419 (N_1419,N_259,N_398);
nor U1420 (N_1420,In_4793,In_904);
and U1421 (N_1421,In_2110,In_4158);
or U1422 (N_1422,In_587,In_1251);
nor U1423 (N_1423,In_3236,In_1751);
nand U1424 (N_1424,In_1569,N_916);
nand U1425 (N_1425,In_1637,In_1425);
xor U1426 (N_1426,In_2835,In_602);
nor U1427 (N_1427,In_3302,In_1815);
nand U1428 (N_1428,In_3840,In_4106);
nor U1429 (N_1429,In_3872,N_926);
and U1430 (N_1430,In_4533,In_1572);
xnor U1431 (N_1431,In_1165,In_1678);
xnor U1432 (N_1432,In_2573,In_2189);
nand U1433 (N_1433,In_2704,In_730);
xor U1434 (N_1434,In_2418,In_1846);
nand U1435 (N_1435,In_4418,N_735);
or U1436 (N_1436,In_2891,In_388);
and U1437 (N_1437,In_4772,In_3727);
xnor U1438 (N_1438,In_3290,In_1599);
nor U1439 (N_1439,N_349,In_612);
nor U1440 (N_1440,In_3625,In_1840);
nand U1441 (N_1441,In_2154,In_1500);
nand U1442 (N_1442,In_4406,In_4355);
nand U1443 (N_1443,In_4659,N_292);
nand U1444 (N_1444,N_395,In_657);
nand U1445 (N_1445,N_447,In_3034);
or U1446 (N_1446,In_7,In_1940);
xnor U1447 (N_1447,N_892,In_3173);
nand U1448 (N_1448,In_3096,In_4553);
nor U1449 (N_1449,In_3390,In_2778);
xor U1450 (N_1450,In_4427,In_3949);
or U1451 (N_1451,N_238,In_398);
and U1452 (N_1452,In_210,In_3944);
nand U1453 (N_1453,N_130,In_4432);
nor U1454 (N_1454,In_3002,In_4467);
nand U1455 (N_1455,In_3815,In_1000);
or U1456 (N_1456,In_3994,N_217);
nand U1457 (N_1457,In_1524,In_3932);
nand U1458 (N_1458,In_2945,In_1422);
nor U1459 (N_1459,N_142,In_1747);
nand U1460 (N_1460,N_68,In_2535);
nand U1461 (N_1461,In_2864,In_161);
nand U1462 (N_1462,In_377,In_484);
or U1463 (N_1463,In_1097,In_3931);
xor U1464 (N_1464,N_756,In_1845);
nor U1465 (N_1465,In_2045,N_624);
nand U1466 (N_1466,In_1899,N_871);
and U1467 (N_1467,N_197,N_209);
or U1468 (N_1468,In_3575,In_913);
nand U1469 (N_1469,N_960,In_3483);
nor U1470 (N_1470,In_302,In_4521);
xnor U1471 (N_1471,In_2341,In_3850);
and U1472 (N_1472,N_123,In_3543);
or U1473 (N_1473,In_1475,In_4723);
or U1474 (N_1474,In_337,N_55);
nand U1475 (N_1475,In_1628,In_4765);
and U1476 (N_1476,In_601,In_1930);
nand U1477 (N_1477,N_780,In_39);
or U1478 (N_1478,In_1675,In_4895);
nand U1479 (N_1479,In_1011,In_2685);
nor U1480 (N_1480,In_230,In_4309);
nor U1481 (N_1481,In_3380,In_2283);
xnor U1482 (N_1482,In_2504,N_525);
xor U1483 (N_1483,In_2868,N_314);
xnor U1484 (N_1484,In_3319,In_158);
or U1485 (N_1485,In_2250,In_3496);
nor U1486 (N_1486,N_573,In_2238);
xnor U1487 (N_1487,In_3017,In_2722);
nand U1488 (N_1488,In_333,N_169);
and U1489 (N_1489,In_2897,In_3272);
xnor U1490 (N_1490,In_2385,In_2993);
nor U1491 (N_1491,In_4375,In_3767);
or U1492 (N_1492,In_4795,In_764);
or U1493 (N_1493,In_873,N_446);
and U1494 (N_1494,In_4823,N_526);
or U1495 (N_1495,In_1261,N_596);
xor U1496 (N_1496,In_4215,In_4205);
xnor U1497 (N_1497,N_183,In_382);
nor U1498 (N_1498,In_3855,In_3867);
xor U1499 (N_1499,In_2460,In_1570);
xnor U1500 (N_1500,In_4796,In_3672);
or U1501 (N_1501,In_1826,In_2334);
nor U1502 (N_1502,N_300,In_2082);
nand U1503 (N_1503,In_3557,In_1687);
or U1504 (N_1504,In_1636,N_324);
nand U1505 (N_1505,N_754,In_4084);
or U1506 (N_1506,In_3154,In_3291);
xnor U1507 (N_1507,N_334,N_712);
and U1508 (N_1508,In_312,In_1801);
nand U1509 (N_1509,In_2185,In_1269);
xnor U1510 (N_1510,N_59,N_726);
nand U1511 (N_1511,In_3537,N_692);
or U1512 (N_1512,N_546,N_765);
nand U1513 (N_1513,In_4626,In_2789);
xnor U1514 (N_1514,In_172,In_2739);
or U1515 (N_1515,In_2072,In_4414);
nand U1516 (N_1516,In_3254,In_1870);
nor U1517 (N_1517,In_3044,N_649);
and U1518 (N_1518,In_2946,In_2349);
or U1519 (N_1519,In_1295,N_133);
nand U1520 (N_1520,N_514,N_968);
nor U1521 (N_1521,N_581,N_731);
xnor U1522 (N_1522,In_1719,In_3439);
and U1523 (N_1523,In_2274,N_651);
or U1524 (N_1524,N_661,In_4304);
or U1525 (N_1525,N_787,In_1440);
and U1526 (N_1526,In_1961,In_4866);
and U1527 (N_1527,N_147,In_4807);
nor U1528 (N_1528,In_2410,In_1860);
and U1529 (N_1529,In_3330,In_2837);
or U1530 (N_1530,In_451,In_2458);
xnor U1531 (N_1531,In_1288,In_135);
or U1532 (N_1532,N_22,In_4754);
and U1533 (N_1533,In_789,In_4890);
and U1534 (N_1534,N_919,N_499);
nand U1535 (N_1535,N_644,In_3527);
nand U1536 (N_1536,In_4317,In_3952);
nor U1537 (N_1537,N_425,In_2276);
nor U1538 (N_1538,In_1390,In_3344);
nor U1539 (N_1539,In_4908,In_2671);
xnor U1540 (N_1540,N_777,In_519);
nor U1541 (N_1541,In_3621,N_51);
or U1542 (N_1542,N_791,In_3098);
nor U1543 (N_1543,In_3040,In_4900);
or U1544 (N_1544,N_116,N_815);
and U1545 (N_1545,In_4777,In_4942);
xnor U1546 (N_1546,N_132,In_2042);
and U1547 (N_1547,In_1077,In_3758);
and U1548 (N_1548,N_716,N_52);
nor U1549 (N_1549,In_3503,In_3449);
xor U1550 (N_1550,In_3924,In_463);
nor U1551 (N_1551,In_3989,In_2917);
xnor U1552 (N_1552,In_282,In_1856);
xnor U1553 (N_1553,In_3688,In_441);
nand U1554 (N_1554,In_4845,In_4011);
xor U1555 (N_1555,In_229,N_591);
nand U1556 (N_1556,In_1060,In_1506);
xnor U1557 (N_1557,N_981,In_3468);
nor U1558 (N_1558,In_970,In_2597);
and U1559 (N_1559,N_13,In_4856);
or U1560 (N_1560,N_400,In_1286);
xor U1561 (N_1561,N_903,In_874);
nor U1562 (N_1562,In_4392,In_493);
and U1563 (N_1563,In_2588,N_333);
and U1564 (N_1564,In_2008,In_3092);
nor U1565 (N_1565,In_223,In_4867);
or U1566 (N_1566,In_3765,In_3480);
nor U1567 (N_1567,N_164,In_2087);
xnor U1568 (N_1568,In_3838,In_3938);
xnor U1569 (N_1569,N_951,In_1988);
nand U1570 (N_1570,In_3629,In_512);
or U1571 (N_1571,In_3433,In_1117);
nor U1572 (N_1572,In_650,In_1722);
or U1573 (N_1573,In_3517,In_4384);
nor U1574 (N_1574,In_4947,In_4721);
xor U1575 (N_1575,In_4277,In_1293);
xnor U1576 (N_1576,In_2057,In_2605);
xor U1577 (N_1577,In_4227,N_598);
nand U1578 (N_1578,In_2074,In_2670);
or U1579 (N_1579,In_4641,N_930);
and U1580 (N_1580,In_3252,In_4713);
nor U1581 (N_1581,In_1618,In_4117);
and U1582 (N_1582,In_1258,In_300);
or U1583 (N_1583,In_2428,In_3325);
or U1584 (N_1584,N_187,In_4043);
or U1585 (N_1585,In_3345,In_4924);
nor U1586 (N_1586,In_2175,In_4766);
and U1587 (N_1587,In_886,In_4759);
nand U1588 (N_1588,In_4296,N_769);
nand U1589 (N_1589,In_2448,N_23);
nand U1590 (N_1590,In_1017,In_4091);
or U1591 (N_1591,In_1691,In_3279);
nor U1592 (N_1592,In_101,In_1023);
or U1593 (N_1593,N_449,N_937);
nor U1594 (N_1594,In_1146,In_3693);
and U1595 (N_1595,In_363,N_623);
xor U1596 (N_1596,In_3769,In_2362);
xnor U1597 (N_1597,In_3820,N_329);
and U1598 (N_1598,N_444,In_2323);
xor U1599 (N_1599,N_363,In_2911);
nand U1600 (N_1600,In_1263,In_2757);
and U1601 (N_1601,In_3041,In_3167);
xnor U1602 (N_1602,N_143,In_343);
and U1603 (N_1603,N_118,In_1509);
xor U1604 (N_1604,In_3177,In_4025);
xor U1605 (N_1605,In_3972,In_3511);
and U1606 (N_1606,In_1361,In_1811);
and U1607 (N_1607,In_961,In_4397);
xor U1608 (N_1608,In_3873,In_1115);
nor U1609 (N_1609,In_2169,N_234);
nand U1610 (N_1610,In_3871,In_2765);
nor U1611 (N_1611,In_4673,In_2844);
nor U1612 (N_1612,In_4448,N_206);
or U1613 (N_1613,In_4295,In_2031);
nand U1614 (N_1614,In_734,In_2674);
and U1615 (N_1615,N_604,In_1074);
or U1616 (N_1616,In_2184,N_590);
and U1617 (N_1617,In_1574,In_1398);
nand U1618 (N_1618,In_3386,N_429);
xor U1619 (N_1619,In_2641,In_976);
xnor U1620 (N_1620,In_794,N_688);
nor U1621 (N_1621,N_672,In_1646);
and U1622 (N_1622,In_3578,In_4532);
and U1623 (N_1623,In_491,In_1437);
nor U1624 (N_1624,In_1623,In_1651);
nand U1625 (N_1625,In_753,N_233);
xnor U1626 (N_1626,In_3766,In_4270);
nor U1627 (N_1627,In_1740,N_778);
and U1628 (N_1628,N_194,In_2668);
nand U1629 (N_1629,In_3569,N_935);
or U1630 (N_1630,N_622,In_2995);
or U1631 (N_1631,In_1585,N_141);
nand U1632 (N_1632,N_200,N_437);
xnor U1633 (N_1633,In_1185,N_584);
xor U1634 (N_1634,In_2580,In_3024);
or U1635 (N_1635,In_2381,In_1121);
nor U1636 (N_1636,In_2475,In_2637);
nor U1637 (N_1637,In_3920,In_6);
or U1638 (N_1638,In_3647,In_2823);
and U1639 (N_1639,In_2236,In_4652);
or U1640 (N_1640,In_2005,In_698);
nor U1641 (N_1641,N_345,In_2499);
and U1642 (N_1642,N_270,In_769);
xor U1643 (N_1643,In_3801,In_2047);
nand U1644 (N_1644,In_3743,In_2894);
xor U1645 (N_1645,N_723,In_2193);
or U1646 (N_1646,N_464,N_889);
nor U1647 (N_1647,In_4735,N_995);
or U1648 (N_1648,In_3875,In_1911);
nand U1649 (N_1649,N_557,In_4380);
xor U1650 (N_1650,In_4159,N_852);
nand U1651 (N_1651,N_841,In_3811);
nand U1652 (N_1652,In_151,In_4592);
nand U1653 (N_1653,N_248,In_811);
nor U1654 (N_1654,In_81,N_122);
and U1655 (N_1655,In_4558,In_981);
and U1656 (N_1656,In_4083,In_783);
or U1657 (N_1657,N_668,In_414);
and U1658 (N_1658,In_4692,In_1612);
nand U1659 (N_1659,N_659,N_831);
nor U1660 (N_1660,N_450,In_1584);
or U1661 (N_1661,In_626,In_882);
and U1662 (N_1662,In_2988,In_1368);
nand U1663 (N_1663,In_1833,N_263);
xor U1664 (N_1664,In_3965,N_971);
or U1665 (N_1665,In_4072,In_4677);
xnor U1666 (N_1666,In_4020,In_2317);
nand U1667 (N_1667,N_739,N_230);
nand U1668 (N_1668,In_2326,In_505);
xnor U1669 (N_1669,In_155,In_1458);
and U1670 (N_1670,N_753,In_1191);
or U1671 (N_1671,In_4957,In_2614);
xor U1672 (N_1672,In_883,N_178);
and U1673 (N_1673,In_191,N_702);
nand U1674 (N_1674,N_650,In_2113);
or U1675 (N_1675,In_478,In_2958);
nand U1676 (N_1676,In_2804,In_897);
nor U1677 (N_1677,N_313,N_743);
xor U1678 (N_1678,In_4666,N_1);
xnor U1679 (N_1679,In_2635,In_2938);
or U1680 (N_1680,N_832,In_4851);
or U1681 (N_1681,N_838,In_4202);
xnor U1682 (N_1682,N_191,In_1428);
xnor U1683 (N_1683,In_1363,In_4519);
and U1684 (N_1684,N_980,In_106);
or U1685 (N_1685,N_840,In_926);
xor U1686 (N_1686,N_749,In_583);
nand U1687 (N_1687,In_4805,In_604);
nand U1688 (N_1688,In_2511,In_3805);
and U1689 (N_1689,N_876,In_2291);
or U1690 (N_1690,N_914,In_2461);
or U1691 (N_1691,In_2922,In_264);
nor U1692 (N_1692,N_351,In_1632);
and U1693 (N_1693,In_500,N_172);
and U1694 (N_1694,In_103,In_143);
and U1695 (N_1695,In_63,In_4307);
nor U1696 (N_1696,In_2473,In_1044);
xnor U1697 (N_1697,In_1857,In_4152);
or U1698 (N_1698,In_571,In_4113);
or U1699 (N_1699,In_233,In_3914);
nand U1700 (N_1700,N_278,In_771);
nor U1701 (N_1701,N_261,N_158);
nor U1702 (N_1702,N_675,In_756);
xor U1703 (N_1703,In_1022,In_4246);
nand U1704 (N_1704,N_992,In_4346);
xnor U1705 (N_1705,N_369,In_3043);
and U1706 (N_1706,N_879,N_126);
or U1707 (N_1707,In_3091,In_1886);
and U1708 (N_1708,In_1734,In_137);
nor U1709 (N_1709,N_216,N_696);
nor U1710 (N_1710,In_992,In_1181);
and U1711 (N_1711,In_3942,In_1328);
nand U1712 (N_1712,N_375,In_1898);
nor U1713 (N_1713,In_1264,N_88);
or U1714 (N_1714,N_988,N_664);
or U1715 (N_1715,In_4575,In_3487);
or U1716 (N_1716,In_803,In_4261);
and U1717 (N_1717,In_1306,N_888);
and U1718 (N_1718,N_847,N_806);
or U1719 (N_1719,In_2148,In_2214);
or U1720 (N_1720,In_3067,In_1441);
xnor U1721 (N_1721,In_738,In_2650);
and U1722 (N_1722,In_1517,In_4008);
and U1723 (N_1723,N_528,In_563);
and U1724 (N_1724,N_171,In_48);
xnor U1725 (N_1725,N_9,In_498);
or U1726 (N_1726,In_2697,In_1041);
nand U1727 (N_1727,In_2130,In_4130);
and U1728 (N_1728,In_497,In_1197);
xnor U1729 (N_1729,In_3045,In_3747);
nand U1730 (N_1730,N_326,In_3648);
nand U1731 (N_1731,N_775,In_2275);
or U1732 (N_1732,In_2626,In_4196);
nand U1733 (N_1733,In_4615,In_13);
nand U1734 (N_1734,In_4453,In_2101);
xor U1735 (N_1735,In_2145,In_385);
nor U1736 (N_1736,In_4932,N_823);
or U1737 (N_1737,In_765,In_1482);
or U1738 (N_1738,In_1250,In_114);
nand U1739 (N_1739,In_2581,In_3624);
nand U1740 (N_1740,N_185,In_1541);
or U1741 (N_1741,In_474,N_657);
nor U1742 (N_1742,In_2200,In_125);
nand U1743 (N_1743,N_759,In_3779);
nand U1744 (N_1744,In_231,In_2035);
or U1745 (N_1745,N_503,In_4449);
and U1746 (N_1746,In_3265,In_3898);
xor U1747 (N_1747,N_518,N_846);
nor U1748 (N_1748,In_4314,In_3909);
nand U1749 (N_1749,N_117,In_560);
nor U1750 (N_1750,In_4211,In_2430);
nand U1751 (N_1751,In_4004,In_4738);
nor U1752 (N_1752,In_3618,In_4568);
nand U1753 (N_1753,In_3666,N_114);
xnor U1754 (N_1754,In_2395,N_271);
nor U1755 (N_1755,In_32,N_501);
nand U1756 (N_1756,In_660,In_1531);
nand U1757 (N_1757,In_2260,In_1052);
nand U1758 (N_1758,N_660,In_3059);
nand U1759 (N_1759,N_372,In_858);
xnor U1760 (N_1760,In_3268,In_2090);
nor U1761 (N_1761,In_2615,In_335);
nand U1762 (N_1762,In_4169,In_58);
or U1763 (N_1763,In_52,In_2933);
and U1764 (N_1764,In_902,In_4188);
nand U1765 (N_1765,N_505,In_717);
nor U1766 (N_1766,In_2180,In_383);
nor U1767 (N_1767,In_787,N_894);
nand U1768 (N_1768,In_445,In_1248);
nand U1769 (N_1769,N_111,In_3893);
nor U1770 (N_1770,In_4177,N_703);
xor U1771 (N_1771,In_2407,In_4006);
nor U1772 (N_1772,In_2419,In_1108);
nand U1773 (N_1773,In_359,In_2888);
nor U1774 (N_1774,N_500,N_938);
nor U1775 (N_1775,N_468,In_2578);
xor U1776 (N_1776,In_2807,In_2384);
nor U1777 (N_1777,N_966,In_3722);
xnor U1778 (N_1778,N_39,N_729);
and U1779 (N_1779,In_599,In_1684);
and U1780 (N_1780,In_731,N_374);
and U1781 (N_1781,N_461,In_4570);
nor U1782 (N_1782,In_4614,In_3388);
or U1783 (N_1783,In_2570,In_1965);
xnor U1784 (N_1784,In_1132,In_3935);
nand U1785 (N_1785,N_383,In_1396);
or U1786 (N_1786,In_1225,In_1891);
or U1787 (N_1787,N_738,In_4120);
nand U1788 (N_1788,In_773,In_244);
and U1789 (N_1789,N_493,In_180);
xnor U1790 (N_1790,In_691,In_3093);
or U1791 (N_1791,N_583,In_2094);
xor U1792 (N_1792,In_1384,In_3237);
and U1793 (N_1793,In_4149,N_177);
xor U1794 (N_1794,In_1356,In_1549);
and U1795 (N_1795,N_139,In_4857);
and U1796 (N_1796,In_3056,In_2646);
xnor U1797 (N_1797,N_762,In_4401);
and U1798 (N_1798,N_15,In_3588);
or U1799 (N_1799,N_682,In_3825);
or U1800 (N_1800,In_4849,In_606);
nand U1801 (N_1801,N_697,N_0);
nor U1802 (N_1802,In_2278,In_2996);
and U1803 (N_1803,N_843,N_32);
nand U1804 (N_1804,In_862,N_428);
nor U1805 (N_1805,In_1661,N_182);
nor U1806 (N_1806,In_1365,In_3610);
nand U1807 (N_1807,In_1742,N_253);
and U1808 (N_1808,In_1176,In_3012);
xor U1809 (N_1809,In_204,In_3191);
and U1810 (N_1810,In_817,In_2241);
nand U1811 (N_1811,In_2210,In_3996);
and U1812 (N_1812,In_4899,In_1730);
or U1813 (N_1813,In_4821,In_1841);
xnor U1814 (N_1814,In_1304,In_799);
nor U1815 (N_1815,N_954,N_537);
xnor U1816 (N_1816,In_1798,In_1836);
or U1817 (N_1817,In_2132,In_472);
nor U1818 (N_1818,In_165,In_1161);
or U1819 (N_1819,In_4737,In_2447);
and U1820 (N_1820,N_316,N_956);
xor U1821 (N_1821,In_4178,In_1501);
nand U1822 (N_1822,In_929,In_4909);
or U1823 (N_1823,In_4640,N_472);
or U1824 (N_1824,In_2799,In_3643);
nor U1825 (N_1825,In_297,N_272);
and U1826 (N_1826,N_850,N_28);
or U1827 (N_1827,N_773,In_3115);
nor U1828 (N_1828,In_295,In_2491);
or U1829 (N_1829,In_3828,N_370);
or U1830 (N_1830,In_4232,In_2965);
nand U1831 (N_1831,N_531,In_1947);
and U1832 (N_1832,N_315,N_26);
nor U1833 (N_1833,In_1879,N_382);
and U1834 (N_1834,In_556,N_266);
and U1835 (N_1835,In_1816,In_2251);
or U1836 (N_1836,In_3716,In_2416);
or U1837 (N_1837,In_3829,In_4040);
or U1838 (N_1838,In_4124,In_2109);
xor U1839 (N_1839,In_2111,N_519);
and U1840 (N_1840,In_291,N_737);
xor U1841 (N_1841,In_3641,In_1699);
xor U1842 (N_1842,N_418,In_141);
and U1843 (N_1843,In_462,N_341);
xor U1844 (N_1844,In_2336,In_481);
and U1845 (N_1845,In_2513,In_620);
nand U1846 (N_1846,In_365,In_345);
xor U1847 (N_1847,In_3323,In_2383);
xnor U1848 (N_1848,N_506,In_3941);
xor U1849 (N_1849,In_3593,In_4433);
or U1850 (N_1850,In_4887,In_2654);
nand U1851 (N_1851,N_744,In_4711);
xnor U1852 (N_1852,In_4187,In_2267);
and U1853 (N_1853,In_593,In_2402);
and U1854 (N_1854,N_407,In_525);
nand U1855 (N_1855,In_2625,In_384);
and U1856 (N_1856,In_3136,N_239);
xor U1857 (N_1857,In_2117,In_321);
xor U1858 (N_1858,In_1391,In_93);
and U1859 (N_1859,In_2364,In_1949);
and U1860 (N_1860,In_1727,In_4672);
nor U1861 (N_1861,N_711,In_178);
xor U1862 (N_1862,In_2150,In_2119);
nand U1863 (N_1863,In_1907,In_4901);
or U1864 (N_1864,N_693,In_251);
or U1865 (N_1865,In_2648,In_648);
or U1866 (N_1866,In_515,In_3874);
nand U1867 (N_1867,In_2443,N_599);
xnor U1868 (N_1868,In_2484,In_1704);
nor U1869 (N_1869,N_963,N_710);
xor U1870 (N_1870,In_4396,In_4507);
nand U1871 (N_1871,In_1749,N_434);
xor U1872 (N_1872,In_2634,N_318);
nor U1873 (N_1873,In_1029,In_4503);
xor U1874 (N_1874,N_559,In_3551);
nand U1875 (N_1875,In_3235,N_213);
nand U1876 (N_1876,In_1138,In_662);
xnor U1877 (N_1877,N_610,N_484);
and U1878 (N_1878,In_4669,N_653);
nor U1879 (N_1879,In_3847,N_92);
or U1880 (N_1880,N_128,N_813);
and U1881 (N_1881,In_46,In_1128);
nor U1882 (N_1882,In_1119,In_754);
nor U1883 (N_1883,N_18,In_1654);
and U1884 (N_1884,N_811,In_2058);
xor U1885 (N_1885,In_1495,In_201);
xor U1886 (N_1886,In_1689,In_4370);
and U1887 (N_1887,In_4444,N_121);
nand U1888 (N_1888,In_4955,In_482);
xnor U1889 (N_1889,In_1380,In_3103);
nand U1890 (N_1890,In_4762,In_3457);
nor U1891 (N_1891,N_150,In_4057);
or U1892 (N_1892,In_1922,In_249);
xnor U1893 (N_1893,In_3476,N_535);
and U1894 (N_1894,In_4873,In_1615);
nand U1895 (N_1895,N_805,In_4678);
or U1896 (N_1896,In_3054,In_1031);
xor U1897 (N_1897,In_615,In_3460);
xnor U1898 (N_1898,In_347,In_3415);
nor U1899 (N_1899,In_1779,N_311);
nand U1900 (N_1900,In_3519,In_3241);
xor U1901 (N_1901,In_409,In_2295);
or U1902 (N_1902,N_957,In_3401);
nor U1903 (N_1903,In_318,In_3150);
nor U1904 (N_1904,In_755,N_58);
and U1905 (N_1905,In_1192,In_3886);
nand U1906 (N_1906,In_3166,In_4727);
or U1907 (N_1907,In_4993,In_4036);
xor U1908 (N_1908,In_1075,In_2369);
nor U1909 (N_1909,In_2771,In_417);
nand U1910 (N_1910,N_670,In_4353);
nor U1911 (N_1911,In_3725,N_890);
nand U1912 (N_1912,In_396,In_4714);
nor U1913 (N_1913,N_2,In_1666);
nand U1914 (N_1914,N_392,In_3233);
nand U1915 (N_1915,In_2761,N_332);
xnor U1916 (N_1916,In_870,In_3523);
and U1917 (N_1917,In_2237,In_120);
xnor U1918 (N_1918,In_1169,N_317);
nor U1919 (N_1919,In_2457,In_1677);
or U1920 (N_1920,In_327,In_1490);
and U1921 (N_1921,In_812,In_1669);
and U1922 (N_1922,In_2120,In_3642);
xor U1923 (N_1923,In_2265,In_2711);
and U1924 (N_1924,In_763,N_157);
or U1925 (N_1925,In_2010,In_3807);
nand U1926 (N_1926,In_4756,In_3271);
xor U1927 (N_1927,N_543,In_1150);
or U1928 (N_1928,In_646,In_2466);
or U1929 (N_1929,In_1663,N_199);
nor U1930 (N_1930,N_867,In_2164);
xnor U1931 (N_1931,In_3628,In_496);
or U1932 (N_1932,In_2322,In_1492);
and U1933 (N_1933,In_3383,In_1061);
xnor U1934 (N_1934,In_4755,In_4026);
nand U1935 (N_1935,In_3248,In_3213);
xor U1936 (N_1936,In_4123,In_1336);
or U1937 (N_1937,N_490,In_4151);
nor U1938 (N_1938,N_45,In_3555);
xor U1939 (N_1939,In_565,In_749);
nor U1940 (N_1940,In_3616,In_1794);
nor U1941 (N_1941,In_1968,N_608);
and U1942 (N_1942,N_897,N_560);
or U1943 (N_1943,In_1731,In_104);
xor U1944 (N_1944,In_979,N_478);
nor U1945 (N_1945,In_4868,In_3242);
xor U1946 (N_1946,In_4841,In_4344);
xor U1947 (N_1947,N_409,In_694);
xor U1948 (N_1948,In_3312,In_4905);
or U1949 (N_1949,N_12,In_1282);
xor U1950 (N_1950,In_3658,N_586);
and U1951 (N_1951,In_1568,In_837);
xor U1952 (N_1952,In_1485,In_3285);
nor U1953 (N_1953,N_880,In_1759);
xor U1954 (N_1954,In_376,In_2071);
nor U1955 (N_1955,N_145,In_724);
xor U1956 (N_1956,N_286,In_1600);
and U1957 (N_1957,In_4716,In_3203);
nand U1958 (N_1958,N_339,In_3216);
and U1959 (N_1959,N_96,In_4602);
nand U1960 (N_1960,In_116,In_2118);
xnor U1961 (N_1961,In_3895,In_3677);
or U1962 (N_1962,In_4241,In_4345);
or U1963 (N_1963,In_881,In_2289);
or U1964 (N_1964,In_4194,In_3458);
nand U1965 (N_1965,N_463,N_210);
xnor U1966 (N_1966,N_264,In_3856);
nand U1967 (N_1967,In_2775,In_4334);
and U1968 (N_1968,In_1200,In_4736);
or U1969 (N_1969,In_3839,In_2303);
nand U1970 (N_1970,N_854,In_963);
and U1971 (N_1971,In_4980,N_836);
nand U1972 (N_1972,N_38,N_618);
and U1973 (N_1973,In_2287,In_4826);
nor U1974 (N_1974,In_142,N_849);
and U1975 (N_1975,In_4590,In_4778);
xnor U1976 (N_1976,In_3736,In_186);
and U1977 (N_1977,In_4658,N_97);
and U1978 (N_1978,N_215,In_1659);
nand U1979 (N_1979,In_2695,In_2791);
and U1980 (N_1980,In_1080,In_3497);
and U1981 (N_1981,In_2836,In_331);
or U1982 (N_1982,In_2143,In_1091);
nand U1983 (N_1983,In_4413,In_1297);
xor U1984 (N_1984,In_1927,In_1279);
xor U1985 (N_1985,In_1946,N_377);
nand U1986 (N_1986,In_3587,In_1018);
or U1987 (N_1987,N_33,In_3891);
xor U1988 (N_1988,In_1148,In_299);
xor U1989 (N_1989,N_273,In_905);
xor U1990 (N_1990,N_445,N_27);
nor U1991 (N_1991,N_572,In_2603);
nor U1992 (N_1992,N_325,In_2947);
nor U1993 (N_1993,In_4894,In_4303);
xor U1994 (N_1994,In_997,In_2798);
nand U1995 (N_1995,N_839,In_820);
nor U1996 (N_1996,In_2764,N_845);
and U1997 (N_1997,In_1190,In_2172);
nor U1998 (N_1998,In_1301,In_3065);
and U1999 (N_1999,N_577,In_3740);
and U2000 (N_2000,N_1025,N_1389);
nor U2001 (N_2001,In_1376,N_1911);
nand U2002 (N_2002,In_3567,In_3201);
xor U2003 (N_2003,N_1063,In_4251);
nor U2004 (N_2004,In_706,N_1076);
nand U2005 (N_2005,In_31,In_3684);
xnor U2006 (N_2006,N_1992,In_1785);
or U2007 (N_2007,In_735,N_1386);
and U2008 (N_2008,In_758,N_1127);
nor U2009 (N_2009,N_1355,N_1701);
nand U2010 (N_2010,In_486,N_1308);
nor U2011 (N_2011,N_1198,N_707);
nor U2012 (N_2012,N_837,In_846);
or U2013 (N_2013,N_948,N_137);
xor U2014 (N_2014,In_4926,N_1404);
xor U2015 (N_2015,In_3143,N_301);
nor U2016 (N_2016,In_3014,In_3591);
nand U2017 (N_2017,N_1834,N_1618);
and U2018 (N_2018,In_759,In_4995);
nor U2019 (N_2019,In_747,In_117);
nor U2020 (N_2020,In_273,N_1362);
xor U2021 (N_2021,In_2168,In_3211);
and U2022 (N_2022,N_1828,In_1240);
and U2023 (N_2023,N_1210,In_3525);
nor U2024 (N_2024,In_3724,In_1848);
xnor U2025 (N_2025,N_380,In_3791);
nor U2026 (N_2026,N_1407,In_1578);
nand U2027 (N_2027,N_878,In_3500);
xnor U2028 (N_2028,In_1406,N_155);
nand U2029 (N_2029,In_4435,In_1595);
and U2030 (N_2030,N_1186,In_3474);
xnor U2031 (N_2031,N_482,N_120);
nand U2032 (N_2032,N_1239,In_2585);
and U2033 (N_2033,In_4145,In_1320);
and U2034 (N_2034,N_1642,In_2339);
and U2035 (N_2035,In_4512,In_290);
and U2036 (N_2036,N_1468,N_597);
xor U2037 (N_2037,In_1196,N_1034);
or U2038 (N_2038,N_1709,N_1016);
nor U2039 (N_2039,N_1622,In_4378);
or U2040 (N_2040,In_2987,In_3830);
nand U2041 (N_2041,N_1839,In_407);
xnor U2042 (N_2042,In_153,N_1744);
and U2043 (N_2043,N_1509,In_156);
or U2044 (N_2044,N_1360,N_1393);
xnor U2045 (N_2045,In_4074,N_976);
nor U2046 (N_2046,In_358,N_1026);
and U2047 (N_2047,N_1082,In_2793);
and U2048 (N_2048,N_1143,N_1817);
nor U2049 (N_2049,In_4373,N_366);
nor U2050 (N_2050,In_1153,In_2229);
and U2051 (N_2051,In_3432,In_281);
nand U2052 (N_2052,N_1685,In_3046);
or U2053 (N_2053,N_1876,N_1124);
xor U2054 (N_2054,In_3945,In_3366);
and U2055 (N_2055,N_1242,N_616);
xor U2056 (N_2056,N_1168,In_2041);
xor U2057 (N_2057,N_416,N_1254);
or U2058 (N_2058,In_791,N_553);
xnor U2059 (N_2059,N_131,N_932);
or U2060 (N_2060,In_3946,In_3294);
or U2061 (N_2061,N_1314,In_3413);
and U2062 (N_2062,N_1062,In_3374);
nand U2063 (N_2063,In_4959,In_967);
nand U2064 (N_2064,N_684,In_841);
nand U2065 (N_2065,In_3379,In_3582);
nand U2066 (N_2066,N_567,In_4012);
and U2067 (N_2067,N_1437,N_303);
or U2068 (N_2068,In_4320,N_1281);
nor U2069 (N_2069,N_1189,In_4547);
nor U2070 (N_2070,In_647,N_1222);
xor U2071 (N_2071,N_1994,N_1448);
and U2072 (N_2072,N_284,N_1800);
nand U2073 (N_2073,In_2574,N_1167);
xnor U2074 (N_2074,In_2929,N_76);
nor U2075 (N_2075,In_38,In_4039);
nand U2076 (N_2076,N_1496,In_3360);
xnor U2077 (N_2077,N_1234,In_4585);
nor U2078 (N_2078,N_1029,N_1451);
and U2079 (N_2079,N_1636,In_1214);
nand U2080 (N_2080,N_1096,N_955);
nor U2081 (N_2081,In_305,N_1379);
xnor U2082 (N_2082,In_2992,In_2703);
nor U2083 (N_2083,N_112,N_1273);
or U2084 (N_2084,N_1781,In_3270);
xor U2085 (N_2085,N_1401,N_294);
nor U2086 (N_2086,In_3425,N_415);
and U2087 (N_2087,In_2016,N_1780);
and U2088 (N_2088,In_3698,N_1521);
xor U2089 (N_2089,N_307,N_802);
nor U2090 (N_2090,In_4877,In_2717);
or U2091 (N_2091,In_2516,N_1741);
nand U2092 (N_2092,In_3554,N_678);
nand U2093 (N_2093,N_1993,N_1942);
nor U2094 (N_2094,N_1660,In_775);
or U2095 (N_2095,In_328,In_964);
nand U2096 (N_2096,In_2889,In_4985);
nor U2097 (N_2097,N_848,N_750);
nand U2098 (N_2098,N_1873,N_1647);
nand U2099 (N_2099,N_480,In_4879);
nor U2100 (N_2100,In_4338,N_1330);
and U2101 (N_2101,In_1058,N_1978);
and U2102 (N_2102,N_1558,N_985);
xor U2103 (N_2103,In_3153,N_1846);
or U2104 (N_2104,In_1791,N_1571);
xor U2105 (N_2105,N_1732,In_2398);
nand U2106 (N_2106,In_3783,N_1742);
and U2107 (N_2107,In_2028,N_1818);
nor U2108 (N_2108,In_349,In_4726);
nor U2109 (N_2109,N_426,In_2070);
nor U2110 (N_2110,N_1444,In_4624);
xor U2111 (N_2111,In_2171,N_1918);
xnor U2112 (N_2112,In_891,N_231);
or U2113 (N_2113,In_3165,In_1338);
nor U2114 (N_2114,In_1640,N_1632);
or U2115 (N_2115,In_4053,N_790);
nand U2116 (N_2116,In_1851,N_186);
nor U2117 (N_2117,In_2414,N_1698);
xnor U2118 (N_2118,N_1083,N_1888);
and U2119 (N_2119,In_670,N_442);
xnor U2120 (N_2120,In_845,In_3481);
and U2121 (N_2121,N_1339,In_2839);
nand U2122 (N_2122,N_725,In_3863);
xor U2123 (N_2123,In_639,N_1900);
and U2124 (N_2124,N_1365,N_459);
nand U2125 (N_2125,N_1551,In_1657);
xor U2126 (N_2126,N_1865,N_421);
xor U2127 (N_2127,N_62,In_700);
xor U2128 (N_2128,N_360,N_1678);
and U2129 (N_2129,N_1080,N_1680);
nand U2130 (N_2130,In_4536,In_1184);
nor U2131 (N_2131,In_235,N_1181);
or U2132 (N_2132,In_3702,In_2989);
nor U2133 (N_2133,In_3627,N_1756);
or U2134 (N_2134,N_30,N_1165);
or U2135 (N_2135,N_1373,In_1820);
and U2136 (N_2136,In_4657,N_1141);
nor U2137 (N_2137,N_1052,In_640);
nor U2138 (N_2138,In_2271,In_4943);
xor U2139 (N_2139,N_676,In_4951);
nor U2140 (N_2140,N_1072,In_2643);
xnor U2141 (N_2141,N_343,N_1208);
or U2142 (N_2142,In_1706,N_950);
nor U2143 (N_2143,N_1842,In_2669);
nor U2144 (N_2144,In_655,In_4854);
or U2145 (N_2145,In_529,In_3943);
and U2146 (N_2146,N_1172,N_1486);
and U2147 (N_2147,In_4741,In_4186);
or U2148 (N_2148,N_1270,In_4218);
xor U2149 (N_2149,In_2040,In_1212);
nand U2150 (N_2150,N_534,N_1795);
nor U2151 (N_2151,In_1754,N_989);
or U2152 (N_2152,N_1441,N_1623);
xor U2153 (N_2153,In_2477,In_2693);
nor U2154 (N_2154,N_1729,N_1023);
nor U2155 (N_2155,N_545,N_1798);
nor U2156 (N_2156,N_1537,In_1757);
or U2157 (N_2157,N_1728,In_2151);
xor U2158 (N_2158,N_1555,In_2331);
nor U2159 (N_2159,N_1580,In_2333);
or U2160 (N_2160,N_1439,N_1387);
xor U2161 (N_2161,In_1499,In_2372);
xnor U2162 (N_2162,N_1582,In_4518);
or U2163 (N_2163,In_4603,N_807);
xnor U2164 (N_2164,N_1803,In_4724);
nand U2165 (N_2165,N_1436,In_3412);
or U2166 (N_2166,N_513,In_4623);
or U2167 (N_2167,N_1306,In_3731);
and U2168 (N_2168,N_477,N_1249);
and U2169 (N_2169,In_4085,N_900);
nand U2170 (N_2170,N_176,N_1774);
or U2171 (N_2171,In_3287,In_1717);
xnor U2172 (N_2172,In_3470,In_2126);
nand U2173 (N_2173,N_1205,In_3156);
or U2174 (N_2174,N_474,N_1746);
nor U2175 (N_2175,In_3749,N_1032);
xor U2176 (N_2176,In_3300,In_220);
xor U2177 (N_2177,N_1670,In_815);
xnor U2178 (N_2178,N_1101,N_196);
nor U2179 (N_2179,In_2730,N_1870);
nor U2180 (N_2180,In_2396,N_1117);
nand U2181 (N_2181,In_888,In_1335);
and U2182 (N_2182,N_1227,In_4732);
xnor U2183 (N_2183,N_1821,In_605);
nor U2184 (N_2184,In_894,In_4510);
nand U2185 (N_2185,N_1119,In_298);
xor U2186 (N_2186,In_3180,N_1121);
and U2187 (N_2187,N_1786,In_1985);
nand U2188 (N_2188,In_2065,In_2434);
or U2189 (N_2189,In_1188,N_1138);
nand U2190 (N_2190,N_1563,N_1986);
nand U2191 (N_2191,In_2990,N_881);
nor U2192 (N_2192,In_3016,N_1000);
xor U2193 (N_2193,N_188,In_1418);
and U2194 (N_2194,In_3039,In_1701);
nor U2195 (N_2195,In_1347,In_2882);
nand U2196 (N_2196,N_718,N_1321);
or U2197 (N_2197,In_2543,N_1287);
nand U2198 (N_2198,N_1500,In_4102);
or U2199 (N_2199,N_1750,In_4936);
nand U2200 (N_2200,In_108,N_1323);
and U2201 (N_2201,N_1816,N_630);
nor U2202 (N_2202,N_799,In_2486);
or U2203 (N_2203,N_1326,N_1552);
nand U2204 (N_2204,N_1519,In_1991);
or U2205 (N_2205,N_554,N_991);
and U2206 (N_2206,In_1561,N_134);
and U2207 (N_2207,N_1699,In_3361);
and U2208 (N_2208,N_1714,In_1002);
and U2209 (N_2209,N_1629,N_1440);
and U2210 (N_2210,In_2895,In_2733);
or U2211 (N_2211,In_4142,N_1009);
xor U2212 (N_2212,N_683,In_4748);
xor U2213 (N_2213,In_75,N_891);
or U2214 (N_2214,N_1408,In_4840);
xnor U2215 (N_2215,N_786,In_2809);
and U2216 (N_2216,N_1140,N_1898);
and U2217 (N_2217,In_167,N_602);
nor U2218 (N_2218,In_364,In_916);
and U2219 (N_2219,N_1535,N_575);
nand U2220 (N_2220,N_16,N_1160);
nand U2221 (N_2221,N_1850,In_1923);
xnor U2222 (N_2222,In_4385,In_3653);
xor U2223 (N_2223,In_2623,N_54);
nand U2224 (N_2224,N_1224,N_1147);
xnor U2225 (N_2225,N_1293,N_1458);
or U2226 (N_2226,N_1645,In_4463);
or U2227 (N_2227,In_3667,In_2152);
xor U2228 (N_2228,N_613,In_1912);
xnor U2229 (N_2229,N_308,In_4164);
or U2230 (N_2230,In_3897,N_1202);
nand U2231 (N_2231,In_4685,In_2432);
nand U2232 (N_2232,In_1033,In_3158);
nor U2233 (N_2233,N_1216,N_1536);
nand U2234 (N_2234,In_2934,In_2357);
or U2235 (N_2235,N_1087,In_4478);
and U2236 (N_2236,In_4139,In_3075);
and U2237 (N_2237,In_1280,N_250);
nand U2238 (N_2238,In_3999,In_4753);
and U2239 (N_2239,N_1358,N_1429);
and U2240 (N_2240,In_3416,In_1218);
nor U2241 (N_2241,N_1997,N_1724);
and U2242 (N_2242,N_1206,N_411);
nor U2243 (N_2243,N_996,N_1664);
xnor U2244 (N_2244,N_1823,In_361);
or U2245 (N_2245,In_1958,In_4325);
and U2246 (N_2246,N_1768,N_818);
and U2247 (N_2247,N_727,N_1995);
nand U2248 (N_2248,In_2644,In_3518);
or U2249 (N_2249,N_1723,N_800);
nand U2250 (N_2250,N_496,N_1073);
nand U2251 (N_2251,N_1592,In_4561);
nand U2252 (N_2252,In_3212,In_4179);
and U2253 (N_2253,N_1331,In_403);
nand U2254 (N_2254,In_1461,N_1018);
xor U2255 (N_2255,N_1395,In_4361);
xnor U2256 (N_2256,In_187,N_883);
and U2257 (N_2257,In_1573,N_751);
or U2258 (N_2258,In_211,N_105);
xor U2259 (N_2259,In_4168,N_1132);
nand U2260 (N_2260,In_1157,N_456);
xor U2261 (N_2261,N_282,In_2404);
nand U2262 (N_2262,N_1303,In_3936);
nor U2263 (N_2263,N_1765,In_4824);
and U2264 (N_2264,In_1388,In_1489);
xnor U2265 (N_2265,N_1950,In_219);
or U2266 (N_2266,In_1213,In_2787);
nor U2267 (N_2267,N_540,In_3114);
nor U2268 (N_2268,In_1479,N_1882);
nand U2269 (N_2269,N_640,N_1556);
nor U2270 (N_2270,N_1484,N_8);
and U2271 (N_2271,In_2161,N_1548);
nor U2272 (N_2272,In_3238,N_1871);
and U2273 (N_2273,In_152,In_1558);
nand U2274 (N_2274,In_3488,N_1253);
nor U2275 (N_2275,N_585,In_1462);
xnor U2276 (N_2276,N_929,In_1813);
nor U2277 (N_2277,N_202,In_4485);
and U2278 (N_2278,N_1430,In_3710);
xnor U2279 (N_2279,In_1592,N_510);
nand U2280 (N_2280,In_552,In_4316);
nor U2281 (N_2281,N_190,In_3009);
or U2282 (N_2282,N_1098,N_1738);
nand U2283 (N_2283,In_790,In_668);
xor U2284 (N_2284,N_574,In_2021);
nor U2285 (N_2285,N_1754,N_1004);
nor U2286 (N_2286,N_1859,In_1546);
or U2287 (N_2287,N_1843,In_1009);
and U2288 (N_2288,In_1497,In_3025);
or U2289 (N_2289,N_700,N_987);
nor U2290 (N_2290,In_3350,In_4195);
nand U2291 (N_2291,In_4636,In_2621);
nor U2292 (N_2292,N_1184,In_2294);
nor U2293 (N_2293,N_652,In_3953);
or U2294 (N_2294,N_14,In_974);
and U2295 (N_2295,In_2718,N_1513);
nand U2296 (N_2296,N_1256,N_1973);
xnor U2297 (N_2297,N_1945,In_1224);
nor U2298 (N_2298,In_4321,N_830);
xor U2299 (N_2299,In_2157,In_2079);
xnor U2300 (N_2300,In_4318,In_736);
xor U2301 (N_2301,In_2738,In_801);
nor U2302 (N_2302,In_3293,In_3787);
or U2303 (N_2303,N_1193,In_3410);
nor U2304 (N_2304,In_2155,In_1332);
nor U2305 (N_2305,N_1782,N_1039);
or U2306 (N_2306,N_699,N_1185);
and U2307 (N_2307,In_2803,N_1835);
and U2308 (N_2308,N_1611,In_4258);
nand U2309 (N_2309,N_1111,In_3446);
or U2310 (N_2310,N_1413,N_1409);
and U2311 (N_2311,N_361,N_1244);
and U2312 (N_2312,N_828,N_924);
nor U2313 (N_2313,N_243,In_1311);
and U2314 (N_2314,In_4844,In_721);
nor U2315 (N_2315,In_3763,N_1110);
or U2316 (N_2316,N_1099,N_1764);
nor U2317 (N_2317,N_1802,In_4037);
nor U2318 (N_2318,In_3338,In_1980);
nor U2319 (N_2319,In_303,In_2720);
nor U2320 (N_2320,N_1020,N_1229);
nor U2321 (N_2321,In_921,N_1204);
and U2322 (N_2322,In_3646,In_3459);
and U2323 (N_2323,N_964,N_887);
and U2324 (N_2324,N_1731,N_1109);
nor U2325 (N_2325,N_479,N_1421);
nor U2326 (N_2326,N_520,N_1905);
nor U2327 (N_2327,N_229,N_804);
and U2328 (N_2328,In_4994,N_1616);
xor U2329 (N_2329,N_547,In_869);
nor U2330 (N_2330,N_1403,In_3959);
or U2331 (N_2331,In_418,N_90);
nor U2332 (N_2332,In_2514,In_2592);
nor U2333 (N_2333,N_1653,In_959);
nor U2334 (N_2334,N_1758,N_1418);
or U2335 (N_2335,N_814,In_1385);
and U2336 (N_2336,In_549,In_1880);
xnor U2337 (N_2337,In_2050,In_585);
or U2338 (N_2338,N_1872,In_3411);
or U2339 (N_2339,In_596,N_1338);
or U2340 (N_2340,N_730,N_1473);
or U2341 (N_2341,N_1848,In_4122);
or U2342 (N_2342,In_1667,N_7);
or U2343 (N_2343,N_767,N_642);
nand U2344 (N_2344,N_1820,N_1690);
nand U2345 (N_2345,In_1863,In_3818);
nand U2346 (N_2346,N_1874,N_1116);
and U2347 (N_2347,N_1959,N_1603);
or U2348 (N_2348,N_1917,In_4548);
nor U2349 (N_2349,N_1976,N_825);
nand U2350 (N_2350,N_1295,In_4066);
xor U2351 (N_2351,N_1385,N_379);
and U2352 (N_2352,N_146,In_1733);
and U2353 (N_2353,In_833,N_834);
nand U2354 (N_2354,In_3031,In_2826);
or U2355 (N_2355,In_2358,In_2233);
nor U2356 (N_2356,N_1767,N_1516);
xnor U2357 (N_2357,N_1836,In_3939);
or U2358 (N_2358,N_19,N_1019);
or U2359 (N_2359,N_1470,In_3668);
xnor U2360 (N_2360,N_915,In_2219);
nand U2361 (N_2361,In_4217,In_2485);
nor U2362 (N_2362,In_1588,N_441);
and U2363 (N_2363,N_1639,N_1845);
xor U2364 (N_2364,N_106,N_340);
xnor U2365 (N_2365,In_2877,N_1028);
or U2366 (N_2366,N_1231,N_240);
xor U2367 (N_2367,N_1190,N_1922);
or U2368 (N_2368,N_167,N_1203);
nor U2369 (N_2369,N_1094,N_1179);
or U2370 (N_2370,In_996,In_701);
and U2371 (N_2371,In_1349,In_1685);
or U2372 (N_2372,N_119,In_3880);
nor U2373 (N_2373,N_1493,N_685);
and U2374 (N_2374,In_2024,In_1256);
xnor U2375 (N_2375,In_265,N_1488);
nand U2376 (N_2376,N_20,N_1902);
xor U2377 (N_2377,N_1627,N_1027);
nor U2378 (N_2378,N_321,In_825);
nand U2379 (N_2379,N_569,N_260);
xor U2380 (N_2380,In_14,In_3678);
or U2381 (N_2381,In_4108,N_984);
xor U2382 (N_2382,N_69,In_1470);
nand U2383 (N_2383,N_1352,N_1588);
or U2384 (N_2384,In_2948,In_3473);
and U2385 (N_2385,In_466,N_226);
xnor U2386 (N_2386,In_4664,In_1594);
nor U2387 (N_2387,N_1183,N_204);
xnor U2388 (N_2388,In_380,In_61);
xor U2389 (N_2389,N_1753,In_2673);
nor U2390 (N_2390,In_1764,N_1745);
nand U2391 (N_2391,In_4041,N_1598);
nand U2392 (N_2392,In_2831,N_1417);
xnor U2393 (N_2393,N_1703,N_1152);
nand U2394 (N_2394,N_1380,N_1097);
nand U2395 (N_2395,In_1239,In_793);
or U2396 (N_2396,N_1941,N_1050);
nand U2397 (N_2397,N_1024,N_1469);
and U2398 (N_2398,In_4479,In_4509);
and U2399 (N_2399,In_621,In_1642);
xnor U2400 (N_2400,N_978,N_1763);
nand U2401 (N_2401,In_1881,N_1880);
nor U2402 (N_2402,N_1163,In_1453);
nand U2403 (N_2403,In_3682,N_1526);
nand U2404 (N_2404,In_4850,N_1384);
and U2405 (N_2405,In_3144,N_1672);
or U2406 (N_2406,In_2503,In_569);
nor U2407 (N_2407,In_4302,In_4638);
nor U2408 (N_2408,In_43,In_2078);
or U2409 (N_2409,In_4708,N_1483);
and U2410 (N_2410,In_600,N_1241);
nor U2411 (N_2411,In_2346,N_1498);
xnor U2412 (N_2412,N_1675,In_368);
nand U2413 (N_2413,N_65,N_1649);
nor U2414 (N_2414,N_1378,N_1171);
xor U2415 (N_2415,N_451,N_746);
nand U2416 (N_2416,In_2089,In_4100);
nand U2417 (N_2417,In_504,In_2924);
and U2418 (N_2418,N_365,N_1607);
or U2419 (N_2419,In_1278,N_717);
xnor U2420 (N_2420,In_4348,N_1071);
or U2421 (N_2421,In_4054,In_3821);
nor U2422 (N_2422,N_1879,In_4143);
or U2423 (N_2423,In_4886,In_2701);
xnor U2424 (N_2424,N_346,N_1161);
nor U2425 (N_2425,In_4771,In_2631);
nand U2426 (N_2426,N_972,In_145);
and U2427 (N_2427,N_492,In_3462);
and U2428 (N_2428,In_3466,N_53);
nand U2429 (N_2429,N_1681,In_2753);
and U2430 (N_2430,N_348,In_3430);
nand U2431 (N_2431,N_1734,N_1103);
and U2432 (N_2432,N_485,In_2454);
and U2433 (N_2433,N_1972,N_288);
nand U2434 (N_2434,In_1611,N_1946);
or U2435 (N_2435,In_28,N_89);
nand U2436 (N_2436,In_4696,N_551);
or U2437 (N_2437,In_832,N_1382);
nand U2438 (N_2438,N_1534,In_1602);
or U2439 (N_2439,In_4559,N_1658);
nand U2440 (N_2440,In_1322,In_4059);
or U2441 (N_2441,In_1158,N_779);
xnor U2442 (N_2442,In_2875,N_1329);
and U2443 (N_2443,N_1875,In_4488);
nand U2444 (N_2444,N_1878,In_465);
xor U2445 (N_2445,In_1649,In_3023);
xor U2446 (N_2446,In_4878,N_1079);
xor U2447 (N_2447,N_1532,In_3137);
xor U2448 (N_2448,In_4647,N_523);
xor U2449 (N_2449,In_952,In_1446);
or U2450 (N_2450,N_1896,N_1559);
nor U2451 (N_2451,N_439,In_2820);
nand U2452 (N_2452,N_1262,N_1688);
xnor U2453 (N_2453,In_1933,N_977);
and U2454 (N_2454,N_1300,N_1144);
nand U2455 (N_2455,In_4388,In_3172);
xor U2456 (N_2456,N_295,N_1497);
or U2457 (N_2457,In_2337,N_1086);
xnor U2458 (N_2458,N_605,N_1751);
nand U2459 (N_2459,N_144,In_3395);
xnor U2460 (N_2460,In_1658,In_4071);
and U2461 (N_2461,In_4368,N_733);
nand U2462 (N_2462,In_3051,N_1324);
or U2463 (N_2463,N_1517,In_3391);
nor U2464 (N_2464,N_851,In_2147);
and U2465 (N_2465,In_3615,In_1234);
and U2466 (N_2466,N_1676,In_2801);
nand U2467 (N_2467,In_580,In_1078);
and U2468 (N_2468,N_1869,N_285);
or U2469 (N_2469,In_3255,N_1313);
nand U2470 (N_2470,N_1529,In_3346);
or U2471 (N_2471,In_2602,In_2097);
and U2472 (N_2472,In_1830,N_1838);
or U2473 (N_2473,In_3876,In_1154);
or U2474 (N_2474,In_1139,N_1433);
nor U2475 (N_2475,N_443,In_4018);
and U2476 (N_2476,N_386,In_1046);
nand U2477 (N_2477,In_2325,N_1695);
or U2478 (N_2478,In_1631,In_4744);
nand U2479 (N_2479,In_4853,In_927);
xor U2480 (N_2480,N_1543,N_587);
and U2481 (N_2481,N_1354,In_1781);
and U2482 (N_2482,N_1065,N_1810);
nor U2483 (N_2483,In_3267,N_220);
and U2484 (N_2484,In_3202,In_3771);
and U2485 (N_2485,In_624,N_1969);
or U2486 (N_2486,In_292,In_1847);
or U2487 (N_2487,In_2142,N_1220);
or U2488 (N_2488,In_4000,In_2112);
nor U2489 (N_2489,In_900,N_1343);
or U2490 (N_2490,In_423,In_2997);
or U2491 (N_2491,In_2060,N_502);
or U2492 (N_2492,In_1537,In_4511);
and U2493 (N_2493,N_909,In_744);
xnor U2494 (N_2494,In_1035,N_269);
nand U2495 (N_2495,In_1389,In_760);
xnor U2496 (N_2496,In_2526,N_795);
nor U2497 (N_2497,N_1506,N_768);
or U2498 (N_2498,N_1507,N_1335);
xor U2499 (N_2499,In_534,N_1075);
xor U2500 (N_2500,In_2114,In_4101);
or U2501 (N_2501,In_3431,In_371);
nand U2502 (N_2502,N_221,N_1667);
nand U2503 (N_2503,N_1615,In_3660);
nor U2504 (N_2504,In_456,In_3247);
or U2505 (N_2505,In_675,N_517);
xnor U2506 (N_2506,N_1717,In_3777);
nand U2507 (N_2507,In_4050,In_1140);
and U2508 (N_2508,N_452,N_1078);
or U2509 (N_2509,In_1550,N_1868);
xnor U2510 (N_2510,N_268,N_741);
nor U2511 (N_2511,In_4092,N_797);
or U2512 (N_2512,In_3604,N_56);
nor U2513 (N_2513,In_1303,N_1791);
nor U2514 (N_2514,N_151,N_1022);
or U2515 (N_2515,N_706,N_1739);
nand U2516 (N_2516,In_3209,N_1567);
nand U2517 (N_2517,In_261,N_1466);
nand U2518 (N_2518,N_1936,In_4468);
and U2519 (N_2519,N_1064,In_3860);
or U2520 (N_2520,In_2462,N_1304);
nand U2521 (N_2521,In_501,N_1769);
or U2522 (N_2522,In_2228,In_2427);
nor U2523 (N_2523,In_4896,In_4333);
and U2524 (N_2524,In_2345,N_1612);
xnor U2525 (N_2525,N_1494,In_3260);
nor U2526 (N_2526,In_4430,In_2930);
nor U2527 (N_2527,N_1949,In_508);
xnor U2528 (N_2528,In_99,In_4064);
xnor U2529 (N_2529,In_676,In_1343);
or U2530 (N_2530,In_2439,In_4710);
nand U2531 (N_2531,In_346,N_297);
nand U2532 (N_2532,In_3042,N_1712);
nor U2533 (N_2533,N_1298,In_3246);
nand U2534 (N_2534,N_1561,In_2825);
nand U2535 (N_2535,In_4387,N_1427);
nand U2536 (N_2536,In_661,In_4459);
or U2537 (N_2537,In_4199,N_1638);
and U2538 (N_2538,In_4801,In_4313);
and U2539 (N_2539,N_1396,In_4230);
nor U2540 (N_2540,In_971,In_1613);
nand U2541 (N_2541,N_1916,In_1633);
and U2542 (N_2542,In_2415,N_1459);
xnor U2543 (N_2543,N_1760,N_1655);
xor U2544 (N_2544,In_1808,N_201);
and U2545 (N_2545,In_1377,N_866);
and U2546 (N_2546,In_2177,N_1170);
xnor U2547 (N_2547,N_1963,In_1086);
nor U2548 (N_2548,In_3249,In_2544);
and U2549 (N_2549,In_4530,In_544);
and U2550 (N_2550,In_1556,In_1945);
nand U2551 (N_2551,N_969,N_1748);
and U2552 (N_2552,N_1926,In_1193);
nor U2553 (N_2553,In_4618,In_2254);
xor U2554 (N_2554,In_2871,In_419);
nor U2555 (N_2555,In_3289,In_2743);
or U2556 (N_2556,N_1633,In_3584);
or U2557 (N_2557,N_1217,N_939);
xor U2558 (N_2558,In_3928,In_4319);
nor U2559 (N_2559,In_3489,N_784);
xor U2560 (N_2560,In_1202,N_1771);
xnor U2561 (N_2561,In_1999,N_1031);
and U2562 (N_2562,N_1708,N_1424);
or U2563 (N_2563,In_294,N_299);
nand U2564 (N_2564,N_1490,N_222);
nand U2565 (N_2565,In_1943,N_1472);
nor U2566 (N_2566,N_136,N_1414);
nand U2567 (N_2567,N_1277,In_1472);
and U2568 (N_2568,N_1620,N_1539);
nor U2569 (N_2569,In_1267,In_4044);
nand U2570 (N_2570,In_3119,N_1398);
or U2571 (N_2571,In_2806,In_568);
or U2572 (N_2572,In_2133,In_1939);
xor U2573 (N_2573,N_1041,In_3036);
nor U2574 (N_2574,In_2792,In_2572);
xnor U2575 (N_2575,N_1337,N_1937);
and U2576 (N_2576,N_1663,In_2207);
xor U2577 (N_2577,N_853,In_183);
nor U2578 (N_2578,N_1434,N_1679);
nand U2579 (N_2579,In_3742,N_404);
or U2580 (N_2580,N_1809,In_2985);
nand U2581 (N_2581,In_4574,N_1617);
nor U2582 (N_2582,N_17,In_1050);
xor U2583 (N_2583,In_623,In_87);
or U2584 (N_2584,In_2749,N_181);
or U2585 (N_2585,N_1861,In_499);
xnor U2586 (N_2586,In_2262,N_1697);
or U2587 (N_2587,In_2752,N_1431);
nor U2588 (N_2588,N_154,N_1822);
or U2589 (N_2589,In_3080,N_1252);
nand U2590 (N_2590,In_4243,N_1452);
nand U2591 (N_2591,In_1520,N_1736);
or U2592 (N_2592,N_986,N_1173);
nor U2593 (N_2593,In_4431,In_3752);
or U2594 (N_2594,In_1563,In_1583);
and U2595 (N_2595,In_3884,N_1689);
or U2596 (N_2596,In_3223,In_97);
nor U2597 (N_2597,In_2705,In_1208);
or U2598 (N_2598,N_1877,In_2468);
and U2599 (N_2599,N_1453,In_2174);
and U2600 (N_2600,In_3981,In_2554);
nor U2601 (N_2601,In_3079,N_353);
or U2602 (N_2602,In_3453,In_3146);
nand U2603 (N_2603,In_4591,In_844);
or U2604 (N_2604,N_1347,In_2378);
nor U2605 (N_2605,In_3526,In_4619);
nand U2606 (N_2606,N_1364,N_1626);
nor U2607 (N_2607,In_436,In_4712);
or U2608 (N_2608,In_2421,In_3078);
nor U2609 (N_2609,In_1941,N_1783);
nand U2610 (N_2610,In_2166,In_1625);
nand U2611 (N_2611,In_3922,In_540);
and U2612 (N_2612,In_3963,In_4489);
nand U2613 (N_2613,N_1333,N_1650);
nor U2614 (N_2614,In_3286,In_509);
xor U2615 (N_2615,In_4332,N_211);
xor U2616 (N_2616,N_1463,In_3010);
nand U2617 (N_2617,In_1567,In_2202);
xnor U2618 (N_2618,N_720,In_3400);
or U2619 (N_2619,N_1797,N_1464);
nor U2620 (N_2620,In_4607,N_1999);
xnor U2621 (N_2621,N_1899,In_3907);
nor U2622 (N_2622,N_860,N_1977);
nor U2623 (N_2623,In_2727,N_408);
nand U2624 (N_2624,In_2455,In_3806);
and U2625 (N_2625,N_135,In_713);
nor U2626 (N_2626,N_1212,In_3696);
or U2627 (N_2627,N_1807,In_1362);
nand U2628 (N_2628,N_170,N_347);
xor U2629 (N_2629,In_1976,In_1962);
and U2630 (N_2630,N_49,In_228);
or U2631 (N_2631,In_672,In_872);
nand U2632 (N_2632,In_1409,N_1457);
nand U2633 (N_2633,N_227,N_1108);
nand U2634 (N_2634,In_2843,In_1109);
xnor U2635 (N_2635,N_350,N_709);
nor U2636 (N_2636,N_1796,N_1608);
or U2637 (N_2637,N_687,In_3687);
and U2638 (N_2638,N_1970,In_1438);
nand U2639 (N_2639,In_1532,N_1938);
nand U2640 (N_2640,In_1862,In_3452);
nor U2641 (N_2641,In_3513,In_18);
nor U2642 (N_2642,N_1187,In_4534);
nand U2643 (N_2643,N_162,In_3419);
or U2644 (N_2644,N_1886,In_4751);
xor U2645 (N_2645,In_659,N_1508);
nor U2646 (N_2646,In_3728,N_438);
nand U2647 (N_2647,N_1017,In_1671);
nand U2648 (N_2648,N_1118,In_4455);
and U2649 (N_2649,In_2441,In_1638);
and U2650 (N_2650,In_4209,N_863);
and U2651 (N_2651,In_1966,N_1960);
nand U2652 (N_2652,N_579,In_2872);
xor U2653 (N_2653,N_1399,N_1827);
or U2654 (N_2654,In_3902,N_1299);
nor U2655 (N_2655,In_885,In_2478);
and U2656 (N_2656,N_1196,In_1553);
or U2657 (N_2657,In_4949,N_257);
or U2658 (N_2658,N_1353,In_4747);
xnor U2659 (N_2659,N_1952,In_4763);
and U2660 (N_2660,N_140,N_1684);
nand U2661 (N_2661,In_2225,In_3170);
nand U2662 (N_2662,N_1302,N_1049);
and U2663 (N_2663,N_1388,In_4312);
xnor U2664 (N_2664,In_2025,In_76);
or U2665 (N_2665,N_530,In_2467);
nor U2666 (N_2666,N_1007,In_4934);
nor U2667 (N_2667,N_1799,N_1855);
and U2668 (N_2668,N_1996,In_1668);
xnor U2669 (N_2669,In_4910,N_1266);
nand U2670 (N_2670,In_4471,N_1102);
and U2671 (N_2671,In_2417,In_969);
nand U2672 (N_2672,In_663,In_100);
and U2673 (N_2673,N_1282,N_701);
nor U2674 (N_2674,In_4170,N_1200);
and U2675 (N_2675,N_1178,In_1614);
xnor U2676 (N_2676,In_47,In_2510);
xnor U2677 (N_2677,In_2401,N_715);
or U2678 (N_2678,In_784,N_1478);
nor U2679 (N_2679,N_782,In_807);
nand U2680 (N_2680,In_2923,In_2667);
nand U2681 (N_2681,In_453,N_1283);
nand U2682 (N_2682,N_1126,N_1344);
nand U2683 (N_2683,N_72,In_589);
xor U2684 (N_2684,N_465,In_2314);
nand U2685 (N_2685,In_1787,N_1761);
or U2686 (N_2686,In_258,In_4238);
nor U2687 (N_2687,In_1410,In_2998);
and U2688 (N_2688,N_595,In_1143);
xnor U2689 (N_2689,N_1935,N_1133);
nand U2690 (N_2690,N_1665,In_3324);
or U2691 (N_2691,In_402,N_1909);
and U2692 (N_2692,In_1871,N_1565);
xor U2693 (N_2693,In_3099,N_1849);
xnor U2694 (N_2694,In_268,In_692);
xor U2695 (N_2695,N_1966,N_1280);
xor U2696 (N_2696,N_1166,In_1290);
nand U2697 (N_2697,N_1258,N_1940);
xor U2698 (N_2698,In_686,In_4746);
or U2699 (N_2699,In_3664,N_549);
or U2700 (N_2700,In_4914,In_1049);
or U2701 (N_2701,N_1260,In_994);
nor U2702 (N_2702,N_1438,In_2009);
nand U2703 (N_2703,In_4405,In_1104);
nand U2704 (N_2704,N_1276,In_4495);
nor U2705 (N_2705,In_1211,N_601);
or U2706 (N_2706,N_1271,N_1621);
nand U2707 (N_2707,N_1228,In_2309);
xor U2708 (N_2708,In_924,N_1250);
or U2709 (N_2709,In_4073,N_1965);
xnor U2710 (N_2710,N_1135,N_302);
xnor U2711 (N_2711,N_1934,In_3508);
nand U2712 (N_2712,N_865,In_226);
nand U2713 (N_2713,In_275,N_1491);
nor U2714 (N_2714,In_1877,In_3814);
nor U2715 (N_2715,N_1289,N_920);
or U2716 (N_2716,N_1805,N_634);
xor U2717 (N_2717,N_1720,In_202);
xnor U2718 (N_2718,In_3995,N_1602);
or U2719 (N_2719,In_1723,N_46);
and U2720 (N_2720,In_1152,N_1342);
nor U2721 (N_2721,N_1814,N_1345);
and U2722 (N_2722,In_3389,N_1422);
xor U2723 (N_2723,In_96,N_1288);
or U2724 (N_2724,In_1014,In_399);
nor U2725 (N_2725,In_3579,N_609);
or U2726 (N_2726,N_1328,In_4273);
nor U2727 (N_2727,N_1197,N_1854);
xnor U2728 (N_2728,In_2136,In_1494);
or U2729 (N_2729,In_3451,N_1221);
or U2730 (N_2730,In_3726,N_246);
nor U2731 (N_2731,N_1528,In_4228);
nor U2732 (N_2732,N_1243,In_4776);
xor U2733 (N_2733,N_1752,N_742);
and U2734 (N_2734,In_828,N_1363);
or U2735 (N_2735,N_1566,In_2684);
nor U2736 (N_2736,In_1610,N_1844);
xor U2737 (N_2737,N_47,In_4987);
or U2738 (N_2738,In_677,N_1346);
or U2739 (N_2739,In_90,In_4458);
or U2740 (N_2740,N_50,N_1255);
xor U2741 (N_2741,In_4679,N_1716);
or U2742 (N_2742,N_1933,In_255);
nor U2743 (N_2743,N_1511,N_385);
and U2744 (N_2744,N_312,N_387);
xor U2745 (N_2745,In_1887,In_2907);
or U2746 (N_2746,N_1495,N_486);
nor U2747 (N_2747,In_4160,N_646);
nor U2748 (N_2748,In_2104,In_876);
and U2749 (N_2749,In_3700,In_1227);
xor U2750 (N_2750,N_905,N_1053);
and U2751 (N_2751,N_1462,N_1001);
and U2752 (N_2752,N_1913,In_4920);
nor U2753 (N_2753,N_410,N_1445);
xor U2754 (N_2754,N_1214,N_1148);
nand U2755 (N_2755,N_576,N_1696);
nor U2756 (N_2756,N_1852,N_236);
xor U2757 (N_2757,In_1639,In_2666);
nor U2758 (N_2758,N_1177,N_728);
and U2759 (N_2759,N_74,In_1235);
and U2760 (N_2760,N_1014,In_447);
and U2761 (N_2761,In_1591,N_1901);
and U2762 (N_2762,N_1371,In_2660);
or U2763 (N_2763,In_1603,In_3);
xnor U2764 (N_2764,N_770,In_1114);
nand U2765 (N_2765,N_925,In_4200);
xnor U2766 (N_2766,In_634,In_3685);
nand U2767 (N_2767,N_397,In_193);
nor U2768 (N_2768,N_125,N_1238);
and U2769 (N_2769,N_103,In_4023);
nand U2770 (N_2770,N_1903,N_1785);
nand U2771 (N_2771,In_3866,In_995);
xnor U2772 (N_2772,N_1201,N_1069);
nand U2773 (N_2773,In_1415,In_4474);
and U2774 (N_2774,N_304,In_3778);
and U2775 (N_2775,N_1394,N_338);
nor U2776 (N_2776,N_1188,In_1562);
nor U2777 (N_2777,N_249,N_1883);
xor U2778 (N_2778,In_699,In_3553);
and U2779 (N_2779,N_619,N_908);
or U2780 (N_2780,In_1712,In_1231);
nand U2781 (N_2781,In_896,In_3720);
xnor U2782 (N_2782,In_2522,N_1248);
nor U2783 (N_2783,In_839,N_1356);
xor U2784 (N_2784,N_1410,In_2884);
xor U2785 (N_2785,N_344,In_4016);
nor U2786 (N_2786,In_340,In_797);
nand U2787 (N_2787,N_1659,In_2124);
nor U2788 (N_2788,N_413,N_1291);
or U2789 (N_2789,In_252,In_4978);
xnor U2790 (N_2790,N_4,In_3217);
and U2791 (N_2791,N_899,In_4056);
nand U2792 (N_2792,N_600,In_842);
nor U2793 (N_2793,N_1547,N_1586);
nor U2794 (N_2794,In_428,N_1893);
nand U2795 (N_2795,N_1784,N_6);
or U2796 (N_2796,N_1630,N_1856);
or U2797 (N_2797,N_1021,In_1445);
nand U2798 (N_2798,N_810,In_2940);
or U2799 (N_2799,N_1981,N_1577);
nor U2800 (N_2800,N_352,N_877);
nand U2801 (N_2801,In_919,In_2678);
nor U2802 (N_2802,N_1153,In_991);
and U2803 (N_2803,In_309,N_677);
xor U2804 (N_2804,N_1593,N_1081);
xor U2805 (N_2805,In_2744,In_2344);
nand U2806 (N_2806,In_696,In_4451);
and U2807 (N_2807,N_1369,N_262);
xor U2808 (N_2808,N_1247,In_4543);
or U2809 (N_2809,N_812,In_4808);
or U2810 (N_2810,N_1157,N_1705);
nand U2811 (N_2811,In_4197,In_4482);
nand U2812 (N_2812,N_1290,In_2746);
nand U2813 (N_2813,In_776,In_4537);
xor U2814 (N_2814,In_1160,In_83);
or U2815 (N_2815,In_1268,In_1559);
and U2816 (N_2816,N_1296,In_4262);
nor U2817 (N_2817,In_3463,N_396);
and U2818 (N_2818,In_834,N_1095);
xnor U2819 (N_2819,N_1568,In_3331);
xnor U2820 (N_2820,In_4667,In_4150);
xnor U2821 (N_2821,N_1625,In_2983);
nor U2822 (N_2822,In_4562,In_3885);
xor U2823 (N_2823,N_1770,In_49);
and U2824 (N_2824,In_91,N_1884);
or U2825 (N_2825,In_4625,N_57);
nor U2826 (N_2826,N_566,N_1562);
or U2827 (N_2827,N_1112,In_3837);
nor U2828 (N_2828,In_2338,N_1002);
or U2829 (N_2829,N_1815,In_703);
and U2830 (N_2830,N_918,N_1546);
nor U2831 (N_2831,In_1473,N_1985);
nand U2832 (N_2832,N_1641,In_1179);
nor U2833 (N_2833,In_3502,In_2069);
xor U2834 (N_2834,In_2505,In_4522);
nand U2835 (N_2835,In_113,N_1060);
or U2836 (N_2836,N_704,In_4131);
nand U2837 (N_2837,N_1156,In_485);
nand U2838 (N_2838,N_1091,In_494);
or U2839 (N_2839,N_1553,In_4298);
xnor U2840 (N_2840,In_3109,N_884);
nand U2841 (N_2841,In_366,In_2269);
and U2842 (N_2842,In_2724,N_1435);
nor U2843 (N_2843,N_792,In_3037);
or U2844 (N_2844,In_1648,In_3171);
xnor U2845 (N_2845,In_439,In_2719);
or U2846 (N_2846,N_1375,N_356);
nand U2847 (N_2847,N_803,In_1130);
and U2848 (N_2848,N_1927,N_740);
and U2849 (N_2849,N_1668,N_975);
xnor U2850 (N_2850,N_1376,In_2527);
xnor U2851 (N_2851,N_1778,N_734);
nand U2852 (N_2852,In_208,N_10);
or U2853 (N_2853,N_1011,In_4260);
or U2854 (N_2854,N_322,In_468);
nand U2855 (N_2855,In_437,N_405);
xnor U2856 (N_2856,N_469,In_3060);
xor U2857 (N_2857,In_3261,In_3961);
and U2858 (N_2858,In_2001,N_1476);
and U2859 (N_2859,N_504,In_3581);
xnor U2860 (N_2860,N_75,N_237);
nor U2861 (N_2861,N_1987,N_1826);
nor U2862 (N_2862,N_1162,N_663);
or U2863 (N_2863,N_1005,N_1545);
nand U2864 (N_2864,N_1853,In_1771);
nor U2865 (N_2865,In_2586,N_1549);
or U2866 (N_2866,N_550,In_1059);
or U2867 (N_2867,In_4911,N_36);
nor U2868 (N_2868,In_4291,N_1841);
or U2869 (N_2869,N_1051,In_1403);
xnor U2870 (N_2870,N_1572,In_1711);
nor U2871 (N_2871,In_3869,N_1599);
and U2872 (N_2872,In_1824,In_3421);
xor U2873 (N_2873,In_4119,In_865);
or U2874 (N_2874,N_1106,In_1882);
xor U2875 (N_2875,N_1953,In_4717);
nand U2876 (N_2876,In_2925,N_1657);
and U2877 (N_2877,N_544,N_1232);
and U2878 (N_2878,In_270,N_611);
nor U2879 (N_2879,N_1361,In_4687);
nor U2880 (N_2880,In_2908,In_3694);
and U2881 (N_2881,N_189,In_1921);
or U2882 (N_2882,In_4357,In_269);
and U2883 (N_2883,In_3775,N_1585);
nand U2884 (N_2884,In_633,In_2011);
nand U2885 (N_2885,In_3774,In_4990);
nand U2886 (N_2886,In_1660,N_1787);
nor U2887 (N_2887,N_1857,In_1284);
and U2888 (N_2888,In_126,In_1330);
and U2889 (N_2889,N_857,N_1406);
nand U2890 (N_2890,N_1793,In_3542);
xnor U2891 (N_2891,In_3846,N_681);
nand U2892 (N_2892,In_637,N_1426);
nor U2893 (N_2893,N_1213,N_1904);
xor U2894 (N_2894,In_2525,N_1357);
and U2895 (N_2895,In_586,N_952);
or U2896 (N_2896,N_529,In_2208);
xnor U2897 (N_2897,N_1656,In_852);
nand U2898 (N_2898,In_3630,In_4268);
and U2899 (N_2899,N_1704,N_1801);
or U2900 (N_2900,N_1492,In_4573);
nand U2901 (N_2901,In_3174,In_1997);
nor U2902 (N_2902,In_510,In_4645);
nand U2903 (N_2903,In_3901,In_348);
xor U2904 (N_2904,N_1145,N_327);
nor U2905 (N_2905,N_643,N_1584);
and U2906 (N_2906,N_422,In_2092);
nor U2907 (N_2907,In_3262,In_2051);
and U2908 (N_2908,In_980,N_1640);
nand U2909 (N_2909,In_131,In_2160);
nor U2910 (N_2910,N_79,N_1530);
or U2911 (N_2911,N_1485,In_3633);
xor U2912 (N_2912,N_93,In_2188);
xnor U2913 (N_2913,In_2212,N_1596);
xor U2914 (N_2914,N_835,In_4979);
nor U2915 (N_2915,In_2470,In_3032);
xor U2916 (N_2916,In_3882,In_1319);
nand U2917 (N_2917,In_1118,In_1266);
nor U2918 (N_2918,In_1859,In_2986);
xnor U2919 (N_2919,In_2370,N_1367);
xnor U2920 (N_2920,N_1077,N_1867);
nor U2921 (N_2921,N_1840,In_1507);
nor U2922 (N_2922,N_1043,In_1483);
and U2923 (N_2923,In_4456,In_3199);
nor U2924 (N_2924,In_3636,In_3712);
xor U2925 (N_2925,In_4125,In_330);
and U2926 (N_2926,In_2974,N_1325);
or U2927 (N_2927,N_983,In_1321);
nor U2928 (N_2928,N_564,N_1811);
nand U2929 (N_2929,N_1951,In_3753);
nand U2930 (N_2930,In_687,In_2020);
nor U2931 (N_2931,N_1939,In_2854);
nor U2932 (N_2932,N_558,N_736);
xnor U2933 (N_2933,N_1540,N_1998);
xnor U2934 (N_2934,In_2125,In_814);
xnor U2935 (N_2935,N_548,N_1792);
nand U2936 (N_2936,N_1315,N_1847);
nand U2937 (N_2937,N_1037,N_1691);
nand U2938 (N_2938,N_198,N_1044);
nor U2939 (N_2939,N_419,N_1146);
nand U2940 (N_2940,N_859,N_1693);
and U2941 (N_2941,N_1230,N_592);
xor U2942 (N_2942,N_1601,N_1637);
nand U2943 (N_2943,In_4207,In_2562);
and U2944 (N_2944,N_319,In_256);
and U2945 (N_2945,In_3917,N_1390);
xnor U2946 (N_2946,In_4001,N_244);
xor U2947 (N_2947,N_1215,N_399);
or U2948 (N_2948,N_603,In_4155);
or U2949 (N_2949,N_109,N_1415);
and U2950 (N_2950,In_479,In_1542);
or U2951 (N_2951,In_2961,N_1958);
nor U2952 (N_2952,N_1522,In_708);
and U2953 (N_2953,N_1610,In_3590);
nor U2954 (N_2954,In_850,In_582);
nor U2955 (N_2955,In_917,In_2975);
xor U2956 (N_2956,N_1722,In_3790);
nor U2957 (N_2957,N_1139,In_3649);
nand U2958 (N_2958,N_516,N_1432);
and U2959 (N_2959,In_4470,N_1948);
nor U2960 (N_2960,In_1478,N_1154);
or U2961 (N_2961,N_1336,N_941);
and U2962 (N_2962,N_1662,In_1873);
or U2963 (N_2963,In_20,N_1643);
or U2964 (N_2964,In_3064,In_1521);
and U2965 (N_2965,N_1199,N_1673);
nor U2966 (N_2966,N_1310,In_999);
nand U2967 (N_2967,N_1068,In_2690);
xor U2968 (N_2968,In_1680,N_3);
and U2969 (N_2969,N_1105,N_115);
and U2970 (N_2970,N_362,In_3723);
nor U2971 (N_2971,N_936,In_3536);
and U2972 (N_2972,N_1512,N_1392);
nor U2973 (N_2973,In_2706,In_3050);
nand U2974 (N_2974,N_1164,N_394);
xor U2975 (N_2975,In_1555,In_2382);
xnor U2976 (N_2976,N_515,N_1499);
and U2977 (N_2977,N_1743,N_949);
xnor U2978 (N_2978,In_1903,N_781);
or U2979 (N_2979,In_1257,N_1058);
nor U2980 (N_2980,N_1461,In_4407);
nand U2981 (N_2981,In_982,N_808);
xor U2982 (N_2982,N_1481,In_3505);
or U2983 (N_2983,N_1825,N_1450);
or U2984 (N_2984,N_37,In_1828);
nor U2985 (N_2985,N_1442,N_1925);
xnor U2986 (N_2986,N_911,In_751);
nand U2987 (N_2987,In_4992,In_2984);
nand U2988 (N_2988,N_1134,N_1887);
nand U2989 (N_2989,N_1515,In_2300);
or U2990 (N_2990,N_43,N_875);
or U2991 (N_2991,N_1635,N_1735);
or U2992 (N_2992,In_4461,In_1401);
nor U2993 (N_2993,In_4128,N_1416);
or U2994 (N_2994,In_2312,N_207);
and U2995 (N_2995,N_1219,In_1259);
nand U2996 (N_2996,N_641,N_774);
or U2997 (N_2997,N_1707,N_1150);
nor U2998 (N_2998,In_3768,N_1122);
or U2999 (N_2999,N_1504,In_2480);
nor U3000 (N_3000,N_2200,N_757);
nand U3001 (N_3001,N_940,N_2932);
and U3002 (N_3002,N_2487,N_2139);
nor U3003 (N_3003,N_1864,N_2961);
nand U3004 (N_3004,N_2651,N_2928);
nand U3005 (N_3005,N_1411,N_862);
nor U3006 (N_3006,N_1114,N_1824);
nand U3007 (N_3007,N_2413,N_944);
xor U3008 (N_3008,In_2582,N_1501);
and U3009 (N_3009,N_2155,In_1397);
or U3010 (N_3010,In_4917,N_2904);
and U3011 (N_3011,In_3799,N_2105);
or U3012 (N_3012,In_149,N_2809);
nand U3013 (N_3013,N_2181,N_1912);
nand U3014 (N_3014,N_1525,N_1070);
nor U3015 (N_3015,N_1209,N_2398);
xor U3016 (N_3016,In_1364,In_3906);
nor U3017 (N_3017,N_2660,N_274);
or U3018 (N_3018,In_3612,N_1003);
nor U3019 (N_3019,In_649,In_3329);
nand U3020 (N_3020,In_1195,In_317);
nand U3021 (N_3021,In_4837,N_2521);
nor U3022 (N_3022,In_4846,N_615);
xnor U3023 (N_3023,N_166,N_2441);
nor U3024 (N_3024,In_1908,In_1222);
nand U3025 (N_3025,N_2842,In_4182);
and U3026 (N_3026,N_2983,In_836);
nand U3027 (N_3027,N_2254,N_2871);
or U3028 (N_3028,N_2552,N_1048);
nand U3029 (N_3029,N_440,N_1726);
or U3030 (N_3030,N_2722,In_1589);
nand U3031 (N_3031,N_2699,In_2351);
nand U3032 (N_3032,N_1046,In_1823);
xor U3033 (N_3033,In_21,In_3011);
and U3034 (N_3034,N_2801,N_2050);
xor U3035 (N_3035,N_481,N_819);
nand U3036 (N_3036,N_2352,N_2889);
nor U3037 (N_3037,N_2112,N_2161);
or U3038 (N_3038,N_1159,N_2193);
nor U3039 (N_3039,N_2629,N_1120);
or U3040 (N_3040,N_1142,N_2601);
nand U3041 (N_3041,N_71,In_3447);
nand U3042 (N_3042,N_631,In_2397);
nor U3043 (N_3043,N_2078,In_4454);
nor U3044 (N_3044,N_2779,N_2606);
xor U3045 (N_3045,N_942,N_2704);
and U3046 (N_3046,N_2018,In_669);
nand U3047 (N_3047,N_2729,N_1318);
and U3048 (N_3048,N_2369,N_2147);
and U3049 (N_3049,N_2271,In_174);
nor U3050 (N_3050,In_4088,In_4411);
or U3051 (N_3051,N_2348,N_2676);
or U3052 (N_3052,N_174,N_2100);
and U3053 (N_3053,N_2357,N_2617);
nand U3054 (N_3054,N_2519,In_2105);
nand U3055 (N_3055,In_4013,In_2802);
xnor U3056 (N_3056,In_2280,N_2577);
and U3057 (N_3057,In_1285,N_2144);
xnor U3058 (N_3058,N_2364,N_2775);
or U3059 (N_3059,N_1631,In_2596);
nor U3060 (N_3060,N_2071,N_1984);
nor U3061 (N_3061,N_1837,N_1762);
and U3062 (N_3062,In_1374,N_2136);
and U3063 (N_3063,N_1652,N_2732);
xnor U3064 (N_3064,N_2120,In_1769);
and U3065 (N_3065,N_1038,N_1446);
or U3066 (N_3066,In_1142,N_2907);
and U3067 (N_3067,N_2150,N_1383);
and U3068 (N_3068,N_2879,N_2500);
or U3069 (N_3069,N_2745,N_2448);
and U3070 (N_3070,In_1223,N_138);
or U3071 (N_3071,In_3441,N_289);
xor U3072 (N_3072,N_1502,N_2310);
or U3073 (N_3073,N_1013,N_1619);
or U3074 (N_3074,In_4069,N_2894);
nand U3075 (N_3075,N_2657,N_2276);
nor U3076 (N_3076,In_40,N_902);
or U3077 (N_3077,N_2965,N_1920);
xnor U3078 (N_3078,N_2232,N_1895);
nand U3079 (N_3079,N_2472,N_245);
xnor U3080 (N_3080,N_1351,In_1748);
nor U3081 (N_3081,N_1510,N_1862);
and U3082 (N_3082,N_2003,N_2399);
xnor U3083 (N_3083,N_1240,In_2960);
nor U3084 (N_3084,N_2687,N_2291);
nor U3085 (N_3085,N_2851,N_2517);
xor U3086 (N_3086,N_2949,In_3095);
xnor U3087 (N_3087,In_4838,N_2114);
nand U3088 (N_3088,N_1316,N_2571);
and U3089 (N_3089,N_1480,N_679);
or U3090 (N_3090,N_2402,In_4165);
or U3091 (N_3091,N_2567,N_1591);
nor U3092 (N_3092,N_1085,N_1514);
nand U3093 (N_3093,N_1123,N_2469);
nor U3094 (N_3094,N_910,In_393);
nand U3095 (N_3095,N_2036,N_2383);
xnor U3096 (N_3096,In_4804,N_2211);
or U3097 (N_3097,N_1957,N_2757);
nor U3098 (N_3098,N_2059,In_42);
xnor U3099 (N_3099,N_2490,In_2636);
nand U3100 (N_3100,N_2848,N_1819);
and U3101 (N_3101,N_817,N_1010);
nor U3102 (N_3102,N_1964,N_1278);
or U3103 (N_3103,N_2578,N_1628);
xor U3104 (N_3104,In_429,N_2828);
and U3105 (N_3105,In_171,In_4257);
and U3106 (N_3106,N_1340,In_3560);
and U3107 (N_3107,N_2605,In_4544);
or U3108 (N_3108,In_2512,In_645);
nand U3109 (N_3109,N_1008,N_1381);
nor U3110 (N_3110,In_3111,N_627);
nor U3111 (N_3111,N_406,N_2381);
xor U3112 (N_3112,N_2066,In_1064);
nand U3113 (N_3113,N_2432,N_2429);
nand U3114 (N_3114,N_2716,N_690);
or U3115 (N_3115,N_1113,N_2602);
xnor U3116 (N_3116,N_1858,N_2881);
nor U3117 (N_3117,N_2248,N_2055);
nor U3118 (N_3118,N_2479,N_2234);
xnor U3119 (N_3119,N_2409,In_307);
xnor U3120 (N_3120,N_1980,N_2088);
and U3121 (N_3121,In_3780,N_2591);
and U3122 (N_3122,In_638,N_2482);
or U3123 (N_3123,N_102,N_2223);
nand U3124 (N_3124,In_1309,In_808);
or U3125 (N_3125,N_2192,N_555);
xnor U3126 (N_3126,In_4051,N_2467);
nor U3127 (N_3127,In_4493,In_1459);
or U3128 (N_3128,In_2471,N_2878);
and U3129 (N_3129,N_108,N_655);
nor U3130 (N_3130,N_695,In_2647);
and U3131 (N_3131,In_3175,N_2781);
xor U3132 (N_3132,N_2721,N_2177);
nor U3133 (N_3133,N_2195,N_2309);
nand U3134 (N_3134,N_2044,N_1775);
nor U3135 (N_3135,N_2133,In_2449);
xor U3136 (N_3136,N_1263,N_2864);
nor U3137 (N_3137,N_556,N_752);
nor U3138 (N_3138,N_2401,N_1055);
xnor U3139 (N_3139,In_4289,In_609);
and U3140 (N_3140,N_1225,N_2786);
nand U3141 (N_3141,N_2021,N_2374);
xor U3142 (N_3142,In_1047,N_218);
xor U3143 (N_3143,N_2987,N_1733);
and U3144 (N_3144,N_483,N_251);
xnor U3145 (N_3145,N_1669,N_2094);
xor U3146 (N_3146,N_1806,N_1503);
and U3147 (N_3147,N_2324,In_2476);
nor U3148 (N_3148,N_1921,N_2640);
nand U3149 (N_3149,N_2958,N_1275);
or U3150 (N_3150,In_941,N_2408);
nand U3151 (N_3151,N_2772,N_2559);
or U3152 (N_3152,N_2977,N_2307);
and U3153 (N_3153,N_629,N_1402);
xnor U3154 (N_3154,N_2865,N_2516);
nand U3155 (N_3155,N_2321,N_2116);
nor U3156 (N_3156,N_462,N_2385);
or U3157 (N_3157,N_2455,N_2734);
nand U3158 (N_3158,N_2030,N_2344);
nand U3159 (N_3159,N_1047,In_1814);
or U3160 (N_3160,N_163,N_214);
nand U3161 (N_3161,In_2557,N_2111);
xor U3162 (N_3162,N_2818,N_2284);
nand U3163 (N_3163,N_2471,N_2572);
and U3164 (N_3164,N_2663,In_4417);
nand U3165 (N_3165,N_1035,N_34);
nor U3166 (N_3166,In_2561,N_1812);
nand U3167 (N_3167,N_2157,N_2224);
nor U3168 (N_3168,N_2944,N_1412);
nand U3169 (N_3169,In_2893,N_2043);
and U3170 (N_3170,N_1067,N_2658);
and U3171 (N_3171,N_2117,In_805);
xor U3172 (N_3172,N_2635,N_1851);
nor U3173 (N_3173,N_2045,In_3022);
and U3174 (N_3174,N_2178,In_2252);
xor U3175 (N_3175,N_2866,N_2236);
nor U3176 (N_3176,N_2146,N_2199);
xor U3177 (N_3177,In_3894,N_2885);
xnor U3178 (N_3178,In_1134,N_2491);
nor U3179 (N_3179,N_2870,N_1341);
nor U3180 (N_3180,N_2038,In_3824);
xnor U3181 (N_3181,N_2082,N_1467);
xnor U3182 (N_3182,N_2953,N_2085);
nor U3183 (N_3183,N_2218,N_2679);
xnor U3184 (N_3184,N_2266,N_2047);
and U3185 (N_3185,In_357,In_4376);
xor U3186 (N_3186,N_2544,N_2267);
xnor U3187 (N_3187,In_3842,N_2072);
nand U3188 (N_3188,N_2711,N_2168);
xnor U3189 (N_3189,N_1554,In_3102);
or U3190 (N_3190,N_1990,N_2574);
and U3191 (N_3191,N_1988,In_1900);
or U3192 (N_3192,N_1956,In_3546);
or U3193 (N_3193,N_1646,N_2361);
or U3194 (N_3194,N_2615,In_3695);
nor U3195 (N_3195,N_2091,In_2692);
or U3196 (N_3196,N_2214,N_2566);
xor U3197 (N_3197,N_2620,N_2262);
and U3198 (N_3198,In_4594,N_2329);
or U3199 (N_3199,N_2210,N_2924);
and U3200 (N_3200,In_374,N_1066);
and U3201 (N_3201,N_2610,N_2843);
xor U3202 (N_3202,N_2543,In_1236);
and U3203 (N_3203,N_2684,N_2918);
xnor U3204 (N_3204,In_922,N_2697);
xor U3205 (N_3205,N_2034,N_2302);
xnor U3206 (N_3206,N_1654,N_2733);
nor U3207 (N_3207,N_2215,N_2850);
and U3208 (N_3208,N_2555,N_2283);
xnor U3209 (N_3209,In_175,N_2826);
xnor U3210 (N_3210,N_2993,N_2176);
xnor U3211 (N_3211,N_2138,In_960);
nand U3212 (N_3212,N_2581,N_1962);
nand U3213 (N_3213,N_2354,N_1334);
and U3214 (N_3214,N_2783,In_3393);
and U3215 (N_3215,N_2217,N_1766);
or U3216 (N_3216,N_2647,N_2394);
nor U3217 (N_3217,In_1683,N_2418);
and U3218 (N_3218,N_2009,N_2474);
or U3219 (N_3219,In_928,In_4822);
and U3220 (N_3220,In_1775,N_1056);
or U3221 (N_3221,N_2836,In_1340);
xor U3222 (N_3222,N_2747,N_2109);
or U3223 (N_3223,N_2057,N_2189);
nand U3224 (N_3224,N_1700,N_2815);
and U3225 (N_3225,N_2511,N_2565);
and U3226 (N_3226,N_2728,N_2718);
xor U3227 (N_3227,N_2494,N_1130);
nand U3228 (N_3228,N_35,In_1457);
or U3229 (N_3229,N_2506,N_2410);
nand U3230 (N_3230,N_2868,In_1738);
xnor U3231 (N_3231,N_2143,In_4419);
nand U3232 (N_3232,N_2631,In_4790);
nor U3233 (N_3233,N_893,N_2664);
nand U3234 (N_3234,In_352,N_2792);
xor U3235 (N_3235,N_2159,N_1889);
nand U3236 (N_3236,In_1065,N_2089);
nor U3237 (N_3237,In_3599,In_3133);
xor U3238 (N_3238,N_2252,In_3550);
xor U3239 (N_3239,In_408,N_2513);
nor U3240 (N_3240,N_1661,In_2413);
nor U3241 (N_3241,N_2892,In_977);
or U3242 (N_3242,N_2514,In_2360);
xor U3243 (N_3243,N_2332,N_487);
or U3244 (N_3244,N_2717,N_2065);
xor U3245 (N_3245,N_2293,In_386);
and U3246 (N_3246,N_2073,In_4882);
and U3247 (N_3247,In_3007,In_4787);
nand U3248 (N_3248,N_1115,N_427);
or U3249 (N_3249,In_848,N_2744);
xor U3250 (N_3250,N_2345,In_4627);
nand U3251 (N_3251,N_2202,N_2263);
nand U3252 (N_3252,N_2915,N_1040);
or U3253 (N_3253,N_1910,N_432);
xor U3254 (N_3254,In_1474,N_2954);
xor U3255 (N_3255,N_1609,N_1425);
or U3256 (N_3256,N_2972,N_2392);
nand U3257 (N_3257,In_1030,N_2788);
and U3258 (N_3258,N_1686,N_2001);
and U3259 (N_3259,N_1897,N_2537);
xnor U3260 (N_3260,In_25,In_1673);
nand U3261 (N_3261,N_2896,N_2101);
and U3262 (N_3262,In_4423,In_3797);
and U3263 (N_3263,In_603,N_2327);
xor U3264 (N_3264,N_2260,N_2760);
nor U3265 (N_3265,N_2685,N_2698);
nand U3266 (N_3266,N_1955,N_2827);
nand U3267 (N_3267,N_2430,N_1477);
and U3268 (N_3268,N_1687,N_2964);
and U3269 (N_3269,In_176,N_2741);
xnor U3270 (N_3270,N_1455,N_2346);
and U3271 (N_3271,N_1725,N_2301);
nor U3272 (N_3272,In_4786,N_2576);
xnor U3273 (N_3273,N_1235,In_2290);
and U3274 (N_3274,N_2447,N_2835);
or U3275 (N_3275,In_3733,In_618);
or U3276 (N_3276,N_2326,N_2011);
or U3277 (N_3277,N_1284,N_874);
and U3278 (N_3278,In_782,N_2287);
xor U3279 (N_3279,N_2151,N_2626);
or U3280 (N_3280,N_2451,In_3117);
xnor U3281 (N_3281,N_2377,N_2528);
or U3282 (N_3282,In_654,N_2259);
nand U3283 (N_3283,N_2808,N_2015);
and U3284 (N_3284,N_2190,N_2093);
nand U3285 (N_3285,N_2110,N_2280);
or U3286 (N_3286,N_2683,N_2300);
xnor U3287 (N_3287,N_533,N_1030);
and U3288 (N_3288,N_2863,N_2033);
and U3289 (N_3289,N_2008,In_1544);
nand U3290 (N_3290,In_1149,N_2053);
or U3291 (N_3291,N_1891,N_2812);
and U3292 (N_3292,In_4842,N_2235);
xnor U3293 (N_3293,In_4484,N_1370);
or U3294 (N_3294,N_2304,N_2592);
or U3295 (N_3295,N_2205,In_554);
nand U3296 (N_3296,N_826,N_2213);
nor U3297 (N_3297,N_2726,N_2063);
or U3298 (N_3298,In_2653,N_2092);
nor U3299 (N_3299,N_962,In_1112);
or U3300 (N_3300,N_2405,N_1292);
nor U3301 (N_3301,In_3598,N_2173);
xnor U3302 (N_3302,N_1175,N_713);
and U3303 (N_3303,N_2462,N_2947);
and U3304 (N_3304,N_2194,N_1892);
or U3305 (N_3305,N_1311,N_1136);
nor U3306 (N_3306,N_2534,N_2943);
nor U3307 (N_3307,N_829,N_2648);
or U3308 (N_3308,In_85,In_1954);
and U3309 (N_3309,N_2265,In_3532);
or U3310 (N_3310,N_2415,In_697);
nand U3311 (N_3311,N_2570,N_2963);
or U3312 (N_3312,N_2170,In_1105);
nor U3313 (N_3313,N_498,N_2356);
nor U3314 (N_3314,N_2123,In_729);
nor U3315 (N_3315,N_2162,N_1245);
nand U3316 (N_3316,N_2623,N_2495);
nor U3317 (N_3317,In_4404,In_1538);
nor U3318 (N_3318,N_2504,N_2861);
xor U3319 (N_3319,In_1275,In_1774);
or U3320 (N_3320,In_4989,N_2703);
and U3321 (N_3321,N_898,N_2427);
nor U3322 (N_3322,In_818,In_267);
xor U3323 (N_3323,In_907,N_2338);
nand U3324 (N_3324,N_1740,N_2695);
or U3325 (N_3325,N_2128,N_612);
nand U3326 (N_3326,N_2542,N_2376);
or U3327 (N_3327,N_2803,N_2670);
xor U3328 (N_3328,N_2665,N_2594);
xnor U3329 (N_3329,N_2891,N_2119);
or U3330 (N_3330,N_2137,N_1374);
or U3331 (N_3331,N_2207,N_2539);
xnor U3332 (N_3332,N_2874,N_1589);
nor U3333 (N_3333,In_864,N_2970);
and U3334 (N_3334,N_2942,In_3190);
nand U3335 (N_3335,N_2282,In_4098);
xor U3336 (N_3336,In_2723,N_2593);
and U3337 (N_3337,N_2323,N_1931);
xnor U3338 (N_3338,N_1366,N_2669);
and U3339 (N_3339,N_2791,N_1947);
or U3340 (N_3340,N_2035,N_2811);
nor U3341 (N_3341,N_2156,In_236);
or U3342 (N_3342,N_2169,N_2492);
xor U3343 (N_3343,N_2245,N_2054);
xor U3344 (N_3344,In_2805,N_2069);
nand U3345 (N_3345,In_4815,N_2274);
or U3346 (N_3346,N_1033,N_1449);
or U3347 (N_3347,N_1319,In_4105);
xnor U3348 (N_3348,In_4649,N_1368);
xnor U3349 (N_3349,N_1261,N_104);
nor U3350 (N_3350,In_4715,N_2366);
and U3351 (N_3351,In_4299,In_22);
nor U3352 (N_3352,N_2797,In_1700);
and U3353 (N_3353,N_2127,N_1613);
nand U3354 (N_3354,N_2032,N_2832);
nor U3355 (N_3355,N_923,N_2062);
nor U3356 (N_3356,N_2520,N_2955);
or U3357 (N_3357,N_2705,N_2857);
or U3358 (N_3358,N_2556,N_2923);
and U3359 (N_3359,In_1944,N_2877);
nor U3360 (N_3360,N_2095,N_1576);
and U3361 (N_3361,N_2436,N_2439);
nand U3362 (N_3362,N_931,In_3967);
nor U3363 (N_3363,N_1194,In_1702);
xor U3364 (N_3364,In_3472,N_1456);
nor U3365 (N_3365,N_1831,N_1420);
nor U3366 (N_3366,N_1579,N_1149);
or U3367 (N_3367,In_3239,N_2502);
xor U3368 (N_3368,In_1713,N_2279);
xnor U3369 (N_3369,N_1207,In_3903);
xor U3370 (N_3370,In_664,N_2061);
nand U3371 (N_3371,N_928,In_1756);
nand U3372 (N_3372,N_2793,N_2740);
nor U3373 (N_3373,N_1129,N_2386);
nor U3374 (N_3374,N_2087,In_195);
and U3375 (N_3375,N_2355,N_2463);
and U3376 (N_3376,N_2946,N_2024);
and U3377 (N_3377,N_2749,N_2643);
nor U3378 (N_3378,In_394,N_1104);
nand U3379 (N_3379,N_1218,N_2773);
xor U3380 (N_3380,In_2846,In_3422);
nand U3381 (N_3381,In_1818,In_2403);
or U3382 (N_3382,N_1789,In_1486);
or U3383 (N_3383,N_2373,N_2540);
xnor U3384 (N_3384,N_686,N_2501);
and U3385 (N_3385,N_2056,N_2017);
xor U3386 (N_3386,N_2614,N_1531);
nor U3387 (N_3387,N_571,N_2124);
nand U3388 (N_3388,In_2633,N_1474);
xnor U3389 (N_3389,N_2297,N_2046);
nand U3390 (N_3390,N_788,N_2546);
nor U3391 (N_3391,N_1211,In_4063);
or U3392 (N_3392,N_388,In_4885);
and U3393 (N_3393,In_3070,N_2612);
and U3394 (N_3394,In_4282,N_2179);
xnor U3395 (N_3395,N_2299,N_2959);
nand U3396 (N_3396,N_2662,N_2988);
or U3397 (N_3397,N_1475,N_1092);
xnor U3398 (N_3398,In_2665,N_1093);
nand U3399 (N_3399,In_1992,N_1574);
nand U3400 (N_3400,N_2600,N_2351);
nor U3401 (N_3401,N_2701,N_2421);
or U3402 (N_3402,N_2925,In_2915);
or U3403 (N_3403,In_1843,In_4347);
and U3404 (N_3404,In_4930,N_1569);
nand U3405 (N_3405,N_2917,N_1223);
nor U3406 (N_3406,N_1542,In_2354);
xnor U3407 (N_3407,N_2666,N_1648);
or U3408 (N_3408,In_2595,N_2039);
nor U3409 (N_3409,N_2590,N_2633);
nand U3410 (N_3410,N_2473,In_4833);
nor U3411 (N_3411,In_2914,N_2644);
xor U3412 (N_3412,In_4644,N_2807);
or U3413 (N_3413,N_2437,N_2919);
and U3414 (N_3414,N_2362,N_982);
and U3415 (N_3415,In_3734,N_2368);
nand U3416 (N_3416,In_578,N_2731);
and U3417 (N_3417,In_4212,N_2422);
or U3418 (N_3418,In_2937,In_2887);
nor U3419 (N_3419,In_2679,N_2389);
xor U3420 (N_3420,N_1605,N_2185);
xnor U3421 (N_3421,N_2702,N_2859);
nand U3422 (N_3422,In_562,N_2649);
xnor U3423 (N_3423,In_513,N_2029);
nand U3424 (N_3424,In_2400,N_2375);
nand U3425 (N_3425,N_2535,In_3597);
and U3426 (N_3426,N_2706,In_2613);
nand U3427 (N_3427,N_2028,In_3304);
nor U3428 (N_3428,N_1692,N_2712);
nand U3429 (N_3429,N_2247,In_1974);
nor U3430 (N_3430,N_1666,N_719);
nor U3431 (N_3431,N_2659,N_2774);
nor U3432 (N_3432,N_2273,N_2997);
xnor U3433 (N_3433,N_2588,In_2496);
nand U3434 (N_3434,N_2844,In_1082);
or U3435 (N_3435,N_1349,N_2583);
and U3436 (N_3436,N_2998,N_2524);
nand U3437 (N_3437,In_4740,N_2145);
nor U3438 (N_3438,N_2785,N_2990);
xor U3439 (N_3439,N_2975,N_2691);
or U3440 (N_3440,N_2261,N_1644);
nor U3441 (N_3441,N_2553,N_2358);
or U3442 (N_3442,N_2384,N_2686);
nor U3443 (N_3443,In_3947,N_78);
xnor U3444 (N_3444,In_1783,N_2342);
xnor U3445 (N_3445,N_1405,N_1191);
and U3446 (N_3446,In_3403,N_2425);
nand U3447 (N_3447,N_2823,In_2951);
nor U3448 (N_3448,N_2720,N_2503);
nor U3449 (N_3449,N_582,N_2126);
xnor U3450 (N_3450,N_2076,N_2325);
xnor U3451 (N_3451,In_2848,N_2052);
nor U3452 (N_3452,In_2231,N_2238);
nand U3453 (N_3453,N_771,N_2370);
and U3454 (N_3454,N_2926,In_722);
and U3455 (N_3455,N_1131,N_2319);
nand U3456 (N_3456,In_1172,In_2093);
nand U3457 (N_3457,In_4671,In_1004);
nand U3458 (N_3458,N_2305,N_2667);
and U3459 (N_3459,N_2505,In_1272);
and U3460 (N_3460,N_2027,N_2158);
or U3461 (N_3461,In_2006,In_4239);
nor U3462 (N_3462,In_2179,N_2674);
xor U3463 (N_3463,N_2512,N_148);
or U3464 (N_3464,N_219,N_1541);
nor U3465 (N_3465,N_2316,N_2315);
xnor U3466 (N_3466,N_2653,In_4103);
and U3467 (N_3467,N_2440,N_2481);
nand U3468 (N_3468,N_2444,In_1995);
or U3469 (N_3469,N_402,N_2846);
nand U3470 (N_3470,N_959,In_4300);
nand U3471 (N_3471,N_2849,In_1452);
nand U3472 (N_3472,N_1233,In_4620);
and U3473 (N_3473,N_2771,In_3980);
and U3474 (N_3474,N_2945,N_2118);
and U3475 (N_3475,In_132,N_2595);
xnor U3476 (N_3476,N_2777,N_1788);
or U3477 (N_3477,N_1036,N_1297);
and U3478 (N_3478,N_1943,N_2575);
nor U3479 (N_3479,In_4399,N_2515);
nand U3480 (N_3480,In_527,N_1721);
xor U3481 (N_3481,In_2786,N_2637);
nor U3482 (N_3482,N_2584,N_2580);
nand U3483 (N_3483,N_1968,In_4848);
and U3484 (N_3484,N_2937,N_2755);
and U3485 (N_3485,N_2743,N_1777);
nand U3486 (N_3486,N_1169,N_2897);
xor U3487 (N_3487,N_1155,N_2768);
xnor U3488 (N_3488,N_2051,N_2221);
nor U3489 (N_3489,In_795,In_3356);
xor U3490 (N_3490,In_4203,N_2328);
xor U3491 (N_3491,N_2335,N_821);
or U3492 (N_3492,In_1865,N_2693);
or U3493 (N_3493,N_86,N_2025);
or U3494 (N_3494,N_2639,N_2830);
nand U3495 (N_3495,N_1538,N_904);
or U3496 (N_3496,N_1772,In_1986);
nand U3497 (N_3497,In_2563,In_2821);
nand U3498 (N_3498,N_401,N_310);
nand U3499 (N_3499,N_2411,N_2858);
nor U3500 (N_3500,N_2312,N_2995);
xor U3501 (N_3501,In_3442,In_2324);
nand U3502 (N_3502,In_4235,N_2187);
and U3503 (N_3503,In_4081,In_1245);
and U3504 (N_3504,N_1730,N_2388);
nand U3505 (N_3505,N_2228,N_156);
and U3506 (N_3506,N_789,In_3563);
nor U3507 (N_3507,In_4520,N_2317);
nand U3508 (N_3508,N_2625,N_1713);
and U3509 (N_3509,N_2869,N_2875);
xor U3510 (N_3510,N_1808,N_2350);
nor U3511 (N_3511,N_2353,N_2986);
and U3512 (N_3512,N_2470,N_2821);
xnor U3513 (N_3513,N_1727,N_2269);
nand U3514 (N_3514,N_673,N_2241);
nand U3515 (N_3515,N_2498,N_2714);
nor U3516 (N_3516,N_2457,N_2081);
nor U3517 (N_3517,N_2167,In_2978);
or U3518 (N_3518,N_2887,N_2900);
xor U3519 (N_3519,In_4045,N_1317);
nand U3520 (N_3520,N_2313,In_3198);
xor U3521 (N_3521,N_2776,N_2250);
and U3522 (N_3522,N_2817,N_2951);
nand U3523 (N_3523,N_1779,In_3205);
xor U3524 (N_3524,N_48,N_2006);
xor U3525 (N_3525,N_2735,In_3793);
xnor U3526 (N_3526,In_3475,N_2754);
and U3527 (N_3527,N_2890,N_2912);
and U3528 (N_3528,N_2102,N_2761);
and U3529 (N_3529,N_2762,N_2525);
or U3530 (N_3530,N_2333,N_287);
and U3531 (N_3531,N_2216,N_2070);
nand U3532 (N_3532,N_2845,N_1908);
nor U3533 (N_3533,N_2867,N_2860);
nand U3534 (N_3534,N_2883,N_328);
and U3535 (N_3535,N_1471,In_3359);
nand U3536 (N_3536,In_311,N_2778);
or U3537 (N_3537,N_2022,N_2707);
nor U3538 (N_3538,N_588,N_2379);
or U3539 (N_3539,N_2412,N_2013);
or U3540 (N_3540,N_1587,N_2725);
nor U3541 (N_3541,N_242,N_2708);
or U3542 (N_3542,In_1630,N_2852);
nor U3543 (N_3543,N_371,In_454);
nand U3544 (N_3544,N_2507,N_2191);
and U3545 (N_3545,N_160,N_2564);
xnor U3546 (N_3546,N_2222,N_2480);
xor U3547 (N_3547,N_2627,N_113);
xor U3548 (N_3548,N_2406,In_1789);
or U3549 (N_3549,N_2604,N_1606);
or U3550 (N_3550,N_2624,N_2753);
xor U3551 (N_3551,In_4981,N_1059);
and U3552 (N_3552,N_2948,N_1924);
nor U3553 (N_3553,N_1320,N_2862);
nor U3554 (N_3554,N_2608,In_1204);
xor U3555 (N_3555,N_2719,N_2692);
nor U3556 (N_3556,N_2748,N_2973);
nor U3557 (N_3557,N_2700,N_2652);
xor U3558 (N_3558,In_1341,N_2978);
or U3559 (N_3559,In_313,N_1176);
nor U3560 (N_3560,N_2931,In_4941);
or U3561 (N_3561,N_1928,N_2152);
nand U3562 (N_3562,N_638,N_1259);
or U3563 (N_3563,In_4531,N_2042);
nor U3564 (N_3564,N_2286,In_3541);
or U3565 (N_3565,N_2014,N_2483);
nand U3566 (N_3566,N_2086,N_2709);
xor U3567 (N_3567,N_2336,In_3918);
nand U3568 (N_3568,N_1581,N_2906);
nand U3569 (N_3569,N_2730,N_2174);
and U3570 (N_3570,In_2055,In_1964);
and U3571 (N_3571,In_1604,N_2518);
nand U3572 (N_3572,In_1842,In_2796);
nor U3573 (N_3573,N_2395,N_1944);
or U3574 (N_3574,In_4785,In_3151);
or U3575 (N_3575,In_1582,N_2468);
and U3576 (N_3576,N_2486,In_3305);
xnor U3577 (N_3577,In_598,N_2763);
nor U3578 (N_3578,N_2837,N_1711);
and U3579 (N_3579,N_2510,N_617);
xnor U3580 (N_3580,In_3018,In_4847);
nand U3581 (N_3581,N_858,N_2230);
nand U3582 (N_3582,In_1034,N_2204);
and U3583 (N_3583,N_2289,In_577);
and U3584 (N_3584,In_3284,N_2622);
nor U3585 (N_3585,N_2229,N_2854);
or U3586 (N_3586,N_2814,N_2538);
and U3587 (N_3587,N_2723,N_2295);
nor U3588 (N_3588,In_246,N_2872);
nor U3589 (N_3589,N_2678,N_2431);
and U3590 (N_3590,In_1918,N_2910);
nand U3591 (N_3591,N_2303,N_2340);
or U3592 (N_3592,In_2758,N_993);
or U3593 (N_3593,N_2466,N_2239);
and U3594 (N_3594,N_1269,In_4457);
xor U3595 (N_3595,N_2278,N_2097);
nand U3596 (N_3596,In_3580,N_2688);
nor U3597 (N_3597,N_2423,N_1089);
nor U3598 (N_3598,N_1237,N_29);
or U3599 (N_3599,In_2715,N_708);
or U3600 (N_3600,N_1180,In_3729);
xnor U3601 (N_3601,In_2313,N_2950);
nand U3602 (N_3602,N_2453,N_149);
nand U3603 (N_3603,N_2681,N_2888);
and U3604 (N_3604,In_1465,N_2598);
nor U3605 (N_3605,In_4315,N_2140);
nand U3606 (N_3606,N_2272,N_2290);
xor U3607 (N_3607,N_277,N_2378);
and U3608 (N_3608,N_1719,In_1906);
or U3609 (N_3609,N_2582,N_2339);
or U3610 (N_3610,In_3655,N_2668);
nor U3611 (N_3611,N_1447,N_654);
nor U3612 (N_3612,N_809,N_1575);
xor U3613 (N_3613,N_2090,N_2449);
nand U3614 (N_3614,N_2132,N_2751);
and U3615 (N_3615,N_2655,N_2488);
or U3616 (N_3616,N_2789,N_1597);
nand U3617 (N_3617,In_1566,N_1084);
or U3618 (N_3618,N_1863,N_1914);
and U3619 (N_3619,N_2971,In_3110);
xnor U3620 (N_3620,N_2798,N_2306);
xor U3621 (N_3621,N_2450,In_1745);
or U3622 (N_3622,N_2991,N_2884);
nand U3623 (N_3623,N_2294,N_2314);
nand U3624 (N_3624,N_1107,N_2936);
xnor U3625 (N_3625,N_2079,In_1763);
or U3626 (N_3626,N_83,In_2577);
nor U3627 (N_3627,In_1373,N_2838);
nor U3628 (N_3628,N_1518,N_2249);
nand U3629 (N_3629,N_1544,In_3231);
xor U3630 (N_3630,N_2929,N_2382);
xor U3631 (N_3631,In_3910,N_2209);
or U3632 (N_3632,N_1583,N_2125);
or U3633 (N_3633,N_2257,N_2589);
nand U3634 (N_3634,N_542,N_2527);
and U3635 (N_3635,In_3690,N_895);
nor U3636 (N_3636,N_1312,N_2285);
nor U3637 (N_3637,N_2484,N_2049);
nor U3638 (N_3638,In_4129,In_2195);
nor U3639 (N_3639,In_2609,In_1123);
nor U3640 (N_3640,In_4415,N_1359);
xnor U3641 (N_3641,In_2131,N_2246);
or U3642 (N_3642,In_92,In_3558);
xnor U3643 (N_3643,N_1505,In_4285);
nor U3644 (N_3644,N_1400,N_2206);
nand U3645 (N_3645,N_1264,In_1696);
nand U3646 (N_3646,N_2220,N_2645);
xor U3647 (N_3647,N_2920,N_359);
and U3648 (N_3648,N_2255,In_2774);
and U3649 (N_3649,In_2687,In_2536);
nor U3650 (N_3650,N_578,N_127);
and U3651 (N_3651,N_2921,In_2273);
nor U3652 (N_3652,N_2320,N_2672);
or U3653 (N_3653,In_4604,In_3975);
nor U3654 (N_3654,N_293,N_2532);
or U3655 (N_3655,N_2795,In_719);
xnor U3656 (N_3656,N_2968,N_2400);
xor U3657 (N_3657,N_2318,N_2476);
xor U3658 (N_3658,N_2840,N_2736);
and U3659 (N_3659,In_1953,In_1708);
xnor U3660 (N_3660,N_1012,In_3116);
xnor U3661 (N_3661,N_2898,N_2096);
xor U3662 (N_3662,N_2288,N_2341);
or U3663 (N_3663,N_2813,N_2359);
or U3664 (N_3664,In_2198,In_4933);
xor U3665 (N_3665,N_563,N_2816);
xnor U3666 (N_3666,N_2154,N_1932);
and U3667 (N_3667,N_2550,N_2935);
nand U3668 (N_3668,N_2084,N_2497);
or U3669 (N_3669,N_2677,N_2541);
nor U3670 (N_3670,N_1578,N_1570);
or U3671 (N_3671,N_2060,N_1694);
and U3672 (N_3672,N_2080,In_2735);
nor U3673 (N_3673,N_2270,In_2610);
xnor U3674 (N_3674,In_1674,In_2589);
and U3675 (N_3675,N_1600,N_2927);
and U3676 (N_3676,N_2557,N_1397);
or U3677 (N_3677,N_2616,N_2464);
nand U3678 (N_3678,N_2240,N_2938);
xor U3679 (N_3679,N_2974,In_2436);
xor U3680 (N_3680,N_2882,N_2456);
or U3681 (N_3681,N_290,N_2019);
nand U3682 (N_3682,N_2012,In_3606);
xnor U3683 (N_3683,In_4689,In_446);
and U3684 (N_3684,N_2142,N_2587);
nand U3685 (N_3685,N_2914,N_2434);
and U3686 (N_3686,N_1894,N_2208);
nor U3687 (N_3687,N_2969,N_1971);
xor U3688 (N_3688,In_3498,N_1757);
nor U3689 (N_3689,N_1045,N_1624);
or U3690 (N_3690,In_545,N_98);
or U3691 (N_3691,N_2569,N_2508);
or U3692 (N_3692,In_859,N_2275);
or U3693 (N_3693,N_291,N_2548);
xnor U3694 (N_3694,In_4903,In_4024);
and U3695 (N_3695,N_714,N_2810);
nand U3696 (N_3696,N_2212,N_1604);
and U3697 (N_3697,In_3645,In_128);
and U3698 (N_3698,N_2628,N_2585);
and U3699 (N_3699,N_2180,In_283);
nor U3700 (N_3700,N_2104,N_2886);
nand U3701 (N_3701,In_4998,N_2067);
xnor U3702 (N_3702,N_1074,N_2172);
and U3703 (N_3703,N_2638,N_2227);
and U3704 (N_3704,N_2281,N_2308);
nor U3705 (N_3705,N_1158,N_2459);
or U3706 (N_3706,In_390,In_2277);
xor U3707 (N_3707,N_2184,N_2829);
nor U3708 (N_3708,In_511,N_844);
nor U3709 (N_3709,N_2820,In_1124);
or U3710 (N_3710,N_2976,In_1959);
or U3711 (N_3711,N_1564,In_745);
xor U3712 (N_3712,N_2251,N_368);
xor U3713 (N_3713,N_2551,N_2106);
and U3714 (N_3714,N_1677,N_2903);
nand U3715 (N_3715,N_2182,N_2183);
xor U3716 (N_3716,N_2048,N_2545);
xor U3717 (N_3717,N_2802,N_674);
and U3718 (N_3718,In_4486,N_2523);
nor U3719 (N_3719,N_1377,In_4034);
and U3720 (N_3720,In_1167,In_4545);
xor U3721 (N_3721,In_4093,N_2893);
nor U3722 (N_3722,N_2393,N_1285);
nor U3723 (N_3723,N_2148,In_130);
or U3724 (N_3724,N_1465,N_470);
xnor U3725 (N_3725,N_1885,N_2244);
and U3726 (N_3726,N_2020,N_2298);
nor U3727 (N_3727,N_2646,In_3607);
or U3728 (N_3728,N_2609,N_1674);
nor U3729 (N_3729,N_2496,N_2416);
xnor U3730 (N_3730,N_2599,N_2129);
or U3731 (N_3731,In_2506,In_955);
nor U3732 (N_3732,N_2984,In_1243);
nor U3733 (N_3733,N_2980,In_1872);
or U3734 (N_3734,N_1804,In_2869);
nor U3735 (N_3735,N_1137,In_2107);
or U3736 (N_3736,N_1906,N_2996);
nor U3737 (N_3737,In_2000,N_2438);
or U3738 (N_3738,In_3713,N_2680);
and U3739 (N_3739,N_488,N_1776);
and U3740 (N_3740,N_2465,N_2769);
nand U3741 (N_3741,N_2075,N_2454);
nand U3742 (N_3742,N_2420,N_1267);
nand U3743 (N_3743,N_2985,In_1493);
nand U3744 (N_3744,N_2767,N_1794);
nand U3745 (N_3745,N_2347,N_2404);
or U3746 (N_3746,N_2107,In_3081);
and U3747 (N_3747,N_1423,N_2746);
and U3748 (N_3748,N_2752,N_1557);
nand U3749 (N_3749,In_539,N_376);
xor U3750 (N_3750,In_3185,In_3535);
nand U3751 (N_3751,N_1236,N_593);
xor U3752 (N_3752,In_4005,N_2163);
nand U3753 (N_3753,N_129,In_2363);
nor U3754 (N_3754,N_2458,In_1233);
nand U3755 (N_3755,In_2066,N_2911);
xnor U3756 (N_3756,N_2160,N_2800);
nor U3757 (N_3757,N_2579,N_235);
nand U3758 (N_3758,In_3911,N_2682);
xnor U3759 (N_3759,N_2371,N_2630);
nand U3760 (N_3760,N_2784,N_1195);
nor U3761 (N_3761,N_2825,N_527);
or U3762 (N_3762,N_256,N_2258);
nand U3763 (N_3763,N_2122,N_1128);
nor U3764 (N_3764,N_2621,In_1924);
nor U3765 (N_3765,N_1125,N_2099);
and U3766 (N_3766,In_10,N_2586);
and U3767 (N_3767,N_1265,N_1015);
nor U3768 (N_3768,N_2934,In_4374);
and U3769 (N_3769,N_1246,In_1619);
nand U3770 (N_3770,N_1706,N_1881);
and U3771 (N_3771,In_2508,In_35);
xor U3772 (N_3772,In_4483,N_2715);
xnor U3773 (N_3773,N_1747,N_2337);
nand U3774 (N_3774,N_1702,In_2052);
and U3775 (N_3775,N_2141,N_2478);
and U3776 (N_3776,N_532,N_1651);
xor U3777 (N_3777,In_1476,N_2656);
xor U3778 (N_3778,N_2264,N_2536);
xnor U3779 (N_3779,N_448,N_2445);
nand U3780 (N_3780,N_2509,N_2895);
and U3781 (N_3781,N_1391,In_3104);
or U3782 (N_3782,N_2613,N_999);
nor U3783 (N_3783,N_2956,In_4356);
nor U3784 (N_3784,In_4172,In_4997);
nand U3785 (N_3785,In_3308,In_216);
and U3786 (N_3786,N_1226,N_1590);
nor U3787 (N_3787,N_1718,N_2833);
nor U3788 (N_3788,N_2758,N_152);
or U3789 (N_3789,N_2522,N_2433);
nand U3790 (N_3790,N_1759,N_1832);
nor U3791 (N_3791,N_2966,N_330);
or U3792 (N_3792,N_990,N_2226);
nand U3793 (N_3793,N_2782,N_2607);
nor U3794 (N_3794,N_2558,N_2770);
xnor U3795 (N_3795,In_3132,N_2654);
nand U3796 (N_3796,N_946,N_2634);
xnor U3797 (N_3797,In_4352,N_1755);
nand U3798 (N_3798,N_2737,N_2452);
xor U3799 (N_3799,N_2530,N_2999);
xor U3800 (N_3800,In_194,N_2077);
or U3801 (N_3801,In_786,N_917);
or U3802 (N_3802,N_1715,N_2822);
nand U3803 (N_3803,N_2750,N_524);
xor U3804 (N_3804,N_436,In_748);
nand U3805 (N_3805,N_2790,N_2499);
and U3806 (N_3806,N_2203,N_2913);
nor U3807 (N_3807,N_2387,In_1216);
nor U3808 (N_3808,N_2115,In_2905);
xnor U3809 (N_3809,In_4408,N_2435);
xor U3810 (N_3810,N_1307,N_2780);
xnor U3811 (N_3811,N_2930,N_1829);
xor U3812 (N_3812,N_669,In_1802);
and U3813 (N_3813,N_2407,N_801);
nand U3814 (N_3814,N_2002,N_1100);
or U3815 (N_3815,N_2957,N_2010);
nand U3816 (N_3816,In_1307,N_1443);
and U3817 (N_3817,N_2967,In_2604);
nand U3818 (N_3818,N_2529,N_2916);
xor U3819 (N_3819,N_1550,N_2661);
nand U3820 (N_3820,N_1454,N_2992);
xnor U3821 (N_3821,N_168,In_4496);
xnor U3822 (N_3822,In_1597,In_3997);
and U3823 (N_3823,In_2777,In_1718);
or U3824 (N_3824,N_2560,N_431);
nor U3825 (N_3825,N_2603,N_1460);
nor U3826 (N_3826,N_2642,In_4308);
nor U3827 (N_3827,N_2135,In_1072);
xor U3828 (N_3828,N_2819,N_1274);
nor U3829 (N_3829,N_1860,N_1930);
nor U3830 (N_3830,N_224,N_2764);
and U3831 (N_3831,N_2016,In_2487);
nor U3832 (N_3832,N_1975,N_2296);
or U3833 (N_3833,N_2806,N_2219);
nor U3834 (N_3834,N_2253,In_4089);
nor U3835 (N_3835,In_4042,In_2781);
xnor U3836 (N_3836,N_758,N_357);
nand U3837 (N_3837,In_1750,N_2292);
nand U3838 (N_3838,N_2902,N_2979);
nor U3839 (N_3839,N_1923,N_1907);
or U3840 (N_3840,N_1151,N_2675);
xor U3841 (N_3841,N_2805,N_906);
nand U3842 (N_3842,N_2909,N_2493);
nand U3843 (N_3843,N_1006,N_1634);
or U3844 (N_3844,N_2611,N_2694);
nor U3845 (N_3845,In_287,N_2197);
nor U3846 (N_3846,In_434,N_2330);
and U3847 (N_3847,N_1866,N_99);
or U3848 (N_3848,N_1272,In_3494);
xor U3849 (N_3849,In_3182,N_2083);
or U3850 (N_3850,N_1322,N_724);
nor U3851 (N_3851,N_1683,In_387);
xor U3852 (N_3852,N_947,In_4248);
or U3853 (N_3853,N_1991,N_2696);
nand U3854 (N_3854,In_3789,N_2031);
xnor U3855 (N_3855,N_2796,N_1301);
nand U3856 (N_3856,In_1066,N_1482);
nor U3857 (N_3857,In_4541,In_1812);
or U3858 (N_3858,N_2641,N_1279);
nand U3859 (N_3859,N_1830,N_1967);
xnor U3860 (N_3860,N_2113,N_1813);
and U3861 (N_3861,In_1039,In_4181);
or U3862 (N_3862,In_3978,In_2083);
and U3863 (N_3863,N_2742,N_1989);
xor U3864 (N_3864,N_433,N_2799);
nor U3865 (N_3865,N_2787,N_2981);
or U3866 (N_3866,N_1929,N_2547);
nor U3867 (N_3867,N_2690,N_1090);
and U3868 (N_3868,N_1524,N_2322);
or U3869 (N_3869,N_2632,N_228);
and U3870 (N_3870,N_2130,In_3107);
and U3871 (N_3871,N_2153,In_473);
and U3872 (N_3872,N_1332,In_4284);
nand U3873 (N_3873,In_3225,In_656);
xor U3874 (N_3874,N_25,N_2242);
and U3875 (N_3875,N_2074,In_1026);
nor U3876 (N_3876,In_4290,N_1919);
or U3877 (N_3877,N_2460,N_1479);
nor U3878 (N_3878,N_507,N_1573);
nand U3879 (N_3879,N_1428,In_1089);
nor U3880 (N_3880,N_1671,N_2372);
xnor U3881 (N_3881,N_2414,N_1251);
xor U3882 (N_3882,N_1915,N_489);
nand U3883 (N_3883,N_2673,In_4699);
and U3884 (N_3884,N_2461,In_4283);
xnor U3885 (N_3885,N_1327,N_2856);
or U3886 (N_3886,In_3183,N_913);
nand U3887 (N_3887,In_1938,N_2941);
or U3888 (N_3888,N_2596,N_1773);
or U3889 (N_3889,N_1305,In_1533);
xnor U3890 (N_3890,N_1268,N_2424);
nor U3891 (N_3891,In_2760,N_2134);
and U3892 (N_3892,N_2108,In_102);
and U3893 (N_3893,N_2403,N_1489);
and U3894 (N_3894,N_2171,In_4884);
and U3895 (N_3895,In_4803,N_2225);
nor U3896 (N_3896,In_2257,N_2563);
and U3897 (N_3897,In_72,N_2597);
and U3898 (N_3898,N_2442,N_192);
xnor U3899 (N_3899,N_2040,N_722);
and U3900 (N_3900,N_2485,N_1961);
xor U3901 (N_3901,N_2243,N_2037);
and U3902 (N_3902,N_2026,N_2876);
nand U3903 (N_3903,N_1594,N_1954);
or U3904 (N_3904,N_1192,N_85);
or U3905 (N_3905,In_1141,N_1061);
or U3906 (N_3906,In_2158,N_2396);
xnor U3907 (N_3907,N_2068,N_1520);
nor U3908 (N_3908,N_2360,In_2159);
or U3909 (N_3909,N_2713,N_2231);
nor U3910 (N_3910,N_1372,N_2824);
nand U3911 (N_3911,N_2121,N_1527);
xnor U3912 (N_3912,N_2004,N_2901);
or U3913 (N_3913,N_2334,N_2847);
nor U3914 (N_3914,N_721,N_2233);
nand U3915 (N_3915,N_2568,N_1737);
xnor U3916 (N_3916,N_2196,N_2853);
and U3917 (N_3917,In_2022,N_2933);
and U3918 (N_3918,N_2477,In_4523);
or U3919 (N_3919,N_2727,N_2618);
nand U3920 (N_3920,N_2804,N_1533);
or U3921 (N_3921,N_184,N_2554);
xor U3922 (N_3922,N_536,In_1622);
or U3923 (N_3923,N_2831,N_2188);
nand U3924 (N_3924,N_2443,N_2237);
or U3925 (N_3925,N_2636,In_3538);
xnor U3926 (N_3926,N_2164,In_1093);
and U3927 (N_3927,In_4927,N_1286);
nor U3928 (N_3928,N_2873,N_2922);
or U3929 (N_3929,N_2331,N_2103);
xor U3930 (N_3930,N_2899,In_792);
xnor U3931 (N_3931,N_2311,N_2994);
nor U3932 (N_3932,N_2165,N_2198);
and U3933 (N_3933,N_2561,N_2489);
or U3934 (N_3934,N_417,N_2419);
nand U3935 (N_3935,N_2940,N_1057);
xnor U3936 (N_3936,N_1890,In_3397);
nand U3937 (N_3937,N_2365,N_2839);
or U3938 (N_3938,N_2005,N_2363);
and U3939 (N_3939,N_1710,N_2671);
nor U3940 (N_3940,In_112,N_2908);
or U3941 (N_3941,N_1294,N_2064);
nor U3942 (N_3942,N_2834,In_3164);
or U3943 (N_3943,N_2962,In_4082);
nor U3944 (N_3944,N_2960,N_1974);
and U3945 (N_3945,N_2549,N_2759);
nor U3946 (N_3946,In_4256,N_2256);
nor U3947 (N_3947,N_2391,N_2023);
nor U3948 (N_3948,N_2417,In_1502);
xnor U3949 (N_3949,N_2880,N_342);
nand U3950 (N_3950,N_1350,N_2131);
nand U3951 (N_3951,N_2739,In_2845);
or U3952 (N_3952,N_1833,In_4450);
xor U3953 (N_3953,N_2268,N_255);
nor U3954 (N_3954,In_2530,N_2765);
nor U3955 (N_3955,N_2952,In_4148);
nand U3956 (N_3956,N_2689,N_1182);
or U3957 (N_3957,N_2367,N_2619);
or U3958 (N_3958,N_1523,N_2526);
xnor U3959 (N_3959,N_2390,In_2353);
and U3960 (N_3960,N_1595,N_491);
xnor U3961 (N_3961,In_3001,N_2000);
nor U3962 (N_3962,N_2277,N_1614);
and U3963 (N_3963,N_63,N_1749);
or U3964 (N_3964,N_1054,In_4055);
or U3965 (N_3965,N_2855,In_3368);
and U3966 (N_3966,N_1979,N_1419);
nor U3967 (N_3967,N_2186,N_2989);
nor U3968 (N_3968,N_2738,N_2428);
and U3969 (N_3969,N_1560,In_257);
nor U3970 (N_3970,N_2446,N_1257);
or U3971 (N_3971,In_2318,N_1088);
or U3972 (N_3972,N_2475,N_1348);
or U3973 (N_3973,In_2963,N_1982);
xnor U3974 (N_3974,N_2426,N_1983);
nor U3975 (N_3975,N_2007,N_2710);
nand U3976 (N_3976,N_2058,In_3071);
or U3977 (N_3977,N_2349,N_2166);
and U3978 (N_3978,N_539,In_901);
xor U3979 (N_3979,N_2794,N_2724);
nand U3980 (N_3980,N_2397,N_2201);
or U3981 (N_3981,In_3363,N_2175);
nand U3982 (N_3982,N_2939,In_4988);
nor U3983 (N_3983,N_2149,In_739);
nor U3984 (N_3984,N_886,N_1487);
nor U3985 (N_3985,In_918,N_2982);
nor U3986 (N_3986,In_401,In_2879);
or U3987 (N_3987,N_2098,N_2766);
nand U3988 (N_3988,N_1174,N_979);
nand U3989 (N_3989,N_2380,N_1682);
xnor U3990 (N_3990,In_1327,N_1309);
xnor U3991 (N_3991,N_864,In_3970);
xor U3992 (N_3992,N_2841,N_2343);
nor U3993 (N_3993,N_2533,N_2562);
nand U3994 (N_3994,In_978,N_1042);
nor U3995 (N_3995,N_1790,N_2573);
nor U3996 (N_3996,N_2756,N_335);
nor U3997 (N_3997,In_2587,N_2905);
nor U3998 (N_3998,N_124,N_2041);
nand U3999 (N_3999,N_2531,N_2650);
xnor U4000 (N_4000,N_3897,N_3376);
xor U4001 (N_4001,N_3605,N_3824);
or U4002 (N_4002,N_3227,N_3805);
or U4003 (N_4003,N_3513,N_3670);
and U4004 (N_4004,N_3747,N_3398);
nor U4005 (N_4005,N_3384,N_3644);
and U4006 (N_4006,N_3952,N_3516);
or U4007 (N_4007,N_3000,N_3892);
xor U4008 (N_4008,N_3649,N_3068);
nor U4009 (N_4009,N_3962,N_3258);
nor U4010 (N_4010,N_3333,N_3680);
xnor U4011 (N_4011,N_3428,N_3083);
nand U4012 (N_4012,N_3861,N_3691);
xor U4013 (N_4013,N_3566,N_3880);
xor U4014 (N_4014,N_3731,N_3545);
nor U4015 (N_4015,N_3431,N_3441);
xnor U4016 (N_4016,N_3915,N_3445);
or U4017 (N_4017,N_3647,N_3882);
nor U4018 (N_4018,N_3130,N_3623);
and U4019 (N_4019,N_3865,N_3180);
and U4020 (N_4020,N_3923,N_3251);
nand U4021 (N_4021,N_3341,N_3032);
nand U4022 (N_4022,N_3521,N_3507);
or U4023 (N_4023,N_3075,N_3693);
nand U4024 (N_4024,N_3673,N_3813);
xor U4025 (N_4025,N_3448,N_3451);
and U4026 (N_4026,N_3781,N_3095);
xnor U4027 (N_4027,N_3348,N_3728);
nand U4028 (N_4028,N_3264,N_3675);
nor U4029 (N_4029,N_3209,N_3662);
or U4030 (N_4030,N_3734,N_3161);
or U4031 (N_4031,N_3113,N_3655);
nor U4032 (N_4032,N_3912,N_3479);
and U4033 (N_4033,N_3919,N_3529);
xnor U4034 (N_4034,N_3242,N_3198);
nand U4035 (N_4035,N_3235,N_3754);
xor U4036 (N_4036,N_3014,N_3374);
nor U4037 (N_4037,N_3855,N_3640);
nand U4038 (N_4038,N_3031,N_3353);
nor U4039 (N_4039,N_3920,N_3648);
nand U4040 (N_4040,N_3142,N_3186);
or U4041 (N_4041,N_3932,N_3899);
nand U4042 (N_4042,N_3409,N_3695);
nand U4043 (N_4043,N_3045,N_3148);
nand U4044 (N_4044,N_3558,N_3913);
or U4045 (N_4045,N_3028,N_3766);
xor U4046 (N_4046,N_3056,N_3346);
and U4047 (N_4047,N_3723,N_3534);
nand U4048 (N_4048,N_3547,N_3034);
and U4049 (N_4049,N_3669,N_3291);
or U4050 (N_4050,N_3540,N_3707);
or U4051 (N_4051,N_3119,N_3790);
nor U4052 (N_4052,N_3578,N_3711);
or U4053 (N_4053,N_3159,N_3854);
nor U4054 (N_4054,N_3385,N_3511);
xor U4055 (N_4055,N_3473,N_3342);
or U4056 (N_4056,N_3732,N_3332);
nor U4057 (N_4057,N_3335,N_3817);
nand U4058 (N_4058,N_3340,N_3576);
or U4059 (N_4059,N_3922,N_3461);
nand U4060 (N_4060,N_3350,N_3443);
nand U4061 (N_4061,N_3415,N_3009);
and U4062 (N_4062,N_3188,N_3630);
or U4063 (N_4063,N_3959,N_3049);
nor U4064 (N_4064,N_3979,N_3453);
xnor U4065 (N_4065,N_3042,N_3424);
or U4066 (N_4066,N_3081,N_3687);
nand U4067 (N_4067,N_3846,N_3624);
nand U4068 (N_4068,N_3307,N_3986);
and U4069 (N_4069,N_3877,N_3671);
or U4070 (N_4070,N_3069,N_3071);
nor U4071 (N_4071,N_3229,N_3543);
nor U4072 (N_4072,N_3779,N_3908);
nand U4073 (N_4073,N_3950,N_3668);
or U4074 (N_4074,N_3109,N_3862);
or U4075 (N_4075,N_3809,N_3129);
xor U4076 (N_4076,N_3970,N_3285);
nor U4077 (N_4077,N_3536,N_3866);
nand U4078 (N_4078,N_3017,N_3914);
xor U4079 (N_4079,N_3555,N_3764);
and U4080 (N_4080,N_3606,N_3399);
nand U4081 (N_4081,N_3482,N_3631);
and U4082 (N_4082,N_3506,N_3568);
nor U4083 (N_4083,N_3514,N_3462);
or U4084 (N_4084,N_3369,N_3167);
and U4085 (N_4085,N_3104,N_3894);
nand U4086 (N_4086,N_3233,N_3515);
or U4087 (N_4087,N_3084,N_3173);
and U4088 (N_4088,N_3370,N_3678);
and U4089 (N_4089,N_3190,N_3783);
nor U4090 (N_4090,N_3921,N_3757);
nand U4091 (N_4091,N_3613,N_3300);
or U4092 (N_4092,N_3019,N_3214);
xor U4093 (N_4093,N_3442,N_3978);
nor U4094 (N_4094,N_3013,N_3393);
xor U4095 (N_4095,N_3849,N_3725);
nand U4096 (N_4096,N_3663,N_3860);
or U4097 (N_4097,N_3610,N_3192);
xnor U4098 (N_4098,N_3364,N_3604);
or U4099 (N_4099,N_3762,N_3697);
nor U4100 (N_4100,N_3412,N_3903);
and U4101 (N_4101,N_3588,N_3288);
and U4102 (N_4102,N_3859,N_3268);
or U4103 (N_4103,N_3259,N_3756);
or U4104 (N_4104,N_3904,N_3868);
nand U4105 (N_4105,N_3886,N_3015);
nand U4106 (N_4106,N_3008,N_3537);
or U4107 (N_4107,N_3270,N_3347);
nand U4108 (N_4108,N_3174,N_3121);
nand U4109 (N_4109,N_3949,N_3947);
xnor U4110 (N_4110,N_3772,N_3218);
and U4111 (N_4111,N_3800,N_3468);
and U4112 (N_4112,N_3497,N_3061);
or U4113 (N_4113,N_3330,N_3775);
xnor U4114 (N_4114,N_3591,N_3256);
nor U4115 (N_4115,N_3826,N_3211);
nor U4116 (N_4116,N_3967,N_3538);
nor U4117 (N_4117,N_3394,N_3659);
xnor U4118 (N_4118,N_3802,N_3417);
xor U4119 (N_4119,N_3444,N_3698);
and U4120 (N_4120,N_3753,N_3222);
or U4121 (N_4121,N_3564,N_3688);
xnor U4122 (N_4122,N_3151,N_3498);
and U4123 (N_4123,N_3717,N_3684);
or U4124 (N_4124,N_3063,N_3987);
nor U4125 (N_4125,N_3406,N_3694);
or U4126 (N_4126,N_3664,N_3359);
nand U4127 (N_4127,N_3377,N_3204);
and U4128 (N_4128,N_3484,N_3027);
xnor U4129 (N_4129,N_3542,N_3819);
and U4130 (N_4130,N_3951,N_3085);
xnor U4131 (N_4131,N_3556,N_3585);
and U4132 (N_4132,N_3147,N_3351);
nor U4133 (N_4133,N_3653,N_3677);
nand U4134 (N_4134,N_3365,N_3867);
nand U4135 (N_4135,N_3279,N_3579);
xor U4136 (N_4136,N_3101,N_3029);
or U4137 (N_4137,N_3257,N_3743);
nand U4138 (N_4138,N_3767,N_3210);
nor U4139 (N_4139,N_3102,N_3569);
xor U4140 (N_4140,N_3665,N_3349);
xor U4141 (N_4141,N_3617,N_3789);
and U4142 (N_4142,N_3927,N_3311);
and U4143 (N_4143,N_3980,N_3744);
nor U4144 (N_4144,N_3567,N_3785);
nor U4145 (N_4145,N_3072,N_3713);
xnor U4146 (N_4146,N_3219,N_3963);
nand U4147 (N_4147,N_3007,N_3395);
xor U4148 (N_4148,N_3895,N_3132);
xnor U4149 (N_4149,N_3776,N_3038);
or U4150 (N_4150,N_3551,N_3459);
nand U4151 (N_4151,N_3845,N_3625);
xor U4152 (N_4152,N_3360,N_3638);
or U4153 (N_4153,N_3768,N_3493);
xnor U4154 (N_4154,N_3690,N_3306);
nand U4155 (N_4155,N_3936,N_3244);
nand U4156 (N_4156,N_3124,N_3089);
and U4157 (N_4157,N_3114,N_3305);
nor U4158 (N_4158,N_3831,N_3413);
xor U4159 (N_4159,N_3116,N_3607);
and U4160 (N_4160,N_3082,N_3989);
or U4161 (N_4161,N_3729,N_3530);
xor U4162 (N_4162,N_3247,N_3060);
xnor U4163 (N_4163,N_3463,N_3942);
nor U4164 (N_4164,N_3149,N_3006);
and U4165 (N_4165,N_3573,N_3505);
nand U4166 (N_4166,N_3517,N_3965);
nor U4167 (N_4167,N_3988,N_3944);
or U4168 (N_4168,N_3423,N_3961);
nor U4169 (N_4169,N_3703,N_3827);
and U4170 (N_4170,N_3881,N_3025);
xnor U4171 (N_4171,N_3383,N_3889);
or U4172 (N_4172,N_3336,N_3667);
xnor U4173 (N_4173,N_3076,N_3487);
nand U4174 (N_4174,N_3784,N_3269);
xor U4175 (N_4175,N_3111,N_3548);
nor U4176 (N_4176,N_3199,N_3616);
xnor U4177 (N_4177,N_3798,N_3217);
nor U4178 (N_4178,N_3329,N_3091);
nand U4179 (N_4179,N_3315,N_3324);
and U4180 (N_4180,N_3751,N_3197);
or U4181 (N_4181,N_3552,N_3420);
or U4182 (N_4182,N_3641,N_3887);
and U4183 (N_4183,N_3930,N_3917);
nand U4184 (N_4184,N_3078,N_3208);
nor U4185 (N_4185,N_3550,N_3512);
and U4186 (N_4186,N_3740,N_3157);
xor U4187 (N_4187,N_3561,N_3293);
nor U4188 (N_4188,N_3041,N_3367);
xor U4189 (N_4189,N_3096,N_3544);
and U4190 (N_4190,N_3267,N_3163);
nor U4191 (N_4191,N_3454,N_3411);
or U4192 (N_4192,N_3297,N_3658);
nor U4193 (N_4193,N_3502,N_3274);
nand U4194 (N_4194,N_3175,N_3736);
nor U4195 (N_4195,N_3144,N_3654);
nand U4196 (N_4196,N_3595,N_3287);
or U4197 (N_4197,N_3488,N_3381);
xnor U4198 (N_4198,N_3918,N_3262);
or U4199 (N_4199,N_3464,N_3977);
and U4200 (N_4200,N_3925,N_3309);
and U4201 (N_4201,N_3371,N_3749);
nor U4202 (N_4202,N_3005,N_3997);
nor U4203 (N_4203,N_3250,N_3522);
or U4204 (N_4204,N_3905,N_3489);
nand U4205 (N_4205,N_3098,N_3964);
nand U4206 (N_4206,N_3929,N_3574);
nand U4207 (N_4207,N_3539,N_3765);
and U4208 (N_4208,N_3177,N_3325);
nor U4209 (N_4209,N_3651,N_3194);
and U4210 (N_4210,N_3856,N_3946);
nor U4211 (N_4211,N_3998,N_3793);
xnor U4212 (N_4212,N_3822,N_3686);
or U4213 (N_4213,N_3470,N_3079);
nor U4214 (N_4214,N_3065,N_3777);
and U4215 (N_4215,N_3265,N_3490);
and U4216 (N_4216,N_3883,N_3236);
xnor U4217 (N_4217,N_3338,N_3145);
or U4218 (N_4218,N_3436,N_3853);
or U4219 (N_4219,N_3873,N_3788);
nand U4220 (N_4220,N_3750,N_3266);
nand U4221 (N_4221,N_3408,N_3002);
or U4222 (N_4222,N_3597,N_3879);
and U4223 (N_4223,N_3053,N_3248);
xnor U4224 (N_4224,N_3193,N_3165);
nand U4225 (N_4225,N_3278,N_3143);
nor U4226 (N_4226,N_3601,N_3589);
or U4227 (N_4227,N_3317,N_3123);
xor U4228 (N_4228,N_3639,N_3852);
or U4229 (N_4229,N_3618,N_3742);
or U4230 (N_4230,N_3692,N_3869);
or U4231 (N_4231,N_3480,N_3221);
or U4232 (N_4232,N_3292,N_3811);
or U4233 (N_4233,N_3991,N_3410);
nor U4234 (N_4234,N_3456,N_3559);
nand U4235 (N_4235,N_3902,N_3621);
or U4236 (N_4236,N_3724,N_3020);
nand U4237 (N_4237,N_3135,N_3632);
nor U4238 (N_4238,N_3202,N_3941);
nand U4239 (N_4239,N_3948,N_3253);
nor U4240 (N_4240,N_3619,N_3823);
xor U4241 (N_4241,N_3689,N_3587);
and U4242 (N_4242,N_3429,N_3926);
nand U4243 (N_4243,N_3628,N_3246);
nor U4244 (N_4244,N_3495,N_3735);
or U4245 (N_4245,N_3382,N_3093);
xor U4246 (N_4246,N_3094,N_3825);
and U4247 (N_4247,N_3366,N_3508);
xor U4248 (N_4248,N_3160,N_3661);
or U4249 (N_4249,N_3276,N_3769);
or U4250 (N_4250,N_3755,N_3973);
and U4251 (N_4251,N_3531,N_3074);
or U4252 (N_4252,N_3387,N_3086);
nor U4253 (N_4253,N_3633,N_3252);
nand U4254 (N_4254,N_3206,N_3581);
and U4255 (N_4255,N_3620,N_3791);
nor U4256 (N_4256,N_3810,N_3844);
or U4257 (N_4257,N_3018,N_3611);
nor U4258 (N_4258,N_3491,N_3334);
nand U4259 (N_4259,N_3636,N_3216);
or U4260 (N_4260,N_3720,N_3666);
or U4261 (N_4261,N_3310,N_3139);
or U4262 (N_4262,N_3565,N_3705);
and U4263 (N_4263,N_3935,N_3437);
xor U4264 (N_4264,N_3048,N_3239);
and U4265 (N_4265,N_3737,N_3909);
nand U4266 (N_4266,N_3830,N_3916);
and U4267 (N_4267,N_3739,N_3541);
nor U4268 (N_4268,N_3281,N_3483);
nand U4269 (N_4269,N_3652,N_3820);
and U4270 (N_4270,N_3594,N_3660);
nor U4271 (N_4271,N_3176,N_3115);
and U4272 (N_4272,N_3771,N_3834);
nand U4273 (N_4273,N_3730,N_3504);
nor U4274 (N_4274,N_3486,N_3363);
xor U4275 (N_4275,N_3200,N_3319);
nand U4276 (N_4276,N_3389,N_3064);
xor U4277 (N_4277,N_3168,N_3808);
nand U4278 (N_4278,N_3302,N_3450);
xnor U4279 (N_4279,N_3748,N_3575);
and U4280 (N_4280,N_3476,N_3314);
xnor U4281 (N_4281,N_3975,N_3183);
nand U4282 (N_4282,N_3375,N_3833);
xnor U4283 (N_4283,N_3699,N_3937);
xnor U4284 (N_4284,N_3294,N_3232);
nor U4285 (N_4285,N_3125,N_3758);
and U4286 (N_4286,N_3608,N_3780);
nand U4287 (N_4287,N_3458,N_3153);
xor U4288 (N_4288,N_3501,N_3321);
or U4289 (N_4289,N_3738,N_3847);
nand U4290 (N_4290,N_3931,N_3156);
nand U4291 (N_4291,N_3296,N_3993);
or U4292 (N_4292,N_3596,N_3172);
and U4293 (N_4293,N_3804,N_3234);
nor U4294 (N_4294,N_3299,N_3642);
xnor U4295 (N_4295,N_3354,N_3137);
or U4296 (N_4296,N_3710,N_3843);
and U4297 (N_4297,N_3577,N_3763);
or U4298 (N_4298,N_3622,N_3572);
xnor U4299 (N_4299,N_3220,N_3794);
nand U4300 (N_4300,N_3796,N_3295);
xnor U4301 (N_4301,N_3405,N_3599);
or U4302 (N_4302,N_3418,N_3471);
or U4303 (N_4303,N_3958,N_3178);
and U4304 (N_4304,N_3774,N_3841);
xor U4305 (N_4305,N_3685,N_3391);
or U4306 (N_4306,N_3870,N_3414);
nor U4307 (N_4307,N_3896,N_3968);
and U4308 (N_4308,N_3526,N_3519);
nor U4309 (N_4309,N_3182,N_3778);
nand U4310 (N_4310,N_3672,N_3815);
xnor U4311 (N_4311,N_3535,N_3612);
nand U4312 (N_4312,N_3906,N_3679);
and U4313 (N_4313,N_3615,N_3901);
nor U4314 (N_4314,N_3888,N_3996);
or U4315 (N_4315,N_3924,N_3277);
or U4316 (N_4316,N_3205,N_3650);
or U4317 (N_4317,N_3590,N_3657);
nand U4318 (N_4318,N_3226,N_3390);
and U4319 (N_4319,N_3228,N_3910);
or U4320 (N_4320,N_3890,N_3432);
and U4321 (N_4321,N_3477,N_3171);
nand U4322 (N_4322,N_3062,N_3240);
nor U4323 (N_4323,N_3331,N_3801);
or U4324 (N_4324,N_3362,N_3080);
xor U4325 (N_4325,N_3733,N_3503);
or U4326 (N_4326,N_3701,N_3828);
or U4327 (N_4327,N_3752,N_3003);
xnor U4328 (N_4328,N_3447,N_3110);
nor U4329 (N_4329,N_3582,N_3245);
nand U4330 (N_4330,N_3864,N_3478);
or U4331 (N_4331,N_3718,N_3598);
nor U4332 (N_4332,N_3054,N_3138);
or U4333 (N_4333,N_3273,N_3803);
xnor U4334 (N_4334,N_3033,N_3485);
or U4335 (N_4335,N_3982,N_3092);
xnor U4336 (N_4336,N_3907,N_3626);
and U4337 (N_4337,N_3055,N_3357);
xor U4338 (N_4338,N_3583,N_3380);
nor U4339 (N_4339,N_3593,N_3643);
and U4340 (N_4340,N_3704,N_3396);
xor U4341 (N_4341,N_3806,N_3133);
nor U4342 (N_4342,N_3945,N_3320);
or U4343 (N_4343,N_3821,N_3051);
and U4344 (N_4344,N_3057,N_3702);
xor U4345 (N_4345,N_3795,N_3313);
or U4346 (N_4346,N_3120,N_3570);
xor U4347 (N_4347,N_3955,N_3301);
xnor U4348 (N_4348,N_3837,N_3105);
nor U4349 (N_4349,N_3836,N_3759);
nand U4350 (N_4350,N_3106,N_3397);
nor U4351 (N_4351,N_3434,N_3990);
and U4352 (N_4352,N_3339,N_3134);
and U4353 (N_4353,N_3494,N_3683);
nand U4354 (N_4354,N_3603,N_3184);
nand U4355 (N_4355,N_3358,N_3255);
nor U4356 (N_4356,N_3560,N_3510);
nor U4357 (N_4357,N_3580,N_3562);
xor U4358 (N_4358,N_3934,N_3289);
nor U4359 (N_4359,N_3549,N_3635);
and U4360 (N_4360,N_3885,N_3634);
nand U4361 (N_4361,N_3323,N_3225);
nand U4362 (N_4362,N_3928,N_3981);
nor U4363 (N_4363,N_3893,N_3356);
and U4364 (N_4364,N_3940,N_3345);
and U4365 (N_4365,N_3097,N_3656);
nand U4366 (N_4366,N_3263,N_3976);
or U4367 (N_4367,N_3337,N_3213);
or U4368 (N_4368,N_3999,N_3716);
xor U4369 (N_4369,N_3994,N_3322);
xor U4370 (N_4370,N_3419,N_3047);
and U4371 (N_4371,N_3352,N_3911);
xor U4372 (N_4372,N_3343,N_3773);
nor U4373 (N_4373,N_3088,N_3146);
or U4374 (N_4374,N_3816,N_3674);
nor U4375 (N_4375,N_3974,N_3191);
nor U4376 (N_4376,N_3303,N_3770);
and U4377 (N_4377,N_3455,N_3373);
and U4378 (N_4378,N_3223,N_3957);
xor U4379 (N_4379,N_3117,N_3392);
and U4380 (N_4380,N_3851,N_3022);
or U4381 (N_4381,N_3282,N_3812);
xnor U4382 (N_4382,N_3466,N_3077);
nand U4383 (N_4383,N_3004,N_3835);
xnor U4384 (N_4384,N_3741,N_3637);
or U4385 (N_4385,N_3469,N_3884);
nand U4386 (N_4386,N_3457,N_3761);
and U4387 (N_4387,N_3304,N_3971);
or U4388 (N_4388,N_3708,N_3969);
nor U4389 (N_4389,N_3440,N_3107);
nor U4390 (N_4390,N_3563,N_3727);
xnor U4391 (N_4391,N_3528,N_3839);
or U4392 (N_4392,N_3722,N_3162);
nand U4393 (N_4393,N_3475,N_3433);
xor U4394 (N_4394,N_3953,N_3682);
or U4395 (N_4395,N_3308,N_3011);
nor U4396 (N_4396,N_3627,N_3966);
nand U4397 (N_4397,N_3103,N_3372);
and U4398 (N_4398,N_3271,N_3439);
nand U4399 (N_4399,N_3992,N_3553);
xnor U4400 (N_4400,N_3318,N_3001);
xnor U4401 (N_4401,N_3158,N_3379);
xor U4402 (N_4402,N_3070,N_3629);
nor U4403 (N_4403,N_3016,N_3243);
or U4404 (N_4404,N_3166,N_3136);
xnor U4405 (N_4405,N_3430,N_3189);
xor U4406 (N_4406,N_3407,N_3141);
nand U4407 (N_4407,N_3943,N_3995);
nor U4408 (N_4408,N_3681,N_3024);
or U4409 (N_4409,N_3985,N_3212);
nand U4410 (N_4410,N_3298,N_3118);
xnor U4411 (N_4411,N_3712,N_3355);
nor U4412 (N_4412,N_3122,N_3388);
xor U4413 (N_4413,N_3933,N_3196);
nor U4414 (N_4414,N_3275,N_3878);
and U4415 (N_4415,N_3714,N_3496);
or U4416 (N_4416,N_3128,N_3787);
or U4417 (N_4417,N_3452,N_3066);
nor U4418 (N_4418,N_3972,N_3090);
and U4419 (N_4419,N_3052,N_3900);
and U4420 (N_4420,N_3438,N_3422);
nor U4421 (N_4421,N_3792,N_3261);
or U4422 (N_4422,N_3280,N_3421);
nor U4423 (N_4423,N_3181,N_3040);
nor U4424 (N_4424,N_3012,N_3797);
xnor U4425 (N_4425,N_3249,N_3401);
nand U4426 (N_4426,N_3035,N_3956);
xnor U4427 (N_4427,N_3818,N_3368);
xor U4428 (N_4428,N_3832,N_3215);
or U4429 (N_4429,N_3044,N_3546);
and U4430 (N_4430,N_3312,N_3073);
nand U4431 (N_4431,N_3155,N_3284);
and U4432 (N_4432,N_3316,N_3154);
or U4433 (N_4433,N_3021,N_3030);
nor U4434 (N_4434,N_3416,N_3446);
or U4435 (N_4435,N_3023,N_3840);
nor U4436 (N_4436,N_3960,N_3760);
xor U4437 (N_4437,N_3164,N_3509);
or U4438 (N_4438,N_3518,N_3614);
nor U4439 (N_4439,N_3492,N_3286);
xnor U4440 (N_4440,N_3571,N_3525);
and U4441 (N_4441,N_3726,N_3706);
nor U4442 (N_4442,N_3326,N_3745);
or U4443 (N_4443,N_3108,N_3829);
and U4444 (N_4444,N_3059,N_3481);
or U4445 (N_4445,N_3696,N_3983);
and U4446 (N_4446,N_3426,N_3876);
nand U4447 (N_4447,N_3241,N_3602);
and U4448 (N_4448,N_3891,N_3592);
xor U4449 (N_4449,N_3523,N_3327);
nor U4450 (N_4450,N_3386,N_3533);
or U4451 (N_4451,N_3043,N_3100);
or U4452 (N_4452,N_3554,N_3584);
nor U4453 (N_4453,N_3609,N_3425);
nor U4454 (N_4454,N_3067,N_3871);
nor U4455 (N_4455,N_3254,N_3520);
or U4456 (N_4456,N_3874,N_3195);
or U4457 (N_4457,N_3046,N_3848);
xnor U4458 (N_4458,N_3524,N_3715);
and U4459 (N_4459,N_3039,N_3719);
nor U4460 (N_4460,N_3050,N_3058);
or U4461 (N_4461,N_3814,N_3170);
nor U4462 (N_4462,N_3203,N_3857);
nor U4463 (N_4463,N_3676,N_3435);
and U4464 (N_4464,N_3272,N_3449);
and U4465 (N_4465,N_3150,N_3231);
or U4466 (N_4466,N_3169,N_3127);
xor U4467 (N_4467,N_3875,N_3037);
nand U4468 (N_4468,N_3087,N_3600);
nand U4469 (N_4469,N_3131,N_3586);
and U4470 (N_4470,N_3984,N_3026);
nor U4471 (N_4471,N_3799,N_3427);
or U4472 (N_4472,N_3344,N_3152);
nor U4473 (N_4473,N_3838,N_3179);
xor U4474 (N_4474,N_3201,N_3230);
or U4475 (N_4475,N_3260,N_3404);
nor U4476 (N_4476,N_3112,N_3746);
nand U4477 (N_4477,N_3207,N_3782);
nor U4478 (N_4478,N_3187,N_3010);
nand U4479 (N_4479,N_3185,N_3472);
xor U4480 (N_4480,N_3238,N_3140);
nand U4481 (N_4481,N_3499,N_3872);
nand U4482 (N_4482,N_3467,N_3858);
or U4483 (N_4483,N_3842,N_3527);
nor U4484 (N_4484,N_3402,N_3939);
xor U4485 (N_4485,N_3646,N_3709);
or U4486 (N_4486,N_3361,N_3460);
nand U4487 (N_4487,N_3099,N_3378);
or U4488 (N_4488,N_3237,N_3938);
and U4489 (N_4489,N_3954,N_3898);
or U4490 (N_4490,N_3532,N_3290);
or U4491 (N_4491,N_3400,N_3786);
xnor U4492 (N_4492,N_3283,N_3465);
xnor U4493 (N_4493,N_3850,N_3807);
nand U4494 (N_4494,N_3557,N_3863);
nand U4495 (N_4495,N_3645,N_3224);
or U4496 (N_4496,N_3403,N_3700);
and U4497 (N_4497,N_3328,N_3721);
and U4498 (N_4498,N_3126,N_3036);
or U4499 (N_4499,N_3500,N_3474);
nor U4500 (N_4500,N_3542,N_3545);
or U4501 (N_4501,N_3356,N_3905);
nand U4502 (N_4502,N_3009,N_3238);
nand U4503 (N_4503,N_3366,N_3505);
and U4504 (N_4504,N_3708,N_3909);
nor U4505 (N_4505,N_3009,N_3062);
or U4506 (N_4506,N_3392,N_3175);
or U4507 (N_4507,N_3613,N_3390);
and U4508 (N_4508,N_3842,N_3914);
nand U4509 (N_4509,N_3754,N_3671);
nand U4510 (N_4510,N_3655,N_3983);
nand U4511 (N_4511,N_3008,N_3645);
nor U4512 (N_4512,N_3984,N_3657);
or U4513 (N_4513,N_3072,N_3688);
or U4514 (N_4514,N_3838,N_3233);
and U4515 (N_4515,N_3029,N_3777);
xor U4516 (N_4516,N_3685,N_3482);
and U4517 (N_4517,N_3718,N_3094);
nor U4518 (N_4518,N_3197,N_3707);
nor U4519 (N_4519,N_3831,N_3276);
and U4520 (N_4520,N_3401,N_3449);
and U4521 (N_4521,N_3499,N_3704);
and U4522 (N_4522,N_3002,N_3702);
nand U4523 (N_4523,N_3168,N_3507);
and U4524 (N_4524,N_3025,N_3766);
or U4525 (N_4525,N_3027,N_3323);
xor U4526 (N_4526,N_3667,N_3069);
xnor U4527 (N_4527,N_3362,N_3874);
and U4528 (N_4528,N_3254,N_3301);
or U4529 (N_4529,N_3500,N_3432);
or U4530 (N_4530,N_3508,N_3494);
and U4531 (N_4531,N_3268,N_3470);
nand U4532 (N_4532,N_3528,N_3412);
or U4533 (N_4533,N_3514,N_3216);
xor U4534 (N_4534,N_3873,N_3356);
nor U4535 (N_4535,N_3669,N_3811);
nand U4536 (N_4536,N_3262,N_3095);
nand U4537 (N_4537,N_3229,N_3065);
or U4538 (N_4538,N_3869,N_3130);
xnor U4539 (N_4539,N_3406,N_3437);
and U4540 (N_4540,N_3942,N_3774);
and U4541 (N_4541,N_3077,N_3648);
nand U4542 (N_4542,N_3154,N_3279);
or U4543 (N_4543,N_3811,N_3635);
xor U4544 (N_4544,N_3685,N_3183);
nand U4545 (N_4545,N_3358,N_3849);
nor U4546 (N_4546,N_3290,N_3880);
or U4547 (N_4547,N_3900,N_3261);
nor U4548 (N_4548,N_3338,N_3451);
nand U4549 (N_4549,N_3009,N_3075);
nor U4550 (N_4550,N_3264,N_3605);
xor U4551 (N_4551,N_3968,N_3793);
or U4552 (N_4552,N_3956,N_3175);
or U4553 (N_4553,N_3070,N_3225);
and U4554 (N_4554,N_3039,N_3422);
nand U4555 (N_4555,N_3112,N_3720);
or U4556 (N_4556,N_3459,N_3374);
xnor U4557 (N_4557,N_3646,N_3066);
and U4558 (N_4558,N_3501,N_3680);
xnor U4559 (N_4559,N_3485,N_3362);
nor U4560 (N_4560,N_3103,N_3402);
xor U4561 (N_4561,N_3133,N_3754);
xnor U4562 (N_4562,N_3618,N_3689);
nor U4563 (N_4563,N_3213,N_3589);
nor U4564 (N_4564,N_3765,N_3900);
xor U4565 (N_4565,N_3369,N_3755);
or U4566 (N_4566,N_3284,N_3984);
and U4567 (N_4567,N_3350,N_3608);
xnor U4568 (N_4568,N_3003,N_3084);
xnor U4569 (N_4569,N_3726,N_3836);
nor U4570 (N_4570,N_3629,N_3320);
nand U4571 (N_4571,N_3761,N_3002);
nand U4572 (N_4572,N_3315,N_3200);
or U4573 (N_4573,N_3485,N_3552);
and U4574 (N_4574,N_3933,N_3287);
nand U4575 (N_4575,N_3431,N_3575);
nor U4576 (N_4576,N_3327,N_3531);
and U4577 (N_4577,N_3416,N_3019);
nand U4578 (N_4578,N_3064,N_3391);
xnor U4579 (N_4579,N_3933,N_3235);
xor U4580 (N_4580,N_3152,N_3548);
xor U4581 (N_4581,N_3570,N_3585);
and U4582 (N_4582,N_3170,N_3254);
nor U4583 (N_4583,N_3493,N_3441);
or U4584 (N_4584,N_3750,N_3495);
nor U4585 (N_4585,N_3029,N_3676);
nand U4586 (N_4586,N_3274,N_3863);
xor U4587 (N_4587,N_3593,N_3921);
xnor U4588 (N_4588,N_3439,N_3918);
and U4589 (N_4589,N_3314,N_3803);
nand U4590 (N_4590,N_3545,N_3469);
or U4591 (N_4591,N_3682,N_3773);
and U4592 (N_4592,N_3059,N_3166);
nor U4593 (N_4593,N_3009,N_3096);
xnor U4594 (N_4594,N_3102,N_3649);
or U4595 (N_4595,N_3785,N_3187);
or U4596 (N_4596,N_3460,N_3163);
xor U4597 (N_4597,N_3021,N_3591);
and U4598 (N_4598,N_3328,N_3064);
xor U4599 (N_4599,N_3615,N_3187);
xnor U4600 (N_4600,N_3363,N_3217);
nand U4601 (N_4601,N_3298,N_3523);
nor U4602 (N_4602,N_3047,N_3405);
and U4603 (N_4603,N_3470,N_3792);
or U4604 (N_4604,N_3907,N_3935);
nand U4605 (N_4605,N_3005,N_3057);
nand U4606 (N_4606,N_3484,N_3131);
or U4607 (N_4607,N_3948,N_3114);
or U4608 (N_4608,N_3339,N_3099);
nand U4609 (N_4609,N_3341,N_3215);
xnor U4610 (N_4610,N_3069,N_3015);
nand U4611 (N_4611,N_3526,N_3500);
nor U4612 (N_4612,N_3006,N_3598);
nand U4613 (N_4613,N_3334,N_3904);
nand U4614 (N_4614,N_3567,N_3214);
nor U4615 (N_4615,N_3404,N_3570);
nand U4616 (N_4616,N_3029,N_3882);
nor U4617 (N_4617,N_3931,N_3324);
xor U4618 (N_4618,N_3173,N_3717);
or U4619 (N_4619,N_3236,N_3479);
and U4620 (N_4620,N_3030,N_3726);
or U4621 (N_4621,N_3940,N_3204);
or U4622 (N_4622,N_3772,N_3171);
and U4623 (N_4623,N_3543,N_3560);
and U4624 (N_4624,N_3341,N_3581);
nor U4625 (N_4625,N_3590,N_3381);
xnor U4626 (N_4626,N_3838,N_3952);
nand U4627 (N_4627,N_3797,N_3713);
nand U4628 (N_4628,N_3175,N_3740);
or U4629 (N_4629,N_3737,N_3739);
nor U4630 (N_4630,N_3179,N_3773);
nor U4631 (N_4631,N_3469,N_3525);
nand U4632 (N_4632,N_3265,N_3533);
xor U4633 (N_4633,N_3606,N_3035);
and U4634 (N_4634,N_3524,N_3785);
nor U4635 (N_4635,N_3052,N_3670);
or U4636 (N_4636,N_3038,N_3595);
nor U4637 (N_4637,N_3057,N_3218);
and U4638 (N_4638,N_3115,N_3075);
or U4639 (N_4639,N_3749,N_3397);
xor U4640 (N_4640,N_3457,N_3590);
xor U4641 (N_4641,N_3194,N_3663);
and U4642 (N_4642,N_3877,N_3979);
or U4643 (N_4643,N_3747,N_3586);
xor U4644 (N_4644,N_3551,N_3224);
or U4645 (N_4645,N_3188,N_3646);
xor U4646 (N_4646,N_3498,N_3223);
or U4647 (N_4647,N_3285,N_3749);
nor U4648 (N_4648,N_3705,N_3818);
nor U4649 (N_4649,N_3822,N_3669);
and U4650 (N_4650,N_3989,N_3071);
xnor U4651 (N_4651,N_3868,N_3498);
and U4652 (N_4652,N_3017,N_3083);
nand U4653 (N_4653,N_3533,N_3973);
nor U4654 (N_4654,N_3730,N_3147);
and U4655 (N_4655,N_3089,N_3648);
nand U4656 (N_4656,N_3162,N_3833);
nor U4657 (N_4657,N_3478,N_3743);
xor U4658 (N_4658,N_3976,N_3511);
nor U4659 (N_4659,N_3014,N_3842);
and U4660 (N_4660,N_3930,N_3113);
nor U4661 (N_4661,N_3472,N_3719);
xnor U4662 (N_4662,N_3130,N_3273);
nor U4663 (N_4663,N_3779,N_3754);
xnor U4664 (N_4664,N_3615,N_3601);
xnor U4665 (N_4665,N_3855,N_3831);
xnor U4666 (N_4666,N_3267,N_3250);
and U4667 (N_4667,N_3915,N_3535);
and U4668 (N_4668,N_3538,N_3793);
nor U4669 (N_4669,N_3327,N_3272);
nor U4670 (N_4670,N_3000,N_3691);
nand U4671 (N_4671,N_3967,N_3451);
xor U4672 (N_4672,N_3806,N_3930);
nand U4673 (N_4673,N_3831,N_3524);
nor U4674 (N_4674,N_3999,N_3276);
nand U4675 (N_4675,N_3520,N_3465);
nand U4676 (N_4676,N_3142,N_3180);
and U4677 (N_4677,N_3583,N_3787);
nand U4678 (N_4678,N_3905,N_3775);
xnor U4679 (N_4679,N_3065,N_3789);
xnor U4680 (N_4680,N_3237,N_3445);
nor U4681 (N_4681,N_3987,N_3797);
xnor U4682 (N_4682,N_3249,N_3680);
nand U4683 (N_4683,N_3809,N_3568);
and U4684 (N_4684,N_3227,N_3202);
nor U4685 (N_4685,N_3302,N_3328);
or U4686 (N_4686,N_3031,N_3123);
nor U4687 (N_4687,N_3210,N_3313);
and U4688 (N_4688,N_3618,N_3705);
nor U4689 (N_4689,N_3634,N_3056);
nand U4690 (N_4690,N_3088,N_3725);
nand U4691 (N_4691,N_3560,N_3737);
nand U4692 (N_4692,N_3806,N_3173);
or U4693 (N_4693,N_3880,N_3256);
or U4694 (N_4694,N_3810,N_3373);
xnor U4695 (N_4695,N_3598,N_3970);
and U4696 (N_4696,N_3798,N_3919);
nand U4697 (N_4697,N_3119,N_3445);
and U4698 (N_4698,N_3175,N_3847);
nand U4699 (N_4699,N_3430,N_3095);
and U4700 (N_4700,N_3842,N_3427);
xnor U4701 (N_4701,N_3509,N_3490);
nor U4702 (N_4702,N_3141,N_3185);
xnor U4703 (N_4703,N_3172,N_3476);
or U4704 (N_4704,N_3979,N_3093);
nand U4705 (N_4705,N_3835,N_3465);
or U4706 (N_4706,N_3733,N_3437);
xor U4707 (N_4707,N_3093,N_3197);
and U4708 (N_4708,N_3310,N_3925);
nor U4709 (N_4709,N_3151,N_3408);
xnor U4710 (N_4710,N_3081,N_3036);
nand U4711 (N_4711,N_3096,N_3244);
and U4712 (N_4712,N_3926,N_3130);
nor U4713 (N_4713,N_3634,N_3134);
nand U4714 (N_4714,N_3413,N_3688);
nand U4715 (N_4715,N_3030,N_3393);
and U4716 (N_4716,N_3592,N_3354);
nor U4717 (N_4717,N_3570,N_3769);
xnor U4718 (N_4718,N_3409,N_3969);
or U4719 (N_4719,N_3379,N_3323);
nand U4720 (N_4720,N_3187,N_3362);
nor U4721 (N_4721,N_3918,N_3471);
xor U4722 (N_4722,N_3879,N_3041);
nor U4723 (N_4723,N_3573,N_3977);
xor U4724 (N_4724,N_3337,N_3634);
or U4725 (N_4725,N_3614,N_3525);
or U4726 (N_4726,N_3127,N_3995);
xnor U4727 (N_4727,N_3226,N_3276);
nor U4728 (N_4728,N_3723,N_3862);
nand U4729 (N_4729,N_3411,N_3543);
and U4730 (N_4730,N_3892,N_3016);
xor U4731 (N_4731,N_3153,N_3480);
nand U4732 (N_4732,N_3640,N_3475);
nor U4733 (N_4733,N_3050,N_3941);
and U4734 (N_4734,N_3524,N_3970);
nand U4735 (N_4735,N_3442,N_3697);
xnor U4736 (N_4736,N_3905,N_3197);
xor U4737 (N_4737,N_3839,N_3969);
and U4738 (N_4738,N_3433,N_3194);
nor U4739 (N_4739,N_3945,N_3150);
and U4740 (N_4740,N_3514,N_3535);
nand U4741 (N_4741,N_3084,N_3369);
nand U4742 (N_4742,N_3690,N_3379);
xor U4743 (N_4743,N_3885,N_3654);
xnor U4744 (N_4744,N_3962,N_3072);
and U4745 (N_4745,N_3119,N_3554);
nor U4746 (N_4746,N_3082,N_3481);
and U4747 (N_4747,N_3844,N_3733);
or U4748 (N_4748,N_3834,N_3150);
nor U4749 (N_4749,N_3987,N_3434);
xor U4750 (N_4750,N_3675,N_3309);
xnor U4751 (N_4751,N_3477,N_3623);
xnor U4752 (N_4752,N_3546,N_3138);
or U4753 (N_4753,N_3194,N_3235);
xor U4754 (N_4754,N_3228,N_3006);
nand U4755 (N_4755,N_3385,N_3362);
nor U4756 (N_4756,N_3891,N_3654);
or U4757 (N_4757,N_3278,N_3294);
nor U4758 (N_4758,N_3019,N_3919);
and U4759 (N_4759,N_3017,N_3976);
xor U4760 (N_4760,N_3652,N_3972);
nand U4761 (N_4761,N_3118,N_3268);
and U4762 (N_4762,N_3051,N_3947);
nor U4763 (N_4763,N_3463,N_3776);
xnor U4764 (N_4764,N_3641,N_3386);
and U4765 (N_4765,N_3640,N_3762);
nand U4766 (N_4766,N_3531,N_3131);
xnor U4767 (N_4767,N_3132,N_3425);
nor U4768 (N_4768,N_3017,N_3359);
xnor U4769 (N_4769,N_3859,N_3596);
and U4770 (N_4770,N_3350,N_3999);
xnor U4771 (N_4771,N_3437,N_3031);
and U4772 (N_4772,N_3356,N_3308);
nor U4773 (N_4773,N_3878,N_3090);
or U4774 (N_4774,N_3056,N_3030);
xor U4775 (N_4775,N_3825,N_3913);
nand U4776 (N_4776,N_3625,N_3135);
or U4777 (N_4777,N_3867,N_3182);
nand U4778 (N_4778,N_3048,N_3658);
or U4779 (N_4779,N_3967,N_3322);
or U4780 (N_4780,N_3381,N_3432);
nor U4781 (N_4781,N_3850,N_3473);
xnor U4782 (N_4782,N_3175,N_3039);
nor U4783 (N_4783,N_3599,N_3485);
xnor U4784 (N_4784,N_3781,N_3128);
and U4785 (N_4785,N_3365,N_3881);
or U4786 (N_4786,N_3427,N_3768);
nor U4787 (N_4787,N_3445,N_3296);
nand U4788 (N_4788,N_3530,N_3696);
xor U4789 (N_4789,N_3971,N_3966);
or U4790 (N_4790,N_3981,N_3106);
and U4791 (N_4791,N_3129,N_3716);
nor U4792 (N_4792,N_3467,N_3071);
nor U4793 (N_4793,N_3202,N_3314);
and U4794 (N_4794,N_3403,N_3798);
xnor U4795 (N_4795,N_3823,N_3081);
and U4796 (N_4796,N_3852,N_3481);
xnor U4797 (N_4797,N_3264,N_3067);
or U4798 (N_4798,N_3055,N_3094);
and U4799 (N_4799,N_3461,N_3934);
nor U4800 (N_4800,N_3664,N_3737);
and U4801 (N_4801,N_3127,N_3920);
nor U4802 (N_4802,N_3835,N_3860);
or U4803 (N_4803,N_3063,N_3500);
xnor U4804 (N_4804,N_3065,N_3215);
or U4805 (N_4805,N_3133,N_3826);
nand U4806 (N_4806,N_3007,N_3715);
and U4807 (N_4807,N_3225,N_3788);
nor U4808 (N_4808,N_3338,N_3734);
nor U4809 (N_4809,N_3186,N_3430);
nand U4810 (N_4810,N_3079,N_3378);
or U4811 (N_4811,N_3533,N_3536);
nand U4812 (N_4812,N_3159,N_3446);
xnor U4813 (N_4813,N_3779,N_3012);
xor U4814 (N_4814,N_3276,N_3425);
or U4815 (N_4815,N_3895,N_3224);
and U4816 (N_4816,N_3770,N_3641);
or U4817 (N_4817,N_3715,N_3756);
xnor U4818 (N_4818,N_3964,N_3803);
or U4819 (N_4819,N_3665,N_3260);
nor U4820 (N_4820,N_3835,N_3940);
or U4821 (N_4821,N_3722,N_3818);
nand U4822 (N_4822,N_3477,N_3937);
and U4823 (N_4823,N_3196,N_3057);
nor U4824 (N_4824,N_3258,N_3412);
nand U4825 (N_4825,N_3294,N_3943);
nor U4826 (N_4826,N_3266,N_3646);
nand U4827 (N_4827,N_3808,N_3005);
nand U4828 (N_4828,N_3350,N_3827);
nor U4829 (N_4829,N_3884,N_3863);
and U4830 (N_4830,N_3461,N_3207);
xor U4831 (N_4831,N_3933,N_3635);
or U4832 (N_4832,N_3276,N_3407);
nand U4833 (N_4833,N_3444,N_3979);
nor U4834 (N_4834,N_3727,N_3863);
nand U4835 (N_4835,N_3048,N_3216);
xnor U4836 (N_4836,N_3138,N_3979);
and U4837 (N_4837,N_3591,N_3760);
and U4838 (N_4838,N_3965,N_3329);
and U4839 (N_4839,N_3861,N_3653);
or U4840 (N_4840,N_3053,N_3870);
nand U4841 (N_4841,N_3565,N_3440);
nor U4842 (N_4842,N_3034,N_3065);
and U4843 (N_4843,N_3417,N_3952);
or U4844 (N_4844,N_3304,N_3968);
and U4845 (N_4845,N_3988,N_3392);
or U4846 (N_4846,N_3514,N_3177);
or U4847 (N_4847,N_3640,N_3189);
and U4848 (N_4848,N_3321,N_3323);
nor U4849 (N_4849,N_3930,N_3356);
and U4850 (N_4850,N_3985,N_3085);
xor U4851 (N_4851,N_3378,N_3515);
xor U4852 (N_4852,N_3933,N_3956);
nor U4853 (N_4853,N_3351,N_3141);
nor U4854 (N_4854,N_3172,N_3252);
nand U4855 (N_4855,N_3245,N_3680);
nor U4856 (N_4856,N_3373,N_3430);
or U4857 (N_4857,N_3593,N_3294);
xnor U4858 (N_4858,N_3386,N_3728);
nand U4859 (N_4859,N_3888,N_3477);
xnor U4860 (N_4860,N_3764,N_3651);
nor U4861 (N_4861,N_3578,N_3552);
xor U4862 (N_4862,N_3586,N_3981);
xor U4863 (N_4863,N_3116,N_3624);
xnor U4864 (N_4864,N_3494,N_3522);
or U4865 (N_4865,N_3762,N_3781);
and U4866 (N_4866,N_3529,N_3979);
nor U4867 (N_4867,N_3557,N_3281);
nand U4868 (N_4868,N_3189,N_3061);
xnor U4869 (N_4869,N_3262,N_3270);
xor U4870 (N_4870,N_3829,N_3477);
nand U4871 (N_4871,N_3227,N_3362);
xor U4872 (N_4872,N_3024,N_3769);
xnor U4873 (N_4873,N_3303,N_3158);
nand U4874 (N_4874,N_3116,N_3672);
and U4875 (N_4875,N_3581,N_3867);
nor U4876 (N_4876,N_3362,N_3991);
nand U4877 (N_4877,N_3532,N_3105);
nand U4878 (N_4878,N_3204,N_3259);
xnor U4879 (N_4879,N_3036,N_3216);
or U4880 (N_4880,N_3558,N_3646);
nor U4881 (N_4881,N_3472,N_3372);
and U4882 (N_4882,N_3851,N_3139);
nor U4883 (N_4883,N_3442,N_3639);
nand U4884 (N_4884,N_3744,N_3516);
or U4885 (N_4885,N_3371,N_3733);
and U4886 (N_4886,N_3283,N_3540);
or U4887 (N_4887,N_3973,N_3700);
or U4888 (N_4888,N_3862,N_3023);
or U4889 (N_4889,N_3966,N_3439);
nand U4890 (N_4890,N_3509,N_3940);
nor U4891 (N_4891,N_3686,N_3785);
or U4892 (N_4892,N_3879,N_3846);
xor U4893 (N_4893,N_3269,N_3008);
or U4894 (N_4894,N_3624,N_3637);
xnor U4895 (N_4895,N_3695,N_3100);
and U4896 (N_4896,N_3393,N_3202);
or U4897 (N_4897,N_3062,N_3762);
nand U4898 (N_4898,N_3909,N_3883);
xnor U4899 (N_4899,N_3817,N_3625);
nor U4900 (N_4900,N_3312,N_3152);
or U4901 (N_4901,N_3741,N_3074);
nand U4902 (N_4902,N_3981,N_3150);
or U4903 (N_4903,N_3654,N_3745);
nor U4904 (N_4904,N_3495,N_3325);
or U4905 (N_4905,N_3603,N_3425);
nand U4906 (N_4906,N_3098,N_3799);
nor U4907 (N_4907,N_3709,N_3988);
and U4908 (N_4908,N_3830,N_3738);
xnor U4909 (N_4909,N_3833,N_3849);
and U4910 (N_4910,N_3434,N_3042);
and U4911 (N_4911,N_3372,N_3115);
or U4912 (N_4912,N_3497,N_3410);
or U4913 (N_4913,N_3166,N_3523);
or U4914 (N_4914,N_3239,N_3330);
xor U4915 (N_4915,N_3925,N_3537);
nand U4916 (N_4916,N_3992,N_3041);
nor U4917 (N_4917,N_3220,N_3946);
and U4918 (N_4918,N_3705,N_3872);
xnor U4919 (N_4919,N_3113,N_3224);
or U4920 (N_4920,N_3539,N_3824);
nand U4921 (N_4921,N_3894,N_3957);
xnor U4922 (N_4922,N_3972,N_3724);
or U4923 (N_4923,N_3999,N_3311);
nor U4924 (N_4924,N_3749,N_3790);
nor U4925 (N_4925,N_3086,N_3489);
nand U4926 (N_4926,N_3375,N_3176);
and U4927 (N_4927,N_3780,N_3200);
and U4928 (N_4928,N_3340,N_3181);
nand U4929 (N_4929,N_3797,N_3896);
or U4930 (N_4930,N_3407,N_3557);
nor U4931 (N_4931,N_3448,N_3164);
or U4932 (N_4932,N_3588,N_3448);
or U4933 (N_4933,N_3608,N_3934);
nand U4934 (N_4934,N_3227,N_3799);
nor U4935 (N_4935,N_3409,N_3018);
and U4936 (N_4936,N_3839,N_3615);
nand U4937 (N_4937,N_3978,N_3238);
or U4938 (N_4938,N_3185,N_3289);
nand U4939 (N_4939,N_3803,N_3530);
or U4940 (N_4940,N_3965,N_3019);
nand U4941 (N_4941,N_3479,N_3344);
nand U4942 (N_4942,N_3960,N_3739);
nand U4943 (N_4943,N_3721,N_3062);
nand U4944 (N_4944,N_3165,N_3848);
nand U4945 (N_4945,N_3389,N_3969);
or U4946 (N_4946,N_3691,N_3613);
or U4947 (N_4947,N_3507,N_3721);
nor U4948 (N_4948,N_3387,N_3317);
and U4949 (N_4949,N_3081,N_3416);
or U4950 (N_4950,N_3745,N_3438);
nor U4951 (N_4951,N_3402,N_3613);
nor U4952 (N_4952,N_3573,N_3026);
or U4953 (N_4953,N_3344,N_3129);
and U4954 (N_4954,N_3157,N_3210);
nand U4955 (N_4955,N_3861,N_3724);
or U4956 (N_4956,N_3167,N_3012);
xnor U4957 (N_4957,N_3455,N_3793);
xor U4958 (N_4958,N_3761,N_3463);
and U4959 (N_4959,N_3749,N_3509);
or U4960 (N_4960,N_3706,N_3718);
and U4961 (N_4961,N_3884,N_3254);
nor U4962 (N_4962,N_3712,N_3531);
nand U4963 (N_4963,N_3714,N_3692);
xor U4964 (N_4964,N_3310,N_3849);
or U4965 (N_4965,N_3226,N_3560);
or U4966 (N_4966,N_3011,N_3291);
and U4967 (N_4967,N_3106,N_3262);
xor U4968 (N_4968,N_3583,N_3697);
nand U4969 (N_4969,N_3860,N_3722);
and U4970 (N_4970,N_3518,N_3222);
xnor U4971 (N_4971,N_3983,N_3873);
xor U4972 (N_4972,N_3134,N_3021);
and U4973 (N_4973,N_3584,N_3617);
nor U4974 (N_4974,N_3699,N_3710);
and U4975 (N_4975,N_3804,N_3280);
and U4976 (N_4976,N_3337,N_3093);
and U4977 (N_4977,N_3126,N_3591);
xnor U4978 (N_4978,N_3625,N_3308);
nand U4979 (N_4979,N_3249,N_3825);
nand U4980 (N_4980,N_3918,N_3414);
or U4981 (N_4981,N_3200,N_3008);
and U4982 (N_4982,N_3439,N_3678);
nand U4983 (N_4983,N_3562,N_3265);
and U4984 (N_4984,N_3804,N_3146);
xor U4985 (N_4985,N_3527,N_3871);
xor U4986 (N_4986,N_3125,N_3910);
xnor U4987 (N_4987,N_3482,N_3334);
nor U4988 (N_4988,N_3915,N_3302);
xor U4989 (N_4989,N_3685,N_3380);
xor U4990 (N_4990,N_3886,N_3841);
nand U4991 (N_4991,N_3839,N_3902);
xor U4992 (N_4992,N_3290,N_3174);
or U4993 (N_4993,N_3806,N_3214);
or U4994 (N_4994,N_3993,N_3281);
xnor U4995 (N_4995,N_3897,N_3499);
or U4996 (N_4996,N_3184,N_3703);
or U4997 (N_4997,N_3102,N_3612);
nor U4998 (N_4998,N_3419,N_3356);
nand U4999 (N_4999,N_3310,N_3674);
xor U5000 (N_5000,N_4644,N_4285);
xnor U5001 (N_5001,N_4040,N_4685);
xnor U5002 (N_5002,N_4201,N_4122);
and U5003 (N_5003,N_4664,N_4400);
nor U5004 (N_5004,N_4812,N_4905);
nor U5005 (N_5005,N_4688,N_4099);
nand U5006 (N_5006,N_4411,N_4478);
xor U5007 (N_5007,N_4647,N_4655);
or U5008 (N_5008,N_4728,N_4774);
nor U5009 (N_5009,N_4572,N_4289);
or U5010 (N_5010,N_4301,N_4799);
nor U5011 (N_5011,N_4928,N_4173);
nand U5012 (N_5012,N_4267,N_4456);
xnor U5013 (N_5013,N_4093,N_4243);
or U5014 (N_5014,N_4940,N_4869);
or U5015 (N_5015,N_4382,N_4840);
xnor U5016 (N_5016,N_4253,N_4380);
xnor U5017 (N_5017,N_4896,N_4874);
or U5018 (N_5018,N_4777,N_4074);
nor U5019 (N_5019,N_4439,N_4031);
nand U5020 (N_5020,N_4376,N_4534);
and U5021 (N_5021,N_4174,N_4300);
xor U5022 (N_5022,N_4436,N_4205);
nand U5023 (N_5023,N_4395,N_4689);
or U5024 (N_5024,N_4232,N_4111);
xnor U5025 (N_5025,N_4604,N_4442);
and U5026 (N_5026,N_4349,N_4352);
xnor U5027 (N_5027,N_4561,N_4316);
and U5028 (N_5028,N_4634,N_4729);
or U5029 (N_5029,N_4098,N_4318);
xor U5030 (N_5030,N_4657,N_4748);
nor U5031 (N_5031,N_4623,N_4498);
nand U5032 (N_5032,N_4895,N_4757);
or U5033 (N_5033,N_4533,N_4610);
nor U5034 (N_5034,N_4880,N_4992);
nand U5035 (N_5035,N_4104,N_4017);
or U5036 (N_5036,N_4373,N_4444);
xor U5037 (N_5037,N_4732,N_4161);
or U5038 (N_5038,N_4007,N_4867);
and U5039 (N_5039,N_4250,N_4523);
xnor U5040 (N_5040,N_4365,N_4771);
nand U5041 (N_5041,N_4706,N_4827);
nand U5042 (N_5042,N_4619,N_4203);
nand U5043 (N_5043,N_4509,N_4446);
nor U5044 (N_5044,N_4778,N_4787);
nor U5045 (N_5045,N_4507,N_4605);
or U5046 (N_5046,N_4493,N_4050);
nand U5047 (N_5047,N_4888,N_4396);
or U5048 (N_5048,N_4650,N_4629);
and U5049 (N_5049,N_4700,N_4680);
or U5050 (N_5050,N_4487,N_4183);
nand U5051 (N_5051,N_4035,N_4780);
nand U5052 (N_5052,N_4890,N_4701);
nor U5053 (N_5053,N_4162,N_4249);
nand U5054 (N_5054,N_4548,N_4851);
nor U5055 (N_5055,N_4772,N_4198);
or U5056 (N_5056,N_4437,N_4049);
nor U5057 (N_5057,N_4699,N_4625);
nand U5058 (N_5058,N_4026,N_4483);
nand U5059 (N_5059,N_4255,N_4987);
nor U5060 (N_5060,N_4025,N_4991);
nor U5061 (N_5061,N_4662,N_4043);
xnor U5062 (N_5062,N_4899,N_4990);
nand U5063 (N_5063,N_4052,N_4121);
xnor U5064 (N_5064,N_4838,N_4505);
and U5065 (N_5065,N_4305,N_4546);
nand U5066 (N_5066,N_4597,N_4480);
xor U5067 (N_5067,N_4003,N_4734);
or U5068 (N_5068,N_4583,N_4955);
nand U5069 (N_5069,N_4034,N_4310);
and U5070 (N_5070,N_4745,N_4835);
nand U5071 (N_5071,N_4348,N_4176);
nor U5072 (N_5072,N_4994,N_4138);
nand U5073 (N_5073,N_4753,N_4746);
xnor U5074 (N_5074,N_4918,N_4144);
nor U5075 (N_5075,N_4736,N_4384);
nor U5076 (N_5076,N_4872,N_4343);
xnor U5077 (N_5077,N_4520,N_4394);
and U5078 (N_5078,N_4926,N_4158);
xor U5079 (N_5079,N_4200,N_4627);
and U5080 (N_5080,N_4603,N_4132);
nor U5081 (N_5081,N_4042,N_4039);
and U5082 (N_5082,N_4624,N_4242);
or U5083 (N_5083,N_4543,N_4151);
xor U5084 (N_5084,N_4537,N_4709);
xnor U5085 (N_5085,N_4878,N_4751);
nor U5086 (N_5086,N_4501,N_4140);
nand U5087 (N_5087,N_4081,N_4403);
and U5088 (N_5088,N_4315,N_4054);
or U5089 (N_5089,N_4549,N_4862);
nor U5090 (N_5090,N_4370,N_4328);
or U5091 (N_5091,N_4166,N_4716);
nor U5092 (N_5092,N_4598,N_4186);
nor U5093 (N_5093,N_4526,N_4527);
or U5094 (N_5094,N_4494,N_4209);
nand U5095 (N_5095,N_4086,N_4666);
nand U5096 (N_5096,N_4171,N_4547);
nor U5097 (N_5097,N_4133,N_4968);
nand U5098 (N_5098,N_4196,N_4881);
nor U5099 (N_5099,N_4222,N_4574);
and U5100 (N_5100,N_4317,N_4973);
nand U5101 (N_5101,N_4333,N_4221);
nand U5102 (N_5102,N_4565,N_4539);
or U5103 (N_5103,N_4902,N_4855);
and U5104 (N_5104,N_4006,N_4087);
or U5105 (N_5105,N_4755,N_4649);
nor U5106 (N_5106,N_4635,N_4443);
nand U5107 (N_5107,N_4920,N_4988);
nand U5108 (N_5108,N_4180,N_4454);
or U5109 (N_5109,N_4187,N_4636);
and U5110 (N_5110,N_4225,N_4359);
xnor U5111 (N_5111,N_4207,N_4073);
nand U5112 (N_5112,N_4524,N_4739);
xor U5113 (N_5113,N_4379,N_4354);
xor U5114 (N_5114,N_4460,N_4268);
nor U5115 (N_5115,N_4492,N_4588);
nor U5116 (N_5116,N_4936,N_4149);
or U5117 (N_5117,N_4586,N_4450);
and U5118 (N_5118,N_4233,N_4894);
and U5119 (N_5119,N_4012,N_4361);
or U5120 (N_5120,N_4261,N_4488);
or U5121 (N_5121,N_4793,N_4303);
nand U5122 (N_5122,N_4287,N_4148);
nand U5123 (N_5123,N_4235,N_4847);
and U5124 (N_5124,N_4339,N_4229);
nand U5125 (N_5125,N_4815,N_4891);
nand U5126 (N_5126,N_4027,N_4782);
nand U5127 (N_5127,N_4230,N_4503);
xnor U5128 (N_5128,N_4368,N_4693);
and U5129 (N_5129,N_4977,N_4326);
nor U5130 (N_5130,N_4554,N_4959);
nor U5131 (N_5131,N_4115,N_4032);
and U5132 (N_5132,N_4834,N_4884);
and U5133 (N_5133,N_4848,N_4355);
and U5134 (N_5134,N_4786,N_4946);
and U5135 (N_5135,N_4291,N_4842);
nand U5136 (N_5136,N_4182,N_4455);
and U5137 (N_5137,N_4088,N_4796);
nor U5138 (N_5138,N_4393,N_4259);
xor U5139 (N_5139,N_4651,N_4504);
or U5140 (N_5140,N_4875,N_4925);
nor U5141 (N_5141,N_4475,N_4536);
nor U5142 (N_5142,N_4766,N_4468);
and U5143 (N_5143,N_4404,N_4117);
xor U5144 (N_5144,N_4105,N_4312);
and U5145 (N_5145,N_4298,N_4571);
and U5146 (N_5146,N_4877,N_4294);
and U5147 (N_5147,N_4555,N_4028);
nand U5148 (N_5148,N_4978,N_4691);
nor U5149 (N_5149,N_4570,N_4160);
or U5150 (N_5150,N_4553,N_4791);
and U5151 (N_5151,N_4727,N_4831);
and U5152 (N_5152,N_4417,N_4071);
and U5153 (N_5153,N_4900,N_4500);
and U5154 (N_5154,N_4270,N_4189);
nand U5155 (N_5155,N_4718,N_4731);
xor U5156 (N_5156,N_4841,N_4608);
xor U5157 (N_5157,N_4089,N_4542);
or U5158 (N_5158,N_4190,N_4957);
and U5159 (N_5159,N_4917,N_4418);
xnor U5160 (N_5160,N_4845,N_4750);
nor U5161 (N_5161,N_4515,N_4288);
nand U5162 (N_5162,N_4046,N_4083);
xnor U5163 (N_5163,N_4278,N_4550);
xnor U5164 (N_5164,N_4023,N_4996);
nand U5165 (N_5165,N_4541,N_4613);
nor U5166 (N_5166,N_4449,N_4257);
nor U5167 (N_5167,N_4084,N_4612);
and U5168 (N_5168,N_4065,N_4481);
xnor U5169 (N_5169,N_4128,N_4113);
or U5170 (N_5170,N_4932,N_4724);
and U5171 (N_5171,N_4309,N_4529);
or U5172 (N_5172,N_4414,N_4883);
xor U5173 (N_5173,N_4983,N_4765);
and U5174 (N_5174,N_4470,N_4824);
and U5175 (N_5175,N_4386,N_4663);
nand U5176 (N_5176,N_4425,N_4675);
nor U5177 (N_5177,N_4805,N_4726);
xor U5178 (N_5178,N_4029,N_4614);
nor U5179 (N_5179,N_4090,N_4217);
xor U5180 (N_5180,N_4826,N_4742);
nor U5181 (N_5181,N_4931,N_4281);
and U5182 (N_5182,N_4857,N_4611);
and U5183 (N_5183,N_4764,N_4949);
nand U5184 (N_5184,N_4051,N_4447);
and U5185 (N_5185,N_4882,N_4055);
or U5186 (N_5186,N_4810,N_4179);
and U5187 (N_5187,N_4356,N_4776);
or U5188 (N_5188,N_4756,N_4146);
or U5189 (N_5189,N_4513,N_4016);
nor U5190 (N_5190,N_4781,N_4477);
xor U5191 (N_5191,N_4346,N_4622);
nor U5192 (N_5192,N_4575,N_4423);
nand U5193 (N_5193,N_4410,N_4969);
and U5194 (N_5194,N_4817,N_4590);
and U5195 (N_5195,N_4214,N_4246);
nor U5196 (N_5196,N_4155,N_4206);
xnor U5197 (N_5197,N_4889,N_4276);
xnor U5198 (N_5198,N_4362,N_4019);
nand U5199 (N_5199,N_4697,N_4540);
nor U5200 (N_5200,N_4584,N_4979);
nor U5201 (N_5201,N_4157,N_4737);
or U5202 (N_5202,N_4602,N_4903);
nor U5203 (N_5203,N_4868,N_4342);
or U5204 (N_5204,N_4218,N_4364);
and U5205 (N_5205,N_4741,N_4702);
or U5206 (N_5206,N_4273,N_4599);
or U5207 (N_5207,N_4985,N_4910);
xor U5208 (N_5208,N_4467,N_4525);
nand U5209 (N_5209,N_4713,N_4596);
and U5210 (N_5210,N_4125,N_4405);
nand U5211 (N_5211,N_4951,N_4999);
nor U5212 (N_5212,N_4934,N_4407);
or U5213 (N_5213,N_4929,N_4095);
nand U5214 (N_5214,N_4124,N_4633);
xnor U5215 (N_5215,N_4156,N_4620);
and U5216 (N_5216,N_4448,N_4094);
nand U5217 (N_5217,N_4163,N_4683);
nor U5218 (N_5218,N_4808,N_4334);
and U5219 (N_5219,N_4427,N_4762);
and U5220 (N_5220,N_4272,N_4422);
or U5221 (N_5221,N_4723,N_4415);
and U5222 (N_5222,N_4814,N_4558);
xnor U5223 (N_5223,N_4402,N_4244);
nor U5224 (N_5224,N_4660,N_4357);
and U5225 (N_5225,N_4915,N_4464);
xor U5226 (N_5226,N_4856,N_4181);
or U5227 (N_5227,N_4961,N_4080);
xnor U5228 (N_5228,N_4528,N_4269);
xnor U5229 (N_5229,N_4068,N_4231);
or U5230 (N_5230,N_4307,N_4152);
xor U5231 (N_5231,N_4803,N_4820);
or U5232 (N_5232,N_4299,N_4559);
and U5233 (N_5233,N_4904,N_4811);
nor U5234 (N_5234,N_4632,N_4177);
xor U5235 (N_5235,N_4265,N_4906);
or U5236 (N_5236,N_4168,N_4863);
or U5237 (N_5237,N_4295,N_4564);
and U5238 (N_5238,N_4658,N_4981);
xor U5239 (N_5239,N_4210,N_4530);
nor U5240 (N_5240,N_4406,N_4954);
nand U5241 (N_5241,N_4616,N_4704);
or U5242 (N_5242,N_4953,N_4041);
nand U5243 (N_5243,N_4458,N_4413);
nor U5244 (N_5244,N_4252,N_4788);
and U5245 (N_5245,N_4129,N_4283);
and U5246 (N_5246,N_4577,N_4535);
nor U5247 (N_5247,N_4615,N_4112);
nand U5248 (N_5248,N_4669,N_4850);
nor U5249 (N_5249,N_4639,N_4369);
nand U5250 (N_5250,N_4710,N_4466);
nor U5251 (N_5251,N_4335,N_4784);
or U5252 (N_5252,N_4995,N_4116);
nor U5253 (N_5253,N_4347,N_4589);
xor U5254 (N_5254,N_4871,N_4421);
and U5255 (N_5255,N_4311,N_4677);
nand U5256 (N_5256,N_4075,N_4165);
nor U5257 (N_5257,N_4876,N_4219);
nand U5258 (N_5258,N_4545,N_4107);
nand U5259 (N_5259,N_4637,N_4927);
and U5260 (N_5260,N_4078,N_4816);
xor U5261 (N_5261,N_4594,N_4853);
nand U5262 (N_5262,N_4366,N_4514);
xor U5263 (N_5263,N_4519,N_4248);
nor U5264 (N_5264,N_4392,N_4892);
and U5265 (N_5265,N_4783,N_4818);
and U5266 (N_5266,N_4473,N_4127);
and U5267 (N_5267,N_4412,N_4795);
xnor U5268 (N_5268,N_4486,N_4169);
nand U5269 (N_5269,N_4433,N_4459);
or U5270 (N_5270,N_4997,N_4337);
xor U5271 (N_5271,N_4659,N_4692);
nand U5272 (N_5272,N_4792,N_4479);
and U5273 (N_5273,N_4293,N_4993);
nand U5274 (N_5274,N_4266,N_4371);
xor U5275 (N_5275,N_4937,N_4451);
nor U5276 (N_5276,N_4175,N_4211);
nor U5277 (N_5277,N_4092,N_4846);
nor U5278 (N_5278,N_4794,N_4308);
or U5279 (N_5279,N_4327,N_4005);
nand U5280 (N_5280,N_4282,N_4919);
nor U5281 (N_5281,N_4208,N_4101);
nor U5282 (N_5282,N_4076,N_4557);
nor U5283 (N_5283,N_4070,N_4806);
or U5284 (N_5284,N_4110,N_4164);
or U5285 (N_5285,N_4024,N_4943);
and U5286 (N_5286,N_4798,N_4332);
nand U5287 (N_5287,N_4061,N_4066);
nand U5288 (N_5288,N_4630,N_4409);
nor U5289 (N_5289,N_4383,N_4236);
and U5290 (N_5290,N_4401,N_4617);
nand U5291 (N_5291,N_4199,N_4518);
nor U5292 (N_5292,N_4560,N_4100);
or U5293 (N_5293,N_4930,N_4240);
nor U5294 (N_5294,N_4773,N_4429);
nand U5295 (N_5295,N_4375,N_4744);
nand U5296 (N_5296,N_4237,N_4801);
nand U5297 (N_5297,N_4419,N_4058);
and U5298 (N_5298,N_4829,N_4962);
or U5299 (N_5299,N_4592,N_4462);
and U5300 (N_5300,N_4667,N_4239);
and U5301 (N_5301,N_4472,N_4228);
xnor U5302 (N_5302,N_4956,N_4952);
nor U5303 (N_5303,N_4279,N_4135);
nor U5304 (N_5304,N_4984,N_4922);
nand U5305 (N_5305,N_4463,N_4690);
nor U5306 (N_5306,N_4004,N_4461);
or U5307 (N_5307,N_4976,N_4197);
nand U5308 (N_5308,N_4103,N_4673);
or U5309 (N_5309,N_4573,N_4989);
nand U5310 (N_5310,N_4367,N_4551);
xor U5311 (N_5311,N_4234,N_4566);
nor U5312 (N_5312,N_4313,N_4471);
nand U5313 (N_5313,N_4873,N_4695);
or U5314 (N_5314,N_4424,N_4652);
nor U5315 (N_5315,N_4569,N_4079);
or U5316 (N_5316,N_4011,N_4147);
xnor U5317 (N_5317,N_4185,N_4914);
nor U5318 (N_5318,N_4885,N_4843);
xor U5319 (N_5319,N_4223,N_4331);
nor U5320 (N_5320,N_4887,N_4262);
and U5321 (N_5321,N_4661,N_4057);
and U5322 (N_5322,N_4686,N_4747);
xor U5323 (N_5323,N_4452,N_4714);
or U5324 (N_5324,N_4568,N_4754);
or U5325 (N_5325,N_4769,N_4391);
or U5326 (N_5326,N_4469,N_4531);
xor U5327 (N_5327,N_4302,N_4966);
nor U5328 (N_5328,N_4290,N_4344);
nand U5329 (N_5329,N_4901,N_4581);
xnor U5330 (N_5330,N_4358,N_4607);
and U5331 (N_5331,N_4432,N_4247);
nor U5332 (N_5332,N_4681,N_4397);
and U5333 (N_5333,N_4759,N_4947);
xor U5334 (N_5334,N_4038,N_4251);
nor U5335 (N_5335,N_4002,N_4708);
nor U5336 (N_5336,N_4958,N_4172);
nand U5337 (N_5337,N_4482,N_4712);
nor U5338 (N_5338,N_4859,N_4563);
xor U5339 (N_5339,N_4921,N_4280);
xnor U5340 (N_5340,N_4213,N_4923);
and U5341 (N_5341,N_4552,N_4740);
nand U5342 (N_5342,N_4670,N_4950);
or U5343 (N_5343,N_4085,N_4705);
nand U5344 (N_5344,N_4321,N_4945);
nand U5345 (N_5345,N_4263,N_4067);
and U5346 (N_5346,N_4224,N_4434);
and U5347 (N_5347,N_4621,N_4114);
nand U5348 (N_5348,N_4858,N_4324);
and U5349 (N_5349,N_4329,N_4018);
nor U5350 (N_5350,N_4879,N_4506);
or U5351 (N_5351,N_4194,N_4353);
nand U5352 (N_5352,N_4284,N_4360);
xor U5353 (N_5353,N_4131,N_4532);
or U5354 (N_5354,N_4277,N_4678);
and U5355 (N_5355,N_4656,N_4045);
or U5356 (N_5356,N_4698,N_4687);
and U5357 (N_5357,N_4538,N_4153);
xor U5358 (N_5358,N_4516,N_4142);
nor U5359 (N_5359,N_4033,N_4490);
or U5360 (N_5360,N_4416,N_4001);
or U5361 (N_5361,N_4059,N_4441);
xor U5362 (N_5362,N_4595,N_4696);
or U5363 (N_5363,N_4338,N_4674);
nand U5364 (N_5364,N_4227,N_4886);
nor U5365 (N_5365,N_4913,N_4377);
or U5366 (N_5366,N_4735,N_4502);
nor U5367 (N_5367,N_4264,N_4591);
xnor U5368 (N_5368,N_4522,N_4580);
nand U5369 (N_5369,N_4258,N_4909);
nor U5370 (N_5370,N_4426,N_4865);
or U5371 (N_5371,N_4056,N_4420);
nand U5372 (N_5372,N_4489,N_4106);
xor U5373 (N_5373,N_4319,N_4982);
nor U5374 (N_5374,N_4960,N_4430);
nor U5375 (N_5375,N_4390,N_4567);
and U5376 (N_5376,N_4137,N_4738);
nand U5377 (N_5377,N_4216,N_4053);
nand U5378 (N_5378,N_4760,N_4752);
nand U5379 (N_5379,N_4768,N_4102);
nand U5380 (N_5380,N_4048,N_4167);
or U5381 (N_5381,N_4924,N_4435);
nand U5382 (N_5382,N_4220,N_4109);
and U5383 (N_5383,N_4226,N_4839);
and U5384 (N_5384,N_4517,N_4428);
and U5385 (N_5385,N_4296,N_4306);
nand U5386 (N_5386,N_4643,N_4512);
and U5387 (N_5387,N_4897,N_4665);
nor U5388 (N_5388,N_4378,N_4908);
or U5389 (N_5389,N_4556,N_4861);
and U5390 (N_5390,N_4495,N_4821);
nand U5391 (N_5391,N_4970,N_4314);
or U5392 (N_5392,N_4965,N_4297);
or U5393 (N_5393,N_4123,N_4802);
nor U5394 (N_5394,N_4134,N_4790);
or U5395 (N_5395,N_4485,N_4062);
or U5396 (N_5396,N_4476,N_4126);
nor U5397 (N_5397,N_4797,N_4854);
nor U5398 (N_5398,N_4195,N_4730);
xor U5399 (N_5399,N_4323,N_4941);
nor U5400 (N_5400,N_4626,N_4330);
or U5401 (N_5401,N_4912,N_4544);
xnor U5402 (N_5402,N_4682,N_4743);
and U5403 (N_5403,N_4143,N_4170);
and U5404 (N_5404,N_4204,N_4800);
xnor U5405 (N_5405,N_4648,N_4013);
nor U5406 (N_5406,N_4510,N_4136);
xnor U5407 (N_5407,N_4191,N_4091);
or U5408 (N_5408,N_4837,N_4641);
and U5409 (N_5409,N_4813,N_4082);
nor U5410 (N_5410,N_4438,N_4388);
nor U5411 (N_5411,N_4600,N_4980);
or U5412 (N_5412,N_4372,N_4119);
and U5413 (N_5413,N_4703,N_4351);
nand U5414 (N_5414,N_4188,N_4521);
or U5415 (N_5415,N_4000,N_4037);
nand U5416 (N_5416,N_4150,N_4496);
or U5417 (N_5417,N_4964,N_4638);
nor U5418 (N_5418,N_4178,N_4063);
nand U5419 (N_5419,N_4030,N_4047);
or U5420 (N_5420,N_4767,N_4807);
or U5421 (N_5421,N_4870,N_4381);
or U5422 (N_5422,N_4770,N_4275);
xnor U5423 (N_5423,N_4399,N_4864);
nor U5424 (N_5424,N_4491,N_4508);
xor U5425 (N_5425,N_4036,N_4653);
xnor U5426 (N_5426,N_4893,N_4852);
or U5427 (N_5427,N_4944,N_4916);
nand U5428 (N_5428,N_4907,N_4585);
and U5429 (N_5429,N_4154,N_4733);
xor U5430 (N_5430,N_4484,N_4866);
nor U5431 (N_5431,N_4830,N_4497);
nand U5432 (N_5432,N_4833,N_4322);
and U5433 (N_5433,N_4145,N_4974);
xor U5434 (N_5434,N_4779,N_4245);
or U5435 (N_5435,N_4008,N_4193);
xor U5436 (N_5436,N_4938,N_4933);
nor U5437 (N_5437,N_4679,N_4972);
or U5438 (N_5438,N_4044,N_4325);
xnor U5439 (N_5439,N_4825,N_4654);
or U5440 (N_5440,N_4758,N_4789);
xnor U5441 (N_5441,N_4832,N_4711);
nand U5442 (N_5442,N_4241,N_4350);
nand U5443 (N_5443,N_4587,N_4609);
or U5444 (N_5444,N_4971,N_4823);
nor U5445 (N_5445,N_4139,N_4785);
nand U5446 (N_5446,N_4749,N_4336);
or U5447 (N_5447,N_4120,N_4304);
xnor U5448 (N_5448,N_4986,N_4860);
or U5449 (N_5449,N_4722,N_4911);
xnor U5450 (N_5450,N_4676,N_4398);
nor U5451 (N_5451,N_4385,N_4717);
nand U5452 (N_5452,N_4819,N_4631);
and U5453 (N_5453,N_4671,N_4340);
or U5454 (N_5454,N_4286,N_4009);
and U5455 (N_5455,N_4341,N_4072);
and U5456 (N_5456,N_4271,N_4618);
and U5457 (N_5457,N_4363,N_4967);
xor U5458 (N_5458,N_4836,N_4345);
nor U5459 (N_5459,N_4060,N_4849);
xnor U5460 (N_5460,N_4474,N_4465);
or U5461 (N_5461,N_4064,N_4763);
nor U5462 (N_5462,N_4809,N_4431);
nor U5463 (N_5463,N_4720,N_4254);
and U5464 (N_5464,N_4828,N_4935);
nor U5465 (N_5465,N_4715,N_4292);
or U5466 (N_5466,N_4320,N_4260);
or U5467 (N_5467,N_4184,N_4721);
nor U5468 (N_5468,N_4453,N_4898);
xnor U5469 (N_5469,N_4694,N_4707);
and U5470 (N_5470,N_4387,N_4642);
and U5471 (N_5471,N_4077,N_4130);
nor U5472 (N_5472,N_4645,N_4719);
nor U5473 (N_5473,N_4640,N_4975);
nor U5474 (N_5474,N_4256,N_4822);
or U5475 (N_5475,N_4238,N_4593);
or U5476 (N_5476,N_4141,N_4511);
or U5477 (N_5477,N_4010,N_4069);
xnor U5478 (N_5478,N_4212,N_4646);
nor U5479 (N_5479,N_4020,N_4440);
nand U5480 (N_5480,N_4942,N_4948);
nand U5481 (N_5481,N_4274,N_4998);
xor U5482 (N_5482,N_4684,N_4579);
nor U5483 (N_5483,N_4445,N_4389);
nor U5484 (N_5484,N_4118,N_4761);
or U5485 (N_5485,N_4672,N_4215);
nor U5486 (N_5486,N_4775,N_4014);
nor U5487 (N_5487,N_4844,N_4963);
or U5488 (N_5488,N_4606,N_4015);
xnor U5489 (N_5489,N_4582,N_4939);
or U5490 (N_5490,N_4562,N_4628);
and U5491 (N_5491,N_4108,N_4408);
nor U5492 (N_5492,N_4668,N_4192);
nor U5493 (N_5493,N_4374,N_4202);
xor U5494 (N_5494,N_4159,N_4725);
and U5495 (N_5495,N_4097,N_4578);
nor U5496 (N_5496,N_4804,N_4576);
xor U5497 (N_5497,N_4022,N_4457);
nor U5498 (N_5498,N_4021,N_4499);
xor U5499 (N_5499,N_4601,N_4096);
and U5500 (N_5500,N_4181,N_4813);
nor U5501 (N_5501,N_4157,N_4701);
or U5502 (N_5502,N_4757,N_4066);
or U5503 (N_5503,N_4014,N_4040);
or U5504 (N_5504,N_4138,N_4278);
nand U5505 (N_5505,N_4267,N_4967);
nor U5506 (N_5506,N_4417,N_4211);
or U5507 (N_5507,N_4791,N_4890);
nand U5508 (N_5508,N_4104,N_4603);
xor U5509 (N_5509,N_4500,N_4564);
or U5510 (N_5510,N_4485,N_4991);
nor U5511 (N_5511,N_4600,N_4583);
nand U5512 (N_5512,N_4716,N_4892);
nor U5513 (N_5513,N_4210,N_4307);
and U5514 (N_5514,N_4584,N_4207);
xnor U5515 (N_5515,N_4228,N_4262);
nand U5516 (N_5516,N_4435,N_4980);
nor U5517 (N_5517,N_4057,N_4376);
or U5518 (N_5518,N_4658,N_4121);
xnor U5519 (N_5519,N_4802,N_4292);
nand U5520 (N_5520,N_4307,N_4521);
and U5521 (N_5521,N_4948,N_4590);
and U5522 (N_5522,N_4778,N_4791);
or U5523 (N_5523,N_4872,N_4965);
and U5524 (N_5524,N_4789,N_4991);
or U5525 (N_5525,N_4175,N_4405);
and U5526 (N_5526,N_4172,N_4070);
and U5527 (N_5527,N_4366,N_4557);
nand U5528 (N_5528,N_4431,N_4650);
nand U5529 (N_5529,N_4879,N_4630);
xor U5530 (N_5530,N_4513,N_4777);
xor U5531 (N_5531,N_4740,N_4735);
nand U5532 (N_5532,N_4075,N_4282);
xnor U5533 (N_5533,N_4668,N_4310);
xor U5534 (N_5534,N_4429,N_4206);
nor U5535 (N_5535,N_4412,N_4870);
xor U5536 (N_5536,N_4582,N_4704);
nor U5537 (N_5537,N_4531,N_4375);
nand U5538 (N_5538,N_4402,N_4635);
nand U5539 (N_5539,N_4651,N_4645);
and U5540 (N_5540,N_4596,N_4715);
and U5541 (N_5541,N_4288,N_4487);
nand U5542 (N_5542,N_4732,N_4811);
nand U5543 (N_5543,N_4512,N_4093);
and U5544 (N_5544,N_4141,N_4699);
and U5545 (N_5545,N_4040,N_4430);
and U5546 (N_5546,N_4193,N_4216);
and U5547 (N_5547,N_4985,N_4197);
and U5548 (N_5548,N_4276,N_4722);
nand U5549 (N_5549,N_4863,N_4144);
nand U5550 (N_5550,N_4497,N_4772);
and U5551 (N_5551,N_4708,N_4262);
and U5552 (N_5552,N_4295,N_4126);
nor U5553 (N_5553,N_4051,N_4332);
and U5554 (N_5554,N_4446,N_4884);
or U5555 (N_5555,N_4907,N_4178);
and U5556 (N_5556,N_4055,N_4288);
xnor U5557 (N_5557,N_4389,N_4505);
xnor U5558 (N_5558,N_4022,N_4380);
nor U5559 (N_5559,N_4463,N_4267);
and U5560 (N_5560,N_4927,N_4857);
or U5561 (N_5561,N_4678,N_4646);
or U5562 (N_5562,N_4981,N_4099);
nor U5563 (N_5563,N_4991,N_4740);
and U5564 (N_5564,N_4711,N_4224);
nand U5565 (N_5565,N_4565,N_4060);
and U5566 (N_5566,N_4569,N_4468);
nor U5567 (N_5567,N_4548,N_4180);
nand U5568 (N_5568,N_4062,N_4110);
xnor U5569 (N_5569,N_4098,N_4994);
or U5570 (N_5570,N_4987,N_4506);
and U5571 (N_5571,N_4071,N_4591);
nor U5572 (N_5572,N_4204,N_4880);
nor U5573 (N_5573,N_4633,N_4677);
and U5574 (N_5574,N_4201,N_4760);
xnor U5575 (N_5575,N_4632,N_4046);
and U5576 (N_5576,N_4131,N_4608);
nand U5577 (N_5577,N_4986,N_4197);
and U5578 (N_5578,N_4881,N_4830);
xor U5579 (N_5579,N_4928,N_4900);
and U5580 (N_5580,N_4856,N_4136);
xnor U5581 (N_5581,N_4994,N_4166);
and U5582 (N_5582,N_4870,N_4811);
xor U5583 (N_5583,N_4130,N_4427);
nand U5584 (N_5584,N_4490,N_4755);
or U5585 (N_5585,N_4984,N_4849);
nor U5586 (N_5586,N_4775,N_4920);
nand U5587 (N_5587,N_4133,N_4515);
xor U5588 (N_5588,N_4021,N_4528);
and U5589 (N_5589,N_4918,N_4288);
and U5590 (N_5590,N_4375,N_4688);
or U5591 (N_5591,N_4046,N_4874);
xnor U5592 (N_5592,N_4285,N_4723);
nor U5593 (N_5593,N_4503,N_4940);
and U5594 (N_5594,N_4030,N_4507);
nor U5595 (N_5595,N_4876,N_4923);
nor U5596 (N_5596,N_4565,N_4399);
nand U5597 (N_5597,N_4262,N_4196);
nand U5598 (N_5598,N_4129,N_4287);
and U5599 (N_5599,N_4228,N_4730);
nand U5600 (N_5600,N_4955,N_4438);
nor U5601 (N_5601,N_4883,N_4966);
xor U5602 (N_5602,N_4708,N_4765);
xnor U5603 (N_5603,N_4572,N_4643);
nor U5604 (N_5604,N_4307,N_4600);
xor U5605 (N_5605,N_4796,N_4207);
nand U5606 (N_5606,N_4234,N_4663);
xnor U5607 (N_5607,N_4957,N_4192);
nand U5608 (N_5608,N_4047,N_4606);
xor U5609 (N_5609,N_4445,N_4318);
nand U5610 (N_5610,N_4301,N_4393);
nand U5611 (N_5611,N_4174,N_4685);
xnor U5612 (N_5612,N_4055,N_4280);
and U5613 (N_5613,N_4680,N_4498);
nand U5614 (N_5614,N_4721,N_4787);
nand U5615 (N_5615,N_4943,N_4559);
nor U5616 (N_5616,N_4237,N_4291);
nand U5617 (N_5617,N_4197,N_4129);
or U5618 (N_5618,N_4309,N_4907);
nand U5619 (N_5619,N_4272,N_4915);
nor U5620 (N_5620,N_4223,N_4591);
or U5621 (N_5621,N_4388,N_4792);
and U5622 (N_5622,N_4116,N_4202);
nand U5623 (N_5623,N_4485,N_4746);
xor U5624 (N_5624,N_4328,N_4408);
nor U5625 (N_5625,N_4771,N_4413);
nor U5626 (N_5626,N_4188,N_4237);
nand U5627 (N_5627,N_4660,N_4768);
xnor U5628 (N_5628,N_4072,N_4121);
or U5629 (N_5629,N_4561,N_4953);
or U5630 (N_5630,N_4627,N_4537);
nand U5631 (N_5631,N_4799,N_4769);
and U5632 (N_5632,N_4184,N_4051);
and U5633 (N_5633,N_4632,N_4363);
nand U5634 (N_5634,N_4412,N_4976);
nor U5635 (N_5635,N_4323,N_4004);
nor U5636 (N_5636,N_4066,N_4470);
nor U5637 (N_5637,N_4312,N_4167);
nand U5638 (N_5638,N_4645,N_4916);
nand U5639 (N_5639,N_4923,N_4566);
and U5640 (N_5640,N_4514,N_4556);
nor U5641 (N_5641,N_4216,N_4798);
or U5642 (N_5642,N_4756,N_4742);
nand U5643 (N_5643,N_4746,N_4291);
xnor U5644 (N_5644,N_4612,N_4015);
nand U5645 (N_5645,N_4221,N_4613);
nor U5646 (N_5646,N_4858,N_4344);
and U5647 (N_5647,N_4899,N_4416);
or U5648 (N_5648,N_4921,N_4756);
and U5649 (N_5649,N_4632,N_4829);
nand U5650 (N_5650,N_4408,N_4832);
or U5651 (N_5651,N_4109,N_4036);
or U5652 (N_5652,N_4492,N_4863);
nor U5653 (N_5653,N_4178,N_4424);
xnor U5654 (N_5654,N_4954,N_4335);
and U5655 (N_5655,N_4857,N_4075);
nor U5656 (N_5656,N_4566,N_4364);
nor U5657 (N_5657,N_4142,N_4177);
xnor U5658 (N_5658,N_4919,N_4284);
xor U5659 (N_5659,N_4793,N_4286);
and U5660 (N_5660,N_4811,N_4592);
or U5661 (N_5661,N_4054,N_4506);
nor U5662 (N_5662,N_4339,N_4356);
or U5663 (N_5663,N_4855,N_4324);
nor U5664 (N_5664,N_4787,N_4654);
nor U5665 (N_5665,N_4775,N_4033);
and U5666 (N_5666,N_4990,N_4096);
xor U5667 (N_5667,N_4196,N_4714);
nand U5668 (N_5668,N_4448,N_4632);
and U5669 (N_5669,N_4940,N_4310);
nor U5670 (N_5670,N_4456,N_4369);
or U5671 (N_5671,N_4366,N_4476);
and U5672 (N_5672,N_4032,N_4122);
nand U5673 (N_5673,N_4150,N_4212);
and U5674 (N_5674,N_4988,N_4090);
nand U5675 (N_5675,N_4848,N_4901);
nor U5676 (N_5676,N_4755,N_4051);
nor U5677 (N_5677,N_4790,N_4612);
nor U5678 (N_5678,N_4525,N_4441);
xnor U5679 (N_5679,N_4217,N_4957);
xnor U5680 (N_5680,N_4621,N_4428);
xor U5681 (N_5681,N_4185,N_4547);
nor U5682 (N_5682,N_4041,N_4597);
xor U5683 (N_5683,N_4204,N_4424);
and U5684 (N_5684,N_4903,N_4716);
and U5685 (N_5685,N_4612,N_4028);
or U5686 (N_5686,N_4201,N_4428);
nor U5687 (N_5687,N_4180,N_4885);
nand U5688 (N_5688,N_4660,N_4344);
and U5689 (N_5689,N_4472,N_4846);
nor U5690 (N_5690,N_4825,N_4474);
nand U5691 (N_5691,N_4610,N_4481);
or U5692 (N_5692,N_4782,N_4417);
and U5693 (N_5693,N_4506,N_4115);
xnor U5694 (N_5694,N_4683,N_4268);
and U5695 (N_5695,N_4031,N_4105);
nor U5696 (N_5696,N_4289,N_4375);
or U5697 (N_5697,N_4481,N_4096);
or U5698 (N_5698,N_4457,N_4267);
xnor U5699 (N_5699,N_4242,N_4402);
and U5700 (N_5700,N_4273,N_4649);
or U5701 (N_5701,N_4484,N_4951);
xor U5702 (N_5702,N_4042,N_4889);
nand U5703 (N_5703,N_4006,N_4380);
xnor U5704 (N_5704,N_4650,N_4728);
nand U5705 (N_5705,N_4783,N_4024);
nor U5706 (N_5706,N_4004,N_4155);
xnor U5707 (N_5707,N_4246,N_4011);
or U5708 (N_5708,N_4579,N_4486);
and U5709 (N_5709,N_4708,N_4304);
nor U5710 (N_5710,N_4892,N_4705);
and U5711 (N_5711,N_4508,N_4400);
nand U5712 (N_5712,N_4518,N_4565);
or U5713 (N_5713,N_4954,N_4818);
nor U5714 (N_5714,N_4556,N_4385);
and U5715 (N_5715,N_4034,N_4719);
nor U5716 (N_5716,N_4270,N_4815);
nand U5717 (N_5717,N_4182,N_4213);
and U5718 (N_5718,N_4257,N_4787);
or U5719 (N_5719,N_4650,N_4974);
or U5720 (N_5720,N_4393,N_4203);
or U5721 (N_5721,N_4581,N_4055);
nor U5722 (N_5722,N_4997,N_4114);
nor U5723 (N_5723,N_4121,N_4869);
or U5724 (N_5724,N_4330,N_4717);
or U5725 (N_5725,N_4669,N_4367);
nor U5726 (N_5726,N_4406,N_4419);
xor U5727 (N_5727,N_4157,N_4445);
nor U5728 (N_5728,N_4416,N_4916);
xnor U5729 (N_5729,N_4024,N_4929);
and U5730 (N_5730,N_4222,N_4981);
nand U5731 (N_5731,N_4313,N_4088);
xor U5732 (N_5732,N_4264,N_4702);
nand U5733 (N_5733,N_4268,N_4113);
nand U5734 (N_5734,N_4784,N_4720);
xnor U5735 (N_5735,N_4832,N_4476);
nor U5736 (N_5736,N_4703,N_4781);
or U5737 (N_5737,N_4592,N_4214);
and U5738 (N_5738,N_4605,N_4694);
xor U5739 (N_5739,N_4574,N_4077);
nor U5740 (N_5740,N_4935,N_4433);
xor U5741 (N_5741,N_4610,N_4710);
nor U5742 (N_5742,N_4709,N_4168);
and U5743 (N_5743,N_4112,N_4165);
nor U5744 (N_5744,N_4773,N_4300);
nor U5745 (N_5745,N_4240,N_4215);
nor U5746 (N_5746,N_4888,N_4206);
or U5747 (N_5747,N_4646,N_4766);
or U5748 (N_5748,N_4816,N_4275);
nor U5749 (N_5749,N_4619,N_4021);
or U5750 (N_5750,N_4489,N_4929);
nor U5751 (N_5751,N_4294,N_4878);
or U5752 (N_5752,N_4517,N_4745);
and U5753 (N_5753,N_4969,N_4272);
xor U5754 (N_5754,N_4015,N_4781);
nand U5755 (N_5755,N_4989,N_4728);
or U5756 (N_5756,N_4681,N_4918);
nor U5757 (N_5757,N_4782,N_4852);
or U5758 (N_5758,N_4677,N_4715);
nor U5759 (N_5759,N_4685,N_4715);
nand U5760 (N_5760,N_4223,N_4759);
and U5761 (N_5761,N_4897,N_4615);
nor U5762 (N_5762,N_4229,N_4697);
xnor U5763 (N_5763,N_4999,N_4858);
and U5764 (N_5764,N_4063,N_4427);
and U5765 (N_5765,N_4411,N_4089);
nor U5766 (N_5766,N_4486,N_4493);
or U5767 (N_5767,N_4196,N_4225);
or U5768 (N_5768,N_4516,N_4018);
nor U5769 (N_5769,N_4831,N_4665);
nor U5770 (N_5770,N_4049,N_4384);
nand U5771 (N_5771,N_4730,N_4216);
nand U5772 (N_5772,N_4136,N_4639);
and U5773 (N_5773,N_4083,N_4876);
and U5774 (N_5774,N_4586,N_4959);
xnor U5775 (N_5775,N_4733,N_4938);
or U5776 (N_5776,N_4832,N_4574);
nand U5777 (N_5777,N_4257,N_4358);
nor U5778 (N_5778,N_4764,N_4396);
and U5779 (N_5779,N_4817,N_4343);
nand U5780 (N_5780,N_4255,N_4956);
xor U5781 (N_5781,N_4604,N_4925);
and U5782 (N_5782,N_4045,N_4325);
xnor U5783 (N_5783,N_4863,N_4726);
nor U5784 (N_5784,N_4771,N_4391);
or U5785 (N_5785,N_4974,N_4267);
and U5786 (N_5786,N_4349,N_4645);
nand U5787 (N_5787,N_4186,N_4923);
or U5788 (N_5788,N_4424,N_4208);
xor U5789 (N_5789,N_4442,N_4022);
nand U5790 (N_5790,N_4005,N_4810);
nand U5791 (N_5791,N_4722,N_4325);
or U5792 (N_5792,N_4511,N_4588);
and U5793 (N_5793,N_4445,N_4410);
nor U5794 (N_5794,N_4206,N_4877);
or U5795 (N_5795,N_4662,N_4801);
xor U5796 (N_5796,N_4990,N_4020);
or U5797 (N_5797,N_4875,N_4163);
nor U5798 (N_5798,N_4063,N_4202);
xnor U5799 (N_5799,N_4799,N_4756);
or U5800 (N_5800,N_4998,N_4152);
nor U5801 (N_5801,N_4930,N_4268);
and U5802 (N_5802,N_4374,N_4850);
xnor U5803 (N_5803,N_4391,N_4587);
nor U5804 (N_5804,N_4882,N_4826);
xnor U5805 (N_5805,N_4090,N_4275);
and U5806 (N_5806,N_4739,N_4764);
xor U5807 (N_5807,N_4313,N_4347);
and U5808 (N_5808,N_4912,N_4409);
or U5809 (N_5809,N_4819,N_4677);
nor U5810 (N_5810,N_4778,N_4451);
xor U5811 (N_5811,N_4739,N_4113);
and U5812 (N_5812,N_4097,N_4142);
and U5813 (N_5813,N_4158,N_4433);
nor U5814 (N_5814,N_4058,N_4913);
nor U5815 (N_5815,N_4768,N_4865);
nor U5816 (N_5816,N_4833,N_4355);
nand U5817 (N_5817,N_4094,N_4761);
and U5818 (N_5818,N_4977,N_4777);
nand U5819 (N_5819,N_4781,N_4195);
or U5820 (N_5820,N_4221,N_4175);
and U5821 (N_5821,N_4677,N_4332);
and U5822 (N_5822,N_4191,N_4007);
nor U5823 (N_5823,N_4025,N_4151);
nor U5824 (N_5824,N_4304,N_4963);
and U5825 (N_5825,N_4293,N_4749);
nor U5826 (N_5826,N_4870,N_4356);
and U5827 (N_5827,N_4790,N_4620);
xor U5828 (N_5828,N_4061,N_4012);
or U5829 (N_5829,N_4570,N_4291);
or U5830 (N_5830,N_4075,N_4065);
nor U5831 (N_5831,N_4380,N_4591);
or U5832 (N_5832,N_4424,N_4266);
nor U5833 (N_5833,N_4763,N_4672);
nand U5834 (N_5834,N_4693,N_4630);
xor U5835 (N_5835,N_4391,N_4932);
nor U5836 (N_5836,N_4040,N_4624);
and U5837 (N_5837,N_4143,N_4570);
and U5838 (N_5838,N_4555,N_4397);
nand U5839 (N_5839,N_4936,N_4650);
xor U5840 (N_5840,N_4860,N_4401);
nand U5841 (N_5841,N_4234,N_4077);
and U5842 (N_5842,N_4071,N_4571);
nand U5843 (N_5843,N_4769,N_4952);
and U5844 (N_5844,N_4672,N_4088);
nand U5845 (N_5845,N_4060,N_4582);
nor U5846 (N_5846,N_4503,N_4122);
xor U5847 (N_5847,N_4798,N_4513);
nor U5848 (N_5848,N_4330,N_4341);
nor U5849 (N_5849,N_4940,N_4699);
xnor U5850 (N_5850,N_4776,N_4503);
and U5851 (N_5851,N_4464,N_4740);
and U5852 (N_5852,N_4156,N_4294);
xnor U5853 (N_5853,N_4266,N_4809);
nor U5854 (N_5854,N_4946,N_4959);
nand U5855 (N_5855,N_4149,N_4176);
or U5856 (N_5856,N_4536,N_4858);
and U5857 (N_5857,N_4212,N_4259);
or U5858 (N_5858,N_4736,N_4350);
nor U5859 (N_5859,N_4632,N_4993);
nor U5860 (N_5860,N_4127,N_4289);
nand U5861 (N_5861,N_4407,N_4847);
nand U5862 (N_5862,N_4216,N_4900);
nand U5863 (N_5863,N_4678,N_4169);
nor U5864 (N_5864,N_4714,N_4533);
nor U5865 (N_5865,N_4986,N_4045);
nand U5866 (N_5866,N_4755,N_4489);
xor U5867 (N_5867,N_4676,N_4153);
or U5868 (N_5868,N_4314,N_4521);
and U5869 (N_5869,N_4883,N_4056);
xor U5870 (N_5870,N_4758,N_4028);
and U5871 (N_5871,N_4258,N_4705);
and U5872 (N_5872,N_4945,N_4650);
nand U5873 (N_5873,N_4411,N_4567);
xor U5874 (N_5874,N_4149,N_4322);
nor U5875 (N_5875,N_4157,N_4341);
nor U5876 (N_5876,N_4412,N_4064);
xnor U5877 (N_5877,N_4826,N_4682);
nand U5878 (N_5878,N_4766,N_4012);
xor U5879 (N_5879,N_4472,N_4861);
nand U5880 (N_5880,N_4301,N_4033);
or U5881 (N_5881,N_4869,N_4452);
and U5882 (N_5882,N_4145,N_4850);
xnor U5883 (N_5883,N_4240,N_4066);
and U5884 (N_5884,N_4193,N_4422);
nor U5885 (N_5885,N_4370,N_4073);
nand U5886 (N_5886,N_4646,N_4802);
and U5887 (N_5887,N_4102,N_4885);
or U5888 (N_5888,N_4540,N_4882);
nor U5889 (N_5889,N_4638,N_4888);
nand U5890 (N_5890,N_4907,N_4139);
or U5891 (N_5891,N_4052,N_4723);
xnor U5892 (N_5892,N_4206,N_4066);
xor U5893 (N_5893,N_4494,N_4398);
and U5894 (N_5894,N_4957,N_4979);
nand U5895 (N_5895,N_4417,N_4162);
or U5896 (N_5896,N_4570,N_4372);
and U5897 (N_5897,N_4299,N_4893);
xnor U5898 (N_5898,N_4629,N_4534);
and U5899 (N_5899,N_4190,N_4381);
or U5900 (N_5900,N_4607,N_4757);
or U5901 (N_5901,N_4715,N_4159);
and U5902 (N_5902,N_4052,N_4252);
and U5903 (N_5903,N_4864,N_4760);
nor U5904 (N_5904,N_4330,N_4905);
and U5905 (N_5905,N_4604,N_4361);
nor U5906 (N_5906,N_4213,N_4825);
xor U5907 (N_5907,N_4718,N_4249);
xor U5908 (N_5908,N_4073,N_4749);
and U5909 (N_5909,N_4617,N_4125);
xnor U5910 (N_5910,N_4039,N_4665);
nand U5911 (N_5911,N_4034,N_4170);
nand U5912 (N_5912,N_4800,N_4487);
xor U5913 (N_5913,N_4995,N_4886);
nand U5914 (N_5914,N_4985,N_4522);
nand U5915 (N_5915,N_4558,N_4962);
or U5916 (N_5916,N_4255,N_4257);
xor U5917 (N_5917,N_4421,N_4384);
or U5918 (N_5918,N_4249,N_4657);
nor U5919 (N_5919,N_4908,N_4791);
nand U5920 (N_5920,N_4381,N_4359);
xor U5921 (N_5921,N_4420,N_4664);
nand U5922 (N_5922,N_4841,N_4171);
xnor U5923 (N_5923,N_4267,N_4022);
nor U5924 (N_5924,N_4398,N_4122);
or U5925 (N_5925,N_4579,N_4929);
and U5926 (N_5926,N_4571,N_4873);
xor U5927 (N_5927,N_4455,N_4766);
xnor U5928 (N_5928,N_4282,N_4922);
or U5929 (N_5929,N_4962,N_4597);
or U5930 (N_5930,N_4863,N_4222);
xnor U5931 (N_5931,N_4266,N_4004);
nor U5932 (N_5932,N_4360,N_4572);
xnor U5933 (N_5933,N_4780,N_4845);
xor U5934 (N_5934,N_4075,N_4499);
nor U5935 (N_5935,N_4723,N_4946);
nand U5936 (N_5936,N_4234,N_4935);
nor U5937 (N_5937,N_4285,N_4432);
nand U5938 (N_5938,N_4746,N_4804);
or U5939 (N_5939,N_4390,N_4437);
xnor U5940 (N_5940,N_4447,N_4144);
and U5941 (N_5941,N_4049,N_4205);
or U5942 (N_5942,N_4503,N_4838);
or U5943 (N_5943,N_4785,N_4531);
or U5944 (N_5944,N_4229,N_4453);
or U5945 (N_5945,N_4712,N_4287);
nor U5946 (N_5946,N_4868,N_4995);
nor U5947 (N_5947,N_4700,N_4887);
xnor U5948 (N_5948,N_4484,N_4985);
or U5949 (N_5949,N_4525,N_4243);
and U5950 (N_5950,N_4868,N_4637);
or U5951 (N_5951,N_4302,N_4814);
nand U5952 (N_5952,N_4409,N_4399);
nand U5953 (N_5953,N_4300,N_4217);
nor U5954 (N_5954,N_4274,N_4900);
nand U5955 (N_5955,N_4586,N_4667);
nand U5956 (N_5956,N_4721,N_4255);
and U5957 (N_5957,N_4803,N_4836);
nand U5958 (N_5958,N_4145,N_4082);
or U5959 (N_5959,N_4442,N_4370);
nor U5960 (N_5960,N_4364,N_4935);
and U5961 (N_5961,N_4327,N_4384);
or U5962 (N_5962,N_4033,N_4507);
nand U5963 (N_5963,N_4521,N_4805);
xnor U5964 (N_5964,N_4333,N_4544);
and U5965 (N_5965,N_4637,N_4359);
xor U5966 (N_5966,N_4991,N_4920);
nor U5967 (N_5967,N_4747,N_4035);
xor U5968 (N_5968,N_4844,N_4719);
xor U5969 (N_5969,N_4035,N_4758);
nor U5970 (N_5970,N_4856,N_4925);
xnor U5971 (N_5971,N_4014,N_4690);
and U5972 (N_5972,N_4557,N_4330);
xor U5973 (N_5973,N_4766,N_4796);
and U5974 (N_5974,N_4867,N_4504);
or U5975 (N_5975,N_4382,N_4865);
nor U5976 (N_5976,N_4705,N_4872);
and U5977 (N_5977,N_4084,N_4577);
and U5978 (N_5978,N_4119,N_4168);
and U5979 (N_5979,N_4432,N_4543);
xor U5980 (N_5980,N_4879,N_4042);
and U5981 (N_5981,N_4817,N_4011);
nand U5982 (N_5982,N_4926,N_4925);
nor U5983 (N_5983,N_4024,N_4033);
or U5984 (N_5984,N_4061,N_4357);
xnor U5985 (N_5985,N_4438,N_4794);
nand U5986 (N_5986,N_4194,N_4624);
xor U5987 (N_5987,N_4160,N_4801);
nor U5988 (N_5988,N_4386,N_4868);
nand U5989 (N_5989,N_4474,N_4729);
nand U5990 (N_5990,N_4372,N_4866);
nand U5991 (N_5991,N_4611,N_4100);
nand U5992 (N_5992,N_4242,N_4793);
nor U5993 (N_5993,N_4095,N_4857);
nor U5994 (N_5994,N_4123,N_4454);
nor U5995 (N_5995,N_4060,N_4056);
xor U5996 (N_5996,N_4417,N_4285);
nand U5997 (N_5997,N_4247,N_4585);
nand U5998 (N_5998,N_4964,N_4213);
and U5999 (N_5999,N_4309,N_4380);
and U6000 (N_6000,N_5895,N_5962);
or U6001 (N_6001,N_5545,N_5898);
or U6002 (N_6002,N_5228,N_5498);
or U6003 (N_6003,N_5739,N_5517);
and U6004 (N_6004,N_5082,N_5721);
nor U6005 (N_6005,N_5409,N_5367);
xnor U6006 (N_6006,N_5324,N_5458);
and U6007 (N_6007,N_5877,N_5398);
nand U6008 (N_6008,N_5327,N_5651);
or U6009 (N_6009,N_5885,N_5953);
nor U6010 (N_6010,N_5337,N_5540);
nand U6011 (N_6011,N_5297,N_5930);
xnor U6012 (N_6012,N_5861,N_5014);
nor U6013 (N_6013,N_5243,N_5634);
or U6014 (N_6014,N_5581,N_5947);
nand U6015 (N_6015,N_5328,N_5235);
or U6016 (N_6016,N_5696,N_5810);
and U6017 (N_6017,N_5492,N_5219);
and U6018 (N_6018,N_5640,N_5864);
and U6019 (N_6019,N_5109,N_5035);
nand U6020 (N_6020,N_5795,N_5140);
nor U6021 (N_6021,N_5226,N_5848);
nor U6022 (N_6022,N_5553,N_5549);
or U6023 (N_6023,N_5858,N_5669);
or U6024 (N_6024,N_5387,N_5096);
and U6025 (N_6025,N_5695,N_5786);
xor U6026 (N_6026,N_5763,N_5736);
nand U6027 (N_6027,N_5589,N_5571);
and U6028 (N_6028,N_5712,N_5704);
or U6029 (N_6029,N_5240,N_5299);
and U6030 (N_6030,N_5595,N_5577);
xor U6031 (N_6031,N_5154,N_5605);
xor U6032 (N_6032,N_5175,N_5932);
and U6033 (N_6033,N_5342,N_5356);
and U6034 (N_6034,N_5438,N_5163);
nor U6035 (N_6035,N_5709,N_5705);
nor U6036 (N_6036,N_5307,N_5726);
nand U6037 (N_6037,N_5737,N_5127);
and U6038 (N_6038,N_5809,N_5227);
xnor U6039 (N_6039,N_5940,N_5206);
nor U6040 (N_6040,N_5701,N_5369);
nor U6041 (N_6041,N_5032,N_5754);
nor U6042 (N_6042,N_5828,N_5527);
or U6043 (N_6043,N_5902,N_5732);
nand U6044 (N_6044,N_5454,N_5482);
or U6045 (N_6045,N_5629,N_5178);
and U6046 (N_6046,N_5575,N_5740);
or U6047 (N_6047,N_5661,N_5167);
xnor U6048 (N_6048,N_5086,N_5650);
nor U6049 (N_6049,N_5434,N_5353);
and U6050 (N_6050,N_5120,N_5088);
nor U6051 (N_6051,N_5679,N_5280);
nand U6052 (N_6052,N_5218,N_5480);
or U6053 (N_6053,N_5223,N_5298);
nand U6054 (N_6054,N_5821,N_5474);
nor U6055 (N_6055,N_5863,N_5748);
xnor U6056 (N_6056,N_5804,N_5432);
nor U6057 (N_6057,N_5826,N_5066);
and U6058 (N_6058,N_5142,N_5027);
nor U6059 (N_6059,N_5785,N_5878);
or U6060 (N_6060,N_5245,N_5397);
nor U6061 (N_6061,N_5106,N_5720);
or U6062 (N_6062,N_5100,N_5759);
and U6063 (N_6063,N_5797,N_5293);
nand U6064 (N_6064,N_5666,N_5462);
nand U6065 (N_6065,N_5714,N_5807);
or U6066 (N_6066,N_5522,N_5355);
xnor U6067 (N_6067,N_5215,N_5113);
nand U6068 (N_6068,N_5242,N_5445);
xnor U6069 (N_6069,N_5415,N_5173);
and U6070 (N_6070,N_5915,N_5475);
nand U6071 (N_6071,N_5209,N_5083);
and U6072 (N_6072,N_5541,N_5539);
nand U6073 (N_6073,N_5772,N_5081);
nor U6074 (N_6074,N_5333,N_5039);
nor U6075 (N_6075,N_5444,N_5671);
nand U6076 (N_6076,N_5533,N_5285);
and U6077 (N_6077,N_5344,N_5429);
or U6078 (N_6078,N_5406,N_5188);
and U6079 (N_6079,N_5970,N_5631);
nand U6080 (N_6080,N_5197,N_5053);
and U6081 (N_6081,N_5182,N_5562);
or U6082 (N_6082,N_5788,N_5220);
nor U6083 (N_6083,N_5674,N_5870);
nor U6084 (N_6084,N_5017,N_5390);
nand U6085 (N_6085,N_5329,N_5708);
nor U6086 (N_6086,N_5395,N_5646);
xor U6087 (N_6087,N_5330,N_5055);
xor U6088 (N_6088,N_5413,N_5105);
xor U6089 (N_6089,N_5950,N_5831);
and U6090 (N_6090,N_5079,N_5937);
and U6091 (N_6091,N_5871,N_5888);
xor U6092 (N_6092,N_5874,N_5128);
xnor U6093 (N_6093,N_5452,N_5653);
xor U6094 (N_6094,N_5642,N_5798);
nor U6095 (N_6095,N_5530,N_5180);
and U6096 (N_6096,N_5838,N_5995);
xnor U6097 (N_6097,N_5208,N_5929);
nand U6098 (N_6098,N_5048,N_5352);
nand U6099 (N_6099,N_5762,N_5115);
xnor U6100 (N_6100,N_5384,N_5247);
and U6101 (N_6101,N_5546,N_5499);
nor U6102 (N_6102,N_5590,N_5857);
xor U6103 (N_6103,N_5946,N_5905);
nor U6104 (N_6104,N_5124,N_5588);
and U6105 (N_6105,N_5021,N_5570);
and U6106 (N_6106,N_5845,N_5987);
nand U6107 (N_6107,N_5891,N_5362);
nor U6108 (N_6108,N_5440,N_5442);
nor U6109 (N_6109,N_5951,N_5020);
nand U6110 (N_6110,N_5408,N_5345);
and U6111 (N_6111,N_5896,N_5814);
or U6112 (N_6112,N_5687,N_5407);
and U6113 (N_6113,N_5317,N_5465);
and U6114 (N_6114,N_5622,N_5808);
or U6115 (N_6115,N_5181,N_5820);
nor U6116 (N_6116,N_5998,N_5585);
or U6117 (N_6117,N_5711,N_5664);
or U6118 (N_6118,N_5271,N_5047);
and U6119 (N_6119,N_5824,N_5107);
xor U6120 (N_6120,N_5628,N_5999);
nor U6121 (N_6121,N_5718,N_5412);
xor U6122 (N_6122,N_5636,N_5806);
xor U6123 (N_6123,N_5556,N_5584);
nand U6124 (N_6124,N_5437,N_5090);
nand U6125 (N_6125,N_5359,N_5598);
or U6126 (N_6126,N_5567,N_5506);
xnor U6127 (N_6127,N_5370,N_5341);
or U6128 (N_6128,N_5051,N_5260);
nand U6129 (N_6129,N_5774,N_5684);
nand U6130 (N_6130,N_5006,N_5985);
nand U6131 (N_6131,N_5383,N_5641);
and U6132 (N_6132,N_5485,N_5016);
nor U6133 (N_6133,N_5520,N_5230);
and U6134 (N_6134,N_5665,N_5232);
and U6135 (N_6135,N_5548,N_5061);
nor U6136 (N_6136,N_5979,N_5967);
or U6137 (N_6137,N_5554,N_5859);
or U6138 (N_6138,N_5091,N_5672);
xor U6139 (N_6139,N_5289,N_5840);
or U6140 (N_6140,N_5514,N_5799);
nor U6141 (N_6141,N_5446,N_5033);
nor U6142 (N_6142,N_5168,N_5776);
nor U6143 (N_6143,N_5463,N_5277);
or U6144 (N_6144,N_5964,N_5213);
nand U6145 (N_6145,N_5073,N_5761);
and U6146 (N_6146,N_5210,N_5116);
xnor U6147 (N_6147,N_5880,N_5050);
or U6148 (N_6148,N_5497,N_5717);
xnor U6149 (N_6149,N_5501,N_5379);
nor U6150 (N_6150,N_5537,N_5259);
or U6151 (N_6151,N_5781,N_5371);
nand U6152 (N_6152,N_5723,N_5284);
nand U6153 (N_6153,N_5185,N_5682);
xnor U6154 (N_6154,N_5363,N_5368);
xnor U6155 (N_6155,N_5161,N_5319);
nor U6156 (N_6156,N_5153,N_5195);
nand U6157 (N_6157,N_5900,N_5275);
xnor U6158 (N_6158,N_5198,N_5426);
xor U6159 (N_6159,N_5262,N_5890);
or U6160 (N_6160,N_5155,N_5443);
xnor U6161 (N_6161,N_5816,N_5780);
xnor U6162 (N_6162,N_5270,N_5057);
nor U6163 (N_6163,N_5724,N_5493);
and U6164 (N_6164,N_5557,N_5743);
and U6165 (N_6165,N_5476,N_5959);
and U6166 (N_6166,N_5169,N_5117);
nor U6167 (N_6167,N_5678,N_5040);
or U6168 (N_6168,N_5852,N_5058);
or U6169 (N_6169,N_5677,N_5393);
or U6170 (N_6170,N_5403,N_5199);
or U6171 (N_6171,N_5886,N_5745);
nor U6172 (N_6172,N_5010,N_5749);
nand U6173 (N_6173,N_5157,N_5129);
nor U6174 (N_6174,N_5529,N_5996);
or U6175 (N_6175,N_5281,N_5414);
nor U6176 (N_6176,N_5236,N_5191);
or U6177 (N_6177,N_5734,N_5258);
xor U6178 (N_6178,N_5564,N_5075);
or U6179 (N_6179,N_5957,N_5361);
nor U6180 (N_6180,N_5494,N_5697);
nor U6181 (N_6181,N_5101,N_5680);
or U6182 (N_6182,N_5322,N_5618);
nand U6183 (N_6183,N_5908,N_5536);
nand U6184 (N_6184,N_5201,N_5619);
xor U6185 (N_6185,N_5688,N_5782);
or U6186 (N_6186,N_5958,N_5710);
or U6187 (N_6187,N_5893,N_5867);
xnor U6188 (N_6188,N_5441,N_5378);
xnor U6189 (N_6189,N_5046,N_5971);
xnor U6190 (N_6190,N_5350,N_5349);
nand U6191 (N_6191,N_5733,N_5511);
xnor U6192 (N_6192,N_5818,N_5875);
and U6193 (N_6193,N_5388,N_5925);
or U6194 (N_6194,N_5767,N_5612);
nand U6195 (N_6195,N_5941,N_5757);
nor U6196 (N_6196,N_5843,N_5029);
and U6197 (N_6197,N_5347,N_5062);
xnor U6198 (N_6198,N_5899,N_5574);
nor U6199 (N_6199,N_5800,N_5421);
or U6200 (N_6200,N_5351,N_5264);
nand U6201 (N_6201,N_5862,N_5849);
xor U6202 (N_6202,N_5273,N_5292);
xor U6203 (N_6203,N_5431,N_5791);
nand U6204 (N_6204,N_5756,N_5645);
nand U6205 (N_6205,N_5147,N_5760);
nand U6206 (N_6206,N_5423,N_5894);
nor U6207 (N_6207,N_5531,N_5360);
and U6208 (N_6208,N_5254,N_5248);
and U6209 (N_6209,N_5239,N_5609);
nand U6210 (N_6210,N_5841,N_5479);
nor U6211 (N_6211,N_5794,N_5917);
xor U6212 (N_6212,N_5560,N_5783);
and U6213 (N_6213,N_5948,N_5578);
and U6214 (N_6214,N_5008,N_5011);
or U6215 (N_6215,N_5166,N_5579);
and U6216 (N_6216,N_5960,N_5968);
xnor U6217 (N_6217,N_5662,N_5775);
nand U6218 (N_6218,N_5435,N_5114);
and U6219 (N_6219,N_5741,N_5722);
or U6220 (N_6220,N_5447,N_5138);
nand U6221 (N_6221,N_5150,N_5657);
nand U6222 (N_6222,N_5045,N_5401);
nand U6223 (N_6223,N_5969,N_5026);
xor U6224 (N_6224,N_5563,N_5792);
and U6225 (N_6225,N_5325,N_5933);
nor U6226 (N_6226,N_5132,N_5993);
xor U6227 (N_6227,N_5832,N_5212);
nand U6228 (N_6228,N_5059,N_5921);
and U6229 (N_6229,N_5922,N_5850);
and U6230 (N_6230,N_5707,N_5945);
nand U6231 (N_6231,N_5939,N_5282);
and U6232 (N_6232,N_5827,N_5009);
xnor U6233 (N_6233,N_5255,N_5765);
or U6234 (N_6234,N_5099,N_5131);
xor U6235 (N_6235,N_5448,N_5658);
nand U6236 (N_6236,N_5112,N_5882);
nand U6237 (N_6237,N_5510,N_5813);
xor U6238 (N_6238,N_5747,N_5310);
xor U6239 (N_6239,N_5183,N_5145);
nor U6240 (N_6240,N_5624,N_5189);
xor U6241 (N_6241,N_5716,N_5943);
and U6242 (N_6242,N_5508,N_5685);
xor U6243 (N_6243,N_5121,N_5477);
xnor U6244 (N_6244,N_5233,N_5990);
nand U6245 (N_6245,N_5391,N_5013);
and U6246 (N_6246,N_5926,N_5309);
nand U6247 (N_6247,N_5534,N_5315);
and U6248 (N_6248,N_5135,N_5043);
xnor U6249 (N_6249,N_5952,N_5071);
xor U6250 (N_6250,N_5509,N_5250);
and U6251 (N_6251,N_5222,N_5686);
and U6252 (N_6252,N_5552,N_5382);
and U6253 (N_6253,N_5502,N_5405);
nor U6254 (N_6254,N_5216,N_5399);
and U6255 (N_6255,N_5323,N_5991);
nand U6256 (N_6256,N_5089,N_5287);
or U6257 (N_6257,N_5374,N_5093);
nand U6258 (N_6258,N_5326,N_5253);
or U6259 (N_6259,N_5110,N_5881);
xnor U6260 (N_6260,N_5072,N_5644);
nand U6261 (N_6261,N_5822,N_5229);
and U6262 (N_6262,N_5654,N_5565);
xnor U6263 (N_6263,N_5162,N_5012);
or U6264 (N_6264,N_5944,N_5856);
xor U6265 (N_6265,N_5730,N_5879);
nand U6266 (N_6266,N_5500,N_5972);
nand U6267 (N_6267,N_5989,N_5825);
xor U6268 (N_6268,N_5424,N_5770);
nand U6269 (N_6269,N_5519,N_5267);
and U6270 (N_6270,N_5266,N_5603);
xor U6271 (N_6271,N_5702,N_5528);
or U6272 (N_6272,N_5637,N_5551);
or U6273 (N_6273,N_5425,N_5366);
and U6274 (N_6274,N_5835,N_5975);
nor U6275 (N_6275,N_5468,N_5647);
xor U6276 (N_6276,N_5675,N_5249);
nor U6277 (N_6277,N_5331,N_5296);
nor U6278 (N_6278,N_5801,N_5692);
and U6279 (N_6279,N_5638,N_5942);
or U6280 (N_6280,N_5257,N_5600);
and U6281 (N_6281,N_5887,N_5316);
nand U6282 (N_6282,N_5486,N_5559);
nand U6283 (N_6283,N_5005,N_5586);
or U6284 (N_6284,N_5044,N_5728);
nand U6285 (N_6285,N_5400,N_5418);
nor U6286 (N_6286,N_5211,N_5436);
or U6287 (N_6287,N_5614,N_5773);
or U6288 (N_6288,N_5022,N_5673);
nand U6289 (N_6289,N_5532,N_5752);
or U6290 (N_6290,N_5580,N_5144);
or U6291 (N_6291,N_5286,N_5340);
or U6292 (N_6292,N_5394,N_5676);
xor U6293 (N_6293,N_5847,N_5504);
nor U6294 (N_6294,N_5516,N_5313);
xnor U6295 (N_6295,N_5256,N_5924);
xor U6296 (N_6296,N_5385,N_5689);
and U6297 (N_6297,N_5478,N_5025);
or U6298 (N_6298,N_5171,N_5063);
and U6299 (N_6299,N_5291,N_5335);
nand U6300 (N_6300,N_5419,N_5217);
nor U6301 (N_6301,N_5984,N_5918);
and U6302 (N_6302,N_5148,N_5608);
or U6303 (N_6303,N_5346,N_5583);
or U6304 (N_6304,N_5855,N_5837);
or U6305 (N_6305,N_5034,N_5513);
or U6306 (N_6306,N_5451,N_5238);
nor U6307 (N_6307,N_5372,N_5049);
and U6308 (N_6308,N_5302,N_5572);
nand U6309 (N_6309,N_5244,N_5873);
xnor U6310 (N_6310,N_5237,N_5496);
nor U6311 (N_6311,N_5833,N_5623);
nor U6312 (N_6312,N_5422,N_5002);
or U6313 (N_6313,N_5141,N_5417);
nand U6314 (N_6314,N_5321,N_5865);
or U6315 (N_6315,N_5036,N_5803);
and U6316 (N_6316,N_5184,N_5146);
xnor U6317 (N_6317,N_5334,N_5376);
xnor U6318 (N_6318,N_5410,N_5587);
and U6319 (N_6319,N_5521,N_5526);
nand U6320 (N_6320,N_5544,N_5495);
and U6321 (N_6321,N_5070,N_5118);
nand U6322 (N_6322,N_5593,N_5965);
or U6323 (N_6323,N_5386,N_5300);
or U6324 (N_6324,N_5023,N_5746);
nor U6325 (N_6325,N_5074,N_5224);
xnor U6326 (N_6326,N_5784,N_5077);
and U6327 (N_6327,N_5123,N_5611);
xnor U6328 (N_6328,N_5906,N_5904);
nor U6329 (N_6329,N_5098,N_5613);
or U6330 (N_6330,N_5052,N_5977);
or U6331 (N_6331,N_5320,N_5076);
nor U6332 (N_6332,N_5420,N_5817);
nand U6333 (N_6333,N_5272,N_5992);
or U6334 (N_6334,N_5294,N_5713);
nand U6335 (N_6335,N_5591,N_5796);
nor U6336 (N_6336,N_5974,N_5963);
and U6337 (N_6337,N_5568,N_5318);
or U6338 (N_6338,N_5851,N_5288);
nor U6339 (N_6339,N_5364,N_5469);
nand U6340 (N_6340,N_5177,N_5823);
or U6341 (N_6341,N_5819,N_5876);
nor U6342 (N_6342,N_5159,N_5805);
and U6343 (N_6343,N_5137,N_5706);
nand U6344 (N_6344,N_5719,N_5164);
nand U6345 (N_6345,N_5981,N_5119);
nor U6346 (N_6346,N_5449,N_5471);
or U6347 (N_6347,N_5308,N_5193);
and U6348 (N_6348,N_5986,N_5727);
or U6349 (N_6349,N_5815,N_5225);
and U6350 (N_6350,N_5909,N_5234);
nor U6351 (N_6351,N_5170,N_5165);
and U6352 (N_6352,N_5778,N_5200);
xor U6353 (N_6353,N_5103,N_5381);
or U6354 (N_6354,N_5396,N_5203);
nor U6355 (N_6355,N_5955,N_5648);
nor U6356 (N_6356,N_5742,N_5670);
nor U6357 (N_6357,N_5505,N_5274);
nand U6358 (N_6358,N_5483,N_5625);
nand U6359 (N_6359,N_5457,N_5453);
nand U6360 (N_6360,N_5639,N_5758);
and U6361 (N_6361,N_5404,N_5931);
xnor U6362 (N_6362,N_5868,N_5261);
and U6363 (N_6363,N_5683,N_5617);
nand U6364 (N_6364,N_5460,N_5488);
nand U6365 (N_6365,N_5087,N_5094);
xnor U6366 (N_6366,N_5455,N_5111);
and U6367 (N_6367,N_5897,N_5018);
and U6368 (N_6368,N_5630,N_5392);
xor U6369 (N_6369,N_5542,N_5860);
nand U6370 (N_6370,N_5427,N_5295);
xnor U6371 (N_6371,N_5846,N_5550);
nand U6372 (N_6372,N_5343,N_5842);
nor U6373 (N_6373,N_5064,N_5263);
or U6374 (N_6374,N_5652,N_5973);
xor U6375 (N_6375,N_5901,N_5192);
nor U6376 (N_6376,N_5430,N_5779);
nand U6377 (N_6377,N_5607,N_5204);
nor U6378 (N_6378,N_5348,N_5632);
nor U6379 (N_6379,N_5470,N_5126);
nor U6380 (N_6380,N_5699,N_5616);
and U6381 (N_6381,N_5019,N_5467);
nor U6382 (N_6382,N_5660,N_5411);
xnor U6383 (N_6383,N_5750,N_5731);
nand U6384 (N_6384,N_5172,N_5729);
xor U6385 (N_6385,N_5276,N_5771);
nor U6386 (N_6386,N_5473,N_5949);
xor U6387 (N_6387,N_5836,N_5490);
and U6388 (N_6388,N_5416,N_5872);
and U6389 (N_6389,N_5934,N_5518);
nand U6390 (N_6390,N_5068,N_5663);
nor U6391 (N_6391,N_5635,N_5031);
or U6392 (N_6392,N_5301,N_5283);
nand U6393 (N_6393,N_5489,N_5853);
nor U6394 (N_6394,N_5251,N_5997);
nor U6395 (N_6395,N_5194,N_5214);
xnor U6396 (N_6396,N_5186,N_5938);
or U6397 (N_6397,N_5621,N_5976);
nor U6398 (N_6398,N_5187,N_5994);
xnor U6399 (N_6399,N_5911,N_5919);
nand U6400 (N_6400,N_5834,N_5304);
nor U6401 (N_6401,N_5428,N_5980);
xor U6402 (N_6402,N_5125,N_5681);
xor U6403 (N_6403,N_5656,N_5205);
and U6404 (N_6404,N_5507,N_5491);
or U6405 (N_6405,N_5755,N_5030);
and U6406 (N_6406,N_5555,N_5332);
and U6407 (N_6407,N_5311,N_5789);
nor U6408 (N_6408,N_5561,N_5599);
or U6409 (N_6409,N_5156,N_5606);
xor U6410 (N_6410,N_5389,N_5202);
and U6411 (N_6411,N_5725,N_5978);
nand U6412 (N_6412,N_5484,N_5015);
and U6413 (N_6413,N_5715,N_5450);
or U6414 (N_6414,N_5582,N_5339);
and U6415 (N_6415,N_5854,N_5080);
nor U6416 (N_6416,N_5889,N_5839);
xor U6417 (N_6417,N_5174,N_5338);
and U6418 (N_6418,N_5380,N_5265);
nand U6419 (N_6419,N_5907,N_5538);
nand U6420 (N_6420,N_5768,N_5158);
or U6421 (N_6421,N_5190,N_5626);
nor U6422 (N_6422,N_5751,N_5097);
xor U6423 (N_6423,N_5525,N_5503);
xnor U6424 (N_6424,N_5130,N_5092);
nor U6425 (N_6425,N_5954,N_5573);
nand U6426 (N_6426,N_5472,N_5655);
nor U6427 (N_6427,N_5844,N_5830);
nor U6428 (N_6428,N_5983,N_5354);
and U6429 (N_6429,N_5459,N_5179);
nor U6430 (N_6430,N_5569,N_5602);
nor U6431 (N_6431,N_5693,N_5936);
and U6432 (N_6432,N_5433,N_5143);
and U6433 (N_6433,N_5056,N_5054);
nor U6434 (N_6434,N_5306,N_5892);
or U6435 (N_6435,N_5176,N_5104);
xor U6436 (N_6436,N_5003,N_5535);
and U6437 (N_6437,N_5037,N_5966);
xor U6438 (N_6438,N_5481,N_5790);
nor U6439 (N_6439,N_5793,N_5956);
or U6440 (N_6440,N_5884,N_5903);
xnor U6441 (N_6441,N_5439,N_5649);
or U6442 (N_6442,N_5136,N_5866);
nand U6443 (N_6443,N_5735,N_5547);
and U6444 (N_6444,N_5596,N_5278);
or U6445 (N_6445,N_5038,N_5829);
nand U6446 (N_6446,N_5357,N_5916);
and U6447 (N_6447,N_5358,N_5461);
nand U6448 (N_6448,N_5633,N_5512);
or U6449 (N_6449,N_5961,N_5102);
or U6450 (N_6450,N_5812,N_5777);
or U6451 (N_6451,N_5523,N_5028);
xor U6452 (N_6452,N_5221,N_5627);
and U6453 (N_6453,N_5268,N_5912);
nor U6454 (N_6454,N_5615,N_5269);
nand U6455 (N_6455,N_5466,N_5085);
nand U6456 (N_6456,N_5377,N_5004);
xnor U6457 (N_6457,N_5869,N_5700);
and U6458 (N_6458,N_5365,N_5620);
or U6459 (N_6459,N_5303,N_5659);
and U6460 (N_6460,N_5067,N_5007);
xnor U6461 (N_6461,N_5668,N_5151);
nand U6462 (N_6462,N_5312,N_5766);
xor U6463 (N_6463,N_5456,N_5095);
nand U6464 (N_6464,N_5764,N_5988);
or U6465 (N_6465,N_5576,N_5065);
or U6466 (N_6466,N_5069,N_5914);
and U6467 (N_6467,N_5060,N_5769);
xor U6468 (N_6468,N_5923,N_5935);
nand U6469 (N_6469,N_5515,N_5375);
and U6470 (N_6470,N_5122,N_5290);
nor U6471 (N_6471,N_5787,N_5133);
nand U6472 (N_6472,N_5982,N_5078);
xor U6473 (N_6473,N_5643,N_5691);
or U6474 (N_6474,N_5910,N_5152);
and U6475 (N_6475,N_5305,N_5524);
or U6476 (N_6476,N_5927,N_5883);
or U6477 (N_6477,N_5913,N_5703);
nor U6478 (N_6478,N_5802,N_5231);
and U6479 (N_6479,N_5597,N_5690);
nand U6480 (N_6480,N_5108,N_5241);
and U6481 (N_6481,N_5601,N_5314);
or U6482 (N_6482,N_5160,N_5698);
nand U6483 (N_6483,N_5279,N_5373);
and U6484 (N_6484,N_5134,N_5139);
xnor U6485 (N_6485,N_5694,N_5041);
or U6486 (N_6486,N_5592,N_5001);
xnor U6487 (N_6487,N_5610,N_5402);
nor U6488 (N_6488,N_5594,N_5667);
nand U6489 (N_6489,N_5811,N_5149);
nand U6490 (N_6490,N_5196,N_5042);
or U6491 (N_6491,N_5738,N_5336);
and U6492 (N_6492,N_5928,N_5024);
nand U6493 (N_6493,N_5487,N_5566);
nand U6494 (N_6494,N_5000,N_5604);
nand U6495 (N_6495,N_5207,N_5464);
nor U6496 (N_6496,N_5753,N_5744);
and U6497 (N_6497,N_5558,N_5543);
nand U6498 (N_6498,N_5246,N_5252);
and U6499 (N_6499,N_5084,N_5920);
nor U6500 (N_6500,N_5802,N_5220);
nand U6501 (N_6501,N_5099,N_5856);
nor U6502 (N_6502,N_5772,N_5214);
nor U6503 (N_6503,N_5055,N_5395);
or U6504 (N_6504,N_5903,N_5604);
xor U6505 (N_6505,N_5650,N_5974);
nor U6506 (N_6506,N_5705,N_5620);
nor U6507 (N_6507,N_5936,N_5573);
xnor U6508 (N_6508,N_5546,N_5395);
nand U6509 (N_6509,N_5616,N_5145);
nand U6510 (N_6510,N_5053,N_5266);
or U6511 (N_6511,N_5256,N_5680);
and U6512 (N_6512,N_5680,N_5777);
xnor U6513 (N_6513,N_5370,N_5951);
and U6514 (N_6514,N_5753,N_5119);
nand U6515 (N_6515,N_5753,N_5891);
and U6516 (N_6516,N_5719,N_5395);
and U6517 (N_6517,N_5010,N_5815);
and U6518 (N_6518,N_5243,N_5828);
and U6519 (N_6519,N_5348,N_5428);
or U6520 (N_6520,N_5565,N_5193);
xor U6521 (N_6521,N_5096,N_5715);
and U6522 (N_6522,N_5548,N_5016);
and U6523 (N_6523,N_5824,N_5644);
and U6524 (N_6524,N_5551,N_5850);
xnor U6525 (N_6525,N_5345,N_5365);
and U6526 (N_6526,N_5792,N_5423);
or U6527 (N_6527,N_5386,N_5616);
nand U6528 (N_6528,N_5681,N_5061);
xnor U6529 (N_6529,N_5801,N_5742);
nor U6530 (N_6530,N_5109,N_5213);
or U6531 (N_6531,N_5011,N_5596);
nor U6532 (N_6532,N_5884,N_5919);
or U6533 (N_6533,N_5043,N_5540);
nor U6534 (N_6534,N_5042,N_5771);
and U6535 (N_6535,N_5871,N_5156);
xnor U6536 (N_6536,N_5175,N_5036);
nand U6537 (N_6537,N_5453,N_5687);
or U6538 (N_6538,N_5079,N_5361);
or U6539 (N_6539,N_5649,N_5430);
nand U6540 (N_6540,N_5001,N_5064);
and U6541 (N_6541,N_5112,N_5664);
or U6542 (N_6542,N_5737,N_5295);
xnor U6543 (N_6543,N_5997,N_5458);
or U6544 (N_6544,N_5626,N_5894);
xnor U6545 (N_6545,N_5829,N_5276);
xnor U6546 (N_6546,N_5947,N_5278);
nor U6547 (N_6547,N_5596,N_5366);
xnor U6548 (N_6548,N_5342,N_5754);
nor U6549 (N_6549,N_5532,N_5627);
or U6550 (N_6550,N_5682,N_5913);
nand U6551 (N_6551,N_5974,N_5395);
xnor U6552 (N_6552,N_5704,N_5141);
nor U6553 (N_6553,N_5887,N_5883);
nor U6554 (N_6554,N_5272,N_5176);
and U6555 (N_6555,N_5633,N_5957);
nor U6556 (N_6556,N_5188,N_5481);
nor U6557 (N_6557,N_5629,N_5608);
xnor U6558 (N_6558,N_5621,N_5469);
nor U6559 (N_6559,N_5018,N_5246);
or U6560 (N_6560,N_5069,N_5682);
xor U6561 (N_6561,N_5817,N_5332);
and U6562 (N_6562,N_5953,N_5164);
and U6563 (N_6563,N_5317,N_5704);
nand U6564 (N_6564,N_5167,N_5875);
or U6565 (N_6565,N_5473,N_5315);
and U6566 (N_6566,N_5477,N_5963);
and U6567 (N_6567,N_5841,N_5437);
and U6568 (N_6568,N_5902,N_5828);
and U6569 (N_6569,N_5592,N_5711);
nor U6570 (N_6570,N_5606,N_5201);
and U6571 (N_6571,N_5864,N_5683);
nor U6572 (N_6572,N_5779,N_5633);
nor U6573 (N_6573,N_5361,N_5034);
nor U6574 (N_6574,N_5045,N_5957);
and U6575 (N_6575,N_5285,N_5967);
nand U6576 (N_6576,N_5547,N_5215);
nand U6577 (N_6577,N_5758,N_5606);
and U6578 (N_6578,N_5645,N_5455);
or U6579 (N_6579,N_5211,N_5934);
or U6580 (N_6580,N_5672,N_5531);
and U6581 (N_6581,N_5347,N_5318);
nor U6582 (N_6582,N_5236,N_5549);
and U6583 (N_6583,N_5330,N_5465);
xnor U6584 (N_6584,N_5240,N_5562);
or U6585 (N_6585,N_5216,N_5954);
xnor U6586 (N_6586,N_5715,N_5426);
nand U6587 (N_6587,N_5972,N_5417);
nand U6588 (N_6588,N_5335,N_5301);
xnor U6589 (N_6589,N_5613,N_5422);
and U6590 (N_6590,N_5558,N_5052);
nand U6591 (N_6591,N_5519,N_5487);
nand U6592 (N_6592,N_5814,N_5656);
nor U6593 (N_6593,N_5780,N_5791);
nor U6594 (N_6594,N_5089,N_5477);
nor U6595 (N_6595,N_5179,N_5327);
and U6596 (N_6596,N_5945,N_5364);
xnor U6597 (N_6597,N_5980,N_5556);
nand U6598 (N_6598,N_5543,N_5028);
or U6599 (N_6599,N_5708,N_5697);
and U6600 (N_6600,N_5568,N_5890);
and U6601 (N_6601,N_5079,N_5423);
and U6602 (N_6602,N_5014,N_5395);
nor U6603 (N_6603,N_5444,N_5482);
nand U6604 (N_6604,N_5958,N_5273);
nor U6605 (N_6605,N_5053,N_5484);
and U6606 (N_6606,N_5694,N_5660);
nand U6607 (N_6607,N_5045,N_5157);
and U6608 (N_6608,N_5458,N_5838);
and U6609 (N_6609,N_5126,N_5864);
nand U6610 (N_6610,N_5676,N_5180);
and U6611 (N_6611,N_5242,N_5732);
and U6612 (N_6612,N_5610,N_5419);
or U6613 (N_6613,N_5727,N_5339);
or U6614 (N_6614,N_5451,N_5152);
nor U6615 (N_6615,N_5888,N_5337);
and U6616 (N_6616,N_5147,N_5772);
and U6617 (N_6617,N_5548,N_5888);
or U6618 (N_6618,N_5773,N_5044);
or U6619 (N_6619,N_5343,N_5841);
and U6620 (N_6620,N_5254,N_5055);
nand U6621 (N_6621,N_5819,N_5256);
and U6622 (N_6622,N_5037,N_5556);
and U6623 (N_6623,N_5222,N_5846);
xor U6624 (N_6624,N_5347,N_5389);
and U6625 (N_6625,N_5664,N_5407);
nand U6626 (N_6626,N_5333,N_5939);
nand U6627 (N_6627,N_5574,N_5578);
xnor U6628 (N_6628,N_5389,N_5472);
xor U6629 (N_6629,N_5273,N_5044);
or U6630 (N_6630,N_5095,N_5148);
or U6631 (N_6631,N_5298,N_5400);
nor U6632 (N_6632,N_5930,N_5920);
and U6633 (N_6633,N_5051,N_5783);
nor U6634 (N_6634,N_5586,N_5379);
xor U6635 (N_6635,N_5082,N_5042);
nand U6636 (N_6636,N_5230,N_5580);
xor U6637 (N_6637,N_5055,N_5401);
nand U6638 (N_6638,N_5190,N_5231);
nor U6639 (N_6639,N_5688,N_5031);
and U6640 (N_6640,N_5382,N_5290);
xnor U6641 (N_6641,N_5558,N_5784);
and U6642 (N_6642,N_5559,N_5433);
or U6643 (N_6643,N_5557,N_5754);
nor U6644 (N_6644,N_5183,N_5634);
nor U6645 (N_6645,N_5707,N_5741);
xnor U6646 (N_6646,N_5106,N_5403);
or U6647 (N_6647,N_5286,N_5515);
and U6648 (N_6648,N_5638,N_5455);
or U6649 (N_6649,N_5646,N_5002);
xor U6650 (N_6650,N_5295,N_5913);
and U6651 (N_6651,N_5420,N_5064);
and U6652 (N_6652,N_5066,N_5675);
nor U6653 (N_6653,N_5883,N_5751);
xnor U6654 (N_6654,N_5846,N_5970);
or U6655 (N_6655,N_5694,N_5379);
or U6656 (N_6656,N_5466,N_5277);
xnor U6657 (N_6657,N_5262,N_5545);
and U6658 (N_6658,N_5920,N_5626);
or U6659 (N_6659,N_5512,N_5164);
xor U6660 (N_6660,N_5528,N_5881);
nand U6661 (N_6661,N_5881,N_5844);
or U6662 (N_6662,N_5226,N_5419);
and U6663 (N_6663,N_5692,N_5699);
or U6664 (N_6664,N_5710,N_5246);
or U6665 (N_6665,N_5640,N_5548);
and U6666 (N_6666,N_5840,N_5246);
or U6667 (N_6667,N_5979,N_5571);
or U6668 (N_6668,N_5603,N_5926);
and U6669 (N_6669,N_5833,N_5238);
and U6670 (N_6670,N_5986,N_5595);
or U6671 (N_6671,N_5817,N_5549);
nor U6672 (N_6672,N_5469,N_5533);
nor U6673 (N_6673,N_5895,N_5500);
or U6674 (N_6674,N_5784,N_5912);
nand U6675 (N_6675,N_5855,N_5614);
or U6676 (N_6676,N_5762,N_5408);
or U6677 (N_6677,N_5602,N_5869);
nor U6678 (N_6678,N_5898,N_5662);
nand U6679 (N_6679,N_5846,N_5044);
nand U6680 (N_6680,N_5118,N_5625);
xnor U6681 (N_6681,N_5254,N_5157);
nand U6682 (N_6682,N_5943,N_5813);
and U6683 (N_6683,N_5573,N_5346);
xnor U6684 (N_6684,N_5256,N_5912);
and U6685 (N_6685,N_5744,N_5377);
xnor U6686 (N_6686,N_5525,N_5066);
nor U6687 (N_6687,N_5805,N_5235);
xor U6688 (N_6688,N_5491,N_5315);
xor U6689 (N_6689,N_5064,N_5282);
xor U6690 (N_6690,N_5823,N_5082);
xnor U6691 (N_6691,N_5797,N_5873);
nor U6692 (N_6692,N_5007,N_5032);
and U6693 (N_6693,N_5899,N_5373);
nand U6694 (N_6694,N_5472,N_5803);
nand U6695 (N_6695,N_5066,N_5147);
nor U6696 (N_6696,N_5545,N_5371);
or U6697 (N_6697,N_5908,N_5120);
and U6698 (N_6698,N_5164,N_5657);
xor U6699 (N_6699,N_5997,N_5606);
and U6700 (N_6700,N_5476,N_5410);
nor U6701 (N_6701,N_5842,N_5428);
and U6702 (N_6702,N_5923,N_5656);
and U6703 (N_6703,N_5699,N_5169);
xnor U6704 (N_6704,N_5478,N_5826);
nand U6705 (N_6705,N_5471,N_5860);
or U6706 (N_6706,N_5549,N_5251);
nand U6707 (N_6707,N_5214,N_5033);
nor U6708 (N_6708,N_5179,N_5876);
nor U6709 (N_6709,N_5332,N_5878);
nor U6710 (N_6710,N_5526,N_5536);
nor U6711 (N_6711,N_5229,N_5928);
nor U6712 (N_6712,N_5124,N_5869);
nand U6713 (N_6713,N_5103,N_5535);
nand U6714 (N_6714,N_5439,N_5746);
and U6715 (N_6715,N_5298,N_5221);
and U6716 (N_6716,N_5656,N_5669);
nor U6717 (N_6717,N_5798,N_5956);
and U6718 (N_6718,N_5622,N_5680);
and U6719 (N_6719,N_5345,N_5752);
xnor U6720 (N_6720,N_5910,N_5177);
and U6721 (N_6721,N_5631,N_5186);
or U6722 (N_6722,N_5868,N_5782);
xnor U6723 (N_6723,N_5630,N_5086);
xnor U6724 (N_6724,N_5606,N_5114);
nor U6725 (N_6725,N_5034,N_5137);
nand U6726 (N_6726,N_5521,N_5429);
and U6727 (N_6727,N_5936,N_5075);
and U6728 (N_6728,N_5958,N_5051);
or U6729 (N_6729,N_5944,N_5188);
or U6730 (N_6730,N_5069,N_5304);
and U6731 (N_6731,N_5702,N_5027);
nor U6732 (N_6732,N_5171,N_5475);
nand U6733 (N_6733,N_5523,N_5770);
and U6734 (N_6734,N_5232,N_5285);
xor U6735 (N_6735,N_5132,N_5549);
xnor U6736 (N_6736,N_5385,N_5305);
or U6737 (N_6737,N_5036,N_5835);
nand U6738 (N_6738,N_5588,N_5018);
nand U6739 (N_6739,N_5153,N_5085);
nor U6740 (N_6740,N_5527,N_5738);
and U6741 (N_6741,N_5727,N_5342);
and U6742 (N_6742,N_5305,N_5522);
nand U6743 (N_6743,N_5544,N_5109);
xnor U6744 (N_6744,N_5740,N_5542);
nand U6745 (N_6745,N_5707,N_5397);
nand U6746 (N_6746,N_5379,N_5109);
and U6747 (N_6747,N_5803,N_5137);
and U6748 (N_6748,N_5827,N_5015);
nor U6749 (N_6749,N_5694,N_5611);
or U6750 (N_6750,N_5544,N_5053);
nor U6751 (N_6751,N_5799,N_5788);
nand U6752 (N_6752,N_5842,N_5826);
xnor U6753 (N_6753,N_5769,N_5530);
and U6754 (N_6754,N_5151,N_5369);
or U6755 (N_6755,N_5137,N_5308);
or U6756 (N_6756,N_5631,N_5513);
xor U6757 (N_6757,N_5682,N_5425);
nor U6758 (N_6758,N_5407,N_5643);
or U6759 (N_6759,N_5137,N_5276);
xnor U6760 (N_6760,N_5272,N_5005);
nor U6761 (N_6761,N_5091,N_5562);
and U6762 (N_6762,N_5327,N_5482);
nor U6763 (N_6763,N_5448,N_5443);
and U6764 (N_6764,N_5980,N_5313);
nor U6765 (N_6765,N_5654,N_5061);
nor U6766 (N_6766,N_5250,N_5100);
and U6767 (N_6767,N_5216,N_5058);
and U6768 (N_6768,N_5460,N_5094);
nand U6769 (N_6769,N_5191,N_5656);
or U6770 (N_6770,N_5547,N_5468);
nand U6771 (N_6771,N_5989,N_5126);
xnor U6772 (N_6772,N_5825,N_5107);
or U6773 (N_6773,N_5770,N_5577);
or U6774 (N_6774,N_5673,N_5064);
nand U6775 (N_6775,N_5676,N_5017);
or U6776 (N_6776,N_5584,N_5008);
nand U6777 (N_6777,N_5181,N_5644);
xor U6778 (N_6778,N_5362,N_5281);
nor U6779 (N_6779,N_5837,N_5422);
nor U6780 (N_6780,N_5513,N_5897);
and U6781 (N_6781,N_5888,N_5575);
or U6782 (N_6782,N_5856,N_5627);
or U6783 (N_6783,N_5040,N_5101);
and U6784 (N_6784,N_5814,N_5922);
nand U6785 (N_6785,N_5068,N_5964);
nor U6786 (N_6786,N_5990,N_5841);
nor U6787 (N_6787,N_5149,N_5203);
nand U6788 (N_6788,N_5288,N_5335);
and U6789 (N_6789,N_5160,N_5348);
or U6790 (N_6790,N_5123,N_5033);
and U6791 (N_6791,N_5511,N_5514);
or U6792 (N_6792,N_5151,N_5039);
nand U6793 (N_6793,N_5306,N_5469);
nor U6794 (N_6794,N_5234,N_5556);
and U6795 (N_6795,N_5753,N_5666);
nor U6796 (N_6796,N_5676,N_5872);
nand U6797 (N_6797,N_5597,N_5442);
and U6798 (N_6798,N_5284,N_5506);
and U6799 (N_6799,N_5969,N_5554);
and U6800 (N_6800,N_5854,N_5551);
and U6801 (N_6801,N_5239,N_5584);
or U6802 (N_6802,N_5093,N_5917);
and U6803 (N_6803,N_5220,N_5628);
and U6804 (N_6804,N_5495,N_5937);
xor U6805 (N_6805,N_5134,N_5823);
nor U6806 (N_6806,N_5084,N_5799);
nand U6807 (N_6807,N_5449,N_5414);
nand U6808 (N_6808,N_5583,N_5407);
or U6809 (N_6809,N_5475,N_5424);
nand U6810 (N_6810,N_5319,N_5720);
nand U6811 (N_6811,N_5394,N_5117);
nand U6812 (N_6812,N_5276,N_5176);
nand U6813 (N_6813,N_5272,N_5368);
and U6814 (N_6814,N_5517,N_5268);
nand U6815 (N_6815,N_5690,N_5282);
nand U6816 (N_6816,N_5478,N_5810);
and U6817 (N_6817,N_5390,N_5737);
nor U6818 (N_6818,N_5261,N_5521);
and U6819 (N_6819,N_5452,N_5414);
or U6820 (N_6820,N_5543,N_5866);
or U6821 (N_6821,N_5968,N_5010);
and U6822 (N_6822,N_5930,N_5342);
nor U6823 (N_6823,N_5378,N_5340);
or U6824 (N_6824,N_5916,N_5914);
or U6825 (N_6825,N_5593,N_5714);
and U6826 (N_6826,N_5689,N_5626);
and U6827 (N_6827,N_5901,N_5445);
nand U6828 (N_6828,N_5222,N_5883);
nand U6829 (N_6829,N_5699,N_5695);
xnor U6830 (N_6830,N_5490,N_5382);
and U6831 (N_6831,N_5740,N_5182);
nand U6832 (N_6832,N_5435,N_5622);
or U6833 (N_6833,N_5868,N_5376);
and U6834 (N_6834,N_5827,N_5060);
nand U6835 (N_6835,N_5366,N_5195);
or U6836 (N_6836,N_5997,N_5664);
nand U6837 (N_6837,N_5427,N_5312);
and U6838 (N_6838,N_5480,N_5245);
nor U6839 (N_6839,N_5969,N_5965);
nand U6840 (N_6840,N_5979,N_5292);
nand U6841 (N_6841,N_5453,N_5811);
xor U6842 (N_6842,N_5967,N_5186);
and U6843 (N_6843,N_5150,N_5464);
nor U6844 (N_6844,N_5126,N_5658);
xor U6845 (N_6845,N_5898,N_5916);
xnor U6846 (N_6846,N_5507,N_5261);
nor U6847 (N_6847,N_5302,N_5765);
xnor U6848 (N_6848,N_5003,N_5970);
xnor U6849 (N_6849,N_5494,N_5513);
and U6850 (N_6850,N_5776,N_5056);
xnor U6851 (N_6851,N_5039,N_5161);
nand U6852 (N_6852,N_5022,N_5741);
and U6853 (N_6853,N_5085,N_5504);
nand U6854 (N_6854,N_5835,N_5760);
nor U6855 (N_6855,N_5722,N_5579);
xor U6856 (N_6856,N_5304,N_5542);
nand U6857 (N_6857,N_5485,N_5875);
or U6858 (N_6858,N_5497,N_5317);
nor U6859 (N_6859,N_5585,N_5564);
nor U6860 (N_6860,N_5379,N_5730);
and U6861 (N_6861,N_5061,N_5547);
nor U6862 (N_6862,N_5422,N_5043);
and U6863 (N_6863,N_5705,N_5744);
nor U6864 (N_6864,N_5742,N_5413);
and U6865 (N_6865,N_5978,N_5293);
or U6866 (N_6866,N_5920,N_5363);
xnor U6867 (N_6867,N_5509,N_5859);
xor U6868 (N_6868,N_5046,N_5783);
nand U6869 (N_6869,N_5361,N_5352);
xnor U6870 (N_6870,N_5742,N_5439);
nand U6871 (N_6871,N_5975,N_5261);
and U6872 (N_6872,N_5912,N_5657);
or U6873 (N_6873,N_5645,N_5958);
or U6874 (N_6874,N_5352,N_5118);
and U6875 (N_6875,N_5517,N_5943);
and U6876 (N_6876,N_5981,N_5138);
nand U6877 (N_6877,N_5156,N_5330);
or U6878 (N_6878,N_5290,N_5845);
nand U6879 (N_6879,N_5033,N_5523);
and U6880 (N_6880,N_5683,N_5280);
xnor U6881 (N_6881,N_5268,N_5786);
nor U6882 (N_6882,N_5879,N_5318);
nand U6883 (N_6883,N_5941,N_5400);
xor U6884 (N_6884,N_5441,N_5142);
xor U6885 (N_6885,N_5315,N_5650);
nand U6886 (N_6886,N_5500,N_5419);
or U6887 (N_6887,N_5485,N_5920);
and U6888 (N_6888,N_5493,N_5526);
xor U6889 (N_6889,N_5069,N_5538);
or U6890 (N_6890,N_5189,N_5304);
or U6891 (N_6891,N_5201,N_5182);
or U6892 (N_6892,N_5657,N_5065);
xor U6893 (N_6893,N_5494,N_5560);
nor U6894 (N_6894,N_5359,N_5848);
nor U6895 (N_6895,N_5742,N_5246);
and U6896 (N_6896,N_5819,N_5316);
xnor U6897 (N_6897,N_5114,N_5832);
nand U6898 (N_6898,N_5808,N_5297);
and U6899 (N_6899,N_5569,N_5130);
nor U6900 (N_6900,N_5002,N_5813);
xnor U6901 (N_6901,N_5673,N_5923);
or U6902 (N_6902,N_5721,N_5612);
nand U6903 (N_6903,N_5544,N_5678);
nor U6904 (N_6904,N_5921,N_5994);
or U6905 (N_6905,N_5405,N_5368);
and U6906 (N_6906,N_5786,N_5152);
and U6907 (N_6907,N_5570,N_5897);
nand U6908 (N_6908,N_5379,N_5179);
nor U6909 (N_6909,N_5225,N_5761);
and U6910 (N_6910,N_5924,N_5032);
nand U6911 (N_6911,N_5226,N_5958);
nand U6912 (N_6912,N_5358,N_5913);
xnor U6913 (N_6913,N_5480,N_5762);
and U6914 (N_6914,N_5797,N_5205);
nand U6915 (N_6915,N_5113,N_5077);
xnor U6916 (N_6916,N_5671,N_5191);
xnor U6917 (N_6917,N_5312,N_5430);
and U6918 (N_6918,N_5842,N_5500);
nand U6919 (N_6919,N_5047,N_5481);
nor U6920 (N_6920,N_5077,N_5913);
nor U6921 (N_6921,N_5279,N_5614);
and U6922 (N_6922,N_5278,N_5170);
nand U6923 (N_6923,N_5258,N_5300);
or U6924 (N_6924,N_5623,N_5509);
or U6925 (N_6925,N_5193,N_5260);
nand U6926 (N_6926,N_5733,N_5028);
or U6927 (N_6927,N_5819,N_5337);
or U6928 (N_6928,N_5888,N_5184);
nand U6929 (N_6929,N_5299,N_5736);
and U6930 (N_6930,N_5489,N_5117);
xor U6931 (N_6931,N_5629,N_5003);
nor U6932 (N_6932,N_5022,N_5373);
nor U6933 (N_6933,N_5123,N_5043);
or U6934 (N_6934,N_5969,N_5853);
and U6935 (N_6935,N_5687,N_5082);
nor U6936 (N_6936,N_5611,N_5678);
or U6937 (N_6937,N_5075,N_5847);
or U6938 (N_6938,N_5946,N_5454);
nor U6939 (N_6939,N_5240,N_5600);
or U6940 (N_6940,N_5051,N_5838);
nand U6941 (N_6941,N_5710,N_5314);
and U6942 (N_6942,N_5197,N_5729);
or U6943 (N_6943,N_5808,N_5831);
or U6944 (N_6944,N_5429,N_5533);
nand U6945 (N_6945,N_5594,N_5229);
xor U6946 (N_6946,N_5448,N_5831);
xnor U6947 (N_6947,N_5226,N_5026);
nor U6948 (N_6948,N_5306,N_5308);
nor U6949 (N_6949,N_5598,N_5879);
or U6950 (N_6950,N_5099,N_5892);
xor U6951 (N_6951,N_5048,N_5584);
or U6952 (N_6952,N_5708,N_5225);
and U6953 (N_6953,N_5469,N_5413);
or U6954 (N_6954,N_5246,N_5454);
or U6955 (N_6955,N_5493,N_5509);
nand U6956 (N_6956,N_5708,N_5456);
xor U6957 (N_6957,N_5353,N_5475);
and U6958 (N_6958,N_5030,N_5008);
or U6959 (N_6959,N_5540,N_5303);
nor U6960 (N_6960,N_5697,N_5452);
nor U6961 (N_6961,N_5829,N_5619);
and U6962 (N_6962,N_5276,N_5211);
nand U6963 (N_6963,N_5967,N_5523);
or U6964 (N_6964,N_5962,N_5715);
and U6965 (N_6965,N_5691,N_5970);
nor U6966 (N_6966,N_5431,N_5654);
nand U6967 (N_6967,N_5650,N_5311);
nor U6968 (N_6968,N_5922,N_5993);
and U6969 (N_6969,N_5882,N_5724);
nor U6970 (N_6970,N_5993,N_5056);
xor U6971 (N_6971,N_5693,N_5543);
nand U6972 (N_6972,N_5754,N_5333);
and U6973 (N_6973,N_5480,N_5991);
nand U6974 (N_6974,N_5689,N_5991);
and U6975 (N_6975,N_5331,N_5409);
nand U6976 (N_6976,N_5622,N_5327);
xor U6977 (N_6977,N_5057,N_5287);
nor U6978 (N_6978,N_5125,N_5613);
xnor U6979 (N_6979,N_5059,N_5525);
nand U6980 (N_6980,N_5929,N_5508);
or U6981 (N_6981,N_5737,N_5240);
xnor U6982 (N_6982,N_5839,N_5760);
nand U6983 (N_6983,N_5829,N_5324);
nor U6984 (N_6984,N_5598,N_5982);
and U6985 (N_6985,N_5824,N_5733);
or U6986 (N_6986,N_5553,N_5031);
nand U6987 (N_6987,N_5583,N_5835);
nand U6988 (N_6988,N_5143,N_5572);
and U6989 (N_6989,N_5089,N_5612);
nor U6990 (N_6990,N_5897,N_5103);
xnor U6991 (N_6991,N_5762,N_5424);
nand U6992 (N_6992,N_5807,N_5783);
and U6993 (N_6993,N_5922,N_5431);
and U6994 (N_6994,N_5407,N_5401);
xor U6995 (N_6995,N_5829,N_5789);
xnor U6996 (N_6996,N_5580,N_5460);
nor U6997 (N_6997,N_5451,N_5309);
and U6998 (N_6998,N_5104,N_5395);
xor U6999 (N_6999,N_5612,N_5719);
xnor U7000 (N_7000,N_6629,N_6383);
nor U7001 (N_7001,N_6186,N_6347);
nor U7002 (N_7002,N_6304,N_6093);
or U7003 (N_7003,N_6833,N_6731);
and U7004 (N_7004,N_6732,N_6518);
or U7005 (N_7005,N_6138,N_6752);
nand U7006 (N_7006,N_6169,N_6307);
and U7007 (N_7007,N_6675,N_6358);
or U7008 (N_7008,N_6269,N_6637);
xnor U7009 (N_7009,N_6840,N_6936);
nor U7010 (N_7010,N_6800,N_6508);
or U7011 (N_7011,N_6626,N_6669);
xnor U7012 (N_7012,N_6402,N_6743);
nor U7013 (N_7013,N_6682,N_6444);
or U7014 (N_7014,N_6040,N_6393);
and U7015 (N_7015,N_6948,N_6797);
and U7016 (N_7016,N_6999,N_6815);
or U7017 (N_7017,N_6645,N_6449);
nand U7018 (N_7018,N_6670,N_6477);
or U7019 (N_7019,N_6987,N_6030);
or U7020 (N_7020,N_6514,N_6021);
nor U7021 (N_7021,N_6971,N_6058);
nand U7022 (N_7022,N_6389,N_6211);
xnor U7023 (N_7023,N_6500,N_6312);
nor U7024 (N_7024,N_6893,N_6192);
xnor U7025 (N_7025,N_6061,N_6709);
nand U7026 (N_7026,N_6713,N_6598);
nor U7027 (N_7027,N_6902,N_6397);
nor U7028 (N_7028,N_6217,N_6396);
nand U7029 (N_7029,N_6339,N_6114);
or U7030 (N_7030,N_6676,N_6403);
or U7031 (N_7031,N_6289,N_6585);
nor U7032 (N_7032,N_6411,N_6355);
nor U7033 (N_7033,N_6969,N_6464);
nor U7034 (N_7034,N_6538,N_6554);
or U7035 (N_7035,N_6995,N_6698);
nor U7036 (N_7036,N_6658,N_6290);
nor U7037 (N_7037,N_6672,N_6496);
or U7038 (N_7038,N_6556,N_6539);
nor U7039 (N_7039,N_6441,N_6866);
and U7040 (N_7040,N_6245,N_6070);
or U7041 (N_7041,N_6791,N_6011);
and U7042 (N_7042,N_6793,N_6210);
xor U7043 (N_7043,N_6320,N_6688);
xor U7044 (N_7044,N_6684,N_6907);
xor U7045 (N_7045,N_6116,N_6112);
or U7046 (N_7046,N_6381,N_6949);
xnor U7047 (N_7047,N_6272,N_6858);
nand U7048 (N_7048,N_6031,N_6369);
xor U7049 (N_7049,N_6136,N_6697);
xor U7050 (N_7050,N_6785,N_6377);
nor U7051 (N_7051,N_6313,N_6437);
nand U7052 (N_7052,N_6310,N_6043);
or U7053 (N_7053,N_6264,N_6525);
or U7054 (N_7054,N_6679,N_6699);
nor U7055 (N_7055,N_6729,N_6214);
nor U7056 (N_7056,N_6165,N_6035);
or U7057 (N_7057,N_6753,N_6484);
nand U7058 (N_7058,N_6755,N_6818);
nand U7059 (N_7059,N_6431,N_6053);
nand U7060 (N_7060,N_6008,N_6228);
and U7061 (N_7061,N_6980,N_6929);
nor U7062 (N_7062,N_6895,N_6931);
xor U7063 (N_7063,N_6327,N_6328);
xnor U7064 (N_7064,N_6838,N_6849);
nor U7065 (N_7065,N_6368,N_6975);
nor U7066 (N_7066,N_6692,N_6303);
xor U7067 (N_7067,N_6851,N_6302);
nor U7068 (N_7068,N_6483,N_6480);
or U7069 (N_7069,N_6925,N_6723);
xnor U7070 (N_7070,N_6612,N_6015);
nor U7071 (N_7071,N_6408,N_6592);
or U7072 (N_7072,N_6482,N_6230);
xor U7073 (N_7073,N_6886,N_6125);
xnor U7074 (N_7074,N_6946,N_6638);
nor U7075 (N_7075,N_6549,N_6375);
xnor U7076 (N_7076,N_6152,N_6174);
or U7077 (N_7077,N_6968,N_6776);
nand U7078 (N_7078,N_6773,N_6364);
or U7079 (N_7079,N_6146,N_6453);
xnor U7080 (N_7080,N_6519,N_6560);
nand U7081 (N_7081,N_6502,N_6433);
xnor U7082 (N_7082,N_6241,N_6470);
and U7083 (N_7083,N_6887,N_6494);
nor U7084 (N_7084,N_6610,N_6844);
xor U7085 (N_7085,N_6227,N_6641);
nand U7086 (N_7086,N_6242,N_6129);
nor U7087 (N_7087,N_6478,N_6395);
and U7088 (N_7088,N_6473,N_6287);
nand U7089 (N_7089,N_6181,N_6348);
and U7090 (N_7090,N_6728,N_6790);
and U7091 (N_7091,N_6940,N_6599);
and U7092 (N_7092,N_6526,N_6110);
or U7093 (N_7093,N_6529,N_6106);
nand U7094 (N_7094,N_6663,N_6628);
and U7095 (N_7095,N_6515,N_6250);
or U7096 (N_7096,N_6077,N_6258);
or U7097 (N_7097,N_6363,N_6545);
and U7098 (N_7098,N_6229,N_6039);
or U7099 (N_7099,N_6774,N_6954);
xor U7100 (N_7100,N_6220,N_6288);
nor U7101 (N_7101,N_6633,N_6821);
or U7102 (N_7102,N_6885,N_6680);
or U7103 (N_7103,N_6080,N_6909);
or U7104 (N_7104,N_6894,N_6427);
nor U7105 (N_7105,N_6719,N_6194);
or U7106 (N_7106,N_6247,N_6845);
or U7107 (N_7107,N_6689,N_6499);
or U7108 (N_7108,N_6023,N_6710);
xnor U7109 (N_7109,N_6701,N_6737);
nand U7110 (N_7110,N_6153,N_6051);
and U7111 (N_7111,N_6993,N_6990);
xor U7112 (N_7112,N_6280,N_6118);
or U7113 (N_7113,N_6809,N_6472);
nand U7114 (N_7114,N_6337,N_6371);
nand U7115 (N_7115,N_6385,N_6516);
xor U7116 (N_7116,N_6742,N_6655);
xnor U7117 (N_7117,N_6253,N_6621);
and U7118 (N_7118,N_6798,N_6275);
xnor U7119 (N_7119,N_6782,N_6009);
and U7120 (N_7120,N_6342,N_6081);
nand U7121 (N_7121,N_6501,N_6796);
and U7122 (N_7122,N_6521,N_6561);
xor U7123 (N_7123,N_6088,N_6157);
nor U7124 (N_7124,N_6581,N_6270);
and U7125 (N_7125,N_6222,N_6741);
nand U7126 (N_7126,N_6255,N_6498);
nand U7127 (N_7127,N_6947,N_6038);
nand U7128 (N_7128,N_6533,N_6158);
xor U7129 (N_7129,N_6848,N_6366);
xnor U7130 (N_7130,N_6846,N_6825);
nand U7131 (N_7131,N_6294,N_6187);
or U7132 (N_7132,N_6768,N_6244);
or U7133 (N_7133,N_6465,N_6479);
nand U7134 (N_7134,N_6237,N_6919);
nand U7135 (N_7135,N_6674,N_6295);
nor U7136 (N_7136,N_6787,N_6373);
and U7137 (N_7137,N_6992,N_6817);
xnor U7138 (N_7138,N_6195,N_6197);
xnor U7139 (N_7139,N_6601,N_6073);
xor U7140 (N_7140,N_6092,N_6913);
and U7141 (N_7141,N_6795,N_6273);
nand U7142 (N_7142,N_6151,N_6918);
nor U7143 (N_7143,N_6096,N_6075);
or U7144 (N_7144,N_6634,N_6757);
xor U7145 (N_7145,N_6718,N_6983);
nand U7146 (N_7146,N_6961,N_6362);
nor U7147 (N_7147,N_6962,N_6937);
nand U7148 (N_7148,N_6277,N_6693);
and U7149 (N_7149,N_6350,N_6235);
nor U7150 (N_7150,N_6248,N_6884);
and U7151 (N_7151,N_6301,N_6132);
nor U7152 (N_7152,N_6082,N_6531);
nand U7153 (N_7153,N_6175,N_6715);
and U7154 (N_7154,N_6686,N_6703);
or U7155 (N_7155,N_6520,N_6551);
xor U7156 (N_7156,N_6984,N_6924);
xor U7157 (N_7157,N_6681,N_6857);
and U7158 (N_7158,N_6690,N_6696);
nor U7159 (N_7159,N_6986,N_6841);
or U7160 (N_7160,N_6430,N_6619);
xor U7161 (N_7161,N_6102,N_6950);
and U7162 (N_7162,N_6279,N_6996);
and U7163 (N_7163,N_6346,N_6330);
or U7164 (N_7164,N_6808,N_6193);
xor U7165 (N_7165,N_6588,N_6562);
or U7166 (N_7166,N_6998,N_6813);
xnor U7167 (N_7167,N_6650,N_6758);
nand U7168 (N_7168,N_6204,N_6452);
or U7169 (N_7169,N_6763,N_6378);
or U7170 (N_7170,N_6702,N_6580);
xor U7171 (N_7171,N_6746,N_6865);
nand U7172 (N_7172,N_6890,N_6631);
and U7173 (N_7173,N_6246,N_6010);
xnor U7174 (N_7174,N_6318,N_6127);
nand U7175 (N_7175,N_6391,N_6847);
nand U7176 (N_7176,N_6336,N_6888);
nor U7177 (N_7177,N_6126,N_6636);
xnor U7178 (N_7178,N_6827,N_6232);
nand U7179 (N_7179,N_6955,N_6137);
or U7180 (N_7180,N_6234,N_6830);
xor U7181 (N_7181,N_6673,N_6831);
and U7182 (N_7182,N_6467,N_6879);
xor U7183 (N_7183,N_6299,N_6256);
nand U7184 (N_7184,N_6422,N_6311);
nor U7185 (N_7185,N_6804,N_6022);
nand U7186 (N_7186,N_6874,N_6769);
and U7187 (N_7187,N_6807,N_6324);
nand U7188 (N_7188,N_6268,N_6683);
or U7189 (N_7189,N_6871,N_6407);
or U7190 (N_7190,N_6823,N_6756);
and U7191 (N_7191,N_6872,N_6648);
nor U7192 (N_7192,N_6485,N_6142);
and U7193 (N_7193,N_6777,N_6527);
xnor U7194 (N_7194,N_6343,N_6801);
or U7195 (N_7195,N_6476,N_6083);
xor U7196 (N_7196,N_6661,N_6458);
or U7197 (N_7197,N_6260,N_6664);
xor U7198 (N_7198,N_6259,N_6837);
xnor U7199 (N_7199,N_6180,N_6249);
or U7200 (N_7200,N_6367,N_6542);
and U7201 (N_7201,N_6360,N_6811);
nor U7202 (N_7202,N_6240,N_6783);
nand U7203 (N_7203,N_6802,N_6920);
xor U7204 (N_7204,N_6916,N_6201);
nand U7205 (N_7205,N_6666,N_6861);
xnor U7206 (N_7206,N_6344,N_6466);
or U7207 (N_7207,N_6943,N_6706);
or U7208 (N_7208,N_6432,N_6238);
xnor U7209 (N_7209,N_6912,N_6932);
xor U7210 (N_7210,N_6577,N_6425);
and U7211 (N_7211,N_6141,N_6606);
nand U7212 (N_7212,N_6944,N_6573);
xnor U7213 (N_7213,N_6727,N_6434);
or U7214 (N_7214,N_6001,N_6412);
xor U7215 (N_7215,N_6376,N_6308);
nand U7216 (N_7216,N_6509,N_6394);
nand U7217 (N_7217,N_6066,N_6921);
xnor U7218 (N_7218,N_6503,N_6063);
xor U7219 (N_7219,N_6429,N_6511);
nor U7220 (N_7220,N_6446,N_6747);
nor U7221 (N_7221,N_6196,N_6770);
xnor U7222 (N_7222,N_6794,N_6155);
xnor U7223 (N_7223,N_6159,N_6543);
nor U7224 (N_7224,N_6724,N_6122);
and U7225 (N_7225,N_6869,N_6016);
nor U7226 (N_7226,N_6878,N_6736);
or U7227 (N_7227,N_6421,N_6700);
or U7228 (N_7228,N_6002,N_6605);
and U7229 (N_7229,N_6558,N_6677);
xor U7230 (N_7230,N_6267,N_6130);
nor U7231 (N_7231,N_6590,N_6145);
nand U7232 (N_7232,N_6111,N_6120);
nor U7233 (N_7233,N_6048,N_6251);
xor U7234 (N_7234,N_6037,N_6548);
and U7235 (N_7235,N_6922,N_6915);
and U7236 (N_7236,N_6910,N_6406);
xnor U7237 (N_7237,N_6812,N_6958);
and U7238 (N_7238,N_6544,N_6319);
xnor U7239 (N_7239,N_6474,N_6341);
or U7240 (N_7240,N_6291,N_6517);
nor U7241 (N_7241,N_6261,N_6564);
nand U7242 (N_7242,N_6492,N_6563);
and U7243 (N_7243,N_6711,N_6338);
and U7244 (N_7244,N_6135,N_6060);
and U7245 (N_7245,N_6099,N_6891);
or U7246 (N_7246,N_6027,N_6789);
nand U7247 (N_7247,N_6414,N_6659);
or U7248 (N_7248,N_6717,N_6162);
and U7249 (N_7249,N_6788,N_6978);
nor U7250 (N_7250,N_6832,N_6639);
nand U7251 (N_7251,N_6864,N_6468);
and U7252 (N_7252,N_6625,N_6143);
or U7253 (N_7253,N_6816,N_6855);
and U7254 (N_7254,N_6578,N_6216);
nor U7255 (N_7255,N_6665,N_6438);
and U7256 (N_7256,N_6036,N_6007);
and U7257 (N_7257,N_6772,N_6644);
or U7258 (N_7258,N_6156,N_6184);
nor U7259 (N_7259,N_6939,N_6620);
nand U7260 (N_7260,N_6972,N_6805);
xnor U7261 (N_7261,N_6989,N_6067);
or U7262 (N_7262,N_6456,N_6356);
xnor U7263 (N_7263,N_6224,N_6231);
or U7264 (N_7264,N_6415,N_6780);
xnor U7265 (N_7265,N_6906,N_6370);
and U7266 (N_7266,N_6013,N_6266);
or U7267 (N_7267,N_6775,N_6604);
xor U7268 (N_7268,N_6447,N_6651);
or U7269 (N_7269,N_6078,N_6759);
and U7270 (N_7270,N_6875,N_6019);
nor U7271 (N_7271,N_6765,N_6460);
nand U7272 (N_7272,N_6098,N_6387);
or U7273 (N_7273,N_6766,N_6822);
nor U7274 (N_7274,N_6160,N_6781);
or U7275 (N_7275,N_6147,N_6896);
nor U7276 (N_7276,N_6003,N_6591);
nor U7277 (N_7277,N_6045,N_6380);
nand U7278 (N_7278,N_6000,N_6488);
nand U7279 (N_7279,N_6309,N_6101);
nand U7280 (N_7280,N_6941,N_6392);
xor U7281 (N_7281,N_6055,N_6685);
nor U7282 (N_7282,N_6300,N_6457);
nand U7283 (N_7283,N_6762,N_6882);
xor U7284 (N_7284,N_6439,N_6170);
nor U7285 (N_7285,N_6094,N_6559);
nor U7286 (N_7286,N_6401,N_6462);
nor U7287 (N_7287,N_6965,N_6173);
nor U7288 (N_7288,N_6982,N_6190);
nor U7289 (N_7289,N_6979,N_6574);
nand U7290 (N_7290,N_6469,N_6257);
nor U7291 (N_7291,N_6325,N_6017);
or U7292 (N_7292,N_6738,N_6792);
nor U7293 (N_7293,N_6883,N_6569);
or U7294 (N_7294,N_6981,N_6897);
and U7295 (N_7295,N_6938,N_6451);
nand U7296 (N_7296,N_6933,N_6413);
and U7297 (N_7297,N_6835,N_6900);
and U7298 (N_7298,N_6068,N_6386);
or U7299 (N_7299,N_6935,N_6404);
nand U7300 (N_7300,N_6293,N_6930);
nor U7301 (N_7301,N_6660,N_6536);
xor U7302 (N_7302,N_6163,N_6357);
nor U7303 (N_7303,N_6750,N_6760);
and U7304 (N_7304,N_6047,N_6778);
nand U7305 (N_7305,N_6442,N_6209);
nor U7306 (N_7306,N_6354,N_6254);
nor U7307 (N_7307,N_6589,N_6179);
and U7308 (N_7308,N_6860,N_6623);
and U7309 (N_7309,N_6630,N_6326);
nand U7310 (N_7310,N_6416,N_6115);
xnor U7311 (N_7311,N_6553,N_6877);
nand U7312 (N_7312,N_6786,N_6349);
or U7313 (N_7313,N_6024,N_6547);
nor U7314 (N_7314,N_6957,N_6086);
nor U7315 (N_7315,N_6904,N_6445);
nand U7316 (N_7316,N_6419,N_6207);
nor U7317 (N_7317,N_6108,N_6218);
nor U7318 (N_7318,N_6820,N_6150);
nor U7319 (N_7319,N_6359,N_6905);
nor U7320 (N_7320,N_6934,N_6899);
xor U7321 (N_7321,N_6819,N_6603);
or U7322 (N_7322,N_6927,N_6345);
or U7323 (N_7323,N_6399,N_6046);
xor U7324 (N_7324,N_6198,N_6627);
xor U7325 (N_7325,N_6139,N_6532);
xnor U7326 (N_7326,N_6880,N_6033);
nand U7327 (N_7327,N_6314,N_6405);
or U7328 (N_7328,N_6384,N_6754);
or U7329 (N_7329,N_6191,N_6144);
nand U7330 (N_7330,N_6056,N_6988);
and U7331 (N_7331,N_6353,N_6213);
nor U7332 (N_7332,N_6720,N_6332);
nand U7333 (N_7333,N_6020,N_6656);
and U7334 (N_7334,N_6767,N_6565);
xor U7335 (N_7335,N_6059,N_6164);
nand U7336 (N_7336,N_6870,N_6761);
nor U7337 (N_7337,N_6600,N_6493);
or U7338 (N_7338,N_6635,N_6225);
xor U7339 (N_7339,N_6567,N_6265);
nor U7340 (N_7340,N_6740,N_6582);
nor U7341 (N_7341,N_6495,N_6667);
nor U7342 (N_7342,N_6528,N_6282);
nand U7343 (N_7343,N_6647,N_6298);
nor U7344 (N_7344,N_6124,N_6172);
xnor U7345 (N_7345,N_6974,N_6243);
or U7346 (N_7346,N_6952,N_6486);
nor U7347 (N_7347,N_6642,N_6443);
nand U7348 (N_7348,N_6052,N_6616);
nand U7349 (N_7349,N_6856,N_6951);
or U7350 (N_7350,N_6089,N_6607);
xor U7351 (N_7351,N_6956,N_6892);
xnor U7352 (N_7352,N_6908,N_6140);
xor U7353 (N_7353,N_6006,N_6853);
xor U7354 (N_7354,N_6065,N_6203);
and U7355 (N_7355,N_6123,N_6091);
xor U7356 (N_7356,N_6678,N_6049);
xnor U7357 (N_7357,N_6315,N_6149);
and U7358 (N_7358,N_6862,N_6409);
nand U7359 (N_7359,N_6928,N_6461);
nand U7360 (N_7360,N_6970,N_6707);
or U7361 (N_7361,N_6911,N_6185);
xor U7362 (N_7362,N_6522,N_6044);
xor U7363 (N_7363,N_6881,N_6997);
nor U7364 (N_7364,N_6323,N_6398);
nand U7365 (N_7365,N_6859,N_6352);
xor U7366 (N_7366,N_6923,N_6744);
and U7367 (N_7367,N_6236,N_6057);
nand U7368 (N_7368,N_6283,N_6379);
nand U7369 (N_7369,N_6541,N_6239);
nand U7370 (N_7370,N_6296,N_6100);
and U7371 (N_7371,N_6285,N_6829);
nand U7372 (N_7372,N_6463,N_6608);
and U7373 (N_7373,N_6566,N_6221);
xor U7374 (N_7374,N_6212,N_6104);
and U7375 (N_7375,N_6182,N_6097);
and U7376 (N_7376,N_6652,N_6994);
nor U7377 (N_7377,N_6842,N_6889);
or U7378 (N_7378,N_6552,N_6739);
or U7379 (N_7379,N_6131,N_6568);
nand U7380 (N_7380,N_6103,N_6121);
or U7381 (N_7381,N_6716,N_6424);
nand U7382 (N_7382,N_6459,N_6824);
or U7383 (N_7383,N_6340,N_6205);
nor U7384 (N_7384,N_6177,N_6602);
nor U7385 (N_7385,N_6617,N_6109);
nand U7386 (N_7386,N_6436,N_6032);
nand U7387 (N_7387,N_6417,N_6614);
xor U7388 (N_7388,N_6335,N_6199);
and U7389 (N_7389,N_6784,N_6168);
xnor U7390 (N_7390,N_6977,N_6810);
and U7391 (N_7391,N_6632,N_6618);
nor U7392 (N_7392,N_6189,N_6867);
xor U7393 (N_7393,N_6597,N_6593);
nor U7394 (N_7394,N_6085,N_6722);
xor U7395 (N_7395,N_6535,N_6166);
nand U7396 (N_7396,N_6262,N_6450);
xor U7397 (N_7397,N_6004,N_6555);
and U7398 (N_7398,N_6991,N_6534);
or U7399 (N_7399,N_6726,N_6714);
and U7400 (N_7400,N_6826,N_6671);
xnor U7401 (N_7401,N_6653,N_6624);
or U7402 (N_7402,N_6985,N_6167);
or U7403 (N_7403,N_6803,N_6426);
or U7404 (N_7404,N_6105,N_6557);
or U7405 (N_7405,N_6622,N_6018);
nor U7406 (N_7406,N_6512,N_6615);
xnor U7407 (N_7407,N_6868,N_6183);
nand U7408 (N_7408,N_6361,N_6852);
or U7409 (N_7409,N_6284,N_6148);
or U7410 (N_7410,N_6400,N_6745);
xor U7411 (N_7411,N_6072,N_6223);
nor U7412 (N_7412,N_6490,N_6028);
or U7413 (N_7413,N_6305,N_6054);
and U7414 (N_7414,N_6834,N_6964);
and U7415 (N_7415,N_6725,N_6321);
nand U7416 (N_7416,N_6188,N_6281);
nor U7417 (N_7417,N_6537,N_6587);
nor U7418 (N_7418,N_6041,N_6322);
nor U7419 (N_7419,N_6926,N_6730);
or U7420 (N_7420,N_6643,N_6034);
and U7421 (N_7421,N_6491,N_6901);
and U7422 (N_7422,N_6850,N_6372);
nor U7423 (N_7423,N_6876,N_6540);
nor U7424 (N_7424,N_6297,N_6695);
or U7425 (N_7425,N_6062,N_6200);
nor U7426 (N_7426,N_6410,N_6524);
xor U7427 (N_7427,N_6523,N_6005);
nor U7428 (N_7428,N_6959,N_6117);
or U7429 (N_7429,N_6779,N_6076);
xor U7430 (N_7430,N_6506,N_6276);
nor U7431 (N_7431,N_6095,N_6487);
or U7432 (N_7432,N_6550,N_6571);
nor U7433 (N_7433,N_6583,N_6390);
xnor U7434 (N_7434,N_6012,N_6440);
xor U7435 (N_7435,N_6481,N_6575);
or U7436 (N_7436,N_6814,N_6687);
nand U7437 (N_7437,N_6161,N_6316);
xor U7438 (N_7438,N_6504,N_6691);
and U7439 (N_7439,N_6154,N_6507);
nand U7440 (N_7440,N_6662,N_6286);
nor U7441 (N_7441,N_6735,N_6572);
nor U7442 (N_7442,N_6274,N_6278);
or U7443 (N_7443,N_6646,N_6176);
nand U7444 (N_7444,N_6586,N_6748);
nor U7445 (N_7445,N_6079,N_6084);
nor U7446 (N_7446,N_6042,N_6202);
nand U7447 (N_7447,N_6903,N_6087);
xnor U7448 (N_7448,N_6455,N_6334);
xnor U7449 (N_7449,N_6382,N_6584);
or U7450 (N_7450,N_6963,N_6090);
nand U7451 (N_7451,N_6329,N_6252);
xnor U7452 (N_7452,N_6292,N_6331);
nor U7453 (N_7453,N_6657,N_6505);
and U7454 (N_7454,N_6854,N_6351);
xor U7455 (N_7455,N_6418,N_6107);
and U7456 (N_7456,N_6074,N_6570);
nor U7457 (N_7457,N_6489,N_6839);
and U7458 (N_7458,N_6423,N_6071);
and U7459 (N_7459,N_6863,N_6613);
and U7460 (N_7460,N_6064,N_6233);
nand U7461 (N_7461,N_6128,N_6471);
and U7462 (N_7462,N_6654,N_6206);
xnor U7463 (N_7463,N_6306,N_6806);
and U7464 (N_7464,N_6510,N_6219);
or U7465 (N_7465,N_6178,N_6317);
nor U7466 (N_7466,N_6226,N_6475);
and U7467 (N_7467,N_6611,N_6134);
xnor U7468 (N_7468,N_6365,N_6594);
xor U7469 (N_7469,N_6873,N_6113);
or U7470 (N_7470,N_6171,N_6428);
or U7471 (N_7471,N_6420,N_6942);
or U7472 (N_7472,N_6208,N_6914);
nor U7473 (N_7473,N_6945,N_6215);
nor U7474 (N_7474,N_6976,N_6454);
and U7475 (N_7475,N_6771,N_6953);
and U7476 (N_7476,N_6967,N_6448);
nand U7477 (N_7477,N_6050,N_6751);
and U7478 (N_7478,N_6026,N_6374);
and U7479 (N_7479,N_6576,N_6014);
or U7480 (N_7480,N_6513,N_6333);
nand U7481 (N_7481,N_6960,N_6119);
xor U7482 (N_7482,N_6069,N_6609);
xor U7483 (N_7483,N_6497,N_6029);
xor U7484 (N_7484,N_6708,N_6596);
or U7485 (N_7485,N_6694,N_6843);
or U7486 (N_7486,N_6733,N_6649);
nor U7487 (N_7487,N_6749,N_6828);
xor U7488 (N_7488,N_6721,N_6668);
or U7489 (N_7489,N_6388,N_6973);
nor U7490 (N_7490,N_6799,N_6917);
nor U7491 (N_7491,N_6546,N_6836);
nand U7492 (N_7492,N_6263,N_6579);
and U7493 (N_7493,N_6734,N_6530);
or U7494 (N_7494,N_6435,N_6595);
nor U7495 (N_7495,N_6640,N_6704);
nor U7496 (N_7496,N_6898,N_6712);
and U7497 (N_7497,N_6025,N_6705);
xnor U7498 (N_7498,N_6764,N_6966);
nand U7499 (N_7499,N_6133,N_6271);
nor U7500 (N_7500,N_6480,N_6158);
and U7501 (N_7501,N_6282,N_6038);
xor U7502 (N_7502,N_6666,N_6819);
xor U7503 (N_7503,N_6903,N_6228);
or U7504 (N_7504,N_6001,N_6110);
xnor U7505 (N_7505,N_6335,N_6655);
or U7506 (N_7506,N_6692,N_6895);
xor U7507 (N_7507,N_6763,N_6153);
and U7508 (N_7508,N_6541,N_6245);
nand U7509 (N_7509,N_6414,N_6372);
nor U7510 (N_7510,N_6985,N_6537);
xnor U7511 (N_7511,N_6400,N_6789);
or U7512 (N_7512,N_6626,N_6865);
or U7513 (N_7513,N_6074,N_6695);
xor U7514 (N_7514,N_6220,N_6786);
nor U7515 (N_7515,N_6230,N_6727);
xor U7516 (N_7516,N_6096,N_6168);
or U7517 (N_7517,N_6595,N_6485);
or U7518 (N_7518,N_6931,N_6571);
or U7519 (N_7519,N_6890,N_6283);
and U7520 (N_7520,N_6088,N_6549);
and U7521 (N_7521,N_6816,N_6785);
or U7522 (N_7522,N_6952,N_6181);
xnor U7523 (N_7523,N_6701,N_6240);
nor U7524 (N_7524,N_6310,N_6215);
xnor U7525 (N_7525,N_6428,N_6509);
nand U7526 (N_7526,N_6289,N_6020);
and U7527 (N_7527,N_6391,N_6458);
and U7528 (N_7528,N_6059,N_6742);
and U7529 (N_7529,N_6691,N_6683);
and U7530 (N_7530,N_6841,N_6912);
or U7531 (N_7531,N_6500,N_6624);
and U7532 (N_7532,N_6723,N_6426);
xor U7533 (N_7533,N_6873,N_6049);
nand U7534 (N_7534,N_6136,N_6493);
nand U7535 (N_7535,N_6015,N_6122);
and U7536 (N_7536,N_6807,N_6801);
xor U7537 (N_7537,N_6727,N_6560);
nand U7538 (N_7538,N_6764,N_6223);
nor U7539 (N_7539,N_6222,N_6281);
and U7540 (N_7540,N_6546,N_6615);
nor U7541 (N_7541,N_6613,N_6031);
nand U7542 (N_7542,N_6103,N_6104);
nand U7543 (N_7543,N_6101,N_6883);
nor U7544 (N_7544,N_6142,N_6800);
nor U7545 (N_7545,N_6195,N_6669);
and U7546 (N_7546,N_6328,N_6470);
and U7547 (N_7547,N_6862,N_6960);
nand U7548 (N_7548,N_6217,N_6445);
or U7549 (N_7549,N_6209,N_6783);
nand U7550 (N_7550,N_6255,N_6744);
xnor U7551 (N_7551,N_6442,N_6221);
xor U7552 (N_7552,N_6591,N_6657);
nand U7553 (N_7553,N_6089,N_6563);
or U7554 (N_7554,N_6812,N_6624);
and U7555 (N_7555,N_6808,N_6365);
and U7556 (N_7556,N_6124,N_6317);
and U7557 (N_7557,N_6587,N_6006);
xnor U7558 (N_7558,N_6233,N_6712);
nor U7559 (N_7559,N_6641,N_6456);
and U7560 (N_7560,N_6003,N_6930);
and U7561 (N_7561,N_6620,N_6875);
nand U7562 (N_7562,N_6576,N_6176);
xnor U7563 (N_7563,N_6973,N_6680);
nor U7564 (N_7564,N_6871,N_6254);
and U7565 (N_7565,N_6960,N_6953);
nor U7566 (N_7566,N_6143,N_6784);
or U7567 (N_7567,N_6634,N_6845);
and U7568 (N_7568,N_6572,N_6047);
nand U7569 (N_7569,N_6235,N_6332);
and U7570 (N_7570,N_6656,N_6152);
xor U7571 (N_7571,N_6395,N_6651);
and U7572 (N_7572,N_6827,N_6458);
nand U7573 (N_7573,N_6410,N_6735);
nand U7574 (N_7574,N_6281,N_6359);
nand U7575 (N_7575,N_6770,N_6705);
xor U7576 (N_7576,N_6983,N_6434);
and U7577 (N_7577,N_6970,N_6141);
nor U7578 (N_7578,N_6333,N_6079);
nor U7579 (N_7579,N_6157,N_6142);
or U7580 (N_7580,N_6123,N_6303);
or U7581 (N_7581,N_6610,N_6644);
nor U7582 (N_7582,N_6532,N_6902);
nor U7583 (N_7583,N_6568,N_6390);
nand U7584 (N_7584,N_6531,N_6050);
nor U7585 (N_7585,N_6371,N_6261);
nor U7586 (N_7586,N_6214,N_6298);
or U7587 (N_7587,N_6707,N_6897);
xor U7588 (N_7588,N_6828,N_6177);
nand U7589 (N_7589,N_6933,N_6950);
or U7590 (N_7590,N_6741,N_6139);
or U7591 (N_7591,N_6191,N_6036);
nand U7592 (N_7592,N_6742,N_6931);
xor U7593 (N_7593,N_6392,N_6147);
nand U7594 (N_7594,N_6850,N_6959);
xnor U7595 (N_7595,N_6156,N_6419);
and U7596 (N_7596,N_6923,N_6732);
xnor U7597 (N_7597,N_6156,N_6908);
or U7598 (N_7598,N_6290,N_6003);
or U7599 (N_7599,N_6632,N_6904);
nor U7600 (N_7600,N_6190,N_6676);
nand U7601 (N_7601,N_6576,N_6119);
nand U7602 (N_7602,N_6191,N_6314);
nor U7603 (N_7603,N_6272,N_6824);
nor U7604 (N_7604,N_6277,N_6101);
nor U7605 (N_7605,N_6965,N_6870);
nor U7606 (N_7606,N_6203,N_6913);
nor U7607 (N_7607,N_6542,N_6257);
or U7608 (N_7608,N_6845,N_6098);
nor U7609 (N_7609,N_6156,N_6309);
or U7610 (N_7610,N_6301,N_6895);
and U7611 (N_7611,N_6977,N_6630);
nand U7612 (N_7612,N_6262,N_6279);
or U7613 (N_7613,N_6684,N_6810);
and U7614 (N_7614,N_6523,N_6365);
nand U7615 (N_7615,N_6314,N_6372);
or U7616 (N_7616,N_6961,N_6529);
and U7617 (N_7617,N_6860,N_6674);
or U7618 (N_7618,N_6498,N_6512);
nor U7619 (N_7619,N_6367,N_6973);
or U7620 (N_7620,N_6561,N_6372);
nand U7621 (N_7621,N_6113,N_6850);
nand U7622 (N_7622,N_6240,N_6036);
and U7623 (N_7623,N_6653,N_6189);
and U7624 (N_7624,N_6863,N_6654);
and U7625 (N_7625,N_6173,N_6072);
and U7626 (N_7626,N_6170,N_6588);
or U7627 (N_7627,N_6227,N_6940);
or U7628 (N_7628,N_6425,N_6805);
nand U7629 (N_7629,N_6903,N_6000);
nor U7630 (N_7630,N_6531,N_6934);
or U7631 (N_7631,N_6958,N_6023);
nor U7632 (N_7632,N_6514,N_6046);
xor U7633 (N_7633,N_6730,N_6018);
nand U7634 (N_7634,N_6749,N_6597);
nand U7635 (N_7635,N_6714,N_6253);
nand U7636 (N_7636,N_6957,N_6830);
nand U7637 (N_7637,N_6502,N_6418);
or U7638 (N_7638,N_6977,N_6864);
nand U7639 (N_7639,N_6412,N_6114);
or U7640 (N_7640,N_6388,N_6049);
and U7641 (N_7641,N_6693,N_6770);
and U7642 (N_7642,N_6234,N_6631);
nor U7643 (N_7643,N_6604,N_6324);
xnor U7644 (N_7644,N_6254,N_6910);
nor U7645 (N_7645,N_6901,N_6361);
nand U7646 (N_7646,N_6171,N_6417);
or U7647 (N_7647,N_6942,N_6560);
or U7648 (N_7648,N_6820,N_6240);
nor U7649 (N_7649,N_6312,N_6467);
nor U7650 (N_7650,N_6750,N_6448);
nand U7651 (N_7651,N_6617,N_6946);
or U7652 (N_7652,N_6489,N_6500);
nand U7653 (N_7653,N_6902,N_6210);
or U7654 (N_7654,N_6399,N_6343);
or U7655 (N_7655,N_6632,N_6068);
xor U7656 (N_7656,N_6496,N_6972);
nand U7657 (N_7657,N_6040,N_6600);
and U7658 (N_7658,N_6333,N_6824);
xnor U7659 (N_7659,N_6294,N_6304);
nand U7660 (N_7660,N_6281,N_6731);
and U7661 (N_7661,N_6790,N_6459);
xor U7662 (N_7662,N_6278,N_6912);
nor U7663 (N_7663,N_6012,N_6343);
nor U7664 (N_7664,N_6872,N_6950);
xnor U7665 (N_7665,N_6756,N_6544);
or U7666 (N_7666,N_6704,N_6657);
nand U7667 (N_7667,N_6613,N_6285);
and U7668 (N_7668,N_6896,N_6454);
xnor U7669 (N_7669,N_6874,N_6536);
or U7670 (N_7670,N_6558,N_6932);
or U7671 (N_7671,N_6794,N_6090);
nor U7672 (N_7672,N_6637,N_6296);
xnor U7673 (N_7673,N_6687,N_6906);
nand U7674 (N_7674,N_6366,N_6040);
nor U7675 (N_7675,N_6561,N_6573);
nand U7676 (N_7676,N_6491,N_6997);
xnor U7677 (N_7677,N_6134,N_6509);
xor U7678 (N_7678,N_6968,N_6303);
xor U7679 (N_7679,N_6016,N_6335);
xnor U7680 (N_7680,N_6878,N_6191);
xnor U7681 (N_7681,N_6893,N_6675);
or U7682 (N_7682,N_6777,N_6259);
nand U7683 (N_7683,N_6159,N_6260);
nor U7684 (N_7684,N_6665,N_6041);
and U7685 (N_7685,N_6030,N_6259);
xor U7686 (N_7686,N_6218,N_6458);
nand U7687 (N_7687,N_6744,N_6534);
nand U7688 (N_7688,N_6101,N_6513);
xnor U7689 (N_7689,N_6965,N_6631);
nor U7690 (N_7690,N_6401,N_6514);
and U7691 (N_7691,N_6313,N_6666);
nand U7692 (N_7692,N_6945,N_6150);
and U7693 (N_7693,N_6679,N_6555);
nand U7694 (N_7694,N_6775,N_6106);
nor U7695 (N_7695,N_6775,N_6633);
xor U7696 (N_7696,N_6713,N_6214);
xor U7697 (N_7697,N_6205,N_6912);
nor U7698 (N_7698,N_6874,N_6886);
and U7699 (N_7699,N_6010,N_6410);
nor U7700 (N_7700,N_6021,N_6468);
xor U7701 (N_7701,N_6690,N_6853);
and U7702 (N_7702,N_6551,N_6061);
nand U7703 (N_7703,N_6398,N_6017);
or U7704 (N_7704,N_6250,N_6956);
or U7705 (N_7705,N_6059,N_6049);
nand U7706 (N_7706,N_6123,N_6861);
nand U7707 (N_7707,N_6582,N_6324);
nor U7708 (N_7708,N_6664,N_6778);
nor U7709 (N_7709,N_6458,N_6960);
xor U7710 (N_7710,N_6938,N_6095);
and U7711 (N_7711,N_6715,N_6431);
or U7712 (N_7712,N_6851,N_6476);
xnor U7713 (N_7713,N_6870,N_6876);
nand U7714 (N_7714,N_6903,N_6821);
or U7715 (N_7715,N_6869,N_6307);
or U7716 (N_7716,N_6724,N_6517);
or U7717 (N_7717,N_6065,N_6431);
or U7718 (N_7718,N_6021,N_6133);
nor U7719 (N_7719,N_6065,N_6232);
xnor U7720 (N_7720,N_6941,N_6598);
or U7721 (N_7721,N_6253,N_6125);
nor U7722 (N_7722,N_6949,N_6362);
nand U7723 (N_7723,N_6098,N_6220);
xnor U7724 (N_7724,N_6697,N_6500);
or U7725 (N_7725,N_6232,N_6425);
or U7726 (N_7726,N_6782,N_6413);
nor U7727 (N_7727,N_6630,N_6562);
or U7728 (N_7728,N_6173,N_6471);
and U7729 (N_7729,N_6379,N_6241);
nor U7730 (N_7730,N_6940,N_6742);
and U7731 (N_7731,N_6751,N_6772);
and U7732 (N_7732,N_6526,N_6875);
nor U7733 (N_7733,N_6517,N_6961);
nand U7734 (N_7734,N_6435,N_6296);
nor U7735 (N_7735,N_6870,N_6981);
nor U7736 (N_7736,N_6578,N_6350);
nand U7737 (N_7737,N_6000,N_6825);
nand U7738 (N_7738,N_6611,N_6181);
xnor U7739 (N_7739,N_6296,N_6771);
nor U7740 (N_7740,N_6117,N_6382);
or U7741 (N_7741,N_6372,N_6036);
nand U7742 (N_7742,N_6958,N_6160);
and U7743 (N_7743,N_6536,N_6308);
or U7744 (N_7744,N_6013,N_6098);
nor U7745 (N_7745,N_6361,N_6190);
nand U7746 (N_7746,N_6064,N_6797);
and U7747 (N_7747,N_6625,N_6762);
or U7748 (N_7748,N_6524,N_6579);
nor U7749 (N_7749,N_6785,N_6703);
nor U7750 (N_7750,N_6026,N_6748);
nand U7751 (N_7751,N_6890,N_6786);
xor U7752 (N_7752,N_6460,N_6456);
xnor U7753 (N_7753,N_6637,N_6505);
nor U7754 (N_7754,N_6321,N_6690);
nand U7755 (N_7755,N_6958,N_6662);
nand U7756 (N_7756,N_6547,N_6053);
and U7757 (N_7757,N_6991,N_6504);
nor U7758 (N_7758,N_6533,N_6343);
nor U7759 (N_7759,N_6216,N_6028);
or U7760 (N_7760,N_6636,N_6922);
nor U7761 (N_7761,N_6213,N_6844);
xor U7762 (N_7762,N_6583,N_6318);
xnor U7763 (N_7763,N_6486,N_6235);
and U7764 (N_7764,N_6048,N_6104);
nor U7765 (N_7765,N_6887,N_6943);
nor U7766 (N_7766,N_6743,N_6945);
nand U7767 (N_7767,N_6109,N_6862);
xnor U7768 (N_7768,N_6956,N_6858);
or U7769 (N_7769,N_6843,N_6262);
or U7770 (N_7770,N_6467,N_6197);
nand U7771 (N_7771,N_6584,N_6250);
or U7772 (N_7772,N_6573,N_6245);
nand U7773 (N_7773,N_6230,N_6541);
nor U7774 (N_7774,N_6675,N_6749);
nand U7775 (N_7775,N_6170,N_6680);
or U7776 (N_7776,N_6390,N_6184);
nand U7777 (N_7777,N_6332,N_6303);
or U7778 (N_7778,N_6336,N_6898);
xor U7779 (N_7779,N_6581,N_6285);
xor U7780 (N_7780,N_6522,N_6612);
xor U7781 (N_7781,N_6137,N_6796);
nand U7782 (N_7782,N_6060,N_6653);
nand U7783 (N_7783,N_6839,N_6553);
and U7784 (N_7784,N_6762,N_6547);
nor U7785 (N_7785,N_6951,N_6716);
nor U7786 (N_7786,N_6869,N_6171);
nor U7787 (N_7787,N_6848,N_6469);
nand U7788 (N_7788,N_6135,N_6239);
or U7789 (N_7789,N_6356,N_6548);
nand U7790 (N_7790,N_6285,N_6248);
and U7791 (N_7791,N_6181,N_6405);
nor U7792 (N_7792,N_6419,N_6676);
and U7793 (N_7793,N_6269,N_6792);
and U7794 (N_7794,N_6010,N_6393);
or U7795 (N_7795,N_6252,N_6216);
or U7796 (N_7796,N_6285,N_6986);
xnor U7797 (N_7797,N_6600,N_6800);
or U7798 (N_7798,N_6109,N_6906);
xor U7799 (N_7799,N_6338,N_6385);
xor U7800 (N_7800,N_6574,N_6432);
nand U7801 (N_7801,N_6245,N_6207);
nor U7802 (N_7802,N_6597,N_6213);
nor U7803 (N_7803,N_6680,N_6696);
xnor U7804 (N_7804,N_6495,N_6106);
or U7805 (N_7805,N_6044,N_6192);
xor U7806 (N_7806,N_6434,N_6388);
nand U7807 (N_7807,N_6921,N_6383);
nor U7808 (N_7808,N_6072,N_6984);
nand U7809 (N_7809,N_6993,N_6789);
xnor U7810 (N_7810,N_6351,N_6976);
or U7811 (N_7811,N_6681,N_6472);
xor U7812 (N_7812,N_6968,N_6695);
xor U7813 (N_7813,N_6073,N_6919);
and U7814 (N_7814,N_6935,N_6850);
nor U7815 (N_7815,N_6511,N_6937);
xnor U7816 (N_7816,N_6748,N_6767);
nand U7817 (N_7817,N_6082,N_6928);
nand U7818 (N_7818,N_6227,N_6566);
nor U7819 (N_7819,N_6004,N_6094);
xnor U7820 (N_7820,N_6838,N_6711);
nor U7821 (N_7821,N_6638,N_6894);
nand U7822 (N_7822,N_6820,N_6152);
or U7823 (N_7823,N_6456,N_6337);
xor U7824 (N_7824,N_6217,N_6148);
or U7825 (N_7825,N_6461,N_6768);
or U7826 (N_7826,N_6508,N_6226);
nand U7827 (N_7827,N_6768,N_6258);
xnor U7828 (N_7828,N_6686,N_6506);
xor U7829 (N_7829,N_6276,N_6929);
nand U7830 (N_7830,N_6538,N_6469);
xor U7831 (N_7831,N_6386,N_6412);
xor U7832 (N_7832,N_6982,N_6189);
and U7833 (N_7833,N_6298,N_6582);
nor U7834 (N_7834,N_6023,N_6106);
and U7835 (N_7835,N_6354,N_6340);
xnor U7836 (N_7836,N_6991,N_6489);
or U7837 (N_7837,N_6437,N_6632);
xnor U7838 (N_7838,N_6287,N_6169);
or U7839 (N_7839,N_6088,N_6443);
nand U7840 (N_7840,N_6189,N_6725);
or U7841 (N_7841,N_6977,N_6056);
nor U7842 (N_7842,N_6676,N_6871);
and U7843 (N_7843,N_6281,N_6123);
nand U7844 (N_7844,N_6352,N_6564);
and U7845 (N_7845,N_6040,N_6033);
nand U7846 (N_7846,N_6741,N_6374);
nor U7847 (N_7847,N_6969,N_6386);
xor U7848 (N_7848,N_6598,N_6704);
nor U7849 (N_7849,N_6815,N_6785);
and U7850 (N_7850,N_6169,N_6770);
nand U7851 (N_7851,N_6087,N_6261);
xnor U7852 (N_7852,N_6754,N_6550);
or U7853 (N_7853,N_6426,N_6799);
or U7854 (N_7854,N_6355,N_6286);
nor U7855 (N_7855,N_6822,N_6534);
or U7856 (N_7856,N_6182,N_6048);
nand U7857 (N_7857,N_6368,N_6001);
nor U7858 (N_7858,N_6870,N_6134);
and U7859 (N_7859,N_6720,N_6793);
or U7860 (N_7860,N_6344,N_6040);
nor U7861 (N_7861,N_6934,N_6460);
or U7862 (N_7862,N_6008,N_6637);
xnor U7863 (N_7863,N_6719,N_6937);
nand U7864 (N_7864,N_6982,N_6072);
nand U7865 (N_7865,N_6501,N_6353);
or U7866 (N_7866,N_6828,N_6621);
and U7867 (N_7867,N_6695,N_6872);
and U7868 (N_7868,N_6176,N_6826);
xor U7869 (N_7869,N_6370,N_6188);
nand U7870 (N_7870,N_6259,N_6751);
or U7871 (N_7871,N_6925,N_6236);
xnor U7872 (N_7872,N_6332,N_6696);
nor U7873 (N_7873,N_6553,N_6332);
nor U7874 (N_7874,N_6104,N_6504);
and U7875 (N_7875,N_6654,N_6578);
nand U7876 (N_7876,N_6067,N_6653);
nor U7877 (N_7877,N_6138,N_6675);
or U7878 (N_7878,N_6970,N_6727);
and U7879 (N_7879,N_6634,N_6823);
and U7880 (N_7880,N_6516,N_6648);
nor U7881 (N_7881,N_6258,N_6800);
xnor U7882 (N_7882,N_6849,N_6206);
nor U7883 (N_7883,N_6526,N_6267);
nand U7884 (N_7884,N_6055,N_6248);
nor U7885 (N_7885,N_6519,N_6939);
or U7886 (N_7886,N_6823,N_6063);
xnor U7887 (N_7887,N_6510,N_6292);
nor U7888 (N_7888,N_6030,N_6407);
nand U7889 (N_7889,N_6466,N_6330);
nor U7890 (N_7890,N_6705,N_6805);
nor U7891 (N_7891,N_6319,N_6498);
nor U7892 (N_7892,N_6419,N_6913);
nand U7893 (N_7893,N_6761,N_6611);
and U7894 (N_7894,N_6435,N_6618);
nor U7895 (N_7895,N_6233,N_6368);
xnor U7896 (N_7896,N_6228,N_6666);
or U7897 (N_7897,N_6687,N_6378);
nor U7898 (N_7898,N_6642,N_6230);
nor U7899 (N_7899,N_6381,N_6659);
xnor U7900 (N_7900,N_6263,N_6492);
nor U7901 (N_7901,N_6761,N_6623);
and U7902 (N_7902,N_6240,N_6801);
nand U7903 (N_7903,N_6547,N_6476);
or U7904 (N_7904,N_6922,N_6711);
nor U7905 (N_7905,N_6461,N_6846);
xor U7906 (N_7906,N_6115,N_6177);
nand U7907 (N_7907,N_6237,N_6366);
and U7908 (N_7908,N_6271,N_6770);
or U7909 (N_7909,N_6655,N_6953);
nand U7910 (N_7910,N_6099,N_6277);
nand U7911 (N_7911,N_6760,N_6863);
nor U7912 (N_7912,N_6059,N_6359);
and U7913 (N_7913,N_6522,N_6331);
nand U7914 (N_7914,N_6996,N_6628);
xor U7915 (N_7915,N_6773,N_6382);
nor U7916 (N_7916,N_6500,N_6817);
and U7917 (N_7917,N_6205,N_6389);
nand U7918 (N_7918,N_6978,N_6092);
xor U7919 (N_7919,N_6845,N_6699);
and U7920 (N_7920,N_6731,N_6604);
or U7921 (N_7921,N_6815,N_6344);
nor U7922 (N_7922,N_6015,N_6002);
nand U7923 (N_7923,N_6684,N_6462);
nor U7924 (N_7924,N_6602,N_6862);
and U7925 (N_7925,N_6196,N_6819);
nand U7926 (N_7926,N_6015,N_6993);
nand U7927 (N_7927,N_6173,N_6296);
nor U7928 (N_7928,N_6172,N_6763);
or U7929 (N_7929,N_6161,N_6776);
or U7930 (N_7930,N_6690,N_6323);
xor U7931 (N_7931,N_6585,N_6539);
and U7932 (N_7932,N_6471,N_6816);
nand U7933 (N_7933,N_6814,N_6885);
nand U7934 (N_7934,N_6781,N_6462);
nand U7935 (N_7935,N_6190,N_6774);
xnor U7936 (N_7936,N_6167,N_6183);
or U7937 (N_7937,N_6920,N_6608);
nor U7938 (N_7938,N_6244,N_6648);
nand U7939 (N_7939,N_6299,N_6551);
or U7940 (N_7940,N_6788,N_6916);
or U7941 (N_7941,N_6801,N_6025);
nor U7942 (N_7942,N_6348,N_6844);
nand U7943 (N_7943,N_6910,N_6937);
and U7944 (N_7944,N_6088,N_6507);
nand U7945 (N_7945,N_6434,N_6066);
nand U7946 (N_7946,N_6602,N_6406);
or U7947 (N_7947,N_6843,N_6124);
nor U7948 (N_7948,N_6196,N_6984);
or U7949 (N_7949,N_6341,N_6014);
and U7950 (N_7950,N_6251,N_6630);
nor U7951 (N_7951,N_6494,N_6132);
xnor U7952 (N_7952,N_6266,N_6347);
or U7953 (N_7953,N_6154,N_6572);
xnor U7954 (N_7954,N_6100,N_6517);
xnor U7955 (N_7955,N_6331,N_6981);
or U7956 (N_7956,N_6988,N_6511);
and U7957 (N_7957,N_6956,N_6084);
nor U7958 (N_7958,N_6244,N_6070);
nand U7959 (N_7959,N_6243,N_6355);
nor U7960 (N_7960,N_6258,N_6092);
nor U7961 (N_7961,N_6636,N_6085);
xor U7962 (N_7962,N_6410,N_6748);
xnor U7963 (N_7963,N_6375,N_6742);
nand U7964 (N_7964,N_6985,N_6536);
xor U7965 (N_7965,N_6413,N_6071);
nand U7966 (N_7966,N_6792,N_6675);
nand U7967 (N_7967,N_6556,N_6547);
nor U7968 (N_7968,N_6303,N_6642);
and U7969 (N_7969,N_6298,N_6577);
nand U7970 (N_7970,N_6191,N_6806);
xor U7971 (N_7971,N_6233,N_6249);
xnor U7972 (N_7972,N_6346,N_6231);
nand U7973 (N_7973,N_6652,N_6892);
xor U7974 (N_7974,N_6410,N_6783);
xnor U7975 (N_7975,N_6909,N_6370);
xor U7976 (N_7976,N_6853,N_6259);
or U7977 (N_7977,N_6520,N_6308);
or U7978 (N_7978,N_6634,N_6389);
and U7979 (N_7979,N_6745,N_6575);
xnor U7980 (N_7980,N_6822,N_6106);
and U7981 (N_7981,N_6641,N_6866);
nor U7982 (N_7982,N_6846,N_6069);
xnor U7983 (N_7983,N_6559,N_6329);
or U7984 (N_7984,N_6240,N_6024);
nand U7985 (N_7985,N_6542,N_6675);
xor U7986 (N_7986,N_6756,N_6233);
nand U7987 (N_7987,N_6390,N_6280);
xor U7988 (N_7988,N_6544,N_6127);
and U7989 (N_7989,N_6807,N_6100);
or U7990 (N_7990,N_6850,N_6475);
and U7991 (N_7991,N_6478,N_6713);
nor U7992 (N_7992,N_6176,N_6573);
xnor U7993 (N_7993,N_6261,N_6218);
nand U7994 (N_7994,N_6296,N_6043);
or U7995 (N_7995,N_6038,N_6580);
and U7996 (N_7996,N_6839,N_6245);
nand U7997 (N_7997,N_6519,N_6521);
or U7998 (N_7998,N_6486,N_6217);
and U7999 (N_7999,N_6777,N_6868);
nand U8000 (N_8000,N_7635,N_7498);
nor U8001 (N_8001,N_7594,N_7547);
xnor U8002 (N_8002,N_7868,N_7837);
or U8003 (N_8003,N_7394,N_7926);
nand U8004 (N_8004,N_7006,N_7095);
or U8005 (N_8005,N_7137,N_7172);
nand U8006 (N_8006,N_7236,N_7354);
nand U8007 (N_8007,N_7412,N_7264);
and U8008 (N_8008,N_7950,N_7010);
and U8009 (N_8009,N_7748,N_7334);
nor U8010 (N_8010,N_7793,N_7364);
nand U8011 (N_8011,N_7618,N_7734);
nand U8012 (N_8012,N_7338,N_7715);
xor U8013 (N_8013,N_7575,N_7516);
nand U8014 (N_8014,N_7130,N_7708);
or U8015 (N_8015,N_7439,N_7343);
nor U8016 (N_8016,N_7487,N_7819);
nand U8017 (N_8017,N_7987,N_7102);
nand U8018 (N_8018,N_7722,N_7884);
or U8019 (N_8019,N_7918,N_7802);
nor U8020 (N_8020,N_7815,N_7320);
nor U8021 (N_8021,N_7899,N_7216);
nand U8022 (N_8022,N_7108,N_7652);
and U8023 (N_8023,N_7864,N_7000);
and U8024 (N_8024,N_7304,N_7692);
xnor U8025 (N_8025,N_7186,N_7224);
nand U8026 (N_8026,N_7639,N_7818);
and U8027 (N_8027,N_7374,N_7340);
nand U8028 (N_8028,N_7174,N_7291);
or U8029 (N_8029,N_7105,N_7564);
and U8030 (N_8030,N_7629,N_7830);
nand U8031 (N_8031,N_7984,N_7156);
and U8032 (N_8032,N_7290,N_7164);
or U8033 (N_8033,N_7346,N_7128);
nand U8034 (N_8034,N_7576,N_7067);
or U8035 (N_8035,N_7201,N_7424);
nand U8036 (N_8036,N_7182,N_7154);
and U8037 (N_8037,N_7359,N_7155);
nor U8038 (N_8038,N_7508,N_7854);
or U8039 (N_8039,N_7740,N_7180);
xnor U8040 (N_8040,N_7751,N_7103);
xnor U8041 (N_8041,N_7045,N_7968);
nor U8042 (N_8042,N_7245,N_7727);
xnor U8043 (N_8043,N_7525,N_7608);
or U8044 (N_8044,N_7914,N_7349);
and U8045 (N_8045,N_7044,N_7367);
or U8046 (N_8046,N_7408,N_7161);
and U8047 (N_8047,N_7702,N_7824);
nor U8048 (N_8048,N_7631,N_7726);
nand U8049 (N_8049,N_7207,N_7641);
or U8050 (N_8050,N_7556,N_7669);
nor U8051 (N_8051,N_7241,N_7765);
and U8052 (N_8052,N_7170,N_7462);
nor U8053 (N_8053,N_7208,N_7901);
and U8054 (N_8054,N_7870,N_7780);
or U8055 (N_8055,N_7535,N_7256);
and U8056 (N_8056,N_7269,N_7150);
nand U8057 (N_8057,N_7686,N_7324);
and U8058 (N_8058,N_7568,N_7299);
xor U8059 (N_8059,N_7147,N_7413);
or U8060 (N_8060,N_7353,N_7326);
nand U8061 (N_8061,N_7217,N_7856);
nor U8062 (N_8062,N_7709,N_7908);
or U8063 (N_8063,N_7943,N_7939);
nand U8064 (N_8064,N_7433,N_7769);
nand U8065 (N_8065,N_7764,N_7888);
nor U8066 (N_8066,N_7775,N_7087);
or U8067 (N_8067,N_7820,N_7716);
nor U8068 (N_8068,N_7379,N_7351);
xnor U8069 (N_8069,N_7557,N_7419);
or U8070 (N_8070,N_7430,N_7410);
nor U8071 (N_8071,N_7160,N_7991);
xor U8072 (N_8072,N_7975,N_7759);
or U8073 (N_8073,N_7074,N_7787);
and U8074 (N_8074,N_7189,N_7838);
nor U8075 (N_8075,N_7549,N_7925);
nand U8076 (N_8076,N_7491,N_7645);
or U8077 (N_8077,N_7676,N_7524);
nand U8078 (N_8078,N_7055,N_7121);
nor U8079 (N_8079,N_7052,N_7168);
nor U8080 (N_8080,N_7428,N_7502);
nor U8081 (N_8081,N_7347,N_7065);
xnor U8082 (N_8082,N_7276,N_7543);
nand U8083 (N_8083,N_7527,N_7792);
nand U8084 (N_8084,N_7331,N_7116);
and U8085 (N_8085,N_7546,N_7007);
or U8086 (N_8086,N_7386,N_7484);
and U8087 (N_8087,N_7931,N_7499);
nor U8088 (N_8088,N_7068,N_7253);
xnor U8089 (N_8089,N_7515,N_7021);
xor U8090 (N_8090,N_7570,N_7238);
or U8091 (N_8091,N_7849,N_7483);
nor U8092 (N_8092,N_7023,N_7265);
nand U8093 (N_8093,N_7595,N_7422);
nand U8094 (N_8094,N_7781,N_7619);
nand U8095 (N_8095,N_7418,N_7732);
nor U8096 (N_8096,N_7159,N_7192);
and U8097 (N_8097,N_7848,N_7625);
and U8098 (N_8098,N_7981,N_7202);
and U8099 (N_8099,N_7833,N_7047);
nor U8100 (N_8100,N_7505,N_7540);
nand U8101 (N_8101,N_7602,N_7393);
xnor U8102 (N_8102,N_7254,N_7784);
nor U8103 (N_8103,N_7513,N_7049);
nand U8104 (N_8104,N_7255,N_7048);
xor U8105 (N_8105,N_7778,N_7947);
and U8106 (N_8106,N_7902,N_7395);
nand U8107 (N_8107,N_7867,N_7736);
nand U8108 (N_8108,N_7341,N_7807);
nor U8109 (N_8109,N_7184,N_7800);
nand U8110 (N_8110,N_7927,N_7218);
and U8111 (N_8111,N_7531,N_7475);
xor U8112 (N_8112,N_7315,N_7919);
and U8113 (N_8113,N_7448,N_7081);
xnor U8114 (N_8114,N_7436,N_7753);
and U8115 (N_8115,N_7167,N_7243);
nor U8116 (N_8116,N_7437,N_7973);
and U8117 (N_8117,N_7398,N_7511);
and U8118 (N_8118,N_7790,N_7574);
or U8119 (N_8119,N_7881,N_7698);
xnor U8120 (N_8120,N_7431,N_7674);
nand U8121 (N_8121,N_7089,N_7879);
nor U8122 (N_8122,N_7034,N_7909);
or U8123 (N_8123,N_7522,N_7659);
and U8124 (N_8124,N_7666,N_7862);
or U8125 (N_8125,N_7670,N_7846);
xor U8126 (N_8126,N_7581,N_7385);
and U8127 (N_8127,N_7392,N_7730);
or U8128 (N_8128,N_7755,N_7944);
or U8129 (N_8129,N_7512,N_7969);
and U8130 (N_8130,N_7717,N_7391);
nor U8131 (N_8131,N_7898,N_7058);
nand U8132 (N_8132,N_7093,N_7417);
xnor U8133 (N_8133,N_7090,N_7539);
nor U8134 (N_8134,N_7965,N_7302);
or U8135 (N_8135,N_7173,N_7289);
or U8136 (N_8136,N_7681,N_7146);
nor U8137 (N_8137,N_7588,N_7565);
and U8138 (N_8138,N_7370,N_7195);
nor U8139 (N_8139,N_7980,N_7680);
or U8140 (N_8140,N_7053,N_7177);
or U8141 (N_8141,N_7024,N_7544);
xor U8142 (N_8142,N_7949,N_7842);
nor U8143 (N_8143,N_7012,N_7894);
nand U8144 (N_8144,N_7729,N_7876);
nand U8145 (N_8145,N_7008,N_7311);
nor U8146 (N_8146,N_7637,N_7163);
nor U8147 (N_8147,N_7310,N_7678);
nor U8148 (N_8148,N_7920,N_7528);
xor U8149 (N_8149,N_7461,N_7957);
nor U8150 (N_8150,N_7796,N_7697);
and U8151 (N_8151,N_7282,N_7069);
xnor U8152 (N_8152,N_7509,N_7518);
nor U8153 (N_8153,N_7280,N_7242);
and U8154 (N_8154,N_7750,N_7096);
nor U8155 (N_8155,N_7139,N_7963);
xor U8156 (N_8156,N_7695,N_7308);
and U8157 (N_8157,N_7136,N_7585);
or U8158 (N_8158,N_7803,N_7999);
and U8159 (N_8159,N_7259,N_7294);
xor U8160 (N_8160,N_7873,N_7257);
or U8161 (N_8161,N_7301,N_7450);
xor U8162 (N_8162,N_7878,N_7318);
or U8163 (N_8163,N_7636,N_7406);
or U8164 (N_8164,N_7688,N_7188);
nor U8165 (N_8165,N_7332,N_7384);
nand U8166 (N_8166,N_7996,N_7887);
nand U8167 (N_8167,N_7601,N_7651);
or U8168 (N_8168,N_7438,N_7832);
nand U8169 (N_8169,N_7454,N_7885);
xor U8170 (N_8170,N_7261,N_7123);
nand U8171 (N_8171,N_7031,N_7091);
nor U8172 (N_8172,N_7279,N_7587);
or U8173 (N_8173,N_7329,N_7169);
or U8174 (N_8174,N_7731,N_7610);
nor U8175 (N_8175,N_7986,N_7707);
xor U8176 (N_8176,N_7278,N_7883);
nor U8177 (N_8177,N_7300,N_7114);
xor U8178 (N_8178,N_7761,N_7911);
xor U8179 (N_8179,N_7490,N_7441);
and U8180 (N_8180,N_7791,N_7643);
or U8181 (N_8181,N_7628,N_7309);
or U8182 (N_8182,N_7689,N_7662);
and U8183 (N_8183,N_7344,N_7719);
nor U8184 (N_8184,N_7612,N_7162);
nor U8185 (N_8185,N_7977,N_7327);
or U8186 (N_8186,N_7009,N_7420);
or U8187 (N_8187,N_7252,N_7075);
nor U8188 (N_8188,N_7054,N_7039);
xnor U8189 (N_8189,N_7030,N_7569);
nand U8190 (N_8190,N_7325,N_7051);
xnor U8191 (N_8191,N_7953,N_7733);
xor U8192 (N_8192,N_7185,N_7768);
nor U8193 (N_8193,N_7232,N_7348);
xnor U8194 (N_8194,N_7725,N_7534);
xnor U8195 (N_8195,N_7572,N_7016);
xor U8196 (N_8196,N_7495,N_7665);
nor U8197 (N_8197,N_7801,N_7244);
nor U8198 (N_8198,N_7365,N_7917);
and U8199 (N_8199,N_7335,N_7703);
and U8200 (N_8200,N_7589,N_7964);
nand U8201 (N_8201,N_7827,N_7330);
and U8202 (N_8202,N_7855,N_7035);
or U8203 (N_8203,N_7743,N_7423);
nor U8204 (N_8204,N_7956,N_7099);
or U8205 (N_8205,N_7672,N_7798);
or U8206 (N_8206,N_7111,N_7647);
nor U8207 (N_8207,N_7584,N_7777);
and U8208 (N_8208,N_7464,N_7270);
or U8209 (N_8209,N_7101,N_7122);
or U8210 (N_8210,N_7550,N_7375);
nand U8211 (N_8211,N_7623,N_7193);
nand U8212 (N_8212,N_7795,N_7371);
and U8213 (N_8213,N_7215,N_7277);
xor U8214 (N_8214,N_7140,N_7882);
nor U8215 (N_8215,N_7656,N_7701);
nor U8216 (N_8216,N_7952,N_7083);
and U8217 (N_8217,N_7042,N_7357);
xor U8218 (N_8218,N_7851,N_7812);
and U8219 (N_8219,N_7135,N_7281);
and U8220 (N_8220,N_7298,N_7459);
nor U8221 (N_8221,N_7134,N_7541);
or U8222 (N_8222,N_7226,N_7283);
xnor U8223 (N_8223,N_7323,N_7403);
nand U8224 (N_8224,N_7025,N_7624);
nand U8225 (N_8225,N_7292,N_7814);
xor U8226 (N_8226,N_7985,N_7533);
or U8227 (N_8227,N_7852,N_7747);
and U8228 (N_8228,N_7994,N_7829);
or U8229 (N_8229,N_7721,N_7718);
or U8230 (N_8230,N_7275,N_7183);
or U8231 (N_8231,N_7860,N_7175);
xor U8232 (N_8232,N_7488,N_7032);
and U8233 (N_8233,N_7376,N_7124);
xnor U8234 (N_8234,N_7797,N_7445);
or U8235 (N_8235,N_7783,N_7492);
xor U8236 (N_8236,N_7249,N_7976);
or U8237 (N_8237,N_7699,N_7586);
or U8238 (N_8238,N_7094,N_7532);
nand U8239 (N_8239,N_7455,N_7735);
nand U8240 (N_8240,N_7724,N_7591);
and U8241 (N_8241,N_7457,N_7085);
nor U8242 (N_8242,N_7813,N_7897);
nor U8243 (N_8243,N_7033,N_7345);
nand U8244 (N_8244,N_7452,N_7080);
and U8245 (N_8245,N_7786,N_7003);
nand U8246 (N_8246,N_7421,N_7036);
or U8247 (N_8247,N_7482,N_7132);
nor U8248 (N_8248,N_7723,N_7714);
and U8249 (N_8249,N_7772,N_7517);
xnor U8250 (N_8250,N_7458,N_7928);
nor U8251 (N_8251,N_7079,N_7598);
xor U8252 (N_8252,N_7013,N_7191);
nand U8253 (N_8253,N_7397,N_7742);
xor U8254 (N_8254,N_7141,N_7014);
nor U8255 (N_8255,N_7213,N_7263);
nand U8256 (N_8256,N_7946,N_7836);
or U8257 (N_8257,N_7247,N_7131);
xnor U8258 (N_8258,N_7088,N_7683);
nor U8259 (N_8259,N_7650,N_7358);
and U8260 (N_8260,N_7138,N_7333);
and U8261 (N_8261,N_7178,N_7409);
nand U8262 (N_8262,N_7372,N_7041);
and U8263 (N_8263,N_7932,N_7231);
xnor U8264 (N_8264,N_7362,N_7523);
nand U8265 (N_8265,N_7655,N_7038);
and U8266 (N_8266,N_7223,N_7209);
nand U8267 (N_8267,N_7110,N_7297);
and U8268 (N_8268,N_7869,N_7799);
nor U8269 (N_8269,N_7305,N_7997);
and U8270 (N_8270,N_7577,N_7316);
xor U8271 (N_8271,N_7794,N_7766);
and U8272 (N_8272,N_7537,N_7640);
nor U8273 (N_8273,N_7107,N_7062);
or U8274 (N_8274,N_7339,N_7704);
or U8275 (N_8275,N_7366,N_7990);
and U8276 (N_8276,N_7858,N_7600);
nand U8277 (N_8277,N_7057,N_7971);
and U8278 (N_8278,N_7271,N_7649);
nor U8279 (N_8279,N_7447,N_7922);
xnor U8280 (N_8280,N_7506,N_7974);
xor U8281 (N_8281,N_7615,N_7056);
or U8282 (N_8282,N_7804,N_7738);
or U8283 (N_8283,N_7504,N_7966);
and U8284 (N_8284,N_7752,N_7028);
nand U8285 (N_8285,N_7720,N_7317);
xnor U8286 (N_8286,N_7235,N_7616);
or U8287 (N_8287,N_7446,N_7415);
nand U8288 (N_8288,N_7510,N_7696);
nor U8289 (N_8289,N_7171,N_7229);
nor U8290 (N_8290,N_7970,N_7176);
nor U8291 (N_8291,N_7507,N_7972);
or U8292 (N_8292,N_7501,N_7762);
nor U8293 (N_8293,N_7693,N_7387);
nor U8294 (N_8294,N_7620,N_7126);
or U8295 (N_8295,N_7782,N_7402);
xor U8296 (N_8296,N_7983,N_7097);
or U8297 (N_8297,N_7754,N_7978);
xor U8298 (N_8298,N_7043,N_7109);
and U8299 (N_8299,N_7467,N_7580);
xnor U8300 (N_8300,N_7773,N_7465);
nand U8301 (N_8301,N_7165,N_7685);
or U8302 (N_8302,N_7451,N_7893);
and U8303 (N_8303,N_7605,N_7880);
nor U8304 (N_8304,N_7040,N_7400);
xor U8305 (N_8305,N_7687,N_7660);
xnor U8306 (N_8306,N_7456,N_7352);
xnor U8307 (N_8307,N_7536,N_7874);
nand U8308 (N_8308,N_7166,N_7875);
nand U8309 (N_8309,N_7390,N_7248);
and U8310 (N_8310,N_7214,N_7383);
xor U8311 (N_8311,N_7789,N_7904);
and U8312 (N_8312,N_7921,N_7378);
and U8313 (N_8313,N_7225,N_7181);
nand U8314 (N_8314,N_7825,N_7200);
nand U8315 (N_8315,N_7633,N_7552);
and U8316 (N_8316,N_7322,N_7596);
or U8317 (N_8317,N_7388,N_7399);
or U8318 (N_8318,N_7210,N_7486);
nor U8319 (N_8319,N_7583,N_7896);
nand U8320 (N_8320,N_7788,N_7117);
nand U8321 (N_8321,N_7542,N_7839);
and U8322 (N_8322,N_7905,N_7015);
xor U8323 (N_8323,N_7503,N_7199);
nor U8324 (N_8324,N_7627,N_7816);
or U8325 (N_8325,N_7071,N_7551);
nand U8326 (N_8326,N_7470,N_7671);
and U8327 (N_8327,N_7453,N_7328);
and U8328 (N_8328,N_7287,N_7469);
xnor U8329 (N_8329,N_7196,N_7822);
or U8330 (N_8330,N_7479,N_7076);
xnor U8331 (N_8331,N_7350,N_7219);
and U8332 (N_8332,N_7757,N_7675);
or U8333 (N_8333,N_7712,N_7891);
nand U8334 (N_8334,N_7337,N_7942);
nand U8335 (N_8335,N_7648,N_7306);
xnor U8336 (N_8336,N_7363,N_7677);
or U8337 (N_8337,N_7250,N_7078);
nand U8338 (N_8338,N_7604,N_7405);
nand U8339 (N_8339,N_7653,N_7227);
xnor U8340 (N_8340,N_7237,N_7561);
nand U8341 (N_8341,N_7018,N_7113);
or U8342 (N_8342,N_7001,N_7857);
or U8343 (N_8343,N_7336,N_7937);
nand U8344 (N_8344,N_7027,N_7526);
nand U8345 (N_8345,N_7989,N_7285);
and U8346 (N_8346,N_7520,N_7554);
nor U8347 (N_8347,N_7916,N_7548);
nand U8348 (N_8348,N_7638,N_7466);
and U8349 (N_8349,N_7634,N_7037);
and U8350 (N_8350,N_7560,N_7260);
and U8351 (N_8351,N_7998,N_7861);
xor U8352 (N_8352,N_7940,N_7930);
and U8353 (N_8353,N_7617,N_7321);
nand U8354 (N_8354,N_7553,N_7945);
nand U8355 (N_8355,N_7204,N_7749);
or U8356 (N_8356,N_7485,N_7434);
and U8357 (N_8357,N_7120,N_7955);
or U8358 (N_8358,N_7959,N_7821);
xnor U8359 (N_8359,N_7579,N_7746);
xor U8360 (N_8360,N_7342,N_7086);
and U8361 (N_8361,N_7559,N_7737);
xor U8362 (N_8362,N_7481,N_7935);
nor U8363 (N_8363,N_7682,N_7545);
and U8364 (N_8364,N_7148,N_7658);
nor U8365 (N_8365,N_7050,N_7020);
xor U8366 (N_8366,N_7614,N_7070);
xnor U8367 (N_8367,N_7005,N_7145);
xnor U8368 (N_8368,N_7823,N_7691);
nor U8369 (N_8369,N_7234,N_7938);
and U8370 (N_8370,N_7562,N_7273);
or U8371 (N_8371,N_7826,N_7380);
nand U8372 (N_8372,N_7493,N_7149);
nor U8373 (N_8373,N_7877,N_7739);
nand U8374 (N_8374,N_7632,N_7115);
or U8375 (N_8375,N_7489,N_7473);
nand U8376 (N_8376,N_7142,N_7599);
xnor U8377 (N_8377,N_7098,N_7017);
xor U8378 (N_8378,N_7118,N_7144);
nand U8379 (N_8379,N_7924,N_7841);
nand U8380 (N_8380,N_7664,N_7295);
and U8381 (N_8381,N_7373,N_7060);
and U8382 (N_8382,N_7432,N_7496);
or U8383 (N_8383,N_7381,N_7603);
or U8384 (N_8384,N_7129,N_7845);
and U8385 (N_8385,N_7853,N_7514);
xnor U8386 (N_8386,N_7929,N_7190);
and U8387 (N_8387,N_7611,N_7258);
or U8388 (N_8388,N_7831,N_7694);
nand U8389 (N_8389,N_7889,N_7004);
nand U8390 (N_8390,N_7106,N_7785);
and U8391 (N_8391,N_7377,N_7770);
nand U8392 (N_8392,N_7444,N_7361);
nor U8393 (N_8393,N_7900,N_7435);
or U8394 (N_8394,N_7988,N_7356);
and U8395 (N_8395,N_7205,N_7133);
nor U8396 (N_8396,N_7679,N_7871);
xor U8397 (N_8397,N_7239,N_7745);
xnor U8398 (N_8398,N_7886,N_7982);
nand U8399 (N_8399,N_7396,N_7002);
nor U8400 (N_8400,N_7153,N_7936);
nor U8401 (N_8401,N_7472,N_7859);
or U8402 (N_8402,N_7630,N_7840);
nand U8403 (N_8403,N_7756,N_7157);
nand U8404 (N_8404,N_7828,N_7808);
and U8405 (N_8405,N_7497,N_7246);
or U8406 (N_8406,N_7810,N_7847);
and U8407 (N_8407,N_7892,N_7642);
xnor U8408 (N_8408,N_7179,N_7646);
or U8409 (N_8409,N_7026,N_7284);
or U8410 (N_8410,N_7092,N_7834);
or U8411 (N_8411,N_7890,N_7233);
and U8412 (N_8412,N_7425,N_7519);
nor U8413 (N_8413,N_7104,N_7314);
xor U8414 (N_8414,N_7059,N_7654);
or U8415 (N_8415,N_7622,N_7319);
and U8416 (N_8416,N_7303,N_7268);
nand U8417 (N_8417,N_7913,N_7460);
xnor U8418 (N_8418,N_7606,N_7573);
or U8419 (N_8419,N_7613,N_7066);
nor U8420 (N_8420,N_7993,N_7084);
or U8421 (N_8421,N_7771,N_7933);
xor U8422 (N_8422,N_7073,N_7401);
xnor U8423 (N_8423,N_7835,N_7474);
nor U8424 (N_8424,N_7872,N_7463);
nand U8425 (N_8425,N_7267,N_7843);
and U8426 (N_8426,N_7863,N_7806);
nand U8427 (N_8427,N_7072,N_7151);
and U8428 (N_8428,N_7476,N_7844);
xnor U8429 (N_8429,N_7061,N_7941);
nand U8430 (N_8430,N_7954,N_7906);
nand U8431 (N_8431,N_7220,N_7728);
xnor U8432 (N_8432,N_7212,N_7592);
nand U8433 (N_8433,N_7776,N_7805);
xnor U8434 (N_8434,N_7426,N_7915);
and U8435 (N_8435,N_7995,N_7571);
and U8436 (N_8436,N_7626,N_7684);
nand U8437 (N_8437,N_7152,N_7382);
or U8438 (N_8438,N_7661,N_7673);
nand U8439 (N_8439,N_7979,N_7779);
and U8440 (N_8440,N_7198,N_7538);
and U8441 (N_8441,N_7700,N_7850);
and U8442 (N_8442,N_7230,N_7077);
or U8443 (N_8443,N_7609,N_7910);
nand U8444 (N_8444,N_7967,N_7961);
xnor U8445 (N_8445,N_7019,N_7567);
nand U8446 (N_8446,N_7480,N_7029);
nor U8447 (N_8447,N_7407,N_7923);
and U8448 (N_8448,N_7710,N_7369);
or U8449 (N_8449,N_7865,N_7607);
or U8450 (N_8450,N_7228,N_7951);
nand U8451 (N_8451,N_7934,N_7558);
or U8452 (N_8452,N_7948,N_7760);
nand U8453 (N_8453,N_7266,N_7296);
nor U8454 (N_8454,N_7763,N_7866);
nand U8455 (N_8455,N_7962,N_7063);
and U8456 (N_8456,N_7644,N_7590);
or U8457 (N_8457,N_7443,N_7203);
or U8458 (N_8458,N_7411,N_7706);
and U8459 (N_8459,N_7194,N_7667);
nor U8460 (N_8460,N_7529,N_7197);
nand U8461 (N_8461,N_7471,N_7240);
nand U8462 (N_8462,N_7125,N_7811);
or U8463 (N_8463,N_7500,N_7817);
and U8464 (N_8464,N_7912,N_7578);
and U8465 (N_8465,N_7758,N_7100);
and U8466 (N_8466,N_7442,N_7705);
xor U8467 (N_8467,N_7668,N_7530);
nand U8468 (N_8468,N_7206,N_7468);
and U8469 (N_8469,N_7690,N_7022);
and U8470 (N_8470,N_7360,N_7274);
xor U8471 (N_8471,N_7355,N_7158);
nor U8472 (N_8472,N_7449,N_7414);
nor U8473 (N_8473,N_7221,N_7429);
nor U8474 (N_8474,N_7494,N_7416);
nor U8475 (N_8475,N_7774,N_7809);
nand U8476 (N_8476,N_7389,N_7082);
nor U8477 (N_8477,N_7663,N_7046);
or U8478 (N_8478,N_7477,N_7286);
xor U8479 (N_8479,N_7143,N_7211);
or U8480 (N_8480,N_7440,N_7744);
nor U8481 (N_8481,N_7272,N_7119);
nand U8482 (N_8482,N_7288,N_7907);
nand U8483 (N_8483,N_7251,N_7992);
nand U8484 (N_8484,N_7566,N_7427);
nand U8485 (N_8485,N_7307,N_7582);
nand U8486 (N_8486,N_7555,N_7011);
or U8487 (N_8487,N_7895,N_7127);
xor U8488 (N_8488,N_7621,N_7478);
nand U8489 (N_8489,N_7222,N_7521);
or U8490 (N_8490,N_7312,N_7711);
xor U8491 (N_8491,N_7112,N_7368);
and U8492 (N_8492,N_7767,N_7313);
or U8493 (N_8493,N_7262,N_7657);
nor U8494 (N_8494,N_7187,N_7958);
and U8495 (N_8495,N_7903,N_7597);
xor U8496 (N_8496,N_7293,N_7741);
or U8497 (N_8497,N_7960,N_7593);
nand U8498 (N_8498,N_7713,N_7404);
and U8499 (N_8499,N_7064,N_7563);
xor U8500 (N_8500,N_7434,N_7569);
xor U8501 (N_8501,N_7108,N_7150);
and U8502 (N_8502,N_7201,N_7369);
and U8503 (N_8503,N_7822,N_7204);
xor U8504 (N_8504,N_7563,N_7685);
nor U8505 (N_8505,N_7645,N_7338);
nor U8506 (N_8506,N_7482,N_7947);
nor U8507 (N_8507,N_7155,N_7726);
nor U8508 (N_8508,N_7351,N_7870);
and U8509 (N_8509,N_7177,N_7396);
nor U8510 (N_8510,N_7904,N_7951);
nand U8511 (N_8511,N_7061,N_7859);
or U8512 (N_8512,N_7681,N_7534);
nand U8513 (N_8513,N_7526,N_7044);
or U8514 (N_8514,N_7051,N_7232);
nor U8515 (N_8515,N_7823,N_7318);
and U8516 (N_8516,N_7036,N_7561);
xnor U8517 (N_8517,N_7214,N_7861);
or U8518 (N_8518,N_7576,N_7802);
nor U8519 (N_8519,N_7156,N_7926);
or U8520 (N_8520,N_7629,N_7551);
and U8521 (N_8521,N_7747,N_7715);
nor U8522 (N_8522,N_7222,N_7846);
nand U8523 (N_8523,N_7284,N_7814);
xnor U8524 (N_8524,N_7512,N_7001);
and U8525 (N_8525,N_7114,N_7149);
nand U8526 (N_8526,N_7217,N_7929);
or U8527 (N_8527,N_7589,N_7549);
and U8528 (N_8528,N_7145,N_7865);
or U8529 (N_8529,N_7327,N_7078);
nand U8530 (N_8530,N_7447,N_7046);
nor U8531 (N_8531,N_7838,N_7631);
xnor U8532 (N_8532,N_7797,N_7361);
nor U8533 (N_8533,N_7254,N_7298);
or U8534 (N_8534,N_7166,N_7036);
nand U8535 (N_8535,N_7952,N_7354);
xnor U8536 (N_8536,N_7251,N_7054);
and U8537 (N_8537,N_7476,N_7033);
nor U8538 (N_8538,N_7163,N_7935);
nor U8539 (N_8539,N_7413,N_7778);
nand U8540 (N_8540,N_7757,N_7894);
or U8541 (N_8541,N_7559,N_7058);
and U8542 (N_8542,N_7894,N_7473);
and U8543 (N_8543,N_7115,N_7198);
xor U8544 (N_8544,N_7153,N_7086);
nor U8545 (N_8545,N_7013,N_7048);
or U8546 (N_8546,N_7538,N_7259);
xnor U8547 (N_8547,N_7806,N_7240);
xor U8548 (N_8548,N_7687,N_7709);
nor U8549 (N_8549,N_7075,N_7200);
or U8550 (N_8550,N_7442,N_7217);
nand U8551 (N_8551,N_7462,N_7211);
xnor U8552 (N_8552,N_7362,N_7516);
or U8553 (N_8553,N_7190,N_7632);
and U8554 (N_8554,N_7392,N_7504);
nand U8555 (N_8555,N_7198,N_7933);
xnor U8556 (N_8556,N_7544,N_7428);
nand U8557 (N_8557,N_7318,N_7660);
or U8558 (N_8558,N_7734,N_7662);
nor U8559 (N_8559,N_7900,N_7743);
nor U8560 (N_8560,N_7037,N_7006);
and U8561 (N_8561,N_7718,N_7167);
or U8562 (N_8562,N_7216,N_7099);
nand U8563 (N_8563,N_7625,N_7750);
xnor U8564 (N_8564,N_7661,N_7871);
and U8565 (N_8565,N_7541,N_7035);
and U8566 (N_8566,N_7566,N_7026);
nor U8567 (N_8567,N_7151,N_7602);
and U8568 (N_8568,N_7182,N_7599);
nand U8569 (N_8569,N_7825,N_7394);
nand U8570 (N_8570,N_7814,N_7394);
nand U8571 (N_8571,N_7038,N_7235);
nand U8572 (N_8572,N_7810,N_7064);
or U8573 (N_8573,N_7691,N_7525);
or U8574 (N_8574,N_7841,N_7036);
and U8575 (N_8575,N_7456,N_7340);
nand U8576 (N_8576,N_7036,N_7928);
and U8577 (N_8577,N_7422,N_7114);
nand U8578 (N_8578,N_7322,N_7150);
nor U8579 (N_8579,N_7879,N_7070);
xnor U8580 (N_8580,N_7016,N_7637);
nand U8581 (N_8581,N_7746,N_7816);
nor U8582 (N_8582,N_7318,N_7223);
or U8583 (N_8583,N_7358,N_7993);
xnor U8584 (N_8584,N_7755,N_7629);
and U8585 (N_8585,N_7788,N_7977);
xor U8586 (N_8586,N_7018,N_7030);
and U8587 (N_8587,N_7970,N_7544);
nand U8588 (N_8588,N_7362,N_7359);
xor U8589 (N_8589,N_7794,N_7044);
nor U8590 (N_8590,N_7571,N_7607);
or U8591 (N_8591,N_7226,N_7467);
and U8592 (N_8592,N_7106,N_7479);
xnor U8593 (N_8593,N_7991,N_7479);
or U8594 (N_8594,N_7381,N_7359);
nor U8595 (N_8595,N_7774,N_7090);
and U8596 (N_8596,N_7998,N_7176);
or U8597 (N_8597,N_7308,N_7495);
nand U8598 (N_8598,N_7000,N_7669);
xor U8599 (N_8599,N_7636,N_7655);
nor U8600 (N_8600,N_7265,N_7570);
nor U8601 (N_8601,N_7939,N_7778);
and U8602 (N_8602,N_7781,N_7035);
or U8603 (N_8603,N_7133,N_7316);
nand U8604 (N_8604,N_7277,N_7890);
nor U8605 (N_8605,N_7936,N_7724);
nand U8606 (N_8606,N_7336,N_7620);
xor U8607 (N_8607,N_7596,N_7412);
xnor U8608 (N_8608,N_7816,N_7751);
nor U8609 (N_8609,N_7147,N_7781);
xnor U8610 (N_8610,N_7853,N_7064);
nand U8611 (N_8611,N_7041,N_7928);
xnor U8612 (N_8612,N_7676,N_7642);
nor U8613 (N_8613,N_7539,N_7810);
nor U8614 (N_8614,N_7820,N_7457);
nand U8615 (N_8615,N_7747,N_7876);
nor U8616 (N_8616,N_7385,N_7144);
and U8617 (N_8617,N_7917,N_7581);
nand U8618 (N_8618,N_7082,N_7564);
nor U8619 (N_8619,N_7592,N_7321);
xnor U8620 (N_8620,N_7676,N_7171);
and U8621 (N_8621,N_7612,N_7340);
xor U8622 (N_8622,N_7831,N_7274);
and U8623 (N_8623,N_7121,N_7119);
nor U8624 (N_8624,N_7640,N_7313);
or U8625 (N_8625,N_7092,N_7084);
or U8626 (N_8626,N_7037,N_7762);
nor U8627 (N_8627,N_7751,N_7036);
and U8628 (N_8628,N_7358,N_7625);
or U8629 (N_8629,N_7895,N_7833);
nand U8630 (N_8630,N_7057,N_7661);
nor U8631 (N_8631,N_7634,N_7238);
or U8632 (N_8632,N_7325,N_7904);
or U8633 (N_8633,N_7362,N_7061);
nor U8634 (N_8634,N_7998,N_7033);
nand U8635 (N_8635,N_7366,N_7017);
xor U8636 (N_8636,N_7066,N_7672);
and U8637 (N_8637,N_7963,N_7364);
and U8638 (N_8638,N_7567,N_7501);
nand U8639 (N_8639,N_7099,N_7736);
and U8640 (N_8640,N_7443,N_7694);
nor U8641 (N_8641,N_7449,N_7204);
or U8642 (N_8642,N_7854,N_7175);
nor U8643 (N_8643,N_7884,N_7796);
and U8644 (N_8644,N_7094,N_7420);
and U8645 (N_8645,N_7060,N_7479);
or U8646 (N_8646,N_7059,N_7735);
nand U8647 (N_8647,N_7065,N_7350);
and U8648 (N_8648,N_7032,N_7540);
nor U8649 (N_8649,N_7171,N_7460);
nand U8650 (N_8650,N_7488,N_7184);
and U8651 (N_8651,N_7492,N_7862);
and U8652 (N_8652,N_7737,N_7451);
and U8653 (N_8653,N_7698,N_7660);
or U8654 (N_8654,N_7488,N_7482);
nand U8655 (N_8655,N_7915,N_7802);
nor U8656 (N_8656,N_7814,N_7609);
nor U8657 (N_8657,N_7735,N_7711);
xor U8658 (N_8658,N_7424,N_7308);
or U8659 (N_8659,N_7442,N_7518);
and U8660 (N_8660,N_7303,N_7946);
or U8661 (N_8661,N_7675,N_7537);
xor U8662 (N_8662,N_7091,N_7838);
and U8663 (N_8663,N_7571,N_7566);
and U8664 (N_8664,N_7704,N_7669);
or U8665 (N_8665,N_7946,N_7821);
xor U8666 (N_8666,N_7730,N_7617);
and U8667 (N_8667,N_7503,N_7720);
nor U8668 (N_8668,N_7178,N_7356);
or U8669 (N_8669,N_7171,N_7494);
nand U8670 (N_8670,N_7882,N_7765);
xor U8671 (N_8671,N_7503,N_7285);
and U8672 (N_8672,N_7667,N_7354);
xnor U8673 (N_8673,N_7944,N_7771);
and U8674 (N_8674,N_7152,N_7793);
or U8675 (N_8675,N_7799,N_7473);
and U8676 (N_8676,N_7009,N_7356);
nor U8677 (N_8677,N_7598,N_7421);
nand U8678 (N_8678,N_7629,N_7603);
nor U8679 (N_8679,N_7837,N_7547);
nand U8680 (N_8680,N_7527,N_7020);
nor U8681 (N_8681,N_7815,N_7448);
and U8682 (N_8682,N_7597,N_7495);
nand U8683 (N_8683,N_7621,N_7118);
nand U8684 (N_8684,N_7013,N_7957);
xor U8685 (N_8685,N_7525,N_7886);
nand U8686 (N_8686,N_7296,N_7462);
and U8687 (N_8687,N_7110,N_7253);
nor U8688 (N_8688,N_7387,N_7803);
or U8689 (N_8689,N_7796,N_7687);
nand U8690 (N_8690,N_7209,N_7465);
xnor U8691 (N_8691,N_7799,N_7588);
xor U8692 (N_8692,N_7505,N_7904);
and U8693 (N_8693,N_7244,N_7953);
or U8694 (N_8694,N_7832,N_7082);
or U8695 (N_8695,N_7655,N_7768);
nand U8696 (N_8696,N_7236,N_7155);
nand U8697 (N_8697,N_7254,N_7583);
and U8698 (N_8698,N_7805,N_7257);
or U8699 (N_8699,N_7212,N_7144);
nor U8700 (N_8700,N_7103,N_7042);
nand U8701 (N_8701,N_7490,N_7294);
xnor U8702 (N_8702,N_7089,N_7892);
nor U8703 (N_8703,N_7255,N_7007);
xnor U8704 (N_8704,N_7372,N_7495);
nor U8705 (N_8705,N_7556,N_7691);
nand U8706 (N_8706,N_7676,N_7913);
nand U8707 (N_8707,N_7005,N_7047);
and U8708 (N_8708,N_7591,N_7128);
and U8709 (N_8709,N_7288,N_7098);
xnor U8710 (N_8710,N_7034,N_7540);
nand U8711 (N_8711,N_7452,N_7657);
xnor U8712 (N_8712,N_7461,N_7685);
nand U8713 (N_8713,N_7227,N_7477);
xnor U8714 (N_8714,N_7635,N_7699);
and U8715 (N_8715,N_7479,N_7799);
or U8716 (N_8716,N_7028,N_7153);
nand U8717 (N_8717,N_7997,N_7931);
or U8718 (N_8718,N_7299,N_7049);
nor U8719 (N_8719,N_7566,N_7052);
nand U8720 (N_8720,N_7813,N_7004);
or U8721 (N_8721,N_7308,N_7627);
and U8722 (N_8722,N_7187,N_7562);
and U8723 (N_8723,N_7515,N_7882);
xnor U8724 (N_8724,N_7774,N_7338);
nand U8725 (N_8725,N_7002,N_7959);
or U8726 (N_8726,N_7556,N_7111);
xor U8727 (N_8727,N_7208,N_7373);
nor U8728 (N_8728,N_7005,N_7224);
and U8729 (N_8729,N_7149,N_7612);
nor U8730 (N_8730,N_7085,N_7733);
nand U8731 (N_8731,N_7686,N_7304);
or U8732 (N_8732,N_7365,N_7444);
nand U8733 (N_8733,N_7787,N_7458);
xnor U8734 (N_8734,N_7722,N_7181);
and U8735 (N_8735,N_7847,N_7603);
xnor U8736 (N_8736,N_7689,N_7319);
or U8737 (N_8737,N_7970,N_7815);
xnor U8738 (N_8738,N_7957,N_7773);
xor U8739 (N_8739,N_7564,N_7897);
nor U8740 (N_8740,N_7374,N_7774);
nor U8741 (N_8741,N_7565,N_7283);
nor U8742 (N_8742,N_7988,N_7328);
and U8743 (N_8743,N_7593,N_7531);
or U8744 (N_8744,N_7537,N_7163);
or U8745 (N_8745,N_7984,N_7348);
xor U8746 (N_8746,N_7746,N_7709);
or U8747 (N_8747,N_7046,N_7366);
nand U8748 (N_8748,N_7839,N_7508);
xor U8749 (N_8749,N_7421,N_7738);
or U8750 (N_8750,N_7369,N_7357);
nor U8751 (N_8751,N_7150,N_7129);
or U8752 (N_8752,N_7762,N_7990);
or U8753 (N_8753,N_7705,N_7037);
or U8754 (N_8754,N_7959,N_7717);
nand U8755 (N_8755,N_7646,N_7094);
and U8756 (N_8756,N_7847,N_7660);
nor U8757 (N_8757,N_7629,N_7161);
and U8758 (N_8758,N_7858,N_7523);
and U8759 (N_8759,N_7219,N_7704);
xor U8760 (N_8760,N_7064,N_7102);
or U8761 (N_8761,N_7301,N_7795);
or U8762 (N_8762,N_7982,N_7639);
and U8763 (N_8763,N_7682,N_7850);
and U8764 (N_8764,N_7217,N_7257);
nor U8765 (N_8765,N_7138,N_7794);
nor U8766 (N_8766,N_7071,N_7599);
nand U8767 (N_8767,N_7713,N_7690);
or U8768 (N_8768,N_7453,N_7452);
nand U8769 (N_8769,N_7657,N_7781);
or U8770 (N_8770,N_7642,N_7241);
and U8771 (N_8771,N_7454,N_7934);
and U8772 (N_8772,N_7631,N_7691);
or U8773 (N_8773,N_7693,N_7398);
and U8774 (N_8774,N_7959,N_7425);
xnor U8775 (N_8775,N_7487,N_7284);
nor U8776 (N_8776,N_7819,N_7496);
nor U8777 (N_8777,N_7749,N_7447);
or U8778 (N_8778,N_7931,N_7297);
xor U8779 (N_8779,N_7620,N_7380);
nand U8780 (N_8780,N_7723,N_7757);
nand U8781 (N_8781,N_7864,N_7955);
and U8782 (N_8782,N_7219,N_7970);
nor U8783 (N_8783,N_7973,N_7314);
xnor U8784 (N_8784,N_7592,N_7677);
and U8785 (N_8785,N_7453,N_7350);
xor U8786 (N_8786,N_7014,N_7482);
nor U8787 (N_8787,N_7262,N_7182);
and U8788 (N_8788,N_7381,N_7334);
or U8789 (N_8789,N_7248,N_7661);
or U8790 (N_8790,N_7159,N_7869);
nor U8791 (N_8791,N_7122,N_7291);
and U8792 (N_8792,N_7012,N_7162);
nor U8793 (N_8793,N_7040,N_7620);
xnor U8794 (N_8794,N_7827,N_7966);
and U8795 (N_8795,N_7350,N_7381);
xnor U8796 (N_8796,N_7551,N_7085);
and U8797 (N_8797,N_7098,N_7794);
nand U8798 (N_8798,N_7931,N_7124);
nand U8799 (N_8799,N_7778,N_7228);
or U8800 (N_8800,N_7260,N_7102);
nand U8801 (N_8801,N_7180,N_7349);
or U8802 (N_8802,N_7753,N_7248);
nand U8803 (N_8803,N_7814,N_7590);
nor U8804 (N_8804,N_7638,N_7202);
xnor U8805 (N_8805,N_7265,N_7650);
nand U8806 (N_8806,N_7605,N_7430);
or U8807 (N_8807,N_7311,N_7268);
xnor U8808 (N_8808,N_7062,N_7962);
nand U8809 (N_8809,N_7784,N_7271);
or U8810 (N_8810,N_7381,N_7881);
or U8811 (N_8811,N_7439,N_7224);
xor U8812 (N_8812,N_7754,N_7272);
and U8813 (N_8813,N_7569,N_7304);
xor U8814 (N_8814,N_7811,N_7250);
and U8815 (N_8815,N_7186,N_7552);
nor U8816 (N_8816,N_7024,N_7804);
xnor U8817 (N_8817,N_7291,N_7899);
or U8818 (N_8818,N_7961,N_7064);
or U8819 (N_8819,N_7462,N_7600);
xor U8820 (N_8820,N_7032,N_7041);
or U8821 (N_8821,N_7763,N_7678);
or U8822 (N_8822,N_7016,N_7986);
nor U8823 (N_8823,N_7150,N_7328);
and U8824 (N_8824,N_7133,N_7874);
and U8825 (N_8825,N_7641,N_7414);
xor U8826 (N_8826,N_7917,N_7475);
xnor U8827 (N_8827,N_7237,N_7500);
nor U8828 (N_8828,N_7245,N_7898);
nand U8829 (N_8829,N_7080,N_7365);
or U8830 (N_8830,N_7887,N_7984);
xnor U8831 (N_8831,N_7228,N_7643);
nor U8832 (N_8832,N_7342,N_7735);
and U8833 (N_8833,N_7497,N_7644);
xnor U8834 (N_8834,N_7053,N_7762);
or U8835 (N_8835,N_7699,N_7933);
and U8836 (N_8836,N_7067,N_7230);
and U8837 (N_8837,N_7544,N_7935);
and U8838 (N_8838,N_7360,N_7148);
xor U8839 (N_8839,N_7672,N_7462);
nand U8840 (N_8840,N_7025,N_7132);
nor U8841 (N_8841,N_7983,N_7769);
nor U8842 (N_8842,N_7118,N_7849);
and U8843 (N_8843,N_7247,N_7242);
or U8844 (N_8844,N_7600,N_7022);
nand U8845 (N_8845,N_7680,N_7531);
or U8846 (N_8846,N_7123,N_7082);
nand U8847 (N_8847,N_7346,N_7389);
or U8848 (N_8848,N_7943,N_7852);
or U8849 (N_8849,N_7959,N_7300);
xor U8850 (N_8850,N_7851,N_7864);
xnor U8851 (N_8851,N_7069,N_7151);
or U8852 (N_8852,N_7993,N_7517);
nor U8853 (N_8853,N_7609,N_7512);
xnor U8854 (N_8854,N_7632,N_7775);
and U8855 (N_8855,N_7077,N_7656);
and U8856 (N_8856,N_7360,N_7714);
and U8857 (N_8857,N_7204,N_7119);
xor U8858 (N_8858,N_7400,N_7217);
and U8859 (N_8859,N_7180,N_7795);
nor U8860 (N_8860,N_7225,N_7257);
or U8861 (N_8861,N_7970,N_7943);
and U8862 (N_8862,N_7737,N_7688);
nand U8863 (N_8863,N_7656,N_7456);
and U8864 (N_8864,N_7892,N_7591);
and U8865 (N_8865,N_7959,N_7480);
and U8866 (N_8866,N_7048,N_7916);
and U8867 (N_8867,N_7574,N_7415);
and U8868 (N_8868,N_7878,N_7218);
xor U8869 (N_8869,N_7796,N_7018);
and U8870 (N_8870,N_7122,N_7086);
nor U8871 (N_8871,N_7155,N_7090);
nand U8872 (N_8872,N_7409,N_7619);
nand U8873 (N_8873,N_7793,N_7167);
and U8874 (N_8874,N_7552,N_7489);
or U8875 (N_8875,N_7428,N_7432);
xor U8876 (N_8876,N_7611,N_7987);
nor U8877 (N_8877,N_7573,N_7838);
and U8878 (N_8878,N_7247,N_7237);
nand U8879 (N_8879,N_7155,N_7670);
xor U8880 (N_8880,N_7903,N_7151);
or U8881 (N_8881,N_7389,N_7902);
nor U8882 (N_8882,N_7545,N_7408);
nor U8883 (N_8883,N_7299,N_7446);
xor U8884 (N_8884,N_7218,N_7385);
nor U8885 (N_8885,N_7805,N_7769);
or U8886 (N_8886,N_7454,N_7844);
xnor U8887 (N_8887,N_7889,N_7364);
nor U8888 (N_8888,N_7649,N_7421);
xnor U8889 (N_8889,N_7476,N_7935);
xnor U8890 (N_8890,N_7498,N_7913);
and U8891 (N_8891,N_7177,N_7015);
nor U8892 (N_8892,N_7605,N_7370);
and U8893 (N_8893,N_7584,N_7673);
and U8894 (N_8894,N_7523,N_7997);
or U8895 (N_8895,N_7844,N_7071);
nor U8896 (N_8896,N_7269,N_7496);
and U8897 (N_8897,N_7647,N_7890);
or U8898 (N_8898,N_7665,N_7357);
nand U8899 (N_8899,N_7689,N_7225);
nand U8900 (N_8900,N_7919,N_7224);
and U8901 (N_8901,N_7067,N_7142);
xor U8902 (N_8902,N_7102,N_7725);
xnor U8903 (N_8903,N_7194,N_7630);
xor U8904 (N_8904,N_7413,N_7298);
and U8905 (N_8905,N_7824,N_7098);
nor U8906 (N_8906,N_7336,N_7044);
nand U8907 (N_8907,N_7095,N_7807);
or U8908 (N_8908,N_7942,N_7863);
nand U8909 (N_8909,N_7481,N_7380);
nand U8910 (N_8910,N_7666,N_7930);
or U8911 (N_8911,N_7971,N_7195);
nand U8912 (N_8912,N_7506,N_7122);
or U8913 (N_8913,N_7936,N_7815);
nor U8914 (N_8914,N_7513,N_7815);
and U8915 (N_8915,N_7799,N_7875);
or U8916 (N_8916,N_7586,N_7625);
or U8917 (N_8917,N_7497,N_7703);
and U8918 (N_8918,N_7104,N_7943);
nor U8919 (N_8919,N_7215,N_7561);
nor U8920 (N_8920,N_7539,N_7625);
or U8921 (N_8921,N_7906,N_7117);
or U8922 (N_8922,N_7301,N_7710);
nor U8923 (N_8923,N_7857,N_7771);
nor U8924 (N_8924,N_7127,N_7261);
xor U8925 (N_8925,N_7526,N_7298);
nor U8926 (N_8926,N_7680,N_7915);
xor U8927 (N_8927,N_7909,N_7079);
xor U8928 (N_8928,N_7989,N_7039);
nor U8929 (N_8929,N_7157,N_7029);
or U8930 (N_8930,N_7279,N_7691);
or U8931 (N_8931,N_7171,N_7255);
nor U8932 (N_8932,N_7053,N_7711);
nor U8933 (N_8933,N_7504,N_7756);
nand U8934 (N_8934,N_7529,N_7503);
nor U8935 (N_8935,N_7217,N_7667);
nand U8936 (N_8936,N_7885,N_7571);
or U8937 (N_8937,N_7753,N_7263);
nor U8938 (N_8938,N_7157,N_7627);
nand U8939 (N_8939,N_7198,N_7789);
xnor U8940 (N_8940,N_7250,N_7388);
nand U8941 (N_8941,N_7896,N_7755);
xor U8942 (N_8942,N_7523,N_7218);
xor U8943 (N_8943,N_7001,N_7896);
nor U8944 (N_8944,N_7216,N_7055);
or U8945 (N_8945,N_7981,N_7276);
or U8946 (N_8946,N_7446,N_7102);
nor U8947 (N_8947,N_7108,N_7885);
nor U8948 (N_8948,N_7069,N_7686);
and U8949 (N_8949,N_7841,N_7731);
and U8950 (N_8950,N_7060,N_7971);
nand U8951 (N_8951,N_7458,N_7235);
and U8952 (N_8952,N_7122,N_7859);
nor U8953 (N_8953,N_7680,N_7104);
nor U8954 (N_8954,N_7631,N_7809);
and U8955 (N_8955,N_7647,N_7096);
or U8956 (N_8956,N_7251,N_7764);
nand U8957 (N_8957,N_7065,N_7463);
nand U8958 (N_8958,N_7946,N_7989);
and U8959 (N_8959,N_7739,N_7406);
xnor U8960 (N_8960,N_7815,N_7153);
xor U8961 (N_8961,N_7382,N_7587);
and U8962 (N_8962,N_7174,N_7034);
nand U8963 (N_8963,N_7186,N_7347);
nor U8964 (N_8964,N_7848,N_7281);
nor U8965 (N_8965,N_7527,N_7925);
xor U8966 (N_8966,N_7158,N_7463);
and U8967 (N_8967,N_7102,N_7379);
nor U8968 (N_8968,N_7069,N_7941);
or U8969 (N_8969,N_7811,N_7134);
xor U8970 (N_8970,N_7609,N_7649);
and U8971 (N_8971,N_7191,N_7145);
or U8972 (N_8972,N_7656,N_7603);
nand U8973 (N_8973,N_7692,N_7624);
or U8974 (N_8974,N_7780,N_7989);
xnor U8975 (N_8975,N_7076,N_7030);
nand U8976 (N_8976,N_7494,N_7899);
and U8977 (N_8977,N_7648,N_7498);
or U8978 (N_8978,N_7756,N_7061);
xnor U8979 (N_8979,N_7186,N_7918);
nor U8980 (N_8980,N_7122,N_7851);
nand U8981 (N_8981,N_7527,N_7930);
xor U8982 (N_8982,N_7259,N_7719);
xor U8983 (N_8983,N_7659,N_7444);
and U8984 (N_8984,N_7753,N_7566);
or U8985 (N_8985,N_7336,N_7153);
and U8986 (N_8986,N_7602,N_7254);
nand U8987 (N_8987,N_7006,N_7563);
or U8988 (N_8988,N_7924,N_7036);
xor U8989 (N_8989,N_7778,N_7845);
nor U8990 (N_8990,N_7879,N_7295);
nand U8991 (N_8991,N_7497,N_7884);
or U8992 (N_8992,N_7673,N_7737);
or U8993 (N_8993,N_7824,N_7395);
or U8994 (N_8994,N_7675,N_7974);
nor U8995 (N_8995,N_7107,N_7898);
xnor U8996 (N_8996,N_7691,N_7854);
nor U8997 (N_8997,N_7533,N_7777);
nand U8998 (N_8998,N_7014,N_7744);
xor U8999 (N_8999,N_7804,N_7233);
and U9000 (N_9000,N_8237,N_8907);
and U9001 (N_9001,N_8932,N_8376);
or U9002 (N_9002,N_8930,N_8817);
and U9003 (N_9003,N_8512,N_8878);
and U9004 (N_9004,N_8795,N_8748);
nor U9005 (N_9005,N_8150,N_8152);
and U9006 (N_9006,N_8393,N_8377);
nand U9007 (N_9007,N_8896,N_8790);
or U9008 (N_9008,N_8202,N_8109);
nand U9009 (N_9009,N_8985,N_8833);
xor U9010 (N_9010,N_8205,N_8765);
xor U9011 (N_9011,N_8055,N_8664);
nand U9012 (N_9012,N_8596,N_8616);
and U9013 (N_9013,N_8414,N_8669);
or U9014 (N_9014,N_8742,N_8798);
and U9015 (N_9015,N_8654,N_8372);
or U9016 (N_9016,N_8358,N_8027);
or U9017 (N_9017,N_8291,N_8723);
nand U9018 (N_9018,N_8854,N_8049);
xor U9019 (N_9019,N_8333,N_8701);
and U9020 (N_9020,N_8266,N_8371);
nand U9021 (N_9021,N_8535,N_8452);
nand U9022 (N_9022,N_8784,N_8581);
nor U9023 (N_9023,N_8649,N_8382);
and U9024 (N_9024,N_8147,N_8425);
nor U9025 (N_9025,N_8953,N_8689);
nand U9026 (N_9026,N_8543,N_8011);
or U9027 (N_9027,N_8990,N_8951);
nand U9028 (N_9028,N_8464,N_8920);
nor U9029 (N_9029,N_8656,N_8045);
or U9030 (N_9030,N_8419,N_8006);
nand U9031 (N_9031,N_8568,N_8588);
or U9032 (N_9032,N_8621,N_8565);
xor U9033 (N_9033,N_8753,N_8307);
nor U9034 (N_9034,N_8971,N_8732);
nor U9035 (N_9035,N_8453,N_8767);
and U9036 (N_9036,N_8935,N_8127);
nor U9037 (N_9037,N_8238,N_8904);
xnor U9038 (N_9038,N_8966,N_8631);
and U9039 (N_9039,N_8403,N_8956);
nand U9040 (N_9040,N_8346,N_8420);
or U9041 (N_9041,N_8200,N_8877);
or U9042 (N_9042,N_8937,N_8069);
nor U9043 (N_9043,N_8478,N_8788);
xnor U9044 (N_9044,N_8611,N_8820);
xnor U9045 (N_9045,N_8711,N_8763);
nor U9046 (N_9046,N_8181,N_8949);
nor U9047 (N_9047,N_8265,N_8516);
or U9048 (N_9048,N_8340,N_8702);
xnor U9049 (N_9049,N_8140,N_8410);
nand U9050 (N_9050,N_8633,N_8774);
xnor U9051 (N_9051,N_8899,N_8670);
or U9052 (N_9052,N_8526,N_8350);
xnor U9053 (N_9053,N_8569,N_8038);
and U9054 (N_9054,N_8772,N_8004);
nand U9055 (N_9055,N_8864,N_8706);
and U9056 (N_9056,N_8725,N_8620);
and U9057 (N_9057,N_8406,N_8791);
nand U9058 (N_9058,N_8034,N_8575);
and U9059 (N_9059,N_8020,N_8874);
and U9060 (N_9060,N_8892,N_8037);
and U9061 (N_9061,N_8434,N_8397);
xnor U9062 (N_9062,N_8713,N_8299);
nand U9063 (N_9063,N_8728,N_8680);
or U9064 (N_9064,N_8842,N_8277);
nand U9065 (N_9065,N_8095,N_8586);
and U9066 (N_9066,N_8607,N_8457);
or U9067 (N_9067,N_8635,N_8413);
xor U9068 (N_9068,N_8313,N_8000);
xnor U9069 (N_9069,N_8477,N_8334);
nor U9070 (N_9070,N_8462,N_8982);
and U9071 (N_9071,N_8963,N_8193);
xor U9072 (N_9072,N_8173,N_8059);
and U9073 (N_9073,N_8169,N_8808);
or U9074 (N_9074,N_8960,N_8282);
nand U9075 (N_9075,N_8077,N_8245);
xor U9076 (N_9076,N_8293,N_8514);
nor U9077 (N_9077,N_8928,N_8001);
and U9078 (N_9078,N_8668,N_8244);
xor U9079 (N_9079,N_8578,N_8128);
and U9080 (N_9080,N_8523,N_8459);
and U9081 (N_9081,N_8893,N_8741);
or U9082 (N_9082,N_8972,N_8185);
xnor U9083 (N_9083,N_8112,N_8294);
and U9084 (N_9084,N_8344,N_8673);
nand U9085 (N_9085,N_8021,N_8008);
nand U9086 (N_9086,N_8658,N_8866);
nand U9087 (N_9087,N_8468,N_8463);
and U9088 (N_9088,N_8832,N_8871);
and U9089 (N_9089,N_8143,N_8720);
nand U9090 (N_9090,N_8383,N_8872);
nand U9091 (N_9091,N_8409,N_8641);
nand U9092 (N_9092,N_8879,N_8912);
and U9093 (N_9093,N_8751,N_8280);
nand U9094 (N_9094,N_8639,N_8524);
nor U9095 (N_9095,N_8121,N_8133);
xor U9096 (N_9096,N_8782,N_8646);
xor U9097 (N_9097,N_8992,N_8220);
or U9098 (N_9098,N_8480,N_8848);
xor U9099 (N_9099,N_8215,N_8922);
nand U9100 (N_9100,N_8430,N_8973);
or U9101 (N_9101,N_8540,N_8438);
or U9102 (N_9102,N_8863,N_8253);
or U9103 (N_9103,N_8709,N_8317);
and U9104 (N_9104,N_8472,N_8969);
nand U9105 (N_9105,N_8597,N_8362);
xnor U9106 (N_9106,N_8944,N_8002);
nor U9107 (N_9107,N_8690,N_8623);
xnor U9108 (N_9108,N_8891,N_8529);
or U9109 (N_9109,N_8506,N_8302);
or U9110 (N_9110,N_8638,N_8249);
or U9111 (N_9111,N_8675,N_8336);
nand U9112 (N_9112,N_8954,N_8634);
xnor U9113 (N_9113,N_8769,N_8063);
or U9114 (N_9114,N_8941,N_8589);
and U9115 (N_9115,N_8933,N_8677);
and U9116 (N_9116,N_8549,N_8235);
or U9117 (N_9117,N_8361,N_8338);
or U9118 (N_9118,N_8227,N_8727);
and U9119 (N_9119,N_8895,N_8965);
xnor U9120 (N_9120,N_8945,N_8564);
and U9121 (N_9121,N_8141,N_8913);
nand U9122 (N_9122,N_8595,N_8190);
xor U9123 (N_9123,N_8867,N_8053);
or U9124 (N_9124,N_8601,N_8332);
nand U9125 (N_9125,N_8983,N_8297);
or U9126 (N_9126,N_8417,N_8803);
xnor U9127 (N_9127,N_8476,N_8672);
nand U9128 (N_9128,N_8373,N_8129);
nand U9129 (N_9129,N_8154,N_8756);
nand U9130 (N_9130,N_8217,N_8640);
and U9131 (N_9131,N_8231,N_8988);
xor U9132 (N_9132,N_8805,N_8062);
or U9133 (N_9133,N_8212,N_8281);
nor U9134 (N_9134,N_8651,N_8278);
nand U9135 (N_9135,N_8174,N_8760);
nand U9136 (N_9136,N_8582,N_8726);
nor U9137 (N_9137,N_8657,N_8347);
or U9138 (N_9138,N_8036,N_8903);
or U9139 (N_9139,N_8806,N_8255);
nand U9140 (N_9140,N_8987,N_8525);
or U9141 (N_9141,N_8473,N_8441);
xnor U9142 (N_9142,N_8773,N_8840);
xor U9143 (N_9143,N_8498,N_8243);
and U9144 (N_9144,N_8745,N_8610);
and U9145 (N_9145,N_8576,N_8351);
or U9146 (N_9146,N_8345,N_8697);
xnor U9147 (N_9147,N_8475,N_8593);
nor U9148 (N_9148,N_8974,N_8314);
nor U9149 (N_9149,N_8600,N_8500);
and U9150 (N_9150,N_8734,N_8545);
and U9151 (N_9151,N_8003,N_8510);
and U9152 (N_9152,N_8836,N_8606);
or U9153 (N_9153,N_8260,N_8708);
xor U9154 (N_9154,N_8167,N_8555);
and U9155 (N_9155,N_8934,N_8747);
or U9156 (N_9156,N_8192,N_8938);
nand U9157 (N_9157,N_8749,N_8067);
xor U9158 (N_9158,N_8554,N_8353);
and U9159 (N_9159,N_8149,N_8348);
nor U9160 (N_9160,N_8835,N_8089);
nand U9161 (N_9161,N_8213,N_8915);
and U9162 (N_9162,N_8859,N_8159);
nor U9163 (N_9163,N_8797,N_8444);
or U9164 (N_9164,N_8400,N_8698);
and U9165 (N_9165,N_8496,N_8290);
xnor U9166 (N_9166,N_8630,N_8447);
and U9167 (N_9167,N_8683,N_8225);
xnor U9168 (N_9168,N_8979,N_8070);
xor U9169 (N_9169,N_8997,N_8379);
or U9170 (N_9170,N_8685,N_8076);
and U9171 (N_9171,N_8572,N_8086);
xnor U9172 (N_9172,N_8590,N_8275);
nand U9173 (N_9173,N_8039,N_8718);
nor U9174 (N_9174,N_8531,N_8078);
and U9175 (N_9175,N_8226,N_8684);
nand U9176 (N_9176,N_8497,N_8515);
and U9177 (N_9177,N_8556,N_8776);
or U9178 (N_9178,N_8232,N_8839);
or U9179 (N_9179,N_8705,N_8902);
nor U9180 (N_9180,N_8541,N_8770);
nand U9181 (N_9181,N_8563,N_8768);
nand U9182 (N_9182,N_8183,N_8870);
xor U9183 (N_9183,N_8598,N_8084);
or U9184 (N_9184,N_8522,N_8882);
or U9185 (N_9185,N_8198,N_8612);
nand U9186 (N_9186,N_8827,N_8838);
nand U9187 (N_9187,N_8865,N_8534);
or U9188 (N_9188,N_8771,N_8164);
nand U9189 (N_9189,N_8752,N_8308);
nor U9190 (N_9190,N_8108,N_8355);
or U9191 (N_9191,N_8398,N_8977);
xnor U9192 (N_9192,N_8861,N_8644);
nor U9193 (N_9193,N_8936,N_8663);
nor U9194 (N_9194,N_8330,N_8196);
nor U9195 (N_9195,N_8072,N_8566);
nor U9196 (N_9196,N_8738,N_8144);
nor U9197 (N_9197,N_8214,N_8482);
and U9198 (N_9198,N_8274,N_8599);
or U9199 (N_9199,N_8804,N_8486);
and U9200 (N_9200,N_8811,N_8024);
nor U9201 (N_9201,N_8028,N_8399);
nor U9202 (N_9202,N_8097,N_8585);
or U9203 (N_9203,N_8052,N_8883);
nor U9204 (N_9204,N_8356,N_8079);
nand U9205 (N_9205,N_8740,N_8026);
nand U9206 (N_9206,N_8385,N_8743);
nor U9207 (N_9207,N_8671,N_8010);
or U9208 (N_9208,N_8388,N_8315);
nor U9209 (N_9209,N_8189,N_8815);
or U9210 (N_9210,N_8652,N_8423);
or U9211 (N_9211,N_8170,N_8551);
or U9212 (N_9212,N_8900,N_8256);
or U9213 (N_9213,N_8730,N_8451);
or U9214 (N_9214,N_8123,N_8239);
nand U9215 (N_9215,N_8918,N_8157);
and U9216 (N_9216,N_8416,N_8488);
or U9217 (N_9217,N_8733,N_8208);
or U9218 (N_9218,N_8528,N_8374);
nand U9219 (N_9219,N_8699,N_8342);
and U9220 (N_9220,N_8094,N_8629);
or U9221 (N_9221,N_8536,N_8520);
nor U9222 (N_9222,N_8947,N_8602);
and U9223 (N_9223,N_8659,N_8851);
xnor U9224 (N_9224,N_8396,N_8868);
nor U9225 (N_9225,N_8923,N_8722);
nand U9226 (N_9226,N_8824,N_8359);
xor U9227 (N_9227,N_8502,N_8958);
nor U9228 (N_9228,N_8492,N_8354);
or U9229 (N_9229,N_8199,N_8424);
nor U9230 (N_9230,N_8645,N_8461);
or U9231 (N_9231,N_8318,N_8905);
nor U9232 (N_9232,N_8357,N_8092);
xor U9233 (N_9233,N_8432,N_8624);
xor U9234 (N_9234,N_8775,N_8009);
and U9235 (N_9235,N_8386,N_8096);
nand U9236 (N_9236,N_8494,N_8889);
and U9237 (N_9237,N_8996,N_8898);
nand U9238 (N_9238,N_8537,N_8609);
nor U9239 (N_9239,N_8106,N_8073);
nor U9240 (N_9240,N_8310,N_8044);
nand U9241 (N_9241,N_8201,N_8888);
nand U9242 (N_9242,N_8364,N_8248);
or U9243 (N_9243,N_8802,N_8801);
or U9244 (N_9244,N_8674,N_8178);
nor U9245 (N_9245,N_8687,N_8552);
or U9246 (N_9246,N_8682,N_8270);
or U9247 (N_9247,N_8378,N_8816);
or U9248 (N_9248,N_8766,N_8544);
nand U9249 (N_9249,N_8691,N_8875);
nor U9250 (N_9250,N_8681,N_8269);
or U9251 (N_9251,N_8679,N_8343);
xnor U9252 (N_9252,N_8583,N_8223);
or U9253 (N_9253,N_8104,N_8830);
and U9254 (N_9254,N_8485,N_8114);
or U9255 (N_9255,N_8507,N_8828);
or U9256 (N_9256,N_8577,N_8984);
nor U9257 (N_9257,N_8341,N_8363);
or U9258 (N_9258,N_8643,N_8787);
nor U9259 (N_9259,N_8254,N_8369);
nor U9260 (N_9260,N_8707,N_8739);
nand U9261 (N_9261,N_8825,N_8405);
nor U9262 (N_9262,N_8186,N_8309);
or U9263 (N_9263,N_8242,N_8271);
and U9264 (N_9264,N_8981,N_8050);
nor U9265 (N_9265,N_8925,N_8258);
nand U9266 (N_9266,N_8047,N_8931);
nor U9267 (N_9267,N_8695,N_8735);
or U9268 (N_9268,N_8130,N_8029);
or U9269 (N_9269,N_8926,N_8224);
nand U9270 (N_9270,N_8917,N_8873);
nand U9271 (N_9271,N_8712,N_8176);
and U9272 (N_9272,N_8312,N_8942);
nand U9273 (N_9273,N_8210,N_8043);
and U9274 (N_9274,N_8381,N_8197);
xnor U9275 (N_9275,N_8251,N_8818);
xnor U9276 (N_9276,N_8573,N_8483);
xnor U9277 (N_9277,N_8560,N_8908);
nand U9278 (N_9278,N_8608,N_8513);
xnor U9279 (N_9279,N_8435,N_8618);
or U9280 (N_9280,N_8207,N_8203);
or U9281 (N_9281,N_8324,N_8910);
nand U9282 (N_9282,N_8636,N_8428);
or U9283 (N_9283,N_8012,N_8138);
xnor U9284 (N_9284,N_8440,N_8126);
nand U9285 (N_9285,N_8276,N_8113);
or U9286 (N_9286,N_8155,N_8445);
nor U9287 (N_9287,N_8261,N_8304);
nor U9288 (N_9288,N_8780,N_8470);
or U9289 (N_9289,N_8057,N_8110);
and U9290 (N_9290,N_8853,N_8655);
nand U9291 (N_9291,N_8395,N_8375);
nor U9292 (N_9292,N_8137,N_8604);
nor U9293 (N_9293,N_8474,N_8319);
and U9294 (N_9294,N_8532,N_8994);
nand U9295 (N_9295,N_8490,N_8180);
xor U9296 (N_9296,N_8642,N_8959);
or U9297 (N_9297,N_8267,N_8329);
or U9298 (N_9298,N_8234,N_8964);
xor U9299 (N_9299,N_8731,N_8219);
or U9300 (N_9300,N_8431,N_8132);
and U9301 (N_9301,N_8099,N_8617);
and U9302 (N_9302,N_8857,N_8999);
nand U9303 (N_9303,N_8919,N_8813);
xor U9304 (N_9304,N_8986,N_8032);
xnor U9305 (N_9305,N_8054,N_8301);
nor U9306 (N_9306,N_8163,N_8153);
xnor U9307 (N_9307,N_8561,N_8778);
or U9308 (N_9308,N_8511,N_8172);
nand U9309 (N_9309,N_8710,N_8025);
xnor U9310 (N_9310,N_8911,N_8625);
nand U9311 (N_9311,N_8087,N_8439);
and U9312 (N_9312,N_8829,N_8066);
and U9313 (N_9313,N_8422,N_8794);
nor U9314 (N_9314,N_8111,N_8040);
or U9315 (N_9315,N_8619,N_8562);
or U9316 (N_9316,N_8862,N_8887);
nor U9317 (N_9317,N_8367,N_8796);
or U9318 (N_9318,N_8626,N_8961);
or U9319 (N_9319,N_8100,N_8469);
and U9320 (N_9320,N_8158,N_8807);
nand U9321 (N_9321,N_8437,N_8637);
nor U9322 (N_9322,N_8591,N_8449);
nor U9323 (N_9323,N_8465,N_8320);
nor U9324 (N_9324,N_8648,N_8989);
nand U9325 (N_9325,N_8171,N_8136);
and U9326 (N_9326,N_8594,N_8548);
nor U9327 (N_9327,N_8810,N_8856);
xor U9328 (N_9328,N_8897,N_8407);
and U9329 (N_9329,N_8448,N_8390);
xnor U9330 (N_9330,N_8759,N_8809);
or U9331 (N_9331,N_8075,N_8976);
nor U9332 (N_9332,N_8321,N_8156);
or U9333 (N_9333,N_8325,N_8031);
or U9334 (N_9334,N_8881,N_8443);
and U9335 (N_9335,N_8081,N_8404);
and U9336 (N_9336,N_8826,N_8151);
and U9337 (N_9337,N_8117,N_8454);
and U9338 (N_9338,N_8068,N_8692);
or U9339 (N_9339,N_8940,N_8392);
or U9340 (N_9340,N_8880,N_8284);
and U9341 (N_9341,N_8091,N_8145);
nand U9342 (N_9342,N_8714,N_8134);
nor U9343 (N_9343,N_8924,N_8850);
and U9344 (N_9344,N_8098,N_8122);
nand U9345 (N_9345,N_8283,N_8819);
or U9346 (N_9346,N_8519,N_8305);
or U9347 (N_9347,N_8704,N_8559);
and U9348 (N_9348,N_8613,N_8495);
or U9349 (N_9349,N_8509,N_8391);
nand U9350 (N_9350,N_8546,N_8744);
or U9351 (N_9351,N_8846,N_8105);
or U9352 (N_9352,N_8030,N_8394);
nor U9353 (N_9353,N_8048,N_8950);
nand U9354 (N_9354,N_8119,N_8493);
and U9355 (N_9355,N_8182,N_8131);
and U9356 (N_9356,N_8946,N_8019);
nand U9357 (N_9357,N_8799,N_8187);
nor U9358 (N_9358,N_8884,N_8216);
nand U9359 (N_9359,N_8508,N_8368);
and U9360 (N_9360,N_8855,N_8421);
nor U9361 (N_9361,N_8647,N_8886);
nor U9362 (N_9362,N_8335,N_8328);
xnor U9363 (N_9363,N_8327,N_8539);
or U9364 (N_9364,N_8995,N_8458);
xor U9365 (N_9365,N_8429,N_8750);
nor U9366 (N_9366,N_8139,N_8841);
nand U9367 (N_9367,N_8665,N_8401);
nor U9368 (N_9368,N_8148,N_8300);
and U9369 (N_9369,N_8737,N_8821);
xor U9370 (N_9370,N_8135,N_8614);
nor U9371 (N_9371,N_8688,N_8980);
and U9372 (N_9372,N_8650,N_8781);
xor U9373 (N_9373,N_8957,N_8088);
or U9374 (N_9374,N_8852,N_8627);
nor U9375 (N_9375,N_8298,N_8365);
xnor U9376 (N_9376,N_8653,N_8592);
xnor U9377 (N_9377,N_8177,N_8939);
and U9378 (N_9378,N_8222,N_8455);
nor U9379 (N_9379,N_8311,N_8762);
nand U9380 (N_9380,N_8168,N_8316);
or U9381 (N_9381,N_8264,N_8754);
xor U9382 (N_9382,N_8632,N_8696);
or U9383 (N_9383,N_8736,N_8360);
nor U9384 (N_9384,N_8521,N_8194);
xnor U9385 (N_9385,N_8858,N_8296);
nand U9386 (N_9386,N_8792,N_8703);
or U9387 (N_9387,N_8948,N_8719);
or U9388 (N_9388,N_8501,N_8518);
xnor U9389 (N_9389,N_8427,N_8761);
and U9390 (N_9390,N_8746,N_8757);
nor U9391 (N_9391,N_8058,N_8489);
nor U9392 (N_9392,N_8331,N_8530);
and U9393 (N_9393,N_8694,N_8230);
nand U9394 (N_9394,N_8481,N_8471);
or U9395 (N_9395,N_8579,N_8894);
and U9396 (N_9396,N_8570,N_8380);
or U9397 (N_9397,N_8083,N_8322);
and U9398 (N_9398,N_8188,N_8250);
xnor U9399 (N_9399,N_8571,N_8060);
and U9400 (N_9400,N_8615,N_8056);
or U9401 (N_9401,N_8755,N_8547);
or U9402 (N_9402,N_8777,N_8843);
nand U9403 (N_9403,N_8229,N_8209);
xor U9404 (N_9404,N_8349,N_8370);
xor U9405 (N_9405,N_8890,N_8337);
and U9406 (N_9406,N_8834,N_8259);
nor U9407 (N_9407,N_8538,N_8085);
nand U9408 (N_9408,N_8456,N_8241);
xor U9409 (N_9409,N_8952,N_8678);
and U9410 (N_9410,N_8204,N_8061);
or U9411 (N_9411,N_8285,N_8339);
nand U9412 (N_9412,N_8013,N_8191);
nor U9413 (N_9413,N_8542,N_8268);
nor U9414 (N_9414,N_8246,N_8786);
nand U9415 (N_9415,N_8758,N_8721);
or U9416 (N_9416,N_8273,N_8228);
and U9417 (N_9417,N_8715,N_8517);
or U9418 (N_9418,N_8142,N_8093);
nand U9419 (N_9419,N_8567,N_8785);
and U9420 (N_9420,N_8914,N_8503);
and U9421 (N_9421,N_8844,N_8366);
nor U9422 (N_9422,N_8667,N_8046);
xor U9423 (N_9423,N_8622,N_8323);
or U9424 (N_9424,N_8279,N_8389);
nand U9425 (N_9425,N_8460,N_8411);
nand U9426 (N_9426,N_8415,N_8504);
xnor U9427 (N_9427,N_8433,N_8533);
and U9428 (N_9428,N_8975,N_8005);
nor U9429 (N_9429,N_8837,N_8115);
xor U9430 (N_9430,N_8849,N_8716);
nand U9431 (N_9431,N_8467,N_8218);
nand U9432 (N_9432,N_8287,N_8233);
and U9433 (N_9433,N_8550,N_8175);
xor U9434 (N_9434,N_8018,N_8402);
nor U9435 (N_9435,N_8384,N_8074);
and U9436 (N_9436,N_8724,N_8876);
or U9437 (N_9437,N_8033,N_8901);
or U9438 (N_9438,N_8927,N_8628);
or U9439 (N_9439,N_8118,N_8065);
or U9440 (N_9440,N_8412,N_8184);
nand U9441 (N_9441,N_8295,N_8071);
nor U9442 (N_9442,N_8793,N_8101);
or U9443 (N_9443,N_8426,N_8800);
nand U9444 (N_9444,N_8102,N_8929);
nand U9445 (N_9445,N_8660,N_8450);
or U9446 (N_9446,N_8845,N_8120);
or U9447 (N_9447,N_8446,N_8847);
and U9448 (N_9448,N_8779,N_8955);
or U9449 (N_9449,N_8584,N_8831);
and U9450 (N_9450,N_8812,N_8023);
and U9451 (N_9451,N_8236,N_8035);
or U9452 (N_9452,N_8968,N_8292);
or U9453 (N_9453,N_8967,N_8090);
xor U9454 (N_9454,N_8998,N_8160);
xnor U9455 (N_9455,N_8007,N_8306);
xor U9456 (N_9456,N_8557,N_8042);
or U9457 (N_9457,N_8991,N_8211);
xor U9458 (N_9458,N_8661,N_8558);
nor U9459 (N_9459,N_8921,N_8764);
nand U9460 (N_9460,N_8051,N_8499);
nand U9461 (N_9461,N_8491,N_8303);
and U9462 (N_9462,N_8286,N_8860);
or U9463 (N_9463,N_8165,N_8943);
nand U9464 (N_9464,N_8418,N_8822);
or U9465 (N_9465,N_8387,N_8166);
or U9466 (N_9466,N_8676,N_8603);
xnor U9467 (N_9467,N_8553,N_8814);
or U9468 (N_9468,N_8823,N_8700);
and U9469 (N_9469,N_8662,N_8729);
nor U9470 (N_9470,N_8783,N_8124);
or U9471 (N_9471,N_8247,N_8970);
and U9472 (N_9472,N_8080,N_8962);
xor U9473 (N_9473,N_8527,N_8666);
nor U9474 (N_9474,N_8408,N_8116);
xor U9475 (N_9475,N_8580,N_8587);
or U9476 (N_9476,N_8993,N_8082);
nor U9477 (N_9477,N_8436,N_8146);
or U9478 (N_9478,N_8916,N_8103);
nor U9479 (N_9479,N_8257,N_8466);
nand U9480 (N_9480,N_8125,N_8240);
nand U9481 (N_9481,N_8064,N_8574);
or U9482 (N_9482,N_8484,N_8022);
nor U9483 (N_9483,N_8505,N_8717);
nor U9484 (N_9484,N_8909,N_8017);
and U9485 (N_9485,N_8789,N_8016);
or U9486 (N_9486,N_8487,N_8442);
nand U9487 (N_9487,N_8263,N_8262);
nand U9488 (N_9488,N_8179,N_8288);
or U9489 (N_9489,N_8221,N_8693);
or U9490 (N_9490,N_8978,N_8885);
xor U9491 (N_9491,N_8686,N_8869);
or U9492 (N_9492,N_8195,N_8161);
xnor U9493 (N_9493,N_8289,N_8272);
xnor U9494 (N_9494,N_8352,N_8014);
nor U9495 (N_9495,N_8906,N_8605);
and U9496 (N_9496,N_8107,N_8041);
nand U9497 (N_9497,N_8326,N_8162);
or U9498 (N_9498,N_8479,N_8206);
and U9499 (N_9499,N_8252,N_8015);
xor U9500 (N_9500,N_8072,N_8206);
or U9501 (N_9501,N_8807,N_8957);
or U9502 (N_9502,N_8774,N_8266);
xnor U9503 (N_9503,N_8671,N_8133);
nand U9504 (N_9504,N_8623,N_8833);
xnor U9505 (N_9505,N_8944,N_8796);
or U9506 (N_9506,N_8546,N_8152);
nor U9507 (N_9507,N_8905,N_8658);
nand U9508 (N_9508,N_8335,N_8283);
xor U9509 (N_9509,N_8519,N_8905);
nand U9510 (N_9510,N_8919,N_8475);
nand U9511 (N_9511,N_8275,N_8206);
or U9512 (N_9512,N_8311,N_8791);
and U9513 (N_9513,N_8822,N_8794);
xor U9514 (N_9514,N_8004,N_8372);
nor U9515 (N_9515,N_8730,N_8763);
xnor U9516 (N_9516,N_8248,N_8022);
nor U9517 (N_9517,N_8814,N_8436);
xor U9518 (N_9518,N_8607,N_8392);
nor U9519 (N_9519,N_8222,N_8823);
or U9520 (N_9520,N_8278,N_8100);
xnor U9521 (N_9521,N_8671,N_8223);
and U9522 (N_9522,N_8219,N_8562);
nor U9523 (N_9523,N_8184,N_8612);
xnor U9524 (N_9524,N_8560,N_8578);
nand U9525 (N_9525,N_8500,N_8194);
xor U9526 (N_9526,N_8628,N_8626);
nor U9527 (N_9527,N_8475,N_8479);
and U9528 (N_9528,N_8516,N_8550);
xor U9529 (N_9529,N_8214,N_8113);
nor U9530 (N_9530,N_8739,N_8828);
or U9531 (N_9531,N_8262,N_8189);
or U9532 (N_9532,N_8805,N_8787);
xnor U9533 (N_9533,N_8474,N_8012);
or U9534 (N_9534,N_8429,N_8293);
and U9535 (N_9535,N_8609,N_8807);
or U9536 (N_9536,N_8068,N_8684);
or U9537 (N_9537,N_8767,N_8555);
or U9538 (N_9538,N_8046,N_8226);
and U9539 (N_9539,N_8909,N_8560);
or U9540 (N_9540,N_8610,N_8410);
and U9541 (N_9541,N_8833,N_8926);
and U9542 (N_9542,N_8300,N_8854);
and U9543 (N_9543,N_8666,N_8434);
nor U9544 (N_9544,N_8926,N_8076);
or U9545 (N_9545,N_8413,N_8757);
and U9546 (N_9546,N_8787,N_8304);
xor U9547 (N_9547,N_8166,N_8706);
or U9548 (N_9548,N_8616,N_8131);
nand U9549 (N_9549,N_8580,N_8520);
nor U9550 (N_9550,N_8271,N_8266);
and U9551 (N_9551,N_8011,N_8793);
nand U9552 (N_9552,N_8816,N_8765);
nor U9553 (N_9553,N_8239,N_8002);
and U9554 (N_9554,N_8422,N_8524);
and U9555 (N_9555,N_8821,N_8429);
xnor U9556 (N_9556,N_8728,N_8156);
and U9557 (N_9557,N_8957,N_8856);
xor U9558 (N_9558,N_8232,N_8415);
nand U9559 (N_9559,N_8138,N_8019);
nor U9560 (N_9560,N_8405,N_8333);
or U9561 (N_9561,N_8319,N_8225);
and U9562 (N_9562,N_8088,N_8251);
nand U9563 (N_9563,N_8494,N_8555);
xor U9564 (N_9564,N_8425,N_8418);
nor U9565 (N_9565,N_8446,N_8743);
or U9566 (N_9566,N_8274,N_8264);
nor U9567 (N_9567,N_8597,N_8958);
nand U9568 (N_9568,N_8723,N_8627);
or U9569 (N_9569,N_8186,N_8378);
or U9570 (N_9570,N_8710,N_8640);
nor U9571 (N_9571,N_8598,N_8945);
and U9572 (N_9572,N_8725,N_8318);
and U9573 (N_9573,N_8733,N_8524);
nand U9574 (N_9574,N_8348,N_8104);
nor U9575 (N_9575,N_8120,N_8552);
or U9576 (N_9576,N_8049,N_8259);
nand U9577 (N_9577,N_8689,N_8091);
nand U9578 (N_9578,N_8648,N_8096);
nor U9579 (N_9579,N_8377,N_8428);
nor U9580 (N_9580,N_8084,N_8899);
and U9581 (N_9581,N_8124,N_8748);
nand U9582 (N_9582,N_8639,N_8049);
xor U9583 (N_9583,N_8163,N_8967);
nand U9584 (N_9584,N_8404,N_8079);
and U9585 (N_9585,N_8281,N_8814);
and U9586 (N_9586,N_8060,N_8891);
nor U9587 (N_9587,N_8403,N_8386);
or U9588 (N_9588,N_8063,N_8461);
xnor U9589 (N_9589,N_8927,N_8869);
xor U9590 (N_9590,N_8114,N_8058);
and U9591 (N_9591,N_8496,N_8519);
and U9592 (N_9592,N_8207,N_8806);
nor U9593 (N_9593,N_8549,N_8044);
and U9594 (N_9594,N_8010,N_8433);
nand U9595 (N_9595,N_8384,N_8269);
and U9596 (N_9596,N_8236,N_8031);
nor U9597 (N_9597,N_8955,N_8456);
xnor U9598 (N_9598,N_8939,N_8295);
and U9599 (N_9599,N_8487,N_8019);
nand U9600 (N_9600,N_8408,N_8181);
and U9601 (N_9601,N_8427,N_8277);
or U9602 (N_9602,N_8315,N_8178);
nor U9603 (N_9603,N_8697,N_8702);
and U9604 (N_9604,N_8206,N_8786);
nand U9605 (N_9605,N_8817,N_8354);
nor U9606 (N_9606,N_8419,N_8551);
or U9607 (N_9607,N_8593,N_8556);
or U9608 (N_9608,N_8314,N_8348);
or U9609 (N_9609,N_8583,N_8065);
nor U9610 (N_9610,N_8650,N_8130);
nor U9611 (N_9611,N_8122,N_8100);
and U9612 (N_9612,N_8949,N_8052);
nand U9613 (N_9613,N_8883,N_8166);
or U9614 (N_9614,N_8209,N_8616);
xor U9615 (N_9615,N_8264,N_8992);
nor U9616 (N_9616,N_8967,N_8867);
or U9617 (N_9617,N_8427,N_8689);
or U9618 (N_9618,N_8805,N_8096);
nand U9619 (N_9619,N_8212,N_8029);
nand U9620 (N_9620,N_8592,N_8508);
nor U9621 (N_9621,N_8775,N_8369);
or U9622 (N_9622,N_8772,N_8056);
nand U9623 (N_9623,N_8445,N_8552);
nand U9624 (N_9624,N_8079,N_8565);
nor U9625 (N_9625,N_8114,N_8082);
and U9626 (N_9626,N_8274,N_8708);
and U9627 (N_9627,N_8517,N_8040);
xor U9628 (N_9628,N_8103,N_8390);
nand U9629 (N_9629,N_8433,N_8316);
nand U9630 (N_9630,N_8038,N_8014);
nor U9631 (N_9631,N_8717,N_8825);
nand U9632 (N_9632,N_8695,N_8110);
nor U9633 (N_9633,N_8478,N_8569);
xor U9634 (N_9634,N_8006,N_8724);
nand U9635 (N_9635,N_8279,N_8328);
xnor U9636 (N_9636,N_8887,N_8075);
nor U9637 (N_9637,N_8976,N_8812);
nor U9638 (N_9638,N_8190,N_8932);
nor U9639 (N_9639,N_8458,N_8532);
or U9640 (N_9640,N_8367,N_8891);
and U9641 (N_9641,N_8326,N_8241);
xnor U9642 (N_9642,N_8342,N_8682);
or U9643 (N_9643,N_8662,N_8817);
xnor U9644 (N_9644,N_8982,N_8869);
or U9645 (N_9645,N_8150,N_8843);
nor U9646 (N_9646,N_8997,N_8765);
or U9647 (N_9647,N_8725,N_8070);
nor U9648 (N_9648,N_8232,N_8350);
and U9649 (N_9649,N_8334,N_8336);
nor U9650 (N_9650,N_8387,N_8651);
nor U9651 (N_9651,N_8732,N_8255);
nor U9652 (N_9652,N_8645,N_8074);
and U9653 (N_9653,N_8271,N_8648);
xnor U9654 (N_9654,N_8715,N_8105);
nor U9655 (N_9655,N_8376,N_8721);
xor U9656 (N_9656,N_8461,N_8699);
and U9657 (N_9657,N_8335,N_8853);
xnor U9658 (N_9658,N_8723,N_8427);
nand U9659 (N_9659,N_8852,N_8669);
nor U9660 (N_9660,N_8692,N_8230);
nor U9661 (N_9661,N_8991,N_8693);
or U9662 (N_9662,N_8498,N_8157);
nor U9663 (N_9663,N_8825,N_8863);
nand U9664 (N_9664,N_8061,N_8620);
nand U9665 (N_9665,N_8412,N_8698);
xnor U9666 (N_9666,N_8148,N_8058);
and U9667 (N_9667,N_8010,N_8349);
nand U9668 (N_9668,N_8512,N_8162);
and U9669 (N_9669,N_8978,N_8703);
xnor U9670 (N_9670,N_8799,N_8651);
nand U9671 (N_9671,N_8777,N_8609);
nand U9672 (N_9672,N_8958,N_8727);
or U9673 (N_9673,N_8732,N_8223);
or U9674 (N_9674,N_8681,N_8935);
xor U9675 (N_9675,N_8526,N_8862);
or U9676 (N_9676,N_8952,N_8153);
or U9677 (N_9677,N_8356,N_8421);
nand U9678 (N_9678,N_8400,N_8211);
xor U9679 (N_9679,N_8913,N_8238);
nor U9680 (N_9680,N_8255,N_8555);
and U9681 (N_9681,N_8869,N_8094);
and U9682 (N_9682,N_8515,N_8056);
nand U9683 (N_9683,N_8803,N_8270);
nor U9684 (N_9684,N_8339,N_8843);
xor U9685 (N_9685,N_8190,N_8603);
and U9686 (N_9686,N_8991,N_8790);
nor U9687 (N_9687,N_8619,N_8037);
and U9688 (N_9688,N_8464,N_8535);
xor U9689 (N_9689,N_8741,N_8170);
nor U9690 (N_9690,N_8168,N_8733);
nor U9691 (N_9691,N_8079,N_8579);
or U9692 (N_9692,N_8739,N_8099);
nor U9693 (N_9693,N_8697,N_8979);
or U9694 (N_9694,N_8051,N_8065);
nor U9695 (N_9695,N_8718,N_8993);
nand U9696 (N_9696,N_8542,N_8240);
nor U9697 (N_9697,N_8927,N_8229);
nand U9698 (N_9698,N_8603,N_8697);
and U9699 (N_9699,N_8337,N_8633);
nor U9700 (N_9700,N_8301,N_8541);
nor U9701 (N_9701,N_8979,N_8418);
and U9702 (N_9702,N_8607,N_8322);
xor U9703 (N_9703,N_8058,N_8036);
xnor U9704 (N_9704,N_8904,N_8704);
xor U9705 (N_9705,N_8959,N_8696);
nor U9706 (N_9706,N_8949,N_8178);
nor U9707 (N_9707,N_8243,N_8510);
or U9708 (N_9708,N_8614,N_8024);
and U9709 (N_9709,N_8859,N_8031);
and U9710 (N_9710,N_8125,N_8449);
xor U9711 (N_9711,N_8665,N_8254);
xnor U9712 (N_9712,N_8485,N_8201);
nand U9713 (N_9713,N_8623,N_8520);
nor U9714 (N_9714,N_8614,N_8131);
or U9715 (N_9715,N_8013,N_8121);
xor U9716 (N_9716,N_8385,N_8526);
and U9717 (N_9717,N_8677,N_8186);
and U9718 (N_9718,N_8902,N_8066);
nand U9719 (N_9719,N_8252,N_8077);
and U9720 (N_9720,N_8541,N_8551);
or U9721 (N_9721,N_8712,N_8987);
nand U9722 (N_9722,N_8537,N_8441);
nor U9723 (N_9723,N_8740,N_8792);
nor U9724 (N_9724,N_8008,N_8235);
nor U9725 (N_9725,N_8973,N_8830);
nand U9726 (N_9726,N_8441,N_8857);
nor U9727 (N_9727,N_8182,N_8577);
or U9728 (N_9728,N_8380,N_8977);
or U9729 (N_9729,N_8199,N_8643);
xor U9730 (N_9730,N_8102,N_8484);
xnor U9731 (N_9731,N_8084,N_8034);
and U9732 (N_9732,N_8584,N_8508);
xor U9733 (N_9733,N_8505,N_8812);
xnor U9734 (N_9734,N_8038,N_8025);
nand U9735 (N_9735,N_8192,N_8215);
and U9736 (N_9736,N_8887,N_8262);
and U9737 (N_9737,N_8478,N_8804);
or U9738 (N_9738,N_8286,N_8759);
and U9739 (N_9739,N_8106,N_8285);
nor U9740 (N_9740,N_8190,N_8543);
nor U9741 (N_9741,N_8413,N_8326);
nand U9742 (N_9742,N_8235,N_8123);
nand U9743 (N_9743,N_8848,N_8014);
nor U9744 (N_9744,N_8441,N_8505);
nor U9745 (N_9745,N_8897,N_8779);
xor U9746 (N_9746,N_8909,N_8793);
and U9747 (N_9747,N_8516,N_8645);
and U9748 (N_9748,N_8774,N_8908);
nor U9749 (N_9749,N_8114,N_8497);
nand U9750 (N_9750,N_8993,N_8945);
or U9751 (N_9751,N_8594,N_8243);
and U9752 (N_9752,N_8611,N_8347);
nand U9753 (N_9753,N_8493,N_8601);
nand U9754 (N_9754,N_8034,N_8312);
xor U9755 (N_9755,N_8044,N_8607);
xor U9756 (N_9756,N_8324,N_8387);
nor U9757 (N_9757,N_8101,N_8260);
xnor U9758 (N_9758,N_8939,N_8612);
nand U9759 (N_9759,N_8698,N_8909);
and U9760 (N_9760,N_8442,N_8523);
nand U9761 (N_9761,N_8804,N_8773);
xor U9762 (N_9762,N_8335,N_8310);
xor U9763 (N_9763,N_8101,N_8331);
nor U9764 (N_9764,N_8502,N_8388);
nand U9765 (N_9765,N_8640,N_8657);
or U9766 (N_9766,N_8850,N_8162);
xor U9767 (N_9767,N_8395,N_8361);
nor U9768 (N_9768,N_8496,N_8010);
nand U9769 (N_9769,N_8095,N_8150);
nor U9770 (N_9770,N_8438,N_8232);
and U9771 (N_9771,N_8146,N_8323);
xor U9772 (N_9772,N_8708,N_8940);
or U9773 (N_9773,N_8474,N_8230);
nor U9774 (N_9774,N_8149,N_8974);
xor U9775 (N_9775,N_8856,N_8982);
or U9776 (N_9776,N_8281,N_8115);
and U9777 (N_9777,N_8307,N_8550);
xnor U9778 (N_9778,N_8040,N_8428);
nand U9779 (N_9779,N_8565,N_8259);
nor U9780 (N_9780,N_8558,N_8513);
and U9781 (N_9781,N_8352,N_8691);
xor U9782 (N_9782,N_8637,N_8066);
or U9783 (N_9783,N_8431,N_8741);
nand U9784 (N_9784,N_8470,N_8962);
nor U9785 (N_9785,N_8023,N_8694);
xnor U9786 (N_9786,N_8461,N_8384);
xnor U9787 (N_9787,N_8480,N_8501);
xor U9788 (N_9788,N_8440,N_8757);
and U9789 (N_9789,N_8178,N_8879);
xnor U9790 (N_9790,N_8821,N_8627);
nand U9791 (N_9791,N_8322,N_8012);
nand U9792 (N_9792,N_8720,N_8425);
nand U9793 (N_9793,N_8501,N_8709);
and U9794 (N_9794,N_8236,N_8779);
or U9795 (N_9795,N_8874,N_8657);
nand U9796 (N_9796,N_8923,N_8615);
nand U9797 (N_9797,N_8067,N_8116);
nor U9798 (N_9798,N_8070,N_8001);
nor U9799 (N_9799,N_8711,N_8136);
nor U9800 (N_9800,N_8174,N_8854);
nand U9801 (N_9801,N_8855,N_8846);
and U9802 (N_9802,N_8558,N_8504);
nand U9803 (N_9803,N_8479,N_8137);
and U9804 (N_9804,N_8353,N_8791);
or U9805 (N_9805,N_8880,N_8946);
or U9806 (N_9806,N_8475,N_8713);
and U9807 (N_9807,N_8242,N_8767);
nand U9808 (N_9808,N_8172,N_8334);
or U9809 (N_9809,N_8664,N_8483);
and U9810 (N_9810,N_8242,N_8267);
nor U9811 (N_9811,N_8567,N_8511);
nand U9812 (N_9812,N_8955,N_8999);
nand U9813 (N_9813,N_8259,N_8301);
xnor U9814 (N_9814,N_8605,N_8192);
nand U9815 (N_9815,N_8652,N_8913);
nor U9816 (N_9816,N_8993,N_8677);
nand U9817 (N_9817,N_8054,N_8174);
xnor U9818 (N_9818,N_8077,N_8057);
nor U9819 (N_9819,N_8785,N_8978);
and U9820 (N_9820,N_8568,N_8041);
nor U9821 (N_9821,N_8640,N_8356);
xnor U9822 (N_9822,N_8069,N_8612);
nor U9823 (N_9823,N_8836,N_8108);
or U9824 (N_9824,N_8617,N_8299);
or U9825 (N_9825,N_8591,N_8891);
or U9826 (N_9826,N_8231,N_8797);
nor U9827 (N_9827,N_8078,N_8864);
nand U9828 (N_9828,N_8959,N_8647);
nor U9829 (N_9829,N_8040,N_8989);
nor U9830 (N_9830,N_8115,N_8304);
and U9831 (N_9831,N_8740,N_8115);
or U9832 (N_9832,N_8730,N_8848);
nor U9833 (N_9833,N_8889,N_8544);
and U9834 (N_9834,N_8663,N_8886);
nor U9835 (N_9835,N_8680,N_8375);
and U9836 (N_9836,N_8070,N_8839);
or U9837 (N_9837,N_8279,N_8799);
or U9838 (N_9838,N_8344,N_8751);
or U9839 (N_9839,N_8710,N_8232);
or U9840 (N_9840,N_8494,N_8725);
nand U9841 (N_9841,N_8966,N_8136);
nand U9842 (N_9842,N_8037,N_8822);
and U9843 (N_9843,N_8285,N_8800);
or U9844 (N_9844,N_8793,N_8110);
and U9845 (N_9845,N_8348,N_8073);
nand U9846 (N_9846,N_8366,N_8906);
nand U9847 (N_9847,N_8420,N_8344);
or U9848 (N_9848,N_8543,N_8232);
xnor U9849 (N_9849,N_8901,N_8845);
xor U9850 (N_9850,N_8665,N_8447);
xnor U9851 (N_9851,N_8380,N_8579);
nand U9852 (N_9852,N_8024,N_8590);
nor U9853 (N_9853,N_8387,N_8412);
nand U9854 (N_9854,N_8535,N_8432);
nor U9855 (N_9855,N_8217,N_8509);
nand U9856 (N_9856,N_8347,N_8344);
or U9857 (N_9857,N_8780,N_8670);
xnor U9858 (N_9858,N_8520,N_8638);
and U9859 (N_9859,N_8933,N_8806);
or U9860 (N_9860,N_8435,N_8123);
nor U9861 (N_9861,N_8876,N_8634);
and U9862 (N_9862,N_8498,N_8046);
and U9863 (N_9863,N_8115,N_8520);
nor U9864 (N_9864,N_8750,N_8245);
and U9865 (N_9865,N_8714,N_8352);
or U9866 (N_9866,N_8054,N_8936);
xor U9867 (N_9867,N_8343,N_8063);
nand U9868 (N_9868,N_8933,N_8207);
or U9869 (N_9869,N_8097,N_8481);
nor U9870 (N_9870,N_8000,N_8030);
and U9871 (N_9871,N_8631,N_8345);
or U9872 (N_9872,N_8922,N_8813);
and U9873 (N_9873,N_8905,N_8401);
nand U9874 (N_9874,N_8599,N_8240);
nor U9875 (N_9875,N_8511,N_8387);
or U9876 (N_9876,N_8852,N_8788);
xnor U9877 (N_9877,N_8246,N_8562);
or U9878 (N_9878,N_8022,N_8719);
nor U9879 (N_9879,N_8817,N_8151);
nor U9880 (N_9880,N_8237,N_8227);
nand U9881 (N_9881,N_8349,N_8566);
and U9882 (N_9882,N_8271,N_8596);
nand U9883 (N_9883,N_8831,N_8648);
or U9884 (N_9884,N_8987,N_8828);
nand U9885 (N_9885,N_8593,N_8114);
and U9886 (N_9886,N_8659,N_8318);
and U9887 (N_9887,N_8187,N_8501);
nor U9888 (N_9888,N_8271,N_8852);
xnor U9889 (N_9889,N_8436,N_8680);
or U9890 (N_9890,N_8985,N_8426);
nand U9891 (N_9891,N_8321,N_8718);
nand U9892 (N_9892,N_8972,N_8325);
nand U9893 (N_9893,N_8663,N_8513);
xnor U9894 (N_9894,N_8830,N_8141);
nand U9895 (N_9895,N_8402,N_8733);
and U9896 (N_9896,N_8037,N_8516);
nor U9897 (N_9897,N_8617,N_8540);
xnor U9898 (N_9898,N_8147,N_8677);
or U9899 (N_9899,N_8367,N_8399);
nor U9900 (N_9900,N_8716,N_8689);
nor U9901 (N_9901,N_8306,N_8525);
nor U9902 (N_9902,N_8785,N_8410);
or U9903 (N_9903,N_8239,N_8741);
or U9904 (N_9904,N_8346,N_8442);
nand U9905 (N_9905,N_8237,N_8833);
xnor U9906 (N_9906,N_8422,N_8292);
nor U9907 (N_9907,N_8569,N_8589);
xnor U9908 (N_9908,N_8186,N_8600);
and U9909 (N_9909,N_8149,N_8295);
nor U9910 (N_9910,N_8934,N_8206);
xor U9911 (N_9911,N_8554,N_8350);
and U9912 (N_9912,N_8171,N_8260);
nor U9913 (N_9913,N_8240,N_8667);
and U9914 (N_9914,N_8525,N_8639);
or U9915 (N_9915,N_8626,N_8108);
or U9916 (N_9916,N_8295,N_8905);
and U9917 (N_9917,N_8055,N_8147);
or U9918 (N_9918,N_8906,N_8022);
nand U9919 (N_9919,N_8943,N_8261);
xor U9920 (N_9920,N_8093,N_8524);
xnor U9921 (N_9921,N_8206,N_8569);
nand U9922 (N_9922,N_8303,N_8360);
xor U9923 (N_9923,N_8621,N_8196);
nand U9924 (N_9924,N_8032,N_8292);
nand U9925 (N_9925,N_8098,N_8417);
nor U9926 (N_9926,N_8534,N_8054);
and U9927 (N_9927,N_8772,N_8801);
nand U9928 (N_9928,N_8263,N_8488);
xor U9929 (N_9929,N_8953,N_8594);
or U9930 (N_9930,N_8763,N_8500);
nor U9931 (N_9931,N_8188,N_8373);
and U9932 (N_9932,N_8693,N_8998);
or U9933 (N_9933,N_8820,N_8335);
xnor U9934 (N_9934,N_8486,N_8762);
and U9935 (N_9935,N_8636,N_8389);
and U9936 (N_9936,N_8256,N_8522);
and U9937 (N_9937,N_8845,N_8167);
or U9938 (N_9938,N_8503,N_8012);
nand U9939 (N_9939,N_8993,N_8507);
and U9940 (N_9940,N_8161,N_8489);
and U9941 (N_9941,N_8075,N_8230);
nor U9942 (N_9942,N_8237,N_8486);
or U9943 (N_9943,N_8351,N_8187);
nor U9944 (N_9944,N_8347,N_8251);
xnor U9945 (N_9945,N_8945,N_8774);
xnor U9946 (N_9946,N_8399,N_8279);
nand U9947 (N_9947,N_8226,N_8899);
nand U9948 (N_9948,N_8650,N_8576);
xnor U9949 (N_9949,N_8164,N_8881);
and U9950 (N_9950,N_8372,N_8057);
nand U9951 (N_9951,N_8413,N_8637);
nor U9952 (N_9952,N_8878,N_8395);
or U9953 (N_9953,N_8959,N_8149);
or U9954 (N_9954,N_8744,N_8148);
or U9955 (N_9955,N_8696,N_8785);
nand U9956 (N_9956,N_8815,N_8183);
xnor U9957 (N_9957,N_8060,N_8722);
nand U9958 (N_9958,N_8230,N_8163);
xor U9959 (N_9959,N_8758,N_8531);
nand U9960 (N_9960,N_8668,N_8065);
and U9961 (N_9961,N_8068,N_8869);
xor U9962 (N_9962,N_8673,N_8180);
xnor U9963 (N_9963,N_8424,N_8018);
xnor U9964 (N_9964,N_8249,N_8762);
xor U9965 (N_9965,N_8572,N_8091);
and U9966 (N_9966,N_8677,N_8894);
and U9967 (N_9967,N_8888,N_8137);
and U9968 (N_9968,N_8302,N_8661);
and U9969 (N_9969,N_8817,N_8255);
or U9970 (N_9970,N_8460,N_8108);
or U9971 (N_9971,N_8387,N_8027);
nand U9972 (N_9972,N_8070,N_8398);
or U9973 (N_9973,N_8414,N_8146);
or U9974 (N_9974,N_8681,N_8787);
nand U9975 (N_9975,N_8289,N_8917);
xnor U9976 (N_9976,N_8644,N_8922);
nand U9977 (N_9977,N_8164,N_8781);
and U9978 (N_9978,N_8457,N_8152);
nand U9979 (N_9979,N_8371,N_8363);
nand U9980 (N_9980,N_8944,N_8032);
and U9981 (N_9981,N_8778,N_8440);
and U9982 (N_9982,N_8506,N_8702);
nand U9983 (N_9983,N_8250,N_8995);
nor U9984 (N_9984,N_8061,N_8222);
and U9985 (N_9985,N_8760,N_8638);
nand U9986 (N_9986,N_8751,N_8382);
and U9987 (N_9987,N_8961,N_8255);
nor U9988 (N_9988,N_8500,N_8514);
and U9989 (N_9989,N_8026,N_8782);
or U9990 (N_9990,N_8277,N_8260);
nand U9991 (N_9991,N_8766,N_8727);
nor U9992 (N_9992,N_8161,N_8461);
or U9993 (N_9993,N_8996,N_8195);
nand U9994 (N_9994,N_8763,N_8108);
xor U9995 (N_9995,N_8667,N_8556);
and U9996 (N_9996,N_8555,N_8208);
or U9997 (N_9997,N_8919,N_8686);
and U9998 (N_9998,N_8824,N_8211);
nand U9999 (N_9999,N_8920,N_8020);
nor U10000 (N_10000,N_9927,N_9662);
xor U10001 (N_10001,N_9586,N_9789);
and U10002 (N_10002,N_9482,N_9621);
and U10003 (N_10003,N_9282,N_9368);
and U10004 (N_10004,N_9244,N_9801);
and U10005 (N_10005,N_9934,N_9591);
and U10006 (N_10006,N_9811,N_9148);
and U10007 (N_10007,N_9111,N_9854);
and U10008 (N_10008,N_9096,N_9883);
xnor U10009 (N_10009,N_9067,N_9821);
xnor U10010 (N_10010,N_9397,N_9572);
xnor U10011 (N_10011,N_9108,N_9751);
nand U10012 (N_10012,N_9750,N_9887);
or U10013 (N_10013,N_9851,N_9243);
xnor U10014 (N_10014,N_9036,N_9951);
xor U10015 (N_10015,N_9076,N_9997);
xnor U10016 (N_10016,N_9372,N_9554);
nor U10017 (N_10017,N_9126,N_9375);
or U10018 (N_10018,N_9156,N_9240);
nor U10019 (N_10019,N_9792,N_9710);
nor U10020 (N_10020,N_9944,N_9063);
nand U10021 (N_10021,N_9037,N_9538);
and U10022 (N_10022,N_9190,N_9344);
nor U10023 (N_10023,N_9151,N_9314);
or U10024 (N_10024,N_9549,N_9676);
or U10025 (N_10025,N_9677,N_9866);
nor U10026 (N_10026,N_9465,N_9128);
or U10027 (N_10027,N_9564,N_9589);
xor U10028 (N_10028,N_9288,N_9868);
and U10029 (N_10029,N_9762,N_9026);
xor U10030 (N_10030,N_9226,N_9786);
xnor U10031 (N_10031,N_9100,N_9311);
or U10032 (N_10032,N_9131,N_9115);
nor U10033 (N_10033,N_9628,N_9163);
nor U10034 (N_10034,N_9877,N_9971);
and U10035 (N_10035,N_9203,N_9254);
nand U10036 (N_10036,N_9515,N_9687);
xnor U10037 (N_10037,N_9505,N_9105);
xnor U10038 (N_10038,N_9843,N_9856);
nand U10039 (N_10039,N_9645,N_9988);
nand U10040 (N_10040,N_9656,N_9907);
nor U10041 (N_10041,N_9120,N_9081);
nor U10042 (N_10042,N_9953,N_9438);
xor U10043 (N_10043,N_9297,N_9134);
or U10044 (N_10044,N_9270,N_9747);
nand U10045 (N_10045,N_9954,N_9265);
xnor U10046 (N_10046,N_9818,N_9376);
xor U10047 (N_10047,N_9742,N_9839);
nand U10048 (N_10048,N_9347,N_9999);
nor U10049 (N_10049,N_9822,N_9178);
xor U10050 (N_10050,N_9514,N_9675);
and U10051 (N_10051,N_9929,N_9109);
or U10052 (N_10052,N_9541,N_9247);
nand U10053 (N_10053,N_9443,N_9285);
xor U10054 (N_10054,N_9606,N_9924);
xor U10055 (N_10055,N_9449,N_9977);
or U10056 (N_10056,N_9604,N_9570);
xnor U10057 (N_10057,N_9183,N_9406);
nor U10058 (N_10058,N_9648,N_9850);
and U10059 (N_10059,N_9776,N_9601);
nand U10060 (N_10060,N_9880,N_9536);
or U10061 (N_10061,N_9500,N_9419);
or U10062 (N_10062,N_9364,N_9356);
xor U10063 (N_10063,N_9852,N_9434);
or U10064 (N_10064,N_9415,N_9758);
nor U10065 (N_10065,N_9638,N_9739);
or U10066 (N_10066,N_9292,N_9595);
xnor U10067 (N_10067,N_9813,N_9040);
and U10068 (N_10068,N_9234,N_9989);
nor U10069 (N_10069,N_9272,N_9587);
nor U10070 (N_10070,N_9761,N_9808);
xnor U10071 (N_10071,N_9031,N_9925);
xor U10072 (N_10072,N_9329,N_9597);
nand U10073 (N_10073,N_9567,N_9117);
and U10074 (N_10074,N_9407,N_9412);
or U10075 (N_10075,N_9011,N_9476);
nor U10076 (N_10076,N_9057,N_9909);
or U10077 (N_10077,N_9043,N_9535);
xnor U10078 (N_10078,N_9847,N_9640);
nand U10079 (N_10079,N_9185,N_9295);
xnor U10080 (N_10080,N_9030,N_9655);
xor U10081 (N_10081,N_9623,N_9740);
nor U10082 (N_10082,N_9552,N_9167);
or U10083 (N_10083,N_9339,N_9889);
nor U10084 (N_10084,N_9310,N_9599);
and U10085 (N_10085,N_9672,N_9530);
xor U10086 (N_10086,N_9468,N_9211);
xnor U10087 (N_10087,N_9905,N_9870);
nand U10088 (N_10088,N_9881,N_9408);
nand U10089 (N_10089,N_9200,N_9281);
nor U10090 (N_10090,N_9715,N_9213);
xor U10091 (N_10091,N_9766,N_9534);
xnor U10092 (N_10092,N_9689,N_9634);
and U10093 (N_10093,N_9803,N_9919);
nor U10094 (N_10094,N_9700,N_9336);
and U10095 (N_10095,N_9009,N_9809);
and U10096 (N_10096,N_9838,N_9362);
and U10097 (N_10097,N_9466,N_9106);
nand U10098 (N_10098,N_9738,N_9760);
nand U10099 (N_10099,N_9262,N_9194);
and U10100 (N_10100,N_9216,N_9256);
and U10101 (N_10101,N_9935,N_9901);
nand U10102 (N_10102,N_9135,N_9097);
and U10103 (N_10103,N_9754,N_9475);
nor U10104 (N_10104,N_9635,N_9331);
nand U10105 (N_10105,N_9752,N_9958);
nor U10106 (N_10106,N_9195,N_9725);
nor U10107 (N_10107,N_9410,N_9246);
nand U10108 (N_10108,N_9706,N_9713);
nand U10109 (N_10109,N_9592,N_9721);
nand U10110 (N_10110,N_9420,N_9723);
xnor U10111 (N_10111,N_9957,N_9093);
or U10112 (N_10112,N_9652,N_9326);
nor U10113 (N_10113,N_9551,N_9222);
and U10114 (N_10114,N_9196,N_9678);
xnor U10115 (N_10115,N_9307,N_9986);
and U10116 (N_10116,N_9517,N_9188);
xnor U10117 (N_10117,N_9576,N_9334);
nand U10118 (N_10118,N_9546,N_9969);
or U10119 (N_10119,N_9473,N_9321);
xor U10120 (N_10120,N_9781,N_9278);
nand U10121 (N_10121,N_9817,N_9296);
xor U10122 (N_10122,N_9258,N_9367);
and U10123 (N_10123,N_9668,N_9705);
nand U10124 (N_10124,N_9125,N_9488);
xnor U10125 (N_10125,N_9284,N_9335);
or U10126 (N_10126,N_9699,N_9273);
nand U10127 (N_10127,N_9442,N_9630);
or U10128 (N_10128,N_9756,N_9663);
xnor U10129 (N_10129,N_9757,N_9064);
nor U10130 (N_10130,N_9658,N_9562);
or U10131 (N_10131,N_9123,N_9012);
and U10132 (N_10132,N_9569,N_9206);
xnor U10133 (N_10133,N_9351,N_9038);
nand U10134 (N_10134,N_9348,N_9483);
nor U10135 (N_10135,N_9769,N_9290);
or U10136 (N_10136,N_9926,N_9718);
and U10137 (N_10137,N_9796,N_9414);
nand U10138 (N_10138,N_9902,N_9000);
or U10139 (N_10139,N_9046,N_9617);
or U10140 (N_10140,N_9006,N_9153);
xnor U10141 (N_10141,N_9859,N_9354);
xnor U10142 (N_10142,N_9070,N_9614);
and U10143 (N_10143,N_9886,N_9893);
or U10144 (N_10144,N_9140,N_9379);
or U10145 (N_10145,N_9826,N_9622);
nand U10146 (N_10146,N_9186,N_9479);
nor U10147 (N_10147,N_9771,N_9582);
nor U10148 (N_10148,N_9299,N_9939);
xor U10149 (N_10149,N_9921,N_9054);
nand U10150 (N_10150,N_9118,N_9960);
or U10151 (N_10151,N_9452,N_9943);
or U10152 (N_10152,N_9133,N_9114);
and U10153 (N_10153,N_9615,N_9707);
nand U10154 (N_10154,N_9229,N_9719);
or U10155 (N_10155,N_9914,N_9337);
nor U10156 (N_10156,N_9386,N_9812);
xor U10157 (N_10157,N_9995,N_9268);
xnor U10158 (N_10158,N_9202,N_9059);
xor U10159 (N_10159,N_9523,N_9861);
nor U10160 (N_10160,N_9961,N_9627);
nor U10161 (N_10161,N_9474,N_9230);
or U10162 (N_10162,N_9933,N_9956);
or U10163 (N_10163,N_9704,N_9155);
or U10164 (N_10164,N_9145,N_9127);
nand U10165 (N_10165,N_9895,N_9755);
nor U10166 (N_10166,N_9524,N_9330);
and U10167 (N_10167,N_9333,N_9529);
nand U10168 (N_10168,N_9249,N_9071);
or U10169 (N_10169,N_9637,N_9189);
or U10170 (N_10170,N_9834,N_9875);
nor U10171 (N_10171,N_9355,N_9965);
or U10172 (N_10172,N_9981,N_9144);
and U10173 (N_10173,N_9045,N_9619);
nand U10174 (N_10174,N_9429,N_9942);
or U10175 (N_10175,N_9644,N_9210);
or U10176 (N_10176,N_9426,N_9504);
or U10177 (N_10177,N_9382,N_9481);
or U10178 (N_10178,N_9112,N_9147);
nand U10179 (N_10179,N_9293,N_9065);
or U10180 (N_10180,N_9735,N_9074);
nor U10181 (N_10181,N_9179,N_9277);
and U10182 (N_10182,N_9319,N_9701);
nand U10183 (N_10183,N_9722,N_9802);
and U10184 (N_10184,N_9209,N_9736);
and U10185 (N_10185,N_9346,N_9447);
and U10186 (N_10186,N_9280,N_9132);
nand U10187 (N_10187,N_9358,N_9840);
xor U10188 (N_10188,N_9435,N_9389);
and U10189 (N_10189,N_9805,N_9413);
nor U10190 (N_10190,N_9983,N_9894);
nand U10191 (N_10191,N_9651,N_9323);
or U10192 (N_10192,N_9952,N_9891);
or U10193 (N_10193,N_9159,N_9274);
nor U10194 (N_10194,N_9171,N_9955);
nand U10195 (N_10195,N_9287,N_9425);
nand U10196 (N_10196,N_9494,N_9033);
or U10197 (N_10197,N_9625,N_9398);
xor U10198 (N_10198,N_9936,N_9913);
or U10199 (N_10199,N_9824,N_9403);
xor U10200 (N_10200,N_9142,N_9102);
nor U10201 (N_10201,N_9343,N_9199);
or U10202 (N_10202,N_9309,N_9729);
and U10203 (N_10203,N_9978,N_9568);
and U10204 (N_10204,N_9791,N_9401);
xor U10205 (N_10205,N_9017,N_9322);
nand U10206 (N_10206,N_9578,N_9400);
nor U10207 (N_10207,N_9034,N_9799);
xnor U10208 (N_10208,N_9224,N_9680);
xor U10209 (N_10209,N_9490,N_9657);
nor U10210 (N_10210,N_9828,N_9027);
and U10211 (N_10211,N_9876,N_9260);
and U10212 (N_10212,N_9816,N_9605);
xnor U10213 (N_10213,N_9320,N_9324);
or U10214 (N_10214,N_9841,N_9207);
or U10215 (N_10215,N_9208,N_9968);
xnor U10216 (N_10216,N_9214,N_9363);
and U10217 (N_10217,N_9533,N_9302);
nand U10218 (N_10218,N_9044,N_9394);
nor U10219 (N_10219,N_9069,N_9306);
and U10220 (N_10220,N_9772,N_9888);
nor U10221 (N_10221,N_9787,N_9647);
and U10222 (N_10222,N_9395,N_9584);
nor U10223 (N_10223,N_9906,N_9985);
nand U10224 (N_10224,N_9528,N_9423);
or U10225 (N_10225,N_9350,N_9378);
nor U10226 (N_10226,N_9765,N_9827);
or U10227 (N_10227,N_9823,N_9225);
and U10228 (N_10228,N_9922,N_9055);
and U10229 (N_10229,N_9782,N_9779);
xnor U10230 (N_10230,N_9431,N_9519);
and U10231 (N_10231,N_9377,N_9191);
or U10232 (N_10232,N_9422,N_9365);
or U10233 (N_10233,N_9393,N_9618);
nor U10234 (N_10234,N_9884,N_9015);
and U10235 (N_10235,N_9079,N_9370);
nand U10236 (N_10236,N_9897,N_9231);
or U10237 (N_10237,N_9690,N_9962);
and U10238 (N_10238,N_9094,N_9556);
nand U10239 (N_10239,N_9836,N_9531);
or U10240 (N_10240,N_9165,N_9716);
or U10241 (N_10241,N_9829,N_9478);
nand U10242 (N_10242,N_9869,N_9219);
nor U10243 (N_10243,N_9930,N_9472);
nor U10244 (N_10244,N_9918,N_9172);
and U10245 (N_10245,N_9708,N_9609);
or U10246 (N_10246,N_9237,N_9416);
nand U10247 (N_10247,N_9166,N_9021);
nor U10248 (N_10248,N_9305,N_9205);
or U10249 (N_10249,N_9506,N_9301);
or U10250 (N_10250,N_9542,N_9810);
and U10251 (N_10251,N_9463,N_9255);
and U10252 (N_10252,N_9608,N_9220);
or U10253 (N_10253,N_9402,N_9874);
nor U10254 (N_10254,N_9062,N_9795);
nand U10255 (N_10255,N_9685,N_9325);
or U10256 (N_10256,N_9650,N_9432);
xnor U10257 (N_10257,N_9746,N_9316);
or U10258 (N_10258,N_9169,N_9182);
nand U10259 (N_10259,N_9223,N_9124);
or U10260 (N_10260,N_9469,N_9684);
xor U10261 (N_10261,N_9660,N_9485);
and U10262 (N_10262,N_9724,N_9464);
nor U10263 (N_10263,N_9221,N_9641);
xnor U10264 (N_10264,N_9904,N_9732);
nor U10265 (N_10265,N_9555,N_9399);
nand U10266 (N_10266,N_9252,N_9497);
nand U10267 (N_10267,N_9516,N_9947);
nand U10268 (N_10268,N_9227,N_9238);
nor U10269 (N_10269,N_9215,N_9193);
xnor U10270 (N_10270,N_9137,N_9631);
or U10271 (N_10271,N_9670,N_9058);
and U10272 (N_10272,N_9543,N_9259);
nand U10273 (N_10273,N_9276,N_9427);
nor U10274 (N_10274,N_9987,N_9099);
and U10275 (N_10275,N_9783,N_9571);
and U10276 (N_10276,N_9804,N_9639);
nand U10277 (N_10277,N_9982,N_9257);
nor U10278 (N_10278,N_9232,N_9937);
nand U10279 (N_10279,N_9201,N_9122);
xnor U10280 (N_10280,N_9051,N_9486);
nand U10281 (N_10281,N_9990,N_9770);
or U10282 (N_10282,N_9371,N_9090);
xor U10283 (N_10283,N_9418,N_9430);
and U10284 (N_10284,N_9581,N_9844);
xnor U10285 (N_10285,N_9712,N_9304);
or U10286 (N_10286,N_9973,N_9882);
or U10287 (N_10287,N_9168,N_9073);
xor U10288 (N_10288,N_9768,N_9734);
and U10289 (N_10289,N_9218,N_9161);
xor U10290 (N_10290,N_9912,N_9298);
and U10291 (N_10291,N_9527,N_9948);
or U10292 (N_10292,N_9646,N_9673);
nand U10293 (N_10293,N_9439,N_9610);
and U10294 (N_10294,N_9553,N_9263);
xnor U10295 (N_10295,N_9941,N_9342);
nand U10296 (N_10296,N_9313,N_9717);
and U10297 (N_10297,N_9896,N_9077);
or U10298 (N_10298,N_9373,N_9437);
xnor U10299 (N_10299,N_9518,N_9271);
xnor U10300 (N_10300,N_9773,N_9674);
xor U10301 (N_10301,N_9404,N_9248);
nand U10302 (N_10302,N_9629,N_9136);
or U10303 (N_10303,N_9853,N_9052);
or U10304 (N_10304,N_9993,N_9184);
xnor U10305 (N_10305,N_9825,N_9537);
xnor U10306 (N_10306,N_9042,N_9020);
and U10307 (N_10307,N_9060,N_9477);
nand U10308 (N_10308,N_9975,N_9484);
nor U10309 (N_10309,N_9023,N_9411);
xor U10310 (N_10310,N_9460,N_9967);
or U10311 (N_10311,N_9085,N_9780);
and U10312 (N_10312,N_9019,N_9900);
xor U10313 (N_10313,N_9048,N_9733);
xnor U10314 (N_10314,N_9217,N_9087);
or U10315 (N_10315,N_9139,N_9175);
or U10316 (N_10316,N_9558,N_9387);
and U10317 (N_10317,N_9121,N_9632);
nor U10318 (N_10318,N_9790,N_9970);
nand U10319 (N_10319,N_9286,N_9509);
or U10320 (N_10320,N_9945,N_9696);
and U10321 (N_10321,N_9714,N_9003);
and U10322 (N_10322,N_9830,N_9308);
xnor U10323 (N_10323,N_9462,N_9984);
or U10324 (N_10324,N_9204,N_9300);
nor U10325 (N_10325,N_9119,N_9149);
nand U10326 (N_10326,N_9777,N_9600);
nor U10327 (N_10327,N_9384,N_9080);
or U10328 (N_10328,N_9908,N_9848);
nor U10329 (N_10329,N_9831,N_9594);
xnor U10330 (N_10330,N_9833,N_9459);
xnor U10331 (N_10331,N_9580,N_9158);
nor U10332 (N_10332,N_9759,N_9498);
xnor U10333 (N_10333,N_9095,N_9845);
xnor U10334 (N_10334,N_9078,N_9010);
or U10335 (N_10335,N_9669,N_9775);
and U10336 (N_10336,N_9612,N_9512);
nand U10337 (N_10337,N_9561,N_9745);
nand U10338 (N_10338,N_9560,N_9154);
xnor U10339 (N_10339,N_9920,N_9357);
nand U10340 (N_10340,N_9025,N_9892);
xnor U10341 (N_10341,N_9022,N_9865);
or U10342 (N_10342,N_9047,N_9928);
nand U10343 (N_10343,N_9141,N_9949);
and U10344 (N_10344,N_9005,N_9590);
and U10345 (N_10345,N_9940,N_9879);
and U10346 (N_10346,N_9082,N_9837);
nor U10347 (N_10347,N_9764,N_9340);
or U10348 (N_10348,N_9453,N_9832);
nand U10349 (N_10349,N_9731,N_9267);
and U10350 (N_10350,N_9980,N_9711);
xnor U10351 (N_10351,N_9496,N_9098);
and U10352 (N_10352,N_9860,N_9294);
or U10353 (N_10353,N_9671,N_9103);
or U10354 (N_10354,N_9730,N_9511);
xnor U10355 (N_10355,N_9004,N_9550);
xor U10356 (N_10356,N_9867,N_9616);
and U10357 (N_10357,N_9440,N_9428);
xor U10358 (N_10358,N_9016,N_9013);
nor U10359 (N_10359,N_9075,N_9835);
and U10360 (N_10360,N_9522,N_9441);
and U10361 (N_10361,N_9539,N_9446);
nor U10362 (N_10362,N_9726,N_9233);
nand U10363 (N_10363,N_9380,N_9235);
nor U10364 (N_10364,N_9289,N_9814);
nor U10365 (N_10365,N_9857,N_9050);
or U10366 (N_10366,N_9611,N_9433);
or U10367 (N_10367,N_9667,N_9642);
xnor U10368 (N_10368,N_9236,N_9291);
or U10369 (N_10369,N_9162,N_9788);
and U10370 (N_10370,N_9737,N_9250);
nor U10371 (N_10371,N_9266,N_9513);
xor U10372 (N_10372,N_9931,N_9709);
and U10373 (N_10373,N_9396,N_9526);
and U10374 (N_10374,N_9480,N_9525);
and U10375 (N_10375,N_9327,N_9996);
nor U10376 (N_10376,N_9101,N_9899);
xnor U10377 (N_10377,N_9177,N_9510);
or U10378 (N_10378,N_9487,N_9720);
nand U10379 (N_10379,N_9068,N_9332);
nand U10380 (N_10380,N_9283,N_9181);
nand U10381 (N_10381,N_9061,N_9748);
nand U10382 (N_10382,N_9315,N_9966);
nand U10383 (N_10383,N_9691,N_9603);
nor U10384 (N_10384,N_9702,N_9784);
nand U10385 (N_10385,N_9056,N_9007);
xor U10386 (N_10386,N_9053,N_9493);
nand U10387 (N_10387,N_9176,N_9959);
nor U10388 (N_10388,N_9579,N_9885);
xor U10389 (N_10389,N_9653,N_9878);
and U10390 (N_10390,N_9566,N_9807);
or U10391 (N_10391,N_9692,N_9303);
nand U10392 (N_10392,N_9345,N_9338);
xor U10393 (N_10393,N_9938,N_9846);
or U10394 (N_10394,N_9864,N_9091);
or U10395 (N_10395,N_9502,N_9381);
nor U10396 (N_10396,N_9457,N_9636);
nand U10397 (N_10397,N_9089,N_9820);
and U10398 (N_10398,N_9083,N_9383);
xor U10399 (N_10399,N_9198,N_9574);
or U10400 (N_10400,N_9994,N_9963);
nand U10401 (N_10401,N_9228,N_9778);
or U10402 (N_10402,N_9001,N_9454);
nand U10403 (N_10403,N_9688,N_9898);
and U10404 (N_10404,N_9174,N_9349);
and U10405 (N_10405,N_9014,N_9456);
or U10406 (N_10406,N_9950,N_9458);
nand U10407 (N_10407,N_9436,N_9049);
nand U10408 (N_10408,N_9547,N_9915);
or U10409 (N_10409,N_9008,N_9088);
and U10410 (N_10410,N_9279,N_9819);
nand U10411 (N_10411,N_9470,N_9084);
and U10412 (N_10412,N_9317,N_9557);
xnor U10413 (N_10413,N_9374,N_9659);
and U10414 (N_10414,N_9421,N_9116);
nor U10415 (N_10415,N_9002,N_9596);
nor U10416 (N_10416,N_9753,N_9245);
nand U10417 (N_10417,N_9545,N_9150);
nand U10418 (N_10418,N_9275,N_9575);
xor U10419 (N_10419,N_9681,N_9903);
or U10420 (N_10420,N_9501,N_9445);
nor U10421 (N_10421,N_9110,N_9066);
nor U10422 (N_10422,N_9138,N_9024);
or U10423 (N_10423,N_9583,N_9491);
nor U10424 (N_10424,N_9911,N_9559);
or U10425 (N_10425,N_9683,N_9369);
nor U10426 (N_10426,N_9160,N_9242);
or U10427 (N_10427,N_9686,N_9694);
and U10428 (N_10428,N_9890,N_9264);
xnor U10429 (N_10429,N_9104,N_9624);
and U10430 (N_10430,N_9503,N_9703);
xnor U10431 (N_10431,N_9029,N_9863);
and U10432 (N_10432,N_9409,N_9405);
or U10433 (N_10433,N_9917,N_9107);
nand U10434 (N_10434,N_9682,N_9390);
nand U10435 (N_10435,N_9695,N_9593);
xnor U10436 (N_10436,N_9170,N_9444);
nand U10437 (N_10437,N_9360,N_9749);
or U10438 (N_10438,N_9143,N_9241);
and U10439 (N_10439,N_9312,N_9508);
nand U10440 (N_10440,N_9391,N_9858);
or U10441 (N_10441,N_9620,N_9035);
and U10442 (N_10442,N_9192,N_9113);
nor U10443 (N_10443,N_9613,N_9451);
or U10444 (N_10444,N_9388,N_9910);
nand U10445 (N_10445,N_9173,N_9424);
nand U10446 (N_10446,N_9665,N_9666);
or U10447 (N_10447,N_9212,N_9521);
and U10448 (N_10448,N_9157,N_9573);
nor U10449 (N_10449,N_9946,N_9602);
or U10450 (N_10450,N_9697,N_9520);
or U10451 (N_10451,N_9540,N_9146);
or U10452 (N_10452,N_9793,N_9028);
nand U10453 (N_10453,N_9495,N_9643);
or U10454 (N_10454,N_9018,N_9032);
xor U10455 (N_10455,N_9359,N_9072);
and U10456 (N_10456,N_9366,N_9352);
and U10457 (N_10457,N_9626,N_9964);
nor U10458 (N_10458,N_9800,N_9664);
or U10459 (N_10459,N_9743,N_9251);
nand U10460 (N_10460,N_9489,N_9164);
xnor U10461 (N_10461,N_9798,N_9923);
nand U10462 (N_10462,N_9976,N_9341);
nand U10463 (N_10463,N_9842,N_9548);
xnor U10464 (N_10464,N_9180,N_9361);
nand U10465 (N_10465,N_9318,N_9385);
xnor U10466 (N_10466,N_9197,N_9585);
or U10467 (N_10467,N_9727,N_9565);
and U10468 (N_10468,N_9130,N_9239);
nor U10469 (N_10469,N_9261,N_9086);
or U10470 (N_10470,N_9563,N_9806);
nand U10471 (N_10471,N_9129,N_9499);
or U10472 (N_10472,N_9269,N_9392);
xnor U10473 (N_10473,N_9698,N_9187);
or U10474 (N_10474,N_9633,N_9916);
and U10475 (N_10475,N_9253,N_9661);
nand U10476 (N_10476,N_9932,N_9649);
and U10477 (N_10477,N_9815,N_9577);
and U10478 (N_10478,N_9744,N_9588);
nand U10479 (N_10479,N_9763,N_9862);
and U10480 (N_10480,N_9979,N_9873);
nor U10481 (N_10481,N_9607,N_9492);
xnor U10482 (N_10482,N_9461,N_9467);
and U10483 (N_10483,N_9741,N_9871);
xnor U10484 (N_10484,N_9507,N_9767);
nand U10485 (N_10485,N_9544,N_9039);
or U10486 (N_10486,N_9532,N_9654);
nand U10487 (N_10487,N_9693,N_9353);
and U10488 (N_10488,N_9679,N_9450);
xnor U10489 (N_10489,N_9794,N_9785);
nor U10490 (N_10490,N_9471,N_9417);
nor U10491 (N_10491,N_9855,N_9092);
nand U10492 (N_10492,N_9998,N_9728);
and U10493 (N_10493,N_9991,N_9041);
or U10494 (N_10494,N_9872,N_9152);
xor U10495 (N_10495,N_9448,N_9797);
xor U10496 (N_10496,N_9774,N_9974);
or U10497 (N_10497,N_9849,N_9972);
and U10498 (N_10498,N_9992,N_9328);
or U10499 (N_10499,N_9455,N_9598);
nor U10500 (N_10500,N_9612,N_9836);
nor U10501 (N_10501,N_9176,N_9933);
nor U10502 (N_10502,N_9496,N_9763);
and U10503 (N_10503,N_9858,N_9829);
nor U10504 (N_10504,N_9613,N_9972);
nand U10505 (N_10505,N_9911,N_9570);
nor U10506 (N_10506,N_9443,N_9183);
nor U10507 (N_10507,N_9976,N_9298);
xor U10508 (N_10508,N_9252,N_9445);
nand U10509 (N_10509,N_9093,N_9369);
and U10510 (N_10510,N_9696,N_9586);
nand U10511 (N_10511,N_9442,N_9287);
nor U10512 (N_10512,N_9279,N_9454);
nand U10513 (N_10513,N_9010,N_9780);
xnor U10514 (N_10514,N_9825,N_9040);
xnor U10515 (N_10515,N_9102,N_9788);
nor U10516 (N_10516,N_9724,N_9470);
nor U10517 (N_10517,N_9967,N_9374);
xor U10518 (N_10518,N_9450,N_9158);
and U10519 (N_10519,N_9228,N_9802);
nor U10520 (N_10520,N_9874,N_9046);
nand U10521 (N_10521,N_9297,N_9026);
nor U10522 (N_10522,N_9146,N_9719);
nand U10523 (N_10523,N_9075,N_9375);
xnor U10524 (N_10524,N_9756,N_9326);
nand U10525 (N_10525,N_9874,N_9506);
xor U10526 (N_10526,N_9079,N_9641);
or U10527 (N_10527,N_9264,N_9862);
and U10528 (N_10528,N_9138,N_9344);
nor U10529 (N_10529,N_9546,N_9252);
and U10530 (N_10530,N_9477,N_9853);
or U10531 (N_10531,N_9628,N_9739);
or U10532 (N_10532,N_9567,N_9030);
nor U10533 (N_10533,N_9961,N_9657);
nor U10534 (N_10534,N_9498,N_9144);
or U10535 (N_10535,N_9887,N_9117);
or U10536 (N_10536,N_9708,N_9588);
xor U10537 (N_10537,N_9247,N_9154);
or U10538 (N_10538,N_9374,N_9508);
and U10539 (N_10539,N_9287,N_9515);
and U10540 (N_10540,N_9222,N_9853);
or U10541 (N_10541,N_9765,N_9010);
xor U10542 (N_10542,N_9370,N_9816);
or U10543 (N_10543,N_9183,N_9655);
or U10544 (N_10544,N_9744,N_9662);
or U10545 (N_10545,N_9513,N_9752);
xor U10546 (N_10546,N_9252,N_9342);
nor U10547 (N_10547,N_9981,N_9070);
or U10548 (N_10548,N_9045,N_9039);
and U10549 (N_10549,N_9108,N_9656);
nor U10550 (N_10550,N_9477,N_9969);
nor U10551 (N_10551,N_9754,N_9731);
and U10552 (N_10552,N_9469,N_9413);
nor U10553 (N_10553,N_9395,N_9470);
and U10554 (N_10554,N_9948,N_9026);
xnor U10555 (N_10555,N_9365,N_9441);
nand U10556 (N_10556,N_9805,N_9183);
or U10557 (N_10557,N_9198,N_9669);
and U10558 (N_10558,N_9415,N_9728);
xor U10559 (N_10559,N_9480,N_9026);
nor U10560 (N_10560,N_9295,N_9888);
xnor U10561 (N_10561,N_9910,N_9603);
xnor U10562 (N_10562,N_9174,N_9370);
nor U10563 (N_10563,N_9808,N_9661);
and U10564 (N_10564,N_9224,N_9916);
and U10565 (N_10565,N_9537,N_9905);
xnor U10566 (N_10566,N_9668,N_9698);
nand U10567 (N_10567,N_9908,N_9794);
xnor U10568 (N_10568,N_9254,N_9449);
nor U10569 (N_10569,N_9363,N_9345);
xor U10570 (N_10570,N_9249,N_9833);
nand U10571 (N_10571,N_9327,N_9729);
and U10572 (N_10572,N_9094,N_9232);
xor U10573 (N_10573,N_9711,N_9664);
and U10574 (N_10574,N_9496,N_9769);
xor U10575 (N_10575,N_9709,N_9980);
or U10576 (N_10576,N_9340,N_9014);
xnor U10577 (N_10577,N_9873,N_9774);
and U10578 (N_10578,N_9322,N_9867);
or U10579 (N_10579,N_9776,N_9521);
nor U10580 (N_10580,N_9259,N_9250);
and U10581 (N_10581,N_9312,N_9702);
nand U10582 (N_10582,N_9626,N_9830);
xor U10583 (N_10583,N_9820,N_9044);
or U10584 (N_10584,N_9478,N_9882);
and U10585 (N_10585,N_9370,N_9105);
nor U10586 (N_10586,N_9735,N_9861);
nand U10587 (N_10587,N_9120,N_9442);
nand U10588 (N_10588,N_9643,N_9562);
nor U10589 (N_10589,N_9102,N_9962);
and U10590 (N_10590,N_9520,N_9209);
or U10591 (N_10591,N_9566,N_9090);
and U10592 (N_10592,N_9580,N_9060);
nand U10593 (N_10593,N_9713,N_9979);
or U10594 (N_10594,N_9225,N_9846);
nor U10595 (N_10595,N_9653,N_9852);
nor U10596 (N_10596,N_9304,N_9780);
and U10597 (N_10597,N_9513,N_9300);
xnor U10598 (N_10598,N_9761,N_9464);
nor U10599 (N_10599,N_9178,N_9793);
nand U10600 (N_10600,N_9494,N_9084);
nor U10601 (N_10601,N_9532,N_9150);
or U10602 (N_10602,N_9579,N_9700);
nor U10603 (N_10603,N_9804,N_9076);
nor U10604 (N_10604,N_9935,N_9721);
nand U10605 (N_10605,N_9637,N_9538);
nor U10606 (N_10606,N_9124,N_9770);
xor U10607 (N_10607,N_9678,N_9039);
nor U10608 (N_10608,N_9168,N_9010);
nor U10609 (N_10609,N_9212,N_9047);
nor U10610 (N_10610,N_9110,N_9829);
or U10611 (N_10611,N_9130,N_9947);
and U10612 (N_10612,N_9437,N_9571);
nand U10613 (N_10613,N_9669,N_9186);
nand U10614 (N_10614,N_9036,N_9246);
or U10615 (N_10615,N_9678,N_9485);
nor U10616 (N_10616,N_9325,N_9941);
nand U10617 (N_10617,N_9803,N_9171);
xor U10618 (N_10618,N_9334,N_9483);
nand U10619 (N_10619,N_9468,N_9048);
nor U10620 (N_10620,N_9591,N_9093);
or U10621 (N_10621,N_9722,N_9526);
or U10622 (N_10622,N_9619,N_9169);
and U10623 (N_10623,N_9676,N_9253);
nand U10624 (N_10624,N_9970,N_9672);
nor U10625 (N_10625,N_9212,N_9987);
and U10626 (N_10626,N_9651,N_9274);
or U10627 (N_10627,N_9938,N_9690);
or U10628 (N_10628,N_9241,N_9512);
or U10629 (N_10629,N_9324,N_9058);
nand U10630 (N_10630,N_9695,N_9939);
nor U10631 (N_10631,N_9866,N_9964);
nand U10632 (N_10632,N_9650,N_9338);
and U10633 (N_10633,N_9065,N_9948);
or U10634 (N_10634,N_9085,N_9459);
and U10635 (N_10635,N_9219,N_9533);
nor U10636 (N_10636,N_9924,N_9442);
or U10637 (N_10637,N_9657,N_9455);
nand U10638 (N_10638,N_9853,N_9681);
xor U10639 (N_10639,N_9781,N_9461);
nor U10640 (N_10640,N_9314,N_9697);
and U10641 (N_10641,N_9752,N_9734);
and U10642 (N_10642,N_9101,N_9831);
nand U10643 (N_10643,N_9118,N_9276);
nor U10644 (N_10644,N_9328,N_9829);
nor U10645 (N_10645,N_9686,N_9055);
xnor U10646 (N_10646,N_9495,N_9153);
nand U10647 (N_10647,N_9619,N_9932);
xnor U10648 (N_10648,N_9445,N_9871);
xor U10649 (N_10649,N_9473,N_9172);
xor U10650 (N_10650,N_9962,N_9381);
nor U10651 (N_10651,N_9060,N_9458);
or U10652 (N_10652,N_9040,N_9317);
nor U10653 (N_10653,N_9377,N_9208);
nor U10654 (N_10654,N_9947,N_9571);
nand U10655 (N_10655,N_9089,N_9110);
and U10656 (N_10656,N_9361,N_9309);
xnor U10657 (N_10657,N_9517,N_9861);
and U10658 (N_10658,N_9665,N_9531);
nor U10659 (N_10659,N_9302,N_9146);
nand U10660 (N_10660,N_9562,N_9666);
or U10661 (N_10661,N_9006,N_9941);
nand U10662 (N_10662,N_9179,N_9294);
nor U10663 (N_10663,N_9528,N_9239);
and U10664 (N_10664,N_9851,N_9887);
xnor U10665 (N_10665,N_9867,N_9976);
or U10666 (N_10666,N_9194,N_9260);
nor U10667 (N_10667,N_9310,N_9535);
xor U10668 (N_10668,N_9948,N_9309);
xor U10669 (N_10669,N_9336,N_9658);
xnor U10670 (N_10670,N_9081,N_9998);
or U10671 (N_10671,N_9728,N_9463);
and U10672 (N_10672,N_9896,N_9393);
or U10673 (N_10673,N_9168,N_9799);
nand U10674 (N_10674,N_9512,N_9217);
or U10675 (N_10675,N_9959,N_9467);
and U10676 (N_10676,N_9617,N_9057);
or U10677 (N_10677,N_9078,N_9136);
nand U10678 (N_10678,N_9101,N_9610);
or U10679 (N_10679,N_9745,N_9521);
and U10680 (N_10680,N_9089,N_9142);
nor U10681 (N_10681,N_9242,N_9547);
nand U10682 (N_10682,N_9636,N_9507);
xnor U10683 (N_10683,N_9489,N_9981);
nand U10684 (N_10684,N_9407,N_9065);
xnor U10685 (N_10685,N_9036,N_9940);
and U10686 (N_10686,N_9113,N_9390);
nand U10687 (N_10687,N_9611,N_9373);
nand U10688 (N_10688,N_9661,N_9503);
xor U10689 (N_10689,N_9777,N_9620);
xnor U10690 (N_10690,N_9143,N_9357);
and U10691 (N_10691,N_9280,N_9441);
and U10692 (N_10692,N_9826,N_9142);
xnor U10693 (N_10693,N_9818,N_9365);
and U10694 (N_10694,N_9447,N_9688);
nor U10695 (N_10695,N_9363,N_9525);
and U10696 (N_10696,N_9721,N_9027);
or U10697 (N_10697,N_9549,N_9371);
nor U10698 (N_10698,N_9039,N_9984);
xnor U10699 (N_10699,N_9230,N_9709);
and U10700 (N_10700,N_9667,N_9945);
xnor U10701 (N_10701,N_9392,N_9981);
nand U10702 (N_10702,N_9030,N_9126);
nand U10703 (N_10703,N_9017,N_9890);
and U10704 (N_10704,N_9593,N_9257);
or U10705 (N_10705,N_9721,N_9386);
and U10706 (N_10706,N_9963,N_9598);
and U10707 (N_10707,N_9386,N_9814);
and U10708 (N_10708,N_9918,N_9133);
and U10709 (N_10709,N_9113,N_9115);
nand U10710 (N_10710,N_9230,N_9060);
xnor U10711 (N_10711,N_9117,N_9501);
xnor U10712 (N_10712,N_9605,N_9024);
or U10713 (N_10713,N_9859,N_9924);
nand U10714 (N_10714,N_9900,N_9210);
or U10715 (N_10715,N_9624,N_9549);
or U10716 (N_10716,N_9412,N_9249);
and U10717 (N_10717,N_9268,N_9884);
xnor U10718 (N_10718,N_9852,N_9864);
nor U10719 (N_10719,N_9270,N_9717);
and U10720 (N_10720,N_9055,N_9409);
nor U10721 (N_10721,N_9344,N_9955);
xor U10722 (N_10722,N_9538,N_9358);
xor U10723 (N_10723,N_9759,N_9177);
or U10724 (N_10724,N_9751,N_9524);
nand U10725 (N_10725,N_9014,N_9635);
xnor U10726 (N_10726,N_9665,N_9296);
nor U10727 (N_10727,N_9464,N_9838);
and U10728 (N_10728,N_9933,N_9037);
or U10729 (N_10729,N_9697,N_9819);
or U10730 (N_10730,N_9697,N_9666);
or U10731 (N_10731,N_9283,N_9076);
nor U10732 (N_10732,N_9205,N_9704);
nor U10733 (N_10733,N_9102,N_9349);
or U10734 (N_10734,N_9481,N_9050);
nand U10735 (N_10735,N_9842,N_9916);
nand U10736 (N_10736,N_9328,N_9654);
xnor U10737 (N_10737,N_9391,N_9141);
nand U10738 (N_10738,N_9976,N_9537);
nor U10739 (N_10739,N_9974,N_9367);
and U10740 (N_10740,N_9911,N_9600);
or U10741 (N_10741,N_9953,N_9934);
nor U10742 (N_10742,N_9288,N_9392);
and U10743 (N_10743,N_9979,N_9010);
xor U10744 (N_10744,N_9370,N_9061);
xnor U10745 (N_10745,N_9393,N_9768);
or U10746 (N_10746,N_9320,N_9120);
nor U10747 (N_10747,N_9285,N_9847);
xnor U10748 (N_10748,N_9589,N_9999);
and U10749 (N_10749,N_9264,N_9912);
nand U10750 (N_10750,N_9080,N_9479);
nand U10751 (N_10751,N_9181,N_9973);
xnor U10752 (N_10752,N_9240,N_9375);
nand U10753 (N_10753,N_9210,N_9508);
xor U10754 (N_10754,N_9466,N_9762);
nor U10755 (N_10755,N_9279,N_9784);
xor U10756 (N_10756,N_9422,N_9679);
xnor U10757 (N_10757,N_9280,N_9955);
xor U10758 (N_10758,N_9489,N_9869);
or U10759 (N_10759,N_9574,N_9463);
or U10760 (N_10760,N_9434,N_9425);
nand U10761 (N_10761,N_9534,N_9978);
nor U10762 (N_10762,N_9212,N_9823);
nand U10763 (N_10763,N_9149,N_9110);
nor U10764 (N_10764,N_9644,N_9048);
and U10765 (N_10765,N_9558,N_9526);
and U10766 (N_10766,N_9046,N_9804);
nor U10767 (N_10767,N_9521,N_9847);
nand U10768 (N_10768,N_9945,N_9253);
and U10769 (N_10769,N_9223,N_9379);
and U10770 (N_10770,N_9881,N_9442);
and U10771 (N_10771,N_9218,N_9585);
xor U10772 (N_10772,N_9974,N_9514);
and U10773 (N_10773,N_9140,N_9997);
or U10774 (N_10774,N_9609,N_9187);
and U10775 (N_10775,N_9540,N_9894);
and U10776 (N_10776,N_9372,N_9517);
xor U10777 (N_10777,N_9459,N_9454);
nand U10778 (N_10778,N_9156,N_9973);
nand U10779 (N_10779,N_9418,N_9940);
and U10780 (N_10780,N_9069,N_9206);
xor U10781 (N_10781,N_9664,N_9823);
xor U10782 (N_10782,N_9679,N_9756);
or U10783 (N_10783,N_9694,N_9198);
nor U10784 (N_10784,N_9953,N_9134);
nand U10785 (N_10785,N_9658,N_9959);
and U10786 (N_10786,N_9203,N_9237);
nor U10787 (N_10787,N_9835,N_9506);
nor U10788 (N_10788,N_9177,N_9228);
xnor U10789 (N_10789,N_9845,N_9350);
xor U10790 (N_10790,N_9694,N_9672);
xnor U10791 (N_10791,N_9089,N_9337);
nor U10792 (N_10792,N_9994,N_9574);
or U10793 (N_10793,N_9441,N_9493);
nand U10794 (N_10794,N_9057,N_9469);
and U10795 (N_10795,N_9784,N_9723);
and U10796 (N_10796,N_9922,N_9747);
xor U10797 (N_10797,N_9540,N_9844);
xnor U10798 (N_10798,N_9162,N_9920);
or U10799 (N_10799,N_9138,N_9410);
xnor U10800 (N_10800,N_9750,N_9218);
and U10801 (N_10801,N_9855,N_9369);
nand U10802 (N_10802,N_9932,N_9880);
xor U10803 (N_10803,N_9878,N_9145);
or U10804 (N_10804,N_9735,N_9499);
xor U10805 (N_10805,N_9042,N_9258);
nor U10806 (N_10806,N_9855,N_9765);
or U10807 (N_10807,N_9159,N_9949);
xnor U10808 (N_10808,N_9620,N_9778);
nor U10809 (N_10809,N_9983,N_9315);
nand U10810 (N_10810,N_9950,N_9023);
nand U10811 (N_10811,N_9597,N_9190);
nor U10812 (N_10812,N_9408,N_9474);
xor U10813 (N_10813,N_9654,N_9889);
xnor U10814 (N_10814,N_9396,N_9125);
nand U10815 (N_10815,N_9995,N_9593);
and U10816 (N_10816,N_9834,N_9893);
nor U10817 (N_10817,N_9919,N_9075);
nor U10818 (N_10818,N_9544,N_9213);
and U10819 (N_10819,N_9923,N_9468);
and U10820 (N_10820,N_9596,N_9470);
nand U10821 (N_10821,N_9456,N_9152);
and U10822 (N_10822,N_9428,N_9965);
and U10823 (N_10823,N_9362,N_9625);
nand U10824 (N_10824,N_9322,N_9352);
xor U10825 (N_10825,N_9190,N_9132);
nor U10826 (N_10826,N_9416,N_9156);
xor U10827 (N_10827,N_9481,N_9396);
and U10828 (N_10828,N_9633,N_9493);
nor U10829 (N_10829,N_9504,N_9076);
or U10830 (N_10830,N_9878,N_9002);
or U10831 (N_10831,N_9613,N_9336);
xor U10832 (N_10832,N_9007,N_9549);
nand U10833 (N_10833,N_9522,N_9293);
nor U10834 (N_10834,N_9880,N_9939);
and U10835 (N_10835,N_9334,N_9181);
nand U10836 (N_10836,N_9027,N_9575);
and U10837 (N_10837,N_9168,N_9462);
nand U10838 (N_10838,N_9215,N_9944);
nor U10839 (N_10839,N_9892,N_9179);
or U10840 (N_10840,N_9245,N_9986);
nand U10841 (N_10841,N_9660,N_9400);
nand U10842 (N_10842,N_9963,N_9405);
xor U10843 (N_10843,N_9423,N_9454);
nor U10844 (N_10844,N_9634,N_9991);
nand U10845 (N_10845,N_9485,N_9108);
nor U10846 (N_10846,N_9182,N_9515);
nor U10847 (N_10847,N_9532,N_9039);
xnor U10848 (N_10848,N_9482,N_9316);
nor U10849 (N_10849,N_9191,N_9738);
nand U10850 (N_10850,N_9686,N_9810);
xnor U10851 (N_10851,N_9616,N_9750);
and U10852 (N_10852,N_9754,N_9576);
nand U10853 (N_10853,N_9463,N_9106);
nand U10854 (N_10854,N_9570,N_9818);
xor U10855 (N_10855,N_9197,N_9857);
nor U10856 (N_10856,N_9083,N_9248);
and U10857 (N_10857,N_9137,N_9389);
nor U10858 (N_10858,N_9025,N_9706);
xor U10859 (N_10859,N_9541,N_9228);
xnor U10860 (N_10860,N_9305,N_9611);
nand U10861 (N_10861,N_9733,N_9069);
and U10862 (N_10862,N_9932,N_9645);
nor U10863 (N_10863,N_9431,N_9080);
nor U10864 (N_10864,N_9272,N_9525);
nor U10865 (N_10865,N_9931,N_9140);
nor U10866 (N_10866,N_9703,N_9143);
and U10867 (N_10867,N_9236,N_9528);
and U10868 (N_10868,N_9296,N_9977);
or U10869 (N_10869,N_9764,N_9791);
or U10870 (N_10870,N_9233,N_9727);
or U10871 (N_10871,N_9138,N_9128);
and U10872 (N_10872,N_9532,N_9819);
or U10873 (N_10873,N_9051,N_9744);
nor U10874 (N_10874,N_9885,N_9051);
xnor U10875 (N_10875,N_9486,N_9225);
nor U10876 (N_10876,N_9264,N_9097);
xnor U10877 (N_10877,N_9889,N_9852);
and U10878 (N_10878,N_9591,N_9844);
nor U10879 (N_10879,N_9804,N_9978);
and U10880 (N_10880,N_9565,N_9827);
nor U10881 (N_10881,N_9331,N_9949);
xnor U10882 (N_10882,N_9871,N_9607);
nor U10883 (N_10883,N_9046,N_9619);
nand U10884 (N_10884,N_9206,N_9718);
and U10885 (N_10885,N_9487,N_9120);
nor U10886 (N_10886,N_9261,N_9172);
xor U10887 (N_10887,N_9472,N_9608);
nor U10888 (N_10888,N_9028,N_9042);
xor U10889 (N_10889,N_9162,N_9090);
and U10890 (N_10890,N_9610,N_9070);
and U10891 (N_10891,N_9925,N_9469);
nand U10892 (N_10892,N_9762,N_9515);
nand U10893 (N_10893,N_9545,N_9179);
or U10894 (N_10894,N_9214,N_9015);
nor U10895 (N_10895,N_9898,N_9078);
or U10896 (N_10896,N_9417,N_9312);
nand U10897 (N_10897,N_9192,N_9877);
nand U10898 (N_10898,N_9286,N_9352);
nor U10899 (N_10899,N_9542,N_9661);
nor U10900 (N_10900,N_9816,N_9894);
and U10901 (N_10901,N_9439,N_9598);
nor U10902 (N_10902,N_9771,N_9224);
and U10903 (N_10903,N_9191,N_9089);
or U10904 (N_10904,N_9213,N_9060);
and U10905 (N_10905,N_9193,N_9992);
or U10906 (N_10906,N_9291,N_9339);
nor U10907 (N_10907,N_9257,N_9712);
nor U10908 (N_10908,N_9560,N_9029);
xnor U10909 (N_10909,N_9172,N_9415);
xnor U10910 (N_10910,N_9926,N_9149);
nand U10911 (N_10911,N_9473,N_9887);
nand U10912 (N_10912,N_9067,N_9914);
nor U10913 (N_10913,N_9411,N_9927);
and U10914 (N_10914,N_9604,N_9174);
or U10915 (N_10915,N_9477,N_9787);
and U10916 (N_10916,N_9820,N_9267);
or U10917 (N_10917,N_9699,N_9915);
xnor U10918 (N_10918,N_9954,N_9220);
and U10919 (N_10919,N_9588,N_9913);
and U10920 (N_10920,N_9549,N_9965);
nand U10921 (N_10921,N_9199,N_9665);
or U10922 (N_10922,N_9972,N_9693);
nand U10923 (N_10923,N_9300,N_9569);
or U10924 (N_10924,N_9459,N_9724);
and U10925 (N_10925,N_9382,N_9942);
or U10926 (N_10926,N_9588,N_9902);
and U10927 (N_10927,N_9337,N_9830);
or U10928 (N_10928,N_9142,N_9081);
xor U10929 (N_10929,N_9888,N_9850);
or U10930 (N_10930,N_9373,N_9681);
nand U10931 (N_10931,N_9855,N_9208);
and U10932 (N_10932,N_9637,N_9588);
nor U10933 (N_10933,N_9379,N_9247);
and U10934 (N_10934,N_9530,N_9938);
nand U10935 (N_10935,N_9326,N_9165);
xnor U10936 (N_10936,N_9809,N_9261);
nand U10937 (N_10937,N_9914,N_9804);
nand U10938 (N_10938,N_9588,N_9904);
or U10939 (N_10939,N_9556,N_9798);
nor U10940 (N_10940,N_9133,N_9135);
nand U10941 (N_10941,N_9761,N_9575);
nor U10942 (N_10942,N_9905,N_9696);
nand U10943 (N_10943,N_9011,N_9307);
nor U10944 (N_10944,N_9661,N_9841);
nand U10945 (N_10945,N_9148,N_9323);
or U10946 (N_10946,N_9966,N_9714);
and U10947 (N_10947,N_9557,N_9198);
nand U10948 (N_10948,N_9531,N_9449);
and U10949 (N_10949,N_9145,N_9731);
or U10950 (N_10950,N_9609,N_9255);
or U10951 (N_10951,N_9624,N_9036);
nand U10952 (N_10952,N_9550,N_9962);
or U10953 (N_10953,N_9475,N_9694);
or U10954 (N_10954,N_9157,N_9476);
or U10955 (N_10955,N_9581,N_9790);
and U10956 (N_10956,N_9116,N_9382);
or U10957 (N_10957,N_9058,N_9507);
nor U10958 (N_10958,N_9495,N_9140);
and U10959 (N_10959,N_9894,N_9950);
nor U10960 (N_10960,N_9092,N_9369);
and U10961 (N_10961,N_9024,N_9051);
nor U10962 (N_10962,N_9290,N_9277);
xnor U10963 (N_10963,N_9044,N_9868);
nor U10964 (N_10964,N_9629,N_9627);
xor U10965 (N_10965,N_9927,N_9409);
or U10966 (N_10966,N_9409,N_9725);
and U10967 (N_10967,N_9915,N_9402);
and U10968 (N_10968,N_9678,N_9105);
or U10969 (N_10969,N_9546,N_9578);
or U10970 (N_10970,N_9516,N_9567);
nor U10971 (N_10971,N_9771,N_9384);
xor U10972 (N_10972,N_9460,N_9878);
or U10973 (N_10973,N_9756,N_9252);
or U10974 (N_10974,N_9197,N_9598);
or U10975 (N_10975,N_9777,N_9711);
nand U10976 (N_10976,N_9315,N_9938);
and U10977 (N_10977,N_9504,N_9141);
and U10978 (N_10978,N_9192,N_9888);
and U10979 (N_10979,N_9153,N_9183);
xor U10980 (N_10980,N_9879,N_9818);
and U10981 (N_10981,N_9702,N_9272);
nor U10982 (N_10982,N_9990,N_9257);
xnor U10983 (N_10983,N_9554,N_9846);
and U10984 (N_10984,N_9465,N_9502);
or U10985 (N_10985,N_9786,N_9884);
nor U10986 (N_10986,N_9340,N_9157);
nand U10987 (N_10987,N_9944,N_9087);
nor U10988 (N_10988,N_9991,N_9563);
or U10989 (N_10989,N_9293,N_9033);
and U10990 (N_10990,N_9952,N_9002);
or U10991 (N_10991,N_9704,N_9838);
and U10992 (N_10992,N_9632,N_9092);
and U10993 (N_10993,N_9832,N_9896);
xor U10994 (N_10994,N_9559,N_9072);
and U10995 (N_10995,N_9577,N_9608);
nand U10996 (N_10996,N_9120,N_9425);
and U10997 (N_10997,N_9119,N_9612);
xnor U10998 (N_10998,N_9848,N_9115);
or U10999 (N_10999,N_9856,N_9288);
nor U11000 (N_11000,N_10372,N_10055);
or U11001 (N_11001,N_10200,N_10538);
nand U11002 (N_11002,N_10642,N_10711);
nand U11003 (N_11003,N_10744,N_10277);
nand U11004 (N_11004,N_10085,N_10409);
nand U11005 (N_11005,N_10646,N_10887);
or U11006 (N_11006,N_10480,N_10197);
nand U11007 (N_11007,N_10985,N_10591);
and U11008 (N_11008,N_10247,N_10975);
and U11009 (N_11009,N_10885,N_10267);
nor U11010 (N_11010,N_10496,N_10999);
or U11011 (N_11011,N_10012,N_10500);
xnor U11012 (N_11012,N_10378,N_10922);
xnor U11013 (N_11013,N_10023,N_10196);
xor U11014 (N_11014,N_10424,N_10433);
nand U11015 (N_11015,N_10049,N_10075);
nand U11016 (N_11016,N_10040,N_10261);
xnor U11017 (N_11017,N_10881,N_10849);
xor U11018 (N_11018,N_10166,N_10319);
and U11019 (N_11019,N_10737,N_10215);
nor U11020 (N_11020,N_10537,N_10921);
nor U11021 (N_11021,N_10305,N_10276);
and U11022 (N_11022,N_10046,N_10919);
or U11023 (N_11023,N_10440,N_10416);
nor U11024 (N_11024,N_10381,N_10489);
nor U11025 (N_11025,N_10414,N_10858);
and U11026 (N_11026,N_10723,N_10769);
xor U11027 (N_11027,N_10264,N_10229);
xor U11028 (N_11028,N_10393,N_10340);
xnor U11029 (N_11029,N_10343,N_10253);
nand U11030 (N_11030,N_10826,N_10127);
and U11031 (N_11031,N_10725,N_10084);
xor U11032 (N_11032,N_10133,N_10132);
or U11033 (N_11033,N_10479,N_10525);
xnor U11034 (N_11034,N_10861,N_10526);
nand U11035 (N_11035,N_10336,N_10158);
xor U11036 (N_11036,N_10007,N_10643);
nor U11037 (N_11037,N_10603,N_10659);
or U11038 (N_11038,N_10289,N_10466);
nor U11039 (N_11039,N_10705,N_10086);
or U11040 (N_11040,N_10565,N_10491);
nor U11041 (N_11041,N_10545,N_10419);
nor U11042 (N_11042,N_10557,N_10153);
nor U11043 (N_11043,N_10771,N_10421);
nand U11044 (N_11044,N_10481,N_10806);
nor U11045 (N_11045,N_10331,N_10349);
xor U11046 (N_11046,N_10297,N_10831);
nor U11047 (N_11047,N_10955,N_10426);
and U11048 (N_11048,N_10572,N_10687);
or U11049 (N_11049,N_10190,N_10191);
or U11050 (N_11050,N_10663,N_10815);
nand U11051 (N_11051,N_10594,N_10917);
nor U11052 (N_11052,N_10819,N_10697);
nand U11053 (N_11053,N_10209,N_10904);
nor U11054 (N_11054,N_10674,N_10620);
nand U11055 (N_11055,N_10753,N_10972);
or U11056 (N_11056,N_10380,N_10540);
and U11057 (N_11057,N_10351,N_10784);
and U11058 (N_11058,N_10874,N_10829);
and U11059 (N_11059,N_10721,N_10314);
nor U11060 (N_11060,N_10788,N_10329);
nand U11061 (N_11061,N_10475,N_10022);
nand U11062 (N_11062,N_10997,N_10776);
or U11063 (N_11063,N_10484,N_10050);
nand U11064 (N_11064,N_10004,N_10929);
xor U11065 (N_11065,N_10296,N_10089);
and U11066 (N_11066,N_10931,N_10309);
nor U11067 (N_11067,N_10518,N_10151);
or U11068 (N_11068,N_10768,N_10162);
nand U11069 (N_11069,N_10810,N_10833);
and U11070 (N_11070,N_10080,N_10606);
or U11071 (N_11071,N_10015,N_10945);
nor U11072 (N_11072,N_10923,N_10602);
or U11073 (N_11073,N_10661,N_10676);
nor U11074 (N_11074,N_10495,N_10649);
nor U11075 (N_11075,N_10368,N_10119);
nor U11076 (N_11076,N_10240,N_10412);
or U11077 (N_11077,N_10008,N_10338);
xor U11078 (N_11078,N_10513,N_10939);
nor U11079 (N_11079,N_10730,N_10498);
nand U11080 (N_11080,N_10911,N_10681);
nand U11081 (N_11081,N_10662,N_10246);
xnor U11082 (N_11082,N_10516,N_10515);
nor U11083 (N_11083,N_10154,N_10384);
and U11084 (N_11084,N_10288,N_10183);
or U11085 (N_11085,N_10003,N_10712);
xor U11086 (N_11086,N_10511,N_10417);
nand U11087 (N_11087,N_10088,N_10250);
nor U11088 (N_11088,N_10601,N_10316);
xor U11089 (N_11089,N_10589,N_10069);
nor U11090 (N_11090,N_10122,N_10952);
nor U11091 (N_11091,N_10038,N_10110);
nand U11092 (N_11092,N_10255,N_10212);
and U11093 (N_11093,N_10057,N_10727);
xor U11094 (N_11094,N_10477,N_10766);
nand U11095 (N_11095,N_10418,N_10241);
nand U11096 (N_11096,N_10024,N_10494);
and U11097 (N_11097,N_10270,N_10555);
xnor U11098 (N_11098,N_10666,N_10065);
nor U11099 (N_11099,N_10944,N_10686);
xnor U11100 (N_11100,N_10556,N_10265);
and U11101 (N_11101,N_10560,N_10285);
or U11102 (N_11102,N_10425,N_10693);
or U11103 (N_11103,N_10031,N_10678);
nand U11104 (N_11104,N_10454,N_10840);
nor U11105 (N_11105,N_10871,N_10371);
xor U11106 (N_11106,N_10587,N_10823);
and U11107 (N_11107,N_10432,N_10415);
nor U11108 (N_11108,N_10506,N_10016);
xor U11109 (N_11109,N_10505,N_10547);
xor U11110 (N_11110,N_10868,N_10959);
xnor U11111 (N_11111,N_10568,N_10120);
or U11112 (N_11112,N_10444,N_10449);
and U11113 (N_11113,N_10562,N_10521);
nor U11114 (N_11114,N_10567,N_10395);
xnor U11115 (N_11115,N_10213,N_10458);
xnor U11116 (N_11116,N_10675,N_10585);
nand U11117 (N_11117,N_10825,N_10383);
nor U11118 (N_11118,N_10740,N_10751);
nor U11119 (N_11119,N_10943,N_10244);
and U11120 (N_11120,N_10897,N_10357);
and U11121 (N_11121,N_10018,N_10696);
nand U11122 (N_11122,N_10364,N_10226);
nor U11123 (N_11123,N_10204,N_10382);
xor U11124 (N_11124,N_10118,N_10108);
nor U11125 (N_11125,N_10683,N_10954);
nor U11126 (N_11126,N_10344,N_10062);
and U11127 (N_11127,N_10106,N_10987);
xor U11128 (N_11128,N_10534,N_10875);
nor U11129 (N_11129,N_10558,N_10205);
nand U11130 (N_11130,N_10413,N_10933);
and U11131 (N_11131,N_10081,N_10934);
nor U11132 (N_11132,N_10655,N_10422);
nand U11133 (N_11133,N_10445,N_10463);
and U11134 (N_11134,N_10629,N_10105);
nand U11135 (N_11135,N_10889,N_10907);
and U11136 (N_11136,N_10116,N_10455);
and U11137 (N_11137,N_10682,N_10199);
and U11138 (N_11138,N_10307,N_10656);
xor U11139 (N_11139,N_10546,N_10541);
nor U11140 (N_11140,N_10530,N_10114);
and U11141 (N_11141,N_10953,N_10844);
and U11142 (N_11142,N_10891,N_10869);
nand U11143 (N_11143,N_10836,N_10434);
and U11144 (N_11144,N_10320,N_10017);
nand U11145 (N_11145,N_10402,N_10410);
xnor U11146 (N_11146,N_10045,N_10070);
and U11147 (N_11147,N_10739,N_10803);
xor U11148 (N_11148,N_10715,N_10724);
nor U11149 (N_11149,N_10877,N_10925);
and U11150 (N_11150,N_10779,N_10439);
nand U11151 (N_11151,N_10400,N_10848);
or U11152 (N_11152,N_10369,N_10978);
nor U11153 (N_11153,N_10300,N_10146);
nand U11154 (N_11154,N_10963,N_10326);
or U11155 (N_11155,N_10828,N_10878);
or U11156 (N_11156,N_10935,N_10860);
or U11157 (N_11157,N_10783,N_10755);
nor U11158 (N_11158,N_10450,N_10210);
nand U11159 (N_11159,N_10388,N_10654);
nand U11160 (N_11160,N_10233,N_10128);
xnor U11161 (N_11161,N_10834,N_10202);
or U11162 (N_11162,N_10614,N_10653);
or U11163 (N_11163,N_10669,N_10076);
or U11164 (N_11164,N_10136,N_10778);
or U11165 (N_11165,N_10198,N_10960);
nand U11166 (N_11166,N_10685,N_10028);
xor U11167 (N_11167,N_10671,N_10266);
nor U11168 (N_11168,N_10956,N_10161);
nor U11169 (N_11169,N_10983,N_10262);
or U11170 (N_11170,N_10615,N_10820);
and U11171 (N_11171,N_10613,N_10286);
nand U11172 (N_11172,N_10798,N_10651);
nand U11173 (N_11173,N_10670,N_10673);
or U11174 (N_11174,N_10301,N_10667);
nor U11175 (N_11175,N_10025,N_10068);
nand U11176 (N_11176,N_10504,N_10961);
xor U11177 (N_11177,N_10841,N_10353);
and U11178 (N_11178,N_10358,N_10736);
or U11179 (N_11179,N_10272,N_10814);
nor U11180 (N_11180,N_10313,N_10908);
nand U11181 (N_11181,N_10989,N_10501);
nor U11182 (N_11182,N_10217,N_10630);
nor U11183 (N_11183,N_10333,N_10002);
and U11184 (N_11184,N_10280,N_10957);
nor U11185 (N_11185,N_10838,N_10706);
nor U11186 (N_11186,N_10657,N_10188);
nor U11187 (N_11187,N_10583,N_10124);
nor U11188 (N_11188,N_10728,N_10103);
nor U11189 (N_11189,N_10011,N_10808);
or U11190 (N_11190,N_10531,N_10271);
nand U11191 (N_11191,N_10293,N_10150);
nor U11192 (N_11192,N_10125,N_10554);
xor U11193 (N_11193,N_10453,N_10872);
xor U11194 (N_11194,N_10647,N_10323);
nand U11195 (N_11195,N_10832,N_10180);
nor U11196 (N_11196,N_10291,N_10795);
or U11197 (N_11197,N_10632,N_10472);
and U11198 (N_11198,N_10822,N_10208);
and U11199 (N_11199,N_10184,N_10936);
xor U11200 (N_11200,N_10436,N_10248);
and U11201 (N_11201,N_10139,N_10302);
nand U11202 (N_11202,N_10970,N_10325);
nor U11203 (N_11203,N_10578,N_10112);
or U11204 (N_11204,N_10342,N_10221);
xnor U11205 (N_11205,N_10430,N_10470);
xor U11206 (N_11206,N_10104,N_10734);
nand U11207 (N_11207,N_10030,N_10093);
xor U11208 (N_11208,N_10401,N_10299);
nor U11209 (N_11209,N_10236,N_10597);
and U11210 (N_11210,N_10257,N_10490);
xor U11211 (N_11211,N_10181,N_10054);
nand U11212 (N_11212,N_10042,N_10273);
nor U11213 (N_11213,N_10051,N_10990);
nor U11214 (N_11214,N_10765,N_10846);
and U11215 (N_11215,N_10249,N_10026);
xor U11216 (N_11216,N_10864,N_10126);
and U11217 (N_11217,N_10910,N_10884);
xnor U11218 (N_11218,N_10702,N_10767);
or U11219 (N_11219,N_10304,N_10748);
nand U11220 (N_11220,N_10256,N_10259);
xnor U11221 (N_11221,N_10187,N_10169);
xnor U11222 (N_11222,N_10637,N_10461);
nor U11223 (N_11223,N_10738,N_10993);
nand U11224 (N_11224,N_10636,N_10720);
xor U11225 (N_11225,N_10906,N_10476);
xnor U11226 (N_11226,N_10163,N_10387);
or U11227 (N_11227,N_10034,N_10624);
xnor U11228 (N_11228,N_10497,N_10001);
nand U11229 (N_11229,N_10576,N_10269);
nand U11230 (N_11230,N_10242,N_10660);
xor U11231 (N_11231,N_10763,N_10053);
nor U11232 (N_11232,N_10281,N_10352);
and U11233 (N_11233,N_10980,N_10679);
or U11234 (N_11234,N_10992,N_10579);
xor U11235 (N_11235,N_10334,N_10438);
and U11236 (N_11236,N_10950,N_10695);
nor U11237 (N_11237,N_10524,N_10855);
xor U11238 (N_11238,N_10507,N_10842);
and U11239 (N_11239,N_10648,N_10274);
or U11240 (N_11240,N_10295,N_10598);
xnor U11241 (N_11241,N_10283,N_10621);
nor U11242 (N_11242,N_10969,N_10502);
nor U11243 (N_11243,N_10386,N_10618);
or U11244 (N_11244,N_10684,N_10837);
or U11245 (N_11245,N_10172,N_10867);
xor U11246 (N_11246,N_10292,N_10764);
nand U11247 (N_11247,N_10394,N_10408);
nand U11248 (N_11248,N_10805,N_10704);
nor U11249 (N_11249,N_10596,N_10619);
nand U11250 (N_11250,N_10566,N_10471);
nand U11251 (N_11251,N_10926,N_10830);
xnor U11252 (N_11252,N_10616,N_10611);
or U11253 (N_11253,N_10856,N_10486);
nor U11254 (N_11254,N_10775,N_10014);
or U11255 (N_11255,N_10982,N_10853);
or U11256 (N_11256,N_10117,N_10130);
nand U11257 (N_11257,N_10174,N_10584);
or U11258 (N_11258,N_10577,N_10701);
xor U11259 (N_11259,N_10707,N_10224);
and U11260 (N_11260,N_10799,N_10423);
and U11261 (N_11261,N_10781,N_10123);
or U11262 (N_11262,N_10474,N_10813);
xor U11263 (N_11263,N_10612,N_10882);
or U11264 (N_11264,N_10404,N_10581);
xor U11265 (N_11265,N_10290,N_10569);
or U11266 (N_11266,N_10716,N_10156);
or U11267 (N_11267,N_10145,N_10389);
or U11268 (N_11268,N_10812,N_10090);
or U11269 (N_11269,N_10341,N_10664);
nand U11270 (N_11270,N_10177,N_10376);
nor U11271 (N_11271,N_10355,N_10318);
nand U11272 (N_11272,N_10609,N_10228);
xnor U11273 (N_11273,N_10852,N_10152);
nor U11274 (N_11274,N_10965,N_10564);
nand U11275 (N_11275,N_10189,N_10726);
or U11276 (N_11276,N_10580,N_10735);
nor U11277 (N_11277,N_10998,N_10311);
nand U11278 (N_11278,N_10732,N_10098);
xor U11279 (N_11279,N_10843,N_10227);
xnor U11280 (N_11280,N_10148,N_10942);
and U11281 (N_11281,N_10006,N_10167);
nor U11282 (N_11282,N_10047,N_10550);
and U11283 (N_11283,N_10665,N_10742);
nand U11284 (N_11284,N_10168,N_10220);
or U11285 (N_11285,N_10039,N_10279);
xor U11286 (N_11286,N_10041,N_10809);
nor U11287 (N_11287,N_10312,N_10315);
and U11288 (N_11288,N_10374,N_10429);
nand U11289 (N_11289,N_10464,N_10689);
or U11290 (N_11290,N_10958,N_10443);
nor U11291 (N_11291,N_10298,N_10232);
nor U11292 (N_11292,N_10178,N_10442);
nor U11293 (N_11293,N_10317,N_10811);
xnor U11294 (N_11294,N_10694,N_10032);
or U11295 (N_11295,N_10033,N_10575);
xor U11296 (N_11296,N_10794,N_10847);
nand U11297 (N_11297,N_10573,N_10121);
and U11298 (N_11298,N_10437,N_10308);
nand U11299 (N_11299,N_10517,N_10390);
nand U11300 (N_11300,N_10797,N_10976);
or U11301 (N_11301,N_10078,N_10745);
and U11302 (N_11302,N_10356,N_10892);
or U11303 (N_11303,N_10071,N_10010);
nand U11304 (N_11304,N_10633,N_10157);
and U11305 (N_11305,N_10222,N_10483);
xor U11306 (N_11306,N_10774,N_10456);
or U11307 (N_11307,N_10348,N_10064);
or U11308 (N_11308,N_10100,N_10551);
xnor U11309 (N_11309,N_10918,N_10160);
nor U11310 (N_11310,N_10758,N_10595);
nand U11311 (N_11311,N_10691,N_10337);
nand U11312 (N_11312,N_10129,N_10435);
nor U11313 (N_11313,N_10717,N_10462);
or U11314 (N_11314,N_10218,N_10321);
or U11315 (N_11315,N_10802,N_10863);
nor U11316 (N_11316,N_10235,N_10137);
nand U11317 (N_11317,N_10941,N_10817);
or U11318 (N_11318,N_10328,N_10780);
xor U11319 (N_11319,N_10592,N_10332);
nand U11320 (N_11320,N_10539,N_10967);
xor U11321 (N_11321,N_10680,N_10060);
and U11322 (N_11322,N_10399,N_10593);
and U11323 (N_11323,N_10544,N_10346);
nand U11324 (N_11324,N_10379,N_10009);
xor U11325 (N_11325,N_10913,N_10971);
xnor U11326 (N_11326,N_10747,N_10036);
nand U11327 (N_11327,N_10020,N_10762);
and U11328 (N_11328,N_10512,N_10995);
nor U11329 (N_11329,N_10625,N_10968);
and U11330 (N_11330,N_10005,N_10063);
or U11331 (N_11331,N_10893,N_10948);
and U11332 (N_11332,N_10741,N_10243);
nor U11333 (N_11333,N_10252,N_10446);
and U11334 (N_11334,N_10949,N_10786);
xor U11335 (N_11335,N_10549,N_10688);
or U11336 (N_11336,N_10839,N_10079);
xnor U11337 (N_11337,N_10900,N_10082);
nand U11338 (N_11338,N_10147,N_10940);
or U11339 (N_11339,N_10928,N_10251);
or U11340 (N_11340,N_10193,N_10396);
and U11341 (N_11341,N_10254,N_10772);
and U11342 (N_11342,N_10225,N_10529);
nor U11343 (N_11343,N_10912,N_10807);
xnor U11344 (N_11344,N_10428,N_10310);
or U11345 (N_11345,N_10658,N_10542);
or U11346 (N_11346,N_10219,N_10330);
nor U11347 (N_11347,N_10986,N_10898);
nor U11348 (N_11348,N_10827,N_10909);
nand U11349 (N_11349,N_10520,N_10377);
xnor U11350 (N_11350,N_10991,N_10974);
nand U11351 (N_11351,N_10185,N_10865);
xnor U11352 (N_11352,N_10700,N_10173);
and U11353 (N_11353,N_10508,N_10223);
nand U11354 (N_11354,N_10142,N_10303);
and U11355 (N_11355,N_10306,N_10574);
or U11356 (N_11356,N_10485,N_10366);
or U11357 (N_11357,N_10759,N_10708);
nand U11358 (N_11358,N_10375,N_10533);
xnor U11359 (N_11359,N_10370,N_10835);
nand U11360 (N_11360,N_10092,N_10713);
nand U11361 (N_11361,N_10548,N_10981);
nor U11362 (N_11362,N_10465,N_10522);
xor U11363 (N_11363,N_10690,N_10354);
nand U11364 (N_11364,N_10622,N_10237);
nor U11365 (N_11365,N_10149,N_10095);
nor U11366 (N_11366,N_10626,N_10203);
or U11367 (N_11367,N_10013,N_10818);
xor U11368 (N_11368,N_10373,N_10552);
nor U11369 (N_11369,N_10607,N_10886);
or U11370 (N_11370,N_10350,N_10920);
nor U11371 (N_11371,N_10785,N_10043);
nand U11372 (N_11372,N_10631,N_10140);
nor U11373 (N_11373,N_10111,N_10644);
nand U11374 (N_11374,N_10211,N_10359);
nor U11375 (N_11375,N_10192,N_10851);
nand U11376 (N_11376,N_10527,N_10322);
nor U11377 (N_11377,N_10182,N_10457);
nand U11378 (N_11378,N_10155,N_10946);
nor U11379 (N_11379,N_10459,N_10962);
and U11380 (N_11380,N_10916,N_10469);
and U11381 (N_11381,N_10391,N_10231);
xor U11382 (N_11382,N_10234,N_10411);
nor U11383 (N_11383,N_10294,N_10857);
nand U11384 (N_11384,N_10278,N_10493);
nor U11385 (N_11385,N_10452,N_10873);
xnor U11386 (N_11386,N_10087,N_10789);
and U11387 (N_11387,N_10499,N_10559);
nor U11388 (N_11388,N_10067,N_10195);
nand U11389 (N_11389,N_10441,N_10048);
xnor U11390 (N_11390,N_10509,N_10473);
nand U11391 (N_11391,N_10915,N_10627);
nor U11392 (N_11392,N_10510,N_10268);
nand U11393 (N_11393,N_10335,N_10131);
nor U11394 (N_11394,N_10536,N_10214);
nor U11395 (N_11395,N_10097,N_10107);
xnor U11396 (N_11396,N_10339,N_10777);
and U11397 (N_11397,N_10362,N_10135);
xnor U11398 (N_11398,N_10608,N_10570);
nor U11399 (N_11399,N_10756,N_10914);
xnor U11400 (N_11400,N_10096,N_10757);
xor U11401 (N_11401,N_10927,N_10821);
nor U11402 (N_11402,N_10029,N_10719);
nor U11403 (N_11403,N_10845,N_10263);
or U11404 (N_11404,N_10360,N_10239);
or U11405 (N_11405,N_10397,N_10553);
nor U11406 (N_11406,N_10134,N_10672);
nor U11407 (N_11407,N_10363,N_10590);
and U11408 (N_11408,N_10966,N_10588);
or U11409 (N_11409,N_10345,N_10487);
xnor U11410 (N_11410,N_10245,N_10791);
xor U11411 (N_11411,N_10731,N_10947);
nand U11412 (N_11412,N_10044,N_10407);
nor U11413 (N_11413,N_10870,N_10979);
nor U11414 (N_11414,N_10175,N_10770);
xor U11415 (N_11415,N_10027,N_10066);
nand U11416 (N_11416,N_10994,N_10101);
nand U11417 (N_11417,N_10634,N_10752);
nand U11418 (N_11418,N_10773,N_10523);
xor U11419 (N_11419,N_10447,N_10641);
and U11420 (N_11420,N_10144,N_10790);
or U11421 (N_11421,N_10094,N_10623);
xor U11422 (N_11422,N_10179,N_10021);
or U11423 (N_11423,N_10977,N_10468);
or U11424 (N_11424,N_10467,N_10733);
or U11425 (N_11425,N_10186,N_10932);
nor U11426 (N_11426,N_10938,N_10478);
and U11427 (N_11427,N_10398,N_10115);
and U11428 (N_11428,N_10061,N_10749);
nand U11429 (N_11429,N_10782,N_10514);
nand U11430 (N_11430,N_10746,N_10431);
xor U11431 (N_11431,N_10532,N_10102);
nor U11432 (N_11432,N_10862,N_10109);
nand U11433 (N_11433,N_10099,N_10937);
and U11434 (N_11434,N_10056,N_10652);
or U11435 (N_11435,N_10216,N_10543);
or U11436 (N_11436,N_10367,N_10492);
xor U11437 (N_11437,N_10924,N_10073);
and U11438 (N_11438,N_10638,N_10902);
or U11439 (N_11439,N_10159,N_10074);
xor U11440 (N_11440,N_10176,N_10037);
or U11441 (N_11441,N_10610,N_10035);
nand U11442 (N_11442,N_10899,N_10535);
nor U11443 (N_11443,N_10895,N_10405);
and U11444 (N_11444,N_10519,N_10901);
nand U11445 (N_11445,N_10793,N_10617);
nand U11446 (N_11446,N_10984,N_10668);
nor U11447 (N_11447,N_10692,N_10347);
xor U11448 (N_11448,N_10605,N_10528);
nand U11449 (N_11449,N_10052,N_10760);
xor U11450 (N_11450,N_10194,N_10019);
nor U11451 (N_11451,N_10365,N_10563);
nand U11452 (N_11452,N_10761,N_10604);
nand U11453 (N_11453,N_10427,N_10801);
xnor U11454 (N_11454,N_10930,N_10141);
nor U11455 (N_11455,N_10482,N_10287);
or U11456 (N_11456,N_10571,N_10385);
or U11457 (N_11457,N_10503,N_10628);
nor U11458 (N_11458,N_10677,N_10327);
xor U11459 (N_11459,N_10824,N_10894);
and U11460 (N_11460,N_10743,N_10600);
xnor U11461 (N_11461,N_10164,N_10171);
nor U11462 (N_11462,N_10206,N_10816);
xnor U11463 (N_11463,N_10792,N_10879);
nand U11464 (N_11464,N_10650,N_10905);
xnor U11465 (N_11465,N_10586,N_10361);
xor U11466 (N_11466,N_10903,N_10645);
and U11467 (N_11467,N_10896,N_10488);
and U11468 (N_11468,N_10640,N_10754);
xor U11469 (N_11469,N_10324,N_10714);
nor U11470 (N_11470,N_10170,N_10883);
nor U11471 (N_11471,N_10787,N_10561);
nand U11472 (N_11472,N_10072,N_10850);
xnor U11473 (N_11473,N_10996,N_10973);
nand U11474 (N_11474,N_10258,N_10890);
nand U11475 (N_11475,N_10091,N_10729);
xor U11476 (N_11476,N_10284,N_10207);
nor U11477 (N_11477,N_10639,N_10718);
and U11478 (N_11478,N_10710,N_10201);
or U11479 (N_11479,N_10699,N_10796);
or U11480 (N_11480,N_10635,N_10165);
and U11481 (N_11481,N_10951,N_10460);
or U11482 (N_11482,N_10750,N_10703);
xor U11483 (N_11483,N_10988,N_10238);
nor U11484 (N_11484,N_10866,N_10230);
nand U11485 (N_11485,N_10083,N_10582);
and U11486 (N_11486,N_10275,N_10854);
xor U11487 (N_11487,N_10406,N_10859);
and U11488 (N_11488,N_10000,N_10964);
xnor U11489 (N_11489,N_10888,N_10709);
and U11490 (N_11490,N_10113,N_10260);
xnor U11491 (N_11491,N_10448,N_10282);
nor U11492 (N_11492,N_10392,N_10804);
or U11493 (N_11493,N_10599,N_10420);
xnor U11494 (N_11494,N_10403,N_10059);
and U11495 (N_11495,N_10876,N_10722);
nand U11496 (N_11496,N_10077,N_10880);
and U11497 (N_11497,N_10143,N_10451);
nand U11498 (N_11498,N_10800,N_10698);
and U11499 (N_11499,N_10058,N_10138);
xnor U11500 (N_11500,N_10154,N_10846);
nand U11501 (N_11501,N_10147,N_10771);
and U11502 (N_11502,N_10746,N_10907);
or U11503 (N_11503,N_10859,N_10583);
xor U11504 (N_11504,N_10233,N_10365);
and U11505 (N_11505,N_10821,N_10836);
xor U11506 (N_11506,N_10182,N_10848);
nor U11507 (N_11507,N_10835,N_10542);
nor U11508 (N_11508,N_10338,N_10150);
or U11509 (N_11509,N_10413,N_10908);
or U11510 (N_11510,N_10576,N_10160);
nand U11511 (N_11511,N_10815,N_10366);
and U11512 (N_11512,N_10456,N_10155);
xnor U11513 (N_11513,N_10055,N_10188);
and U11514 (N_11514,N_10913,N_10352);
or U11515 (N_11515,N_10344,N_10503);
and U11516 (N_11516,N_10923,N_10649);
and U11517 (N_11517,N_10362,N_10523);
xnor U11518 (N_11518,N_10508,N_10248);
or U11519 (N_11519,N_10678,N_10624);
and U11520 (N_11520,N_10705,N_10959);
and U11521 (N_11521,N_10534,N_10500);
and U11522 (N_11522,N_10822,N_10919);
and U11523 (N_11523,N_10309,N_10365);
nand U11524 (N_11524,N_10907,N_10490);
nand U11525 (N_11525,N_10357,N_10422);
or U11526 (N_11526,N_10334,N_10824);
nor U11527 (N_11527,N_10090,N_10730);
nand U11528 (N_11528,N_10184,N_10149);
and U11529 (N_11529,N_10890,N_10769);
or U11530 (N_11530,N_10038,N_10387);
nor U11531 (N_11531,N_10831,N_10910);
nand U11532 (N_11532,N_10481,N_10024);
and U11533 (N_11533,N_10621,N_10001);
nand U11534 (N_11534,N_10255,N_10552);
xnor U11535 (N_11535,N_10276,N_10475);
and U11536 (N_11536,N_10934,N_10696);
nor U11537 (N_11537,N_10671,N_10073);
nand U11538 (N_11538,N_10650,N_10502);
nor U11539 (N_11539,N_10511,N_10819);
nor U11540 (N_11540,N_10903,N_10393);
nor U11541 (N_11541,N_10057,N_10080);
nand U11542 (N_11542,N_10581,N_10349);
xor U11543 (N_11543,N_10795,N_10257);
nor U11544 (N_11544,N_10654,N_10066);
and U11545 (N_11545,N_10915,N_10249);
or U11546 (N_11546,N_10915,N_10247);
nand U11547 (N_11547,N_10647,N_10893);
nand U11548 (N_11548,N_10186,N_10240);
or U11549 (N_11549,N_10963,N_10459);
and U11550 (N_11550,N_10337,N_10481);
nor U11551 (N_11551,N_10125,N_10596);
nor U11552 (N_11552,N_10237,N_10372);
nor U11553 (N_11553,N_10685,N_10090);
nor U11554 (N_11554,N_10033,N_10546);
or U11555 (N_11555,N_10343,N_10158);
or U11556 (N_11556,N_10099,N_10818);
nor U11557 (N_11557,N_10179,N_10602);
and U11558 (N_11558,N_10847,N_10730);
xnor U11559 (N_11559,N_10744,N_10350);
nand U11560 (N_11560,N_10834,N_10539);
nand U11561 (N_11561,N_10575,N_10302);
or U11562 (N_11562,N_10627,N_10223);
nor U11563 (N_11563,N_10568,N_10624);
nand U11564 (N_11564,N_10989,N_10239);
and U11565 (N_11565,N_10758,N_10975);
and U11566 (N_11566,N_10930,N_10628);
xnor U11567 (N_11567,N_10905,N_10355);
and U11568 (N_11568,N_10025,N_10474);
xor U11569 (N_11569,N_10141,N_10340);
nand U11570 (N_11570,N_10455,N_10267);
nand U11571 (N_11571,N_10991,N_10565);
xnor U11572 (N_11572,N_10734,N_10139);
xor U11573 (N_11573,N_10263,N_10999);
or U11574 (N_11574,N_10786,N_10579);
nor U11575 (N_11575,N_10701,N_10497);
nand U11576 (N_11576,N_10765,N_10637);
xnor U11577 (N_11577,N_10054,N_10604);
and U11578 (N_11578,N_10627,N_10819);
nand U11579 (N_11579,N_10162,N_10460);
nand U11580 (N_11580,N_10207,N_10019);
or U11581 (N_11581,N_10990,N_10281);
and U11582 (N_11582,N_10666,N_10529);
nand U11583 (N_11583,N_10386,N_10836);
nor U11584 (N_11584,N_10560,N_10916);
nand U11585 (N_11585,N_10813,N_10825);
xor U11586 (N_11586,N_10276,N_10984);
nor U11587 (N_11587,N_10872,N_10966);
xor U11588 (N_11588,N_10337,N_10686);
nand U11589 (N_11589,N_10524,N_10910);
and U11590 (N_11590,N_10119,N_10128);
nor U11591 (N_11591,N_10481,N_10452);
nor U11592 (N_11592,N_10964,N_10821);
nor U11593 (N_11593,N_10969,N_10757);
nor U11594 (N_11594,N_10968,N_10063);
nand U11595 (N_11595,N_10519,N_10272);
and U11596 (N_11596,N_10492,N_10310);
nor U11597 (N_11597,N_10771,N_10319);
or U11598 (N_11598,N_10278,N_10893);
nor U11599 (N_11599,N_10724,N_10183);
xor U11600 (N_11600,N_10750,N_10670);
nor U11601 (N_11601,N_10853,N_10829);
or U11602 (N_11602,N_10329,N_10542);
or U11603 (N_11603,N_10617,N_10561);
nor U11604 (N_11604,N_10596,N_10389);
or U11605 (N_11605,N_10437,N_10764);
or U11606 (N_11606,N_10896,N_10869);
or U11607 (N_11607,N_10027,N_10899);
nor U11608 (N_11608,N_10630,N_10754);
and U11609 (N_11609,N_10902,N_10466);
and U11610 (N_11610,N_10235,N_10287);
and U11611 (N_11611,N_10407,N_10218);
and U11612 (N_11612,N_10188,N_10374);
or U11613 (N_11613,N_10963,N_10846);
nand U11614 (N_11614,N_10330,N_10753);
xnor U11615 (N_11615,N_10198,N_10801);
and U11616 (N_11616,N_10815,N_10759);
and U11617 (N_11617,N_10963,N_10801);
or U11618 (N_11618,N_10164,N_10225);
or U11619 (N_11619,N_10446,N_10746);
or U11620 (N_11620,N_10110,N_10901);
nand U11621 (N_11621,N_10421,N_10640);
or U11622 (N_11622,N_10093,N_10724);
nor U11623 (N_11623,N_10061,N_10741);
nor U11624 (N_11624,N_10438,N_10097);
xor U11625 (N_11625,N_10087,N_10337);
nor U11626 (N_11626,N_10670,N_10156);
nand U11627 (N_11627,N_10319,N_10287);
and U11628 (N_11628,N_10961,N_10064);
xnor U11629 (N_11629,N_10130,N_10984);
nand U11630 (N_11630,N_10342,N_10922);
nor U11631 (N_11631,N_10832,N_10783);
and U11632 (N_11632,N_10428,N_10641);
nor U11633 (N_11633,N_10927,N_10764);
nor U11634 (N_11634,N_10966,N_10948);
nor U11635 (N_11635,N_10271,N_10968);
and U11636 (N_11636,N_10106,N_10017);
nor U11637 (N_11637,N_10173,N_10547);
or U11638 (N_11638,N_10960,N_10332);
and U11639 (N_11639,N_10868,N_10126);
or U11640 (N_11640,N_10578,N_10291);
and U11641 (N_11641,N_10953,N_10522);
and U11642 (N_11642,N_10575,N_10751);
nor U11643 (N_11643,N_10171,N_10218);
nor U11644 (N_11644,N_10994,N_10102);
or U11645 (N_11645,N_10103,N_10694);
nand U11646 (N_11646,N_10757,N_10440);
and U11647 (N_11647,N_10540,N_10161);
xnor U11648 (N_11648,N_10705,N_10988);
xnor U11649 (N_11649,N_10760,N_10677);
nand U11650 (N_11650,N_10261,N_10441);
nand U11651 (N_11651,N_10153,N_10861);
or U11652 (N_11652,N_10464,N_10316);
and U11653 (N_11653,N_10633,N_10253);
or U11654 (N_11654,N_10014,N_10799);
xnor U11655 (N_11655,N_10660,N_10731);
nand U11656 (N_11656,N_10701,N_10026);
or U11657 (N_11657,N_10178,N_10343);
nand U11658 (N_11658,N_10864,N_10653);
nor U11659 (N_11659,N_10695,N_10367);
nor U11660 (N_11660,N_10233,N_10108);
nand U11661 (N_11661,N_10073,N_10572);
or U11662 (N_11662,N_10449,N_10406);
nand U11663 (N_11663,N_10502,N_10307);
xnor U11664 (N_11664,N_10368,N_10237);
xnor U11665 (N_11665,N_10683,N_10685);
nand U11666 (N_11666,N_10512,N_10178);
or U11667 (N_11667,N_10069,N_10606);
nand U11668 (N_11668,N_10170,N_10596);
nor U11669 (N_11669,N_10673,N_10523);
or U11670 (N_11670,N_10267,N_10851);
and U11671 (N_11671,N_10113,N_10067);
and U11672 (N_11672,N_10253,N_10381);
and U11673 (N_11673,N_10184,N_10674);
nor U11674 (N_11674,N_10245,N_10027);
and U11675 (N_11675,N_10148,N_10827);
or U11676 (N_11676,N_10529,N_10460);
xnor U11677 (N_11677,N_10601,N_10616);
or U11678 (N_11678,N_10134,N_10015);
nand U11679 (N_11679,N_10462,N_10616);
or U11680 (N_11680,N_10462,N_10010);
nand U11681 (N_11681,N_10944,N_10715);
nand U11682 (N_11682,N_10205,N_10619);
or U11683 (N_11683,N_10560,N_10312);
nor U11684 (N_11684,N_10235,N_10463);
xnor U11685 (N_11685,N_10924,N_10271);
and U11686 (N_11686,N_10577,N_10933);
nand U11687 (N_11687,N_10567,N_10157);
nand U11688 (N_11688,N_10839,N_10929);
and U11689 (N_11689,N_10341,N_10815);
nor U11690 (N_11690,N_10533,N_10890);
xor U11691 (N_11691,N_10085,N_10695);
nor U11692 (N_11692,N_10265,N_10133);
xor U11693 (N_11693,N_10401,N_10119);
xnor U11694 (N_11694,N_10273,N_10310);
or U11695 (N_11695,N_10480,N_10482);
or U11696 (N_11696,N_10494,N_10895);
xor U11697 (N_11697,N_10730,N_10490);
or U11698 (N_11698,N_10176,N_10356);
or U11699 (N_11699,N_10771,N_10067);
or U11700 (N_11700,N_10329,N_10425);
nand U11701 (N_11701,N_10006,N_10306);
nor U11702 (N_11702,N_10764,N_10049);
xnor U11703 (N_11703,N_10486,N_10441);
nand U11704 (N_11704,N_10444,N_10988);
or U11705 (N_11705,N_10426,N_10198);
nand U11706 (N_11706,N_10857,N_10031);
xnor U11707 (N_11707,N_10863,N_10627);
nand U11708 (N_11708,N_10233,N_10485);
nand U11709 (N_11709,N_10890,N_10801);
xnor U11710 (N_11710,N_10749,N_10139);
and U11711 (N_11711,N_10245,N_10216);
xor U11712 (N_11712,N_10872,N_10254);
or U11713 (N_11713,N_10340,N_10425);
nand U11714 (N_11714,N_10865,N_10462);
nor U11715 (N_11715,N_10682,N_10392);
and U11716 (N_11716,N_10315,N_10164);
or U11717 (N_11717,N_10154,N_10068);
nor U11718 (N_11718,N_10373,N_10048);
nor U11719 (N_11719,N_10839,N_10034);
and U11720 (N_11720,N_10223,N_10091);
nor U11721 (N_11721,N_10516,N_10943);
nor U11722 (N_11722,N_10629,N_10321);
and U11723 (N_11723,N_10483,N_10795);
nand U11724 (N_11724,N_10066,N_10491);
and U11725 (N_11725,N_10379,N_10064);
and U11726 (N_11726,N_10602,N_10214);
xor U11727 (N_11727,N_10935,N_10994);
xnor U11728 (N_11728,N_10670,N_10506);
xnor U11729 (N_11729,N_10212,N_10753);
xor U11730 (N_11730,N_10678,N_10542);
and U11731 (N_11731,N_10851,N_10261);
nand U11732 (N_11732,N_10385,N_10076);
nand U11733 (N_11733,N_10824,N_10601);
nand U11734 (N_11734,N_10755,N_10705);
nand U11735 (N_11735,N_10457,N_10365);
or U11736 (N_11736,N_10047,N_10782);
xnor U11737 (N_11737,N_10515,N_10504);
nor U11738 (N_11738,N_10473,N_10406);
or U11739 (N_11739,N_10310,N_10449);
nand U11740 (N_11740,N_10160,N_10092);
and U11741 (N_11741,N_10600,N_10125);
xnor U11742 (N_11742,N_10739,N_10430);
nand U11743 (N_11743,N_10702,N_10877);
nor U11744 (N_11744,N_10821,N_10724);
nand U11745 (N_11745,N_10771,N_10297);
or U11746 (N_11746,N_10596,N_10864);
xor U11747 (N_11747,N_10378,N_10562);
nand U11748 (N_11748,N_10633,N_10180);
nor U11749 (N_11749,N_10143,N_10897);
nor U11750 (N_11750,N_10002,N_10669);
nand U11751 (N_11751,N_10479,N_10091);
nand U11752 (N_11752,N_10031,N_10838);
or U11753 (N_11753,N_10102,N_10222);
nand U11754 (N_11754,N_10452,N_10060);
and U11755 (N_11755,N_10042,N_10891);
nand U11756 (N_11756,N_10675,N_10776);
nor U11757 (N_11757,N_10313,N_10803);
nand U11758 (N_11758,N_10968,N_10079);
nand U11759 (N_11759,N_10559,N_10439);
or U11760 (N_11760,N_10236,N_10931);
nand U11761 (N_11761,N_10985,N_10460);
nor U11762 (N_11762,N_10070,N_10717);
and U11763 (N_11763,N_10107,N_10386);
and U11764 (N_11764,N_10150,N_10854);
xor U11765 (N_11765,N_10488,N_10361);
or U11766 (N_11766,N_10186,N_10707);
or U11767 (N_11767,N_10647,N_10217);
nor U11768 (N_11768,N_10564,N_10664);
nor U11769 (N_11769,N_10904,N_10025);
xor U11770 (N_11770,N_10408,N_10279);
nor U11771 (N_11771,N_10762,N_10449);
or U11772 (N_11772,N_10890,N_10032);
or U11773 (N_11773,N_10942,N_10664);
nand U11774 (N_11774,N_10196,N_10731);
or U11775 (N_11775,N_10393,N_10449);
nand U11776 (N_11776,N_10437,N_10441);
nor U11777 (N_11777,N_10879,N_10263);
and U11778 (N_11778,N_10555,N_10758);
and U11779 (N_11779,N_10808,N_10508);
nand U11780 (N_11780,N_10734,N_10265);
nand U11781 (N_11781,N_10864,N_10376);
or U11782 (N_11782,N_10078,N_10780);
nor U11783 (N_11783,N_10761,N_10002);
and U11784 (N_11784,N_10379,N_10397);
and U11785 (N_11785,N_10571,N_10691);
nor U11786 (N_11786,N_10231,N_10967);
and U11787 (N_11787,N_10489,N_10321);
nor U11788 (N_11788,N_10415,N_10237);
or U11789 (N_11789,N_10432,N_10521);
nor U11790 (N_11790,N_10907,N_10544);
and U11791 (N_11791,N_10898,N_10165);
or U11792 (N_11792,N_10314,N_10894);
and U11793 (N_11793,N_10168,N_10341);
nand U11794 (N_11794,N_10549,N_10014);
nor U11795 (N_11795,N_10062,N_10892);
nand U11796 (N_11796,N_10764,N_10986);
and U11797 (N_11797,N_10404,N_10403);
or U11798 (N_11798,N_10554,N_10258);
or U11799 (N_11799,N_10187,N_10678);
nor U11800 (N_11800,N_10192,N_10011);
nand U11801 (N_11801,N_10076,N_10888);
nor U11802 (N_11802,N_10247,N_10045);
or U11803 (N_11803,N_10607,N_10395);
nand U11804 (N_11804,N_10480,N_10437);
nand U11805 (N_11805,N_10864,N_10061);
or U11806 (N_11806,N_10074,N_10698);
or U11807 (N_11807,N_10993,N_10115);
nor U11808 (N_11808,N_10239,N_10153);
xnor U11809 (N_11809,N_10799,N_10419);
xnor U11810 (N_11810,N_10506,N_10717);
xnor U11811 (N_11811,N_10427,N_10802);
and U11812 (N_11812,N_10794,N_10211);
nand U11813 (N_11813,N_10549,N_10062);
nand U11814 (N_11814,N_10661,N_10574);
nand U11815 (N_11815,N_10397,N_10533);
and U11816 (N_11816,N_10881,N_10137);
and U11817 (N_11817,N_10335,N_10694);
xnor U11818 (N_11818,N_10706,N_10319);
nor U11819 (N_11819,N_10659,N_10120);
and U11820 (N_11820,N_10066,N_10723);
or U11821 (N_11821,N_10938,N_10950);
nor U11822 (N_11822,N_10075,N_10268);
nor U11823 (N_11823,N_10792,N_10911);
and U11824 (N_11824,N_10374,N_10476);
nand U11825 (N_11825,N_10421,N_10588);
xor U11826 (N_11826,N_10356,N_10138);
nand U11827 (N_11827,N_10352,N_10731);
nor U11828 (N_11828,N_10679,N_10196);
or U11829 (N_11829,N_10921,N_10790);
nor U11830 (N_11830,N_10105,N_10971);
or U11831 (N_11831,N_10209,N_10334);
or U11832 (N_11832,N_10686,N_10024);
and U11833 (N_11833,N_10011,N_10755);
nand U11834 (N_11834,N_10015,N_10235);
nor U11835 (N_11835,N_10645,N_10137);
nand U11836 (N_11836,N_10522,N_10567);
and U11837 (N_11837,N_10263,N_10361);
xor U11838 (N_11838,N_10506,N_10177);
xnor U11839 (N_11839,N_10228,N_10509);
xnor U11840 (N_11840,N_10856,N_10001);
and U11841 (N_11841,N_10793,N_10544);
or U11842 (N_11842,N_10069,N_10819);
nand U11843 (N_11843,N_10676,N_10416);
or U11844 (N_11844,N_10491,N_10782);
or U11845 (N_11845,N_10455,N_10325);
and U11846 (N_11846,N_10295,N_10632);
nor U11847 (N_11847,N_10444,N_10504);
or U11848 (N_11848,N_10232,N_10272);
nand U11849 (N_11849,N_10057,N_10339);
nand U11850 (N_11850,N_10428,N_10743);
and U11851 (N_11851,N_10765,N_10369);
and U11852 (N_11852,N_10581,N_10171);
xnor U11853 (N_11853,N_10002,N_10034);
nor U11854 (N_11854,N_10027,N_10847);
or U11855 (N_11855,N_10458,N_10637);
nor U11856 (N_11856,N_10662,N_10669);
and U11857 (N_11857,N_10529,N_10958);
and U11858 (N_11858,N_10514,N_10185);
and U11859 (N_11859,N_10356,N_10095);
nand U11860 (N_11860,N_10197,N_10481);
xnor U11861 (N_11861,N_10873,N_10971);
or U11862 (N_11862,N_10476,N_10895);
or U11863 (N_11863,N_10236,N_10449);
nor U11864 (N_11864,N_10835,N_10494);
xnor U11865 (N_11865,N_10909,N_10610);
xnor U11866 (N_11866,N_10872,N_10600);
xor U11867 (N_11867,N_10388,N_10005);
and U11868 (N_11868,N_10149,N_10448);
or U11869 (N_11869,N_10182,N_10207);
nand U11870 (N_11870,N_10878,N_10714);
xnor U11871 (N_11871,N_10528,N_10144);
xnor U11872 (N_11872,N_10733,N_10510);
xor U11873 (N_11873,N_10219,N_10007);
nor U11874 (N_11874,N_10058,N_10080);
or U11875 (N_11875,N_10942,N_10491);
nand U11876 (N_11876,N_10503,N_10711);
and U11877 (N_11877,N_10402,N_10103);
and U11878 (N_11878,N_10801,N_10254);
nor U11879 (N_11879,N_10687,N_10212);
nor U11880 (N_11880,N_10724,N_10570);
xor U11881 (N_11881,N_10389,N_10482);
or U11882 (N_11882,N_10302,N_10772);
and U11883 (N_11883,N_10577,N_10221);
and U11884 (N_11884,N_10339,N_10044);
or U11885 (N_11885,N_10222,N_10873);
or U11886 (N_11886,N_10873,N_10207);
or U11887 (N_11887,N_10147,N_10532);
nor U11888 (N_11888,N_10062,N_10390);
nand U11889 (N_11889,N_10247,N_10095);
or U11890 (N_11890,N_10412,N_10041);
nor U11891 (N_11891,N_10666,N_10330);
nand U11892 (N_11892,N_10414,N_10904);
or U11893 (N_11893,N_10551,N_10691);
or U11894 (N_11894,N_10669,N_10083);
xor U11895 (N_11895,N_10269,N_10323);
or U11896 (N_11896,N_10942,N_10945);
nand U11897 (N_11897,N_10457,N_10435);
nand U11898 (N_11898,N_10816,N_10436);
or U11899 (N_11899,N_10647,N_10319);
or U11900 (N_11900,N_10102,N_10040);
nor U11901 (N_11901,N_10590,N_10289);
xor U11902 (N_11902,N_10388,N_10727);
nand U11903 (N_11903,N_10949,N_10326);
xor U11904 (N_11904,N_10137,N_10757);
nand U11905 (N_11905,N_10773,N_10428);
and U11906 (N_11906,N_10894,N_10139);
xor U11907 (N_11907,N_10804,N_10782);
xor U11908 (N_11908,N_10825,N_10610);
nor U11909 (N_11909,N_10789,N_10870);
xor U11910 (N_11910,N_10952,N_10061);
nand U11911 (N_11911,N_10376,N_10591);
nand U11912 (N_11912,N_10684,N_10062);
xnor U11913 (N_11913,N_10962,N_10362);
nand U11914 (N_11914,N_10712,N_10982);
nand U11915 (N_11915,N_10099,N_10159);
nor U11916 (N_11916,N_10464,N_10929);
and U11917 (N_11917,N_10840,N_10954);
xnor U11918 (N_11918,N_10601,N_10508);
and U11919 (N_11919,N_10666,N_10374);
or U11920 (N_11920,N_10434,N_10548);
nor U11921 (N_11921,N_10091,N_10380);
or U11922 (N_11922,N_10597,N_10092);
or U11923 (N_11923,N_10500,N_10359);
or U11924 (N_11924,N_10187,N_10548);
nor U11925 (N_11925,N_10695,N_10139);
xor U11926 (N_11926,N_10705,N_10081);
xor U11927 (N_11927,N_10291,N_10850);
nor U11928 (N_11928,N_10660,N_10756);
and U11929 (N_11929,N_10133,N_10357);
nor U11930 (N_11930,N_10487,N_10376);
or U11931 (N_11931,N_10996,N_10192);
nor U11932 (N_11932,N_10802,N_10295);
nor U11933 (N_11933,N_10064,N_10981);
xor U11934 (N_11934,N_10602,N_10377);
nor U11935 (N_11935,N_10617,N_10445);
or U11936 (N_11936,N_10224,N_10677);
nand U11937 (N_11937,N_10476,N_10034);
nor U11938 (N_11938,N_10107,N_10328);
xnor U11939 (N_11939,N_10357,N_10737);
xnor U11940 (N_11940,N_10740,N_10731);
nor U11941 (N_11941,N_10461,N_10220);
and U11942 (N_11942,N_10759,N_10597);
or U11943 (N_11943,N_10958,N_10357);
xnor U11944 (N_11944,N_10030,N_10364);
nor U11945 (N_11945,N_10237,N_10824);
nor U11946 (N_11946,N_10962,N_10742);
and U11947 (N_11947,N_10679,N_10443);
or U11948 (N_11948,N_10854,N_10719);
nor U11949 (N_11949,N_10802,N_10614);
or U11950 (N_11950,N_10317,N_10537);
nor U11951 (N_11951,N_10392,N_10117);
xnor U11952 (N_11952,N_10761,N_10827);
or U11953 (N_11953,N_10786,N_10259);
xor U11954 (N_11954,N_10120,N_10061);
nand U11955 (N_11955,N_10732,N_10401);
nand U11956 (N_11956,N_10233,N_10576);
and U11957 (N_11957,N_10395,N_10588);
nand U11958 (N_11958,N_10515,N_10138);
and U11959 (N_11959,N_10951,N_10230);
xor U11960 (N_11960,N_10064,N_10624);
nand U11961 (N_11961,N_10490,N_10455);
nor U11962 (N_11962,N_10282,N_10391);
xor U11963 (N_11963,N_10233,N_10552);
nand U11964 (N_11964,N_10218,N_10767);
nand U11965 (N_11965,N_10230,N_10996);
or U11966 (N_11966,N_10820,N_10167);
and U11967 (N_11967,N_10952,N_10108);
xnor U11968 (N_11968,N_10513,N_10350);
or U11969 (N_11969,N_10987,N_10942);
xnor U11970 (N_11970,N_10716,N_10102);
nor U11971 (N_11971,N_10050,N_10751);
nor U11972 (N_11972,N_10162,N_10569);
nand U11973 (N_11973,N_10783,N_10090);
xnor U11974 (N_11974,N_10683,N_10585);
xnor U11975 (N_11975,N_10470,N_10224);
and U11976 (N_11976,N_10142,N_10239);
or U11977 (N_11977,N_10701,N_10862);
xor U11978 (N_11978,N_10857,N_10184);
and U11979 (N_11979,N_10482,N_10922);
nand U11980 (N_11980,N_10520,N_10777);
and U11981 (N_11981,N_10201,N_10258);
xnor U11982 (N_11982,N_10482,N_10588);
nand U11983 (N_11983,N_10465,N_10095);
nand U11984 (N_11984,N_10745,N_10544);
and U11985 (N_11985,N_10812,N_10019);
nor U11986 (N_11986,N_10134,N_10129);
nor U11987 (N_11987,N_10745,N_10150);
or U11988 (N_11988,N_10464,N_10309);
and U11989 (N_11989,N_10067,N_10298);
and U11990 (N_11990,N_10827,N_10699);
nand U11991 (N_11991,N_10939,N_10798);
or U11992 (N_11992,N_10406,N_10424);
xor U11993 (N_11993,N_10441,N_10958);
nand U11994 (N_11994,N_10656,N_10491);
nor U11995 (N_11995,N_10107,N_10781);
nand U11996 (N_11996,N_10128,N_10714);
or U11997 (N_11997,N_10570,N_10383);
nand U11998 (N_11998,N_10941,N_10306);
and U11999 (N_11999,N_10999,N_10125);
nor U12000 (N_12000,N_11793,N_11666);
xnor U12001 (N_12001,N_11124,N_11596);
and U12002 (N_12002,N_11989,N_11484);
or U12003 (N_12003,N_11134,N_11747);
and U12004 (N_12004,N_11859,N_11955);
nand U12005 (N_12005,N_11288,N_11048);
nor U12006 (N_12006,N_11331,N_11084);
nor U12007 (N_12007,N_11910,N_11499);
nor U12008 (N_12008,N_11376,N_11074);
or U12009 (N_12009,N_11758,N_11700);
nor U12010 (N_12010,N_11544,N_11417);
nor U12011 (N_12011,N_11366,N_11297);
nor U12012 (N_12012,N_11834,N_11483);
or U12013 (N_12013,N_11847,N_11335);
or U12014 (N_12014,N_11319,N_11943);
and U12015 (N_12015,N_11628,N_11592);
or U12016 (N_12016,N_11449,N_11980);
nor U12017 (N_12017,N_11810,N_11197);
and U12018 (N_12018,N_11979,N_11919);
nor U12019 (N_12019,N_11768,N_11069);
nand U12020 (N_12020,N_11874,N_11370);
and U12021 (N_12021,N_11873,N_11912);
or U12022 (N_12022,N_11729,N_11017);
or U12023 (N_12023,N_11047,N_11763);
xnor U12024 (N_12024,N_11219,N_11314);
nor U12025 (N_12025,N_11202,N_11339);
or U12026 (N_12026,N_11279,N_11459);
and U12027 (N_12027,N_11389,N_11815);
or U12028 (N_12028,N_11621,N_11665);
and U12029 (N_12029,N_11617,N_11911);
nor U12030 (N_12030,N_11450,N_11591);
nand U12031 (N_12031,N_11467,N_11300);
and U12032 (N_12032,N_11278,N_11864);
nor U12033 (N_12033,N_11368,N_11221);
xor U12034 (N_12034,N_11953,N_11145);
or U12035 (N_12035,N_11462,N_11249);
and U12036 (N_12036,N_11148,N_11528);
and U12037 (N_12037,N_11885,N_11798);
nor U12038 (N_12038,N_11127,N_11647);
xnor U12039 (N_12039,N_11669,N_11492);
nor U12040 (N_12040,N_11143,N_11881);
and U12041 (N_12041,N_11424,N_11745);
nand U12042 (N_12042,N_11854,N_11357);
xor U12043 (N_12043,N_11939,N_11839);
nand U12044 (N_12044,N_11780,N_11915);
nand U12045 (N_12045,N_11120,N_11948);
nor U12046 (N_12046,N_11588,N_11485);
and U12047 (N_12047,N_11493,N_11844);
and U12048 (N_12048,N_11397,N_11056);
nand U12049 (N_12049,N_11900,N_11042);
xnor U12050 (N_12050,N_11648,N_11725);
nor U12051 (N_12051,N_11342,N_11909);
or U12052 (N_12052,N_11287,N_11846);
and U12053 (N_12053,N_11988,N_11585);
and U12054 (N_12054,N_11879,N_11077);
and U12055 (N_12055,N_11014,N_11141);
nand U12056 (N_12056,N_11008,N_11889);
and U12057 (N_12057,N_11573,N_11031);
xnor U12058 (N_12058,N_11777,N_11323);
or U12059 (N_12059,N_11961,N_11905);
nor U12060 (N_12060,N_11371,N_11926);
nor U12061 (N_12061,N_11165,N_11845);
or U12062 (N_12062,N_11868,N_11224);
and U12063 (N_12063,N_11865,N_11950);
nand U12064 (N_12064,N_11749,N_11842);
nor U12065 (N_12065,N_11130,N_11906);
xnor U12066 (N_12066,N_11404,N_11931);
xor U12067 (N_12067,N_11057,N_11916);
nor U12068 (N_12068,N_11536,N_11674);
and U12069 (N_12069,N_11826,N_11550);
xnor U12070 (N_12070,N_11863,N_11533);
and U12071 (N_12071,N_11481,N_11243);
nor U12072 (N_12072,N_11509,N_11754);
or U12073 (N_12073,N_11639,N_11817);
or U12074 (N_12074,N_11814,N_11307);
and U12075 (N_12075,N_11794,N_11626);
or U12076 (N_12076,N_11140,N_11699);
and U12077 (N_12077,N_11242,N_11532);
nor U12078 (N_12078,N_11981,N_11361);
nor U12079 (N_12079,N_11599,N_11809);
or U12080 (N_12080,N_11035,N_11396);
nand U12081 (N_12081,N_11012,N_11313);
xnor U12082 (N_12082,N_11013,N_11748);
nor U12083 (N_12083,N_11354,N_11189);
nor U12084 (N_12084,N_11114,N_11126);
nand U12085 (N_12085,N_11779,N_11121);
and U12086 (N_12086,N_11346,N_11119);
or U12087 (N_12087,N_11066,N_11803);
nor U12088 (N_12088,N_11398,N_11561);
and U12089 (N_12089,N_11386,N_11073);
or U12090 (N_12090,N_11262,N_11791);
and U12091 (N_12091,N_11291,N_11315);
and U12092 (N_12092,N_11995,N_11508);
nand U12093 (N_12093,N_11324,N_11938);
nor U12094 (N_12094,N_11158,N_11717);
xnor U12095 (N_12095,N_11547,N_11616);
nand U12096 (N_12096,N_11843,N_11546);
nor U12097 (N_12097,N_11173,N_11690);
and U12098 (N_12098,N_11043,N_11194);
nand U12099 (N_12099,N_11273,N_11036);
xor U12100 (N_12100,N_11395,N_11682);
nand U12101 (N_12101,N_11106,N_11363);
or U12102 (N_12102,N_11918,N_11125);
or U12103 (N_12103,N_11542,N_11325);
nand U12104 (N_12104,N_11063,N_11782);
or U12105 (N_12105,N_11622,N_11399);
or U12106 (N_12106,N_11082,N_11518);
and U12107 (N_12107,N_11344,N_11551);
and U12108 (N_12108,N_11608,N_11755);
and U12109 (N_12109,N_11799,N_11208);
or U12110 (N_12110,N_11861,N_11226);
xnor U12111 (N_12111,N_11234,N_11466);
nor U12112 (N_12112,N_11212,N_11986);
xor U12113 (N_12113,N_11739,N_11691);
xnor U12114 (N_12114,N_11046,N_11022);
or U12115 (N_12115,N_11445,N_11480);
nor U12116 (N_12116,N_11583,N_11828);
xnor U12117 (N_12117,N_11723,N_11341);
xnor U12118 (N_12118,N_11730,N_11615);
nor U12119 (N_12119,N_11526,N_11316);
or U12120 (N_12120,N_11624,N_11967);
nor U12121 (N_12121,N_11732,N_11963);
nand U12122 (N_12122,N_11892,N_11030);
nand U12123 (N_12123,N_11520,N_11138);
and U12124 (N_12124,N_11813,N_11606);
nand U12125 (N_12125,N_11210,N_11553);
nand U12126 (N_12126,N_11427,N_11860);
xnor U12127 (N_12127,N_11867,N_11137);
or U12128 (N_12128,N_11175,N_11461);
nand U12129 (N_12129,N_11770,N_11964);
xor U12130 (N_12130,N_11973,N_11488);
nand U12131 (N_12131,N_11935,N_11719);
xnor U12132 (N_12132,N_11766,N_11949);
and U12133 (N_12133,N_11517,N_11391);
xor U12134 (N_12134,N_11601,N_11038);
xor U12135 (N_12135,N_11159,N_11771);
xor U12136 (N_12136,N_11235,N_11061);
nand U12137 (N_12137,N_11802,N_11068);
and U12138 (N_12138,N_11196,N_11537);
nor U12139 (N_12139,N_11452,N_11280);
nand U12140 (N_12140,N_11549,N_11166);
or U12141 (N_12141,N_11220,N_11516);
and U12142 (N_12142,N_11060,N_11207);
and U12143 (N_12143,N_11428,N_11992);
nand U12144 (N_12144,N_11205,N_11232);
nor U12145 (N_12145,N_11115,N_11091);
or U12146 (N_12146,N_11922,N_11160);
nand U12147 (N_12147,N_11555,N_11659);
and U12148 (N_12148,N_11439,N_11535);
nand U12149 (N_12149,N_11584,N_11538);
or U12150 (N_12150,N_11942,N_11736);
or U12151 (N_12151,N_11811,N_11654);
nand U12152 (N_12152,N_11971,N_11463);
nand U12153 (N_12153,N_11855,N_11378);
or U12154 (N_12154,N_11470,N_11714);
nor U12155 (N_12155,N_11218,N_11364);
and U12156 (N_12156,N_11193,N_11330);
and U12157 (N_12157,N_11633,N_11681);
nor U12158 (N_12158,N_11925,N_11415);
or U12159 (N_12159,N_11422,N_11675);
and U12160 (N_12160,N_11122,N_11150);
and U12161 (N_12161,N_11656,N_11525);
or U12162 (N_12162,N_11952,N_11495);
xnor U12163 (N_12163,N_11129,N_11029);
and U12164 (N_12164,N_11206,N_11151);
nand U12165 (N_12165,N_11728,N_11959);
nor U12166 (N_12166,N_11848,N_11095);
xor U12167 (N_12167,N_11101,N_11917);
and U12168 (N_12168,N_11618,N_11781);
and U12169 (N_12169,N_11812,N_11001);
and U12170 (N_12170,N_11103,N_11079);
or U12171 (N_12171,N_11365,N_11045);
and U12172 (N_12172,N_11425,N_11712);
nand U12173 (N_12173,N_11414,N_11455);
nor U12174 (N_12174,N_11807,N_11667);
xor U12175 (N_12175,N_11104,N_11083);
and U12176 (N_12176,N_11275,N_11394);
nor U12177 (N_12177,N_11527,N_11559);
nand U12178 (N_12178,N_11946,N_11521);
nor U12179 (N_12179,N_11642,N_11420);
xnor U12180 (N_12180,N_11977,N_11403);
and U12181 (N_12181,N_11698,N_11856);
nand U12182 (N_12182,N_11058,N_11746);
nand U12183 (N_12183,N_11440,N_11572);
xor U12184 (N_12184,N_11002,N_11080);
nand U12185 (N_12185,N_11541,N_11976);
and U12186 (N_12186,N_11759,N_11109);
and U12187 (N_12187,N_11947,N_11568);
or U12188 (N_12188,N_11136,N_11734);
or U12189 (N_12189,N_11767,N_11345);
and U12190 (N_12190,N_11635,N_11178);
nand U12191 (N_12191,N_11737,N_11443);
or U12192 (N_12192,N_11380,N_11116);
or U12193 (N_12193,N_11904,N_11231);
or U12194 (N_12194,N_11164,N_11882);
or U12195 (N_12195,N_11604,N_11523);
xor U12196 (N_12196,N_11962,N_11993);
xnor U12197 (N_12197,N_11418,N_11021);
nor U12198 (N_12198,N_11720,N_11870);
or U12199 (N_12199,N_11410,N_11876);
xnor U12200 (N_12200,N_11306,N_11144);
nand U12201 (N_12201,N_11545,N_11304);
and U12202 (N_12202,N_11695,N_11582);
or U12203 (N_12203,N_11686,N_11914);
nand U12204 (N_12204,N_11227,N_11708);
and U12205 (N_12205,N_11776,N_11460);
xor U12206 (N_12206,N_11658,N_11172);
nand U12207 (N_12207,N_11531,N_11678);
and U12208 (N_12208,N_11849,N_11477);
and U12209 (N_12209,N_11271,N_11374);
and U12210 (N_12210,N_11498,N_11786);
and U12211 (N_12211,N_11603,N_11142);
nand U12212 (N_12212,N_11894,N_11177);
xor U12213 (N_12213,N_11188,N_11586);
or U12214 (N_12214,N_11373,N_11442);
nand U12215 (N_12215,N_11975,N_11750);
xnor U12216 (N_12216,N_11731,N_11774);
xnor U12217 (N_12217,N_11289,N_11796);
and U12218 (N_12218,N_11825,N_11381);
nand U12219 (N_12219,N_11853,N_11349);
or U12220 (N_12220,N_11651,N_11147);
or U12221 (N_12221,N_11321,N_11260);
xor U12222 (N_12222,N_11169,N_11075);
nand U12223 (N_12223,N_11186,N_11097);
and U12224 (N_12224,N_11878,N_11862);
and U12225 (N_12225,N_11240,N_11311);
nand U12226 (N_12226,N_11923,N_11703);
and U12227 (N_12227,N_11710,N_11184);
nor U12228 (N_12228,N_11872,N_11901);
nor U12229 (N_12229,N_11377,N_11757);
or U12230 (N_12230,N_11896,N_11276);
nor U12231 (N_12231,N_11448,N_11434);
nand U12232 (N_12232,N_11217,N_11400);
xor U12233 (N_12233,N_11429,N_11185);
xnor U12234 (N_12234,N_11790,N_11707);
or U12235 (N_12235,N_11643,N_11183);
nand U12236 (N_12236,N_11944,N_11111);
and U12237 (N_12237,N_11436,N_11510);
xnor U12238 (N_12238,N_11741,N_11054);
or U12239 (N_12239,N_11581,N_11577);
nand U12240 (N_12240,N_11662,N_11941);
and U12241 (N_12241,N_11102,N_11494);
or U12242 (N_12242,N_11688,N_11630);
nor U12243 (N_12243,N_11623,N_11500);
and U12244 (N_12244,N_11552,N_11329);
or U12245 (N_12245,N_11457,N_11997);
xnor U12246 (N_12246,N_11836,N_11388);
nand U12247 (N_12247,N_11044,N_11089);
or U12248 (N_12248,N_11530,N_11390);
xnor U12249 (N_12249,N_11762,N_11071);
xnor U12250 (N_12250,N_11562,N_11247);
xor U12251 (N_12251,N_11123,N_11308);
or U12252 (N_12252,N_11170,N_11564);
xnor U12253 (N_12253,N_11884,N_11664);
nand U12254 (N_12254,N_11255,N_11011);
nor U12255 (N_12255,N_11640,N_11360);
nor U12256 (N_12256,N_11792,N_11641);
nor U12257 (N_12257,N_11026,N_11936);
nor U12258 (N_12258,N_11299,N_11246);
nand U12259 (N_12259,N_11627,N_11451);
and U12260 (N_12260,N_11020,N_11524);
and U12261 (N_12261,N_11253,N_11998);
nor U12262 (N_12262,N_11927,N_11567);
and U12263 (N_12263,N_11327,N_11401);
or U12264 (N_12264,N_11515,N_11819);
nand U12265 (N_12265,N_11190,N_11233);
nor U12266 (N_12266,N_11869,N_11668);
nor U12267 (N_12267,N_11358,N_11851);
and U12268 (N_12268,N_11850,N_11180);
or U12269 (N_12269,N_11003,N_11554);
and U12270 (N_12270,N_11877,N_11742);
xnor U12271 (N_12271,N_11818,N_11644);
xor U12272 (N_12272,N_11684,N_11310);
nor U12273 (N_12273,N_11661,N_11801);
or U12274 (N_12274,N_11441,N_11446);
nand U12275 (N_12275,N_11128,N_11468);
nand U12276 (N_12276,N_11954,N_11272);
or U12277 (N_12277,N_11191,N_11489);
or U12278 (N_12278,N_11264,N_11800);
nor U12279 (N_12279,N_11025,N_11174);
or U12280 (N_12280,N_11340,N_11406);
and U12281 (N_12281,N_11829,N_11282);
nand U12282 (N_12282,N_11486,N_11318);
xnor U12283 (N_12283,N_11317,N_11740);
and U12284 (N_12284,N_11795,N_11579);
or U12285 (N_12285,N_11006,N_11804);
or U12286 (N_12286,N_11211,N_11000);
xnor U12287 (N_12287,N_11895,N_11018);
nand U12288 (N_12288,N_11823,N_11689);
xor U12289 (N_12289,N_11407,N_11663);
nor U12290 (N_12290,N_11511,N_11760);
and U12291 (N_12291,N_11744,N_11806);
or U12292 (N_12292,N_11866,N_11437);
xnor U12293 (N_12293,N_11822,N_11702);
and U12294 (N_12294,N_11576,N_11041);
nor U12295 (N_12295,N_11292,N_11356);
xnor U12296 (N_12296,N_11670,N_11419);
or U12297 (N_12297,N_11225,N_11506);
nand U12298 (N_12298,N_11519,N_11685);
nand U12299 (N_12299,N_11118,N_11637);
or U12300 (N_12300,N_11808,N_11204);
nor U12301 (N_12301,N_11093,N_11051);
nor U12302 (N_12302,N_11384,N_11081);
xnor U12303 (N_12303,N_11230,N_11430);
nand U12304 (N_12304,N_11984,N_11574);
or U12305 (N_12305,N_11987,N_11921);
or U12306 (N_12306,N_11298,N_11956);
or U12307 (N_12307,N_11350,N_11969);
or U12308 (N_12308,N_11629,N_11171);
xnor U12309 (N_12309,N_11871,N_11548);
nor U12310 (N_12310,N_11610,N_11652);
nand U12311 (N_12311,N_11367,N_11775);
xnor U12312 (N_12312,N_11268,N_11065);
nand U12313 (N_12313,N_11062,N_11228);
nand U12314 (N_12314,N_11764,N_11203);
nor U12315 (N_12315,N_11891,N_11625);
and U12316 (N_12316,N_11416,N_11858);
and U12317 (N_12317,N_11263,N_11705);
nand U12318 (N_12318,N_11704,N_11250);
nor U12319 (N_12319,N_11229,N_11501);
nand U12320 (N_12320,N_11216,N_11507);
and U12321 (N_12321,N_11985,N_11301);
nand U12322 (N_12322,N_11765,N_11888);
or U12323 (N_12323,N_11679,N_11636);
nor U12324 (N_12324,N_11176,N_11383);
nand U12325 (N_12325,N_11209,N_11088);
nand U12326 (N_12326,N_11650,N_11085);
xnor U12327 (N_12327,N_11478,N_11598);
xnor U12328 (N_12328,N_11072,N_11474);
and U12329 (N_12329,N_11033,N_11653);
xor U12330 (N_12330,N_11199,N_11261);
nand U12331 (N_12331,N_11432,N_11824);
and U12332 (N_12332,N_11351,N_11692);
nor U12333 (N_12333,N_11673,N_11009);
nand U12334 (N_12334,N_11198,N_11886);
and U12335 (N_12335,N_11413,N_11334);
and U12336 (N_12336,N_11497,N_11566);
or U12337 (N_12337,N_11438,N_11490);
or U12338 (N_12338,N_11087,N_11727);
and U12339 (N_12339,N_11099,N_11933);
nand U12340 (N_12340,N_11743,N_11277);
xor U12341 (N_12341,N_11619,N_11464);
or U12342 (N_12342,N_11837,N_11857);
xor U12343 (N_12343,N_11110,N_11290);
nand U12344 (N_12344,N_11722,N_11426);
nor U12345 (N_12345,N_11241,N_11258);
and U12346 (N_12346,N_11213,N_11028);
nor U12347 (N_12347,N_11752,N_11951);
and U12348 (N_12348,N_11179,N_11154);
xnor U12349 (N_12349,N_11902,N_11597);
or U12350 (N_12350,N_11458,N_11605);
or U12351 (N_12351,N_11067,N_11117);
xor U12352 (N_12352,N_11100,N_11965);
xnor U12353 (N_12353,N_11660,N_11472);
and U12354 (N_12354,N_11153,N_11840);
nand U12355 (N_12355,N_11983,N_11718);
nand U12356 (N_12356,N_11274,N_11833);
or U12357 (N_12357,N_11590,N_11254);
and U12358 (N_12358,N_11163,N_11522);
and U12359 (N_12359,N_11303,N_11333);
xnor U12360 (N_12360,N_11789,N_11353);
or U12361 (N_12361,N_11076,N_11267);
or U12362 (N_12362,N_11751,N_11677);
nand U12363 (N_12363,N_11269,N_11676);
nand U12364 (N_12364,N_11096,N_11393);
nor U12365 (N_12365,N_11050,N_11638);
and U12366 (N_12366,N_11402,N_11543);
or U12367 (N_12367,N_11112,N_11680);
and U12368 (N_12368,N_11423,N_11052);
nand U12369 (N_12369,N_11612,N_11600);
or U12370 (N_12370,N_11248,N_11558);
or U12371 (N_12371,N_11835,N_11724);
and U12372 (N_12372,N_11991,N_11570);
and U12373 (N_12373,N_11502,N_11940);
nand U12374 (N_12374,N_11296,N_11907);
xor U12375 (N_12375,N_11156,N_11375);
nor U12376 (N_12376,N_11256,N_11168);
xor U12377 (N_12377,N_11534,N_11696);
xor U12378 (N_12378,N_11015,N_11830);
and U12379 (N_12379,N_11968,N_11305);
nand U12380 (N_12380,N_11982,N_11960);
nand U12381 (N_12381,N_11475,N_11182);
and U12382 (N_12382,N_11631,N_11974);
nor U12383 (N_12383,N_11575,N_11004);
and U12384 (N_12384,N_11343,N_11487);
or U12385 (N_12385,N_11094,N_11970);
and U12386 (N_12386,N_11738,N_11482);
or U12387 (N_12387,N_11034,N_11512);
or U12388 (N_12388,N_11613,N_11369);
nand U12389 (N_12389,N_11222,N_11411);
and U12390 (N_12390,N_11966,N_11785);
nor U12391 (N_12391,N_11338,N_11924);
and U12392 (N_12392,N_11412,N_11958);
and U12393 (N_12393,N_11328,N_11049);
nand U12394 (N_12394,N_11761,N_11713);
nor U12395 (N_12395,N_11563,N_11133);
xor U12396 (N_12396,N_11587,N_11146);
or U12397 (N_12397,N_11937,N_11701);
or U12398 (N_12398,N_11820,N_11105);
xnor U12399 (N_12399,N_11040,N_11281);
nor U12400 (N_12400,N_11244,N_11721);
nor U12401 (N_12401,N_11753,N_11469);
nand U12402 (N_12402,N_11620,N_11898);
or U12403 (N_12403,N_11504,N_11214);
and U12404 (N_12404,N_11920,N_11649);
and U12405 (N_12405,N_11694,N_11609);
or U12406 (N_12406,N_11108,N_11132);
nand U12407 (N_12407,N_11238,N_11706);
nor U12408 (N_12408,N_11726,N_11852);
and U12409 (N_12409,N_11897,N_11201);
and U12410 (N_12410,N_11405,N_11392);
and U12411 (N_12411,N_11805,N_11756);
nor U12412 (N_12412,N_11131,N_11711);
or U12413 (N_12413,N_11037,N_11816);
nor U12414 (N_12414,N_11454,N_11155);
nor U12415 (N_12415,N_11787,N_11135);
and U12416 (N_12416,N_11893,N_11320);
nor U12417 (N_12417,N_11447,N_11362);
nor U12418 (N_12418,N_11880,N_11187);
or U12419 (N_12419,N_11646,N_11589);
xor U12420 (N_12420,N_11539,N_11379);
nor U12421 (N_12421,N_11832,N_11769);
nor U12422 (N_12422,N_11433,N_11778);
nor U12423 (N_12423,N_11252,N_11284);
xnor U12424 (N_12424,N_11514,N_11972);
xor U12425 (N_12425,N_11286,N_11540);
nor U12426 (N_12426,N_11611,N_11294);
nor U12427 (N_12427,N_11347,N_11431);
nor U12428 (N_12428,N_11382,N_11996);
nand U12429 (N_12429,N_11875,N_11479);
nor U12430 (N_12430,N_11657,N_11529);
and U12431 (N_12431,N_11435,N_11978);
or U12432 (N_12432,N_11773,N_11453);
nor U12433 (N_12433,N_11326,N_11053);
or U12434 (N_12434,N_11465,N_11332);
nor U12435 (N_12435,N_11709,N_11064);
nand U12436 (N_12436,N_11655,N_11632);
nor U12437 (N_12437,N_11560,N_11149);
or U12438 (N_12438,N_11309,N_11784);
and U12439 (N_12439,N_11557,N_11283);
or U12440 (N_12440,N_11223,N_11107);
nand U12441 (N_12441,N_11945,N_11285);
or U12442 (N_12442,N_11994,N_11181);
nand U12443 (N_12443,N_11595,N_11571);
or U12444 (N_12444,N_11827,N_11016);
xnor U12445 (N_12445,N_11602,N_11565);
nor U12446 (N_12446,N_11070,N_11783);
and U12447 (N_12447,N_11359,N_11270);
or U12448 (N_12448,N_11990,N_11473);
xor U12449 (N_12449,N_11716,N_11928);
nand U12450 (N_12450,N_11957,N_11594);
nand U12451 (N_12451,N_11312,N_11078);
and U12452 (N_12452,N_11337,N_11302);
nand U12453 (N_12453,N_11239,N_11265);
nand U12454 (N_12454,N_11192,N_11614);
xnor U12455 (N_12455,N_11055,N_11934);
nor U12456 (N_12456,N_11697,N_11090);
and U12457 (N_12457,N_11887,N_11788);
or U12458 (N_12458,N_11913,N_11024);
or U12459 (N_12459,N_11161,N_11797);
or U12460 (N_12460,N_11735,N_11772);
nand U12461 (N_12461,N_11999,N_11336);
or U12462 (N_12462,N_11841,N_11456);
nor U12463 (N_12463,N_11408,N_11113);
or U12464 (N_12464,N_11569,N_11259);
and U12465 (N_12465,N_11491,N_11010);
xor U12466 (N_12466,N_11385,N_11251);
and U12467 (N_12467,N_11930,N_11007);
or U12468 (N_12468,N_11838,N_11580);
nor U12469 (N_12469,N_11513,N_11634);
nand U12470 (N_12470,N_11476,N_11295);
or U12471 (N_12471,N_11821,N_11086);
and U12472 (N_12472,N_11215,N_11903);
or U12473 (N_12473,N_11733,N_11257);
xnor U12474 (N_12474,N_11027,N_11355);
nor U12475 (N_12475,N_11039,N_11929);
xor U12476 (N_12476,N_11245,N_11899);
or U12477 (N_12477,N_11693,N_11387);
nor U12478 (N_12478,N_11496,N_11645);
nor U12479 (N_12479,N_11578,N_11671);
nor U12480 (N_12480,N_11157,N_11908);
nand U12481 (N_12481,N_11162,N_11293);
xnor U12482 (N_12482,N_11715,N_11352);
or U12483 (N_12483,N_11409,N_11023);
nand U12484 (N_12484,N_11200,N_11322);
nor U12485 (N_12485,N_11471,N_11505);
nor U12486 (N_12486,N_11167,N_11593);
nand U12487 (N_12487,N_11883,N_11139);
xor U12488 (N_12488,N_11266,N_11098);
xor U12489 (N_12489,N_11236,N_11683);
and U12490 (N_12490,N_11607,N_11372);
or U12491 (N_12491,N_11348,N_11237);
xor U12492 (N_12492,N_11444,N_11152);
and U12493 (N_12493,N_11059,N_11195);
or U12494 (N_12494,N_11831,N_11421);
nand U12495 (N_12495,N_11556,N_11687);
nor U12496 (N_12496,N_11005,N_11672);
xnor U12497 (N_12497,N_11890,N_11503);
nand U12498 (N_12498,N_11019,N_11092);
and U12499 (N_12499,N_11932,N_11032);
and U12500 (N_12500,N_11754,N_11422);
xor U12501 (N_12501,N_11906,N_11084);
and U12502 (N_12502,N_11184,N_11360);
xor U12503 (N_12503,N_11958,N_11045);
or U12504 (N_12504,N_11918,N_11858);
nor U12505 (N_12505,N_11466,N_11109);
nand U12506 (N_12506,N_11702,N_11446);
nor U12507 (N_12507,N_11231,N_11253);
and U12508 (N_12508,N_11764,N_11945);
and U12509 (N_12509,N_11752,N_11064);
nand U12510 (N_12510,N_11169,N_11359);
nor U12511 (N_12511,N_11289,N_11991);
nand U12512 (N_12512,N_11537,N_11272);
nor U12513 (N_12513,N_11646,N_11058);
nand U12514 (N_12514,N_11752,N_11366);
and U12515 (N_12515,N_11720,N_11726);
nor U12516 (N_12516,N_11770,N_11869);
nor U12517 (N_12517,N_11961,N_11588);
and U12518 (N_12518,N_11639,N_11427);
xnor U12519 (N_12519,N_11503,N_11562);
nand U12520 (N_12520,N_11052,N_11484);
xor U12521 (N_12521,N_11029,N_11522);
nor U12522 (N_12522,N_11993,N_11232);
nor U12523 (N_12523,N_11715,N_11009);
or U12524 (N_12524,N_11071,N_11697);
xor U12525 (N_12525,N_11700,N_11279);
or U12526 (N_12526,N_11666,N_11173);
nor U12527 (N_12527,N_11430,N_11909);
and U12528 (N_12528,N_11054,N_11996);
xor U12529 (N_12529,N_11841,N_11698);
or U12530 (N_12530,N_11348,N_11554);
xor U12531 (N_12531,N_11476,N_11106);
and U12532 (N_12532,N_11823,N_11782);
nor U12533 (N_12533,N_11338,N_11532);
or U12534 (N_12534,N_11585,N_11667);
and U12535 (N_12535,N_11293,N_11021);
xnor U12536 (N_12536,N_11541,N_11746);
or U12537 (N_12537,N_11900,N_11727);
and U12538 (N_12538,N_11015,N_11691);
and U12539 (N_12539,N_11918,N_11140);
nand U12540 (N_12540,N_11037,N_11540);
xnor U12541 (N_12541,N_11158,N_11218);
nand U12542 (N_12542,N_11331,N_11444);
and U12543 (N_12543,N_11210,N_11460);
or U12544 (N_12544,N_11606,N_11635);
nand U12545 (N_12545,N_11169,N_11765);
nor U12546 (N_12546,N_11401,N_11989);
xnor U12547 (N_12547,N_11446,N_11113);
nor U12548 (N_12548,N_11362,N_11999);
xnor U12549 (N_12549,N_11143,N_11002);
nor U12550 (N_12550,N_11713,N_11794);
nand U12551 (N_12551,N_11111,N_11239);
nor U12552 (N_12552,N_11634,N_11049);
or U12553 (N_12553,N_11429,N_11808);
and U12554 (N_12554,N_11705,N_11608);
and U12555 (N_12555,N_11710,N_11099);
and U12556 (N_12556,N_11176,N_11801);
and U12557 (N_12557,N_11371,N_11376);
and U12558 (N_12558,N_11629,N_11103);
and U12559 (N_12559,N_11173,N_11101);
nand U12560 (N_12560,N_11052,N_11861);
and U12561 (N_12561,N_11579,N_11169);
and U12562 (N_12562,N_11964,N_11513);
nor U12563 (N_12563,N_11641,N_11235);
xor U12564 (N_12564,N_11479,N_11374);
xnor U12565 (N_12565,N_11781,N_11388);
nand U12566 (N_12566,N_11092,N_11656);
and U12567 (N_12567,N_11703,N_11272);
nor U12568 (N_12568,N_11582,N_11358);
xnor U12569 (N_12569,N_11039,N_11634);
and U12570 (N_12570,N_11761,N_11632);
and U12571 (N_12571,N_11334,N_11376);
or U12572 (N_12572,N_11472,N_11458);
and U12573 (N_12573,N_11066,N_11020);
and U12574 (N_12574,N_11373,N_11401);
and U12575 (N_12575,N_11783,N_11257);
or U12576 (N_12576,N_11573,N_11115);
and U12577 (N_12577,N_11066,N_11287);
nand U12578 (N_12578,N_11999,N_11226);
or U12579 (N_12579,N_11040,N_11241);
nor U12580 (N_12580,N_11473,N_11350);
and U12581 (N_12581,N_11542,N_11167);
xor U12582 (N_12582,N_11758,N_11655);
nor U12583 (N_12583,N_11859,N_11818);
nor U12584 (N_12584,N_11849,N_11993);
or U12585 (N_12585,N_11632,N_11050);
nand U12586 (N_12586,N_11894,N_11806);
nor U12587 (N_12587,N_11690,N_11681);
nor U12588 (N_12588,N_11343,N_11667);
or U12589 (N_12589,N_11822,N_11057);
and U12590 (N_12590,N_11381,N_11499);
nor U12591 (N_12591,N_11710,N_11281);
nand U12592 (N_12592,N_11898,N_11141);
and U12593 (N_12593,N_11682,N_11783);
and U12594 (N_12594,N_11670,N_11794);
xnor U12595 (N_12595,N_11953,N_11025);
and U12596 (N_12596,N_11700,N_11494);
nand U12597 (N_12597,N_11578,N_11357);
nor U12598 (N_12598,N_11511,N_11335);
or U12599 (N_12599,N_11946,N_11485);
nand U12600 (N_12600,N_11425,N_11059);
xnor U12601 (N_12601,N_11578,N_11116);
nor U12602 (N_12602,N_11073,N_11252);
and U12603 (N_12603,N_11763,N_11744);
xor U12604 (N_12604,N_11015,N_11357);
nand U12605 (N_12605,N_11086,N_11595);
xnor U12606 (N_12606,N_11375,N_11910);
or U12607 (N_12607,N_11878,N_11318);
xnor U12608 (N_12608,N_11614,N_11746);
and U12609 (N_12609,N_11610,N_11694);
and U12610 (N_12610,N_11000,N_11898);
or U12611 (N_12611,N_11946,N_11101);
nor U12612 (N_12612,N_11675,N_11339);
nand U12613 (N_12613,N_11700,N_11019);
xor U12614 (N_12614,N_11630,N_11760);
nand U12615 (N_12615,N_11082,N_11102);
and U12616 (N_12616,N_11133,N_11759);
or U12617 (N_12617,N_11622,N_11339);
nor U12618 (N_12618,N_11310,N_11854);
or U12619 (N_12619,N_11512,N_11631);
nor U12620 (N_12620,N_11402,N_11635);
or U12621 (N_12621,N_11462,N_11679);
nand U12622 (N_12622,N_11299,N_11722);
xnor U12623 (N_12623,N_11325,N_11173);
or U12624 (N_12624,N_11858,N_11472);
or U12625 (N_12625,N_11460,N_11368);
nor U12626 (N_12626,N_11481,N_11257);
nand U12627 (N_12627,N_11655,N_11933);
or U12628 (N_12628,N_11430,N_11148);
xor U12629 (N_12629,N_11929,N_11299);
or U12630 (N_12630,N_11539,N_11867);
nand U12631 (N_12631,N_11977,N_11210);
and U12632 (N_12632,N_11438,N_11135);
nand U12633 (N_12633,N_11796,N_11156);
nand U12634 (N_12634,N_11870,N_11162);
nor U12635 (N_12635,N_11975,N_11172);
nor U12636 (N_12636,N_11463,N_11807);
or U12637 (N_12637,N_11589,N_11065);
nor U12638 (N_12638,N_11199,N_11987);
and U12639 (N_12639,N_11921,N_11692);
or U12640 (N_12640,N_11518,N_11024);
nand U12641 (N_12641,N_11598,N_11762);
or U12642 (N_12642,N_11341,N_11939);
nand U12643 (N_12643,N_11337,N_11759);
and U12644 (N_12644,N_11128,N_11281);
nor U12645 (N_12645,N_11699,N_11500);
nor U12646 (N_12646,N_11269,N_11412);
and U12647 (N_12647,N_11084,N_11045);
nor U12648 (N_12648,N_11945,N_11892);
and U12649 (N_12649,N_11584,N_11343);
xnor U12650 (N_12650,N_11302,N_11300);
or U12651 (N_12651,N_11923,N_11978);
nor U12652 (N_12652,N_11473,N_11956);
and U12653 (N_12653,N_11942,N_11899);
xnor U12654 (N_12654,N_11693,N_11027);
xor U12655 (N_12655,N_11437,N_11592);
and U12656 (N_12656,N_11136,N_11594);
nor U12657 (N_12657,N_11267,N_11838);
and U12658 (N_12658,N_11145,N_11146);
nor U12659 (N_12659,N_11100,N_11742);
nand U12660 (N_12660,N_11321,N_11861);
and U12661 (N_12661,N_11452,N_11148);
or U12662 (N_12662,N_11845,N_11355);
and U12663 (N_12663,N_11321,N_11546);
nand U12664 (N_12664,N_11724,N_11121);
or U12665 (N_12665,N_11854,N_11105);
xnor U12666 (N_12666,N_11265,N_11053);
and U12667 (N_12667,N_11466,N_11678);
nand U12668 (N_12668,N_11539,N_11633);
xnor U12669 (N_12669,N_11707,N_11010);
nor U12670 (N_12670,N_11054,N_11544);
and U12671 (N_12671,N_11055,N_11768);
nor U12672 (N_12672,N_11735,N_11890);
xnor U12673 (N_12673,N_11479,N_11254);
nand U12674 (N_12674,N_11408,N_11304);
and U12675 (N_12675,N_11358,N_11213);
nand U12676 (N_12676,N_11443,N_11118);
nor U12677 (N_12677,N_11723,N_11687);
xnor U12678 (N_12678,N_11879,N_11088);
or U12679 (N_12679,N_11881,N_11480);
nor U12680 (N_12680,N_11983,N_11914);
xor U12681 (N_12681,N_11843,N_11031);
nand U12682 (N_12682,N_11448,N_11277);
and U12683 (N_12683,N_11320,N_11256);
xor U12684 (N_12684,N_11459,N_11857);
or U12685 (N_12685,N_11307,N_11859);
nand U12686 (N_12686,N_11158,N_11950);
xor U12687 (N_12687,N_11910,N_11836);
xor U12688 (N_12688,N_11931,N_11183);
nand U12689 (N_12689,N_11122,N_11506);
xor U12690 (N_12690,N_11566,N_11435);
nand U12691 (N_12691,N_11669,N_11317);
nand U12692 (N_12692,N_11472,N_11758);
and U12693 (N_12693,N_11124,N_11407);
xnor U12694 (N_12694,N_11994,N_11937);
xor U12695 (N_12695,N_11599,N_11098);
nor U12696 (N_12696,N_11669,N_11489);
or U12697 (N_12697,N_11768,N_11744);
xnor U12698 (N_12698,N_11830,N_11058);
nor U12699 (N_12699,N_11222,N_11291);
xnor U12700 (N_12700,N_11855,N_11820);
or U12701 (N_12701,N_11500,N_11926);
nor U12702 (N_12702,N_11019,N_11311);
nand U12703 (N_12703,N_11466,N_11384);
nor U12704 (N_12704,N_11790,N_11397);
and U12705 (N_12705,N_11722,N_11272);
nor U12706 (N_12706,N_11782,N_11530);
xor U12707 (N_12707,N_11094,N_11453);
or U12708 (N_12708,N_11544,N_11437);
nand U12709 (N_12709,N_11874,N_11331);
xor U12710 (N_12710,N_11147,N_11823);
nor U12711 (N_12711,N_11642,N_11587);
nor U12712 (N_12712,N_11968,N_11081);
nor U12713 (N_12713,N_11419,N_11459);
nor U12714 (N_12714,N_11392,N_11253);
xor U12715 (N_12715,N_11511,N_11871);
nand U12716 (N_12716,N_11706,N_11096);
and U12717 (N_12717,N_11139,N_11983);
and U12718 (N_12718,N_11817,N_11735);
nor U12719 (N_12719,N_11804,N_11785);
or U12720 (N_12720,N_11297,N_11634);
nor U12721 (N_12721,N_11323,N_11536);
and U12722 (N_12722,N_11493,N_11922);
nor U12723 (N_12723,N_11494,N_11523);
or U12724 (N_12724,N_11911,N_11748);
and U12725 (N_12725,N_11809,N_11316);
nand U12726 (N_12726,N_11236,N_11139);
or U12727 (N_12727,N_11012,N_11992);
nand U12728 (N_12728,N_11462,N_11117);
xnor U12729 (N_12729,N_11067,N_11558);
and U12730 (N_12730,N_11187,N_11204);
nand U12731 (N_12731,N_11267,N_11435);
xnor U12732 (N_12732,N_11997,N_11724);
nor U12733 (N_12733,N_11602,N_11012);
or U12734 (N_12734,N_11514,N_11119);
nor U12735 (N_12735,N_11947,N_11455);
nor U12736 (N_12736,N_11119,N_11094);
or U12737 (N_12737,N_11427,N_11701);
and U12738 (N_12738,N_11488,N_11165);
xor U12739 (N_12739,N_11238,N_11041);
nand U12740 (N_12740,N_11319,N_11119);
nand U12741 (N_12741,N_11021,N_11903);
and U12742 (N_12742,N_11794,N_11234);
nand U12743 (N_12743,N_11463,N_11241);
and U12744 (N_12744,N_11803,N_11510);
and U12745 (N_12745,N_11787,N_11053);
and U12746 (N_12746,N_11087,N_11251);
nor U12747 (N_12747,N_11741,N_11677);
or U12748 (N_12748,N_11409,N_11493);
xor U12749 (N_12749,N_11624,N_11484);
and U12750 (N_12750,N_11717,N_11230);
or U12751 (N_12751,N_11745,N_11502);
xor U12752 (N_12752,N_11673,N_11476);
xor U12753 (N_12753,N_11524,N_11699);
nand U12754 (N_12754,N_11125,N_11217);
nand U12755 (N_12755,N_11810,N_11063);
xnor U12756 (N_12756,N_11396,N_11938);
nand U12757 (N_12757,N_11555,N_11502);
or U12758 (N_12758,N_11406,N_11168);
and U12759 (N_12759,N_11515,N_11477);
and U12760 (N_12760,N_11437,N_11245);
or U12761 (N_12761,N_11970,N_11329);
nand U12762 (N_12762,N_11262,N_11229);
nor U12763 (N_12763,N_11609,N_11514);
nand U12764 (N_12764,N_11387,N_11911);
nand U12765 (N_12765,N_11371,N_11920);
and U12766 (N_12766,N_11724,N_11587);
xor U12767 (N_12767,N_11927,N_11631);
or U12768 (N_12768,N_11572,N_11468);
nand U12769 (N_12769,N_11919,N_11326);
and U12770 (N_12770,N_11331,N_11868);
nand U12771 (N_12771,N_11159,N_11966);
or U12772 (N_12772,N_11825,N_11409);
nand U12773 (N_12773,N_11918,N_11205);
xnor U12774 (N_12774,N_11140,N_11610);
or U12775 (N_12775,N_11272,N_11088);
or U12776 (N_12776,N_11659,N_11270);
xor U12777 (N_12777,N_11001,N_11089);
xor U12778 (N_12778,N_11795,N_11232);
or U12779 (N_12779,N_11043,N_11779);
or U12780 (N_12780,N_11936,N_11481);
xor U12781 (N_12781,N_11435,N_11508);
and U12782 (N_12782,N_11388,N_11172);
nor U12783 (N_12783,N_11891,N_11729);
nor U12784 (N_12784,N_11231,N_11526);
xnor U12785 (N_12785,N_11002,N_11800);
and U12786 (N_12786,N_11549,N_11394);
xor U12787 (N_12787,N_11407,N_11574);
and U12788 (N_12788,N_11170,N_11337);
xor U12789 (N_12789,N_11496,N_11747);
nand U12790 (N_12790,N_11421,N_11150);
and U12791 (N_12791,N_11990,N_11008);
xor U12792 (N_12792,N_11148,N_11950);
nor U12793 (N_12793,N_11892,N_11801);
nor U12794 (N_12794,N_11460,N_11806);
or U12795 (N_12795,N_11096,N_11852);
xor U12796 (N_12796,N_11749,N_11391);
nand U12797 (N_12797,N_11223,N_11349);
nand U12798 (N_12798,N_11588,N_11399);
nor U12799 (N_12799,N_11350,N_11868);
xor U12800 (N_12800,N_11932,N_11394);
and U12801 (N_12801,N_11840,N_11345);
and U12802 (N_12802,N_11587,N_11993);
nand U12803 (N_12803,N_11363,N_11204);
nor U12804 (N_12804,N_11485,N_11532);
nor U12805 (N_12805,N_11445,N_11596);
xor U12806 (N_12806,N_11944,N_11787);
and U12807 (N_12807,N_11602,N_11834);
nor U12808 (N_12808,N_11451,N_11910);
or U12809 (N_12809,N_11787,N_11731);
nand U12810 (N_12810,N_11470,N_11856);
or U12811 (N_12811,N_11026,N_11103);
xnor U12812 (N_12812,N_11259,N_11458);
or U12813 (N_12813,N_11987,N_11328);
and U12814 (N_12814,N_11452,N_11892);
and U12815 (N_12815,N_11365,N_11991);
nand U12816 (N_12816,N_11722,N_11136);
or U12817 (N_12817,N_11679,N_11148);
nand U12818 (N_12818,N_11980,N_11116);
and U12819 (N_12819,N_11511,N_11447);
xor U12820 (N_12820,N_11711,N_11517);
and U12821 (N_12821,N_11384,N_11610);
nand U12822 (N_12822,N_11343,N_11112);
xnor U12823 (N_12823,N_11587,N_11974);
nand U12824 (N_12824,N_11310,N_11937);
nand U12825 (N_12825,N_11511,N_11697);
nor U12826 (N_12826,N_11069,N_11028);
xor U12827 (N_12827,N_11622,N_11443);
or U12828 (N_12828,N_11945,N_11040);
and U12829 (N_12829,N_11944,N_11376);
nand U12830 (N_12830,N_11457,N_11027);
nand U12831 (N_12831,N_11579,N_11786);
or U12832 (N_12832,N_11549,N_11113);
nor U12833 (N_12833,N_11735,N_11514);
xor U12834 (N_12834,N_11549,N_11146);
nor U12835 (N_12835,N_11344,N_11649);
or U12836 (N_12836,N_11624,N_11435);
xor U12837 (N_12837,N_11325,N_11441);
nand U12838 (N_12838,N_11401,N_11951);
nor U12839 (N_12839,N_11522,N_11040);
and U12840 (N_12840,N_11378,N_11173);
or U12841 (N_12841,N_11400,N_11066);
nor U12842 (N_12842,N_11530,N_11731);
xnor U12843 (N_12843,N_11610,N_11669);
nand U12844 (N_12844,N_11542,N_11816);
xor U12845 (N_12845,N_11411,N_11162);
or U12846 (N_12846,N_11933,N_11645);
or U12847 (N_12847,N_11615,N_11934);
nand U12848 (N_12848,N_11546,N_11743);
or U12849 (N_12849,N_11028,N_11496);
or U12850 (N_12850,N_11065,N_11700);
nor U12851 (N_12851,N_11042,N_11518);
nor U12852 (N_12852,N_11780,N_11895);
nand U12853 (N_12853,N_11253,N_11156);
or U12854 (N_12854,N_11314,N_11156);
and U12855 (N_12855,N_11039,N_11043);
nor U12856 (N_12856,N_11343,N_11582);
xnor U12857 (N_12857,N_11781,N_11437);
or U12858 (N_12858,N_11699,N_11435);
nor U12859 (N_12859,N_11205,N_11347);
nand U12860 (N_12860,N_11926,N_11265);
and U12861 (N_12861,N_11319,N_11504);
and U12862 (N_12862,N_11933,N_11871);
nor U12863 (N_12863,N_11116,N_11813);
xor U12864 (N_12864,N_11216,N_11843);
xnor U12865 (N_12865,N_11335,N_11622);
xnor U12866 (N_12866,N_11005,N_11946);
and U12867 (N_12867,N_11469,N_11313);
nor U12868 (N_12868,N_11618,N_11719);
nor U12869 (N_12869,N_11429,N_11577);
nand U12870 (N_12870,N_11646,N_11482);
and U12871 (N_12871,N_11236,N_11358);
nor U12872 (N_12872,N_11102,N_11397);
nor U12873 (N_12873,N_11178,N_11302);
nor U12874 (N_12874,N_11600,N_11070);
and U12875 (N_12875,N_11805,N_11656);
or U12876 (N_12876,N_11005,N_11547);
nand U12877 (N_12877,N_11499,N_11644);
nor U12878 (N_12878,N_11257,N_11656);
xor U12879 (N_12879,N_11574,N_11097);
xnor U12880 (N_12880,N_11133,N_11501);
nand U12881 (N_12881,N_11672,N_11885);
and U12882 (N_12882,N_11575,N_11567);
or U12883 (N_12883,N_11043,N_11406);
or U12884 (N_12884,N_11040,N_11131);
and U12885 (N_12885,N_11833,N_11126);
nand U12886 (N_12886,N_11692,N_11618);
or U12887 (N_12887,N_11045,N_11412);
nor U12888 (N_12888,N_11256,N_11186);
nand U12889 (N_12889,N_11071,N_11738);
nand U12890 (N_12890,N_11071,N_11885);
and U12891 (N_12891,N_11289,N_11528);
and U12892 (N_12892,N_11757,N_11245);
or U12893 (N_12893,N_11533,N_11669);
or U12894 (N_12894,N_11717,N_11069);
and U12895 (N_12895,N_11421,N_11783);
xnor U12896 (N_12896,N_11974,N_11868);
and U12897 (N_12897,N_11052,N_11742);
xnor U12898 (N_12898,N_11182,N_11564);
nand U12899 (N_12899,N_11328,N_11911);
or U12900 (N_12900,N_11782,N_11462);
nand U12901 (N_12901,N_11730,N_11931);
or U12902 (N_12902,N_11199,N_11305);
and U12903 (N_12903,N_11694,N_11386);
nor U12904 (N_12904,N_11907,N_11929);
xnor U12905 (N_12905,N_11320,N_11092);
xor U12906 (N_12906,N_11437,N_11016);
and U12907 (N_12907,N_11805,N_11356);
nor U12908 (N_12908,N_11816,N_11848);
and U12909 (N_12909,N_11116,N_11800);
xnor U12910 (N_12910,N_11817,N_11860);
xor U12911 (N_12911,N_11888,N_11984);
nor U12912 (N_12912,N_11183,N_11005);
or U12913 (N_12913,N_11073,N_11786);
xor U12914 (N_12914,N_11635,N_11027);
nand U12915 (N_12915,N_11631,N_11865);
or U12916 (N_12916,N_11170,N_11426);
nand U12917 (N_12917,N_11929,N_11656);
or U12918 (N_12918,N_11459,N_11540);
xnor U12919 (N_12919,N_11533,N_11239);
nand U12920 (N_12920,N_11721,N_11500);
and U12921 (N_12921,N_11185,N_11256);
or U12922 (N_12922,N_11747,N_11339);
nand U12923 (N_12923,N_11756,N_11712);
nand U12924 (N_12924,N_11109,N_11611);
nand U12925 (N_12925,N_11703,N_11940);
nor U12926 (N_12926,N_11873,N_11116);
or U12927 (N_12927,N_11044,N_11107);
nand U12928 (N_12928,N_11494,N_11650);
and U12929 (N_12929,N_11581,N_11330);
xor U12930 (N_12930,N_11574,N_11626);
nor U12931 (N_12931,N_11162,N_11847);
nor U12932 (N_12932,N_11012,N_11610);
nand U12933 (N_12933,N_11239,N_11553);
nand U12934 (N_12934,N_11238,N_11959);
xor U12935 (N_12935,N_11391,N_11070);
nor U12936 (N_12936,N_11540,N_11562);
xor U12937 (N_12937,N_11650,N_11232);
xor U12938 (N_12938,N_11345,N_11866);
xnor U12939 (N_12939,N_11407,N_11050);
nor U12940 (N_12940,N_11180,N_11436);
and U12941 (N_12941,N_11479,N_11475);
xor U12942 (N_12942,N_11630,N_11495);
or U12943 (N_12943,N_11516,N_11759);
and U12944 (N_12944,N_11804,N_11045);
nor U12945 (N_12945,N_11217,N_11270);
or U12946 (N_12946,N_11840,N_11036);
nor U12947 (N_12947,N_11459,N_11555);
nand U12948 (N_12948,N_11051,N_11313);
and U12949 (N_12949,N_11482,N_11287);
nor U12950 (N_12950,N_11131,N_11743);
nor U12951 (N_12951,N_11130,N_11451);
or U12952 (N_12952,N_11381,N_11020);
xor U12953 (N_12953,N_11364,N_11766);
and U12954 (N_12954,N_11245,N_11617);
or U12955 (N_12955,N_11536,N_11696);
and U12956 (N_12956,N_11680,N_11577);
xnor U12957 (N_12957,N_11080,N_11236);
xor U12958 (N_12958,N_11101,N_11706);
and U12959 (N_12959,N_11158,N_11971);
xor U12960 (N_12960,N_11826,N_11012);
nand U12961 (N_12961,N_11824,N_11541);
and U12962 (N_12962,N_11533,N_11497);
xor U12963 (N_12963,N_11973,N_11922);
or U12964 (N_12964,N_11744,N_11276);
and U12965 (N_12965,N_11711,N_11003);
or U12966 (N_12966,N_11589,N_11942);
nor U12967 (N_12967,N_11976,N_11568);
nor U12968 (N_12968,N_11750,N_11534);
and U12969 (N_12969,N_11548,N_11814);
xor U12970 (N_12970,N_11913,N_11839);
and U12971 (N_12971,N_11800,N_11848);
and U12972 (N_12972,N_11753,N_11546);
or U12973 (N_12973,N_11509,N_11632);
or U12974 (N_12974,N_11606,N_11018);
or U12975 (N_12975,N_11615,N_11139);
nor U12976 (N_12976,N_11443,N_11922);
nand U12977 (N_12977,N_11724,N_11175);
xor U12978 (N_12978,N_11084,N_11759);
and U12979 (N_12979,N_11491,N_11714);
nand U12980 (N_12980,N_11089,N_11615);
nand U12981 (N_12981,N_11803,N_11235);
xor U12982 (N_12982,N_11073,N_11613);
nor U12983 (N_12983,N_11072,N_11951);
nand U12984 (N_12984,N_11168,N_11586);
xnor U12985 (N_12985,N_11840,N_11308);
nand U12986 (N_12986,N_11978,N_11138);
and U12987 (N_12987,N_11242,N_11514);
xor U12988 (N_12988,N_11319,N_11386);
xnor U12989 (N_12989,N_11802,N_11969);
and U12990 (N_12990,N_11665,N_11230);
xor U12991 (N_12991,N_11223,N_11423);
nand U12992 (N_12992,N_11088,N_11853);
and U12993 (N_12993,N_11165,N_11205);
or U12994 (N_12994,N_11614,N_11031);
nand U12995 (N_12995,N_11366,N_11914);
and U12996 (N_12996,N_11720,N_11328);
nor U12997 (N_12997,N_11192,N_11123);
or U12998 (N_12998,N_11505,N_11287);
nor U12999 (N_12999,N_11917,N_11270);
xor U13000 (N_13000,N_12663,N_12591);
nand U13001 (N_13001,N_12737,N_12958);
nor U13002 (N_13002,N_12478,N_12651);
nor U13003 (N_13003,N_12360,N_12963);
and U13004 (N_13004,N_12610,N_12519);
nand U13005 (N_13005,N_12893,N_12265);
xor U13006 (N_13006,N_12130,N_12144);
nand U13007 (N_13007,N_12169,N_12861);
and U13008 (N_13008,N_12106,N_12939);
nor U13009 (N_13009,N_12086,N_12454);
and U13010 (N_13010,N_12906,N_12312);
xnor U13011 (N_13011,N_12033,N_12921);
or U13012 (N_13012,N_12804,N_12596);
and U13013 (N_13013,N_12530,N_12681);
or U13014 (N_13014,N_12296,N_12287);
and U13015 (N_13015,N_12697,N_12606);
nand U13016 (N_13016,N_12516,N_12167);
nor U13017 (N_13017,N_12676,N_12231);
nand U13018 (N_13018,N_12288,N_12303);
and U13019 (N_13019,N_12613,N_12497);
nand U13020 (N_13020,N_12334,N_12262);
or U13021 (N_13021,N_12221,N_12081);
xor U13022 (N_13022,N_12194,N_12255);
xor U13023 (N_13023,N_12246,N_12784);
and U13024 (N_13024,N_12222,N_12878);
xor U13025 (N_13025,N_12896,N_12252);
and U13026 (N_13026,N_12064,N_12514);
xnor U13027 (N_13027,N_12439,N_12585);
nand U13028 (N_13028,N_12152,N_12306);
xor U13029 (N_13029,N_12540,N_12362);
nand U13030 (N_13030,N_12616,N_12286);
xnor U13031 (N_13031,N_12348,N_12976);
and U13032 (N_13032,N_12128,N_12155);
xor U13033 (N_13033,N_12739,N_12382);
xnor U13034 (N_13034,N_12575,N_12201);
and U13035 (N_13035,N_12883,N_12153);
or U13036 (N_13036,N_12293,N_12176);
and U13037 (N_13037,N_12627,N_12234);
nor U13038 (N_13038,N_12354,N_12694);
or U13039 (N_13039,N_12502,N_12846);
nand U13040 (N_13040,N_12714,N_12538);
xor U13041 (N_13041,N_12477,N_12609);
or U13042 (N_13042,N_12931,N_12586);
xnor U13043 (N_13043,N_12007,N_12436);
xnor U13044 (N_13044,N_12188,N_12889);
and U13045 (N_13045,N_12970,N_12561);
and U13046 (N_13046,N_12603,N_12196);
and U13047 (N_13047,N_12617,N_12839);
and U13048 (N_13048,N_12433,N_12527);
xnor U13049 (N_13049,N_12365,N_12473);
or U13050 (N_13050,N_12395,N_12206);
nor U13051 (N_13051,N_12203,N_12829);
or U13052 (N_13052,N_12393,N_12699);
and U13053 (N_13053,N_12825,N_12069);
xnor U13054 (N_13054,N_12767,N_12210);
and U13055 (N_13055,N_12202,N_12971);
nor U13056 (N_13056,N_12499,N_12453);
xnor U13057 (N_13057,N_12189,N_12353);
nor U13058 (N_13058,N_12728,N_12523);
and U13059 (N_13059,N_12571,N_12492);
nand U13060 (N_13060,N_12930,N_12845);
nor U13061 (N_13061,N_12109,N_12529);
and U13062 (N_13062,N_12779,N_12567);
and U13063 (N_13063,N_12133,N_12823);
or U13064 (N_13064,N_12619,N_12813);
nor U13065 (N_13065,N_12378,N_12107);
or U13066 (N_13066,N_12991,N_12216);
or U13067 (N_13067,N_12654,N_12281);
nor U13068 (N_13068,N_12464,N_12413);
nor U13069 (N_13069,N_12815,N_12257);
and U13070 (N_13070,N_12226,N_12355);
or U13071 (N_13071,N_12366,N_12863);
nand U13072 (N_13072,N_12675,N_12914);
xor U13073 (N_13073,N_12770,N_12483);
nor U13074 (N_13074,N_12981,N_12505);
and U13075 (N_13075,N_12099,N_12230);
nor U13076 (N_13076,N_12294,N_12451);
and U13077 (N_13077,N_12667,N_12199);
nand U13078 (N_13078,N_12219,N_12756);
and U13079 (N_13079,N_12092,N_12562);
xnor U13080 (N_13080,N_12638,N_12072);
xnor U13081 (N_13081,N_12810,N_12361);
nand U13082 (N_13082,N_12791,N_12503);
or U13083 (N_13083,N_12763,N_12108);
nand U13084 (N_13084,N_12052,N_12611);
nor U13085 (N_13085,N_12649,N_12398);
nor U13086 (N_13086,N_12013,N_12924);
nor U13087 (N_13087,N_12993,N_12666);
or U13088 (N_13088,N_12768,N_12305);
xor U13089 (N_13089,N_12528,N_12005);
nor U13090 (N_13090,N_12866,N_12200);
nand U13091 (N_13091,N_12386,N_12336);
or U13092 (N_13092,N_12175,N_12875);
and U13093 (N_13093,N_12022,N_12549);
and U13094 (N_13094,N_12449,N_12380);
xor U13095 (N_13095,N_12693,N_12040);
or U13096 (N_13096,N_12215,N_12351);
or U13097 (N_13097,N_12817,N_12882);
nand U13098 (N_13098,N_12036,N_12080);
nor U13099 (N_13099,N_12788,N_12588);
nand U13100 (N_13100,N_12070,N_12909);
or U13101 (N_13101,N_12626,N_12946);
or U13102 (N_13102,N_12542,N_12570);
xnor U13103 (N_13103,N_12911,N_12011);
or U13104 (N_13104,N_12310,N_12724);
nor U13105 (N_13105,N_12669,N_12923);
and U13106 (N_13106,N_12781,N_12487);
xnor U13107 (N_13107,N_12044,N_12753);
nand U13108 (N_13108,N_12233,N_12488);
xnor U13109 (N_13109,N_12750,N_12621);
xor U13110 (N_13110,N_12998,N_12122);
nor U13111 (N_13111,N_12706,N_12038);
and U13112 (N_13112,N_12146,N_12683);
nand U13113 (N_13113,N_12479,N_12665);
nor U13114 (N_13114,N_12860,N_12944);
nand U13115 (N_13115,N_12560,N_12096);
or U13116 (N_13116,N_12237,N_12115);
and U13117 (N_13117,N_12029,N_12847);
xnor U13118 (N_13118,N_12389,N_12733);
nor U13119 (N_13119,N_12299,N_12563);
nor U13120 (N_13120,N_12006,N_12557);
and U13121 (N_13121,N_12648,N_12954);
nor U13122 (N_13122,N_12774,N_12445);
and U13123 (N_13123,N_12148,N_12668);
and U13124 (N_13124,N_12541,N_12264);
nand U13125 (N_13125,N_12712,N_12343);
nor U13126 (N_13126,N_12721,N_12960);
and U13127 (N_13127,N_12652,N_12061);
or U13128 (N_13128,N_12656,N_12873);
nand U13129 (N_13129,N_12719,N_12165);
xnor U13130 (N_13130,N_12597,N_12495);
and U13131 (N_13131,N_12513,N_12994);
nand U13132 (N_13132,N_12715,N_12802);
nand U13133 (N_13133,N_12278,N_12865);
nand U13134 (N_13134,N_12761,N_12301);
and U13135 (N_13135,N_12441,N_12383);
nand U13136 (N_13136,N_12021,N_12874);
and U13137 (N_13137,N_12250,N_12397);
nor U13138 (N_13138,N_12496,N_12256);
nor U13139 (N_13139,N_12997,N_12512);
xor U13140 (N_13140,N_12127,N_12291);
xnor U13141 (N_13141,N_12213,N_12880);
or U13142 (N_13142,N_12412,N_12717);
nand U13143 (N_13143,N_12628,N_12251);
nand U13144 (N_13144,N_12455,N_12766);
or U13145 (N_13145,N_12826,N_12953);
nor U13146 (N_13146,N_12996,N_12579);
and U13147 (N_13147,N_12375,N_12664);
xor U13148 (N_13148,N_12138,N_12701);
and U13149 (N_13149,N_12623,N_12722);
nor U13150 (N_13150,N_12536,N_12735);
nand U13151 (N_13151,N_12438,N_12025);
nand U13152 (N_13152,N_12710,N_12999);
or U13153 (N_13153,N_12275,N_12049);
or U13154 (N_13154,N_12869,N_12493);
nor U13155 (N_13155,N_12684,N_12045);
nor U13156 (N_13156,N_12647,N_12458);
nor U13157 (N_13157,N_12983,N_12187);
or U13158 (N_13158,N_12595,N_12332);
nand U13159 (N_13159,N_12419,N_12026);
and U13160 (N_13160,N_12709,N_12481);
xor U13161 (N_13161,N_12749,N_12401);
nor U13162 (N_13162,N_12437,N_12908);
or U13163 (N_13163,N_12000,N_12211);
or U13164 (N_13164,N_12593,N_12088);
nand U13165 (N_13165,N_12898,N_12381);
and U13166 (N_13166,N_12129,N_12918);
or U13167 (N_13167,N_12474,N_12225);
and U13168 (N_13168,N_12708,N_12313);
and U13169 (N_13169,N_12830,N_12121);
or U13170 (N_13170,N_12282,N_12720);
and U13171 (N_13171,N_12407,N_12622);
or U13172 (N_13172,N_12420,N_12024);
nor U13173 (N_13173,N_12772,N_12677);
and U13174 (N_13174,N_12066,N_12434);
nand U13175 (N_13175,N_12460,N_12832);
nor U13176 (N_13176,N_12035,N_12387);
and U13177 (N_13177,N_12390,N_12317);
nor U13178 (N_13178,N_12131,N_12309);
xor U13179 (N_13179,N_12682,N_12157);
and U13180 (N_13180,N_12082,N_12158);
xor U13181 (N_13181,N_12102,N_12746);
or U13182 (N_13182,N_12764,N_12110);
nor U13183 (N_13183,N_12584,N_12053);
or U13184 (N_13184,N_12820,N_12349);
and U13185 (N_13185,N_12871,N_12634);
and U13186 (N_13186,N_12164,N_12848);
or U13187 (N_13187,N_12058,N_12150);
and U13188 (N_13188,N_12903,N_12633);
nand U13189 (N_13189,N_12602,N_12039);
and U13190 (N_13190,N_12576,N_12030);
nor U13191 (N_13191,N_12073,N_12448);
or U13192 (N_13192,N_12253,N_12227);
nor U13193 (N_13193,N_12950,N_12350);
and U13194 (N_13194,N_12261,N_12339);
or U13195 (N_13195,N_12104,N_12941);
or U13196 (N_13196,N_12229,N_12247);
nand U13197 (N_13197,N_12819,N_12489);
and U13198 (N_13198,N_12320,N_12808);
nand U13199 (N_13199,N_12377,N_12010);
or U13200 (N_13200,N_12639,N_12315);
and U13201 (N_13201,N_12945,N_12142);
xnor U13202 (N_13202,N_12014,N_12811);
nand U13203 (N_13203,N_12446,N_12966);
nand U13204 (N_13204,N_12969,N_12469);
nand U13205 (N_13205,N_12224,N_12004);
and U13206 (N_13206,N_12032,N_12744);
xor U13207 (N_13207,N_12711,N_12019);
or U13208 (N_13208,N_12145,N_12653);
or U13209 (N_13209,N_12244,N_12457);
or U13210 (N_13210,N_12485,N_12316);
or U13211 (N_13211,N_12057,N_12872);
nand U13212 (N_13212,N_12841,N_12618);
or U13213 (N_13213,N_12300,N_12640);
or U13214 (N_13214,N_12867,N_12174);
or U13215 (N_13215,N_12589,N_12968);
nand U13216 (N_13216,N_12195,N_12192);
or U13217 (N_13217,N_12017,N_12927);
nand U13218 (N_13218,N_12472,N_12135);
and U13219 (N_13219,N_12283,N_12027);
nor U13220 (N_13220,N_12123,N_12277);
and U13221 (N_13221,N_12431,N_12156);
nor U13222 (N_13222,N_12426,N_12417);
nand U13223 (N_13223,N_12120,N_12577);
and U13224 (N_13224,N_12179,N_12323);
xnor U13225 (N_13225,N_12442,N_12661);
nand U13226 (N_13226,N_12427,N_12337);
and U13227 (N_13227,N_12091,N_12751);
or U13228 (N_13228,N_12543,N_12854);
nor U13229 (N_13229,N_12636,N_12974);
or U13230 (N_13230,N_12740,N_12447);
nand U13231 (N_13231,N_12548,N_12624);
and U13232 (N_13232,N_12394,N_12228);
xor U13233 (N_13233,N_12552,N_12553);
or U13234 (N_13234,N_12868,N_12556);
nor U13235 (N_13235,N_12186,N_12786);
nand U13236 (N_13236,N_12385,N_12738);
nor U13237 (N_13237,N_12992,N_12116);
and U13238 (N_13238,N_12776,N_12347);
and U13239 (N_13239,N_12800,N_12071);
xnor U13240 (N_13240,N_12748,N_12391);
and U13241 (N_13241,N_12978,N_12322);
xnor U13242 (N_13242,N_12185,N_12973);
nor U13243 (N_13243,N_12703,N_12181);
xor U13244 (N_13244,N_12218,N_12059);
nor U13245 (N_13245,N_12578,N_12657);
or U13246 (N_13246,N_12067,N_12330);
nand U13247 (N_13247,N_12799,N_12159);
xnor U13248 (N_13248,N_12463,N_12484);
nand U13249 (N_13249,N_12023,N_12644);
or U13250 (N_13250,N_12198,N_12698);
or U13251 (N_13251,N_12405,N_12270);
nand U13252 (N_13252,N_12835,N_12468);
nand U13253 (N_13253,N_12702,N_12335);
nand U13254 (N_13254,N_12151,N_12078);
xor U13255 (N_13255,N_12111,N_12979);
nand U13256 (N_13256,N_12965,N_12525);
nor U13257 (N_13257,N_12807,N_12614);
xor U13258 (N_13258,N_12134,N_12725);
nand U13259 (N_13259,N_12635,N_12881);
xor U13260 (N_13260,N_12295,N_12690);
nand U13261 (N_13261,N_12331,N_12885);
and U13262 (N_13262,N_12857,N_12328);
xnor U13263 (N_13263,N_12118,N_12384);
xnor U13264 (N_13264,N_12902,N_12777);
nand U13265 (N_13265,N_12459,N_12402);
and U13266 (N_13266,N_12732,N_12704);
and U13267 (N_13267,N_12239,N_12430);
or U13268 (N_13268,N_12569,N_12778);
xor U13269 (N_13269,N_12147,N_12173);
or U13270 (N_13270,N_12340,N_12894);
xor U13271 (N_13271,N_12601,N_12506);
and U13272 (N_13272,N_12047,N_12191);
nand U13273 (N_13273,N_12090,N_12510);
and U13274 (N_13274,N_12787,N_12934);
or U13275 (N_13275,N_12897,N_12679);
xor U13276 (N_13276,N_12163,N_12041);
or U13277 (N_13277,N_12550,N_12289);
nand U13278 (N_13278,N_12988,N_12856);
or U13279 (N_13279,N_12539,N_12342);
nand U13280 (N_13280,N_12522,N_12670);
or U13281 (N_13281,N_12326,N_12055);
or U13282 (N_13282,N_12094,N_12743);
xnor U13283 (N_13283,N_12853,N_12048);
xnor U13284 (N_13284,N_12285,N_12357);
and U13285 (N_13285,N_12031,N_12471);
nor U13286 (N_13286,N_12718,N_12678);
xnor U13287 (N_13287,N_12432,N_12917);
nor U13288 (N_13288,N_12534,N_12139);
nor U13289 (N_13289,N_12009,N_12170);
and U13290 (N_13290,N_12223,N_12915);
or U13291 (N_13291,N_12076,N_12374);
xor U13292 (N_13292,N_12642,N_12598);
xor U13293 (N_13293,N_12132,N_12183);
nor U13294 (N_13294,N_12922,N_12916);
nor U13295 (N_13295,N_12535,N_12824);
nand U13296 (N_13296,N_12892,N_12491);
nand U13297 (N_13297,N_12314,N_12212);
nor U13298 (N_13298,N_12920,N_12271);
xor U13299 (N_13299,N_12190,N_12424);
and U13300 (N_13300,N_12466,N_12925);
nand U13301 (N_13301,N_12079,N_12637);
nand U13302 (N_13302,N_12759,N_12537);
nor U13303 (N_13303,N_12870,N_12809);
nor U13304 (N_13304,N_12700,N_12904);
nand U13305 (N_13305,N_12905,N_12369);
and U13306 (N_13306,N_12117,N_12773);
nor U13307 (N_13307,N_12632,N_12936);
nor U13308 (N_13308,N_12643,N_12242);
xor U13309 (N_13309,N_12172,N_12259);
xor U13310 (N_13310,N_12864,N_12838);
and U13311 (N_13311,N_12051,N_12985);
xor U13312 (N_13312,N_12604,N_12370);
xnor U13313 (N_13313,N_12308,N_12028);
xnor U13314 (N_13314,N_12594,N_12008);
xnor U13315 (N_13315,N_12957,N_12077);
nor U13316 (N_13316,N_12607,N_12416);
and U13317 (N_13317,N_12204,N_12418);
nand U13318 (N_13318,N_12042,N_12359);
xor U13319 (N_13319,N_12141,N_12599);
nor U13320 (N_13320,N_12517,N_12947);
xnor U13321 (N_13321,N_12605,N_12758);
or U13322 (N_13322,N_12180,N_12363);
nand U13323 (N_13323,N_12450,N_12741);
nand U13324 (N_13324,N_12161,N_12975);
xor U13325 (N_13325,N_12197,N_12232);
xor U13326 (N_13326,N_12425,N_12840);
xor U13327 (N_13327,N_12429,N_12659);
or U13328 (N_13328,N_12100,N_12646);
and U13329 (N_13329,N_12818,N_12267);
or U13330 (N_13330,N_12687,N_12625);
nor U13331 (N_13331,N_12440,N_12280);
nand U13332 (N_13332,N_12964,N_12327);
xnor U13333 (N_13333,N_12184,N_12736);
nand U13334 (N_13334,N_12695,N_12943);
nor U13335 (N_13335,N_12403,N_12855);
nand U13336 (N_13336,N_12093,N_12089);
nor U13337 (N_13337,N_12980,N_12166);
nor U13338 (N_13338,N_12119,N_12790);
nand U13339 (N_13339,N_12843,N_12012);
xor U13340 (N_13340,N_12063,N_12726);
or U13341 (N_13341,N_12087,N_12559);
and U13342 (N_13342,N_12368,N_12956);
nand U13343 (N_13343,N_12731,N_12062);
nor U13344 (N_13344,N_12962,N_12895);
xor U13345 (N_13345,N_12302,N_12933);
nand U13346 (N_13346,N_12546,N_12050);
xor U13347 (N_13347,N_12849,N_12480);
xor U13348 (N_13348,N_12494,N_12399);
or U13349 (N_13349,N_12124,N_12423);
nand U13350 (N_13350,N_12243,N_12928);
or U13351 (N_13351,N_12113,N_12177);
and U13352 (N_13352,N_12645,N_12400);
xnor U13353 (N_13353,N_12762,N_12713);
and U13354 (N_13354,N_12730,N_12580);
nand U13355 (N_13355,N_12490,N_12511);
nand U13356 (N_13356,N_12796,N_12046);
nand U13357 (N_13357,N_12344,N_12886);
xor U13358 (N_13358,N_12125,N_12723);
or U13359 (N_13359,N_12373,N_12707);
nor U13360 (N_13360,N_12411,N_12408);
and U13361 (N_13361,N_12752,N_12798);
xnor U13362 (N_13362,N_12112,N_12178);
nor U13363 (N_13363,N_12162,N_12097);
xor U13364 (N_13364,N_12615,N_12533);
nand U13365 (N_13365,N_12620,N_12140);
and U13366 (N_13366,N_12217,N_12572);
xnor U13367 (N_13367,N_12887,N_12565);
or U13368 (N_13368,N_12987,N_12745);
nor U13369 (N_13369,N_12755,N_12955);
and U13370 (N_13370,N_12900,N_12075);
xnor U13371 (N_13371,N_12105,N_12236);
nor U13372 (N_13372,N_12443,N_12074);
nand U13373 (N_13373,N_12065,N_12590);
xnor U13374 (N_13374,N_12241,N_12673);
xor U13375 (N_13375,N_12806,N_12269);
or U13376 (N_13376,N_12901,N_12182);
and U13377 (N_13377,N_12587,N_12816);
and U13378 (N_13378,N_12414,N_12558);
nand U13379 (N_13379,N_12521,N_12345);
or U13380 (N_13380,N_12805,N_12783);
or U13381 (N_13381,N_12114,N_12456);
xor U13382 (N_13382,N_12812,N_12691);
nor U13383 (N_13383,N_12476,N_12338);
or U13384 (N_13384,N_12333,N_12899);
xor U13385 (N_13385,N_12003,N_12307);
xnor U13386 (N_13386,N_12043,N_12850);
and U13387 (N_13387,N_12154,N_12890);
nor U13388 (N_13388,N_12524,N_12937);
nand U13389 (N_13389,N_12951,N_12566);
nor U13390 (N_13390,N_12068,N_12801);
nor U13391 (N_13391,N_12465,N_12467);
or U13392 (N_13392,N_12422,N_12324);
and U13393 (N_13393,N_12245,N_12919);
xor U13394 (N_13394,N_12568,N_12083);
or U13395 (N_13395,N_12742,N_12298);
and U13396 (N_13396,N_12470,N_12461);
and U13397 (N_13397,N_12515,N_12103);
or U13398 (N_13398,N_12268,N_12990);
and U13399 (N_13399,N_12989,N_12272);
or U13400 (N_13400,N_12220,N_12564);
xor U13401 (N_13401,N_12935,N_12573);
xnor U13402 (N_13402,N_12891,N_12034);
xor U13403 (N_13403,N_12612,N_12462);
or U13404 (N_13404,N_12160,N_12016);
nand U13405 (N_13405,N_12207,N_12780);
xnor U13406 (N_13406,N_12716,N_12977);
or U13407 (N_13407,N_12392,N_12747);
and U13408 (N_13408,N_12508,N_12085);
and U13409 (N_13409,N_12782,N_12814);
xnor U13410 (N_13410,N_12238,N_12952);
nand U13411 (N_13411,N_12101,N_12696);
and U13412 (N_13412,N_12325,N_12658);
and U13413 (N_13413,N_12608,N_12274);
xor U13414 (N_13414,N_12304,N_12765);
nor U13415 (N_13415,N_12851,N_12193);
or U13416 (N_13416,N_12292,N_12932);
or U13417 (N_13417,N_12692,N_12240);
xnor U13418 (N_13418,N_12982,N_12674);
or U13419 (N_13419,N_12396,N_12406);
and U13420 (N_13420,N_12171,N_12641);
or U13421 (N_13421,N_12942,N_12926);
nand U13422 (N_13422,N_12020,N_12388);
xnor U13423 (N_13423,N_12143,N_12876);
nand U13424 (N_13424,N_12600,N_12822);
xnor U13425 (N_13425,N_12948,N_12002);
nor U13426 (N_13426,N_12486,N_12544);
and U13427 (N_13427,N_12266,N_12907);
nand U13428 (N_13428,N_12168,N_12862);
nand U13429 (N_13429,N_12888,N_12910);
xnor U13430 (N_13430,N_12831,N_12015);
nand U13431 (N_13431,N_12545,N_12311);
nand U13432 (N_13432,N_12341,N_12631);
nor U13433 (N_13433,N_12321,N_12792);
nor U13434 (N_13434,N_12098,N_12984);
xor U13435 (N_13435,N_12581,N_12364);
nand U13436 (N_13436,N_12208,N_12526);
nand U13437 (N_13437,N_12249,N_12518);
or U13438 (N_13438,N_12771,N_12555);
nor U13439 (N_13439,N_12452,N_12444);
nand U13440 (N_13440,N_12729,N_12279);
or U13441 (N_13441,N_12263,N_12273);
and U13442 (N_13442,N_12879,N_12757);
xnor U13443 (N_13443,N_12037,N_12972);
xor U13444 (N_13444,N_12428,N_12769);
or U13445 (N_13445,N_12794,N_12680);
nand U13446 (N_13446,N_12689,N_12372);
xor U13447 (N_13447,N_12410,N_12940);
xnor U13448 (N_13448,N_12507,N_12318);
or U13449 (N_13449,N_12660,N_12912);
xnor U13450 (N_13450,N_12504,N_12376);
nor U13451 (N_13451,N_12126,N_12379);
nand U13452 (N_13452,N_12842,N_12986);
and U13453 (N_13453,N_12859,N_12475);
nor U13454 (N_13454,N_12551,N_12959);
or U13455 (N_13455,N_12662,N_12629);
xor U13456 (N_13456,N_12554,N_12583);
xor U13457 (N_13457,N_12214,N_12967);
nor U13458 (N_13458,N_12509,N_12501);
and U13459 (N_13459,N_12929,N_12995);
nand U13460 (N_13460,N_12795,N_12001);
or U13461 (N_13461,N_12482,N_12297);
nor U13462 (N_13462,N_12352,N_12803);
and U13463 (N_13463,N_12686,N_12961);
nand U13464 (N_13464,N_12060,N_12520);
nor U13465 (N_13465,N_12435,N_12833);
nor U13466 (N_13466,N_12260,N_12785);
nor U13467 (N_13467,N_12913,N_12258);
nand U13468 (N_13468,N_12404,N_12095);
and U13469 (N_13469,N_12836,N_12734);
xnor U13470 (N_13470,N_12630,N_12018);
nor U13471 (N_13471,N_12084,N_12531);
nand U13472 (N_13472,N_12136,N_12235);
xnor U13473 (N_13473,N_12205,N_12371);
xnor U13474 (N_13474,N_12409,N_12793);
nor U13475 (N_13475,N_12149,N_12828);
and U13476 (N_13476,N_12754,N_12532);
or U13477 (N_13477,N_12290,N_12137);
or U13478 (N_13478,N_12650,N_12284);
nor U13479 (N_13479,N_12844,N_12834);
or U13480 (N_13480,N_12672,N_12837);
or U13481 (N_13481,N_12056,N_12421);
or U13482 (N_13482,N_12329,N_12547);
xnor U13483 (N_13483,N_12884,N_12356);
and U13484 (N_13484,N_12358,N_12949);
nand U13485 (N_13485,N_12688,N_12276);
nand U13486 (N_13486,N_12655,N_12705);
xnor U13487 (N_13487,N_12415,N_12498);
or U13488 (N_13488,N_12582,N_12827);
and U13489 (N_13489,N_12852,N_12319);
or U13490 (N_13490,N_12760,N_12877);
nor U13491 (N_13491,N_12858,N_12574);
and U13492 (N_13492,N_12346,N_12248);
xnor U13493 (N_13493,N_12500,N_12797);
or U13494 (N_13494,N_12789,N_12671);
xor U13495 (N_13495,N_12254,N_12592);
xor U13496 (N_13496,N_12054,N_12821);
and U13497 (N_13497,N_12367,N_12938);
or U13498 (N_13498,N_12209,N_12685);
nand U13499 (N_13499,N_12775,N_12727);
nor U13500 (N_13500,N_12549,N_12485);
and U13501 (N_13501,N_12339,N_12616);
nor U13502 (N_13502,N_12843,N_12625);
or U13503 (N_13503,N_12994,N_12241);
nor U13504 (N_13504,N_12202,N_12510);
xor U13505 (N_13505,N_12687,N_12214);
nor U13506 (N_13506,N_12055,N_12011);
nor U13507 (N_13507,N_12492,N_12689);
or U13508 (N_13508,N_12562,N_12271);
xor U13509 (N_13509,N_12295,N_12775);
nand U13510 (N_13510,N_12431,N_12087);
or U13511 (N_13511,N_12714,N_12049);
or U13512 (N_13512,N_12031,N_12734);
nand U13513 (N_13513,N_12913,N_12683);
and U13514 (N_13514,N_12493,N_12644);
or U13515 (N_13515,N_12736,N_12310);
or U13516 (N_13516,N_12468,N_12148);
xor U13517 (N_13517,N_12328,N_12926);
or U13518 (N_13518,N_12090,N_12152);
nor U13519 (N_13519,N_12546,N_12521);
or U13520 (N_13520,N_12794,N_12427);
nand U13521 (N_13521,N_12354,N_12802);
and U13522 (N_13522,N_12830,N_12763);
nor U13523 (N_13523,N_12786,N_12679);
and U13524 (N_13524,N_12191,N_12163);
or U13525 (N_13525,N_12032,N_12091);
nor U13526 (N_13526,N_12088,N_12544);
nand U13527 (N_13527,N_12184,N_12512);
nor U13528 (N_13528,N_12684,N_12682);
xnor U13529 (N_13529,N_12352,N_12553);
xnor U13530 (N_13530,N_12133,N_12485);
nor U13531 (N_13531,N_12546,N_12010);
nand U13532 (N_13532,N_12663,N_12017);
nand U13533 (N_13533,N_12961,N_12885);
or U13534 (N_13534,N_12532,N_12030);
nand U13535 (N_13535,N_12634,N_12368);
nand U13536 (N_13536,N_12995,N_12591);
nand U13537 (N_13537,N_12270,N_12183);
xnor U13538 (N_13538,N_12536,N_12666);
xnor U13539 (N_13539,N_12365,N_12551);
nand U13540 (N_13540,N_12215,N_12692);
nand U13541 (N_13541,N_12630,N_12830);
nand U13542 (N_13542,N_12542,N_12131);
or U13543 (N_13543,N_12345,N_12168);
nor U13544 (N_13544,N_12689,N_12519);
xnor U13545 (N_13545,N_12814,N_12502);
nor U13546 (N_13546,N_12211,N_12397);
nor U13547 (N_13547,N_12031,N_12129);
and U13548 (N_13548,N_12576,N_12553);
or U13549 (N_13549,N_12512,N_12695);
or U13550 (N_13550,N_12758,N_12733);
nand U13551 (N_13551,N_12340,N_12665);
and U13552 (N_13552,N_12693,N_12775);
or U13553 (N_13553,N_12776,N_12087);
and U13554 (N_13554,N_12195,N_12277);
nand U13555 (N_13555,N_12679,N_12290);
nor U13556 (N_13556,N_12802,N_12168);
nand U13557 (N_13557,N_12860,N_12688);
and U13558 (N_13558,N_12038,N_12151);
nand U13559 (N_13559,N_12453,N_12011);
and U13560 (N_13560,N_12672,N_12338);
nand U13561 (N_13561,N_12068,N_12400);
and U13562 (N_13562,N_12455,N_12204);
nand U13563 (N_13563,N_12107,N_12053);
or U13564 (N_13564,N_12618,N_12495);
or U13565 (N_13565,N_12367,N_12513);
xor U13566 (N_13566,N_12425,N_12972);
and U13567 (N_13567,N_12507,N_12575);
and U13568 (N_13568,N_12230,N_12714);
nor U13569 (N_13569,N_12680,N_12058);
xnor U13570 (N_13570,N_12013,N_12066);
xor U13571 (N_13571,N_12879,N_12492);
nand U13572 (N_13572,N_12984,N_12519);
or U13573 (N_13573,N_12274,N_12887);
nor U13574 (N_13574,N_12912,N_12545);
and U13575 (N_13575,N_12137,N_12274);
and U13576 (N_13576,N_12461,N_12822);
and U13577 (N_13577,N_12001,N_12385);
nor U13578 (N_13578,N_12226,N_12708);
and U13579 (N_13579,N_12985,N_12121);
or U13580 (N_13580,N_12081,N_12147);
and U13581 (N_13581,N_12234,N_12742);
nand U13582 (N_13582,N_12878,N_12774);
and U13583 (N_13583,N_12426,N_12011);
nor U13584 (N_13584,N_12805,N_12084);
nor U13585 (N_13585,N_12498,N_12578);
and U13586 (N_13586,N_12959,N_12628);
xnor U13587 (N_13587,N_12951,N_12617);
xnor U13588 (N_13588,N_12072,N_12141);
and U13589 (N_13589,N_12724,N_12905);
xor U13590 (N_13590,N_12173,N_12180);
xor U13591 (N_13591,N_12673,N_12862);
or U13592 (N_13592,N_12851,N_12488);
nor U13593 (N_13593,N_12278,N_12326);
or U13594 (N_13594,N_12300,N_12145);
and U13595 (N_13595,N_12794,N_12599);
and U13596 (N_13596,N_12753,N_12513);
or U13597 (N_13597,N_12127,N_12265);
nor U13598 (N_13598,N_12095,N_12610);
nor U13599 (N_13599,N_12175,N_12918);
or U13600 (N_13600,N_12166,N_12325);
or U13601 (N_13601,N_12076,N_12003);
and U13602 (N_13602,N_12063,N_12111);
nand U13603 (N_13603,N_12084,N_12108);
nor U13604 (N_13604,N_12184,N_12256);
xnor U13605 (N_13605,N_12706,N_12324);
and U13606 (N_13606,N_12115,N_12825);
or U13607 (N_13607,N_12931,N_12430);
xnor U13608 (N_13608,N_12084,N_12360);
xor U13609 (N_13609,N_12640,N_12437);
nand U13610 (N_13610,N_12161,N_12842);
nand U13611 (N_13611,N_12996,N_12097);
nor U13612 (N_13612,N_12102,N_12496);
nand U13613 (N_13613,N_12188,N_12967);
nor U13614 (N_13614,N_12691,N_12955);
and U13615 (N_13615,N_12892,N_12549);
and U13616 (N_13616,N_12546,N_12437);
xor U13617 (N_13617,N_12051,N_12053);
and U13618 (N_13618,N_12022,N_12337);
and U13619 (N_13619,N_12952,N_12184);
nor U13620 (N_13620,N_12306,N_12170);
or U13621 (N_13621,N_12517,N_12588);
xnor U13622 (N_13622,N_12891,N_12079);
xor U13623 (N_13623,N_12662,N_12401);
nor U13624 (N_13624,N_12794,N_12277);
or U13625 (N_13625,N_12040,N_12661);
xor U13626 (N_13626,N_12545,N_12298);
nor U13627 (N_13627,N_12055,N_12788);
and U13628 (N_13628,N_12467,N_12802);
or U13629 (N_13629,N_12539,N_12858);
xor U13630 (N_13630,N_12305,N_12875);
xnor U13631 (N_13631,N_12072,N_12280);
xor U13632 (N_13632,N_12106,N_12554);
and U13633 (N_13633,N_12763,N_12145);
and U13634 (N_13634,N_12204,N_12522);
nand U13635 (N_13635,N_12814,N_12539);
and U13636 (N_13636,N_12401,N_12548);
or U13637 (N_13637,N_12516,N_12726);
nand U13638 (N_13638,N_12641,N_12940);
and U13639 (N_13639,N_12786,N_12252);
nand U13640 (N_13640,N_12136,N_12979);
or U13641 (N_13641,N_12680,N_12675);
xnor U13642 (N_13642,N_12945,N_12128);
nand U13643 (N_13643,N_12900,N_12505);
and U13644 (N_13644,N_12146,N_12238);
xor U13645 (N_13645,N_12323,N_12668);
nand U13646 (N_13646,N_12086,N_12317);
or U13647 (N_13647,N_12036,N_12122);
nand U13648 (N_13648,N_12862,N_12182);
or U13649 (N_13649,N_12392,N_12687);
nor U13650 (N_13650,N_12845,N_12493);
or U13651 (N_13651,N_12664,N_12314);
or U13652 (N_13652,N_12065,N_12511);
xor U13653 (N_13653,N_12793,N_12651);
nor U13654 (N_13654,N_12574,N_12656);
or U13655 (N_13655,N_12718,N_12162);
nand U13656 (N_13656,N_12740,N_12241);
xnor U13657 (N_13657,N_12557,N_12115);
or U13658 (N_13658,N_12733,N_12789);
or U13659 (N_13659,N_12639,N_12165);
nand U13660 (N_13660,N_12393,N_12623);
and U13661 (N_13661,N_12809,N_12933);
nor U13662 (N_13662,N_12790,N_12334);
or U13663 (N_13663,N_12520,N_12589);
xor U13664 (N_13664,N_12863,N_12153);
or U13665 (N_13665,N_12930,N_12068);
nor U13666 (N_13666,N_12423,N_12896);
or U13667 (N_13667,N_12398,N_12865);
and U13668 (N_13668,N_12128,N_12569);
or U13669 (N_13669,N_12716,N_12161);
or U13670 (N_13670,N_12645,N_12320);
or U13671 (N_13671,N_12292,N_12655);
or U13672 (N_13672,N_12117,N_12229);
or U13673 (N_13673,N_12579,N_12920);
and U13674 (N_13674,N_12561,N_12808);
and U13675 (N_13675,N_12595,N_12215);
xnor U13676 (N_13676,N_12816,N_12193);
and U13677 (N_13677,N_12286,N_12413);
or U13678 (N_13678,N_12589,N_12230);
nand U13679 (N_13679,N_12416,N_12988);
xor U13680 (N_13680,N_12250,N_12770);
nor U13681 (N_13681,N_12150,N_12794);
or U13682 (N_13682,N_12017,N_12485);
nand U13683 (N_13683,N_12190,N_12828);
nor U13684 (N_13684,N_12799,N_12585);
nor U13685 (N_13685,N_12074,N_12812);
nor U13686 (N_13686,N_12776,N_12663);
and U13687 (N_13687,N_12719,N_12718);
nor U13688 (N_13688,N_12144,N_12817);
nand U13689 (N_13689,N_12605,N_12776);
or U13690 (N_13690,N_12716,N_12244);
or U13691 (N_13691,N_12412,N_12767);
nor U13692 (N_13692,N_12667,N_12705);
nand U13693 (N_13693,N_12576,N_12166);
or U13694 (N_13694,N_12869,N_12552);
xnor U13695 (N_13695,N_12234,N_12413);
xor U13696 (N_13696,N_12846,N_12937);
nand U13697 (N_13697,N_12147,N_12964);
nand U13698 (N_13698,N_12264,N_12476);
xor U13699 (N_13699,N_12566,N_12934);
xnor U13700 (N_13700,N_12943,N_12918);
xor U13701 (N_13701,N_12332,N_12153);
or U13702 (N_13702,N_12406,N_12719);
and U13703 (N_13703,N_12697,N_12467);
nor U13704 (N_13704,N_12964,N_12620);
xnor U13705 (N_13705,N_12125,N_12703);
nor U13706 (N_13706,N_12237,N_12483);
or U13707 (N_13707,N_12278,N_12283);
xnor U13708 (N_13708,N_12566,N_12906);
nand U13709 (N_13709,N_12843,N_12819);
nand U13710 (N_13710,N_12917,N_12148);
or U13711 (N_13711,N_12857,N_12267);
xnor U13712 (N_13712,N_12431,N_12633);
nor U13713 (N_13713,N_12948,N_12740);
and U13714 (N_13714,N_12065,N_12052);
xor U13715 (N_13715,N_12469,N_12016);
and U13716 (N_13716,N_12250,N_12391);
and U13717 (N_13717,N_12860,N_12420);
nand U13718 (N_13718,N_12089,N_12350);
nand U13719 (N_13719,N_12225,N_12901);
nand U13720 (N_13720,N_12481,N_12485);
xor U13721 (N_13721,N_12325,N_12112);
xnor U13722 (N_13722,N_12678,N_12217);
and U13723 (N_13723,N_12257,N_12463);
nor U13724 (N_13724,N_12596,N_12316);
nor U13725 (N_13725,N_12504,N_12739);
xor U13726 (N_13726,N_12252,N_12625);
nand U13727 (N_13727,N_12414,N_12100);
or U13728 (N_13728,N_12328,N_12319);
nor U13729 (N_13729,N_12871,N_12199);
nand U13730 (N_13730,N_12826,N_12650);
and U13731 (N_13731,N_12784,N_12487);
or U13732 (N_13732,N_12166,N_12733);
nor U13733 (N_13733,N_12298,N_12977);
nand U13734 (N_13734,N_12438,N_12102);
and U13735 (N_13735,N_12526,N_12732);
and U13736 (N_13736,N_12161,N_12707);
and U13737 (N_13737,N_12450,N_12267);
xor U13738 (N_13738,N_12006,N_12528);
xnor U13739 (N_13739,N_12961,N_12347);
xor U13740 (N_13740,N_12456,N_12299);
xor U13741 (N_13741,N_12866,N_12737);
or U13742 (N_13742,N_12325,N_12688);
or U13743 (N_13743,N_12057,N_12763);
and U13744 (N_13744,N_12235,N_12289);
nor U13745 (N_13745,N_12223,N_12831);
and U13746 (N_13746,N_12052,N_12394);
or U13747 (N_13747,N_12869,N_12738);
nor U13748 (N_13748,N_12525,N_12076);
and U13749 (N_13749,N_12053,N_12396);
and U13750 (N_13750,N_12880,N_12556);
and U13751 (N_13751,N_12046,N_12044);
or U13752 (N_13752,N_12663,N_12356);
nand U13753 (N_13753,N_12186,N_12750);
nand U13754 (N_13754,N_12274,N_12521);
or U13755 (N_13755,N_12795,N_12582);
xnor U13756 (N_13756,N_12675,N_12237);
and U13757 (N_13757,N_12991,N_12597);
nand U13758 (N_13758,N_12983,N_12203);
xnor U13759 (N_13759,N_12430,N_12777);
nor U13760 (N_13760,N_12579,N_12508);
xor U13761 (N_13761,N_12238,N_12090);
xor U13762 (N_13762,N_12744,N_12456);
or U13763 (N_13763,N_12437,N_12899);
nor U13764 (N_13764,N_12795,N_12849);
nor U13765 (N_13765,N_12071,N_12692);
and U13766 (N_13766,N_12572,N_12958);
nor U13767 (N_13767,N_12382,N_12477);
and U13768 (N_13768,N_12785,N_12257);
nor U13769 (N_13769,N_12430,N_12980);
xor U13770 (N_13770,N_12205,N_12358);
or U13771 (N_13771,N_12435,N_12404);
and U13772 (N_13772,N_12921,N_12243);
and U13773 (N_13773,N_12376,N_12018);
and U13774 (N_13774,N_12678,N_12219);
nand U13775 (N_13775,N_12037,N_12922);
and U13776 (N_13776,N_12670,N_12705);
nor U13777 (N_13777,N_12831,N_12474);
nand U13778 (N_13778,N_12316,N_12870);
nor U13779 (N_13779,N_12542,N_12147);
nand U13780 (N_13780,N_12572,N_12176);
xor U13781 (N_13781,N_12429,N_12032);
xor U13782 (N_13782,N_12763,N_12357);
or U13783 (N_13783,N_12080,N_12645);
xor U13784 (N_13784,N_12901,N_12928);
nand U13785 (N_13785,N_12994,N_12242);
nand U13786 (N_13786,N_12436,N_12401);
xnor U13787 (N_13787,N_12068,N_12296);
nor U13788 (N_13788,N_12976,N_12616);
and U13789 (N_13789,N_12805,N_12741);
nand U13790 (N_13790,N_12457,N_12581);
or U13791 (N_13791,N_12806,N_12508);
and U13792 (N_13792,N_12422,N_12161);
nand U13793 (N_13793,N_12588,N_12190);
nand U13794 (N_13794,N_12671,N_12618);
nor U13795 (N_13795,N_12223,N_12113);
and U13796 (N_13796,N_12835,N_12503);
nand U13797 (N_13797,N_12125,N_12654);
nand U13798 (N_13798,N_12914,N_12552);
nor U13799 (N_13799,N_12604,N_12722);
or U13800 (N_13800,N_12569,N_12269);
xnor U13801 (N_13801,N_12376,N_12060);
nor U13802 (N_13802,N_12712,N_12663);
or U13803 (N_13803,N_12679,N_12188);
nor U13804 (N_13804,N_12139,N_12753);
xnor U13805 (N_13805,N_12859,N_12710);
and U13806 (N_13806,N_12848,N_12007);
nor U13807 (N_13807,N_12972,N_12524);
nor U13808 (N_13808,N_12647,N_12480);
and U13809 (N_13809,N_12477,N_12290);
nor U13810 (N_13810,N_12595,N_12635);
and U13811 (N_13811,N_12745,N_12844);
xnor U13812 (N_13812,N_12689,N_12589);
nand U13813 (N_13813,N_12010,N_12561);
or U13814 (N_13814,N_12264,N_12170);
xor U13815 (N_13815,N_12533,N_12099);
nand U13816 (N_13816,N_12942,N_12645);
nor U13817 (N_13817,N_12802,N_12379);
or U13818 (N_13818,N_12285,N_12059);
nand U13819 (N_13819,N_12004,N_12833);
or U13820 (N_13820,N_12578,N_12765);
and U13821 (N_13821,N_12708,N_12656);
nand U13822 (N_13822,N_12119,N_12750);
nand U13823 (N_13823,N_12511,N_12389);
nor U13824 (N_13824,N_12875,N_12929);
xor U13825 (N_13825,N_12420,N_12948);
nand U13826 (N_13826,N_12270,N_12641);
xor U13827 (N_13827,N_12417,N_12022);
and U13828 (N_13828,N_12755,N_12974);
nor U13829 (N_13829,N_12048,N_12022);
xor U13830 (N_13830,N_12702,N_12352);
and U13831 (N_13831,N_12187,N_12675);
nand U13832 (N_13832,N_12623,N_12000);
xor U13833 (N_13833,N_12252,N_12274);
and U13834 (N_13834,N_12578,N_12274);
xor U13835 (N_13835,N_12649,N_12296);
or U13836 (N_13836,N_12191,N_12021);
and U13837 (N_13837,N_12202,N_12629);
xnor U13838 (N_13838,N_12066,N_12851);
xnor U13839 (N_13839,N_12373,N_12623);
and U13840 (N_13840,N_12519,N_12940);
and U13841 (N_13841,N_12220,N_12351);
xor U13842 (N_13842,N_12892,N_12328);
nor U13843 (N_13843,N_12403,N_12659);
nand U13844 (N_13844,N_12415,N_12191);
nor U13845 (N_13845,N_12404,N_12310);
or U13846 (N_13846,N_12177,N_12547);
xor U13847 (N_13847,N_12749,N_12131);
nand U13848 (N_13848,N_12694,N_12106);
nand U13849 (N_13849,N_12385,N_12681);
xnor U13850 (N_13850,N_12429,N_12300);
nor U13851 (N_13851,N_12030,N_12811);
nor U13852 (N_13852,N_12589,N_12819);
nor U13853 (N_13853,N_12211,N_12565);
and U13854 (N_13854,N_12406,N_12518);
and U13855 (N_13855,N_12123,N_12483);
or U13856 (N_13856,N_12140,N_12478);
and U13857 (N_13857,N_12905,N_12294);
xnor U13858 (N_13858,N_12304,N_12993);
and U13859 (N_13859,N_12925,N_12570);
and U13860 (N_13860,N_12069,N_12001);
xnor U13861 (N_13861,N_12308,N_12356);
or U13862 (N_13862,N_12673,N_12186);
or U13863 (N_13863,N_12382,N_12554);
and U13864 (N_13864,N_12303,N_12555);
or U13865 (N_13865,N_12313,N_12210);
xor U13866 (N_13866,N_12439,N_12408);
nor U13867 (N_13867,N_12319,N_12169);
nand U13868 (N_13868,N_12977,N_12516);
or U13869 (N_13869,N_12704,N_12751);
or U13870 (N_13870,N_12424,N_12728);
nand U13871 (N_13871,N_12814,N_12390);
and U13872 (N_13872,N_12580,N_12260);
and U13873 (N_13873,N_12036,N_12498);
nand U13874 (N_13874,N_12131,N_12839);
nor U13875 (N_13875,N_12195,N_12129);
nor U13876 (N_13876,N_12984,N_12801);
and U13877 (N_13877,N_12231,N_12590);
or U13878 (N_13878,N_12276,N_12610);
and U13879 (N_13879,N_12832,N_12496);
nand U13880 (N_13880,N_12344,N_12939);
or U13881 (N_13881,N_12394,N_12423);
nand U13882 (N_13882,N_12317,N_12687);
and U13883 (N_13883,N_12570,N_12069);
or U13884 (N_13884,N_12675,N_12167);
xor U13885 (N_13885,N_12046,N_12374);
and U13886 (N_13886,N_12383,N_12878);
nor U13887 (N_13887,N_12210,N_12863);
nand U13888 (N_13888,N_12254,N_12116);
nor U13889 (N_13889,N_12973,N_12809);
xnor U13890 (N_13890,N_12803,N_12817);
or U13891 (N_13891,N_12349,N_12314);
nand U13892 (N_13892,N_12565,N_12542);
nand U13893 (N_13893,N_12420,N_12209);
nor U13894 (N_13894,N_12035,N_12941);
nand U13895 (N_13895,N_12506,N_12364);
nand U13896 (N_13896,N_12342,N_12720);
xor U13897 (N_13897,N_12606,N_12744);
xor U13898 (N_13898,N_12340,N_12934);
or U13899 (N_13899,N_12081,N_12598);
or U13900 (N_13900,N_12580,N_12630);
or U13901 (N_13901,N_12351,N_12750);
xor U13902 (N_13902,N_12171,N_12446);
or U13903 (N_13903,N_12819,N_12782);
nand U13904 (N_13904,N_12503,N_12861);
and U13905 (N_13905,N_12913,N_12521);
and U13906 (N_13906,N_12393,N_12053);
nor U13907 (N_13907,N_12424,N_12422);
and U13908 (N_13908,N_12865,N_12799);
or U13909 (N_13909,N_12463,N_12950);
or U13910 (N_13910,N_12506,N_12814);
and U13911 (N_13911,N_12790,N_12827);
xor U13912 (N_13912,N_12955,N_12836);
nand U13913 (N_13913,N_12570,N_12440);
or U13914 (N_13914,N_12613,N_12208);
nor U13915 (N_13915,N_12997,N_12374);
nand U13916 (N_13916,N_12030,N_12601);
xnor U13917 (N_13917,N_12831,N_12000);
xor U13918 (N_13918,N_12387,N_12065);
and U13919 (N_13919,N_12796,N_12505);
and U13920 (N_13920,N_12503,N_12923);
or U13921 (N_13921,N_12943,N_12356);
or U13922 (N_13922,N_12753,N_12177);
nor U13923 (N_13923,N_12907,N_12040);
nand U13924 (N_13924,N_12429,N_12096);
nor U13925 (N_13925,N_12739,N_12821);
or U13926 (N_13926,N_12921,N_12573);
xor U13927 (N_13927,N_12572,N_12883);
nand U13928 (N_13928,N_12376,N_12714);
nor U13929 (N_13929,N_12084,N_12908);
or U13930 (N_13930,N_12641,N_12803);
nand U13931 (N_13931,N_12222,N_12080);
or U13932 (N_13932,N_12349,N_12494);
or U13933 (N_13933,N_12815,N_12529);
xor U13934 (N_13934,N_12124,N_12347);
nand U13935 (N_13935,N_12540,N_12901);
or U13936 (N_13936,N_12814,N_12394);
or U13937 (N_13937,N_12418,N_12222);
xnor U13938 (N_13938,N_12511,N_12788);
nand U13939 (N_13939,N_12771,N_12022);
nand U13940 (N_13940,N_12224,N_12727);
xnor U13941 (N_13941,N_12831,N_12884);
and U13942 (N_13942,N_12818,N_12865);
and U13943 (N_13943,N_12778,N_12592);
nor U13944 (N_13944,N_12263,N_12850);
or U13945 (N_13945,N_12072,N_12789);
xnor U13946 (N_13946,N_12015,N_12684);
and U13947 (N_13947,N_12103,N_12921);
and U13948 (N_13948,N_12073,N_12851);
nand U13949 (N_13949,N_12807,N_12073);
or U13950 (N_13950,N_12119,N_12317);
and U13951 (N_13951,N_12185,N_12321);
nor U13952 (N_13952,N_12406,N_12443);
or U13953 (N_13953,N_12713,N_12696);
nor U13954 (N_13954,N_12733,N_12441);
or U13955 (N_13955,N_12723,N_12838);
nand U13956 (N_13956,N_12254,N_12676);
nand U13957 (N_13957,N_12976,N_12388);
nor U13958 (N_13958,N_12778,N_12521);
and U13959 (N_13959,N_12005,N_12374);
or U13960 (N_13960,N_12869,N_12850);
or U13961 (N_13961,N_12709,N_12388);
nor U13962 (N_13962,N_12163,N_12747);
nand U13963 (N_13963,N_12797,N_12882);
or U13964 (N_13964,N_12203,N_12018);
nand U13965 (N_13965,N_12330,N_12326);
xor U13966 (N_13966,N_12161,N_12429);
and U13967 (N_13967,N_12906,N_12523);
and U13968 (N_13968,N_12817,N_12451);
or U13969 (N_13969,N_12485,N_12176);
xnor U13970 (N_13970,N_12110,N_12220);
or U13971 (N_13971,N_12684,N_12327);
and U13972 (N_13972,N_12515,N_12970);
or U13973 (N_13973,N_12990,N_12178);
or U13974 (N_13974,N_12286,N_12061);
nand U13975 (N_13975,N_12141,N_12774);
xnor U13976 (N_13976,N_12387,N_12760);
nand U13977 (N_13977,N_12823,N_12428);
and U13978 (N_13978,N_12547,N_12947);
xor U13979 (N_13979,N_12027,N_12701);
nor U13980 (N_13980,N_12829,N_12453);
nand U13981 (N_13981,N_12624,N_12605);
xor U13982 (N_13982,N_12737,N_12056);
nor U13983 (N_13983,N_12373,N_12409);
or U13984 (N_13984,N_12172,N_12616);
and U13985 (N_13985,N_12917,N_12132);
or U13986 (N_13986,N_12263,N_12401);
xnor U13987 (N_13987,N_12810,N_12965);
or U13988 (N_13988,N_12300,N_12449);
and U13989 (N_13989,N_12007,N_12519);
xor U13990 (N_13990,N_12822,N_12260);
xor U13991 (N_13991,N_12712,N_12784);
nor U13992 (N_13992,N_12309,N_12633);
nand U13993 (N_13993,N_12817,N_12853);
or U13994 (N_13994,N_12815,N_12492);
and U13995 (N_13995,N_12463,N_12503);
nor U13996 (N_13996,N_12075,N_12254);
nor U13997 (N_13997,N_12216,N_12008);
and U13998 (N_13998,N_12844,N_12037);
nor U13999 (N_13999,N_12639,N_12582);
and U14000 (N_14000,N_13041,N_13177);
nor U14001 (N_14001,N_13319,N_13506);
nand U14002 (N_14002,N_13308,N_13811);
nor U14003 (N_14003,N_13638,N_13067);
nand U14004 (N_14004,N_13714,N_13281);
xnor U14005 (N_14005,N_13813,N_13136);
nor U14006 (N_14006,N_13210,N_13610);
or U14007 (N_14007,N_13917,N_13590);
or U14008 (N_14008,N_13592,N_13483);
and U14009 (N_14009,N_13407,N_13330);
nand U14010 (N_14010,N_13167,N_13804);
nand U14011 (N_14011,N_13348,N_13669);
xnor U14012 (N_14012,N_13595,N_13773);
nor U14013 (N_14013,N_13869,N_13430);
or U14014 (N_14014,N_13109,N_13049);
xor U14015 (N_14015,N_13116,N_13553);
or U14016 (N_14016,N_13973,N_13013);
xnor U14017 (N_14017,N_13472,N_13708);
and U14018 (N_14018,N_13182,N_13137);
or U14019 (N_14019,N_13089,N_13462);
nor U14020 (N_14020,N_13583,N_13215);
and U14021 (N_14021,N_13873,N_13941);
or U14022 (N_14022,N_13364,N_13436);
nor U14023 (N_14023,N_13535,N_13115);
nor U14024 (N_14024,N_13517,N_13062);
or U14025 (N_14025,N_13198,N_13290);
nor U14026 (N_14026,N_13050,N_13056);
nor U14027 (N_14027,N_13826,N_13850);
or U14028 (N_14028,N_13753,N_13931);
nor U14029 (N_14029,N_13480,N_13523);
nor U14030 (N_14030,N_13699,N_13284);
or U14031 (N_14031,N_13191,N_13539);
or U14032 (N_14032,N_13456,N_13183);
xor U14033 (N_14033,N_13259,N_13149);
xnor U14034 (N_14034,N_13018,N_13060);
xnor U14035 (N_14035,N_13943,N_13048);
and U14036 (N_14036,N_13511,N_13924);
xor U14037 (N_14037,N_13887,N_13971);
or U14038 (N_14038,N_13596,N_13494);
nor U14039 (N_14039,N_13176,N_13522);
nand U14040 (N_14040,N_13527,N_13818);
nand U14041 (N_14041,N_13328,N_13897);
xor U14042 (N_14042,N_13286,N_13620);
and U14043 (N_14043,N_13237,N_13750);
and U14044 (N_14044,N_13489,N_13168);
xor U14045 (N_14045,N_13147,N_13028);
nand U14046 (N_14046,N_13443,N_13758);
and U14047 (N_14047,N_13691,N_13948);
xnor U14048 (N_14048,N_13900,N_13022);
xor U14049 (N_14049,N_13081,N_13894);
nand U14050 (N_14050,N_13731,N_13232);
or U14051 (N_14051,N_13180,N_13497);
or U14052 (N_14052,N_13179,N_13432);
and U14053 (N_14053,N_13678,N_13602);
xor U14054 (N_14054,N_13275,N_13188);
or U14055 (N_14055,N_13248,N_13085);
or U14056 (N_14056,N_13297,N_13304);
and U14057 (N_14057,N_13142,N_13547);
nand U14058 (N_14058,N_13730,N_13800);
xnor U14059 (N_14059,N_13847,N_13615);
nor U14060 (N_14060,N_13040,N_13208);
or U14061 (N_14061,N_13078,N_13203);
nand U14062 (N_14062,N_13352,N_13556);
nand U14063 (N_14063,N_13760,N_13575);
nand U14064 (N_14064,N_13710,N_13171);
or U14065 (N_14065,N_13947,N_13907);
xor U14066 (N_14066,N_13829,N_13353);
xor U14067 (N_14067,N_13026,N_13487);
or U14068 (N_14068,N_13564,N_13193);
or U14069 (N_14069,N_13054,N_13955);
or U14070 (N_14070,N_13791,N_13832);
nor U14071 (N_14071,N_13543,N_13295);
and U14072 (N_14072,N_13382,N_13502);
xnor U14073 (N_14073,N_13055,N_13102);
xor U14074 (N_14074,N_13902,N_13032);
nor U14075 (N_14075,N_13733,N_13439);
nand U14076 (N_14076,N_13127,N_13743);
or U14077 (N_14077,N_13244,N_13589);
or U14078 (N_14078,N_13676,N_13314);
xor U14079 (N_14079,N_13420,N_13510);
xnor U14080 (N_14080,N_13234,N_13036);
nor U14081 (N_14081,N_13076,N_13698);
nand U14082 (N_14082,N_13812,N_13482);
or U14083 (N_14083,N_13819,N_13378);
nor U14084 (N_14084,N_13607,N_13920);
xor U14085 (N_14085,N_13192,N_13618);
nor U14086 (N_14086,N_13571,N_13519);
and U14087 (N_14087,N_13991,N_13937);
xnor U14088 (N_14088,N_13389,N_13910);
xnor U14089 (N_14089,N_13379,N_13993);
nand U14090 (N_14090,N_13435,N_13512);
nor U14091 (N_14091,N_13383,N_13119);
nor U14092 (N_14092,N_13122,N_13186);
or U14093 (N_14093,N_13662,N_13656);
and U14094 (N_14094,N_13222,N_13940);
or U14095 (N_14095,N_13767,N_13741);
and U14096 (N_14096,N_13452,N_13331);
xnor U14097 (N_14097,N_13141,N_13311);
xnor U14098 (N_14098,N_13132,N_13987);
nand U14099 (N_14099,N_13031,N_13852);
or U14100 (N_14100,N_13928,N_13488);
nor U14101 (N_14101,N_13732,N_13632);
nand U14102 (N_14102,N_13005,N_13358);
nor U14103 (N_14103,N_13516,N_13751);
or U14104 (N_14104,N_13762,N_13793);
nor U14105 (N_14105,N_13004,N_13694);
and U14106 (N_14106,N_13112,N_13289);
nor U14107 (N_14107,N_13303,N_13672);
nor U14108 (N_14108,N_13396,N_13916);
and U14109 (N_14109,N_13969,N_13939);
or U14110 (N_14110,N_13737,N_13010);
nor U14111 (N_14111,N_13460,N_13992);
or U14112 (N_14112,N_13027,N_13270);
nor U14113 (N_14113,N_13346,N_13824);
nand U14114 (N_14114,N_13957,N_13219);
nand U14115 (N_14115,N_13283,N_13810);
or U14116 (N_14116,N_13989,N_13377);
xnor U14117 (N_14117,N_13318,N_13356);
or U14118 (N_14118,N_13084,N_13809);
xnor U14119 (N_14119,N_13034,N_13463);
xnor U14120 (N_14120,N_13256,N_13059);
xnor U14121 (N_14121,N_13133,N_13785);
or U14122 (N_14122,N_13474,N_13313);
nand U14123 (N_14123,N_13808,N_13475);
and U14124 (N_14124,N_13601,N_13674);
xor U14125 (N_14125,N_13301,N_13425);
and U14126 (N_14126,N_13650,N_13250);
nor U14127 (N_14127,N_13169,N_13798);
and U14128 (N_14128,N_13229,N_13901);
nand U14129 (N_14129,N_13172,N_13552);
xor U14130 (N_14130,N_13603,N_13082);
and U14131 (N_14131,N_13926,N_13268);
nor U14132 (N_14132,N_13934,N_13675);
or U14133 (N_14133,N_13775,N_13706);
nand U14134 (N_14134,N_13230,N_13306);
nand U14135 (N_14135,N_13503,N_13406);
nor U14136 (N_14136,N_13424,N_13994);
nor U14137 (N_14137,N_13000,N_13677);
nor U14138 (N_14138,N_13189,N_13044);
xor U14139 (N_14139,N_13039,N_13799);
nor U14140 (N_14140,N_13144,N_13337);
nor U14141 (N_14141,N_13562,N_13763);
nor U14142 (N_14142,N_13140,N_13114);
nand U14143 (N_14143,N_13185,N_13093);
and U14144 (N_14144,N_13954,N_13980);
xor U14145 (N_14145,N_13685,N_13163);
and U14146 (N_14146,N_13849,N_13944);
xor U14147 (N_14147,N_13438,N_13164);
nor U14148 (N_14148,N_13431,N_13293);
xor U14149 (N_14149,N_13912,N_13448);
nand U14150 (N_14150,N_13083,N_13146);
or U14151 (N_14151,N_13045,N_13716);
nand U14152 (N_14152,N_13573,N_13752);
nand U14153 (N_14153,N_13009,N_13249);
xor U14154 (N_14154,N_13789,N_13046);
xnor U14155 (N_14155,N_13243,N_13047);
xor U14156 (N_14156,N_13123,N_13367);
nand U14157 (N_14157,N_13768,N_13405);
and U14158 (N_14158,N_13484,N_13029);
xnor U14159 (N_14159,N_13101,N_13659);
and U14160 (N_14160,N_13679,N_13441);
xnor U14161 (N_14161,N_13058,N_13651);
nor U14162 (N_14162,N_13722,N_13375);
nand U14163 (N_14163,N_13366,N_13950);
nand U14164 (N_14164,N_13534,N_13844);
nor U14165 (N_14165,N_13953,N_13196);
nand U14166 (N_14166,N_13876,N_13225);
nand U14167 (N_14167,N_13823,N_13922);
xnor U14168 (N_14168,N_13066,N_13423);
or U14169 (N_14169,N_13074,N_13889);
or U14170 (N_14170,N_13972,N_13559);
nand U14171 (N_14171,N_13279,N_13199);
nor U14172 (N_14172,N_13715,N_13326);
and U14173 (N_14173,N_13492,N_13509);
xnor U14174 (N_14174,N_13445,N_13086);
nand U14175 (N_14175,N_13979,N_13365);
nor U14176 (N_14176,N_13689,N_13749);
nand U14177 (N_14177,N_13363,N_13576);
or U14178 (N_14178,N_13621,N_13064);
nor U14179 (N_14179,N_13288,N_13828);
nor U14180 (N_14180,N_13848,N_13568);
xnor U14181 (N_14181,N_13412,N_13857);
xnor U14182 (N_14182,N_13440,N_13106);
nor U14183 (N_14183,N_13877,N_13051);
nand U14184 (N_14184,N_13187,N_13946);
and U14185 (N_14185,N_13012,N_13280);
or U14186 (N_14186,N_13345,N_13017);
xor U14187 (N_14187,N_13342,N_13411);
and U14188 (N_14188,N_13645,N_13956);
or U14189 (N_14189,N_13967,N_13960);
or U14190 (N_14190,N_13644,N_13218);
nor U14191 (N_14191,N_13663,N_13421);
nor U14192 (N_14192,N_13719,N_13360);
nand U14193 (N_14193,N_13403,N_13988);
xnor U14194 (N_14194,N_13121,N_13817);
xnor U14195 (N_14195,N_13129,N_13336);
xor U14196 (N_14196,N_13742,N_13666);
nand U14197 (N_14197,N_13764,N_13837);
xor U14198 (N_14198,N_13409,N_13518);
nand U14199 (N_14199,N_13200,N_13267);
nand U14200 (N_14200,N_13376,N_13317);
xor U14201 (N_14201,N_13524,N_13744);
or U14202 (N_14202,N_13619,N_13238);
nor U14203 (N_14203,N_13725,N_13052);
nor U14204 (N_14204,N_13467,N_13766);
or U14205 (N_14205,N_13696,N_13305);
xor U14206 (N_14206,N_13624,N_13613);
and U14207 (N_14207,N_13778,N_13830);
or U14208 (N_14208,N_13614,N_13588);
xor U14209 (N_14209,N_13385,N_13854);
and U14210 (N_14210,N_13531,N_13608);
xor U14211 (N_14211,N_13549,N_13653);
and U14212 (N_14212,N_13871,N_13158);
nor U14213 (N_14213,N_13961,N_13966);
nand U14214 (N_14214,N_13867,N_13661);
xor U14215 (N_14215,N_13491,N_13151);
nand U14216 (N_14216,N_13388,N_13555);
and U14217 (N_14217,N_13104,N_13473);
nor U14218 (N_14218,N_13888,N_13839);
xnor U14219 (N_14219,N_13560,N_13780);
xor U14220 (N_14220,N_13231,N_13860);
or U14221 (N_14221,N_13011,N_13736);
and U14222 (N_14222,N_13533,N_13938);
and U14223 (N_14223,N_13466,N_13657);
xnor U14224 (N_14224,N_13513,N_13214);
xor U14225 (N_14225,N_13984,N_13194);
nor U14226 (N_14226,N_13242,N_13429);
and U14227 (N_14227,N_13680,N_13983);
or U14228 (N_14228,N_13251,N_13859);
nand U14229 (N_14229,N_13855,N_13341);
nor U14230 (N_14230,N_13415,N_13393);
xor U14231 (N_14231,N_13368,N_13501);
or U14232 (N_14232,N_13628,N_13410);
xor U14233 (N_14233,N_13264,N_13557);
or U14234 (N_14234,N_13670,N_13373);
nand U14235 (N_14235,N_13520,N_13468);
nor U14236 (N_14236,N_13801,N_13426);
nor U14237 (N_14237,N_13577,N_13038);
nand U14238 (N_14238,N_13478,N_13007);
nor U14239 (N_14239,N_13963,N_13063);
xor U14240 (N_14240,N_13880,N_13371);
nor U14241 (N_14241,N_13327,N_13515);
nand U14242 (N_14242,N_13874,N_13913);
or U14243 (N_14243,N_13355,N_13687);
xnor U14244 (N_14244,N_13858,N_13496);
and U14245 (N_14245,N_13145,N_13779);
or U14246 (N_14246,N_13160,N_13395);
nand U14247 (N_14247,N_13374,N_13761);
nor U14248 (N_14248,N_13092,N_13580);
and U14249 (N_14249,N_13197,N_13444);
or U14250 (N_14250,N_13254,N_13921);
xor U14251 (N_14251,N_13500,N_13490);
nor U14252 (N_14252,N_13759,N_13591);
nor U14253 (N_14253,N_13235,N_13241);
xor U14254 (N_14254,N_13636,N_13831);
and U14255 (N_14255,N_13097,N_13099);
nand U14256 (N_14256,N_13587,N_13386);
nor U14257 (N_14257,N_13300,N_13833);
nand U14258 (N_14258,N_13864,N_13959);
nand U14259 (N_14259,N_13999,N_13970);
xnor U14260 (N_14260,N_13566,N_13397);
nand U14261 (N_14261,N_13124,N_13755);
nor U14262 (N_14262,N_13709,N_13205);
or U14263 (N_14263,N_13226,N_13126);
or U14264 (N_14264,N_13545,N_13053);
or U14265 (N_14265,N_13820,N_13540);
and U14266 (N_14266,N_13446,N_13339);
nor U14267 (N_14267,N_13875,N_13143);
nor U14268 (N_14268,N_13274,N_13713);
xor U14269 (N_14269,N_13729,N_13184);
nand U14270 (N_14270,N_13043,N_13227);
xor U14271 (N_14271,N_13673,N_13181);
nor U14272 (N_14272,N_13261,N_13681);
or U14273 (N_14273,N_13903,N_13015);
and U14274 (N_14274,N_13285,N_13890);
and U14275 (N_14275,N_13981,N_13521);
or U14276 (N_14276,N_13025,N_13906);
or U14277 (N_14277,N_13629,N_13175);
or U14278 (N_14278,N_13493,N_13335);
nand U14279 (N_14279,N_13643,N_13447);
xnor U14280 (N_14280,N_13221,N_13206);
nand U14281 (N_14281,N_13927,N_13792);
or U14282 (N_14282,N_13686,N_13077);
or U14283 (N_14283,N_13597,N_13257);
or U14284 (N_14284,N_13929,N_13951);
and U14285 (N_14285,N_13770,N_13451);
xnor U14286 (N_14286,N_13612,N_13434);
nor U14287 (N_14287,N_13351,N_13100);
nor U14288 (N_14288,N_13795,N_13886);
nand U14289 (N_14289,N_13370,N_13006);
xnor U14290 (N_14290,N_13247,N_13418);
or U14291 (N_14291,N_13882,N_13647);
nor U14292 (N_14292,N_13417,N_13098);
or U14293 (N_14293,N_13162,N_13428);
or U14294 (N_14294,N_13135,N_13756);
nor U14295 (N_14295,N_13195,N_13498);
or U14296 (N_14296,N_13905,N_13223);
nand U14297 (N_14297,N_13148,N_13682);
nand U14298 (N_14298,N_13582,N_13641);
or U14299 (N_14299,N_13605,N_13457);
xor U14300 (N_14300,N_13945,N_13623);
or U14301 (N_14301,N_13296,N_13978);
and U14302 (N_14302,N_13975,N_13538);
and U14303 (N_14303,N_13726,N_13783);
xor U14304 (N_14304,N_13541,N_13325);
xnor U14305 (N_14305,N_13505,N_13340);
nor U14306 (N_14306,N_13724,N_13035);
or U14307 (N_14307,N_13625,N_13637);
or U14308 (N_14308,N_13668,N_13787);
or U14309 (N_14309,N_13246,N_13727);
xor U14310 (N_14310,N_13061,N_13861);
nor U14311 (N_14311,N_13703,N_13486);
and U14312 (N_14312,N_13578,N_13454);
nor U14313 (N_14313,N_13458,N_13350);
and U14314 (N_14314,N_13822,N_13019);
nor U14315 (N_14315,N_13631,N_13170);
or U14316 (N_14316,N_13413,N_13260);
nor U14317 (N_14317,N_13125,N_13885);
nand U14318 (N_14318,N_13307,N_13344);
nand U14319 (N_14319,N_13033,N_13479);
and U14320 (N_14320,N_13204,N_13131);
nor U14321 (N_14321,N_13788,N_13211);
xor U14322 (N_14322,N_13648,N_13532);
nor U14323 (N_14323,N_13707,N_13400);
nor U14324 (N_14324,N_13095,N_13606);
xnor U14325 (N_14325,N_13654,N_13797);
and U14326 (N_14326,N_13834,N_13233);
or U14327 (N_14327,N_13658,N_13572);
or U14328 (N_14328,N_13117,N_13477);
and U14329 (N_14329,N_13693,N_13369);
nand U14330 (N_14330,N_13087,N_13359);
or U14331 (N_14331,N_13544,N_13842);
nor U14332 (N_14332,N_13273,N_13481);
nor U14333 (N_14333,N_13914,N_13807);
nor U14334 (N_14334,N_13329,N_13190);
nor U14335 (N_14335,N_13271,N_13723);
xor U14336 (N_14336,N_13622,N_13495);
xor U14337 (N_14337,N_13827,N_13213);
nor U14338 (N_14338,N_13459,N_13918);
nand U14339 (N_14339,N_13150,N_13001);
xnor U14340 (N_14340,N_13630,N_13702);
xor U14341 (N_14341,N_13008,N_13825);
xor U14342 (N_14342,N_13633,N_13245);
xor U14343 (N_14343,N_13646,N_13757);
nor U14344 (N_14344,N_13514,N_13253);
or U14345 (N_14345,N_13090,N_13224);
xnor U14346 (N_14346,N_13700,N_13546);
nor U14347 (N_14347,N_13754,N_13739);
nand U14348 (N_14348,N_13923,N_13806);
nand U14349 (N_14349,N_13649,N_13042);
nand U14350 (N_14350,N_13201,N_13096);
nand U14351 (N_14351,N_13252,N_13909);
nand U14352 (N_14352,N_13952,N_13688);
or U14353 (N_14353,N_13391,N_13016);
nand U14354 (N_14354,N_13617,N_13173);
nor U14355 (N_14355,N_13915,N_13165);
xnor U14356 (N_14356,N_13402,N_13471);
nor U14357 (N_14357,N_13153,N_13394);
nand U14358 (N_14358,N_13962,N_13536);
or U14359 (N_14359,N_13997,N_13239);
and U14360 (N_14360,N_13380,N_13690);
or U14361 (N_14361,N_13684,N_13118);
xor U14362 (N_14362,N_13387,N_13504);
or U14363 (N_14363,N_13639,N_13712);
or U14364 (N_14364,N_13734,N_13816);
and U14365 (N_14365,N_13128,N_13349);
xor U14366 (N_14366,N_13728,N_13266);
or U14367 (N_14367,N_13416,N_13652);
and U14368 (N_14368,N_13020,N_13419);
nand U14369 (N_14369,N_13277,N_13476);
nor U14370 (N_14370,N_13990,N_13265);
xor U14371 (N_14371,N_13720,N_13878);
and U14372 (N_14372,N_13600,N_13316);
or U14373 (N_14373,N_13073,N_13784);
nand U14374 (N_14374,N_13071,N_13558);
and U14375 (N_14375,N_13701,N_13786);
nand U14376 (N_14376,N_13161,N_13695);
or U14377 (N_14377,N_13398,N_13986);
nor U14378 (N_14378,N_13781,N_13642);
nor U14379 (N_14379,N_13110,N_13958);
nor U14380 (N_14380,N_13347,N_13507);
nor U14381 (N_14381,N_13068,N_13870);
nand U14382 (N_14382,N_13977,N_13469);
nor U14383 (N_14383,N_13212,N_13088);
nor U14384 (N_14384,N_13401,N_13292);
xor U14385 (N_14385,N_13548,N_13079);
nor U14386 (N_14386,N_13841,N_13838);
nand U14387 (N_14387,N_13911,N_13014);
and U14388 (N_14388,N_13771,N_13738);
nor U14389 (N_14389,N_13103,N_13333);
and U14390 (N_14390,N_13616,N_13278);
nand U14391 (N_14391,N_13627,N_13711);
nand U14392 (N_14392,N_13671,N_13790);
or U14393 (N_14393,N_13299,N_13872);
nor U14394 (N_14394,N_13803,N_13207);
nand U14395 (N_14395,N_13372,N_13156);
nand U14396 (N_14396,N_13057,N_13263);
or U14397 (N_14397,N_13626,N_13777);
or U14398 (N_14398,N_13065,N_13209);
nand U14399 (N_14399,N_13091,N_13414);
xnor U14400 (N_14400,N_13357,N_13321);
or U14401 (N_14401,N_13765,N_13134);
xor U14402 (N_14402,N_13310,N_13932);
nor U14403 (N_14403,N_13846,N_13107);
and U14404 (N_14404,N_13717,N_13996);
xor U14405 (N_14405,N_13465,N_13868);
nand U14406 (N_14406,N_13598,N_13745);
nand U14407 (N_14407,N_13139,N_13262);
and U14408 (N_14408,N_13105,N_13069);
or U14409 (N_14409,N_13904,N_13399);
or U14410 (N_14410,N_13282,N_13236);
and U14411 (N_14411,N_13152,N_13721);
nand U14412 (N_14412,N_13269,N_13362);
nand U14413 (N_14413,N_13354,N_13692);
nand U14414 (N_14414,N_13735,N_13879);
nor U14415 (N_14415,N_13499,N_13113);
nor U14416 (N_14416,N_13704,N_13567);
xnor U14417 (N_14417,N_13843,N_13856);
and U14418 (N_14418,N_13998,N_13525);
nor U14419 (N_14419,N_13772,N_13974);
or U14420 (N_14420,N_13746,N_13272);
and U14421 (N_14421,N_13166,N_13574);
nand U14422 (N_14422,N_13111,N_13528);
or U14423 (N_14423,N_13949,N_13381);
or U14424 (N_14424,N_13740,N_13258);
and U14425 (N_14425,N_13291,N_13569);
nor U14426 (N_14426,N_13774,N_13794);
xor U14427 (N_14427,N_13485,N_13526);
and U14428 (N_14428,N_13030,N_13453);
nand U14429 (N_14429,N_13866,N_13667);
or U14430 (N_14430,N_13565,N_13542);
nand U14431 (N_14431,N_13120,N_13899);
or U14432 (N_14432,N_13202,N_13935);
nor U14433 (N_14433,N_13220,N_13585);
nand U14434 (N_14434,N_13461,N_13718);
xor U14435 (N_14435,N_13217,N_13862);
nor U14436 (N_14436,N_13508,N_13964);
nor U14437 (N_14437,N_13815,N_13240);
xnor U14438 (N_14438,N_13450,N_13361);
or U14439 (N_14439,N_13130,N_13898);
nor U14440 (N_14440,N_13315,N_13343);
nand U14441 (N_14441,N_13561,N_13072);
and U14442 (N_14442,N_13155,N_13995);
and U14443 (N_14443,N_13570,N_13863);
and U14444 (N_14444,N_13925,N_13108);
nand U14445 (N_14445,N_13427,N_13896);
and U14446 (N_14446,N_13640,N_13579);
and U14447 (N_14447,N_13455,N_13529);
and U14448 (N_14448,N_13604,N_13891);
xor U14449 (N_14449,N_13634,N_13985);
and U14450 (N_14450,N_13174,N_13982);
nand U14451 (N_14451,N_13594,N_13021);
xor U14452 (N_14452,N_13023,N_13747);
nand U14453 (N_14453,N_13611,N_13748);
and U14454 (N_14454,N_13323,N_13930);
and U14455 (N_14455,N_13390,N_13593);
nor U14456 (N_14456,N_13835,N_13881);
xnor U14457 (N_14457,N_13554,N_13437);
or U14458 (N_14458,N_13584,N_13530);
nand U14459 (N_14459,N_13893,N_13216);
nand U14460 (N_14460,N_13563,N_13802);
and U14461 (N_14461,N_13840,N_13895);
nor U14462 (N_14462,N_13294,N_13853);
or U14463 (N_14463,N_13965,N_13635);
and U14464 (N_14464,N_13159,N_13255);
or U14465 (N_14465,N_13884,N_13933);
xor U14466 (N_14466,N_13942,N_13024);
xor U14467 (N_14467,N_13865,N_13609);
xnor U14468 (N_14468,N_13094,N_13883);
or U14469 (N_14469,N_13287,N_13776);
xnor U14470 (N_14470,N_13154,N_13919);
xor U14471 (N_14471,N_13298,N_13080);
xor U14472 (N_14472,N_13908,N_13782);
or U14473 (N_14473,N_13228,N_13334);
or U14474 (N_14474,N_13178,N_13892);
and U14475 (N_14475,N_13586,N_13551);
and U14476 (N_14476,N_13550,N_13422);
nand U14477 (N_14477,N_13037,N_13660);
xor U14478 (N_14478,N_13324,N_13449);
or U14479 (N_14479,N_13599,N_13442);
nand U14480 (N_14480,N_13138,N_13075);
nor U14481 (N_14481,N_13070,N_13976);
and U14482 (N_14482,N_13683,N_13309);
or U14483 (N_14483,N_13302,N_13157);
or U14484 (N_14484,N_13003,N_13312);
xnor U14485 (N_14485,N_13769,N_13664);
and U14486 (N_14486,N_13665,N_13384);
xnor U14487 (N_14487,N_13002,N_13845);
nand U14488 (N_14488,N_13338,N_13276);
or U14489 (N_14489,N_13470,N_13836);
or U14490 (N_14490,N_13705,N_13464);
xor U14491 (N_14491,N_13322,N_13655);
nand U14492 (N_14492,N_13697,N_13332);
nand U14493 (N_14493,N_13537,N_13404);
nand U14494 (N_14494,N_13392,N_13320);
or U14495 (N_14495,N_13851,N_13408);
or U14496 (N_14496,N_13814,N_13581);
nand U14497 (N_14497,N_13805,N_13968);
nand U14498 (N_14498,N_13936,N_13433);
and U14499 (N_14499,N_13821,N_13796);
xor U14500 (N_14500,N_13966,N_13205);
and U14501 (N_14501,N_13254,N_13771);
and U14502 (N_14502,N_13545,N_13662);
or U14503 (N_14503,N_13584,N_13377);
and U14504 (N_14504,N_13244,N_13058);
and U14505 (N_14505,N_13635,N_13146);
or U14506 (N_14506,N_13435,N_13826);
xnor U14507 (N_14507,N_13987,N_13064);
or U14508 (N_14508,N_13955,N_13776);
xor U14509 (N_14509,N_13584,N_13547);
and U14510 (N_14510,N_13931,N_13631);
and U14511 (N_14511,N_13540,N_13667);
xnor U14512 (N_14512,N_13143,N_13630);
and U14513 (N_14513,N_13454,N_13815);
nor U14514 (N_14514,N_13098,N_13995);
and U14515 (N_14515,N_13532,N_13402);
nor U14516 (N_14516,N_13362,N_13772);
xor U14517 (N_14517,N_13019,N_13525);
nand U14518 (N_14518,N_13629,N_13910);
nor U14519 (N_14519,N_13726,N_13250);
nand U14520 (N_14520,N_13654,N_13249);
nor U14521 (N_14521,N_13978,N_13680);
or U14522 (N_14522,N_13618,N_13907);
nand U14523 (N_14523,N_13756,N_13719);
xor U14524 (N_14524,N_13427,N_13536);
nand U14525 (N_14525,N_13560,N_13155);
and U14526 (N_14526,N_13000,N_13870);
and U14527 (N_14527,N_13002,N_13394);
or U14528 (N_14528,N_13063,N_13267);
nor U14529 (N_14529,N_13350,N_13713);
or U14530 (N_14530,N_13968,N_13880);
and U14531 (N_14531,N_13250,N_13617);
nand U14532 (N_14532,N_13633,N_13771);
nor U14533 (N_14533,N_13523,N_13871);
xnor U14534 (N_14534,N_13931,N_13114);
and U14535 (N_14535,N_13402,N_13397);
nand U14536 (N_14536,N_13429,N_13202);
or U14537 (N_14537,N_13237,N_13510);
and U14538 (N_14538,N_13141,N_13127);
or U14539 (N_14539,N_13001,N_13357);
and U14540 (N_14540,N_13583,N_13795);
nand U14541 (N_14541,N_13797,N_13454);
or U14542 (N_14542,N_13842,N_13798);
nand U14543 (N_14543,N_13815,N_13047);
xor U14544 (N_14544,N_13095,N_13919);
or U14545 (N_14545,N_13385,N_13574);
xor U14546 (N_14546,N_13132,N_13793);
xor U14547 (N_14547,N_13664,N_13038);
xnor U14548 (N_14548,N_13223,N_13919);
xnor U14549 (N_14549,N_13471,N_13074);
nand U14550 (N_14550,N_13307,N_13122);
and U14551 (N_14551,N_13928,N_13599);
nor U14552 (N_14552,N_13740,N_13834);
nor U14553 (N_14553,N_13033,N_13247);
xor U14554 (N_14554,N_13555,N_13561);
xor U14555 (N_14555,N_13379,N_13319);
xor U14556 (N_14556,N_13502,N_13094);
and U14557 (N_14557,N_13233,N_13274);
and U14558 (N_14558,N_13283,N_13063);
and U14559 (N_14559,N_13945,N_13745);
or U14560 (N_14560,N_13678,N_13322);
or U14561 (N_14561,N_13878,N_13215);
or U14562 (N_14562,N_13927,N_13791);
or U14563 (N_14563,N_13258,N_13945);
xor U14564 (N_14564,N_13435,N_13859);
xnor U14565 (N_14565,N_13829,N_13039);
and U14566 (N_14566,N_13551,N_13027);
and U14567 (N_14567,N_13368,N_13607);
nor U14568 (N_14568,N_13929,N_13642);
nand U14569 (N_14569,N_13458,N_13479);
or U14570 (N_14570,N_13368,N_13126);
and U14571 (N_14571,N_13507,N_13431);
nor U14572 (N_14572,N_13111,N_13582);
nor U14573 (N_14573,N_13239,N_13291);
nand U14574 (N_14574,N_13100,N_13466);
xnor U14575 (N_14575,N_13280,N_13078);
nand U14576 (N_14576,N_13209,N_13140);
xor U14577 (N_14577,N_13701,N_13780);
or U14578 (N_14578,N_13898,N_13843);
xor U14579 (N_14579,N_13465,N_13625);
and U14580 (N_14580,N_13988,N_13674);
or U14581 (N_14581,N_13230,N_13585);
xor U14582 (N_14582,N_13444,N_13277);
nand U14583 (N_14583,N_13525,N_13443);
nor U14584 (N_14584,N_13284,N_13358);
or U14585 (N_14585,N_13304,N_13366);
xor U14586 (N_14586,N_13390,N_13023);
nand U14587 (N_14587,N_13729,N_13598);
nor U14588 (N_14588,N_13171,N_13249);
or U14589 (N_14589,N_13804,N_13335);
nor U14590 (N_14590,N_13693,N_13925);
xor U14591 (N_14591,N_13080,N_13032);
nand U14592 (N_14592,N_13090,N_13830);
xnor U14593 (N_14593,N_13221,N_13153);
nor U14594 (N_14594,N_13465,N_13038);
xnor U14595 (N_14595,N_13452,N_13937);
xnor U14596 (N_14596,N_13768,N_13666);
or U14597 (N_14597,N_13741,N_13543);
and U14598 (N_14598,N_13326,N_13859);
nand U14599 (N_14599,N_13434,N_13829);
and U14600 (N_14600,N_13781,N_13687);
xnor U14601 (N_14601,N_13939,N_13944);
and U14602 (N_14602,N_13201,N_13617);
xor U14603 (N_14603,N_13469,N_13697);
xor U14604 (N_14604,N_13560,N_13905);
nand U14605 (N_14605,N_13957,N_13947);
and U14606 (N_14606,N_13545,N_13303);
nor U14607 (N_14607,N_13052,N_13554);
nor U14608 (N_14608,N_13918,N_13221);
and U14609 (N_14609,N_13300,N_13232);
and U14610 (N_14610,N_13298,N_13443);
nand U14611 (N_14611,N_13646,N_13616);
and U14612 (N_14612,N_13514,N_13660);
or U14613 (N_14613,N_13887,N_13478);
or U14614 (N_14614,N_13599,N_13841);
nor U14615 (N_14615,N_13036,N_13619);
nor U14616 (N_14616,N_13874,N_13705);
or U14617 (N_14617,N_13111,N_13873);
xor U14618 (N_14618,N_13897,N_13744);
nor U14619 (N_14619,N_13754,N_13508);
and U14620 (N_14620,N_13669,N_13748);
or U14621 (N_14621,N_13988,N_13089);
nor U14622 (N_14622,N_13371,N_13643);
nor U14623 (N_14623,N_13512,N_13293);
nor U14624 (N_14624,N_13066,N_13127);
xor U14625 (N_14625,N_13357,N_13566);
or U14626 (N_14626,N_13968,N_13980);
xnor U14627 (N_14627,N_13514,N_13349);
or U14628 (N_14628,N_13296,N_13299);
xor U14629 (N_14629,N_13844,N_13490);
nand U14630 (N_14630,N_13338,N_13496);
and U14631 (N_14631,N_13400,N_13526);
nand U14632 (N_14632,N_13422,N_13939);
and U14633 (N_14633,N_13683,N_13624);
and U14634 (N_14634,N_13759,N_13314);
and U14635 (N_14635,N_13500,N_13729);
or U14636 (N_14636,N_13601,N_13524);
nand U14637 (N_14637,N_13894,N_13238);
and U14638 (N_14638,N_13028,N_13341);
nand U14639 (N_14639,N_13116,N_13960);
xor U14640 (N_14640,N_13685,N_13793);
nor U14641 (N_14641,N_13464,N_13442);
nor U14642 (N_14642,N_13623,N_13943);
or U14643 (N_14643,N_13684,N_13264);
xnor U14644 (N_14644,N_13248,N_13105);
or U14645 (N_14645,N_13262,N_13848);
xnor U14646 (N_14646,N_13123,N_13577);
xnor U14647 (N_14647,N_13309,N_13743);
nor U14648 (N_14648,N_13204,N_13537);
or U14649 (N_14649,N_13800,N_13348);
xnor U14650 (N_14650,N_13571,N_13170);
or U14651 (N_14651,N_13994,N_13568);
nand U14652 (N_14652,N_13563,N_13186);
nand U14653 (N_14653,N_13041,N_13654);
and U14654 (N_14654,N_13462,N_13598);
nor U14655 (N_14655,N_13352,N_13220);
and U14656 (N_14656,N_13065,N_13327);
and U14657 (N_14657,N_13410,N_13466);
nor U14658 (N_14658,N_13737,N_13376);
or U14659 (N_14659,N_13219,N_13090);
or U14660 (N_14660,N_13320,N_13359);
nor U14661 (N_14661,N_13257,N_13376);
nand U14662 (N_14662,N_13619,N_13763);
nand U14663 (N_14663,N_13914,N_13855);
nor U14664 (N_14664,N_13470,N_13130);
nand U14665 (N_14665,N_13908,N_13485);
xnor U14666 (N_14666,N_13237,N_13189);
nand U14667 (N_14667,N_13749,N_13565);
or U14668 (N_14668,N_13026,N_13319);
nand U14669 (N_14669,N_13551,N_13318);
nor U14670 (N_14670,N_13004,N_13610);
and U14671 (N_14671,N_13415,N_13432);
xor U14672 (N_14672,N_13419,N_13186);
and U14673 (N_14673,N_13896,N_13003);
nor U14674 (N_14674,N_13519,N_13790);
and U14675 (N_14675,N_13545,N_13998);
nor U14676 (N_14676,N_13723,N_13702);
xnor U14677 (N_14677,N_13780,N_13886);
nor U14678 (N_14678,N_13301,N_13436);
xnor U14679 (N_14679,N_13613,N_13742);
or U14680 (N_14680,N_13986,N_13497);
or U14681 (N_14681,N_13208,N_13996);
or U14682 (N_14682,N_13701,N_13109);
nand U14683 (N_14683,N_13212,N_13011);
nand U14684 (N_14684,N_13083,N_13060);
and U14685 (N_14685,N_13733,N_13919);
nor U14686 (N_14686,N_13738,N_13833);
nor U14687 (N_14687,N_13420,N_13152);
and U14688 (N_14688,N_13176,N_13453);
xnor U14689 (N_14689,N_13555,N_13723);
xnor U14690 (N_14690,N_13607,N_13123);
nand U14691 (N_14691,N_13125,N_13034);
nor U14692 (N_14692,N_13903,N_13652);
and U14693 (N_14693,N_13049,N_13166);
nand U14694 (N_14694,N_13805,N_13203);
nor U14695 (N_14695,N_13150,N_13175);
nand U14696 (N_14696,N_13189,N_13421);
or U14697 (N_14697,N_13666,N_13526);
xnor U14698 (N_14698,N_13935,N_13209);
nand U14699 (N_14699,N_13862,N_13766);
or U14700 (N_14700,N_13202,N_13191);
or U14701 (N_14701,N_13627,N_13868);
nor U14702 (N_14702,N_13580,N_13172);
or U14703 (N_14703,N_13235,N_13748);
nand U14704 (N_14704,N_13258,N_13183);
nand U14705 (N_14705,N_13122,N_13867);
xor U14706 (N_14706,N_13204,N_13855);
or U14707 (N_14707,N_13460,N_13150);
nor U14708 (N_14708,N_13262,N_13267);
nand U14709 (N_14709,N_13249,N_13940);
nand U14710 (N_14710,N_13585,N_13857);
nor U14711 (N_14711,N_13464,N_13510);
nor U14712 (N_14712,N_13819,N_13390);
xnor U14713 (N_14713,N_13876,N_13926);
xor U14714 (N_14714,N_13585,N_13407);
nand U14715 (N_14715,N_13630,N_13773);
nor U14716 (N_14716,N_13359,N_13938);
nand U14717 (N_14717,N_13568,N_13884);
nor U14718 (N_14718,N_13323,N_13833);
or U14719 (N_14719,N_13355,N_13493);
xnor U14720 (N_14720,N_13895,N_13940);
nand U14721 (N_14721,N_13802,N_13465);
nor U14722 (N_14722,N_13996,N_13534);
xor U14723 (N_14723,N_13582,N_13543);
and U14724 (N_14724,N_13073,N_13246);
nand U14725 (N_14725,N_13538,N_13823);
or U14726 (N_14726,N_13652,N_13356);
xor U14727 (N_14727,N_13679,N_13851);
and U14728 (N_14728,N_13355,N_13956);
nand U14729 (N_14729,N_13571,N_13695);
or U14730 (N_14730,N_13793,N_13402);
xor U14731 (N_14731,N_13067,N_13372);
or U14732 (N_14732,N_13816,N_13119);
xnor U14733 (N_14733,N_13977,N_13407);
nor U14734 (N_14734,N_13938,N_13561);
nor U14735 (N_14735,N_13602,N_13154);
nor U14736 (N_14736,N_13243,N_13030);
nor U14737 (N_14737,N_13318,N_13285);
nand U14738 (N_14738,N_13876,N_13772);
xnor U14739 (N_14739,N_13678,N_13419);
xor U14740 (N_14740,N_13037,N_13545);
nand U14741 (N_14741,N_13324,N_13497);
nor U14742 (N_14742,N_13350,N_13822);
or U14743 (N_14743,N_13045,N_13464);
nor U14744 (N_14744,N_13206,N_13018);
xnor U14745 (N_14745,N_13772,N_13884);
or U14746 (N_14746,N_13285,N_13416);
and U14747 (N_14747,N_13382,N_13512);
xnor U14748 (N_14748,N_13048,N_13582);
nand U14749 (N_14749,N_13188,N_13612);
xor U14750 (N_14750,N_13985,N_13710);
nand U14751 (N_14751,N_13265,N_13152);
or U14752 (N_14752,N_13170,N_13879);
nor U14753 (N_14753,N_13740,N_13524);
nand U14754 (N_14754,N_13966,N_13125);
or U14755 (N_14755,N_13344,N_13870);
or U14756 (N_14756,N_13440,N_13091);
and U14757 (N_14757,N_13654,N_13950);
and U14758 (N_14758,N_13468,N_13769);
nor U14759 (N_14759,N_13260,N_13360);
and U14760 (N_14760,N_13767,N_13260);
xor U14761 (N_14761,N_13080,N_13217);
nand U14762 (N_14762,N_13657,N_13166);
and U14763 (N_14763,N_13777,N_13994);
xor U14764 (N_14764,N_13542,N_13254);
and U14765 (N_14765,N_13826,N_13853);
and U14766 (N_14766,N_13131,N_13287);
and U14767 (N_14767,N_13558,N_13983);
nor U14768 (N_14768,N_13783,N_13893);
xor U14769 (N_14769,N_13891,N_13557);
nor U14770 (N_14770,N_13059,N_13115);
nand U14771 (N_14771,N_13318,N_13544);
nor U14772 (N_14772,N_13666,N_13825);
and U14773 (N_14773,N_13759,N_13473);
and U14774 (N_14774,N_13975,N_13500);
or U14775 (N_14775,N_13020,N_13806);
xnor U14776 (N_14776,N_13830,N_13475);
nand U14777 (N_14777,N_13993,N_13917);
and U14778 (N_14778,N_13217,N_13774);
nand U14779 (N_14779,N_13406,N_13806);
nor U14780 (N_14780,N_13216,N_13954);
xnor U14781 (N_14781,N_13125,N_13585);
nand U14782 (N_14782,N_13536,N_13617);
nand U14783 (N_14783,N_13861,N_13614);
xor U14784 (N_14784,N_13626,N_13455);
or U14785 (N_14785,N_13974,N_13966);
xnor U14786 (N_14786,N_13107,N_13338);
and U14787 (N_14787,N_13515,N_13536);
or U14788 (N_14788,N_13166,N_13116);
or U14789 (N_14789,N_13778,N_13317);
nand U14790 (N_14790,N_13976,N_13730);
and U14791 (N_14791,N_13273,N_13996);
or U14792 (N_14792,N_13614,N_13566);
and U14793 (N_14793,N_13616,N_13526);
and U14794 (N_14794,N_13949,N_13767);
nor U14795 (N_14795,N_13364,N_13824);
or U14796 (N_14796,N_13494,N_13004);
nand U14797 (N_14797,N_13926,N_13269);
nor U14798 (N_14798,N_13226,N_13944);
nand U14799 (N_14799,N_13622,N_13819);
and U14800 (N_14800,N_13921,N_13829);
and U14801 (N_14801,N_13345,N_13752);
or U14802 (N_14802,N_13755,N_13982);
xor U14803 (N_14803,N_13582,N_13812);
and U14804 (N_14804,N_13522,N_13393);
and U14805 (N_14805,N_13154,N_13712);
or U14806 (N_14806,N_13504,N_13801);
or U14807 (N_14807,N_13217,N_13758);
and U14808 (N_14808,N_13286,N_13510);
nand U14809 (N_14809,N_13698,N_13052);
or U14810 (N_14810,N_13895,N_13380);
or U14811 (N_14811,N_13685,N_13231);
or U14812 (N_14812,N_13704,N_13199);
and U14813 (N_14813,N_13879,N_13412);
and U14814 (N_14814,N_13763,N_13914);
xor U14815 (N_14815,N_13782,N_13622);
nand U14816 (N_14816,N_13513,N_13986);
xor U14817 (N_14817,N_13993,N_13718);
nand U14818 (N_14818,N_13139,N_13633);
xnor U14819 (N_14819,N_13190,N_13355);
or U14820 (N_14820,N_13955,N_13283);
xnor U14821 (N_14821,N_13401,N_13738);
and U14822 (N_14822,N_13043,N_13978);
nor U14823 (N_14823,N_13832,N_13078);
xnor U14824 (N_14824,N_13396,N_13586);
and U14825 (N_14825,N_13119,N_13263);
nor U14826 (N_14826,N_13370,N_13326);
and U14827 (N_14827,N_13271,N_13535);
xor U14828 (N_14828,N_13845,N_13082);
and U14829 (N_14829,N_13264,N_13501);
or U14830 (N_14830,N_13415,N_13488);
nor U14831 (N_14831,N_13417,N_13853);
xor U14832 (N_14832,N_13102,N_13037);
nor U14833 (N_14833,N_13680,N_13671);
nand U14834 (N_14834,N_13762,N_13554);
and U14835 (N_14835,N_13749,N_13360);
xnor U14836 (N_14836,N_13887,N_13858);
xor U14837 (N_14837,N_13495,N_13343);
nand U14838 (N_14838,N_13600,N_13369);
nand U14839 (N_14839,N_13068,N_13709);
or U14840 (N_14840,N_13479,N_13211);
nor U14841 (N_14841,N_13636,N_13016);
nor U14842 (N_14842,N_13142,N_13913);
nor U14843 (N_14843,N_13873,N_13692);
nand U14844 (N_14844,N_13124,N_13224);
nor U14845 (N_14845,N_13177,N_13482);
nand U14846 (N_14846,N_13233,N_13763);
xnor U14847 (N_14847,N_13880,N_13657);
nand U14848 (N_14848,N_13367,N_13039);
and U14849 (N_14849,N_13349,N_13709);
or U14850 (N_14850,N_13013,N_13860);
and U14851 (N_14851,N_13532,N_13062);
xor U14852 (N_14852,N_13882,N_13964);
or U14853 (N_14853,N_13808,N_13763);
nor U14854 (N_14854,N_13478,N_13077);
nor U14855 (N_14855,N_13442,N_13202);
and U14856 (N_14856,N_13447,N_13335);
xor U14857 (N_14857,N_13314,N_13085);
nand U14858 (N_14858,N_13434,N_13849);
nor U14859 (N_14859,N_13291,N_13136);
xnor U14860 (N_14860,N_13625,N_13377);
nand U14861 (N_14861,N_13819,N_13459);
xnor U14862 (N_14862,N_13575,N_13085);
nor U14863 (N_14863,N_13975,N_13571);
nand U14864 (N_14864,N_13161,N_13409);
and U14865 (N_14865,N_13682,N_13179);
xnor U14866 (N_14866,N_13373,N_13705);
nor U14867 (N_14867,N_13661,N_13071);
and U14868 (N_14868,N_13736,N_13531);
or U14869 (N_14869,N_13440,N_13397);
or U14870 (N_14870,N_13117,N_13175);
nor U14871 (N_14871,N_13878,N_13829);
and U14872 (N_14872,N_13596,N_13974);
nand U14873 (N_14873,N_13539,N_13141);
xnor U14874 (N_14874,N_13747,N_13191);
xnor U14875 (N_14875,N_13801,N_13145);
xor U14876 (N_14876,N_13199,N_13003);
xnor U14877 (N_14877,N_13413,N_13280);
nand U14878 (N_14878,N_13172,N_13326);
nor U14879 (N_14879,N_13505,N_13468);
nand U14880 (N_14880,N_13983,N_13902);
and U14881 (N_14881,N_13840,N_13428);
nor U14882 (N_14882,N_13903,N_13894);
xor U14883 (N_14883,N_13222,N_13655);
nor U14884 (N_14884,N_13685,N_13225);
xor U14885 (N_14885,N_13435,N_13111);
nor U14886 (N_14886,N_13545,N_13585);
nor U14887 (N_14887,N_13566,N_13414);
xor U14888 (N_14888,N_13142,N_13752);
nand U14889 (N_14889,N_13512,N_13804);
nor U14890 (N_14890,N_13930,N_13891);
xnor U14891 (N_14891,N_13197,N_13253);
nor U14892 (N_14892,N_13407,N_13293);
and U14893 (N_14893,N_13869,N_13261);
and U14894 (N_14894,N_13001,N_13852);
nand U14895 (N_14895,N_13134,N_13188);
xor U14896 (N_14896,N_13953,N_13944);
xnor U14897 (N_14897,N_13304,N_13981);
xnor U14898 (N_14898,N_13548,N_13619);
nor U14899 (N_14899,N_13924,N_13395);
nand U14900 (N_14900,N_13140,N_13369);
nor U14901 (N_14901,N_13538,N_13573);
nor U14902 (N_14902,N_13650,N_13933);
and U14903 (N_14903,N_13502,N_13552);
and U14904 (N_14904,N_13511,N_13784);
xnor U14905 (N_14905,N_13987,N_13204);
nor U14906 (N_14906,N_13272,N_13510);
and U14907 (N_14907,N_13520,N_13572);
nand U14908 (N_14908,N_13932,N_13672);
nand U14909 (N_14909,N_13647,N_13005);
xor U14910 (N_14910,N_13122,N_13312);
nor U14911 (N_14911,N_13886,N_13107);
nand U14912 (N_14912,N_13719,N_13031);
xnor U14913 (N_14913,N_13831,N_13998);
and U14914 (N_14914,N_13605,N_13580);
xnor U14915 (N_14915,N_13345,N_13482);
xnor U14916 (N_14916,N_13303,N_13490);
or U14917 (N_14917,N_13587,N_13720);
xor U14918 (N_14918,N_13880,N_13464);
nand U14919 (N_14919,N_13230,N_13254);
nand U14920 (N_14920,N_13374,N_13690);
and U14921 (N_14921,N_13361,N_13647);
or U14922 (N_14922,N_13407,N_13119);
and U14923 (N_14923,N_13754,N_13606);
nand U14924 (N_14924,N_13412,N_13334);
nand U14925 (N_14925,N_13346,N_13675);
nor U14926 (N_14926,N_13867,N_13165);
and U14927 (N_14927,N_13477,N_13125);
xnor U14928 (N_14928,N_13460,N_13063);
nor U14929 (N_14929,N_13607,N_13964);
nor U14930 (N_14930,N_13357,N_13327);
nor U14931 (N_14931,N_13257,N_13628);
and U14932 (N_14932,N_13784,N_13937);
and U14933 (N_14933,N_13841,N_13906);
nand U14934 (N_14934,N_13886,N_13883);
and U14935 (N_14935,N_13171,N_13205);
nor U14936 (N_14936,N_13101,N_13204);
and U14937 (N_14937,N_13082,N_13505);
nor U14938 (N_14938,N_13029,N_13385);
and U14939 (N_14939,N_13621,N_13117);
nand U14940 (N_14940,N_13684,N_13132);
and U14941 (N_14941,N_13259,N_13363);
and U14942 (N_14942,N_13784,N_13785);
or U14943 (N_14943,N_13916,N_13165);
nor U14944 (N_14944,N_13096,N_13599);
xnor U14945 (N_14945,N_13594,N_13153);
nor U14946 (N_14946,N_13288,N_13361);
and U14947 (N_14947,N_13731,N_13594);
xor U14948 (N_14948,N_13027,N_13696);
nand U14949 (N_14949,N_13917,N_13604);
nor U14950 (N_14950,N_13193,N_13881);
nand U14951 (N_14951,N_13184,N_13104);
and U14952 (N_14952,N_13931,N_13466);
nand U14953 (N_14953,N_13632,N_13303);
and U14954 (N_14954,N_13734,N_13836);
xnor U14955 (N_14955,N_13895,N_13937);
and U14956 (N_14956,N_13470,N_13966);
xor U14957 (N_14957,N_13428,N_13678);
or U14958 (N_14958,N_13836,N_13171);
nand U14959 (N_14959,N_13943,N_13067);
and U14960 (N_14960,N_13797,N_13555);
nor U14961 (N_14961,N_13016,N_13692);
or U14962 (N_14962,N_13820,N_13741);
xnor U14963 (N_14963,N_13917,N_13425);
nand U14964 (N_14964,N_13402,N_13725);
nand U14965 (N_14965,N_13863,N_13421);
or U14966 (N_14966,N_13098,N_13595);
xnor U14967 (N_14967,N_13041,N_13970);
xnor U14968 (N_14968,N_13857,N_13570);
and U14969 (N_14969,N_13761,N_13073);
or U14970 (N_14970,N_13332,N_13733);
nor U14971 (N_14971,N_13993,N_13811);
and U14972 (N_14972,N_13543,N_13488);
xnor U14973 (N_14973,N_13493,N_13549);
and U14974 (N_14974,N_13052,N_13280);
nand U14975 (N_14975,N_13242,N_13593);
xor U14976 (N_14976,N_13702,N_13822);
nand U14977 (N_14977,N_13081,N_13896);
nand U14978 (N_14978,N_13103,N_13666);
or U14979 (N_14979,N_13945,N_13905);
xnor U14980 (N_14980,N_13580,N_13961);
or U14981 (N_14981,N_13086,N_13822);
xnor U14982 (N_14982,N_13463,N_13900);
xor U14983 (N_14983,N_13664,N_13419);
xor U14984 (N_14984,N_13668,N_13556);
nor U14985 (N_14985,N_13280,N_13638);
nand U14986 (N_14986,N_13218,N_13869);
nand U14987 (N_14987,N_13996,N_13524);
nand U14988 (N_14988,N_13184,N_13705);
xor U14989 (N_14989,N_13628,N_13077);
xor U14990 (N_14990,N_13913,N_13733);
or U14991 (N_14991,N_13292,N_13536);
or U14992 (N_14992,N_13411,N_13760);
nor U14993 (N_14993,N_13047,N_13197);
xor U14994 (N_14994,N_13518,N_13596);
nor U14995 (N_14995,N_13148,N_13236);
nand U14996 (N_14996,N_13615,N_13234);
nand U14997 (N_14997,N_13573,N_13396);
or U14998 (N_14998,N_13795,N_13581);
and U14999 (N_14999,N_13506,N_13910);
xor U15000 (N_15000,N_14878,N_14472);
xnor U15001 (N_15001,N_14858,N_14937);
or U15002 (N_15002,N_14998,N_14514);
nand U15003 (N_15003,N_14535,N_14265);
and U15004 (N_15004,N_14188,N_14690);
or U15005 (N_15005,N_14442,N_14641);
nand U15006 (N_15006,N_14577,N_14439);
and U15007 (N_15007,N_14278,N_14488);
and U15008 (N_15008,N_14664,N_14213);
and U15009 (N_15009,N_14525,N_14899);
nor U15010 (N_15010,N_14548,N_14801);
and U15011 (N_15011,N_14348,N_14350);
nor U15012 (N_15012,N_14663,N_14087);
nand U15013 (N_15013,N_14136,N_14179);
or U15014 (N_15014,N_14702,N_14571);
or U15015 (N_15015,N_14028,N_14304);
xnor U15016 (N_15016,N_14709,N_14695);
xnor U15017 (N_15017,N_14845,N_14515);
nand U15018 (N_15018,N_14119,N_14673);
or U15019 (N_15019,N_14569,N_14629);
nand U15020 (N_15020,N_14961,N_14250);
nor U15021 (N_15021,N_14008,N_14814);
xor U15022 (N_15022,N_14681,N_14753);
or U15023 (N_15023,N_14138,N_14716);
or U15024 (N_15024,N_14780,N_14026);
or U15025 (N_15025,N_14286,N_14077);
or U15026 (N_15026,N_14643,N_14881);
nand U15027 (N_15027,N_14254,N_14052);
xnor U15028 (N_15028,N_14965,N_14579);
xnor U15029 (N_15029,N_14104,N_14169);
nor U15030 (N_15030,N_14076,N_14595);
nand U15031 (N_15031,N_14870,N_14591);
or U15032 (N_15032,N_14742,N_14366);
or U15033 (N_15033,N_14701,N_14612);
or U15034 (N_15034,N_14996,N_14691);
or U15035 (N_15035,N_14649,N_14338);
xor U15036 (N_15036,N_14640,N_14380);
or U15037 (N_15037,N_14171,N_14270);
nor U15038 (N_15038,N_14703,N_14602);
and U15039 (N_15039,N_14167,N_14279);
and U15040 (N_15040,N_14575,N_14345);
or U15041 (N_15041,N_14693,N_14244);
nor U15042 (N_15042,N_14872,N_14971);
nand U15043 (N_15043,N_14409,N_14337);
or U15044 (N_15044,N_14622,N_14538);
xor U15045 (N_15045,N_14420,N_14769);
nand U15046 (N_15046,N_14053,N_14465);
or U15047 (N_15047,N_14853,N_14717);
or U15048 (N_15048,N_14707,N_14658);
and U15049 (N_15049,N_14929,N_14540);
nor U15050 (N_15050,N_14372,N_14137);
nand U15051 (N_15051,N_14726,N_14711);
nand U15052 (N_15052,N_14837,N_14761);
and U15053 (N_15053,N_14947,N_14125);
or U15054 (N_15054,N_14386,N_14978);
nand U15055 (N_15055,N_14782,N_14039);
nor U15056 (N_15056,N_14257,N_14309);
xnor U15057 (N_15057,N_14061,N_14071);
xnor U15058 (N_15058,N_14308,N_14745);
or U15059 (N_15059,N_14223,N_14128);
nor U15060 (N_15060,N_14048,N_14666);
nor U15061 (N_15061,N_14009,N_14486);
xnor U15062 (N_15062,N_14100,N_14470);
xnor U15063 (N_15063,N_14868,N_14075);
nor U15064 (N_15064,N_14564,N_14850);
nand U15065 (N_15065,N_14124,N_14245);
and U15066 (N_15066,N_14995,N_14820);
or U15067 (N_15067,N_14299,N_14408);
xor U15068 (N_15068,N_14434,N_14404);
or U15069 (N_15069,N_14976,N_14297);
nor U15070 (N_15070,N_14558,N_14949);
and U15071 (N_15071,N_14143,N_14480);
or U15072 (N_15072,N_14598,N_14093);
xnor U15073 (N_15073,N_14054,N_14997);
or U15074 (N_15074,N_14960,N_14799);
xnor U15075 (N_15075,N_14990,N_14594);
or U15076 (N_15076,N_14865,N_14301);
and U15077 (N_15077,N_14530,N_14802);
nand U15078 (N_15078,N_14553,N_14552);
nand U15079 (N_15079,N_14962,N_14029);
xnor U15080 (N_15080,N_14199,N_14583);
nand U15081 (N_15081,N_14477,N_14628);
nor U15082 (N_15082,N_14163,N_14164);
nand U15083 (N_15083,N_14444,N_14060);
and U15084 (N_15084,N_14202,N_14980);
nand U15085 (N_15085,N_14102,N_14925);
and U15086 (N_15086,N_14776,N_14954);
xor U15087 (N_15087,N_14050,N_14534);
xnor U15088 (N_15088,N_14344,N_14280);
xor U15089 (N_15089,N_14021,N_14118);
and U15090 (N_15090,N_14375,N_14400);
nand U15091 (N_15091,N_14362,N_14633);
xor U15092 (N_15092,N_14310,N_14051);
and U15093 (N_15093,N_14792,N_14522);
or U15094 (N_15094,N_14547,N_14618);
and U15095 (N_15095,N_14098,N_14632);
or U15096 (N_15096,N_14490,N_14927);
nand U15097 (N_15097,N_14388,N_14267);
nand U15098 (N_15098,N_14959,N_14296);
and U15099 (N_15099,N_14590,N_14221);
nand U15100 (N_15100,N_14469,N_14336);
nor U15101 (N_15101,N_14183,N_14032);
and U15102 (N_15102,N_14821,N_14011);
xnor U15103 (N_15103,N_14023,N_14003);
and U15104 (N_15104,N_14110,N_14824);
nor U15105 (N_15105,N_14974,N_14127);
nand U15106 (N_15106,N_14610,N_14706);
nor U15107 (N_15107,N_14920,N_14638);
xor U15108 (N_15108,N_14678,N_14361);
xnor U15109 (N_15109,N_14004,N_14405);
nor U15110 (N_15110,N_14047,N_14207);
nand U15111 (N_15111,N_14097,N_14580);
nor U15112 (N_15112,N_14750,N_14479);
or U15113 (N_15113,N_14608,N_14027);
nor U15114 (N_15114,N_14928,N_14222);
nand U15115 (N_15115,N_14787,N_14812);
or U15116 (N_15116,N_14290,N_14190);
xnor U15117 (N_15117,N_14732,N_14363);
or U15118 (N_15118,N_14563,N_14392);
and U15119 (N_15119,N_14603,N_14680);
and U15120 (N_15120,N_14121,N_14091);
or U15121 (N_15121,N_14880,N_14172);
xnor U15122 (N_15122,N_14274,N_14305);
or U15123 (N_15123,N_14253,N_14752);
nor U15124 (N_15124,N_14228,N_14421);
or U15125 (N_15125,N_14161,N_14034);
nand U15126 (N_15126,N_14911,N_14945);
xor U15127 (N_15127,N_14331,N_14891);
xnor U15128 (N_15128,N_14260,N_14330);
and U15129 (N_15129,N_14746,N_14148);
and U15130 (N_15130,N_14166,N_14539);
nand U15131 (N_15131,N_14294,N_14651);
xor U15132 (N_15132,N_14625,N_14120);
nor U15133 (N_15133,N_14191,N_14374);
nand U15134 (N_15134,N_14587,N_14645);
and U15135 (N_15135,N_14243,N_14289);
and U15136 (N_15136,N_14939,N_14885);
xor U15137 (N_15137,N_14755,N_14617);
and U15138 (N_15138,N_14454,N_14378);
xnor U15139 (N_15139,N_14144,N_14869);
nor U15140 (N_15140,N_14342,N_14777);
nand U15141 (N_15141,N_14614,N_14074);
xor U15142 (N_15142,N_14145,N_14770);
xor U15143 (N_15143,N_14201,N_14528);
nor U15144 (N_15144,N_14391,N_14482);
xor U15145 (N_15145,N_14655,N_14358);
and U15146 (N_15146,N_14266,N_14578);
and U15147 (N_15147,N_14227,N_14063);
nor U15148 (N_15148,N_14926,N_14963);
or U15149 (N_15149,N_14284,N_14269);
xnor U15150 (N_15150,N_14857,N_14133);
nor U15151 (N_15151,N_14807,N_14537);
xnor U15152 (N_15152,N_14012,N_14854);
and U15153 (N_15153,N_14679,N_14197);
xnor U15154 (N_15154,N_14355,N_14401);
and U15155 (N_15155,N_14365,N_14674);
nor U15156 (N_15156,N_14452,N_14943);
nor U15157 (N_15157,N_14830,N_14554);
nor U15158 (N_15158,N_14533,N_14735);
nor U15159 (N_15159,N_14057,N_14806);
nand U15160 (N_15160,N_14886,N_14462);
and U15161 (N_15161,N_14433,N_14379);
xnor U15162 (N_15162,N_14123,N_14968);
nand U15163 (N_15163,N_14767,N_14083);
xor U15164 (N_15164,N_14696,N_14248);
and U15165 (N_15165,N_14653,N_14644);
or U15166 (N_15166,N_14018,N_14500);
or U15167 (N_15167,N_14080,N_14036);
and U15168 (N_15168,N_14605,N_14017);
or U15169 (N_15169,N_14852,N_14209);
xor U15170 (N_15170,N_14743,N_14985);
and U15171 (N_15171,N_14252,N_14065);
or U15172 (N_15172,N_14423,N_14217);
nand U15173 (N_15173,N_14323,N_14417);
nand U15174 (N_15174,N_14210,N_14727);
nand U15175 (N_15175,N_14892,N_14182);
xor U15176 (N_15176,N_14883,N_14152);
nand U15177 (N_15177,N_14263,N_14038);
nand U15178 (N_15178,N_14156,N_14347);
nand U15179 (N_15179,N_14668,N_14520);
nor U15180 (N_15180,N_14768,N_14849);
nor U15181 (N_15181,N_14736,N_14991);
or U15182 (N_15182,N_14131,N_14446);
xor U15183 (N_15183,N_14975,N_14095);
nand U15184 (N_15184,N_14982,N_14001);
or U15185 (N_15185,N_14030,N_14352);
and U15186 (N_15186,N_14863,N_14069);
xnor U15187 (N_15187,N_14196,N_14509);
nor U15188 (N_15188,N_14271,N_14597);
xor U15189 (N_15189,N_14897,N_14329);
or U15190 (N_15190,N_14198,N_14627);
xnor U15191 (N_15191,N_14112,N_14403);
and U15192 (N_15192,N_14316,N_14983);
nor U15193 (N_15193,N_14848,N_14831);
and U15194 (N_15194,N_14778,N_14715);
and U15195 (N_15195,N_14445,N_14635);
nand U15196 (N_15196,N_14654,N_14382);
and U15197 (N_15197,N_14957,N_14946);
and U15198 (N_15198,N_14122,N_14238);
and U15199 (N_15199,N_14114,N_14970);
xnor U15200 (N_15200,N_14942,N_14451);
nand U15201 (N_15201,N_14804,N_14557);
nand U15202 (N_15202,N_14178,N_14295);
and U15203 (N_15203,N_14239,N_14321);
xnor U15204 (N_15204,N_14904,N_14896);
or U15205 (N_15205,N_14541,N_14312);
xor U15206 (N_15206,N_14428,N_14613);
nand U15207 (N_15207,N_14411,N_14019);
or U15208 (N_15208,N_14272,N_14035);
or U15209 (N_15209,N_14619,N_14022);
nor U15210 (N_15210,N_14879,N_14670);
and U15211 (N_15211,N_14549,N_14399);
nand U15212 (N_15212,N_14322,N_14986);
or U15213 (N_15213,N_14934,N_14773);
or U15214 (N_15214,N_14532,N_14418);
nor U15215 (N_15215,N_14758,N_14556);
xnor U15216 (N_15216,N_14431,N_14484);
nor U15217 (N_15217,N_14785,N_14453);
nand U15218 (N_15218,N_14842,N_14893);
xor U15219 (N_15219,N_14958,N_14841);
nor U15220 (N_15220,N_14206,N_14165);
nor U15221 (N_15221,N_14684,N_14987);
nand U15222 (N_15222,N_14024,N_14364);
nor U15223 (N_15223,N_14694,N_14918);
xor U15224 (N_15224,N_14458,N_14461);
and U15225 (N_15225,N_14573,N_14456);
nand U15226 (N_15226,N_14059,N_14040);
nand U15227 (N_15227,N_14584,N_14818);
xnor U15228 (N_15228,N_14952,N_14449);
nand U15229 (N_15229,N_14944,N_14220);
nand U15230 (N_15230,N_14994,N_14231);
xor U15231 (N_15231,N_14713,N_14218);
xnor U15232 (N_15232,N_14318,N_14977);
and U15233 (N_15233,N_14236,N_14874);
nor U15234 (N_15234,N_14734,N_14676);
nand U15235 (N_15235,N_14055,N_14705);
or U15236 (N_15236,N_14168,N_14682);
xor U15237 (N_15237,N_14073,N_14828);
nor U15238 (N_15238,N_14771,N_14407);
and U15239 (N_15239,N_14793,N_14789);
or U15240 (N_15240,N_14692,N_14173);
or U15241 (N_15241,N_14887,N_14543);
nand U15242 (N_15242,N_14459,N_14393);
and U15243 (N_15243,N_14314,N_14287);
or U15244 (N_15244,N_14313,N_14176);
and U15245 (N_15245,N_14941,N_14056);
nand U15246 (N_15246,N_14013,N_14630);
nor U15247 (N_15247,N_14846,N_14839);
and U15248 (N_15248,N_14216,N_14795);
or U15249 (N_15249,N_14699,N_14468);
nand U15250 (N_15250,N_14636,N_14650);
nand U15251 (N_15251,N_14607,N_14066);
nand U15252 (N_15252,N_14599,N_14096);
nand U15253 (N_15253,N_14187,N_14246);
xnor U15254 (N_15254,N_14744,N_14276);
or U15255 (N_15255,N_14800,N_14416);
xor U15256 (N_15256,N_14268,N_14389);
nor U15257 (N_15257,N_14819,N_14910);
or U15258 (N_15258,N_14835,N_14387);
and U15259 (N_15259,N_14130,N_14760);
and U15260 (N_15260,N_14988,N_14147);
xor U15261 (N_15261,N_14720,N_14425);
nor U15262 (N_15262,N_14448,N_14808);
or U15263 (N_15263,N_14495,N_14510);
or U15264 (N_15264,N_14142,N_14798);
xnor U15265 (N_15265,N_14476,N_14058);
nor U15266 (N_15266,N_14647,N_14981);
nand U15267 (N_15267,N_14240,N_14085);
and U15268 (N_15268,N_14501,N_14346);
xnor U15269 (N_15269,N_14508,N_14581);
nor U15270 (N_15270,N_14162,N_14150);
xor U15271 (N_15271,N_14483,N_14786);
nor U15272 (N_15272,N_14412,N_14621);
nand U15273 (N_15273,N_14235,N_14545);
nor U15274 (N_15274,N_14157,N_14894);
or U15275 (N_15275,N_14840,N_14261);
and U15276 (N_15276,N_14247,N_14672);
nand U15277 (N_15277,N_14797,N_14328);
xor U15278 (N_15278,N_14567,N_14396);
or U15279 (N_15279,N_14908,N_14205);
nand U15280 (N_15280,N_14493,N_14503);
nor U15281 (N_15281,N_14349,N_14419);
nor U15282 (N_15282,N_14049,N_14637);
or U15283 (N_15283,N_14738,N_14566);
and U15284 (N_15284,N_14794,N_14507);
or U15285 (N_15285,N_14394,N_14722);
nand U15286 (N_15286,N_14922,N_14487);
or U15287 (N_15287,N_14115,N_14357);
or U15288 (N_15288,N_14385,N_14914);
nor U15289 (N_15289,N_14989,N_14781);
and U15290 (N_15290,N_14415,N_14611);
nand U15291 (N_15291,N_14596,N_14025);
xnor U15292 (N_15292,N_14436,N_14192);
nand U15293 (N_15293,N_14332,N_14565);
and U15294 (N_15294,N_14273,N_14160);
and U15295 (N_15295,N_14838,N_14721);
nand U15296 (N_15296,N_14950,N_14249);
and U15297 (N_15297,N_14117,N_14135);
and U15298 (N_15298,N_14440,N_14042);
nand U15299 (N_15299,N_14754,N_14282);
xor U15300 (N_15300,N_14531,N_14233);
and U15301 (N_15301,N_14826,N_14642);
xnor U15302 (N_15302,N_14226,N_14311);
xor U15303 (N_15303,N_14572,N_14103);
and U15304 (N_15304,N_14546,N_14241);
or U15305 (N_15305,N_14438,N_14367);
and U15306 (N_15306,N_14652,N_14866);
and U15307 (N_15307,N_14827,N_14570);
xor U15308 (N_15308,N_14370,N_14523);
and U15309 (N_15309,N_14457,N_14327);
and U15310 (N_15310,N_14817,N_14749);
and U15311 (N_15311,N_14764,N_14888);
or U15312 (N_15312,N_14099,N_14876);
and U15313 (N_15313,N_14302,N_14626);
nand U15314 (N_15314,N_14882,N_14158);
nand U15315 (N_15315,N_14474,N_14536);
xnor U15316 (N_15316,N_14710,N_14973);
nand U15317 (N_15317,N_14219,N_14656);
or U15318 (N_15318,N_14551,N_14002);
or U15319 (N_15319,N_14759,N_14146);
nand U15320 (N_15320,N_14725,N_14923);
or U15321 (N_15321,N_14843,N_14810);
and U15322 (N_15322,N_14214,N_14194);
and U15323 (N_15323,N_14341,N_14561);
xnor U15324 (N_15324,N_14498,N_14443);
xor U15325 (N_15325,N_14964,N_14154);
xor U15326 (N_15326,N_14659,N_14984);
nor U15327 (N_15327,N_14813,N_14521);
nor U15328 (N_15328,N_14847,N_14718);
xnor U15329 (N_15329,N_14390,N_14067);
or U15330 (N_15330,N_14262,N_14141);
or U15331 (N_15331,N_14747,N_14657);
nor U15332 (N_15332,N_14519,N_14855);
or U15333 (N_15333,N_14559,N_14719);
and U15334 (N_15334,N_14784,N_14485);
xor U15335 (N_15335,N_14092,N_14860);
nor U15336 (N_15336,N_14938,N_14615);
or U15337 (N_15337,N_14708,N_14140);
and U15338 (N_15338,N_14966,N_14756);
xor U15339 (N_15339,N_14258,N_14397);
or U15340 (N_15340,N_14242,N_14697);
and U15341 (N_15341,N_14285,N_14275);
xor U15342 (N_15342,N_14741,N_14867);
and U15343 (N_15343,N_14862,N_14516);
and U15344 (N_15344,N_14730,N_14829);
nor U15345 (N_15345,N_14478,N_14467);
xnor U15346 (N_15346,N_14951,N_14592);
xnor U15347 (N_15347,N_14105,N_14319);
nor U15348 (N_15348,N_14933,N_14511);
nor U15349 (N_15349,N_14307,N_14757);
nor U15350 (N_15350,N_14502,N_14422);
and U15351 (N_15351,N_14291,N_14335);
and U15352 (N_15352,N_14739,N_14832);
xor U15353 (N_15353,N_14953,N_14609);
and U15354 (N_15354,N_14139,N_14844);
and U15355 (N_15355,N_14714,N_14373);
xor U15356 (N_15356,N_14203,N_14174);
nand U15357 (N_15357,N_14298,N_14079);
nand U15358 (N_15358,N_14334,N_14212);
and U15359 (N_15359,N_14359,N_14568);
nor U15360 (N_15360,N_14116,N_14687);
and U15361 (N_15361,N_14698,N_14935);
xor U15362 (N_15362,N_14134,N_14689);
nor U15363 (N_15363,N_14512,N_14898);
xnor U15364 (N_15364,N_14072,N_14384);
xor U15365 (N_15365,N_14089,N_14895);
nor U15366 (N_15366,N_14324,N_14661);
nand U15367 (N_15367,N_14620,N_14046);
and U15368 (N_15368,N_14993,N_14326);
xnor U15369 (N_15369,N_14475,N_14129);
nand U15370 (N_15370,N_14410,N_14921);
nor U15371 (N_15371,N_14671,N_14159);
and U15372 (N_15372,N_14700,N_14413);
or U15373 (N_15373,N_14070,N_14731);
or U15374 (N_15374,N_14940,N_14779);
and U15375 (N_15375,N_14429,N_14224);
nand U15376 (N_15376,N_14489,N_14936);
xor U15377 (N_15377,N_14772,N_14177);
xor U15378 (N_15378,N_14729,N_14712);
nor U15379 (N_15379,N_14014,N_14232);
or U15380 (N_15380,N_14504,N_14234);
xnor U15381 (N_15381,N_14109,N_14082);
or U15382 (N_15382,N_14437,N_14081);
xnor U15383 (N_15383,N_14353,N_14460);
nor U15384 (N_15384,N_14306,N_14343);
nand U15385 (N_15385,N_14424,N_14185);
nand U15386 (N_15386,N_14704,N_14907);
xnor U15387 (N_15387,N_14441,N_14809);
nor U15388 (N_15388,N_14293,N_14499);
and U15389 (N_15389,N_14170,N_14873);
nand U15390 (N_15390,N_14288,N_14916);
or U15391 (N_15391,N_14524,N_14588);
or U15392 (N_15392,N_14277,N_14631);
nand U15393 (N_15393,N_14186,N_14251);
xor U15394 (N_15394,N_14932,N_14010);
nor U15395 (N_15395,N_14015,N_14041);
and U15396 (N_15396,N_14601,N_14016);
nand U15397 (N_15397,N_14204,N_14766);
nand U15398 (N_15398,N_14317,N_14931);
and U15399 (N_15399,N_14924,N_14149);
nor U15400 (N_15400,N_14634,N_14667);
nand U15401 (N_15401,N_14877,N_14856);
and U15402 (N_15402,N_14200,N_14919);
xnor U15403 (N_15403,N_14669,N_14912);
nand U15404 (N_15404,N_14044,N_14972);
nor U15405 (N_15405,N_14303,N_14414);
nor U15406 (N_15406,N_14639,N_14435);
or U15407 (N_15407,N_14045,N_14368);
or U15408 (N_15408,N_14450,N_14471);
and U15409 (N_15409,N_14683,N_14775);
nand U15410 (N_15410,N_14007,N_14237);
nand U15411 (N_15411,N_14589,N_14426);
xnor U15412 (N_15412,N_14113,N_14031);
nand U15413 (N_15413,N_14126,N_14230);
nor U15414 (N_15414,N_14215,N_14383);
and U15415 (N_15415,N_14111,N_14723);
xor U15416 (N_15416,N_14796,N_14427);
xnor U15417 (N_15417,N_14062,N_14751);
or U15418 (N_15418,N_14481,N_14193);
nand U15419 (N_15419,N_14555,N_14132);
nand U15420 (N_15420,N_14675,N_14466);
nand U15421 (N_15421,N_14834,N_14225);
xor U15422 (N_15422,N_14623,N_14805);
and U15423 (N_15423,N_14562,N_14956);
or U15424 (N_15424,N_14320,N_14889);
nand U15425 (N_15425,N_14665,N_14180);
or U15426 (N_15426,N_14815,N_14208);
xnor U15427 (N_15427,N_14184,N_14903);
and U15428 (N_15428,N_14582,N_14395);
nor U15429 (N_15429,N_14542,N_14833);
or U15430 (N_15430,N_14822,N_14506);
nor U15431 (N_15431,N_14432,N_14748);
nand U15432 (N_15432,N_14181,N_14930);
xor U15433 (N_15433,N_14685,N_14340);
xnor U15434 (N_15434,N_14108,N_14491);
or U15435 (N_15435,N_14774,N_14259);
and U15436 (N_15436,N_14955,N_14724);
and U15437 (N_15437,N_14300,N_14969);
nor U15438 (N_15438,N_14043,N_14371);
xnor U15439 (N_15439,N_14464,N_14356);
and U15440 (N_15440,N_14740,N_14861);
nand U15441 (N_15441,N_14106,N_14900);
xnor U15442 (N_15442,N_14967,N_14902);
nand U15443 (N_15443,N_14377,N_14406);
xnor U15444 (N_15444,N_14086,N_14544);
xor U15445 (N_15445,N_14518,N_14783);
or U15446 (N_15446,N_14576,N_14593);
or U15447 (N_15447,N_14788,N_14677);
or U15448 (N_15448,N_14915,N_14517);
and U15449 (N_15449,N_14586,N_14529);
or U15450 (N_15450,N_14463,N_14948);
nor U15451 (N_15451,N_14616,N_14255);
nand U15452 (N_15452,N_14803,N_14823);
nand U15453 (N_15453,N_14884,N_14333);
nor U15454 (N_15454,N_14790,N_14354);
xnor U15455 (N_15455,N_14864,N_14351);
xor U15456 (N_15456,N_14000,N_14585);
or U15457 (N_15457,N_14550,N_14513);
xor U15458 (N_15458,N_14688,N_14256);
nor U15459 (N_15459,N_14737,N_14037);
and U15460 (N_15460,N_14526,N_14816);
xnor U15461 (N_15461,N_14527,N_14381);
nor U15462 (N_15462,N_14624,N_14153);
and U15463 (N_15463,N_14068,N_14006);
nand U15464 (N_15464,N_14505,N_14917);
or U15465 (N_15465,N_14497,N_14020);
or U15466 (N_15466,N_14992,N_14890);
nand U15467 (N_15467,N_14005,N_14686);
and U15468 (N_15468,N_14211,N_14175);
and U15469 (N_15469,N_14825,N_14339);
nand U15470 (N_15470,N_14763,N_14728);
and U15471 (N_15471,N_14560,N_14264);
nand U15472 (N_15472,N_14078,N_14901);
nor U15473 (N_15473,N_14369,N_14155);
or U15474 (N_15474,N_14871,N_14851);
and U15475 (N_15475,N_14376,N_14473);
nand U15476 (N_15476,N_14084,N_14859);
nor U15477 (N_15477,N_14151,N_14033);
nand U15478 (N_15478,N_14979,N_14090);
nand U15479 (N_15479,N_14600,N_14292);
and U15480 (N_15480,N_14836,N_14905);
nand U15481 (N_15481,N_14195,N_14064);
nor U15482 (N_15482,N_14447,N_14492);
xor U15483 (N_15483,N_14455,N_14315);
nand U15484 (N_15484,N_14606,N_14494);
nand U15485 (N_15485,N_14875,N_14189);
nor U15486 (N_15486,N_14909,N_14811);
or U15487 (N_15487,N_14398,N_14999);
nand U15488 (N_15488,N_14762,N_14283);
or U15489 (N_15489,N_14791,N_14662);
nand U15490 (N_15490,N_14094,N_14646);
xnor U15491 (N_15491,N_14325,N_14281);
nand U15492 (N_15492,N_14088,N_14574);
and U15493 (N_15493,N_14101,N_14733);
nand U15494 (N_15494,N_14496,N_14913);
nand U15495 (N_15495,N_14660,N_14229);
nand U15496 (N_15496,N_14604,N_14107);
or U15497 (N_15497,N_14765,N_14430);
xnor U15498 (N_15498,N_14402,N_14648);
or U15499 (N_15499,N_14360,N_14906);
nand U15500 (N_15500,N_14937,N_14734);
or U15501 (N_15501,N_14695,N_14758);
nor U15502 (N_15502,N_14000,N_14874);
or U15503 (N_15503,N_14904,N_14177);
nand U15504 (N_15504,N_14123,N_14628);
xnor U15505 (N_15505,N_14152,N_14040);
and U15506 (N_15506,N_14003,N_14318);
or U15507 (N_15507,N_14196,N_14279);
xnor U15508 (N_15508,N_14366,N_14621);
and U15509 (N_15509,N_14256,N_14916);
nor U15510 (N_15510,N_14202,N_14918);
and U15511 (N_15511,N_14344,N_14017);
xor U15512 (N_15512,N_14560,N_14887);
nor U15513 (N_15513,N_14061,N_14101);
and U15514 (N_15514,N_14427,N_14139);
nand U15515 (N_15515,N_14870,N_14484);
or U15516 (N_15516,N_14309,N_14643);
or U15517 (N_15517,N_14240,N_14487);
xnor U15518 (N_15518,N_14984,N_14480);
nand U15519 (N_15519,N_14521,N_14990);
xor U15520 (N_15520,N_14488,N_14498);
xnor U15521 (N_15521,N_14382,N_14976);
nor U15522 (N_15522,N_14131,N_14488);
nor U15523 (N_15523,N_14086,N_14024);
xor U15524 (N_15524,N_14717,N_14184);
nand U15525 (N_15525,N_14866,N_14956);
and U15526 (N_15526,N_14070,N_14508);
and U15527 (N_15527,N_14676,N_14161);
and U15528 (N_15528,N_14910,N_14182);
nor U15529 (N_15529,N_14505,N_14466);
xnor U15530 (N_15530,N_14859,N_14770);
nor U15531 (N_15531,N_14543,N_14414);
nand U15532 (N_15532,N_14853,N_14193);
nand U15533 (N_15533,N_14902,N_14325);
nor U15534 (N_15534,N_14218,N_14766);
xnor U15535 (N_15535,N_14605,N_14427);
xor U15536 (N_15536,N_14417,N_14393);
xnor U15537 (N_15537,N_14098,N_14677);
nor U15538 (N_15538,N_14472,N_14495);
nor U15539 (N_15539,N_14822,N_14929);
xnor U15540 (N_15540,N_14352,N_14360);
nor U15541 (N_15541,N_14837,N_14972);
or U15542 (N_15542,N_14204,N_14337);
nor U15543 (N_15543,N_14023,N_14751);
and U15544 (N_15544,N_14865,N_14911);
and U15545 (N_15545,N_14408,N_14629);
nand U15546 (N_15546,N_14000,N_14781);
nand U15547 (N_15547,N_14753,N_14057);
xnor U15548 (N_15548,N_14602,N_14744);
nand U15549 (N_15549,N_14060,N_14656);
or U15550 (N_15550,N_14191,N_14129);
or U15551 (N_15551,N_14157,N_14384);
xnor U15552 (N_15552,N_14883,N_14381);
xnor U15553 (N_15553,N_14967,N_14783);
and U15554 (N_15554,N_14405,N_14139);
xor U15555 (N_15555,N_14233,N_14143);
xor U15556 (N_15556,N_14461,N_14959);
or U15557 (N_15557,N_14775,N_14187);
and U15558 (N_15558,N_14095,N_14509);
nand U15559 (N_15559,N_14808,N_14843);
or U15560 (N_15560,N_14522,N_14731);
or U15561 (N_15561,N_14047,N_14630);
nand U15562 (N_15562,N_14971,N_14694);
nand U15563 (N_15563,N_14144,N_14488);
nand U15564 (N_15564,N_14933,N_14440);
or U15565 (N_15565,N_14932,N_14608);
nor U15566 (N_15566,N_14829,N_14341);
nand U15567 (N_15567,N_14658,N_14654);
nand U15568 (N_15568,N_14521,N_14503);
or U15569 (N_15569,N_14187,N_14085);
and U15570 (N_15570,N_14725,N_14490);
and U15571 (N_15571,N_14295,N_14736);
nand U15572 (N_15572,N_14535,N_14476);
or U15573 (N_15573,N_14297,N_14794);
nor U15574 (N_15574,N_14911,N_14555);
or U15575 (N_15575,N_14456,N_14314);
xnor U15576 (N_15576,N_14922,N_14793);
nand U15577 (N_15577,N_14499,N_14743);
and U15578 (N_15578,N_14061,N_14605);
xnor U15579 (N_15579,N_14043,N_14784);
nand U15580 (N_15580,N_14491,N_14407);
nor U15581 (N_15581,N_14586,N_14725);
nor U15582 (N_15582,N_14535,N_14377);
nand U15583 (N_15583,N_14492,N_14389);
xor U15584 (N_15584,N_14234,N_14727);
nor U15585 (N_15585,N_14277,N_14420);
and U15586 (N_15586,N_14649,N_14400);
and U15587 (N_15587,N_14039,N_14849);
xor U15588 (N_15588,N_14138,N_14323);
nor U15589 (N_15589,N_14420,N_14287);
and U15590 (N_15590,N_14075,N_14785);
and U15591 (N_15591,N_14035,N_14677);
or U15592 (N_15592,N_14816,N_14650);
nor U15593 (N_15593,N_14666,N_14439);
nor U15594 (N_15594,N_14350,N_14957);
or U15595 (N_15595,N_14068,N_14109);
nor U15596 (N_15596,N_14268,N_14064);
nand U15597 (N_15597,N_14816,N_14287);
xor U15598 (N_15598,N_14164,N_14618);
nor U15599 (N_15599,N_14236,N_14910);
and U15600 (N_15600,N_14602,N_14331);
and U15601 (N_15601,N_14912,N_14421);
xnor U15602 (N_15602,N_14190,N_14578);
nand U15603 (N_15603,N_14933,N_14416);
nand U15604 (N_15604,N_14109,N_14030);
nor U15605 (N_15605,N_14830,N_14992);
or U15606 (N_15606,N_14118,N_14202);
xnor U15607 (N_15607,N_14790,N_14799);
nor U15608 (N_15608,N_14153,N_14500);
nand U15609 (N_15609,N_14990,N_14489);
nand U15610 (N_15610,N_14684,N_14620);
nor U15611 (N_15611,N_14153,N_14130);
xnor U15612 (N_15612,N_14201,N_14784);
or U15613 (N_15613,N_14225,N_14621);
nor U15614 (N_15614,N_14188,N_14139);
nor U15615 (N_15615,N_14560,N_14685);
and U15616 (N_15616,N_14197,N_14140);
xnor U15617 (N_15617,N_14829,N_14042);
nand U15618 (N_15618,N_14447,N_14378);
nor U15619 (N_15619,N_14982,N_14901);
nand U15620 (N_15620,N_14532,N_14202);
and U15621 (N_15621,N_14586,N_14942);
nor U15622 (N_15622,N_14355,N_14079);
xnor U15623 (N_15623,N_14234,N_14768);
and U15624 (N_15624,N_14363,N_14042);
nand U15625 (N_15625,N_14609,N_14880);
or U15626 (N_15626,N_14584,N_14163);
nand U15627 (N_15627,N_14319,N_14490);
or U15628 (N_15628,N_14166,N_14313);
xnor U15629 (N_15629,N_14167,N_14390);
and U15630 (N_15630,N_14800,N_14934);
nand U15631 (N_15631,N_14249,N_14036);
nor U15632 (N_15632,N_14197,N_14967);
nand U15633 (N_15633,N_14853,N_14216);
nor U15634 (N_15634,N_14706,N_14828);
and U15635 (N_15635,N_14527,N_14442);
xor U15636 (N_15636,N_14202,N_14841);
nor U15637 (N_15637,N_14361,N_14482);
and U15638 (N_15638,N_14635,N_14859);
nand U15639 (N_15639,N_14005,N_14347);
nor U15640 (N_15640,N_14770,N_14554);
or U15641 (N_15641,N_14267,N_14653);
xnor U15642 (N_15642,N_14142,N_14185);
xor U15643 (N_15643,N_14106,N_14639);
xnor U15644 (N_15644,N_14536,N_14499);
and U15645 (N_15645,N_14905,N_14773);
or U15646 (N_15646,N_14432,N_14774);
xnor U15647 (N_15647,N_14432,N_14393);
and U15648 (N_15648,N_14892,N_14633);
nand U15649 (N_15649,N_14754,N_14292);
nor U15650 (N_15650,N_14020,N_14108);
nand U15651 (N_15651,N_14330,N_14834);
nand U15652 (N_15652,N_14992,N_14775);
and U15653 (N_15653,N_14822,N_14791);
nor U15654 (N_15654,N_14647,N_14448);
xor U15655 (N_15655,N_14593,N_14309);
and U15656 (N_15656,N_14087,N_14226);
or U15657 (N_15657,N_14688,N_14450);
nand U15658 (N_15658,N_14874,N_14569);
and U15659 (N_15659,N_14288,N_14964);
or U15660 (N_15660,N_14619,N_14214);
xnor U15661 (N_15661,N_14248,N_14946);
nor U15662 (N_15662,N_14022,N_14414);
xor U15663 (N_15663,N_14116,N_14231);
nor U15664 (N_15664,N_14321,N_14005);
or U15665 (N_15665,N_14306,N_14166);
or U15666 (N_15666,N_14921,N_14485);
xor U15667 (N_15667,N_14027,N_14383);
xnor U15668 (N_15668,N_14583,N_14828);
nand U15669 (N_15669,N_14468,N_14657);
nand U15670 (N_15670,N_14344,N_14011);
xor U15671 (N_15671,N_14374,N_14982);
and U15672 (N_15672,N_14357,N_14102);
xor U15673 (N_15673,N_14542,N_14565);
nor U15674 (N_15674,N_14304,N_14742);
xor U15675 (N_15675,N_14860,N_14798);
and U15676 (N_15676,N_14108,N_14570);
nor U15677 (N_15677,N_14682,N_14748);
xnor U15678 (N_15678,N_14528,N_14670);
and U15679 (N_15679,N_14652,N_14584);
nor U15680 (N_15680,N_14723,N_14214);
xnor U15681 (N_15681,N_14608,N_14966);
xnor U15682 (N_15682,N_14269,N_14258);
and U15683 (N_15683,N_14581,N_14754);
and U15684 (N_15684,N_14850,N_14765);
nand U15685 (N_15685,N_14375,N_14188);
nor U15686 (N_15686,N_14335,N_14664);
and U15687 (N_15687,N_14574,N_14922);
nand U15688 (N_15688,N_14845,N_14059);
xnor U15689 (N_15689,N_14751,N_14493);
and U15690 (N_15690,N_14757,N_14463);
xor U15691 (N_15691,N_14150,N_14009);
nand U15692 (N_15692,N_14004,N_14398);
nand U15693 (N_15693,N_14672,N_14115);
xor U15694 (N_15694,N_14209,N_14168);
or U15695 (N_15695,N_14288,N_14719);
xor U15696 (N_15696,N_14040,N_14732);
or U15697 (N_15697,N_14502,N_14217);
and U15698 (N_15698,N_14583,N_14319);
xnor U15699 (N_15699,N_14551,N_14605);
or U15700 (N_15700,N_14821,N_14394);
and U15701 (N_15701,N_14281,N_14191);
nor U15702 (N_15702,N_14715,N_14287);
or U15703 (N_15703,N_14146,N_14361);
xnor U15704 (N_15704,N_14352,N_14060);
or U15705 (N_15705,N_14296,N_14432);
nor U15706 (N_15706,N_14090,N_14390);
nor U15707 (N_15707,N_14015,N_14658);
xnor U15708 (N_15708,N_14629,N_14164);
xnor U15709 (N_15709,N_14498,N_14575);
nand U15710 (N_15710,N_14114,N_14003);
nor U15711 (N_15711,N_14875,N_14922);
xor U15712 (N_15712,N_14849,N_14169);
xnor U15713 (N_15713,N_14619,N_14784);
and U15714 (N_15714,N_14882,N_14553);
or U15715 (N_15715,N_14411,N_14349);
xnor U15716 (N_15716,N_14820,N_14921);
or U15717 (N_15717,N_14189,N_14428);
xnor U15718 (N_15718,N_14921,N_14930);
and U15719 (N_15719,N_14950,N_14170);
nand U15720 (N_15720,N_14159,N_14265);
nand U15721 (N_15721,N_14958,N_14582);
or U15722 (N_15722,N_14030,N_14648);
nand U15723 (N_15723,N_14605,N_14556);
or U15724 (N_15724,N_14446,N_14289);
and U15725 (N_15725,N_14513,N_14922);
nand U15726 (N_15726,N_14373,N_14634);
and U15727 (N_15727,N_14494,N_14235);
and U15728 (N_15728,N_14224,N_14206);
and U15729 (N_15729,N_14260,N_14110);
nand U15730 (N_15730,N_14806,N_14703);
nor U15731 (N_15731,N_14342,N_14789);
xor U15732 (N_15732,N_14734,N_14707);
xor U15733 (N_15733,N_14556,N_14249);
nand U15734 (N_15734,N_14655,N_14580);
or U15735 (N_15735,N_14665,N_14065);
and U15736 (N_15736,N_14311,N_14630);
and U15737 (N_15737,N_14377,N_14046);
xor U15738 (N_15738,N_14681,N_14810);
nor U15739 (N_15739,N_14473,N_14031);
and U15740 (N_15740,N_14646,N_14930);
nor U15741 (N_15741,N_14975,N_14577);
or U15742 (N_15742,N_14792,N_14363);
and U15743 (N_15743,N_14451,N_14265);
or U15744 (N_15744,N_14385,N_14734);
nor U15745 (N_15745,N_14482,N_14331);
or U15746 (N_15746,N_14006,N_14230);
nand U15747 (N_15747,N_14104,N_14732);
nor U15748 (N_15748,N_14919,N_14803);
nand U15749 (N_15749,N_14933,N_14712);
or U15750 (N_15750,N_14604,N_14638);
xnor U15751 (N_15751,N_14853,N_14642);
and U15752 (N_15752,N_14062,N_14012);
and U15753 (N_15753,N_14126,N_14619);
xnor U15754 (N_15754,N_14628,N_14314);
or U15755 (N_15755,N_14784,N_14973);
nand U15756 (N_15756,N_14770,N_14378);
nand U15757 (N_15757,N_14374,N_14037);
nand U15758 (N_15758,N_14965,N_14408);
xnor U15759 (N_15759,N_14614,N_14885);
and U15760 (N_15760,N_14911,N_14183);
xor U15761 (N_15761,N_14529,N_14662);
or U15762 (N_15762,N_14391,N_14712);
nor U15763 (N_15763,N_14911,N_14790);
nor U15764 (N_15764,N_14756,N_14879);
nor U15765 (N_15765,N_14251,N_14796);
nand U15766 (N_15766,N_14624,N_14572);
or U15767 (N_15767,N_14605,N_14941);
nand U15768 (N_15768,N_14579,N_14463);
xnor U15769 (N_15769,N_14394,N_14795);
and U15770 (N_15770,N_14454,N_14396);
or U15771 (N_15771,N_14186,N_14926);
nand U15772 (N_15772,N_14643,N_14920);
nand U15773 (N_15773,N_14407,N_14144);
xor U15774 (N_15774,N_14050,N_14600);
xor U15775 (N_15775,N_14881,N_14735);
nand U15776 (N_15776,N_14356,N_14008);
xnor U15777 (N_15777,N_14374,N_14205);
and U15778 (N_15778,N_14887,N_14450);
or U15779 (N_15779,N_14398,N_14986);
nand U15780 (N_15780,N_14207,N_14673);
nor U15781 (N_15781,N_14451,N_14287);
xor U15782 (N_15782,N_14491,N_14038);
nand U15783 (N_15783,N_14430,N_14112);
xnor U15784 (N_15784,N_14571,N_14352);
xor U15785 (N_15785,N_14708,N_14837);
nand U15786 (N_15786,N_14858,N_14546);
nor U15787 (N_15787,N_14644,N_14446);
or U15788 (N_15788,N_14447,N_14075);
or U15789 (N_15789,N_14229,N_14313);
nor U15790 (N_15790,N_14525,N_14764);
xnor U15791 (N_15791,N_14265,N_14604);
xor U15792 (N_15792,N_14494,N_14579);
nand U15793 (N_15793,N_14608,N_14586);
nand U15794 (N_15794,N_14901,N_14872);
nor U15795 (N_15795,N_14625,N_14987);
and U15796 (N_15796,N_14618,N_14028);
and U15797 (N_15797,N_14627,N_14292);
nor U15798 (N_15798,N_14834,N_14510);
nor U15799 (N_15799,N_14009,N_14494);
xor U15800 (N_15800,N_14299,N_14082);
nand U15801 (N_15801,N_14031,N_14372);
or U15802 (N_15802,N_14130,N_14971);
nand U15803 (N_15803,N_14118,N_14650);
and U15804 (N_15804,N_14404,N_14640);
or U15805 (N_15805,N_14620,N_14147);
nor U15806 (N_15806,N_14805,N_14924);
nand U15807 (N_15807,N_14007,N_14348);
or U15808 (N_15808,N_14062,N_14625);
xor U15809 (N_15809,N_14546,N_14335);
and U15810 (N_15810,N_14346,N_14992);
xor U15811 (N_15811,N_14418,N_14105);
nand U15812 (N_15812,N_14037,N_14415);
nand U15813 (N_15813,N_14917,N_14688);
or U15814 (N_15814,N_14530,N_14636);
and U15815 (N_15815,N_14691,N_14187);
and U15816 (N_15816,N_14856,N_14819);
nand U15817 (N_15817,N_14149,N_14685);
xnor U15818 (N_15818,N_14052,N_14059);
nor U15819 (N_15819,N_14640,N_14295);
nor U15820 (N_15820,N_14592,N_14893);
and U15821 (N_15821,N_14460,N_14800);
and U15822 (N_15822,N_14051,N_14272);
xnor U15823 (N_15823,N_14327,N_14519);
xnor U15824 (N_15824,N_14069,N_14496);
nor U15825 (N_15825,N_14133,N_14967);
xnor U15826 (N_15826,N_14269,N_14327);
nor U15827 (N_15827,N_14502,N_14254);
xor U15828 (N_15828,N_14900,N_14514);
nand U15829 (N_15829,N_14501,N_14213);
nand U15830 (N_15830,N_14981,N_14116);
nor U15831 (N_15831,N_14665,N_14727);
or U15832 (N_15832,N_14811,N_14369);
or U15833 (N_15833,N_14674,N_14244);
xnor U15834 (N_15834,N_14563,N_14578);
or U15835 (N_15835,N_14098,N_14785);
nand U15836 (N_15836,N_14781,N_14766);
nand U15837 (N_15837,N_14963,N_14822);
nor U15838 (N_15838,N_14787,N_14190);
nand U15839 (N_15839,N_14178,N_14833);
nor U15840 (N_15840,N_14131,N_14584);
nor U15841 (N_15841,N_14802,N_14526);
and U15842 (N_15842,N_14846,N_14894);
nor U15843 (N_15843,N_14817,N_14140);
xor U15844 (N_15844,N_14640,N_14926);
xor U15845 (N_15845,N_14201,N_14083);
nand U15846 (N_15846,N_14041,N_14602);
nor U15847 (N_15847,N_14679,N_14993);
nand U15848 (N_15848,N_14113,N_14073);
nor U15849 (N_15849,N_14275,N_14414);
nor U15850 (N_15850,N_14510,N_14514);
nand U15851 (N_15851,N_14570,N_14587);
and U15852 (N_15852,N_14611,N_14840);
nor U15853 (N_15853,N_14939,N_14752);
nor U15854 (N_15854,N_14347,N_14354);
or U15855 (N_15855,N_14370,N_14177);
nor U15856 (N_15856,N_14490,N_14177);
xnor U15857 (N_15857,N_14473,N_14318);
and U15858 (N_15858,N_14823,N_14699);
or U15859 (N_15859,N_14983,N_14857);
or U15860 (N_15860,N_14900,N_14052);
nor U15861 (N_15861,N_14290,N_14358);
nor U15862 (N_15862,N_14896,N_14877);
and U15863 (N_15863,N_14592,N_14484);
xnor U15864 (N_15864,N_14885,N_14244);
nor U15865 (N_15865,N_14756,N_14402);
and U15866 (N_15866,N_14833,N_14831);
nand U15867 (N_15867,N_14531,N_14758);
and U15868 (N_15868,N_14114,N_14348);
and U15869 (N_15869,N_14925,N_14295);
nor U15870 (N_15870,N_14572,N_14702);
xor U15871 (N_15871,N_14290,N_14568);
or U15872 (N_15872,N_14542,N_14769);
xnor U15873 (N_15873,N_14132,N_14676);
xnor U15874 (N_15874,N_14754,N_14518);
or U15875 (N_15875,N_14272,N_14702);
nand U15876 (N_15876,N_14755,N_14113);
nand U15877 (N_15877,N_14074,N_14134);
xnor U15878 (N_15878,N_14803,N_14665);
xor U15879 (N_15879,N_14715,N_14741);
nand U15880 (N_15880,N_14358,N_14023);
nand U15881 (N_15881,N_14276,N_14070);
or U15882 (N_15882,N_14975,N_14906);
nor U15883 (N_15883,N_14156,N_14325);
nor U15884 (N_15884,N_14536,N_14528);
and U15885 (N_15885,N_14313,N_14388);
nand U15886 (N_15886,N_14828,N_14399);
nor U15887 (N_15887,N_14956,N_14772);
or U15888 (N_15888,N_14579,N_14681);
xnor U15889 (N_15889,N_14785,N_14676);
or U15890 (N_15890,N_14936,N_14545);
and U15891 (N_15891,N_14829,N_14588);
nand U15892 (N_15892,N_14660,N_14245);
nor U15893 (N_15893,N_14308,N_14394);
and U15894 (N_15894,N_14099,N_14082);
nor U15895 (N_15895,N_14244,N_14246);
and U15896 (N_15896,N_14297,N_14367);
and U15897 (N_15897,N_14055,N_14850);
and U15898 (N_15898,N_14073,N_14456);
nor U15899 (N_15899,N_14245,N_14397);
and U15900 (N_15900,N_14666,N_14160);
nand U15901 (N_15901,N_14735,N_14985);
nor U15902 (N_15902,N_14709,N_14938);
nor U15903 (N_15903,N_14469,N_14204);
or U15904 (N_15904,N_14912,N_14816);
xnor U15905 (N_15905,N_14006,N_14902);
and U15906 (N_15906,N_14463,N_14784);
xor U15907 (N_15907,N_14056,N_14733);
nor U15908 (N_15908,N_14861,N_14482);
xnor U15909 (N_15909,N_14190,N_14847);
and U15910 (N_15910,N_14706,N_14716);
nand U15911 (N_15911,N_14370,N_14674);
xnor U15912 (N_15912,N_14548,N_14290);
nand U15913 (N_15913,N_14249,N_14030);
xor U15914 (N_15914,N_14550,N_14997);
nor U15915 (N_15915,N_14119,N_14720);
xnor U15916 (N_15916,N_14996,N_14569);
nor U15917 (N_15917,N_14853,N_14584);
xnor U15918 (N_15918,N_14170,N_14528);
or U15919 (N_15919,N_14917,N_14333);
or U15920 (N_15920,N_14861,N_14637);
and U15921 (N_15921,N_14218,N_14602);
and U15922 (N_15922,N_14128,N_14398);
or U15923 (N_15923,N_14252,N_14374);
and U15924 (N_15924,N_14942,N_14750);
and U15925 (N_15925,N_14404,N_14311);
nand U15926 (N_15926,N_14613,N_14043);
nor U15927 (N_15927,N_14696,N_14066);
nor U15928 (N_15928,N_14716,N_14512);
xor U15929 (N_15929,N_14441,N_14426);
nand U15930 (N_15930,N_14303,N_14775);
nor U15931 (N_15931,N_14870,N_14027);
and U15932 (N_15932,N_14375,N_14836);
or U15933 (N_15933,N_14632,N_14600);
nand U15934 (N_15934,N_14522,N_14940);
xor U15935 (N_15935,N_14490,N_14738);
or U15936 (N_15936,N_14452,N_14881);
and U15937 (N_15937,N_14893,N_14616);
nand U15938 (N_15938,N_14672,N_14844);
xnor U15939 (N_15939,N_14696,N_14261);
or U15940 (N_15940,N_14628,N_14438);
nand U15941 (N_15941,N_14851,N_14312);
and U15942 (N_15942,N_14263,N_14422);
or U15943 (N_15943,N_14680,N_14852);
and U15944 (N_15944,N_14306,N_14499);
or U15945 (N_15945,N_14674,N_14548);
nand U15946 (N_15946,N_14447,N_14340);
nor U15947 (N_15947,N_14652,N_14841);
nor U15948 (N_15948,N_14148,N_14471);
xnor U15949 (N_15949,N_14233,N_14596);
nand U15950 (N_15950,N_14835,N_14404);
xnor U15951 (N_15951,N_14855,N_14302);
nor U15952 (N_15952,N_14163,N_14129);
nand U15953 (N_15953,N_14643,N_14045);
and U15954 (N_15954,N_14948,N_14353);
nand U15955 (N_15955,N_14738,N_14335);
and U15956 (N_15956,N_14214,N_14291);
and U15957 (N_15957,N_14598,N_14899);
xor U15958 (N_15958,N_14592,N_14300);
and U15959 (N_15959,N_14341,N_14461);
and U15960 (N_15960,N_14929,N_14302);
and U15961 (N_15961,N_14403,N_14003);
nand U15962 (N_15962,N_14358,N_14415);
nand U15963 (N_15963,N_14290,N_14124);
nand U15964 (N_15964,N_14065,N_14042);
xor U15965 (N_15965,N_14243,N_14526);
nand U15966 (N_15966,N_14784,N_14857);
or U15967 (N_15967,N_14276,N_14798);
xnor U15968 (N_15968,N_14304,N_14403);
xor U15969 (N_15969,N_14666,N_14961);
and U15970 (N_15970,N_14979,N_14448);
and U15971 (N_15971,N_14457,N_14463);
and U15972 (N_15972,N_14195,N_14053);
nand U15973 (N_15973,N_14229,N_14355);
nand U15974 (N_15974,N_14679,N_14251);
nand U15975 (N_15975,N_14073,N_14704);
and U15976 (N_15976,N_14463,N_14199);
or U15977 (N_15977,N_14152,N_14227);
and U15978 (N_15978,N_14722,N_14626);
nand U15979 (N_15979,N_14598,N_14933);
nand U15980 (N_15980,N_14862,N_14732);
and U15981 (N_15981,N_14245,N_14357);
or U15982 (N_15982,N_14995,N_14059);
or U15983 (N_15983,N_14259,N_14106);
nand U15984 (N_15984,N_14316,N_14073);
and U15985 (N_15985,N_14531,N_14551);
nand U15986 (N_15986,N_14052,N_14833);
and U15987 (N_15987,N_14551,N_14371);
nand U15988 (N_15988,N_14680,N_14901);
nand U15989 (N_15989,N_14994,N_14901);
nor U15990 (N_15990,N_14321,N_14102);
xor U15991 (N_15991,N_14767,N_14861);
and U15992 (N_15992,N_14633,N_14333);
xnor U15993 (N_15993,N_14816,N_14969);
nor U15994 (N_15994,N_14553,N_14757);
nand U15995 (N_15995,N_14223,N_14900);
xnor U15996 (N_15996,N_14063,N_14622);
nand U15997 (N_15997,N_14714,N_14662);
xnor U15998 (N_15998,N_14237,N_14717);
or U15999 (N_15999,N_14764,N_14372);
nor U16000 (N_16000,N_15234,N_15887);
nand U16001 (N_16001,N_15121,N_15308);
or U16002 (N_16002,N_15881,N_15662);
xnor U16003 (N_16003,N_15224,N_15686);
nor U16004 (N_16004,N_15975,N_15115);
or U16005 (N_16005,N_15884,N_15671);
xor U16006 (N_16006,N_15725,N_15506);
xor U16007 (N_16007,N_15715,N_15325);
xor U16008 (N_16008,N_15533,N_15741);
or U16009 (N_16009,N_15582,N_15519);
and U16010 (N_16010,N_15163,N_15626);
nor U16011 (N_16011,N_15013,N_15299);
nor U16012 (N_16012,N_15432,N_15988);
nand U16013 (N_16013,N_15553,N_15610);
and U16014 (N_16014,N_15555,N_15266);
nand U16015 (N_16015,N_15260,N_15226);
and U16016 (N_16016,N_15052,N_15390);
nand U16017 (N_16017,N_15602,N_15098);
xor U16018 (N_16018,N_15225,N_15682);
or U16019 (N_16019,N_15567,N_15197);
nand U16020 (N_16020,N_15433,N_15763);
or U16021 (N_16021,N_15985,N_15687);
and U16022 (N_16022,N_15600,N_15864);
and U16023 (N_16023,N_15191,N_15304);
nor U16024 (N_16024,N_15425,N_15713);
and U16025 (N_16025,N_15323,N_15385);
nand U16026 (N_16026,N_15938,N_15246);
nand U16027 (N_16027,N_15669,N_15300);
nor U16028 (N_16028,N_15535,N_15134);
and U16029 (N_16029,N_15587,N_15783);
nand U16030 (N_16030,N_15484,N_15603);
xor U16031 (N_16031,N_15078,N_15059);
xor U16032 (N_16032,N_15905,N_15672);
nand U16033 (N_16033,N_15086,N_15024);
xnor U16034 (N_16034,N_15062,N_15638);
nor U16035 (N_16035,N_15696,N_15812);
or U16036 (N_16036,N_15799,N_15992);
xnor U16037 (N_16037,N_15747,N_15824);
and U16038 (N_16038,N_15361,N_15096);
and U16039 (N_16039,N_15190,N_15220);
and U16040 (N_16040,N_15186,N_15819);
nor U16041 (N_16041,N_15601,N_15316);
xnor U16042 (N_16042,N_15693,N_15146);
or U16043 (N_16043,N_15127,N_15100);
nand U16044 (N_16044,N_15818,N_15754);
and U16045 (N_16045,N_15435,N_15635);
and U16046 (N_16046,N_15952,N_15289);
nor U16047 (N_16047,N_15281,N_15064);
nand U16048 (N_16048,N_15558,N_15643);
or U16049 (N_16049,N_15792,N_15674);
xnor U16050 (N_16050,N_15108,N_15159);
and U16051 (N_16051,N_15875,N_15920);
nor U16052 (N_16052,N_15764,N_15423);
and U16053 (N_16053,N_15489,N_15837);
and U16054 (N_16054,N_15835,N_15876);
and U16055 (N_16055,N_15080,N_15073);
xor U16056 (N_16056,N_15481,N_15175);
and U16057 (N_16057,N_15898,N_15907);
nand U16058 (N_16058,N_15228,N_15443);
nand U16059 (N_16059,N_15951,N_15298);
and U16060 (N_16060,N_15156,N_15749);
and U16061 (N_16061,N_15014,N_15598);
or U16062 (N_16062,N_15158,N_15960);
and U16063 (N_16063,N_15499,N_15744);
and U16064 (N_16064,N_15613,N_15734);
or U16065 (N_16065,N_15315,N_15070);
nor U16066 (N_16066,N_15929,N_15294);
xnor U16067 (N_16067,N_15384,N_15195);
nor U16068 (N_16068,N_15169,N_15502);
nor U16069 (N_16069,N_15660,N_15366);
nand U16070 (N_16070,N_15531,N_15415);
nor U16071 (N_16071,N_15599,N_15871);
and U16072 (N_16072,N_15846,N_15196);
nor U16073 (N_16073,N_15775,N_15591);
xnor U16074 (N_16074,N_15051,N_15509);
nand U16075 (N_16075,N_15751,N_15140);
or U16076 (N_16076,N_15337,N_15117);
nor U16077 (N_16077,N_15869,N_15945);
or U16078 (N_16078,N_15360,N_15546);
nor U16079 (N_16079,N_15351,N_15834);
nand U16080 (N_16080,N_15788,N_15075);
or U16081 (N_16081,N_15795,N_15202);
nor U16082 (N_16082,N_15068,N_15465);
nor U16083 (N_16083,N_15828,N_15577);
xor U16084 (N_16084,N_15194,N_15547);
or U16085 (N_16085,N_15910,N_15394);
xnor U16086 (N_16086,N_15785,N_15437);
nor U16087 (N_16087,N_15615,N_15408);
or U16088 (N_16088,N_15641,N_15072);
xnor U16089 (N_16089,N_15411,N_15549);
or U16090 (N_16090,N_15185,N_15798);
nand U16091 (N_16091,N_15244,N_15673);
nor U16092 (N_16092,N_15991,N_15652);
xor U16093 (N_16093,N_15939,N_15733);
and U16094 (N_16094,N_15885,N_15625);
and U16095 (N_16095,N_15612,N_15439);
or U16096 (N_16096,N_15786,N_15892);
xor U16097 (N_16097,N_15103,N_15369);
xnor U16098 (N_16098,N_15797,N_15681);
or U16099 (N_16099,N_15500,N_15604);
and U16100 (N_16100,N_15926,N_15596);
xnor U16101 (N_16101,N_15130,N_15995);
or U16102 (N_16102,N_15275,N_15557);
nor U16103 (N_16103,N_15243,N_15329);
xor U16104 (N_16104,N_15843,N_15621);
nand U16105 (N_16105,N_15324,N_15262);
and U16106 (N_16106,N_15357,N_15987);
and U16107 (N_16107,N_15911,N_15405);
xor U16108 (N_16108,N_15962,N_15398);
nand U16109 (N_16109,N_15507,N_15208);
and U16110 (N_16110,N_15627,N_15344);
nand U16111 (N_16111,N_15376,N_15964);
xnor U16112 (N_16112,N_15336,N_15999);
or U16113 (N_16113,N_15946,N_15654);
or U16114 (N_16114,N_15565,N_15285);
xnor U16115 (N_16115,N_15313,N_15728);
or U16116 (N_16116,N_15665,N_15503);
nor U16117 (N_16117,N_15750,N_15559);
nor U16118 (N_16118,N_15003,N_15766);
and U16119 (N_16119,N_15033,N_15584);
xnor U16120 (N_16120,N_15517,N_15233);
and U16121 (N_16121,N_15414,N_15594);
nand U16122 (N_16122,N_15343,N_15990);
nand U16123 (N_16123,N_15804,N_15690);
and U16124 (N_16124,N_15542,N_15501);
nor U16125 (N_16125,N_15381,N_15157);
nor U16126 (N_16126,N_15066,N_15396);
and U16127 (N_16127,N_15286,N_15495);
nor U16128 (N_16128,N_15706,N_15753);
and U16129 (N_16129,N_15189,N_15280);
nor U16130 (N_16130,N_15407,N_15755);
and U16131 (N_16131,N_15203,N_15950);
or U16132 (N_16132,N_15365,N_15354);
and U16133 (N_16133,N_15181,N_15133);
xor U16134 (N_16134,N_15044,N_15772);
and U16135 (N_16135,N_15368,N_15522);
nand U16136 (N_16136,N_15406,N_15049);
and U16137 (N_16137,N_15231,N_15145);
and U16138 (N_16138,N_15017,N_15077);
or U16139 (N_16139,N_15434,N_15107);
nor U16140 (N_16140,N_15923,N_15160);
nor U16141 (N_16141,N_15402,N_15504);
or U16142 (N_16142,N_15057,N_15431);
nor U16143 (N_16143,N_15685,N_15109);
nor U16144 (N_16144,N_15401,N_15328);
or U16145 (N_16145,N_15105,N_15055);
xnor U16146 (N_16146,N_15870,N_15832);
xnor U16147 (N_16147,N_15742,N_15271);
or U16148 (N_16148,N_15114,N_15416);
nor U16149 (N_16149,N_15241,N_15449);
nand U16150 (N_16150,N_15878,N_15664);
xor U16151 (N_16151,N_15184,N_15250);
and U16152 (N_16152,N_15642,N_15427);
and U16153 (N_16153,N_15781,N_15460);
nor U16154 (N_16154,N_15239,N_15016);
and U16155 (N_16155,N_15091,N_15063);
nand U16156 (N_16156,N_15321,N_15392);
nand U16157 (N_16157,N_15462,N_15041);
or U16158 (N_16158,N_15815,N_15482);
nand U16159 (N_16159,N_15167,N_15010);
nand U16160 (N_16160,N_15668,N_15757);
xor U16161 (N_16161,N_15071,N_15767);
xor U16162 (N_16162,N_15479,N_15274);
nand U16163 (N_16163,N_15839,N_15378);
or U16164 (N_16164,N_15088,N_15931);
xnor U16165 (N_16165,N_15128,N_15058);
xnor U16166 (N_16166,N_15735,N_15768);
nand U16167 (N_16167,N_15363,N_15796);
nand U16168 (N_16168,N_15386,N_15709);
or U16169 (N_16169,N_15617,N_15729);
xor U16170 (N_16170,N_15453,N_15291);
xnor U16171 (N_16171,N_15035,N_15417);
and U16172 (N_16172,N_15147,N_15464);
xnor U16173 (N_16173,N_15498,N_15698);
and U16174 (N_16174,N_15578,N_15083);
xor U16175 (N_16175,N_15649,N_15833);
and U16176 (N_16176,N_15647,N_15045);
nor U16177 (N_16177,N_15135,N_15817);
nand U16178 (N_16178,N_15912,N_15803);
nand U16179 (N_16179,N_15322,N_15777);
and U16180 (N_16180,N_15341,N_15173);
nand U16181 (N_16181,N_15830,N_15183);
xnor U16182 (N_16182,N_15983,N_15862);
nand U16183 (N_16183,N_15572,N_15571);
or U16184 (N_16184,N_15981,N_15537);
and U16185 (N_16185,N_15890,N_15512);
xnor U16186 (N_16186,N_15927,N_15521);
and U16187 (N_16187,N_15093,N_15886);
xnor U16188 (N_16188,N_15025,N_15844);
nand U16189 (N_16189,N_15277,N_15111);
or U16190 (N_16190,N_15831,N_15721);
nand U16191 (N_16191,N_15182,N_15825);
nand U16192 (N_16192,N_15663,N_15094);
nand U16193 (N_16193,N_15561,N_15305);
nand U16194 (N_16194,N_15099,N_15644);
or U16195 (N_16195,N_15042,N_15544);
or U16196 (N_16196,N_15312,N_15932);
nor U16197 (N_16197,N_15568,N_15165);
nand U16198 (N_16198,N_15659,N_15873);
nor U16199 (N_16199,N_15908,N_15539);
nor U16200 (N_16200,N_15015,N_15467);
nand U16201 (N_16201,N_15614,N_15726);
xor U16202 (N_16202,N_15670,N_15515);
and U16203 (N_16203,N_15554,N_15773);
xnor U16204 (N_16204,N_15667,N_15152);
nand U16205 (N_16205,N_15865,N_15958);
nand U16206 (N_16206,N_15680,N_15252);
nor U16207 (N_16207,N_15588,N_15897);
or U16208 (N_16208,N_15925,N_15556);
nand U16209 (N_16209,N_15004,N_15560);
nor U16210 (N_16210,N_15123,N_15288);
and U16211 (N_16211,N_15762,N_15466);
and U16212 (N_16212,N_15235,N_15845);
or U16213 (N_16213,N_15776,N_15586);
nand U16214 (N_16214,N_15919,N_15653);
and U16215 (N_16215,N_15139,N_15257);
xor U16216 (N_16216,N_15894,N_15155);
nor U16217 (N_16217,N_15278,N_15081);
and U16218 (N_16218,N_15545,N_15311);
nor U16219 (N_16219,N_15880,N_15816);
nor U16220 (N_16220,N_15697,N_15348);
nand U16221 (N_16221,N_15475,N_15223);
or U16222 (N_16222,N_15811,N_15863);
or U16223 (N_16223,N_15924,N_15276);
and U16224 (N_16224,N_15023,N_15616);
nand U16225 (N_16225,N_15028,N_15389);
and U16226 (N_16226,N_15419,N_15860);
and U16227 (N_16227,N_15903,N_15037);
or U16228 (N_16228,N_15956,N_15930);
nor U16229 (N_16229,N_15214,N_15756);
or U16230 (N_16230,N_15205,N_15000);
and U16231 (N_16231,N_15452,N_15760);
and U16232 (N_16232,N_15583,N_15349);
or U16233 (N_16233,N_15372,N_15765);
and U16234 (N_16234,N_15151,N_15144);
nor U16235 (N_16235,N_15790,N_15532);
or U16236 (N_16236,N_15566,N_15352);
and U16237 (N_16237,N_15794,N_15961);
and U16238 (N_16238,N_15529,N_15948);
nor U16239 (N_16239,N_15718,N_15605);
xor U16240 (N_16240,N_15192,N_15856);
nand U16241 (N_16241,N_15122,N_15889);
and U16242 (N_16242,N_15232,N_15441);
nand U16243 (N_16243,N_15330,N_15410);
nor U16244 (N_16244,N_15236,N_15269);
or U16245 (N_16245,N_15284,N_15178);
nand U16246 (N_16246,N_15116,N_15993);
or U16247 (N_16247,N_15267,N_15575);
nor U16248 (N_16248,N_15069,N_15550);
and U16249 (N_16249,N_15179,N_15353);
or U16250 (N_16250,N_15034,N_15711);
nand U16251 (N_16251,N_15978,N_15618);
nand U16252 (N_16252,N_15838,N_15253);
nand U16253 (N_16253,N_15563,N_15740);
nor U16254 (N_16254,N_15371,N_15695);
xnor U16255 (N_16255,N_15082,N_15675);
xor U16256 (N_16256,N_15850,N_15902);
nand U16257 (N_16257,N_15129,N_15046);
and U16258 (N_16258,N_15332,N_15388);
or U16259 (N_16259,N_15119,N_15018);
xor U16260 (N_16260,N_15730,N_15261);
xnor U16261 (N_16261,N_15331,N_15074);
nor U16262 (N_16262,N_15868,N_15085);
and U16263 (N_16263,N_15256,N_15719);
and U16264 (N_16264,N_15678,N_15518);
and U16265 (N_16265,N_15895,N_15769);
or U16266 (N_16266,N_15210,N_15356);
nor U16267 (N_16267,N_15534,N_15774);
or U16268 (N_16268,N_15858,N_15326);
and U16269 (N_16269,N_15562,N_15496);
and U16270 (N_16270,N_15944,N_15030);
nand U16271 (N_16271,N_15691,N_15714);
or U16272 (N_16272,N_15976,N_15597);
or U16273 (N_16273,N_15009,N_15374);
nand U16274 (N_16274,N_15700,N_15891);
or U16275 (N_16275,N_15188,N_15959);
or U16276 (N_16276,N_15972,N_15632);
or U16277 (N_16277,N_15272,N_15318);
and U16278 (N_16278,N_15636,N_15842);
and U16279 (N_16279,N_15126,N_15631);
nand U16280 (N_16280,N_15997,N_15822);
nand U16281 (N_16281,N_15217,N_15808);
nor U16282 (N_16282,N_15297,N_15821);
xor U16283 (N_16283,N_15254,N_15901);
nand U16284 (N_16284,N_15655,N_15784);
or U16285 (N_16285,N_15040,N_15780);
xor U16286 (N_16286,N_15031,N_15989);
xnor U16287 (N_16287,N_15412,N_15514);
nor U16288 (N_16288,N_15132,N_15650);
or U16289 (N_16289,N_15963,N_15393);
nand U16290 (N_16290,N_15180,N_15490);
or U16291 (N_16291,N_15176,N_15986);
or U16292 (N_16292,N_15268,N_15720);
and U16293 (N_16293,N_15350,N_15153);
nor U16294 (N_16294,N_15065,N_15483);
nor U16295 (N_16295,N_15421,N_15806);
nand U16296 (N_16296,N_15826,N_15974);
xnor U16297 (N_16297,N_15849,N_15474);
or U16298 (N_16298,N_15221,N_15943);
xor U16299 (N_16299,N_15888,N_15488);
nor U16300 (N_16300,N_15448,N_15273);
xnor U16301 (N_16301,N_15589,N_15658);
nand U16302 (N_16302,N_15438,N_15476);
and U16303 (N_16303,N_15789,N_15209);
xor U16304 (N_16304,N_15026,N_15251);
xor U16305 (N_16305,N_15552,N_15306);
xnor U16306 (N_16306,N_15307,N_15342);
nand U16307 (N_16307,N_15637,N_15020);
nand U16308 (N_16308,N_15270,N_15731);
xnor U16309 (N_16309,N_15087,N_15279);
and U16310 (N_16310,N_15984,N_15480);
xnor U16311 (N_16311,N_15904,N_15934);
nor U16312 (N_16312,N_15543,N_15827);
or U16313 (N_16313,N_15216,N_15079);
or U16314 (N_16314,N_15712,N_15882);
or U16315 (N_16315,N_15861,N_15229);
or U16316 (N_16316,N_15168,N_15061);
xor U16317 (N_16317,N_15648,N_15101);
xor U16318 (N_16318,N_15630,N_15036);
nor U16319 (N_16319,N_15928,N_15199);
and U16320 (N_16320,N_15526,N_15998);
and U16321 (N_16321,N_15592,N_15782);
nor U16322 (N_16322,N_15362,N_15440);
or U16323 (N_16323,N_15380,N_15634);
xor U16324 (N_16324,N_15006,N_15138);
xor U16325 (N_16325,N_15131,N_15463);
and U16326 (N_16326,N_15201,N_15611);
xor U16327 (N_16327,N_15089,N_15112);
nor U16328 (N_16328,N_15420,N_15444);
nor U16329 (N_16329,N_15541,N_15053);
or U16330 (N_16330,N_15258,N_15980);
nor U16331 (N_16331,N_15092,N_15704);
and U16332 (N_16332,N_15955,N_15487);
or U16333 (N_16333,N_15513,N_15486);
or U16334 (N_16334,N_15745,N_15248);
nor U16335 (N_16335,N_15623,N_15265);
xor U16336 (N_16336,N_15872,N_15346);
and U16337 (N_16337,N_15802,N_15581);
xnor U16338 (N_16338,N_15450,N_15966);
nand U16339 (N_16339,N_15629,N_15564);
xor U16340 (N_16340,N_15056,N_15633);
or U16341 (N_16341,N_15090,N_15174);
xnor U16342 (N_16342,N_15198,N_15739);
or U16343 (N_16343,N_15149,N_15125);
nand U16344 (N_16344,N_15110,N_15358);
or U16345 (N_16345,N_15370,N_15387);
xnor U16346 (N_16346,N_15607,N_15150);
nand U16347 (N_16347,N_15805,N_15900);
or U16348 (N_16348,N_15238,N_15005);
and U16349 (N_16349,N_15048,N_15227);
nor U16350 (N_16350,N_15778,N_15723);
xnor U16351 (N_16351,N_15367,N_15468);
xnor U16352 (N_16352,N_15397,N_15640);
or U16353 (N_16353,N_15338,N_15836);
and U16354 (N_16354,N_15207,N_15177);
xnor U16355 (N_16355,N_15866,N_15829);
xor U16356 (N_16356,N_15508,N_15230);
xnor U16357 (N_16357,N_15317,N_15454);
and U16358 (N_16358,N_15761,N_15877);
and U16359 (N_16359,N_15237,N_15800);
nand U16360 (N_16360,N_15104,N_15124);
and U16361 (N_16361,N_15528,N_15413);
xnor U16362 (N_16362,N_15801,N_15259);
and U16363 (N_16363,N_15717,N_15050);
xor U16364 (N_16364,N_15187,N_15841);
and U16365 (N_16365,N_15937,N_15979);
or U16366 (N_16366,N_15791,N_15255);
and U16367 (N_16367,N_15540,N_15002);
or U16368 (N_16368,N_15922,N_15851);
or U16369 (N_16369,N_15738,N_15573);
xor U16370 (N_16370,N_15579,N_15164);
or U16371 (N_16371,N_15120,N_15580);
xor U16372 (N_16372,N_15935,N_15688);
nor U16373 (N_16373,N_15770,N_15333);
nor U16374 (N_16374,N_15585,N_15684);
xor U16375 (N_16375,N_15524,N_15595);
nand U16376 (N_16376,N_15345,N_15947);
xnor U16377 (N_16377,N_15067,N_15456);
nand U16378 (N_16378,N_15677,N_15970);
nand U16379 (N_16379,N_15879,N_15106);
xor U16380 (N_16380,N_15705,N_15240);
and U16381 (N_16381,N_15022,N_15309);
nor U16382 (N_16382,N_15491,N_15752);
or U16383 (N_16383,N_15222,N_15445);
or U16384 (N_16384,N_15622,N_15787);
xnor U16385 (N_16385,N_15170,N_15969);
nand U16386 (N_16386,N_15218,N_15293);
or U16387 (N_16387,N_15551,N_15651);
nand U16388 (N_16388,N_15359,N_15823);
or U16389 (N_16389,N_15054,N_15097);
xor U16390 (N_16390,N_15472,N_15424);
nor U16391 (N_16391,N_15478,N_15339);
nor U16392 (N_16392,N_15971,N_15458);
nor U16393 (N_16393,N_15692,N_15683);
and U16394 (N_16394,N_15736,N_15936);
nand U16395 (N_16395,N_15166,N_15249);
nand U16396 (N_16396,N_15699,N_15027);
nand U16397 (N_16397,N_15530,N_15859);
xor U16398 (N_16398,N_15290,N_15942);
nand U16399 (N_16399,N_15032,N_15430);
and U16400 (N_16400,N_15143,N_15949);
xor U16401 (N_16401,N_15007,N_15918);
nand U16402 (N_16402,N_15820,N_15377);
or U16403 (N_16403,N_15883,N_15493);
xor U16404 (N_16404,N_15807,N_15608);
or U16405 (N_16405,N_15382,N_15282);
nor U16406 (N_16406,N_15335,N_15505);
nand U16407 (N_16407,N_15447,N_15302);
nand U16408 (N_16408,N_15391,N_15855);
or U16409 (N_16409,N_15793,N_15245);
or U16410 (N_16410,N_15727,N_15840);
xor U16411 (N_16411,N_15494,N_15909);
or U16412 (N_16412,N_15206,N_15355);
nand U16413 (N_16413,N_15403,N_15570);
or U16414 (N_16414,N_15076,N_15060);
or U16415 (N_16415,N_15142,N_15940);
and U16416 (N_16416,N_15301,N_15264);
xnor U16417 (N_16417,N_15899,N_15538);
or U16418 (N_16418,N_15242,N_15676);
xor U16419 (N_16419,N_15646,N_15574);
nor U16420 (N_16420,N_15593,N_15708);
or U16421 (N_16421,N_15485,N_15215);
xor U16422 (N_16422,N_15400,N_15470);
or U16423 (N_16423,N_15536,N_15896);
xnor U16424 (N_16424,N_15283,N_15471);
nor U16425 (N_16425,N_15497,N_15047);
or U16426 (N_16426,N_15263,N_15038);
xnor U16427 (N_16427,N_15019,N_15477);
xnor U16428 (N_16428,N_15347,N_15141);
nand U16429 (N_16429,N_15619,N_15914);
or U16430 (N_16430,N_15809,N_15247);
or U16431 (N_16431,N_15666,N_15212);
xor U16432 (N_16432,N_15941,N_15710);
xnor U16433 (N_16433,N_15996,N_15893);
and U16434 (N_16434,N_15200,N_15933);
or U16435 (N_16435,N_15913,N_15171);
and U16436 (N_16436,N_15161,N_15810);
xor U16437 (N_16437,N_15399,N_15606);
nand U16438 (N_16438,N_15193,N_15701);
and U16439 (N_16439,N_15314,N_15375);
nor U16440 (N_16440,N_15523,N_15982);
xnor U16441 (N_16441,N_15520,N_15915);
nand U16442 (N_16442,N_15814,N_15527);
and U16443 (N_16443,N_15154,N_15748);
xnor U16444 (N_16444,N_15418,N_15848);
xnor U16445 (N_16445,N_15921,N_15813);
and U16446 (N_16446,N_15404,N_15008);
nand U16447 (N_16447,N_15379,N_15296);
xor U16448 (N_16448,N_15473,N_15364);
xor U16449 (N_16449,N_15451,N_15724);
and U16450 (N_16450,N_15694,N_15867);
xor U16451 (N_16451,N_15967,N_15383);
or U16452 (N_16452,N_15422,N_15510);
xnor U16453 (N_16453,N_15426,N_15576);
or U16454 (N_16454,N_15287,N_15994);
and U16455 (N_16455,N_15340,N_15639);
and U16456 (N_16456,N_15771,N_15118);
xor U16457 (N_16457,N_15461,N_15436);
xnor U16458 (N_16458,N_15459,N_15716);
and U16459 (N_16459,N_15511,N_15954);
nor U16460 (N_16460,N_15852,N_15084);
xor U16461 (N_16461,N_15702,N_15303);
or U16462 (N_16462,N_15095,N_15136);
or U16463 (N_16463,N_15525,N_15620);
or U16464 (N_16464,N_15137,N_15039);
or U16465 (N_16465,N_15732,N_15548);
xnor U16466 (N_16466,N_15722,N_15957);
xnor U16467 (N_16467,N_15029,N_15707);
and U16468 (N_16468,N_15211,N_15043);
xor U16469 (N_16469,N_15457,N_15492);
and U16470 (N_16470,N_15737,N_15609);
nor U16471 (N_16471,N_15746,N_15916);
nor U16472 (N_16472,N_15292,N_15428);
and U16473 (N_16473,N_15906,N_15516);
nor U16474 (N_16474,N_15968,N_15689);
nor U16475 (N_16475,N_15429,N_15148);
nand U16476 (N_16476,N_15446,N_15624);
xnor U16477 (N_16477,N_15011,N_15743);
nor U16478 (N_16478,N_15334,N_15012);
or U16479 (N_16479,N_15977,N_15656);
xnor U16480 (N_16480,N_15319,N_15162);
or U16481 (N_16481,N_15442,N_15409);
nor U16482 (N_16482,N_15857,N_15759);
and U16483 (N_16483,N_15590,N_15628);
nor U16484 (N_16484,N_15001,N_15703);
xor U16485 (N_16485,N_15213,N_15953);
xnor U16486 (N_16486,N_15874,N_15854);
nand U16487 (N_16487,N_15219,N_15320);
xnor U16488 (N_16488,N_15973,N_15758);
xnor U16489 (N_16489,N_15204,N_15327);
nor U16490 (N_16490,N_15847,N_15779);
nor U16491 (N_16491,N_15373,N_15102);
nor U16492 (N_16492,N_15569,N_15172);
nor U16493 (N_16493,N_15645,N_15917);
or U16494 (N_16494,N_15853,N_15661);
xor U16495 (N_16495,N_15965,N_15395);
or U16496 (N_16496,N_15657,N_15469);
xor U16497 (N_16497,N_15113,N_15455);
nor U16498 (N_16498,N_15310,N_15679);
nand U16499 (N_16499,N_15295,N_15021);
xnor U16500 (N_16500,N_15774,N_15270);
and U16501 (N_16501,N_15524,N_15276);
and U16502 (N_16502,N_15824,N_15649);
or U16503 (N_16503,N_15973,N_15081);
and U16504 (N_16504,N_15812,N_15860);
and U16505 (N_16505,N_15779,N_15448);
or U16506 (N_16506,N_15559,N_15622);
xor U16507 (N_16507,N_15666,N_15107);
nor U16508 (N_16508,N_15846,N_15966);
nor U16509 (N_16509,N_15707,N_15014);
or U16510 (N_16510,N_15973,N_15731);
nand U16511 (N_16511,N_15238,N_15479);
or U16512 (N_16512,N_15866,N_15303);
and U16513 (N_16513,N_15105,N_15926);
xnor U16514 (N_16514,N_15656,N_15852);
or U16515 (N_16515,N_15395,N_15126);
and U16516 (N_16516,N_15978,N_15066);
or U16517 (N_16517,N_15499,N_15473);
or U16518 (N_16518,N_15203,N_15008);
nor U16519 (N_16519,N_15879,N_15399);
nor U16520 (N_16520,N_15981,N_15393);
xor U16521 (N_16521,N_15807,N_15294);
and U16522 (N_16522,N_15328,N_15914);
nor U16523 (N_16523,N_15697,N_15277);
and U16524 (N_16524,N_15667,N_15873);
or U16525 (N_16525,N_15746,N_15035);
nand U16526 (N_16526,N_15230,N_15174);
or U16527 (N_16527,N_15336,N_15258);
nor U16528 (N_16528,N_15090,N_15294);
or U16529 (N_16529,N_15879,N_15288);
and U16530 (N_16530,N_15617,N_15487);
and U16531 (N_16531,N_15199,N_15331);
nand U16532 (N_16532,N_15630,N_15305);
xor U16533 (N_16533,N_15621,N_15099);
and U16534 (N_16534,N_15652,N_15414);
xor U16535 (N_16535,N_15017,N_15918);
and U16536 (N_16536,N_15828,N_15119);
nand U16537 (N_16537,N_15730,N_15499);
nand U16538 (N_16538,N_15797,N_15066);
xnor U16539 (N_16539,N_15687,N_15617);
or U16540 (N_16540,N_15977,N_15234);
and U16541 (N_16541,N_15337,N_15682);
and U16542 (N_16542,N_15000,N_15889);
or U16543 (N_16543,N_15313,N_15482);
and U16544 (N_16544,N_15283,N_15621);
xnor U16545 (N_16545,N_15362,N_15762);
and U16546 (N_16546,N_15125,N_15856);
nor U16547 (N_16547,N_15879,N_15913);
xnor U16548 (N_16548,N_15064,N_15839);
or U16549 (N_16549,N_15484,N_15211);
xor U16550 (N_16550,N_15403,N_15928);
and U16551 (N_16551,N_15911,N_15269);
xor U16552 (N_16552,N_15943,N_15136);
nor U16553 (N_16553,N_15903,N_15172);
or U16554 (N_16554,N_15273,N_15445);
and U16555 (N_16555,N_15042,N_15732);
xnor U16556 (N_16556,N_15309,N_15684);
xnor U16557 (N_16557,N_15612,N_15300);
or U16558 (N_16558,N_15607,N_15554);
nand U16559 (N_16559,N_15051,N_15224);
nand U16560 (N_16560,N_15999,N_15740);
and U16561 (N_16561,N_15705,N_15951);
nor U16562 (N_16562,N_15680,N_15128);
nand U16563 (N_16563,N_15305,N_15855);
or U16564 (N_16564,N_15305,N_15816);
xor U16565 (N_16565,N_15023,N_15946);
xnor U16566 (N_16566,N_15117,N_15931);
or U16567 (N_16567,N_15357,N_15954);
nand U16568 (N_16568,N_15420,N_15911);
nor U16569 (N_16569,N_15699,N_15278);
nand U16570 (N_16570,N_15549,N_15696);
or U16571 (N_16571,N_15871,N_15529);
nand U16572 (N_16572,N_15844,N_15265);
or U16573 (N_16573,N_15362,N_15693);
nand U16574 (N_16574,N_15785,N_15522);
and U16575 (N_16575,N_15109,N_15198);
xor U16576 (N_16576,N_15411,N_15750);
or U16577 (N_16577,N_15324,N_15655);
and U16578 (N_16578,N_15738,N_15142);
nand U16579 (N_16579,N_15097,N_15721);
nor U16580 (N_16580,N_15189,N_15106);
nor U16581 (N_16581,N_15299,N_15341);
nor U16582 (N_16582,N_15290,N_15860);
nand U16583 (N_16583,N_15642,N_15917);
or U16584 (N_16584,N_15129,N_15970);
xnor U16585 (N_16585,N_15122,N_15654);
nor U16586 (N_16586,N_15594,N_15776);
and U16587 (N_16587,N_15410,N_15241);
nor U16588 (N_16588,N_15892,N_15399);
xor U16589 (N_16589,N_15564,N_15227);
or U16590 (N_16590,N_15650,N_15123);
or U16591 (N_16591,N_15593,N_15108);
or U16592 (N_16592,N_15883,N_15647);
nand U16593 (N_16593,N_15913,N_15850);
or U16594 (N_16594,N_15652,N_15523);
or U16595 (N_16595,N_15607,N_15747);
nand U16596 (N_16596,N_15793,N_15865);
xor U16597 (N_16597,N_15236,N_15695);
and U16598 (N_16598,N_15504,N_15625);
xor U16599 (N_16599,N_15249,N_15974);
and U16600 (N_16600,N_15939,N_15390);
nand U16601 (N_16601,N_15317,N_15776);
and U16602 (N_16602,N_15925,N_15944);
xnor U16603 (N_16603,N_15202,N_15272);
xor U16604 (N_16604,N_15434,N_15774);
or U16605 (N_16605,N_15145,N_15564);
or U16606 (N_16606,N_15414,N_15386);
nand U16607 (N_16607,N_15737,N_15080);
nand U16608 (N_16608,N_15674,N_15960);
xor U16609 (N_16609,N_15863,N_15568);
or U16610 (N_16610,N_15217,N_15730);
xor U16611 (N_16611,N_15498,N_15099);
or U16612 (N_16612,N_15827,N_15023);
nand U16613 (N_16613,N_15070,N_15551);
and U16614 (N_16614,N_15838,N_15452);
nand U16615 (N_16615,N_15959,N_15537);
nor U16616 (N_16616,N_15548,N_15343);
xor U16617 (N_16617,N_15199,N_15560);
and U16618 (N_16618,N_15481,N_15796);
xor U16619 (N_16619,N_15808,N_15260);
nand U16620 (N_16620,N_15586,N_15850);
and U16621 (N_16621,N_15656,N_15500);
and U16622 (N_16622,N_15168,N_15113);
xnor U16623 (N_16623,N_15593,N_15495);
nand U16624 (N_16624,N_15163,N_15467);
nand U16625 (N_16625,N_15547,N_15766);
or U16626 (N_16626,N_15591,N_15913);
nor U16627 (N_16627,N_15244,N_15479);
xor U16628 (N_16628,N_15678,N_15890);
or U16629 (N_16629,N_15546,N_15713);
nand U16630 (N_16630,N_15628,N_15269);
or U16631 (N_16631,N_15695,N_15372);
or U16632 (N_16632,N_15303,N_15506);
nand U16633 (N_16633,N_15607,N_15980);
or U16634 (N_16634,N_15059,N_15565);
nor U16635 (N_16635,N_15602,N_15756);
nand U16636 (N_16636,N_15266,N_15551);
and U16637 (N_16637,N_15515,N_15115);
xnor U16638 (N_16638,N_15714,N_15134);
and U16639 (N_16639,N_15917,N_15060);
nand U16640 (N_16640,N_15955,N_15553);
nor U16641 (N_16641,N_15773,N_15942);
nor U16642 (N_16642,N_15116,N_15284);
nor U16643 (N_16643,N_15061,N_15023);
or U16644 (N_16644,N_15960,N_15945);
nor U16645 (N_16645,N_15645,N_15698);
nand U16646 (N_16646,N_15207,N_15877);
nand U16647 (N_16647,N_15045,N_15105);
or U16648 (N_16648,N_15895,N_15809);
xor U16649 (N_16649,N_15529,N_15962);
nand U16650 (N_16650,N_15078,N_15778);
nor U16651 (N_16651,N_15798,N_15093);
nand U16652 (N_16652,N_15694,N_15726);
xnor U16653 (N_16653,N_15316,N_15509);
nor U16654 (N_16654,N_15585,N_15073);
nand U16655 (N_16655,N_15368,N_15013);
xor U16656 (N_16656,N_15389,N_15461);
nand U16657 (N_16657,N_15771,N_15457);
xnor U16658 (N_16658,N_15402,N_15043);
or U16659 (N_16659,N_15083,N_15229);
or U16660 (N_16660,N_15906,N_15571);
and U16661 (N_16661,N_15471,N_15812);
nand U16662 (N_16662,N_15755,N_15263);
and U16663 (N_16663,N_15769,N_15048);
nor U16664 (N_16664,N_15698,N_15914);
nor U16665 (N_16665,N_15751,N_15846);
nor U16666 (N_16666,N_15147,N_15404);
nand U16667 (N_16667,N_15740,N_15636);
nand U16668 (N_16668,N_15619,N_15732);
and U16669 (N_16669,N_15095,N_15000);
xnor U16670 (N_16670,N_15705,N_15639);
nor U16671 (N_16671,N_15738,N_15474);
nor U16672 (N_16672,N_15706,N_15347);
xnor U16673 (N_16673,N_15613,N_15899);
or U16674 (N_16674,N_15718,N_15627);
and U16675 (N_16675,N_15426,N_15928);
or U16676 (N_16676,N_15947,N_15211);
and U16677 (N_16677,N_15075,N_15763);
and U16678 (N_16678,N_15959,N_15666);
nand U16679 (N_16679,N_15714,N_15716);
nand U16680 (N_16680,N_15451,N_15860);
xor U16681 (N_16681,N_15778,N_15303);
or U16682 (N_16682,N_15016,N_15261);
nor U16683 (N_16683,N_15911,N_15273);
and U16684 (N_16684,N_15171,N_15596);
nor U16685 (N_16685,N_15480,N_15047);
and U16686 (N_16686,N_15747,N_15962);
and U16687 (N_16687,N_15988,N_15115);
or U16688 (N_16688,N_15293,N_15274);
and U16689 (N_16689,N_15042,N_15473);
and U16690 (N_16690,N_15844,N_15823);
xnor U16691 (N_16691,N_15110,N_15833);
or U16692 (N_16692,N_15755,N_15246);
nor U16693 (N_16693,N_15003,N_15243);
nor U16694 (N_16694,N_15023,N_15772);
nor U16695 (N_16695,N_15310,N_15140);
and U16696 (N_16696,N_15153,N_15106);
or U16697 (N_16697,N_15965,N_15396);
and U16698 (N_16698,N_15428,N_15613);
nand U16699 (N_16699,N_15770,N_15147);
or U16700 (N_16700,N_15571,N_15021);
or U16701 (N_16701,N_15522,N_15669);
nor U16702 (N_16702,N_15430,N_15538);
or U16703 (N_16703,N_15649,N_15409);
nor U16704 (N_16704,N_15584,N_15209);
nand U16705 (N_16705,N_15744,N_15332);
nand U16706 (N_16706,N_15464,N_15646);
or U16707 (N_16707,N_15511,N_15826);
nor U16708 (N_16708,N_15947,N_15019);
and U16709 (N_16709,N_15764,N_15486);
nor U16710 (N_16710,N_15709,N_15629);
xor U16711 (N_16711,N_15187,N_15239);
nand U16712 (N_16712,N_15385,N_15871);
or U16713 (N_16713,N_15865,N_15597);
or U16714 (N_16714,N_15622,N_15369);
xnor U16715 (N_16715,N_15093,N_15153);
xor U16716 (N_16716,N_15553,N_15348);
xnor U16717 (N_16717,N_15168,N_15585);
xnor U16718 (N_16718,N_15050,N_15826);
or U16719 (N_16719,N_15531,N_15649);
or U16720 (N_16720,N_15302,N_15042);
and U16721 (N_16721,N_15988,N_15652);
and U16722 (N_16722,N_15199,N_15828);
xnor U16723 (N_16723,N_15570,N_15483);
nor U16724 (N_16724,N_15531,N_15105);
xor U16725 (N_16725,N_15317,N_15792);
or U16726 (N_16726,N_15914,N_15920);
and U16727 (N_16727,N_15447,N_15778);
nand U16728 (N_16728,N_15366,N_15941);
nor U16729 (N_16729,N_15019,N_15762);
and U16730 (N_16730,N_15746,N_15838);
or U16731 (N_16731,N_15174,N_15474);
xor U16732 (N_16732,N_15379,N_15080);
nand U16733 (N_16733,N_15291,N_15433);
nor U16734 (N_16734,N_15628,N_15305);
nand U16735 (N_16735,N_15252,N_15523);
nor U16736 (N_16736,N_15836,N_15819);
nor U16737 (N_16737,N_15051,N_15355);
or U16738 (N_16738,N_15447,N_15029);
xor U16739 (N_16739,N_15721,N_15905);
nand U16740 (N_16740,N_15942,N_15465);
nand U16741 (N_16741,N_15002,N_15405);
or U16742 (N_16742,N_15412,N_15032);
nor U16743 (N_16743,N_15759,N_15059);
or U16744 (N_16744,N_15066,N_15070);
xnor U16745 (N_16745,N_15990,N_15168);
xnor U16746 (N_16746,N_15410,N_15770);
xor U16747 (N_16747,N_15904,N_15467);
xor U16748 (N_16748,N_15538,N_15780);
or U16749 (N_16749,N_15439,N_15945);
and U16750 (N_16750,N_15676,N_15942);
xor U16751 (N_16751,N_15318,N_15956);
and U16752 (N_16752,N_15023,N_15649);
and U16753 (N_16753,N_15758,N_15727);
xnor U16754 (N_16754,N_15207,N_15569);
nor U16755 (N_16755,N_15429,N_15749);
xnor U16756 (N_16756,N_15158,N_15144);
nand U16757 (N_16757,N_15338,N_15678);
nand U16758 (N_16758,N_15986,N_15924);
and U16759 (N_16759,N_15701,N_15514);
nand U16760 (N_16760,N_15650,N_15439);
nand U16761 (N_16761,N_15606,N_15774);
and U16762 (N_16762,N_15605,N_15908);
or U16763 (N_16763,N_15072,N_15974);
or U16764 (N_16764,N_15773,N_15753);
xnor U16765 (N_16765,N_15178,N_15297);
or U16766 (N_16766,N_15688,N_15005);
xor U16767 (N_16767,N_15205,N_15782);
nor U16768 (N_16768,N_15139,N_15156);
nor U16769 (N_16769,N_15658,N_15698);
and U16770 (N_16770,N_15362,N_15269);
and U16771 (N_16771,N_15945,N_15925);
or U16772 (N_16772,N_15852,N_15308);
nand U16773 (N_16773,N_15822,N_15703);
nor U16774 (N_16774,N_15279,N_15689);
xnor U16775 (N_16775,N_15003,N_15705);
xnor U16776 (N_16776,N_15920,N_15726);
or U16777 (N_16777,N_15293,N_15665);
nand U16778 (N_16778,N_15544,N_15847);
nor U16779 (N_16779,N_15905,N_15753);
xor U16780 (N_16780,N_15730,N_15454);
xnor U16781 (N_16781,N_15766,N_15896);
xnor U16782 (N_16782,N_15633,N_15102);
nand U16783 (N_16783,N_15594,N_15492);
xor U16784 (N_16784,N_15474,N_15332);
xnor U16785 (N_16785,N_15445,N_15285);
nor U16786 (N_16786,N_15635,N_15094);
or U16787 (N_16787,N_15789,N_15959);
nor U16788 (N_16788,N_15793,N_15132);
nor U16789 (N_16789,N_15824,N_15821);
or U16790 (N_16790,N_15304,N_15848);
nor U16791 (N_16791,N_15828,N_15806);
nor U16792 (N_16792,N_15065,N_15823);
xnor U16793 (N_16793,N_15802,N_15863);
nor U16794 (N_16794,N_15338,N_15520);
xor U16795 (N_16795,N_15358,N_15387);
and U16796 (N_16796,N_15567,N_15459);
nor U16797 (N_16797,N_15569,N_15317);
nand U16798 (N_16798,N_15378,N_15549);
and U16799 (N_16799,N_15859,N_15362);
nor U16800 (N_16800,N_15079,N_15544);
and U16801 (N_16801,N_15925,N_15204);
and U16802 (N_16802,N_15444,N_15253);
xor U16803 (N_16803,N_15378,N_15913);
nor U16804 (N_16804,N_15789,N_15666);
or U16805 (N_16805,N_15067,N_15979);
xnor U16806 (N_16806,N_15349,N_15342);
and U16807 (N_16807,N_15569,N_15457);
nand U16808 (N_16808,N_15236,N_15469);
xnor U16809 (N_16809,N_15168,N_15519);
nor U16810 (N_16810,N_15881,N_15623);
and U16811 (N_16811,N_15339,N_15141);
or U16812 (N_16812,N_15424,N_15137);
xnor U16813 (N_16813,N_15428,N_15974);
or U16814 (N_16814,N_15977,N_15910);
nand U16815 (N_16815,N_15345,N_15840);
nand U16816 (N_16816,N_15125,N_15543);
xor U16817 (N_16817,N_15470,N_15036);
nand U16818 (N_16818,N_15229,N_15885);
or U16819 (N_16819,N_15998,N_15204);
nor U16820 (N_16820,N_15399,N_15862);
and U16821 (N_16821,N_15759,N_15653);
nor U16822 (N_16822,N_15990,N_15334);
nand U16823 (N_16823,N_15548,N_15114);
nor U16824 (N_16824,N_15700,N_15542);
xnor U16825 (N_16825,N_15762,N_15352);
nor U16826 (N_16826,N_15006,N_15461);
nor U16827 (N_16827,N_15298,N_15356);
nand U16828 (N_16828,N_15132,N_15466);
or U16829 (N_16829,N_15908,N_15837);
xor U16830 (N_16830,N_15242,N_15358);
and U16831 (N_16831,N_15103,N_15729);
nand U16832 (N_16832,N_15894,N_15557);
xnor U16833 (N_16833,N_15654,N_15915);
nand U16834 (N_16834,N_15802,N_15912);
and U16835 (N_16835,N_15039,N_15870);
nor U16836 (N_16836,N_15922,N_15086);
xor U16837 (N_16837,N_15268,N_15415);
nor U16838 (N_16838,N_15364,N_15510);
nand U16839 (N_16839,N_15824,N_15179);
or U16840 (N_16840,N_15965,N_15155);
xnor U16841 (N_16841,N_15385,N_15003);
xor U16842 (N_16842,N_15040,N_15558);
nor U16843 (N_16843,N_15947,N_15429);
or U16844 (N_16844,N_15808,N_15414);
and U16845 (N_16845,N_15635,N_15749);
xor U16846 (N_16846,N_15269,N_15361);
or U16847 (N_16847,N_15242,N_15023);
and U16848 (N_16848,N_15778,N_15786);
or U16849 (N_16849,N_15636,N_15212);
nor U16850 (N_16850,N_15779,N_15467);
nand U16851 (N_16851,N_15280,N_15713);
nor U16852 (N_16852,N_15095,N_15111);
and U16853 (N_16853,N_15986,N_15960);
xor U16854 (N_16854,N_15511,N_15423);
and U16855 (N_16855,N_15701,N_15958);
nand U16856 (N_16856,N_15707,N_15175);
nand U16857 (N_16857,N_15610,N_15431);
nor U16858 (N_16858,N_15614,N_15938);
or U16859 (N_16859,N_15271,N_15420);
or U16860 (N_16860,N_15247,N_15757);
nand U16861 (N_16861,N_15752,N_15001);
nor U16862 (N_16862,N_15008,N_15602);
xnor U16863 (N_16863,N_15507,N_15184);
and U16864 (N_16864,N_15182,N_15882);
xor U16865 (N_16865,N_15771,N_15605);
nand U16866 (N_16866,N_15832,N_15737);
nor U16867 (N_16867,N_15302,N_15506);
xor U16868 (N_16868,N_15391,N_15824);
nor U16869 (N_16869,N_15359,N_15288);
nand U16870 (N_16870,N_15460,N_15082);
nor U16871 (N_16871,N_15324,N_15343);
nand U16872 (N_16872,N_15623,N_15871);
nand U16873 (N_16873,N_15486,N_15127);
nand U16874 (N_16874,N_15231,N_15643);
xor U16875 (N_16875,N_15005,N_15417);
nand U16876 (N_16876,N_15579,N_15851);
and U16877 (N_16877,N_15191,N_15619);
and U16878 (N_16878,N_15560,N_15543);
xor U16879 (N_16879,N_15259,N_15378);
xor U16880 (N_16880,N_15996,N_15085);
and U16881 (N_16881,N_15902,N_15455);
or U16882 (N_16882,N_15966,N_15171);
or U16883 (N_16883,N_15734,N_15298);
nor U16884 (N_16884,N_15093,N_15776);
nand U16885 (N_16885,N_15171,N_15433);
nand U16886 (N_16886,N_15312,N_15603);
and U16887 (N_16887,N_15037,N_15796);
xor U16888 (N_16888,N_15528,N_15678);
or U16889 (N_16889,N_15436,N_15964);
or U16890 (N_16890,N_15428,N_15107);
and U16891 (N_16891,N_15367,N_15146);
xor U16892 (N_16892,N_15632,N_15582);
or U16893 (N_16893,N_15479,N_15288);
nor U16894 (N_16894,N_15582,N_15894);
xor U16895 (N_16895,N_15032,N_15282);
and U16896 (N_16896,N_15053,N_15346);
xor U16897 (N_16897,N_15426,N_15602);
or U16898 (N_16898,N_15416,N_15247);
and U16899 (N_16899,N_15025,N_15379);
nor U16900 (N_16900,N_15882,N_15333);
nor U16901 (N_16901,N_15207,N_15894);
or U16902 (N_16902,N_15299,N_15029);
and U16903 (N_16903,N_15749,N_15651);
and U16904 (N_16904,N_15597,N_15829);
and U16905 (N_16905,N_15212,N_15697);
or U16906 (N_16906,N_15214,N_15345);
nor U16907 (N_16907,N_15782,N_15495);
or U16908 (N_16908,N_15884,N_15613);
nor U16909 (N_16909,N_15831,N_15078);
and U16910 (N_16910,N_15381,N_15757);
nor U16911 (N_16911,N_15902,N_15102);
or U16912 (N_16912,N_15868,N_15396);
or U16913 (N_16913,N_15246,N_15541);
nor U16914 (N_16914,N_15999,N_15411);
xor U16915 (N_16915,N_15642,N_15756);
and U16916 (N_16916,N_15245,N_15676);
xor U16917 (N_16917,N_15746,N_15653);
and U16918 (N_16918,N_15742,N_15200);
xor U16919 (N_16919,N_15682,N_15392);
nor U16920 (N_16920,N_15794,N_15954);
and U16921 (N_16921,N_15091,N_15707);
nand U16922 (N_16922,N_15332,N_15200);
nand U16923 (N_16923,N_15397,N_15405);
and U16924 (N_16924,N_15622,N_15001);
nand U16925 (N_16925,N_15689,N_15202);
and U16926 (N_16926,N_15008,N_15605);
or U16927 (N_16927,N_15298,N_15030);
nand U16928 (N_16928,N_15106,N_15200);
or U16929 (N_16929,N_15393,N_15365);
and U16930 (N_16930,N_15877,N_15227);
nand U16931 (N_16931,N_15657,N_15510);
or U16932 (N_16932,N_15214,N_15134);
xor U16933 (N_16933,N_15889,N_15841);
nor U16934 (N_16934,N_15912,N_15473);
and U16935 (N_16935,N_15582,N_15793);
nand U16936 (N_16936,N_15481,N_15007);
nand U16937 (N_16937,N_15443,N_15122);
or U16938 (N_16938,N_15643,N_15302);
nor U16939 (N_16939,N_15975,N_15812);
or U16940 (N_16940,N_15042,N_15091);
or U16941 (N_16941,N_15496,N_15748);
nor U16942 (N_16942,N_15672,N_15902);
and U16943 (N_16943,N_15217,N_15068);
nor U16944 (N_16944,N_15849,N_15956);
and U16945 (N_16945,N_15662,N_15179);
xor U16946 (N_16946,N_15280,N_15203);
and U16947 (N_16947,N_15427,N_15152);
and U16948 (N_16948,N_15464,N_15638);
xor U16949 (N_16949,N_15830,N_15921);
xor U16950 (N_16950,N_15258,N_15752);
or U16951 (N_16951,N_15904,N_15774);
and U16952 (N_16952,N_15719,N_15084);
nand U16953 (N_16953,N_15283,N_15640);
and U16954 (N_16954,N_15650,N_15935);
or U16955 (N_16955,N_15827,N_15021);
and U16956 (N_16956,N_15419,N_15753);
and U16957 (N_16957,N_15177,N_15475);
and U16958 (N_16958,N_15508,N_15488);
nor U16959 (N_16959,N_15217,N_15965);
nand U16960 (N_16960,N_15603,N_15913);
and U16961 (N_16961,N_15351,N_15157);
xor U16962 (N_16962,N_15023,N_15777);
or U16963 (N_16963,N_15168,N_15663);
or U16964 (N_16964,N_15071,N_15824);
nor U16965 (N_16965,N_15995,N_15005);
or U16966 (N_16966,N_15610,N_15619);
xnor U16967 (N_16967,N_15061,N_15732);
nand U16968 (N_16968,N_15548,N_15415);
and U16969 (N_16969,N_15586,N_15671);
nor U16970 (N_16970,N_15164,N_15273);
nand U16971 (N_16971,N_15435,N_15358);
nor U16972 (N_16972,N_15245,N_15836);
nand U16973 (N_16973,N_15869,N_15838);
and U16974 (N_16974,N_15853,N_15672);
nor U16975 (N_16975,N_15847,N_15245);
nand U16976 (N_16976,N_15154,N_15365);
nand U16977 (N_16977,N_15549,N_15971);
or U16978 (N_16978,N_15155,N_15598);
or U16979 (N_16979,N_15610,N_15615);
or U16980 (N_16980,N_15824,N_15195);
nand U16981 (N_16981,N_15378,N_15165);
nand U16982 (N_16982,N_15450,N_15890);
nand U16983 (N_16983,N_15292,N_15748);
or U16984 (N_16984,N_15955,N_15892);
or U16985 (N_16985,N_15084,N_15247);
or U16986 (N_16986,N_15417,N_15332);
nand U16987 (N_16987,N_15210,N_15908);
or U16988 (N_16988,N_15133,N_15577);
nor U16989 (N_16989,N_15059,N_15637);
or U16990 (N_16990,N_15244,N_15522);
nand U16991 (N_16991,N_15547,N_15906);
xor U16992 (N_16992,N_15483,N_15309);
xnor U16993 (N_16993,N_15245,N_15749);
nor U16994 (N_16994,N_15724,N_15145);
xor U16995 (N_16995,N_15616,N_15335);
xor U16996 (N_16996,N_15659,N_15916);
or U16997 (N_16997,N_15455,N_15734);
or U16998 (N_16998,N_15760,N_15923);
nor U16999 (N_16999,N_15662,N_15321);
nor U17000 (N_17000,N_16300,N_16887);
nand U17001 (N_17001,N_16313,N_16306);
or U17002 (N_17002,N_16374,N_16603);
xnor U17003 (N_17003,N_16153,N_16639);
xnor U17004 (N_17004,N_16742,N_16420);
or U17005 (N_17005,N_16921,N_16509);
or U17006 (N_17006,N_16382,N_16483);
or U17007 (N_17007,N_16668,N_16323);
nand U17008 (N_17008,N_16385,N_16314);
and U17009 (N_17009,N_16284,N_16293);
nor U17010 (N_17010,N_16452,N_16858);
and U17011 (N_17011,N_16677,N_16753);
nor U17012 (N_17012,N_16368,N_16772);
nor U17013 (N_17013,N_16156,N_16891);
and U17014 (N_17014,N_16130,N_16854);
nand U17015 (N_17015,N_16715,N_16451);
nand U17016 (N_17016,N_16612,N_16598);
or U17017 (N_17017,N_16683,N_16722);
or U17018 (N_17018,N_16619,N_16568);
nor U17019 (N_17019,N_16661,N_16594);
nor U17020 (N_17020,N_16209,N_16925);
or U17021 (N_17021,N_16946,N_16103);
xnor U17022 (N_17022,N_16795,N_16411);
or U17023 (N_17023,N_16519,N_16131);
nand U17024 (N_17024,N_16232,N_16225);
nor U17025 (N_17025,N_16345,N_16947);
nor U17026 (N_17026,N_16790,N_16062);
nor U17027 (N_17027,N_16309,N_16781);
and U17028 (N_17028,N_16839,N_16029);
or U17029 (N_17029,N_16535,N_16750);
and U17030 (N_17030,N_16855,N_16964);
nor U17031 (N_17031,N_16364,N_16104);
nor U17032 (N_17032,N_16129,N_16278);
nand U17033 (N_17033,N_16813,N_16967);
nand U17034 (N_17034,N_16810,N_16558);
xor U17035 (N_17035,N_16554,N_16154);
xor U17036 (N_17036,N_16424,N_16695);
xnor U17037 (N_17037,N_16560,N_16935);
xnor U17038 (N_17038,N_16920,N_16767);
xnor U17039 (N_17039,N_16807,N_16146);
xnor U17040 (N_17040,N_16237,N_16408);
xnor U17041 (N_17041,N_16114,N_16570);
nand U17042 (N_17042,N_16550,N_16938);
nor U17043 (N_17043,N_16493,N_16692);
nand U17044 (N_17044,N_16797,N_16096);
or U17045 (N_17045,N_16526,N_16418);
and U17046 (N_17046,N_16291,N_16128);
xnor U17047 (N_17047,N_16516,N_16874);
or U17048 (N_17048,N_16914,N_16965);
and U17049 (N_17049,N_16702,N_16466);
nand U17050 (N_17050,N_16663,N_16456);
nor U17051 (N_17051,N_16758,N_16630);
or U17052 (N_17052,N_16700,N_16143);
xor U17053 (N_17053,N_16703,N_16489);
nor U17054 (N_17054,N_16913,N_16377);
or U17055 (N_17055,N_16744,N_16281);
xnor U17056 (N_17056,N_16206,N_16730);
or U17057 (N_17057,N_16735,N_16267);
or U17058 (N_17058,N_16575,N_16358);
and U17059 (N_17059,N_16419,N_16680);
and U17060 (N_17060,N_16490,N_16701);
nand U17061 (N_17061,N_16273,N_16361);
xnor U17062 (N_17062,N_16595,N_16982);
nand U17063 (N_17063,N_16567,N_16572);
or U17064 (N_17064,N_16997,N_16097);
and U17065 (N_17065,N_16067,N_16876);
or U17066 (N_17066,N_16537,N_16244);
nor U17067 (N_17067,N_16823,N_16638);
and U17068 (N_17068,N_16211,N_16510);
and U17069 (N_17069,N_16410,N_16402);
and U17070 (N_17070,N_16773,N_16287);
xnor U17071 (N_17071,N_16939,N_16307);
and U17072 (N_17072,N_16474,N_16963);
nand U17073 (N_17073,N_16923,N_16806);
nor U17074 (N_17074,N_16936,N_16039);
or U17075 (N_17075,N_16138,N_16221);
and U17076 (N_17076,N_16427,N_16401);
and U17077 (N_17077,N_16593,N_16829);
and U17078 (N_17078,N_16447,N_16094);
or U17079 (N_17079,N_16018,N_16833);
and U17080 (N_17080,N_16940,N_16149);
or U17081 (N_17081,N_16251,N_16768);
and U17082 (N_17082,N_16738,N_16249);
or U17083 (N_17083,N_16125,N_16999);
and U17084 (N_17084,N_16969,N_16332);
and U17085 (N_17085,N_16849,N_16126);
xnor U17086 (N_17086,N_16384,N_16988);
xnor U17087 (N_17087,N_16328,N_16588);
and U17088 (N_17088,N_16532,N_16369);
nor U17089 (N_17089,N_16205,N_16437);
nand U17090 (N_17090,N_16670,N_16405);
or U17091 (N_17091,N_16687,N_16892);
or U17092 (N_17092,N_16116,N_16301);
and U17093 (N_17093,N_16805,N_16587);
or U17094 (N_17094,N_16137,N_16170);
nor U17095 (N_17095,N_16983,N_16718);
or U17096 (N_17096,N_16083,N_16778);
nand U17097 (N_17097,N_16743,N_16416);
or U17098 (N_17098,N_16217,N_16981);
and U17099 (N_17099,N_16848,N_16446);
and U17100 (N_17100,N_16178,N_16118);
nand U17101 (N_17101,N_16055,N_16023);
or U17102 (N_17102,N_16478,N_16366);
and U17103 (N_17103,N_16499,N_16404);
xnor U17104 (N_17104,N_16783,N_16615);
nor U17105 (N_17105,N_16792,N_16780);
nor U17106 (N_17106,N_16026,N_16580);
nand U17107 (N_17107,N_16257,N_16801);
xor U17108 (N_17108,N_16106,N_16247);
xnor U17109 (N_17109,N_16196,N_16471);
and U17110 (N_17110,N_16423,N_16144);
xor U17111 (N_17111,N_16037,N_16763);
nand U17112 (N_17112,N_16911,N_16065);
nor U17113 (N_17113,N_16534,N_16505);
xnor U17114 (N_17114,N_16539,N_16367);
xor U17115 (N_17115,N_16406,N_16658);
xnor U17116 (N_17116,N_16190,N_16748);
nand U17117 (N_17117,N_16354,N_16803);
nand U17118 (N_17118,N_16950,N_16871);
nor U17119 (N_17119,N_16504,N_16228);
xor U17120 (N_17120,N_16540,N_16652);
and U17121 (N_17121,N_16990,N_16977);
nand U17122 (N_17122,N_16253,N_16684);
or U17123 (N_17123,N_16769,N_16460);
nand U17124 (N_17124,N_16704,N_16559);
and U17125 (N_17125,N_16996,N_16252);
or U17126 (N_17126,N_16953,N_16045);
nor U17127 (N_17127,N_16458,N_16941);
xor U17128 (N_17128,N_16186,N_16787);
or U17129 (N_17129,N_16850,N_16616);
nor U17130 (N_17130,N_16283,N_16095);
or U17131 (N_17131,N_16525,N_16432);
nand U17132 (N_17132,N_16583,N_16169);
nor U17133 (N_17133,N_16047,N_16290);
nand U17134 (N_17134,N_16012,N_16811);
and U17135 (N_17135,N_16127,N_16245);
and U17136 (N_17136,N_16676,N_16959);
and U17137 (N_17137,N_16714,N_16394);
or U17138 (N_17138,N_16573,N_16207);
nand U17139 (N_17139,N_16980,N_16521);
xor U17140 (N_17140,N_16098,N_16482);
nor U17141 (N_17141,N_16148,N_16870);
and U17142 (N_17142,N_16948,N_16958);
nand U17143 (N_17143,N_16238,N_16896);
nor U17144 (N_17144,N_16187,N_16317);
and U17145 (N_17145,N_16229,N_16142);
xor U17146 (N_17146,N_16929,N_16707);
xnor U17147 (N_17147,N_16720,N_16756);
nor U17148 (N_17148,N_16117,N_16362);
or U17149 (N_17149,N_16476,N_16020);
nand U17150 (N_17150,N_16224,N_16865);
xor U17151 (N_17151,N_16285,N_16017);
xor U17152 (N_17152,N_16475,N_16721);
nor U17153 (N_17153,N_16181,N_16694);
and U17154 (N_17154,N_16544,N_16623);
xnor U17155 (N_17155,N_16949,N_16183);
xor U17156 (N_17156,N_16841,N_16336);
nand U17157 (N_17157,N_16355,N_16121);
or U17158 (N_17158,N_16705,N_16133);
or U17159 (N_17159,N_16011,N_16465);
nor U17160 (N_17160,N_16412,N_16193);
nand U17161 (N_17161,N_16024,N_16837);
nand U17162 (N_17162,N_16524,N_16847);
xnor U17163 (N_17163,N_16533,N_16264);
xor U17164 (N_17164,N_16302,N_16150);
nor U17165 (N_17165,N_16034,N_16500);
nand U17166 (N_17166,N_16932,N_16576);
xor U17167 (N_17167,N_16088,N_16254);
xnor U17168 (N_17168,N_16972,N_16216);
xor U17169 (N_17169,N_16889,N_16242);
or U17170 (N_17170,N_16726,N_16513);
and U17171 (N_17171,N_16713,N_16966);
xnor U17172 (N_17172,N_16443,N_16734);
nand U17173 (N_17173,N_16777,N_16370);
nand U17174 (N_17174,N_16799,N_16072);
nor U17175 (N_17175,N_16809,N_16485);
xnor U17176 (N_17176,N_16994,N_16888);
and U17177 (N_17177,N_16454,N_16657);
and U17178 (N_17178,N_16484,N_16357);
nand U17179 (N_17179,N_16863,N_16134);
and U17180 (N_17180,N_16698,N_16873);
and U17181 (N_17181,N_16884,N_16076);
and U17182 (N_17182,N_16538,N_16943);
nor U17183 (N_17183,N_16340,N_16041);
or U17184 (N_17184,N_16299,N_16472);
nand U17185 (N_17185,N_16189,N_16227);
and U17186 (N_17186,N_16162,N_16650);
xor U17187 (N_17187,N_16344,N_16415);
and U17188 (N_17188,N_16656,N_16312);
xnor U17189 (N_17189,N_16165,N_16877);
nor U17190 (N_17190,N_16802,N_16511);
or U17191 (N_17191,N_16015,N_16102);
or U17192 (N_17192,N_16733,N_16388);
xor U17193 (N_17193,N_16099,N_16172);
or U17194 (N_17194,N_16425,N_16686);
nand U17195 (N_17195,N_16068,N_16602);
xor U17196 (N_17196,N_16845,N_16185);
and U17197 (N_17197,N_16961,N_16449);
or U17198 (N_17198,N_16915,N_16897);
xor U17199 (N_17199,N_16000,N_16448);
xnor U17200 (N_17200,N_16275,N_16671);
or U17201 (N_17201,N_16399,N_16978);
and U17202 (N_17202,N_16584,N_16581);
nand U17203 (N_17203,N_16331,N_16001);
xnor U17204 (N_17204,N_16334,N_16577);
nor U17205 (N_17205,N_16856,N_16298);
or U17206 (N_17206,N_16723,N_16634);
nand U17207 (N_17207,N_16201,N_16578);
and U17208 (N_17208,N_16033,N_16842);
nor U17209 (N_17209,N_16151,N_16880);
or U17210 (N_17210,N_16708,N_16645);
or U17211 (N_17211,N_16157,N_16392);
or U17212 (N_17212,N_16168,N_16112);
xor U17213 (N_17213,N_16779,N_16642);
nand U17214 (N_17214,N_16831,N_16900);
or U17215 (N_17215,N_16327,N_16840);
or U17216 (N_17216,N_16646,N_16360);
nand U17217 (N_17217,N_16022,N_16916);
nand U17218 (N_17218,N_16755,N_16400);
xor U17219 (N_17219,N_16240,N_16725);
xnor U17220 (N_17220,N_16804,N_16564);
nand U17221 (N_17221,N_16667,N_16107);
or U17222 (N_17222,N_16295,N_16235);
xnor U17223 (N_17223,N_16473,N_16325);
and U17224 (N_17224,N_16551,N_16776);
nor U17225 (N_17225,N_16699,N_16766);
nand U17226 (N_17226,N_16737,N_16497);
and U17227 (N_17227,N_16494,N_16906);
xor U17228 (N_17228,N_16363,N_16825);
nor U17229 (N_17229,N_16100,N_16625);
nor U17230 (N_17230,N_16883,N_16260);
or U17231 (N_17231,N_16122,N_16395);
or U17232 (N_17232,N_16009,N_16674);
or U17233 (N_17233,N_16591,N_16732);
nand U17234 (N_17234,N_16901,N_16164);
nor U17235 (N_17235,N_16775,N_16324);
nor U17236 (N_17236,N_16786,N_16596);
or U17237 (N_17237,N_16241,N_16455);
nand U17238 (N_17238,N_16908,N_16860);
or U17239 (N_17239,N_16010,N_16202);
nand U17240 (N_17240,N_16651,N_16341);
and U17241 (N_17241,N_16294,N_16785);
nor U17242 (N_17242,N_16422,N_16115);
nand U17243 (N_17243,N_16933,N_16007);
nor U17244 (N_17244,N_16266,N_16035);
or U17245 (N_17245,N_16962,N_16822);
xor U17246 (N_17246,N_16794,N_16431);
nor U17247 (N_17247,N_16059,N_16259);
nor U17248 (N_17248,N_16407,N_16263);
nor U17249 (N_17249,N_16827,N_16751);
or U17250 (N_17250,N_16426,N_16330);
nor U17251 (N_17251,N_16176,N_16464);
nand U17252 (N_17252,N_16074,N_16951);
and U17253 (N_17253,N_16016,N_16859);
nor U17254 (N_17254,N_16706,N_16739);
nor U17255 (N_17255,N_16957,N_16869);
xnor U17256 (N_17256,N_16728,N_16665);
or U17257 (N_17257,N_16119,N_16653);
nor U17258 (N_17258,N_16073,N_16789);
or U17259 (N_17259,N_16907,N_16905);
nor U17260 (N_17260,N_16373,N_16614);
nand U17261 (N_17261,N_16673,N_16672);
nor U17262 (N_17262,N_16878,N_16381);
or U17263 (N_17263,N_16643,N_16712);
or U17264 (N_17264,N_16648,N_16279);
and U17265 (N_17265,N_16389,N_16346);
and U17266 (N_17266,N_16640,N_16043);
or U17267 (N_17267,N_16895,N_16882);
xor U17268 (N_17268,N_16879,N_16140);
and U17269 (N_17269,N_16993,N_16711);
or U17270 (N_17270,N_16246,N_16480);
nand U17271 (N_17271,N_16761,N_16231);
and U17272 (N_17272,N_16042,N_16163);
nor U17273 (N_17273,N_16214,N_16005);
and U17274 (N_17274,N_16199,N_16380);
nand U17275 (N_17275,N_16740,N_16036);
or U17276 (N_17276,N_16061,N_16468);
nand U17277 (N_17277,N_16028,N_16203);
nor U17278 (N_17278,N_16991,N_16080);
nor U17279 (N_17279,N_16433,N_16147);
and U17280 (N_17280,N_16944,N_16215);
and U17281 (N_17281,N_16132,N_16089);
nand U17282 (N_17282,N_16436,N_16729);
and U17283 (N_17283,N_16501,N_16812);
or U17284 (N_17284,N_16265,N_16716);
xor U17285 (N_17285,N_16498,N_16457);
and U17286 (N_17286,N_16788,N_16815);
xnor U17287 (N_17287,N_16180,N_16867);
and U17288 (N_17288,N_16152,N_16335);
and U17289 (N_17289,N_16430,N_16931);
xnor U17290 (N_17290,N_16838,N_16784);
and U17291 (N_17291,N_16862,N_16754);
nand U17292 (N_17292,N_16014,N_16664);
nand U17293 (N_17293,N_16890,N_16543);
xor U17294 (N_17294,N_16428,N_16269);
and U17295 (N_17295,N_16338,N_16629);
and U17296 (N_17296,N_16613,N_16391);
nand U17297 (N_17297,N_16379,N_16030);
and U17298 (N_17298,N_16208,N_16542);
xnor U17299 (N_17299,N_16678,N_16904);
and U17300 (N_17300,N_16681,N_16626);
or U17301 (N_17301,N_16469,N_16912);
or U17302 (N_17302,N_16851,N_16566);
nor U17303 (N_17303,N_16624,N_16124);
nor U17304 (N_17304,N_16320,N_16998);
nor U17305 (N_17305,N_16002,N_16976);
or U17306 (N_17306,N_16610,N_16968);
nor U17307 (N_17307,N_16038,N_16166);
and U17308 (N_17308,N_16343,N_16297);
and U17309 (N_17309,N_16601,N_16796);
nand U17310 (N_17310,N_16606,N_16903);
nor U17311 (N_17311,N_16770,N_16282);
nand U17312 (N_17312,N_16173,N_16919);
xor U17313 (N_17313,N_16523,N_16937);
or U17314 (N_17314,N_16622,N_16375);
or U17315 (N_17315,N_16063,N_16258);
or U17316 (N_17316,N_16492,N_16442);
and U17317 (N_17317,N_16226,N_16844);
xnor U17318 (N_17318,N_16262,N_16852);
nor U17319 (N_17319,N_16371,N_16204);
or U17320 (N_17320,N_16421,N_16696);
xor U17321 (N_17321,N_16496,N_16111);
xor U17322 (N_17322,N_16049,N_16644);
nor U17323 (N_17323,N_16618,N_16691);
or U17324 (N_17324,N_16818,N_16192);
or U17325 (N_17325,N_16835,N_16989);
or U17326 (N_17326,N_16349,N_16508);
xnor U17327 (N_17327,N_16086,N_16308);
nor U17328 (N_17328,N_16372,N_16814);
nor U17329 (N_17329,N_16548,N_16082);
nor U17330 (N_17330,N_16556,N_16893);
or U17331 (N_17331,N_16502,N_16270);
nand U17332 (N_17332,N_16316,N_16329);
xnor U17333 (N_17333,N_16477,N_16321);
or U17334 (N_17334,N_16633,N_16326);
xnor U17335 (N_17335,N_16585,N_16945);
xnor U17336 (N_17336,N_16710,N_16597);
nor U17337 (N_17337,N_16296,N_16599);
nand U17338 (N_17338,N_16288,N_16177);
nor U17339 (N_17339,N_16467,N_16025);
xor U17340 (N_17340,N_16857,N_16960);
nand U17341 (N_17341,N_16386,N_16736);
or U17342 (N_17342,N_16158,N_16987);
nand U17343 (N_17343,N_16182,N_16974);
nand U17344 (N_17344,N_16175,N_16752);
or U17345 (N_17345,N_16574,N_16236);
xor U17346 (N_17346,N_16188,N_16481);
nand U17347 (N_17347,N_16760,N_16463);
xor U17348 (N_17348,N_16075,N_16955);
or U17349 (N_17349,N_16435,N_16620);
nor U17350 (N_17350,N_16090,N_16289);
or U17351 (N_17351,N_16557,N_16070);
and U17352 (N_17352,N_16444,N_16579);
nor U17353 (N_17353,N_16654,N_16984);
xor U17354 (N_17354,N_16649,N_16954);
and U17355 (N_17355,N_16046,N_16636);
nor U17356 (N_17356,N_16834,N_16396);
and U17357 (N_17357,N_16004,N_16210);
xnor U17358 (N_17358,N_16611,N_16495);
nor U17359 (N_17359,N_16110,N_16079);
or U17360 (N_17360,N_16604,N_16975);
xnor U17361 (N_17361,N_16135,N_16052);
or U17362 (N_17362,N_16414,N_16662);
nor U17363 (N_17363,N_16348,N_16197);
or U17364 (N_17364,N_16592,N_16487);
xnor U17365 (N_17365,N_16462,N_16569);
xnor U17366 (N_17366,N_16184,N_16413);
nor U17367 (N_17367,N_16479,N_16136);
nand U17368 (N_17368,N_16219,N_16220);
nor U17369 (N_17369,N_16924,N_16627);
or U17370 (N_17370,N_16899,N_16562);
or U17371 (N_17371,N_16549,N_16351);
nor U17372 (N_17372,N_16223,N_16440);
and U17373 (N_17373,N_16319,N_16350);
nand U17374 (N_17374,N_16546,N_16830);
xor U17375 (N_17375,N_16040,N_16459);
or U17376 (N_17376,N_16057,N_16843);
xor U17377 (N_17377,N_16641,N_16545);
nand U17378 (N_17378,N_16439,N_16048);
xnor U17379 (N_17379,N_16085,N_16697);
nor U17380 (N_17380,N_16992,N_16727);
nand U17381 (N_17381,N_16305,N_16450);
xor U17382 (N_17382,N_16749,N_16084);
xor U17383 (N_17383,N_16488,N_16970);
nor U17384 (N_17384,N_16491,N_16200);
nor U17385 (N_17385,N_16058,N_16167);
nand U17386 (N_17386,N_16066,N_16621);
and U17387 (N_17387,N_16782,N_16311);
nor U17388 (N_17388,N_16861,N_16218);
xor U17389 (N_17389,N_16635,N_16666);
xnor U17390 (N_17390,N_16682,N_16222);
nor U17391 (N_17391,N_16926,N_16304);
and U17392 (N_17392,N_16902,N_16213);
and U17393 (N_17393,N_16376,N_16605);
nor U17394 (N_17394,N_16986,N_16515);
and U17395 (N_17395,N_16280,N_16409);
or U17396 (N_17396,N_16179,N_16764);
and U17397 (N_17397,N_16745,N_16171);
nor U17398 (N_17398,N_16832,N_16589);
xor U17399 (N_17399,N_16105,N_16816);
xnor U17400 (N_17400,N_16875,N_16255);
nor U17401 (N_17401,N_16318,N_16631);
or U17402 (N_17402,N_16031,N_16159);
or U17403 (N_17403,N_16292,N_16675);
or U17404 (N_17404,N_16952,N_16693);
or U17405 (N_17405,N_16250,N_16141);
or U17406 (N_17406,N_16013,N_16774);
and U17407 (N_17407,N_16113,N_16243);
nor U17408 (N_17408,N_16234,N_16885);
or U17409 (N_17409,N_16365,N_16660);
nand U17410 (N_17410,N_16268,N_16719);
nand U17411 (N_17411,N_16536,N_16517);
or U17412 (N_17412,N_16918,N_16690);
nor U17413 (N_17413,N_16541,N_16195);
and U17414 (N_17414,N_16689,N_16390);
and U17415 (N_17415,N_16868,N_16310);
nand U17416 (N_17416,N_16765,N_16383);
or U17417 (N_17417,N_16529,N_16194);
or U17418 (N_17418,N_16826,N_16909);
nor U17419 (N_17419,N_16590,N_16942);
nand U17420 (N_17420,N_16438,N_16659);
xnor U17421 (N_17421,N_16820,N_16518);
and U17422 (N_17422,N_16808,N_16359);
nor U17423 (N_17423,N_16092,N_16277);
nor U17424 (N_17424,N_16056,N_16506);
nand U17425 (N_17425,N_16928,N_16429);
or U17426 (N_17426,N_16724,N_16337);
or U17427 (N_17427,N_16342,N_16356);
nor U17428 (N_17428,N_16417,N_16050);
or U17429 (N_17429,N_16637,N_16378);
nor U17430 (N_17430,N_16757,N_16528);
or U17431 (N_17431,N_16824,N_16019);
nand U17432 (N_17432,N_16393,N_16160);
xor U17433 (N_17433,N_16565,N_16434);
nor U17434 (N_17434,N_16685,N_16817);
and U17435 (N_17435,N_16741,N_16387);
nor U17436 (N_17436,N_16995,N_16607);
nor U17437 (N_17437,N_16552,N_16339);
xor U17438 (N_17438,N_16800,N_16617);
nor U17439 (N_17439,N_16979,N_16791);
and U17440 (N_17440,N_16239,N_16248);
xnor U17441 (N_17441,N_16044,N_16647);
nor U17442 (N_17442,N_16161,N_16828);
and U17443 (N_17443,N_16403,N_16212);
nor U17444 (N_17444,N_16233,N_16322);
or U17445 (N_17445,N_16709,N_16553);
nand U17446 (N_17446,N_16453,N_16032);
nor U17447 (N_17447,N_16441,N_16060);
and U17448 (N_17448,N_16917,N_16191);
nand U17449 (N_17449,N_16486,N_16898);
nor U17450 (N_17450,N_16563,N_16628);
nand U17451 (N_17451,N_16520,N_16120);
or U17452 (N_17452,N_16717,N_16108);
or U17453 (N_17453,N_16333,N_16819);
nor U17454 (N_17454,N_16793,N_16922);
or U17455 (N_17455,N_16139,N_16461);
or U17456 (N_17456,N_16398,N_16971);
xnor U17457 (N_17457,N_16821,N_16078);
xnor U17458 (N_17458,N_16101,N_16527);
xnor U17459 (N_17459,N_16272,N_16145);
xor U17460 (N_17460,N_16093,N_16276);
nand U17461 (N_17461,N_16522,N_16027);
xnor U17462 (N_17462,N_16230,N_16655);
nand U17463 (N_17463,N_16198,N_16747);
or U17464 (N_17464,N_16051,N_16956);
or U17465 (N_17465,N_16530,N_16561);
nor U17466 (N_17466,N_16006,N_16872);
xnor U17467 (N_17467,N_16846,N_16445);
nand U17468 (N_17468,N_16985,N_16669);
or U17469 (N_17469,N_16347,N_16746);
nor U17470 (N_17470,N_16512,N_16927);
and U17471 (N_17471,N_16771,N_16064);
nand U17472 (N_17472,N_16608,N_16547);
xor U17473 (N_17473,N_16762,N_16109);
and U17474 (N_17474,N_16836,N_16054);
or U17475 (N_17475,N_16600,N_16759);
and U17476 (N_17476,N_16353,N_16053);
or U17477 (N_17477,N_16087,N_16003);
and U17478 (N_17478,N_16174,N_16688);
nor U17479 (N_17479,N_16886,N_16571);
nor U17480 (N_17480,N_16397,N_16866);
and U17481 (N_17481,N_16555,N_16582);
nor U17482 (N_17482,N_16256,N_16503);
nor U17483 (N_17483,N_16123,N_16271);
or U17484 (N_17484,N_16081,N_16632);
xor U17485 (N_17485,N_16731,N_16514);
nand U17486 (N_17486,N_16069,N_16973);
and U17487 (N_17487,N_16470,N_16261);
nor U17488 (N_17488,N_16315,N_16077);
and U17489 (N_17489,N_16091,N_16894);
nor U17490 (N_17490,N_16303,N_16798);
nand U17491 (N_17491,N_16609,N_16071);
nor U17492 (N_17492,N_16155,N_16930);
nand U17493 (N_17493,N_16531,N_16507);
or U17494 (N_17494,N_16352,N_16881);
nor U17495 (N_17495,N_16586,N_16910);
and U17496 (N_17496,N_16008,N_16274);
nor U17497 (N_17497,N_16934,N_16853);
or U17498 (N_17498,N_16679,N_16864);
or U17499 (N_17499,N_16286,N_16021);
or U17500 (N_17500,N_16706,N_16195);
or U17501 (N_17501,N_16813,N_16425);
nor U17502 (N_17502,N_16943,N_16323);
xnor U17503 (N_17503,N_16323,N_16079);
nand U17504 (N_17504,N_16582,N_16294);
xor U17505 (N_17505,N_16612,N_16311);
and U17506 (N_17506,N_16603,N_16861);
or U17507 (N_17507,N_16570,N_16581);
or U17508 (N_17508,N_16191,N_16328);
nand U17509 (N_17509,N_16211,N_16470);
nor U17510 (N_17510,N_16502,N_16372);
nand U17511 (N_17511,N_16596,N_16918);
nor U17512 (N_17512,N_16093,N_16048);
and U17513 (N_17513,N_16508,N_16902);
and U17514 (N_17514,N_16448,N_16169);
nand U17515 (N_17515,N_16997,N_16093);
nor U17516 (N_17516,N_16437,N_16230);
and U17517 (N_17517,N_16702,N_16685);
or U17518 (N_17518,N_16615,N_16127);
and U17519 (N_17519,N_16858,N_16347);
and U17520 (N_17520,N_16591,N_16018);
xnor U17521 (N_17521,N_16900,N_16680);
or U17522 (N_17522,N_16927,N_16209);
nor U17523 (N_17523,N_16196,N_16558);
nor U17524 (N_17524,N_16001,N_16877);
or U17525 (N_17525,N_16062,N_16691);
nand U17526 (N_17526,N_16276,N_16448);
or U17527 (N_17527,N_16847,N_16699);
or U17528 (N_17528,N_16948,N_16917);
or U17529 (N_17529,N_16295,N_16206);
nor U17530 (N_17530,N_16037,N_16771);
xnor U17531 (N_17531,N_16176,N_16724);
xnor U17532 (N_17532,N_16835,N_16574);
nor U17533 (N_17533,N_16913,N_16544);
nand U17534 (N_17534,N_16492,N_16938);
and U17535 (N_17535,N_16889,N_16415);
and U17536 (N_17536,N_16949,N_16087);
xnor U17537 (N_17537,N_16545,N_16539);
or U17538 (N_17538,N_16408,N_16390);
or U17539 (N_17539,N_16224,N_16867);
xnor U17540 (N_17540,N_16912,N_16304);
xnor U17541 (N_17541,N_16859,N_16549);
nand U17542 (N_17542,N_16366,N_16504);
nor U17543 (N_17543,N_16156,N_16538);
and U17544 (N_17544,N_16461,N_16684);
and U17545 (N_17545,N_16300,N_16360);
and U17546 (N_17546,N_16571,N_16917);
nand U17547 (N_17547,N_16465,N_16185);
xnor U17548 (N_17548,N_16453,N_16857);
xor U17549 (N_17549,N_16330,N_16755);
and U17550 (N_17550,N_16855,N_16328);
or U17551 (N_17551,N_16143,N_16233);
and U17552 (N_17552,N_16508,N_16523);
nor U17553 (N_17553,N_16819,N_16203);
and U17554 (N_17554,N_16788,N_16126);
or U17555 (N_17555,N_16249,N_16861);
xnor U17556 (N_17556,N_16552,N_16071);
and U17557 (N_17557,N_16224,N_16086);
nand U17558 (N_17558,N_16727,N_16977);
xor U17559 (N_17559,N_16588,N_16639);
and U17560 (N_17560,N_16288,N_16145);
or U17561 (N_17561,N_16460,N_16024);
nand U17562 (N_17562,N_16841,N_16857);
xnor U17563 (N_17563,N_16358,N_16662);
and U17564 (N_17564,N_16874,N_16008);
nor U17565 (N_17565,N_16419,N_16739);
and U17566 (N_17566,N_16488,N_16718);
nand U17567 (N_17567,N_16356,N_16475);
nand U17568 (N_17568,N_16052,N_16104);
nand U17569 (N_17569,N_16582,N_16913);
or U17570 (N_17570,N_16966,N_16354);
or U17571 (N_17571,N_16095,N_16526);
nor U17572 (N_17572,N_16310,N_16603);
xor U17573 (N_17573,N_16095,N_16752);
nand U17574 (N_17574,N_16723,N_16608);
and U17575 (N_17575,N_16120,N_16641);
xor U17576 (N_17576,N_16035,N_16271);
nor U17577 (N_17577,N_16860,N_16201);
or U17578 (N_17578,N_16039,N_16222);
nor U17579 (N_17579,N_16000,N_16323);
xor U17580 (N_17580,N_16149,N_16360);
nor U17581 (N_17581,N_16847,N_16041);
nand U17582 (N_17582,N_16259,N_16695);
nand U17583 (N_17583,N_16925,N_16325);
or U17584 (N_17584,N_16548,N_16489);
and U17585 (N_17585,N_16012,N_16456);
xor U17586 (N_17586,N_16153,N_16377);
and U17587 (N_17587,N_16704,N_16551);
and U17588 (N_17588,N_16311,N_16369);
xor U17589 (N_17589,N_16362,N_16364);
or U17590 (N_17590,N_16154,N_16217);
xor U17591 (N_17591,N_16033,N_16816);
or U17592 (N_17592,N_16952,N_16296);
xor U17593 (N_17593,N_16895,N_16816);
xnor U17594 (N_17594,N_16873,N_16964);
and U17595 (N_17595,N_16242,N_16448);
nor U17596 (N_17596,N_16043,N_16618);
or U17597 (N_17597,N_16443,N_16212);
xor U17598 (N_17598,N_16016,N_16109);
or U17599 (N_17599,N_16021,N_16104);
xnor U17600 (N_17600,N_16075,N_16203);
xor U17601 (N_17601,N_16309,N_16038);
and U17602 (N_17602,N_16646,N_16096);
xor U17603 (N_17603,N_16885,N_16493);
nand U17604 (N_17604,N_16748,N_16409);
nand U17605 (N_17605,N_16903,N_16006);
xor U17606 (N_17606,N_16469,N_16580);
or U17607 (N_17607,N_16089,N_16243);
and U17608 (N_17608,N_16680,N_16164);
xnor U17609 (N_17609,N_16499,N_16269);
nand U17610 (N_17610,N_16575,N_16644);
and U17611 (N_17611,N_16497,N_16995);
nor U17612 (N_17612,N_16180,N_16763);
xor U17613 (N_17613,N_16886,N_16657);
xnor U17614 (N_17614,N_16220,N_16348);
nand U17615 (N_17615,N_16814,N_16845);
nor U17616 (N_17616,N_16455,N_16933);
xor U17617 (N_17617,N_16387,N_16038);
xor U17618 (N_17618,N_16422,N_16224);
nor U17619 (N_17619,N_16004,N_16684);
nor U17620 (N_17620,N_16151,N_16907);
or U17621 (N_17621,N_16818,N_16311);
xnor U17622 (N_17622,N_16093,N_16396);
xnor U17623 (N_17623,N_16594,N_16876);
and U17624 (N_17624,N_16389,N_16990);
and U17625 (N_17625,N_16959,N_16886);
xnor U17626 (N_17626,N_16610,N_16662);
nand U17627 (N_17627,N_16035,N_16117);
xor U17628 (N_17628,N_16965,N_16784);
or U17629 (N_17629,N_16111,N_16010);
xnor U17630 (N_17630,N_16082,N_16251);
nand U17631 (N_17631,N_16607,N_16443);
and U17632 (N_17632,N_16941,N_16920);
and U17633 (N_17633,N_16770,N_16593);
nand U17634 (N_17634,N_16302,N_16945);
xnor U17635 (N_17635,N_16172,N_16932);
xnor U17636 (N_17636,N_16527,N_16033);
xor U17637 (N_17637,N_16484,N_16506);
or U17638 (N_17638,N_16400,N_16672);
nor U17639 (N_17639,N_16952,N_16490);
or U17640 (N_17640,N_16996,N_16265);
and U17641 (N_17641,N_16990,N_16435);
and U17642 (N_17642,N_16197,N_16810);
xnor U17643 (N_17643,N_16476,N_16483);
or U17644 (N_17644,N_16207,N_16683);
or U17645 (N_17645,N_16223,N_16916);
or U17646 (N_17646,N_16216,N_16052);
or U17647 (N_17647,N_16869,N_16476);
nor U17648 (N_17648,N_16351,N_16027);
nand U17649 (N_17649,N_16288,N_16834);
and U17650 (N_17650,N_16483,N_16071);
xor U17651 (N_17651,N_16517,N_16521);
or U17652 (N_17652,N_16740,N_16281);
nor U17653 (N_17653,N_16263,N_16828);
and U17654 (N_17654,N_16239,N_16965);
and U17655 (N_17655,N_16426,N_16082);
and U17656 (N_17656,N_16184,N_16726);
xor U17657 (N_17657,N_16526,N_16066);
and U17658 (N_17658,N_16809,N_16114);
and U17659 (N_17659,N_16288,N_16549);
or U17660 (N_17660,N_16705,N_16318);
nand U17661 (N_17661,N_16437,N_16059);
nor U17662 (N_17662,N_16055,N_16710);
xor U17663 (N_17663,N_16007,N_16291);
and U17664 (N_17664,N_16258,N_16040);
and U17665 (N_17665,N_16577,N_16545);
or U17666 (N_17666,N_16834,N_16531);
nor U17667 (N_17667,N_16997,N_16552);
xnor U17668 (N_17668,N_16416,N_16070);
nand U17669 (N_17669,N_16018,N_16535);
xnor U17670 (N_17670,N_16093,N_16590);
or U17671 (N_17671,N_16095,N_16540);
nand U17672 (N_17672,N_16899,N_16166);
and U17673 (N_17673,N_16783,N_16049);
nand U17674 (N_17674,N_16619,N_16195);
nor U17675 (N_17675,N_16870,N_16257);
nor U17676 (N_17676,N_16156,N_16531);
nor U17677 (N_17677,N_16422,N_16898);
xor U17678 (N_17678,N_16958,N_16101);
nand U17679 (N_17679,N_16014,N_16248);
nor U17680 (N_17680,N_16830,N_16928);
nand U17681 (N_17681,N_16812,N_16385);
and U17682 (N_17682,N_16792,N_16565);
xor U17683 (N_17683,N_16734,N_16434);
or U17684 (N_17684,N_16199,N_16564);
nor U17685 (N_17685,N_16707,N_16199);
and U17686 (N_17686,N_16395,N_16073);
nor U17687 (N_17687,N_16452,N_16266);
nand U17688 (N_17688,N_16329,N_16143);
and U17689 (N_17689,N_16860,N_16199);
nor U17690 (N_17690,N_16231,N_16405);
nor U17691 (N_17691,N_16954,N_16060);
nor U17692 (N_17692,N_16927,N_16553);
nand U17693 (N_17693,N_16747,N_16343);
and U17694 (N_17694,N_16037,N_16372);
and U17695 (N_17695,N_16243,N_16743);
nor U17696 (N_17696,N_16810,N_16692);
nand U17697 (N_17697,N_16159,N_16857);
nand U17698 (N_17698,N_16409,N_16614);
nor U17699 (N_17699,N_16515,N_16583);
xnor U17700 (N_17700,N_16597,N_16911);
nor U17701 (N_17701,N_16121,N_16422);
nand U17702 (N_17702,N_16528,N_16938);
and U17703 (N_17703,N_16699,N_16440);
nor U17704 (N_17704,N_16739,N_16491);
and U17705 (N_17705,N_16270,N_16758);
xnor U17706 (N_17706,N_16047,N_16124);
and U17707 (N_17707,N_16592,N_16469);
and U17708 (N_17708,N_16225,N_16888);
nand U17709 (N_17709,N_16105,N_16618);
or U17710 (N_17710,N_16392,N_16541);
or U17711 (N_17711,N_16187,N_16633);
nor U17712 (N_17712,N_16886,N_16387);
xnor U17713 (N_17713,N_16270,N_16386);
nand U17714 (N_17714,N_16386,N_16078);
nand U17715 (N_17715,N_16386,N_16639);
xor U17716 (N_17716,N_16865,N_16630);
xor U17717 (N_17717,N_16520,N_16895);
and U17718 (N_17718,N_16973,N_16041);
and U17719 (N_17719,N_16275,N_16554);
and U17720 (N_17720,N_16337,N_16540);
and U17721 (N_17721,N_16389,N_16197);
nor U17722 (N_17722,N_16278,N_16744);
nand U17723 (N_17723,N_16418,N_16827);
xor U17724 (N_17724,N_16589,N_16995);
nor U17725 (N_17725,N_16511,N_16306);
and U17726 (N_17726,N_16003,N_16357);
or U17727 (N_17727,N_16803,N_16843);
xor U17728 (N_17728,N_16761,N_16855);
xor U17729 (N_17729,N_16059,N_16206);
nor U17730 (N_17730,N_16958,N_16860);
nand U17731 (N_17731,N_16304,N_16276);
and U17732 (N_17732,N_16634,N_16052);
nand U17733 (N_17733,N_16046,N_16540);
and U17734 (N_17734,N_16035,N_16779);
xor U17735 (N_17735,N_16609,N_16236);
and U17736 (N_17736,N_16879,N_16035);
nor U17737 (N_17737,N_16970,N_16752);
nor U17738 (N_17738,N_16028,N_16135);
and U17739 (N_17739,N_16478,N_16786);
xor U17740 (N_17740,N_16784,N_16311);
xor U17741 (N_17741,N_16054,N_16680);
and U17742 (N_17742,N_16458,N_16919);
xor U17743 (N_17743,N_16938,N_16647);
xor U17744 (N_17744,N_16684,N_16031);
nand U17745 (N_17745,N_16425,N_16417);
or U17746 (N_17746,N_16751,N_16339);
nand U17747 (N_17747,N_16320,N_16940);
and U17748 (N_17748,N_16975,N_16227);
or U17749 (N_17749,N_16065,N_16318);
nor U17750 (N_17750,N_16603,N_16721);
nand U17751 (N_17751,N_16286,N_16765);
nor U17752 (N_17752,N_16013,N_16997);
or U17753 (N_17753,N_16666,N_16290);
or U17754 (N_17754,N_16048,N_16425);
and U17755 (N_17755,N_16356,N_16678);
nor U17756 (N_17756,N_16601,N_16906);
and U17757 (N_17757,N_16027,N_16474);
xnor U17758 (N_17758,N_16365,N_16875);
nor U17759 (N_17759,N_16564,N_16436);
and U17760 (N_17760,N_16530,N_16546);
and U17761 (N_17761,N_16822,N_16005);
or U17762 (N_17762,N_16790,N_16359);
nor U17763 (N_17763,N_16291,N_16751);
and U17764 (N_17764,N_16617,N_16682);
and U17765 (N_17765,N_16687,N_16697);
or U17766 (N_17766,N_16939,N_16127);
and U17767 (N_17767,N_16396,N_16363);
nand U17768 (N_17768,N_16952,N_16411);
nand U17769 (N_17769,N_16424,N_16104);
xor U17770 (N_17770,N_16138,N_16761);
or U17771 (N_17771,N_16891,N_16019);
nor U17772 (N_17772,N_16695,N_16843);
nor U17773 (N_17773,N_16273,N_16602);
xor U17774 (N_17774,N_16222,N_16947);
or U17775 (N_17775,N_16150,N_16825);
or U17776 (N_17776,N_16067,N_16294);
or U17777 (N_17777,N_16678,N_16666);
and U17778 (N_17778,N_16136,N_16959);
xor U17779 (N_17779,N_16515,N_16989);
and U17780 (N_17780,N_16328,N_16948);
nor U17781 (N_17781,N_16148,N_16035);
nor U17782 (N_17782,N_16250,N_16753);
nor U17783 (N_17783,N_16909,N_16216);
or U17784 (N_17784,N_16004,N_16074);
nor U17785 (N_17785,N_16406,N_16158);
or U17786 (N_17786,N_16006,N_16473);
nor U17787 (N_17787,N_16220,N_16711);
nand U17788 (N_17788,N_16779,N_16489);
or U17789 (N_17789,N_16300,N_16959);
nor U17790 (N_17790,N_16112,N_16973);
nand U17791 (N_17791,N_16369,N_16877);
nor U17792 (N_17792,N_16613,N_16710);
xnor U17793 (N_17793,N_16999,N_16670);
and U17794 (N_17794,N_16100,N_16781);
nand U17795 (N_17795,N_16974,N_16693);
xor U17796 (N_17796,N_16111,N_16666);
and U17797 (N_17797,N_16394,N_16526);
nand U17798 (N_17798,N_16969,N_16656);
or U17799 (N_17799,N_16261,N_16408);
xnor U17800 (N_17800,N_16774,N_16335);
nor U17801 (N_17801,N_16998,N_16532);
and U17802 (N_17802,N_16404,N_16012);
nor U17803 (N_17803,N_16625,N_16955);
nor U17804 (N_17804,N_16106,N_16492);
or U17805 (N_17805,N_16882,N_16186);
or U17806 (N_17806,N_16290,N_16471);
nand U17807 (N_17807,N_16240,N_16753);
and U17808 (N_17808,N_16085,N_16382);
xor U17809 (N_17809,N_16233,N_16280);
and U17810 (N_17810,N_16234,N_16380);
and U17811 (N_17811,N_16564,N_16472);
and U17812 (N_17812,N_16490,N_16852);
nand U17813 (N_17813,N_16305,N_16135);
or U17814 (N_17814,N_16856,N_16773);
and U17815 (N_17815,N_16263,N_16621);
or U17816 (N_17816,N_16489,N_16600);
or U17817 (N_17817,N_16089,N_16019);
nor U17818 (N_17818,N_16062,N_16882);
xnor U17819 (N_17819,N_16112,N_16066);
nand U17820 (N_17820,N_16757,N_16700);
xnor U17821 (N_17821,N_16835,N_16543);
nand U17822 (N_17822,N_16797,N_16855);
nand U17823 (N_17823,N_16937,N_16253);
nand U17824 (N_17824,N_16528,N_16965);
or U17825 (N_17825,N_16428,N_16052);
xnor U17826 (N_17826,N_16479,N_16939);
xor U17827 (N_17827,N_16819,N_16630);
or U17828 (N_17828,N_16269,N_16843);
or U17829 (N_17829,N_16607,N_16529);
and U17830 (N_17830,N_16587,N_16053);
and U17831 (N_17831,N_16656,N_16028);
xnor U17832 (N_17832,N_16290,N_16421);
nand U17833 (N_17833,N_16911,N_16567);
and U17834 (N_17834,N_16608,N_16972);
and U17835 (N_17835,N_16823,N_16493);
and U17836 (N_17836,N_16142,N_16265);
nand U17837 (N_17837,N_16300,N_16749);
or U17838 (N_17838,N_16687,N_16999);
xor U17839 (N_17839,N_16999,N_16958);
nand U17840 (N_17840,N_16143,N_16947);
xnor U17841 (N_17841,N_16774,N_16942);
and U17842 (N_17842,N_16763,N_16514);
xor U17843 (N_17843,N_16197,N_16085);
nand U17844 (N_17844,N_16613,N_16876);
or U17845 (N_17845,N_16085,N_16703);
or U17846 (N_17846,N_16565,N_16354);
or U17847 (N_17847,N_16619,N_16487);
nand U17848 (N_17848,N_16165,N_16432);
nand U17849 (N_17849,N_16378,N_16486);
nor U17850 (N_17850,N_16993,N_16841);
and U17851 (N_17851,N_16438,N_16506);
nor U17852 (N_17852,N_16179,N_16703);
and U17853 (N_17853,N_16081,N_16671);
nor U17854 (N_17854,N_16993,N_16023);
nor U17855 (N_17855,N_16945,N_16535);
and U17856 (N_17856,N_16523,N_16811);
nor U17857 (N_17857,N_16448,N_16043);
nand U17858 (N_17858,N_16446,N_16254);
nand U17859 (N_17859,N_16984,N_16820);
nand U17860 (N_17860,N_16822,N_16196);
xor U17861 (N_17861,N_16822,N_16073);
nand U17862 (N_17862,N_16224,N_16952);
nand U17863 (N_17863,N_16709,N_16800);
or U17864 (N_17864,N_16917,N_16464);
nand U17865 (N_17865,N_16153,N_16371);
xnor U17866 (N_17866,N_16608,N_16875);
and U17867 (N_17867,N_16947,N_16734);
nand U17868 (N_17868,N_16521,N_16853);
or U17869 (N_17869,N_16115,N_16796);
nand U17870 (N_17870,N_16126,N_16269);
nor U17871 (N_17871,N_16544,N_16415);
nor U17872 (N_17872,N_16100,N_16467);
and U17873 (N_17873,N_16876,N_16437);
or U17874 (N_17874,N_16589,N_16023);
or U17875 (N_17875,N_16143,N_16229);
xor U17876 (N_17876,N_16375,N_16189);
nand U17877 (N_17877,N_16718,N_16861);
nand U17878 (N_17878,N_16597,N_16079);
nor U17879 (N_17879,N_16060,N_16999);
and U17880 (N_17880,N_16314,N_16257);
nor U17881 (N_17881,N_16848,N_16314);
nand U17882 (N_17882,N_16585,N_16973);
nor U17883 (N_17883,N_16725,N_16534);
nand U17884 (N_17884,N_16257,N_16928);
nor U17885 (N_17885,N_16257,N_16566);
nor U17886 (N_17886,N_16072,N_16278);
nor U17887 (N_17887,N_16275,N_16045);
and U17888 (N_17888,N_16468,N_16971);
nand U17889 (N_17889,N_16534,N_16113);
xnor U17890 (N_17890,N_16464,N_16868);
nand U17891 (N_17891,N_16207,N_16243);
xor U17892 (N_17892,N_16086,N_16842);
xor U17893 (N_17893,N_16580,N_16260);
or U17894 (N_17894,N_16332,N_16294);
nor U17895 (N_17895,N_16655,N_16032);
or U17896 (N_17896,N_16275,N_16377);
nand U17897 (N_17897,N_16395,N_16014);
or U17898 (N_17898,N_16603,N_16290);
nand U17899 (N_17899,N_16542,N_16638);
and U17900 (N_17900,N_16311,N_16980);
or U17901 (N_17901,N_16263,N_16479);
xnor U17902 (N_17902,N_16775,N_16079);
nand U17903 (N_17903,N_16051,N_16727);
nand U17904 (N_17904,N_16008,N_16536);
nand U17905 (N_17905,N_16912,N_16098);
xnor U17906 (N_17906,N_16203,N_16213);
or U17907 (N_17907,N_16169,N_16764);
nor U17908 (N_17908,N_16900,N_16903);
and U17909 (N_17909,N_16212,N_16740);
or U17910 (N_17910,N_16572,N_16613);
or U17911 (N_17911,N_16835,N_16349);
and U17912 (N_17912,N_16652,N_16803);
nand U17913 (N_17913,N_16334,N_16279);
or U17914 (N_17914,N_16518,N_16364);
nor U17915 (N_17915,N_16723,N_16160);
and U17916 (N_17916,N_16600,N_16090);
nor U17917 (N_17917,N_16024,N_16141);
nor U17918 (N_17918,N_16010,N_16721);
nand U17919 (N_17919,N_16250,N_16076);
and U17920 (N_17920,N_16890,N_16419);
nor U17921 (N_17921,N_16667,N_16044);
nor U17922 (N_17922,N_16455,N_16419);
xor U17923 (N_17923,N_16002,N_16070);
nor U17924 (N_17924,N_16672,N_16708);
and U17925 (N_17925,N_16843,N_16159);
and U17926 (N_17926,N_16298,N_16956);
or U17927 (N_17927,N_16815,N_16039);
nor U17928 (N_17928,N_16941,N_16408);
or U17929 (N_17929,N_16373,N_16564);
xnor U17930 (N_17930,N_16351,N_16048);
xor U17931 (N_17931,N_16555,N_16369);
xor U17932 (N_17932,N_16248,N_16445);
and U17933 (N_17933,N_16274,N_16648);
xnor U17934 (N_17934,N_16638,N_16696);
and U17935 (N_17935,N_16500,N_16618);
and U17936 (N_17936,N_16491,N_16678);
nor U17937 (N_17937,N_16342,N_16984);
and U17938 (N_17938,N_16400,N_16131);
nand U17939 (N_17939,N_16251,N_16037);
nor U17940 (N_17940,N_16587,N_16279);
and U17941 (N_17941,N_16175,N_16655);
nor U17942 (N_17942,N_16920,N_16927);
xnor U17943 (N_17943,N_16681,N_16858);
and U17944 (N_17944,N_16017,N_16701);
and U17945 (N_17945,N_16229,N_16170);
nor U17946 (N_17946,N_16798,N_16825);
nand U17947 (N_17947,N_16091,N_16867);
and U17948 (N_17948,N_16755,N_16939);
or U17949 (N_17949,N_16862,N_16202);
and U17950 (N_17950,N_16683,N_16762);
nand U17951 (N_17951,N_16625,N_16918);
nor U17952 (N_17952,N_16700,N_16755);
nor U17953 (N_17953,N_16382,N_16043);
nor U17954 (N_17954,N_16484,N_16099);
nand U17955 (N_17955,N_16694,N_16846);
xor U17956 (N_17956,N_16216,N_16444);
nand U17957 (N_17957,N_16272,N_16134);
nand U17958 (N_17958,N_16254,N_16758);
and U17959 (N_17959,N_16796,N_16012);
xnor U17960 (N_17960,N_16195,N_16841);
nand U17961 (N_17961,N_16802,N_16484);
nor U17962 (N_17962,N_16384,N_16702);
xor U17963 (N_17963,N_16719,N_16305);
nand U17964 (N_17964,N_16237,N_16503);
or U17965 (N_17965,N_16021,N_16981);
xor U17966 (N_17966,N_16806,N_16504);
xor U17967 (N_17967,N_16976,N_16900);
or U17968 (N_17968,N_16951,N_16841);
nand U17969 (N_17969,N_16397,N_16561);
nor U17970 (N_17970,N_16642,N_16445);
xor U17971 (N_17971,N_16675,N_16808);
or U17972 (N_17972,N_16537,N_16402);
and U17973 (N_17973,N_16395,N_16658);
or U17974 (N_17974,N_16610,N_16616);
nand U17975 (N_17975,N_16439,N_16694);
xor U17976 (N_17976,N_16879,N_16319);
or U17977 (N_17977,N_16580,N_16046);
nor U17978 (N_17978,N_16137,N_16885);
nand U17979 (N_17979,N_16252,N_16398);
nor U17980 (N_17980,N_16222,N_16864);
nand U17981 (N_17981,N_16404,N_16803);
or U17982 (N_17982,N_16770,N_16747);
and U17983 (N_17983,N_16464,N_16793);
nand U17984 (N_17984,N_16625,N_16768);
and U17985 (N_17985,N_16949,N_16656);
xor U17986 (N_17986,N_16306,N_16694);
nand U17987 (N_17987,N_16521,N_16973);
xnor U17988 (N_17988,N_16320,N_16125);
xor U17989 (N_17989,N_16502,N_16321);
xor U17990 (N_17990,N_16498,N_16727);
or U17991 (N_17991,N_16026,N_16688);
xnor U17992 (N_17992,N_16512,N_16274);
nand U17993 (N_17993,N_16788,N_16978);
and U17994 (N_17994,N_16820,N_16949);
nor U17995 (N_17995,N_16195,N_16361);
and U17996 (N_17996,N_16291,N_16188);
and U17997 (N_17997,N_16387,N_16808);
or U17998 (N_17998,N_16188,N_16557);
nor U17999 (N_17999,N_16052,N_16077);
or U18000 (N_18000,N_17116,N_17612);
nand U18001 (N_18001,N_17954,N_17328);
nand U18002 (N_18002,N_17296,N_17835);
nor U18003 (N_18003,N_17550,N_17971);
nand U18004 (N_18004,N_17016,N_17360);
nand U18005 (N_18005,N_17912,N_17668);
and U18006 (N_18006,N_17739,N_17066);
nor U18007 (N_18007,N_17135,N_17243);
nand U18008 (N_18008,N_17123,N_17485);
and U18009 (N_18009,N_17888,N_17103);
or U18010 (N_18010,N_17689,N_17295);
or U18011 (N_18011,N_17254,N_17958);
nor U18012 (N_18012,N_17967,N_17253);
xor U18013 (N_18013,N_17705,N_17868);
or U18014 (N_18014,N_17655,N_17547);
nand U18015 (N_18015,N_17068,N_17911);
xor U18016 (N_18016,N_17285,N_17316);
nand U18017 (N_18017,N_17884,N_17021);
nand U18018 (N_18018,N_17206,N_17466);
xor U18019 (N_18019,N_17190,N_17162);
and U18020 (N_18020,N_17684,N_17405);
and U18021 (N_18021,N_17771,N_17386);
xor U18022 (N_18022,N_17286,N_17957);
or U18023 (N_18023,N_17460,N_17783);
xor U18024 (N_18024,N_17026,N_17311);
or U18025 (N_18025,N_17453,N_17422);
and U18026 (N_18026,N_17304,N_17011);
nand U18027 (N_18027,N_17604,N_17455);
and U18028 (N_18028,N_17701,N_17621);
nor U18029 (N_18029,N_17831,N_17279);
nor U18030 (N_18030,N_17309,N_17504);
xor U18031 (N_18031,N_17688,N_17737);
xor U18032 (N_18032,N_17534,N_17139);
nor U18033 (N_18033,N_17980,N_17978);
xnor U18034 (N_18034,N_17015,N_17115);
xnor U18035 (N_18035,N_17355,N_17467);
xnor U18036 (N_18036,N_17923,N_17763);
xnor U18037 (N_18037,N_17395,N_17002);
or U18038 (N_18038,N_17663,N_17171);
nor U18039 (N_18039,N_17693,N_17306);
nand U18040 (N_18040,N_17438,N_17833);
nor U18041 (N_18041,N_17148,N_17132);
nand U18042 (N_18042,N_17137,N_17027);
nor U18043 (N_18043,N_17210,N_17671);
nand U18044 (N_18044,N_17380,N_17756);
nand U18045 (N_18045,N_17432,N_17987);
xor U18046 (N_18046,N_17562,N_17617);
or U18047 (N_18047,N_17326,N_17824);
xor U18048 (N_18048,N_17303,N_17790);
xor U18049 (N_18049,N_17310,N_17155);
xnor U18050 (N_18050,N_17752,N_17322);
nor U18051 (N_18051,N_17158,N_17567);
and U18052 (N_18052,N_17594,N_17998);
or U18053 (N_18053,N_17102,N_17493);
or U18054 (N_18054,N_17964,N_17968);
and U18055 (N_18055,N_17639,N_17633);
nand U18056 (N_18056,N_17029,N_17289);
nand U18057 (N_18057,N_17513,N_17876);
or U18058 (N_18058,N_17004,N_17863);
or U18059 (N_18059,N_17544,N_17898);
and U18060 (N_18060,N_17675,N_17627);
or U18061 (N_18061,N_17110,N_17268);
nor U18062 (N_18062,N_17409,N_17895);
xnor U18063 (N_18063,N_17425,N_17629);
nor U18064 (N_18064,N_17064,N_17271);
xnor U18065 (N_18065,N_17174,N_17529);
or U18066 (N_18066,N_17691,N_17489);
or U18067 (N_18067,N_17151,N_17204);
nor U18068 (N_18068,N_17855,N_17554);
or U18069 (N_18069,N_17112,N_17682);
nand U18070 (N_18070,N_17336,N_17556);
or U18071 (N_18071,N_17757,N_17664);
nand U18072 (N_18072,N_17749,N_17194);
xnor U18073 (N_18073,N_17244,N_17878);
nor U18074 (N_18074,N_17973,N_17219);
or U18075 (N_18075,N_17651,N_17284);
xnor U18076 (N_18076,N_17372,N_17085);
nand U18077 (N_18077,N_17804,N_17665);
xor U18078 (N_18078,N_17062,N_17972);
and U18079 (N_18079,N_17381,N_17732);
nor U18080 (N_18080,N_17090,N_17871);
and U18081 (N_18081,N_17505,N_17839);
and U18082 (N_18082,N_17560,N_17748);
nor U18083 (N_18083,N_17055,N_17608);
nand U18084 (N_18084,N_17374,N_17974);
or U18085 (N_18085,N_17492,N_17041);
nand U18086 (N_18086,N_17030,N_17514);
or U18087 (N_18087,N_17028,N_17789);
and U18088 (N_18088,N_17905,N_17107);
or U18089 (N_18089,N_17775,N_17557);
xor U18090 (N_18090,N_17497,N_17673);
or U18091 (N_18091,N_17001,N_17901);
or U18092 (N_18092,N_17262,N_17251);
nand U18093 (N_18093,N_17843,N_17018);
nand U18094 (N_18094,N_17654,N_17945);
and U18095 (N_18095,N_17765,N_17942);
or U18096 (N_18096,N_17357,N_17081);
nor U18097 (N_18097,N_17502,N_17390);
nor U18098 (N_18098,N_17379,N_17653);
or U18099 (N_18099,N_17335,N_17480);
or U18100 (N_18100,N_17862,N_17152);
xnor U18101 (N_18101,N_17844,N_17010);
or U18102 (N_18102,N_17203,N_17334);
xor U18103 (N_18103,N_17387,N_17166);
and U18104 (N_18104,N_17549,N_17017);
nor U18105 (N_18105,N_17005,N_17879);
xnor U18106 (N_18106,N_17385,N_17722);
and U18107 (N_18107,N_17988,N_17614);
nor U18108 (N_18108,N_17875,N_17074);
or U18109 (N_18109,N_17444,N_17404);
nand U18110 (N_18110,N_17412,N_17872);
nor U18111 (N_18111,N_17788,N_17350);
nor U18112 (N_18112,N_17128,N_17590);
or U18113 (N_18113,N_17431,N_17161);
and U18114 (N_18114,N_17578,N_17511);
nor U18115 (N_18115,N_17223,N_17235);
nor U18116 (N_18116,N_17365,N_17642);
xor U18117 (N_18117,N_17240,N_17234);
and U18118 (N_18118,N_17414,N_17776);
and U18119 (N_18119,N_17450,N_17220);
or U18120 (N_18120,N_17817,N_17777);
nand U18121 (N_18121,N_17167,N_17353);
nor U18122 (N_18122,N_17506,N_17288);
or U18123 (N_18123,N_17227,N_17424);
xnor U18124 (N_18124,N_17138,N_17532);
nor U18125 (N_18125,N_17212,N_17451);
or U18126 (N_18126,N_17163,N_17834);
xor U18127 (N_18127,N_17782,N_17870);
xnor U18128 (N_18128,N_17827,N_17293);
nor U18129 (N_18129,N_17358,N_17057);
or U18130 (N_18130,N_17142,N_17091);
or U18131 (N_18131,N_17180,N_17826);
nor U18132 (N_18132,N_17221,N_17156);
nand U18133 (N_18133,N_17486,N_17263);
xnor U18134 (N_18134,N_17815,N_17426);
xnor U18135 (N_18135,N_17904,N_17430);
nand U18136 (N_18136,N_17478,N_17956);
nand U18137 (N_18137,N_17986,N_17040);
or U18138 (N_18138,N_17000,N_17969);
nand U18139 (N_18139,N_17553,N_17452);
and U18140 (N_18140,N_17393,N_17126);
xor U18141 (N_18141,N_17264,N_17809);
nor U18142 (N_18142,N_17766,N_17046);
xor U18143 (N_18143,N_17743,N_17267);
nand U18144 (N_18144,N_17299,N_17742);
or U18145 (N_18145,N_17545,N_17519);
nand U18146 (N_18146,N_17507,N_17169);
and U18147 (N_18147,N_17145,N_17172);
or U18148 (N_18148,N_17441,N_17370);
and U18149 (N_18149,N_17571,N_17265);
nor U18150 (N_18150,N_17908,N_17022);
or U18151 (N_18151,N_17178,N_17146);
or U18152 (N_18152,N_17993,N_17242);
xnor U18153 (N_18153,N_17119,N_17900);
and U18154 (N_18154,N_17320,N_17858);
or U18155 (N_18155,N_17952,N_17736);
xnor U18156 (N_18156,N_17063,N_17628);
xnor U18157 (N_18157,N_17187,N_17710);
or U18158 (N_18158,N_17061,N_17930);
xnor U18159 (N_18159,N_17587,N_17352);
nor U18160 (N_18160,N_17052,N_17764);
and U18161 (N_18161,N_17185,N_17925);
or U18162 (N_18162,N_17601,N_17417);
nand U18163 (N_18163,N_17546,N_17369);
and U18164 (N_18164,N_17857,N_17821);
nand U18165 (N_18165,N_17927,N_17241);
xor U18166 (N_18166,N_17965,N_17232);
xnor U18167 (N_18167,N_17491,N_17106);
nand U18168 (N_18168,N_17727,N_17347);
or U18169 (N_18169,N_17769,N_17421);
xnor U18170 (N_18170,N_17854,N_17632);
and U18171 (N_18171,N_17012,N_17464);
nor U18172 (N_18172,N_17881,N_17373);
or U18173 (N_18173,N_17596,N_17818);
xnor U18174 (N_18174,N_17315,N_17044);
nand U18175 (N_18175,N_17468,N_17979);
nor U18176 (N_18176,N_17256,N_17585);
nor U18177 (N_18177,N_17449,N_17798);
xor U18178 (N_18178,N_17848,N_17456);
nand U18179 (N_18179,N_17894,N_17032);
nor U18180 (N_18180,N_17861,N_17282);
xor U18181 (N_18181,N_17448,N_17056);
nand U18182 (N_18182,N_17877,N_17067);
nand U18183 (N_18183,N_17494,N_17570);
xnor U18184 (N_18184,N_17740,N_17312);
nor U18185 (N_18185,N_17410,N_17255);
and U18186 (N_18186,N_17995,N_17209);
or U18187 (N_18187,N_17428,N_17362);
nor U18188 (N_18188,N_17569,N_17563);
xor U18189 (N_18189,N_17860,N_17591);
and U18190 (N_18190,N_17233,N_17774);
xor U18191 (N_18191,N_17198,N_17709);
or U18192 (N_18192,N_17528,N_17784);
nor U18193 (N_18193,N_17940,N_17555);
and U18194 (N_18194,N_17989,N_17400);
nor U18195 (N_18195,N_17699,N_17222);
and U18196 (N_18196,N_17572,N_17313);
or U18197 (N_18197,N_17048,N_17593);
or U18198 (N_18198,N_17082,N_17565);
or U18199 (N_18199,N_17586,N_17100);
and U18200 (N_18200,N_17683,N_17948);
xnor U18201 (N_18201,N_17348,N_17401);
or U18202 (N_18202,N_17919,N_17333);
nor U18203 (N_18203,N_17666,N_17245);
or U18204 (N_18204,N_17298,N_17674);
and U18205 (N_18205,N_17483,N_17893);
or U18206 (N_18206,N_17238,N_17340);
nand U18207 (N_18207,N_17823,N_17733);
nor U18208 (N_18208,N_17626,N_17484);
or U18209 (N_18209,N_17907,N_17439);
xor U18210 (N_18210,N_17805,N_17630);
and U18211 (N_18211,N_17548,N_17584);
and U18212 (N_18212,N_17523,N_17734);
xnor U18213 (N_18213,N_17407,N_17435);
or U18214 (N_18214,N_17867,N_17076);
nand U18215 (N_18215,N_17196,N_17924);
nor U18216 (N_18216,N_17885,N_17897);
xor U18217 (N_18217,N_17157,N_17475);
nor U18218 (N_18218,N_17595,N_17273);
and U18219 (N_18219,N_17257,N_17915);
and U18220 (N_18220,N_17199,N_17249);
or U18221 (N_18221,N_17516,N_17853);
nor U18222 (N_18222,N_17324,N_17966);
xnor U18223 (N_18223,N_17738,N_17800);
nand U18224 (N_18224,N_17944,N_17625);
and U18225 (N_18225,N_17208,N_17521);
xor U18226 (N_18226,N_17133,N_17501);
nor U18227 (N_18227,N_17276,N_17050);
or U18228 (N_18228,N_17711,N_17721);
xor U18229 (N_18229,N_17088,N_17291);
nor U18230 (N_18230,N_17399,N_17811);
nand U18231 (N_18231,N_17496,N_17136);
xnor U18232 (N_18232,N_17213,N_17247);
nand U18233 (N_18233,N_17205,N_17419);
nor U18234 (N_18234,N_17896,N_17454);
or U18235 (N_18235,N_17660,N_17903);
xor U18236 (N_18236,N_17105,N_17606);
nand U18237 (N_18237,N_17624,N_17246);
nor U18238 (N_18238,N_17436,N_17325);
and U18239 (N_18239,N_17101,N_17075);
xor U18240 (N_18240,N_17389,N_17820);
and U18241 (N_18241,N_17724,N_17281);
nand U18242 (N_18242,N_17184,N_17640);
nor U18243 (N_18243,N_17008,N_17648);
and U18244 (N_18244,N_17023,N_17943);
or U18245 (N_18245,N_17471,N_17195);
xor U18246 (N_18246,N_17723,N_17356);
or U18247 (N_18247,N_17706,N_17149);
nor U18248 (N_18248,N_17164,N_17343);
nor U18249 (N_18249,N_17941,N_17846);
and U18250 (N_18250,N_17394,N_17672);
and U18251 (N_18251,N_17269,N_17397);
and U18252 (N_18252,N_17165,N_17230);
or U18253 (N_18253,N_17891,N_17602);
and U18254 (N_18254,N_17482,N_17787);
and U18255 (N_18255,N_17495,N_17909);
and U18256 (N_18256,N_17170,N_17802);
and U18257 (N_18257,N_17917,N_17791);
or U18258 (N_18258,N_17715,N_17535);
or U18259 (N_18259,N_17186,N_17037);
or U18260 (N_18260,N_17479,N_17473);
nor U18261 (N_18261,N_17702,N_17814);
xor U18262 (N_18262,N_17677,N_17889);
nand U18263 (N_18263,N_17508,N_17990);
nand U18264 (N_18264,N_17582,N_17260);
and U18265 (N_18265,N_17098,N_17321);
nor U18266 (N_18266,N_17551,N_17690);
xor U18267 (N_18267,N_17134,N_17836);
or U18268 (N_18268,N_17961,N_17197);
and U18269 (N_18269,N_17543,N_17476);
or U18270 (N_18270,N_17936,N_17982);
and U18271 (N_18271,N_17792,N_17914);
xnor U18272 (N_18272,N_17842,N_17883);
nor U18273 (N_18273,N_17713,N_17697);
and U18274 (N_18274,N_17175,N_17457);
or U18275 (N_18275,N_17994,N_17498);
or U18276 (N_18276,N_17647,N_17955);
nor U18277 (N_18277,N_17735,N_17490);
xnor U18278 (N_18278,N_17122,N_17488);
or U18279 (N_18279,N_17038,N_17160);
or U18280 (N_18280,N_17616,N_17211);
xor U18281 (N_18281,N_17034,N_17750);
xor U18282 (N_18282,N_17499,N_17121);
or U18283 (N_18283,N_17459,N_17662);
xnor U18284 (N_18284,N_17089,N_17573);
or U18285 (N_18285,N_17079,N_17849);
nand U18286 (N_18286,N_17415,N_17345);
nor U18287 (N_18287,N_17856,N_17806);
nand U18288 (N_18288,N_17359,N_17314);
and U18289 (N_18289,N_17111,N_17947);
nor U18290 (N_18290,N_17880,N_17692);
or U18291 (N_18291,N_17047,N_17985);
xor U18292 (N_18292,N_17418,N_17083);
and U18293 (N_18293,N_17442,N_17780);
xnor U18294 (N_18294,N_17200,N_17997);
xnor U18295 (N_18295,N_17841,N_17916);
xnor U18296 (N_18296,N_17719,N_17959);
nand U18297 (N_18297,N_17413,N_17071);
and U18298 (N_18298,N_17618,N_17224);
xor U18299 (N_18299,N_17741,N_17698);
and U18300 (N_18300,N_17851,N_17762);
nor U18301 (N_18301,N_17579,N_17920);
xnor U18302 (N_18302,N_17013,N_17058);
or U18303 (N_18303,N_17770,N_17746);
nand U18304 (N_18304,N_17822,N_17096);
and U18305 (N_18305,N_17368,N_17793);
nand U18306 (N_18306,N_17622,N_17109);
xnor U18307 (N_18307,N_17694,N_17500);
and U18308 (N_18308,N_17963,N_17613);
nor U18309 (N_18309,N_17686,N_17619);
nor U18310 (N_18310,N_17087,N_17445);
nor U18311 (N_18311,N_17576,N_17751);
or U18312 (N_18312,N_17785,N_17275);
and U18313 (N_18313,N_17019,N_17667);
nand U18314 (N_18314,N_17077,N_17643);
nand U18315 (N_18315,N_17847,N_17669);
nor U18316 (N_18316,N_17049,N_17641);
and U18317 (N_18317,N_17351,N_17716);
nor U18318 (N_18318,N_17065,N_17656);
nand U18319 (N_18319,N_17635,N_17154);
nor U18320 (N_18320,N_17946,N_17939);
nor U18321 (N_18321,N_17129,N_17150);
nor U18322 (N_18322,N_17294,N_17465);
and U18323 (N_18323,N_17589,N_17527);
and U18324 (N_18324,N_17364,N_17583);
nor U18325 (N_18325,N_17599,N_17533);
nand U18326 (N_18326,N_17192,N_17302);
and U18327 (N_18327,N_17918,N_17531);
nand U18328 (N_18328,N_17657,N_17097);
and U18329 (N_18329,N_17886,N_17039);
nor U18330 (N_18330,N_17007,N_17773);
nand U18331 (N_18331,N_17960,N_17929);
and U18332 (N_18332,N_17095,N_17252);
or U18333 (N_18333,N_17280,N_17910);
nor U18334 (N_18334,N_17346,N_17761);
xor U18335 (N_18335,N_17976,N_17443);
nor U18336 (N_18336,N_17215,N_17932);
xor U18337 (N_18337,N_17104,N_17283);
nor U18338 (N_18338,N_17634,N_17859);
and U18339 (N_18339,N_17564,N_17094);
nor U18340 (N_18340,N_17708,N_17024);
and U18341 (N_18341,N_17006,N_17829);
nor U18342 (N_18342,N_17922,N_17795);
nor U18343 (N_18343,N_17339,N_17864);
nor U18344 (N_18344,N_17411,N_17687);
xnor U18345 (N_18345,N_17403,N_17600);
nand U18346 (N_18346,N_17631,N_17638);
xnor U18347 (N_18347,N_17779,N_17678);
xor U18348 (N_18348,N_17649,N_17539);
nand U18349 (N_18349,N_17882,N_17680);
or U18350 (N_18350,N_17093,N_17045);
xnor U18351 (N_18351,N_17926,N_17537);
or U18352 (N_18352,N_17383,N_17873);
xnor U18353 (N_18353,N_17266,N_17825);
nand U18354 (N_18354,N_17290,N_17540);
nand U18355 (N_18355,N_17679,N_17031);
and U18356 (N_18356,N_17819,N_17226);
nand U18357 (N_18357,N_17130,N_17392);
or U18358 (N_18358,N_17838,N_17588);
or U18359 (N_18359,N_17182,N_17278);
or U18360 (N_18360,N_17366,N_17561);
nor U18361 (N_18361,N_17509,N_17518);
xor U18362 (N_18362,N_17938,N_17704);
xnor U18363 (N_18363,N_17297,N_17636);
nand U18364 (N_18364,N_17461,N_17272);
nor U18365 (N_18365,N_17033,N_17906);
nand U18366 (N_18366,N_17218,N_17510);
and U18367 (N_18367,N_17072,N_17141);
or U18368 (N_18368,N_17832,N_17440);
xnor U18369 (N_18369,N_17469,N_17623);
nor U18370 (N_18370,N_17183,N_17931);
or U18371 (N_18371,N_17341,N_17522);
nor U18372 (N_18372,N_17707,N_17610);
nor U18373 (N_18373,N_17217,N_17808);
xnor U18374 (N_18374,N_17597,N_17114);
and U18375 (N_18375,N_17147,N_17384);
nor U18376 (N_18376,N_17338,N_17928);
nand U18377 (N_18377,N_17670,N_17755);
nor U18378 (N_18378,N_17250,N_17201);
nor U18379 (N_18379,N_17899,N_17977);
nor U18380 (N_18380,N_17080,N_17685);
xor U18381 (N_18381,N_17934,N_17237);
nor U18382 (N_18382,N_17845,N_17301);
and U18383 (N_18383,N_17396,N_17813);
nand U18384 (N_18384,N_17463,N_17801);
and U18385 (N_18385,N_17951,N_17287);
nand U18386 (N_18386,N_17371,N_17503);
xnor U18387 (N_18387,N_17159,N_17828);
and U18388 (N_18388,N_17053,N_17117);
nand U18389 (N_18389,N_17458,N_17377);
nand U18390 (N_18390,N_17131,N_17520);
nor U18391 (N_18391,N_17307,N_17542);
nor U18392 (N_18392,N_17429,N_17344);
xnor U18393 (N_18393,N_17330,N_17308);
and U18394 (N_18394,N_17574,N_17474);
or U18395 (N_18395,N_17176,N_17331);
xor U18396 (N_18396,N_17446,N_17258);
xnor U18397 (N_18397,N_17376,N_17481);
or U18398 (N_18398,N_17420,N_17652);
and U18399 (N_18399,N_17092,N_17318);
nor U18400 (N_18400,N_17730,N_17953);
and U18401 (N_18401,N_17659,N_17402);
xor U18402 (N_18402,N_17069,N_17866);
or U18403 (N_18403,N_17717,N_17536);
xor U18404 (N_18404,N_17332,N_17337);
nand U18405 (N_18405,N_17433,N_17729);
nor U18406 (N_18406,N_17714,N_17799);
or U18407 (N_18407,N_17720,N_17996);
or U18408 (N_18408,N_17611,N_17984);
nand U18409 (N_18409,N_17173,N_17270);
or U18410 (N_18410,N_17970,N_17645);
or U18411 (N_18411,N_17681,N_17487);
or U18412 (N_18412,N_17292,N_17051);
nand U18413 (N_18413,N_17837,N_17768);
xor U18414 (N_18414,N_17869,N_17525);
nor U18415 (N_18415,N_17323,N_17259);
nor U18416 (N_18416,N_17181,N_17042);
nor U18417 (N_18417,N_17615,N_17300);
xnor U18418 (N_18418,N_17388,N_17526);
or U18419 (N_18419,N_17517,N_17744);
nor U18420 (N_18420,N_17747,N_17981);
xor U18421 (N_18421,N_17225,N_17228);
nor U18422 (N_18422,N_17598,N_17999);
nand U18423 (N_18423,N_17797,N_17812);
nor U18424 (N_18424,N_17472,N_17363);
xor U18425 (N_18425,N_17070,N_17575);
and U18426 (N_18426,N_17124,N_17512);
nand U18427 (N_18427,N_17462,N_17609);
xor U18428 (N_18428,N_17696,N_17317);
nand U18429 (N_18429,N_17661,N_17605);
nand U18430 (N_18430,N_17153,N_17214);
or U18431 (N_18431,N_17580,N_17207);
xor U18432 (N_18432,N_17767,N_17753);
and U18433 (N_18433,N_17025,N_17718);
nand U18434 (N_18434,N_17786,N_17035);
nor U18435 (N_18435,N_17437,N_17108);
nor U18436 (N_18436,N_17423,N_17188);
or U18437 (N_18437,N_17329,N_17731);
nor U18438 (N_18438,N_17398,N_17796);
and U18439 (N_18439,N_17231,N_17607);
and U18440 (N_18440,N_17014,N_17391);
and U18441 (N_18441,N_17375,N_17541);
and U18442 (N_18442,N_17378,N_17118);
xor U18443 (N_18443,N_17202,N_17020);
nand U18444 (N_18444,N_17887,N_17676);
nor U18445 (N_18445,N_17191,N_17216);
or U18446 (N_18446,N_17754,N_17725);
or U18447 (N_18447,N_17319,N_17892);
or U18448 (N_18448,N_17874,N_17229);
nor U18449 (N_18449,N_17760,N_17143);
and U18450 (N_18450,N_17515,N_17361);
nand U18451 (N_18451,N_17530,N_17470);
and U18452 (N_18452,N_17447,N_17658);
and U18453 (N_18453,N_17581,N_17646);
nand U18454 (N_18454,N_17902,N_17703);
nor U18455 (N_18455,N_17477,N_17239);
xor U18456 (N_18456,N_17758,N_17305);
xor U18457 (N_18457,N_17695,N_17078);
nor U18458 (N_18458,N_17248,N_17277);
nor U18459 (N_18459,N_17794,N_17524);
or U18460 (N_18460,N_17059,N_17084);
nand U18461 (N_18461,N_17538,N_17193);
and U18462 (N_18462,N_17342,N_17558);
or U18463 (N_18463,N_17803,N_17644);
nor U18464 (N_18464,N_17168,N_17382);
nand U18465 (N_18465,N_17772,N_17850);
xnor U18466 (N_18466,N_17852,N_17086);
or U18467 (N_18467,N_17144,N_17726);
nor U18468 (N_18468,N_17434,N_17810);
nor U18469 (N_18469,N_17933,N_17349);
or U18470 (N_18470,N_17113,N_17950);
and U18471 (N_18471,N_17603,N_17043);
and U18472 (N_18472,N_17983,N_17949);
nor U18473 (N_18473,N_17427,N_17620);
nand U18474 (N_18474,N_17921,N_17759);
xor U18475 (N_18475,N_17189,N_17728);
and U18476 (N_18476,N_17781,N_17778);
nor U18477 (N_18477,N_17592,N_17962);
nor U18478 (N_18478,N_17036,N_17816);
or U18479 (N_18479,N_17650,N_17073);
nand U18480 (N_18480,N_17807,N_17568);
or U18481 (N_18481,N_17865,N_17261);
and U18482 (N_18482,N_17120,N_17992);
or U18483 (N_18483,N_17003,N_17179);
nand U18484 (N_18484,N_17416,N_17712);
nand U18485 (N_18485,N_17913,N_17099);
xor U18486 (N_18486,N_17552,N_17406);
and U18487 (N_18487,N_17700,N_17054);
nand U18488 (N_18488,N_17559,N_17577);
nor U18489 (N_18489,N_17274,N_17935);
nor U18490 (N_18490,N_17127,N_17840);
nor U18491 (N_18491,N_17140,N_17060);
and U18492 (N_18492,N_17890,N_17177);
nor U18493 (N_18493,N_17637,N_17566);
nor U18494 (N_18494,N_17367,N_17745);
and U18495 (N_18495,N_17991,N_17009);
xor U18496 (N_18496,N_17125,N_17408);
and U18497 (N_18497,N_17236,N_17937);
or U18498 (N_18498,N_17975,N_17327);
nand U18499 (N_18499,N_17830,N_17354);
nand U18500 (N_18500,N_17437,N_17575);
xor U18501 (N_18501,N_17993,N_17450);
xor U18502 (N_18502,N_17157,N_17211);
xor U18503 (N_18503,N_17360,N_17364);
or U18504 (N_18504,N_17792,N_17374);
xor U18505 (N_18505,N_17569,N_17425);
and U18506 (N_18506,N_17505,N_17942);
nand U18507 (N_18507,N_17871,N_17281);
or U18508 (N_18508,N_17762,N_17779);
or U18509 (N_18509,N_17585,N_17677);
nand U18510 (N_18510,N_17146,N_17666);
or U18511 (N_18511,N_17131,N_17985);
and U18512 (N_18512,N_17075,N_17799);
xor U18513 (N_18513,N_17505,N_17864);
and U18514 (N_18514,N_17058,N_17060);
nand U18515 (N_18515,N_17435,N_17989);
nor U18516 (N_18516,N_17530,N_17514);
and U18517 (N_18517,N_17793,N_17680);
or U18518 (N_18518,N_17080,N_17276);
nand U18519 (N_18519,N_17053,N_17894);
nand U18520 (N_18520,N_17307,N_17406);
and U18521 (N_18521,N_17107,N_17146);
xnor U18522 (N_18522,N_17501,N_17157);
and U18523 (N_18523,N_17888,N_17185);
nand U18524 (N_18524,N_17925,N_17608);
xor U18525 (N_18525,N_17361,N_17313);
xnor U18526 (N_18526,N_17252,N_17186);
nor U18527 (N_18527,N_17715,N_17091);
xnor U18528 (N_18528,N_17843,N_17498);
nor U18529 (N_18529,N_17795,N_17589);
xnor U18530 (N_18530,N_17976,N_17822);
or U18531 (N_18531,N_17260,N_17884);
nor U18532 (N_18532,N_17238,N_17505);
nand U18533 (N_18533,N_17140,N_17402);
and U18534 (N_18534,N_17313,N_17899);
nor U18535 (N_18535,N_17518,N_17876);
nor U18536 (N_18536,N_17866,N_17253);
nor U18537 (N_18537,N_17152,N_17204);
and U18538 (N_18538,N_17682,N_17612);
and U18539 (N_18539,N_17375,N_17185);
nand U18540 (N_18540,N_17573,N_17007);
and U18541 (N_18541,N_17318,N_17451);
nand U18542 (N_18542,N_17478,N_17233);
nand U18543 (N_18543,N_17254,N_17508);
nand U18544 (N_18544,N_17044,N_17668);
and U18545 (N_18545,N_17756,N_17700);
or U18546 (N_18546,N_17906,N_17391);
nand U18547 (N_18547,N_17021,N_17697);
nand U18548 (N_18548,N_17047,N_17085);
nor U18549 (N_18549,N_17888,N_17847);
or U18550 (N_18550,N_17759,N_17914);
or U18551 (N_18551,N_17217,N_17532);
or U18552 (N_18552,N_17804,N_17380);
nand U18553 (N_18553,N_17201,N_17156);
nand U18554 (N_18554,N_17537,N_17520);
nand U18555 (N_18555,N_17985,N_17193);
nand U18556 (N_18556,N_17358,N_17016);
nor U18557 (N_18557,N_17263,N_17723);
and U18558 (N_18558,N_17283,N_17076);
and U18559 (N_18559,N_17061,N_17308);
or U18560 (N_18560,N_17509,N_17513);
nand U18561 (N_18561,N_17486,N_17908);
and U18562 (N_18562,N_17671,N_17572);
xor U18563 (N_18563,N_17156,N_17210);
nor U18564 (N_18564,N_17329,N_17000);
or U18565 (N_18565,N_17986,N_17882);
or U18566 (N_18566,N_17658,N_17711);
nand U18567 (N_18567,N_17018,N_17889);
or U18568 (N_18568,N_17745,N_17971);
xor U18569 (N_18569,N_17575,N_17826);
xnor U18570 (N_18570,N_17942,N_17013);
and U18571 (N_18571,N_17260,N_17844);
or U18572 (N_18572,N_17810,N_17091);
nand U18573 (N_18573,N_17118,N_17856);
xor U18574 (N_18574,N_17232,N_17178);
xor U18575 (N_18575,N_17352,N_17463);
or U18576 (N_18576,N_17671,N_17747);
or U18577 (N_18577,N_17185,N_17990);
nand U18578 (N_18578,N_17690,N_17863);
xor U18579 (N_18579,N_17702,N_17695);
and U18580 (N_18580,N_17941,N_17001);
and U18581 (N_18581,N_17511,N_17927);
xnor U18582 (N_18582,N_17431,N_17840);
nor U18583 (N_18583,N_17953,N_17334);
nor U18584 (N_18584,N_17303,N_17858);
xor U18585 (N_18585,N_17614,N_17424);
nand U18586 (N_18586,N_17571,N_17871);
nand U18587 (N_18587,N_17367,N_17905);
nor U18588 (N_18588,N_17666,N_17356);
or U18589 (N_18589,N_17140,N_17695);
and U18590 (N_18590,N_17015,N_17820);
or U18591 (N_18591,N_17783,N_17915);
nand U18592 (N_18592,N_17900,N_17682);
nor U18593 (N_18593,N_17113,N_17731);
xnor U18594 (N_18594,N_17857,N_17248);
and U18595 (N_18595,N_17397,N_17957);
nand U18596 (N_18596,N_17259,N_17548);
and U18597 (N_18597,N_17042,N_17000);
and U18598 (N_18598,N_17409,N_17925);
nand U18599 (N_18599,N_17738,N_17662);
and U18600 (N_18600,N_17485,N_17002);
xor U18601 (N_18601,N_17331,N_17235);
or U18602 (N_18602,N_17741,N_17687);
and U18603 (N_18603,N_17363,N_17396);
nor U18604 (N_18604,N_17865,N_17278);
and U18605 (N_18605,N_17208,N_17389);
and U18606 (N_18606,N_17760,N_17160);
xor U18607 (N_18607,N_17241,N_17474);
nand U18608 (N_18608,N_17622,N_17794);
nor U18609 (N_18609,N_17148,N_17542);
nor U18610 (N_18610,N_17303,N_17194);
or U18611 (N_18611,N_17843,N_17197);
and U18612 (N_18612,N_17070,N_17450);
xnor U18613 (N_18613,N_17100,N_17274);
nand U18614 (N_18614,N_17785,N_17798);
nor U18615 (N_18615,N_17280,N_17465);
or U18616 (N_18616,N_17437,N_17941);
or U18617 (N_18617,N_17365,N_17521);
nand U18618 (N_18618,N_17874,N_17423);
nor U18619 (N_18619,N_17270,N_17189);
xor U18620 (N_18620,N_17283,N_17385);
nand U18621 (N_18621,N_17305,N_17074);
and U18622 (N_18622,N_17974,N_17442);
xnor U18623 (N_18623,N_17712,N_17199);
nor U18624 (N_18624,N_17386,N_17984);
or U18625 (N_18625,N_17113,N_17648);
nand U18626 (N_18626,N_17843,N_17203);
nand U18627 (N_18627,N_17903,N_17324);
or U18628 (N_18628,N_17537,N_17400);
xor U18629 (N_18629,N_17829,N_17680);
or U18630 (N_18630,N_17090,N_17439);
nor U18631 (N_18631,N_17248,N_17654);
nor U18632 (N_18632,N_17742,N_17995);
and U18633 (N_18633,N_17603,N_17909);
nor U18634 (N_18634,N_17853,N_17604);
or U18635 (N_18635,N_17097,N_17969);
and U18636 (N_18636,N_17266,N_17286);
or U18637 (N_18637,N_17610,N_17890);
nor U18638 (N_18638,N_17969,N_17362);
or U18639 (N_18639,N_17052,N_17119);
and U18640 (N_18640,N_17352,N_17610);
nor U18641 (N_18641,N_17212,N_17326);
xor U18642 (N_18642,N_17311,N_17231);
xnor U18643 (N_18643,N_17040,N_17849);
and U18644 (N_18644,N_17011,N_17335);
nand U18645 (N_18645,N_17979,N_17447);
xor U18646 (N_18646,N_17898,N_17512);
and U18647 (N_18647,N_17063,N_17922);
and U18648 (N_18648,N_17898,N_17055);
xor U18649 (N_18649,N_17614,N_17691);
or U18650 (N_18650,N_17591,N_17678);
nor U18651 (N_18651,N_17413,N_17998);
and U18652 (N_18652,N_17821,N_17501);
nor U18653 (N_18653,N_17832,N_17093);
or U18654 (N_18654,N_17015,N_17879);
or U18655 (N_18655,N_17969,N_17072);
xor U18656 (N_18656,N_17583,N_17297);
xor U18657 (N_18657,N_17144,N_17635);
and U18658 (N_18658,N_17425,N_17181);
nor U18659 (N_18659,N_17271,N_17437);
nor U18660 (N_18660,N_17644,N_17780);
and U18661 (N_18661,N_17291,N_17903);
nand U18662 (N_18662,N_17678,N_17714);
nand U18663 (N_18663,N_17004,N_17605);
nand U18664 (N_18664,N_17523,N_17786);
or U18665 (N_18665,N_17353,N_17507);
nand U18666 (N_18666,N_17593,N_17007);
or U18667 (N_18667,N_17981,N_17654);
and U18668 (N_18668,N_17268,N_17055);
or U18669 (N_18669,N_17691,N_17091);
nand U18670 (N_18670,N_17898,N_17156);
or U18671 (N_18671,N_17146,N_17639);
nor U18672 (N_18672,N_17010,N_17526);
nand U18673 (N_18673,N_17896,N_17982);
and U18674 (N_18674,N_17648,N_17092);
nor U18675 (N_18675,N_17478,N_17384);
and U18676 (N_18676,N_17702,N_17365);
xor U18677 (N_18677,N_17420,N_17245);
nand U18678 (N_18678,N_17621,N_17750);
nand U18679 (N_18679,N_17772,N_17529);
or U18680 (N_18680,N_17367,N_17179);
or U18681 (N_18681,N_17931,N_17298);
nand U18682 (N_18682,N_17069,N_17427);
or U18683 (N_18683,N_17787,N_17251);
nand U18684 (N_18684,N_17536,N_17674);
and U18685 (N_18685,N_17369,N_17517);
or U18686 (N_18686,N_17177,N_17352);
nor U18687 (N_18687,N_17908,N_17424);
nor U18688 (N_18688,N_17394,N_17648);
nor U18689 (N_18689,N_17902,N_17171);
xor U18690 (N_18690,N_17383,N_17871);
nor U18691 (N_18691,N_17574,N_17784);
nand U18692 (N_18692,N_17550,N_17455);
nand U18693 (N_18693,N_17030,N_17265);
or U18694 (N_18694,N_17334,N_17296);
and U18695 (N_18695,N_17816,N_17826);
or U18696 (N_18696,N_17813,N_17022);
nand U18697 (N_18697,N_17388,N_17669);
and U18698 (N_18698,N_17320,N_17569);
or U18699 (N_18699,N_17576,N_17750);
nor U18700 (N_18700,N_17302,N_17355);
nand U18701 (N_18701,N_17280,N_17438);
nand U18702 (N_18702,N_17805,N_17948);
or U18703 (N_18703,N_17942,N_17778);
nand U18704 (N_18704,N_17271,N_17808);
or U18705 (N_18705,N_17121,N_17317);
or U18706 (N_18706,N_17620,N_17915);
nand U18707 (N_18707,N_17468,N_17706);
nor U18708 (N_18708,N_17822,N_17232);
nand U18709 (N_18709,N_17614,N_17184);
nor U18710 (N_18710,N_17048,N_17338);
nand U18711 (N_18711,N_17291,N_17604);
nor U18712 (N_18712,N_17507,N_17567);
and U18713 (N_18713,N_17977,N_17848);
and U18714 (N_18714,N_17618,N_17677);
xnor U18715 (N_18715,N_17308,N_17515);
xor U18716 (N_18716,N_17171,N_17478);
or U18717 (N_18717,N_17638,N_17983);
nand U18718 (N_18718,N_17225,N_17977);
nand U18719 (N_18719,N_17303,N_17951);
and U18720 (N_18720,N_17742,N_17625);
or U18721 (N_18721,N_17708,N_17438);
and U18722 (N_18722,N_17048,N_17283);
and U18723 (N_18723,N_17100,N_17441);
and U18724 (N_18724,N_17294,N_17858);
xor U18725 (N_18725,N_17117,N_17962);
nand U18726 (N_18726,N_17191,N_17406);
nand U18727 (N_18727,N_17341,N_17676);
or U18728 (N_18728,N_17970,N_17424);
and U18729 (N_18729,N_17570,N_17637);
nor U18730 (N_18730,N_17834,N_17341);
nor U18731 (N_18731,N_17875,N_17640);
nand U18732 (N_18732,N_17087,N_17883);
xor U18733 (N_18733,N_17688,N_17128);
nand U18734 (N_18734,N_17570,N_17474);
or U18735 (N_18735,N_17208,N_17617);
nand U18736 (N_18736,N_17065,N_17524);
nand U18737 (N_18737,N_17857,N_17587);
and U18738 (N_18738,N_17628,N_17534);
and U18739 (N_18739,N_17897,N_17814);
xnor U18740 (N_18740,N_17412,N_17335);
nand U18741 (N_18741,N_17368,N_17635);
nand U18742 (N_18742,N_17180,N_17027);
xnor U18743 (N_18743,N_17585,N_17962);
and U18744 (N_18744,N_17862,N_17474);
nand U18745 (N_18745,N_17039,N_17910);
xor U18746 (N_18746,N_17580,N_17193);
nand U18747 (N_18747,N_17039,N_17978);
xor U18748 (N_18748,N_17846,N_17660);
xor U18749 (N_18749,N_17011,N_17241);
xor U18750 (N_18750,N_17304,N_17199);
nand U18751 (N_18751,N_17185,N_17776);
or U18752 (N_18752,N_17281,N_17659);
nand U18753 (N_18753,N_17422,N_17777);
nor U18754 (N_18754,N_17857,N_17806);
nand U18755 (N_18755,N_17199,N_17184);
nor U18756 (N_18756,N_17951,N_17313);
and U18757 (N_18757,N_17977,N_17327);
nand U18758 (N_18758,N_17579,N_17229);
and U18759 (N_18759,N_17313,N_17014);
nor U18760 (N_18760,N_17857,N_17279);
or U18761 (N_18761,N_17321,N_17257);
xnor U18762 (N_18762,N_17160,N_17429);
xor U18763 (N_18763,N_17242,N_17521);
and U18764 (N_18764,N_17786,N_17363);
nor U18765 (N_18765,N_17731,N_17956);
nand U18766 (N_18766,N_17498,N_17942);
nand U18767 (N_18767,N_17874,N_17064);
or U18768 (N_18768,N_17233,N_17810);
nor U18769 (N_18769,N_17055,N_17246);
and U18770 (N_18770,N_17812,N_17325);
nand U18771 (N_18771,N_17475,N_17825);
nand U18772 (N_18772,N_17028,N_17950);
and U18773 (N_18773,N_17931,N_17490);
or U18774 (N_18774,N_17130,N_17906);
or U18775 (N_18775,N_17663,N_17306);
or U18776 (N_18776,N_17037,N_17726);
nand U18777 (N_18777,N_17289,N_17276);
and U18778 (N_18778,N_17153,N_17850);
or U18779 (N_18779,N_17012,N_17661);
and U18780 (N_18780,N_17983,N_17639);
nand U18781 (N_18781,N_17040,N_17128);
or U18782 (N_18782,N_17468,N_17002);
and U18783 (N_18783,N_17928,N_17358);
nor U18784 (N_18784,N_17941,N_17216);
or U18785 (N_18785,N_17527,N_17721);
nand U18786 (N_18786,N_17736,N_17385);
nor U18787 (N_18787,N_17435,N_17079);
nand U18788 (N_18788,N_17859,N_17932);
xnor U18789 (N_18789,N_17597,N_17800);
nand U18790 (N_18790,N_17908,N_17351);
and U18791 (N_18791,N_17495,N_17720);
xor U18792 (N_18792,N_17609,N_17544);
and U18793 (N_18793,N_17800,N_17179);
nand U18794 (N_18794,N_17529,N_17051);
xnor U18795 (N_18795,N_17253,N_17448);
nand U18796 (N_18796,N_17359,N_17057);
nor U18797 (N_18797,N_17190,N_17389);
or U18798 (N_18798,N_17397,N_17953);
nand U18799 (N_18799,N_17359,N_17662);
nor U18800 (N_18800,N_17870,N_17518);
nand U18801 (N_18801,N_17223,N_17453);
xnor U18802 (N_18802,N_17198,N_17657);
nor U18803 (N_18803,N_17644,N_17291);
and U18804 (N_18804,N_17749,N_17649);
nand U18805 (N_18805,N_17395,N_17296);
xor U18806 (N_18806,N_17429,N_17118);
xor U18807 (N_18807,N_17556,N_17331);
nor U18808 (N_18808,N_17178,N_17448);
xor U18809 (N_18809,N_17065,N_17672);
xnor U18810 (N_18810,N_17362,N_17412);
nand U18811 (N_18811,N_17585,N_17666);
nor U18812 (N_18812,N_17263,N_17275);
and U18813 (N_18813,N_17491,N_17018);
xnor U18814 (N_18814,N_17531,N_17933);
nor U18815 (N_18815,N_17888,N_17157);
nor U18816 (N_18816,N_17087,N_17945);
and U18817 (N_18817,N_17061,N_17564);
nor U18818 (N_18818,N_17393,N_17688);
and U18819 (N_18819,N_17951,N_17612);
nand U18820 (N_18820,N_17409,N_17061);
xnor U18821 (N_18821,N_17962,N_17071);
xnor U18822 (N_18822,N_17049,N_17228);
nor U18823 (N_18823,N_17058,N_17138);
nor U18824 (N_18824,N_17537,N_17999);
or U18825 (N_18825,N_17870,N_17195);
and U18826 (N_18826,N_17244,N_17066);
nor U18827 (N_18827,N_17987,N_17232);
xnor U18828 (N_18828,N_17622,N_17925);
nor U18829 (N_18829,N_17964,N_17358);
or U18830 (N_18830,N_17977,N_17516);
nor U18831 (N_18831,N_17911,N_17147);
xor U18832 (N_18832,N_17374,N_17478);
and U18833 (N_18833,N_17703,N_17540);
or U18834 (N_18834,N_17409,N_17974);
and U18835 (N_18835,N_17601,N_17195);
nand U18836 (N_18836,N_17857,N_17534);
nand U18837 (N_18837,N_17568,N_17379);
and U18838 (N_18838,N_17923,N_17380);
nand U18839 (N_18839,N_17118,N_17112);
nor U18840 (N_18840,N_17648,N_17632);
nand U18841 (N_18841,N_17911,N_17021);
and U18842 (N_18842,N_17533,N_17657);
or U18843 (N_18843,N_17454,N_17881);
or U18844 (N_18844,N_17986,N_17968);
nand U18845 (N_18845,N_17097,N_17258);
nand U18846 (N_18846,N_17357,N_17306);
nand U18847 (N_18847,N_17893,N_17231);
nor U18848 (N_18848,N_17100,N_17807);
or U18849 (N_18849,N_17877,N_17577);
and U18850 (N_18850,N_17737,N_17517);
and U18851 (N_18851,N_17208,N_17214);
or U18852 (N_18852,N_17985,N_17843);
or U18853 (N_18853,N_17589,N_17850);
or U18854 (N_18854,N_17314,N_17681);
and U18855 (N_18855,N_17980,N_17048);
and U18856 (N_18856,N_17541,N_17608);
nor U18857 (N_18857,N_17445,N_17018);
or U18858 (N_18858,N_17455,N_17025);
xnor U18859 (N_18859,N_17665,N_17756);
nor U18860 (N_18860,N_17855,N_17995);
or U18861 (N_18861,N_17807,N_17564);
nand U18862 (N_18862,N_17593,N_17306);
nor U18863 (N_18863,N_17483,N_17206);
nand U18864 (N_18864,N_17415,N_17735);
nand U18865 (N_18865,N_17057,N_17697);
nor U18866 (N_18866,N_17923,N_17477);
nand U18867 (N_18867,N_17202,N_17602);
nand U18868 (N_18868,N_17209,N_17785);
nand U18869 (N_18869,N_17703,N_17216);
xor U18870 (N_18870,N_17162,N_17878);
nand U18871 (N_18871,N_17275,N_17929);
xor U18872 (N_18872,N_17302,N_17487);
and U18873 (N_18873,N_17095,N_17603);
xor U18874 (N_18874,N_17163,N_17195);
and U18875 (N_18875,N_17218,N_17060);
nor U18876 (N_18876,N_17091,N_17320);
xnor U18877 (N_18877,N_17939,N_17064);
or U18878 (N_18878,N_17827,N_17184);
or U18879 (N_18879,N_17594,N_17790);
xnor U18880 (N_18880,N_17223,N_17073);
nand U18881 (N_18881,N_17170,N_17134);
and U18882 (N_18882,N_17575,N_17076);
and U18883 (N_18883,N_17224,N_17969);
nand U18884 (N_18884,N_17065,N_17183);
or U18885 (N_18885,N_17658,N_17273);
nand U18886 (N_18886,N_17229,N_17319);
nor U18887 (N_18887,N_17440,N_17271);
nand U18888 (N_18888,N_17293,N_17846);
and U18889 (N_18889,N_17563,N_17070);
and U18890 (N_18890,N_17983,N_17453);
or U18891 (N_18891,N_17377,N_17786);
nor U18892 (N_18892,N_17041,N_17725);
and U18893 (N_18893,N_17799,N_17954);
nor U18894 (N_18894,N_17636,N_17769);
xor U18895 (N_18895,N_17193,N_17031);
nor U18896 (N_18896,N_17369,N_17944);
xor U18897 (N_18897,N_17746,N_17419);
xor U18898 (N_18898,N_17202,N_17581);
xnor U18899 (N_18899,N_17395,N_17377);
xor U18900 (N_18900,N_17859,N_17776);
or U18901 (N_18901,N_17596,N_17160);
xor U18902 (N_18902,N_17017,N_17020);
xnor U18903 (N_18903,N_17984,N_17442);
and U18904 (N_18904,N_17770,N_17197);
and U18905 (N_18905,N_17886,N_17426);
nand U18906 (N_18906,N_17546,N_17553);
and U18907 (N_18907,N_17072,N_17346);
and U18908 (N_18908,N_17512,N_17959);
nand U18909 (N_18909,N_17224,N_17648);
xor U18910 (N_18910,N_17038,N_17123);
nand U18911 (N_18911,N_17307,N_17531);
nor U18912 (N_18912,N_17388,N_17130);
xor U18913 (N_18913,N_17299,N_17524);
xor U18914 (N_18914,N_17454,N_17337);
or U18915 (N_18915,N_17221,N_17736);
and U18916 (N_18916,N_17042,N_17685);
and U18917 (N_18917,N_17581,N_17113);
xor U18918 (N_18918,N_17730,N_17570);
xor U18919 (N_18919,N_17601,N_17737);
nand U18920 (N_18920,N_17104,N_17255);
and U18921 (N_18921,N_17067,N_17764);
or U18922 (N_18922,N_17547,N_17310);
or U18923 (N_18923,N_17060,N_17298);
nor U18924 (N_18924,N_17076,N_17052);
xor U18925 (N_18925,N_17103,N_17848);
xor U18926 (N_18926,N_17502,N_17512);
and U18927 (N_18927,N_17006,N_17047);
or U18928 (N_18928,N_17174,N_17177);
and U18929 (N_18929,N_17753,N_17287);
nand U18930 (N_18930,N_17252,N_17601);
or U18931 (N_18931,N_17617,N_17723);
and U18932 (N_18932,N_17235,N_17224);
nor U18933 (N_18933,N_17791,N_17772);
xnor U18934 (N_18934,N_17227,N_17156);
xor U18935 (N_18935,N_17718,N_17773);
or U18936 (N_18936,N_17187,N_17907);
nor U18937 (N_18937,N_17764,N_17041);
or U18938 (N_18938,N_17481,N_17561);
nor U18939 (N_18939,N_17874,N_17176);
and U18940 (N_18940,N_17097,N_17475);
nand U18941 (N_18941,N_17612,N_17945);
nand U18942 (N_18942,N_17005,N_17933);
xnor U18943 (N_18943,N_17516,N_17966);
nand U18944 (N_18944,N_17050,N_17446);
nand U18945 (N_18945,N_17335,N_17569);
and U18946 (N_18946,N_17831,N_17099);
nor U18947 (N_18947,N_17410,N_17375);
nand U18948 (N_18948,N_17755,N_17616);
nor U18949 (N_18949,N_17235,N_17807);
nand U18950 (N_18950,N_17688,N_17434);
nor U18951 (N_18951,N_17503,N_17080);
xnor U18952 (N_18952,N_17690,N_17882);
xnor U18953 (N_18953,N_17376,N_17189);
xnor U18954 (N_18954,N_17241,N_17918);
or U18955 (N_18955,N_17963,N_17066);
nor U18956 (N_18956,N_17639,N_17446);
and U18957 (N_18957,N_17396,N_17469);
xnor U18958 (N_18958,N_17758,N_17163);
and U18959 (N_18959,N_17303,N_17943);
nand U18960 (N_18960,N_17268,N_17426);
nor U18961 (N_18961,N_17334,N_17292);
and U18962 (N_18962,N_17247,N_17727);
xnor U18963 (N_18963,N_17152,N_17937);
nor U18964 (N_18964,N_17887,N_17778);
or U18965 (N_18965,N_17087,N_17824);
xnor U18966 (N_18966,N_17944,N_17655);
or U18967 (N_18967,N_17131,N_17218);
nand U18968 (N_18968,N_17749,N_17905);
or U18969 (N_18969,N_17090,N_17847);
nand U18970 (N_18970,N_17725,N_17274);
or U18971 (N_18971,N_17578,N_17536);
and U18972 (N_18972,N_17108,N_17979);
nor U18973 (N_18973,N_17092,N_17150);
xnor U18974 (N_18974,N_17642,N_17239);
nand U18975 (N_18975,N_17709,N_17505);
nor U18976 (N_18976,N_17543,N_17477);
and U18977 (N_18977,N_17493,N_17127);
nand U18978 (N_18978,N_17376,N_17020);
or U18979 (N_18979,N_17119,N_17634);
and U18980 (N_18980,N_17618,N_17847);
or U18981 (N_18981,N_17493,N_17803);
nand U18982 (N_18982,N_17348,N_17463);
nand U18983 (N_18983,N_17429,N_17488);
nand U18984 (N_18984,N_17972,N_17892);
or U18985 (N_18985,N_17642,N_17551);
and U18986 (N_18986,N_17843,N_17909);
nor U18987 (N_18987,N_17677,N_17829);
or U18988 (N_18988,N_17656,N_17243);
or U18989 (N_18989,N_17639,N_17603);
or U18990 (N_18990,N_17262,N_17882);
nor U18991 (N_18991,N_17896,N_17108);
and U18992 (N_18992,N_17427,N_17219);
xnor U18993 (N_18993,N_17586,N_17256);
and U18994 (N_18994,N_17692,N_17039);
or U18995 (N_18995,N_17695,N_17254);
xnor U18996 (N_18996,N_17551,N_17970);
or U18997 (N_18997,N_17626,N_17161);
and U18998 (N_18998,N_17796,N_17482);
or U18999 (N_18999,N_17747,N_17616);
nor U19000 (N_19000,N_18085,N_18434);
nand U19001 (N_19001,N_18951,N_18754);
and U19002 (N_19002,N_18809,N_18119);
nor U19003 (N_19003,N_18051,N_18839);
nand U19004 (N_19004,N_18682,N_18654);
nor U19005 (N_19005,N_18784,N_18231);
nor U19006 (N_19006,N_18385,N_18848);
and U19007 (N_19007,N_18121,N_18732);
nand U19008 (N_19008,N_18803,N_18959);
and U19009 (N_19009,N_18221,N_18915);
xor U19010 (N_19010,N_18762,N_18199);
or U19011 (N_19011,N_18403,N_18257);
nor U19012 (N_19012,N_18646,N_18826);
xnor U19013 (N_19013,N_18426,N_18308);
and U19014 (N_19014,N_18091,N_18154);
xor U19015 (N_19015,N_18755,N_18453);
and U19016 (N_19016,N_18787,N_18550);
nand U19017 (N_19017,N_18963,N_18381);
nand U19018 (N_19018,N_18602,N_18499);
nor U19019 (N_19019,N_18105,N_18948);
or U19020 (N_19020,N_18374,N_18026);
nor U19021 (N_19021,N_18817,N_18876);
or U19022 (N_19022,N_18413,N_18759);
and U19023 (N_19023,N_18421,N_18081);
and U19024 (N_19024,N_18920,N_18225);
or U19025 (N_19025,N_18684,N_18238);
or U19026 (N_19026,N_18962,N_18856);
and U19027 (N_19027,N_18693,N_18987);
or U19028 (N_19028,N_18635,N_18446);
nand U19029 (N_19029,N_18389,N_18651);
xnor U19030 (N_19030,N_18407,N_18571);
xor U19031 (N_19031,N_18997,N_18983);
nor U19032 (N_19032,N_18266,N_18899);
nor U19033 (N_19033,N_18758,N_18484);
nand U19034 (N_19034,N_18598,N_18780);
nand U19035 (N_19035,N_18515,N_18017);
xor U19036 (N_19036,N_18361,N_18069);
nand U19037 (N_19037,N_18551,N_18717);
xnor U19038 (N_19038,N_18622,N_18675);
nand U19039 (N_19039,N_18212,N_18104);
nand U19040 (N_19040,N_18898,N_18103);
and U19041 (N_19041,N_18127,N_18993);
nand U19042 (N_19042,N_18362,N_18269);
xor U19043 (N_19043,N_18541,N_18241);
nand U19044 (N_19044,N_18366,N_18882);
and U19045 (N_19045,N_18331,N_18152);
xnor U19046 (N_19046,N_18353,N_18042);
nand U19047 (N_19047,N_18073,N_18520);
or U19048 (N_19048,N_18650,N_18735);
nor U19049 (N_19049,N_18981,N_18877);
xor U19050 (N_19050,N_18427,N_18686);
and U19051 (N_19051,N_18075,N_18343);
or U19052 (N_19052,N_18246,N_18796);
and U19053 (N_19053,N_18628,N_18388);
xnor U19054 (N_19054,N_18102,N_18275);
nand U19055 (N_19055,N_18857,N_18038);
xnor U19056 (N_19056,N_18814,N_18953);
or U19057 (N_19057,N_18866,N_18138);
xnor U19058 (N_19058,N_18536,N_18701);
nor U19059 (N_19059,N_18947,N_18451);
or U19060 (N_19060,N_18317,N_18841);
nand U19061 (N_19061,N_18371,N_18255);
xnor U19062 (N_19062,N_18170,N_18032);
xor U19063 (N_19063,N_18113,N_18924);
and U19064 (N_19064,N_18641,N_18433);
xnor U19065 (N_19065,N_18593,N_18891);
xor U19066 (N_19066,N_18428,N_18088);
nor U19067 (N_19067,N_18647,N_18505);
nand U19068 (N_19068,N_18829,N_18538);
nor U19069 (N_19069,N_18100,N_18155);
or U19070 (N_19070,N_18128,N_18132);
nor U19071 (N_19071,N_18709,N_18853);
and U19072 (N_19072,N_18554,N_18063);
xor U19073 (N_19073,N_18933,N_18697);
nand U19074 (N_19074,N_18098,N_18872);
nor U19075 (N_19075,N_18849,N_18776);
or U19076 (N_19076,N_18844,N_18518);
nor U19077 (N_19077,N_18498,N_18464);
nand U19078 (N_19078,N_18478,N_18035);
xor U19079 (N_19079,N_18577,N_18001);
nor U19080 (N_19080,N_18354,N_18120);
xor U19081 (N_19081,N_18587,N_18367);
nor U19082 (N_19082,N_18846,N_18752);
nor U19083 (N_19083,N_18307,N_18114);
and U19084 (N_19084,N_18357,N_18086);
xnor U19085 (N_19085,N_18481,N_18182);
or U19086 (N_19086,N_18047,N_18563);
or U19087 (N_19087,N_18410,N_18880);
nor U19088 (N_19088,N_18019,N_18881);
and U19089 (N_19089,N_18268,N_18486);
nand U19090 (N_19090,N_18277,N_18319);
xnor U19091 (N_19091,N_18286,N_18117);
nand U19092 (N_19092,N_18629,N_18724);
and U19093 (N_19093,N_18733,N_18420);
or U19094 (N_19094,N_18688,N_18992);
nand U19095 (N_19095,N_18958,N_18581);
nor U19096 (N_19096,N_18150,N_18730);
xnor U19097 (N_19097,N_18249,N_18557);
xnor U19098 (N_19098,N_18873,N_18202);
or U19099 (N_19099,N_18626,N_18471);
or U19100 (N_19100,N_18183,N_18502);
or U19101 (N_19101,N_18350,N_18850);
and U19102 (N_19102,N_18671,N_18594);
and U19103 (N_19103,N_18312,N_18140);
nor U19104 (N_19104,N_18384,N_18111);
nand U19105 (N_19105,N_18614,N_18309);
or U19106 (N_19106,N_18175,N_18519);
and U19107 (N_19107,N_18835,N_18833);
and U19108 (N_19108,N_18544,N_18721);
or U19109 (N_19109,N_18610,N_18136);
and U19110 (N_19110,N_18698,N_18004);
and U19111 (N_19111,N_18251,N_18665);
nand U19112 (N_19112,N_18674,N_18692);
xor U19113 (N_19113,N_18763,N_18879);
and U19114 (N_19114,N_18886,N_18009);
nor U19115 (N_19115,N_18049,N_18176);
and U19116 (N_19116,N_18524,N_18852);
xnor U19117 (N_19117,N_18445,N_18438);
nor U19118 (N_19118,N_18909,N_18971);
xnor U19119 (N_19119,N_18097,N_18562);
nor U19120 (N_19120,N_18482,N_18028);
nor U19121 (N_19121,N_18585,N_18930);
xnor U19122 (N_19122,N_18437,N_18363);
or U19123 (N_19123,N_18168,N_18156);
and U19124 (N_19124,N_18235,N_18072);
nor U19125 (N_19125,N_18099,N_18859);
nand U19126 (N_19126,N_18704,N_18939);
and U19127 (N_19127,N_18213,N_18193);
xor U19128 (N_19128,N_18510,N_18552);
xor U19129 (N_19129,N_18321,N_18443);
or U19130 (N_19130,N_18813,N_18060);
or U19131 (N_19131,N_18087,N_18601);
or U19132 (N_19132,N_18964,N_18984);
xor U19133 (N_19133,N_18294,N_18261);
or U19134 (N_19134,N_18200,N_18477);
nand U19135 (N_19135,N_18301,N_18095);
nand U19136 (N_19136,N_18638,N_18122);
nor U19137 (N_19137,N_18253,N_18021);
nor U19138 (N_19138,N_18897,N_18995);
nor U19139 (N_19139,N_18494,N_18956);
nand U19140 (N_19140,N_18018,N_18262);
nor U19141 (N_19141,N_18123,N_18861);
nand U19142 (N_19142,N_18435,N_18912);
xor U19143 (N_19143,N_18497,N_18398);
nor U19144 (N_19144,N_18133,N_18436);
and U19145 (N_19145,N_18927,N_18643);
xnor U19146 (N_19146,N_18712,N_18273);
xor U19147 (N_19147,N_18240,N_18228);
xor U19148 (N_19148,N_18224,N_18474);
or U19149 (N_19149,N_18694,N_18961);
nor U19150 (N_19150,N_18400,N_18816);
or U19151 (N_19151,N_18592,N_18089);
or U19152 (N_19152,N_18279,N_18823);
xor U19153 (N_19153,N_18973,N_18239);
nand U19154 (N_19154,N_18488,N_18655);
xnor U19155 (N_19155,N_18146,N_18864);
nor U19156 (N_19156,N_18621,N_18575);
or U19157 (N_19157,N_18292,N_18349);
nand U19158 (N_19158,N_18931,N_18719);
or U19159 (N_19159,N_18925,N_18226);
nor U19160 (N_19160,N_18907,N_18387);
and U19161 (N_19161,N_18600,N_18703);
or U19162 (N_19162,N_18046,N_18157);
xnor U19163 (N_19163,N_18667,N_18523);
nor U19164 (N_19164,N_18738,N_18782);
nand U19165 (N_19165,N_18599,N_18247);
or U19166 (N_19166,N_18854,N_18574);
xnor U19167 (N_19167,N_18534,N_18302);
and U19168 (N_19168,N_18408,N_18805);
nand U19169 (N_19169,N_18663,N_18528);
nand U19170 (N_19170,N_18611,N_18492);
and U19171 (N_19171,N_18910,N_18586);
nor U19172 (N_19172,N_18061,N_18661);
or U19173 (N_19173,N_18386,N_18397);
and U19174 (N_19174,N_18040,N_18680);
nor U19175 (N_19175,N_18632,N_18209);
and U19176 (N_19176,N_18589,N_18695);
nand U19177 (N_19177,N_18820,N_18162);
nor U19178 (N_19178,N_18053,N_18000);
nor U19179 (N_19179,N_18144,N_18802);
nand U19180 (N_19180,N_18940,N_18934);
nor U19181 (N_19181,N_18896,N_18358);
nand U19182 (N_19182,N_18489,N_18690);
and U19183 (N_19183,N_18423,N_18818);
nand U19184 (N_19184,N_18596,N_18198);
xnor U19185 (N_19185,N_18618,N_18360);
nand U19186 (N_19186,N_18744,N_18804);
and U19187 (N_19187,N_18998,N_18245);
nand U19188 (N_19188,N_18994,N_18475);
and U19189 (N_19189,N_18346,N_18705);
or U19190 (N_19190,N_18625,N_18783);
or U19191 (N_19191,N_18707,N_18822);
or U19192 (N_19192,N_18210,N_18798);
nor U19193 (N_19193,N_18570,N_18828);
xor U19194 (N_19194,N_18941,N_18553);
and U19195 (N_19195,N_18027,N_18821);
or U19196 (N_19196,N_18236,N_18379);
and U19197 (N_19197,N_18616,N_18189);
nand U19198 (N_19198,N_18406,N_18677);
and U19199 (N_19199,N_18967,N_18149);
or U19200 (N_19200,N_18003,N_18756);
nor U19201 (N_19201,N_18270,N_18214);
or U19202 (N_19202,N_18480,N_18883);
nand U19203 (N_19203,N_18578,N_18008);
xnor U19204 (N_19204,N_18186,N_18159);
nor U19205 (N_19205,N_18380,N_18250);
nand U19206 (N_19206,N_18867,N_18615);
or U19207 (N_19207,N_18169,N_18532);
nor U19208 (N_19208,N_18917,N_18448);
and U19209 (N_19209,N_18888,N_18281);
or U19210 (N_19210,N_18761,N_18539);
nand U19211 (N_19211,N_18276,N_18630);
or U19212 (N_19212,N_18944,N_18267);
or U19213 (N_19213,N_18161,N_18955);
xor U19214 (N_19214,N_18352,N_18711);
or U19215 (N_19215,N_18383,N_18968);
xor U19216 (N_19216,N_18504,N_18710);
and U19217 (N_19217,N_18942,N_18952);
nor U19218 (N_19218,N_18364,N_18836);
and U19219 (N_19219,N_18860,N_18056);
or U19220 (N_19220,N_18179,N_18633);
xnor U19221 (N_19221,N_18229,N_18837);
xor U19222 (N_19222,N_18370,N_18439);
or U19223 (N_19223,N_18414,N_18048);
xnor U19224 (N_19224,N_18237,N_18310);
xor U19225 (N_19225,N_18351,N_18065);
or U19226 (N_19226,N_18449,N_18691);
nand U19227 (N_19227,N_18298,N_18219);
nor U19228 (N_19228,N_18007,N_18749);
nor U19229 (N_19229,N_18634,N_18772);
xnor U19230 (N_19230,N_18868,N_18143);
nand U19231 (N_19231,N_18954,N_18679);
xor U19232 (N_19232,N_18535,N_18166);
and U19233 (N_19233,N_18324,N_18187);
and U19234 (N_19234,N_18583,N_18005);
xor U19235 (N_19235,N_18607,N_18045);
or U19236 (N_19236,N_18232,N_18068);
xor U19237 (N_19237,N_18450,N_18767);
nor U19238 (N_19238,N_18845,N_18503);
xnor U19239 (N_19239,N_18858,N_18681);
nand U19240 (N_19240,N_18177,N_18293);
or U19241 (N_19241,N_18530,N_18750);
nand U19242 (N_19242,N_18299,N_18115);
xnor U19243 (N_19243,N_18922,N_18558);
xnor U19244 (N_19244,N_18597,N_18440);
or U19245 (N_19245,N_18878,N_18141);
or U19246 (N_19246,N_18982,N_18466);
xor U19247 (N_19247,N_18274,N_18781);
nor U19248 (N_19248,N_18769,N_18648);
xnor U19249 (N_19249,N_18030,N_18071);
and U19250 (N_19250,N_18545,N_18430);
and U19251 (N_19251,N_18945,N_18057);
nand U19252 (N_19252,N_18425,N_18230);
or U19253 (N_19253,N_18173,N_18472);
xnor U19254 (N_19254,N_18569,N_18637);
xnor U19255 (N_19255,N_18672,N_18893);
and U19256 (N_19256,N_18206,N_18770);
xnor U19257 (N_19257,N_18799,N_18044);
nand U19258 (N_19258,N_18424,N_18334);
xor U19259 (N_19259,N_18623,N_18470);
nor U19260 (N_19260,N_18264,N_18295);
nand U19261 (N_19261,N_18333,N_18404);
xor U19262 (N_19262,N_18673,N_18521);
xnor U19263 (N_19263,N_18741,N_18130);
xor U19264 (N_19264,N_18743,N_18092);
or U19265 (N_19265,N_18313,N_18792);
or U19266 (N_19266,N_18957,N_18617);
or U19267 (N_19267,N_18344,N_18107);
and U19268 (N_19268,N_18723,N_18024);
nor U19269 (N_19269,N_18476,N_18365);
xnor U19270 (N_19270,N_18727,N_18506);
or U19271 (N_19271,N_18700,N_18522);
and U19272 (N_19272,N_18547,N_18254);
nand U19273 (N_19273,N_18659,N_18300);
nand U19274 (N_19274,N_18559,N_18288);
and U19275 (N_19275,N_18025,N_18341);
or U19276 (N_19276,N_18928,N_18272);
nor U19277 (N_19277,N_18533,N_18218);
or U19278 (N_19278,N_18077,N_18969);
and U19279 (N_19279,N_18980,N_18336);
nand U19280 (N_19280,N_18487,N_18171);
and U19281 (N_19281,N_18417,N_18718);
xor U19282 (N_19282,N_18495,N_18582);
nand U19283 (N_19283,N_18014,N_18282);
nor U19284 (N_19284,N_18566,N_18908);
nor U19285 (N_19285,N_18819,N_18320);
or U19286 (N_19286,N_18283,N_18285);
and U19287 (N_19287,N_18702,N_18514);
nand U19288 (N_19288,N_18913,N_18936);
nor U19289 (N_19289,N_18062,N_18517);
and U19290 (N_19290,N_18863,N_18181);
nor U19291 (N_19291,N_18560,N_18184);
nor U19292 (N_19292,N_18568,N_18670);
nand U19293 (N_19293,N_18946,N_18023);
or U19294 (N_19294,N_18619,N_18603);
xnor U19295 (N_19295,N_18479,N_18919);
or U19296 (N_19296,N_18656,N_18167);
nand U19297 (N_19297,N_18851,N_18865);
xor U19298 (N_19298,N_18824,N_18271);
xor U19299 (N_19299,N_18855,N_18706);
xnor U19300 (N_19300,N_18631,N_18079);
or U19301 (N_19301,N_18485,N_18010);
xor U19302 (N_19302,N_18305,N_18794);
and U19303 (N_19303,N_18605,N_18084);
nor U19304 (N_19304,N_18842,N_18016);
nor U19305 (N_19305,N_18037,N_18429);
nand U19306 (N_19306,N_18106,N_18033);
nor U19307 (N_19307,N_18444,N_18699);
nor U19308 (N_19308,N_18064,N_18252);
nor U19309 (N_19309,N_18258,N_18290);
nor U19310 (N_19310,N_18059,N_18676);
nor U19311 (N_19311,N_18359,N_18223);
nand U19312 (N_19312,N_18895,N_18929);
or U19313 (N_19313,N_18134,N_18368);
nand U19314 (N_19314,N_18843,N_18938);
nor U19315 (N_19315,N_18043,N_18467);
nand U19316 (N_19316,N_18500,N_18034);
nor U19317 (N_19317,N_18652,N_18297);
xor U19318 (N_19318,N_18180,N_18260);
nor U19319 (N_19319,N_18287,N_18462);
nor U19320 (N_19320,N_18543,N_18172);
or U19321 (N_19321,N_18685,N_18527);
xnor U19322 (N_19322,N_18259,N_18979);
xor U19323 (N_19323,N_18020,N_18052);
or U19324 (N_19324,N_18431,N_18999);
and U19325 (N_19325,N_18160,N_18960);
xor U19326 (N_19326,N_18204,N_18070);
and U19327 (N_19327,N_18325,N_18966);
or U19328 (N_19328,N_18894,N_18190);
or U19329 (N_19329,N_18788,N_18725);
or U19330 (N_19330,N_18461,N_18082);
nand U19331 (N_19331,N_18728,N_18716);
and U19332 (N_19332,N_18165,N_18509);
xnor U19333 (N_19333,N_18567,N_18548);
or U19334 (N_19334,N_18139,N_18454);
or U19335 (N_19335,N_18764,N_18375);
or U19336 (N_19336,N_18011,N_18986);
nor U19337 (N_19337,N_18904,N_18330);
nand U19338 (N_19338,N_18965,N_18263);
xor U19339 (N_19339,N_18163,N_18457);
nor U19340 (N_19340,N_18194,N_18396);
xnor U19341 (N_19341,N_18278,N_18142);
nand U19342 (N_19342,N_18327,N_18174);
nand U19343 (N_19343,N_18771,N_18790);
nand U19344 (N_19344,N_18572,N_18496);
nor U19345 (N_19345,N_18542,N_18409);
and U19346 (N_19346,N_18284,N_18831);
and U19347 (N_19347,N_18664,N_18036);
nand U19348 (N_19348,N_18076,N_18722);
and U19349 (N_19349,N_18595,N_18129);
nand U19350 (N_19350,N_18977,N_18126);
xor U19351 (N_19351,N_18714,N_18192);
or U19352 (N_19352,N_18653,N_18215);
or U19353 (N_19353,N_18540,N_18148);
nand U19354 (N_19354,N_18789,N_18207);
nor U19355 (N_19355,N_18892,N_18768);
and U19356 (N_19356,N_18797,N_18561);
nand U19357 (N_19357,N_18576,N_18393);
or U19358 (N_19358,N_18609,N_18525);
and U19359 (N_19359,N_18074,N_18734);
or U19360 (N_19360,N_18657,N_18584);
nor U19361 (N_19361,N_18645,N_18490);
xor U19362 (N_19362,N_18890,N_18348);
or U19363 (N_19363,N_18329,N_18369);
nand U19364 (N_19364,N_18248,N_18748);
nor U19365 (N_19365,N_18322,N_18713);
xnor U19366 (N_19366,N_18415,N_18620);
xnor U19367 (N_19367,N_18151,N_18736);
or U19368 (N_19368,N_18950,N_18949);
nor U19369 (N_19369,N_18658,N_18546);
and U19370 (N_19370,N_18473,N_18501);
nand U19371 (N_19371,N_18978,N_18678);
and U19372 (N_19372,N_18468,N_18564);
and U19373 (N_19373,N_18145,N_18990);
and U19374 (N_19374,N_18887,N_18164);
xor U19375 (N_19375,N_18339,N_18234);
xor U19376 (N_19376,N_18627,N_18916);
or U19377 (N_19377,N_18318,N_18080);
nand U19378 (N_19378,N_18178,N_18906);
or U19379 (N_19379,N_18459,N_18591);
and U19380 (N_19380,N_18465,N_18903);
xor U19381 (N_19381,N_18800,N_18382);
nor U19382 (N_19382,N_18217,N_18777);
nor U19383 (N_19383,N_18233,N_18394);
xnor U19384 (N_19384,N_18315,N_18041);
xor U19385 (N_19385,N_18751,N_18093);
nor U19386 (N_19386,N_18469,N_18642);
and U19387 (N_19387,N_18411,N_18884);
nor U19388 (N_19388,N_18911,N_18205);
nand U19389 (N_19389,N_18289,N_18323);
xnor U19390 (N_19390,N_18304,N_18280);
xnor U19391 (N_19391,N_18116,N_18242);
nor U19392 (N_19392,N_18644,N_18937);
or U19393 (N_19393,N_18015,N_18779);
xnor U19394 (N_19394,N_18432,N_18050);
and U19395 (N_19395,N_18083,N_18483);
or U19396 (N_19396,N_18067,N_18090);
nor U19397 (N_19397,N_18066,N_18606);
xor U19398 (N_19398,N_18373,N_18416);
and U19399 (N_19399,N_18185,N_18793);
and U19400 (N_19400,N_18096,N_18402);
nand U19401 (N_19401,N_18296,N_18801);
xnor U19402 (N_19402,N_18778,N_18862);
nor U19403 (N_19403,N_18991,N_18588);
nor U19404 (N_19404,N_18493,N_18774);
xnor U19405 (N_19405,N_18840,N_18316);
or U19406 (N_19406,N_18377,N_18002);
xor U19407 (N_19407,N_18507,N_18401);
nor U19408 (N_19408,N_18742,N_18112);
nor U19409 (N_19409,N_18511,N_18405);
nor U19410 (N_19410,N_18125,N_18356);
and U19411 (N_19411,N_18078,N_18055);
and U19412 (N_19412,N_18869,N_18147);
nor U19413 (N_19413,N_18660,N_18378);
nand U19414 (N_19414,N_18791,N_18195);
or U19415 (N_19415,N_18815,N_18972);
nand U19416 (N_19416,N_18669,N_18244);
nand U19417 (N_19417,N_18765,N_18608);
or U19418 (N_19418,N_18460,N_18031);
nand U19419 (N_19419,N_18834,N_18108);
nor U19420 (N_19420,N_18976,N_18786);
nor U19421 (N_19421,N_18188,N_18452);
nand U19422 (N_19422,N_18419,N_18757);
xnor U19423 (N_19423,N_18689,N_18211);
nor U19424 (N_19424,N_18395,N_18639);
nor U19425 (N_19425,N_18926,N_18731);
nand U19426 (N_19426,N_18442,N_18158);
nand U19427 (N_19427,N_18109,N_18974);
nand U19428 (N_19428,N_18975,N_18889);
xnor U19429 (N_19429,N_18827,N_18491);
nand U19430 (N_19430,N_18555,N_18590);
or U19431 (N_19431,N_18243,N_18737);
nand U19432 (N_19432,N_18874,N_18516);
or U19433 (N_19433,N_18191,N_18013);
xor U19434 (N_19434,N_18326,N_18314);
and U19435 (N_19435,N_18807,N_18135);
xor U19436 (N_19436,N_18022,N_18729);
and U19437 (N_19437,N_18549,N_18447);
nand U19438 (N_19438,N_18604,N_18338);
or U19439 (N_19439,N_18012,N_18376);
or U19440 (N_19440,N_18512,N_18463);
and U19441 (N_19441,N_18666,N_18345);
xor U19442 (N_19442,N_18832,N_18613);
xnor U19443 (N_19443,N_18640,N_18458);
nor U19444 (N_19444,N_18683,N_18935);
xor U19445 (N_19445,N_18885,N_18773);
and U19446 (N_19446,N_18914,N_18918);
or U19447 (N_19447,N_18332,N_18636);
xnor U19448 (N_19448,N_18222,N_18612);
or U19449 (N_19449,N_18775,N_18203);
xor U19450 (N_19450,N_18726,N_18811);
and U19451 (N_19451,N_18227,N_18039);
nor U19452 (N_19452,N_18537,N_18812);
nand U19453 (N_19453,N_18306,N_18905);
nor U19454 (N_19454,N_18391,N_18988);
and U19455 (N_19455,N_18337,N_18335);
nand U19456 (N_19456,N_18342,N_18708);
and U19457 (N_19457,N_18399,N_18220);
nor U19458 (N_19458,N_18901,N_18943);
or U19459 (N_19459,N_18649,N_18870);
xor U19460 (N_19460,N_18216,N_18662);
nor U19461 (N_19461,N_18900,N_18875);
nor U19462 (N_19462,N_18565,N_18830);
nand U19463 (N_19463,N_18256,N_18902);
nor U19464 (N_19464,N_18412,N_18328);
xnor U19465 (N_19465,N_18556,N_18580);
nand U19466 (N_19466,N_18124,N_18668);
nand U19467 (N_19467,N_18970,N_18531);
and U19468 (N_19468,N_18094,N_18624);
nand U19469 (N_19469,N_18996,N_18760);
xor U19470 (N_19470,N_18513,N_18392);
or U19471 (N_19471,N_18372,N_18196);
nand U19472 (N_19472,N_18871,N_18110);
xor U19473 (N_19473,N_18785,N_18390);
or U19474 (N_19474,N_18932,N_18303);
nor U19475 (N_19475,N_18508,N_18746);
and U19476 (N_19476,N_18441,N_18208);
nor U19477 (N_19477,N_18825,N_18806);
nand U19478 (N_19478,N_18101,N_18573);
and U19479 (N_19479,N_18745,N_18265);
or U19480 (N_19480,N_18747,N_18422);
or U19481 (N_19481,N_18838,N_18985);
xor U19482 (N_19482,N_18006,N_18696);
nand U19483 (N_19483,N_18118,N_18355);
nand U19484 (N_19484,N_18197,N_18311);
nand U19485 (N_19485,N_18456,N_18740);
xnor U19486 (N_19486,N_18058,N_18054);
nand U19487 (N_19487,N_18529,N_18753);
nor U19488 (N_19488,N_18810,N_18201);
nor U19489 (N_19489,N_18340,N_18921);
and U19490 (N_19490,N_18153,N_18989);
xor U19491 (N_19491,N_18715,N_18291);
and U19492 (N_19492,N_18808,N_18526);
or U19493 (N_19493,N_18687,N_18455);
xnor U19494 (N_19494,N_18029,N_18137);
xor U19495 (N_19495,N_18847,N_18347);
nor U19496 (N_19496,N_18795,N_18739);
or U19497 (N_19497,N_18766,N_18131);
and U19498 (N_19498,N_18720,N_18923);
xor U19499 (N_19499,N_18579,N_18418);
or U19500 (N_19500,N_18847,N_18288);
or U19501 (N_19501,N_18313,N_18116);
nor U19502 (N_19502,N_18717,N_18337);
and U19503 (N_19503,N_18824,N_18795);
or U19504 (N_19504,N_18585,N_18348);
nor U19505 (N_19505,N_18623,N_18323);
nand U19506 (N_19506,N_18602,N_18974);
nor U19507 (N_19507,N_18194,N_18862);
and U19508 (N_19508,N_18323,N_18645);
nand U19509 (N_19509,N_18876,N_18856);
and U19510 (N_19510,N_18956,N_18864);
and U19511 (N_19511,N_18625,N_18446);
and U19512 (N_19512,N_18478,N_18033);
nor U19513 (N_19513,N_18825,N_18182);
or U19514 (N_19514,N_18965,N_18031);
nand U19515 (N_19515,N_18000,N_18720);
nand U19516 (N_19516,N_18975,N_18712);
or U19517 (N_19517,N_18059,N_18480);
or U19518 (N_19518,N_18856,N_18817);
nor U19519 (N_19519,N_18722,N_18209);
nor U19520 (N_19520,N_18956,N_18730);
and U19521 (N_19521,N_18698,N_18712);
xor U19522 (N_19522,N_18409,N_18574);
and U19523 (N_19523,N_18913,N_18812);
nand U19524 (N_19524,N_18297,N_18934);
xor U19525 (N_19525,N_18707,N_18112);
xnor U19526 (N_19526,N_18908,N_18620);
xor U19527 (N_19527,N_18374,N_18780);
or U19528 (N_19528,N_18678,N_18216);
nand U19529 (N_19529,N_18530,N_18545);
nor U19530 (N_19530,N_18674,N_18451);
and U19531 (N_19531,N_18882,N_18121);
xnor U19532 (N_19532,N_18170,N_18433);
or U19533 (N_19533,N_18791,N_18258);
nand U19534 (N_19534,N_18520,N_18912);
nor U19535 (N_19535,N_18712,N_18696);
and U19536 (N_19536,N_18382,N_18621);
xnor U19537 (N_19537,N_18435,N_18290);
nor U19538 (N_19538,N_18747,N_18930);
and U19539 (N_19539,N_18204,N_18173);
and U19540 (N_19540,N_18590,N_18042);
nor U19541 (N_19541,N_18812,N_18085);
nor U19542 (N_19542,N_18547,N_18717);
xnor U19543 (N_19543,N_18785,N_18259);
nor U19544 (N_19544,N_18731,N_18105);
nand U19545 (N_19545,N_18559,N_18056);
nand U19546 (N_19546,N_18634,N_18592);
nor U19547 (N_19547,N_18430,N_18890);
and U19548 (N_19548,N_18734,N_18937);
or U19549 (N_19549,N_18940,N_18565);
xor U19550 (N_19550,N_18606,N_18169);
and U19551 (N_19551,N_18225,N_18581);
and U19552 (N_19552,N_18662,N_18160);
or U19553 (N_19553,N_18963,N_18768);
or U19554 (N_19554,N_18015,N_18990);
or U19555 (N_19555,N_18221,N_18704);
and U19556 (N_19556,N_18747,N_18430);
or U19557 (N_19557,N_18135,N_18714);
nand U19558 (N_19558,N_18646,N_18474);
and U19559 (N_19559,N_18461,N_18472);
nor U19560 (N_19560,N_18591,N_18861);
and U19561 (N_19561,N_18196,N_18644);
nand U19562 (N_19562,N_18805,N_18006);
nor U19563 (N_19563,N_18474,N_18722);
or U19564 (N_19564,N_18996,N_18269);
and U19565 (N_19565,N_18622,N_18889);
nor U19566 (N_19566,N_18181,N_18886);
nand U19567 (N_19567,N_18098,N_18066);
or U19568 (N_19568,N_18208,N_18830);
xnor U19569 (N_19569,N_18922,N_18779);
and U19570 (N_19570,N_18710,N_18818);
nand U19571 (N_19571,N_18154,N_18528);
or U19572 (N_19572,N_18140,N_18515);
nor U19573 (N_19573,N_18667,N_18755);
nor U19574 (N_19574,N_18727,N_18315);
nand U19575 (N_19575,N_18812,N_18389);
nor U19576 (N_19576,N_18291,N_18728);
nand U19577 (N_19577,N_18410,N_18939);
nor U19578 (N_19578,N_18037,N_18293);
nand U19579 (N_19579,N_18038,N_18234);
or U19580 (N_19580,N_18799,N_18296);
nand U19581 (N_19581,N_18977,N_18609);
nor U19582 (N_19582,N_18254,N_18119);
xnor U19583 (N_19583,N_18348,N_18024);
and U19584 (N_19584,N_18942,N_18946);
nor U19585 (N_19585,N_18921,N_18811);
nor U19586 (N_19586,N_18237,N_18355);
xor U19587 (N_19587,N_18667,N_18502);
or U19588 (N_19588,N_18006,N_18617);
or U19589 (N_19589,N_18259,N_18338);
nand U19590 (N_19590,N_18675,N_18522);
xnor U19591 (N_19591,N_18677,N_18364);
or U19592 (N_19592,N_18090,N_18692);
and U19593 (N_19593,N_18583,N_18370);
or U19594 (N_19594,N_18173,N_18991);
or U19595 (N_19595,N_18935,N_18982);
or U19596 (N_19596,N_18896,N_18814);
or U19597 (N_19597,N_18611,N_18141);
nand U19598 (N_19598,N_18676,N_18998);
and U19599 (N_19599,N_18130,N_18183);
nand U19600 (N_19600,N_18425,N_18392);
xor U19601 (N_19601,N_18799,N_18074);
or U19602 (N_19602,N_18107,N_18164);
and U19603 (N_19603,N_18924,N_18901);
and U19604 (N_19604,N_18982,N_18993);
nand U19605 (N_19605,N_18718,N_18736);
nand U19606 (N_19606,N_18424,N_18141);
xor U19607 (N_19607,N_18747,N_18538);
nor U19608 (N_19608,N_18760,N_18221);
and U19609 (N_19609,N_18952,N_18912);
and U19610 (N_19610,N_18374,N_18082);
and U19611 (N_19611,N_18011,N_18173);
nand U19612 (N_19612,N_18839,N_18805);
xnor U19613 (N_19613,N_18161,N_18850);
xnor U19614 (N_19614,N_18165,N_18524);
and U19615 (N_19615,N_18012,N_18839);
or U19616 (N_19616,N_18029,N_18273);
or U19617 (N_19617,N_18211,N_18678);
or U19618 (N_19618,N_18589,N_18433);
and U19619 (N_19619,N_18987,N_18126);
nor U19620 (N_19620,N_18745,N_18836);
nand U19621 (N_19621,N_18217,N_18837);
and U19622 (N_19622,N_18222,N_18444);
xor U19623 (N_19623,N_18306,N_18566);
xnor U19624 (N_19624,N_18911,N_18637);
nand U19625 (N_19625,N_18891,N_18621);
and U19626 (N_19626,N_18080,N_18860);
xnor U19627 (N_19627,N_18112,N_18004);
nor U19628 (N_19628,N_18145,N_18729);
nand U19629 (N_19629,N_18873,N_18859);
and U19630 (N_19630,N_18429,N_18822);
or U19631 (N_19631,N_18755,N_18959);
and U19632 (N_19632,N_18099,N_18622);
or U19633 (N_19633,N_18802,N_18319);
xor U19634 (N_19634,N_18736,N_18539);
nor U19635 (N_19635,N_18603,N_18324);
or U19636 (N_19636,N_18056,N_18344);
xor U19637 (N_19637,N_18048,N_18467);
nor U19638 (N_19638,N_18242,N_18158);
and U19639 (N_19639,N_18235,N_18936);
xnor U19640 (N_19640,N_18739,N_18109);
xor U19641 (N_19641,N_18202,N_18992);
and U19642 (N_19642,N_18759,N_18864);
xor U19643 (N_19643,N_18562,N_18821);
or U19644 (N_19644,N_18974,N_18440);
nand U19645 (N_19645,N_18481,N_18446);
xnor U19646 (N_19646,N_18939,N_18350);
and U19647 (N_19647,N_18825,N_18044);
and U19648 (N_19648,N_18879,N_18195);
and U19649 (N_19649,N_18510,N_18263);
nor U19650 (N_19650,N_18936,N_18798);
xnor U19651 (N_19651,N_18125,N_18470);
nand U19652 (N_19652,N_18518,N_18136);
nand U19653 (N_19653,N_18652,N_18378);
or U19654 (N_19654,N_18697,N_18227);
xnor U19655 (N_19655,N_18102,N_18340);
or U19656 (N_19656,N_18062,N_18646);
nor U19657 (N_19657,N_18048,N_18390);
xor U19658 (N_19658,N_18337,N_18834);
nor U19659 (N_19659,N_18104,N_18434);
nor U19660 (N_19660,N_18612,N_18931);
nor U19661 (N_19661,N_18791,N_18629);
nand U19662 (N_19662,N_18109,N_18362);
nand U19663 (N_19663,N_18236,N_18544);
and U19664 (N_19664,N_18669,N_18942);
or U19665 (N_19665,N_18700,N_18996);
nand U19666 (N_19666,N_18264,N_18796);
nor U19667 (N_19667,N_18344,N_18406);
nand U19668 (N_19668,N_18748,N_18052);
or U19669 (N_19669,N_18450,N_18624);
nor U19670 (N_19670,N_18021,N_18723);
nand U19671 (N_19671,N_18973,N_18786);
nand U19672 (N_19672,N_18442,N_18958);
nor U19673 (N_19673,N_18615,N_18228);
and U19674 (N_19674,N_18727,N_18687);
xor U19675 (N_19675,N_18287,N_18787);
or U19676 (N_19676,N_18599,N_18671);
and U19677 (N_19677,N_18882,N_18611);
xor U19678 (N_19678,N_18414,N_18389);
xor U19679 (N_19679,N_18940,N_18015);
nor U19680 (N_19680,N_18303,N_18826);
xor U19681 (N_19681,N_18507,N_18597);
xnor U19682 (N_19682,N_18932,N_18133);
or U19683 (N_19683,N_18500,N_18346);
xnor U19684 (N_19684,N_18505,N_18890);
nor U19685 (N_19685,N_18587,N_18422);
or U19686 (N_19686,N_18303,N_18371);
nor U19687 (N_19687,N_18912,N_18342);
or U19688 (N_19688,N_18076,N_18882);
nor U19689 (N_19689,N_18587,N_18501);
or U19690 (N_19690,N_18469,N_18917);
nor U19691 (N_19691,N_18766,N_18220);
nor U19692 (N_19692,N_18896,N_18410);
nand U19693 (N_19693,N_18392,N_18822);
xnor U19694 (N_19694,N_18921,N_18102);
or U19695 (N_19695,N_18087,N_18003);
nor U19696 (N_19696,N_18532,N_18117);
xnor U19697 (N_19697,N_18993,N_18335);
and U19698 (N_19698,N_18265,N_18161);
xor U19699 (N_19699,N_18958,N_18057);
or U19700 (N_19700,N_18273,N_18301);
and U19701 (N_19701,N_18157,N_18113);
and U19702 (N_19702,N_18971,N_18389);
nand U19703 (N_19703,N_18181,N_18096);
xor U19704 (N_19704,N_18898,N_18821);
xnor U19705 (N_19705,N_18870,N_18760);
xnor U19706 (N_19706,N_18514,N_18645);
nor U19707 (N_19707,N_18228,N_18065);
nor U19708 (N_19708,N_18419,N_18304);
or U19709 (N_19709,N_18122,N_18471);
nor U19710 (N_19710,N_18638,N_18356);
nand U19711 (N_19711,N_18454,N_18930);
or U19712 (N_19712,N_18952,N_18713);
nand U19713 (N_19713,N_18909,N_18695);
nand U19714 (N_19714,N_18173,N_18014);
xnor U19715 (N_19715,N_18143,N_18065);
nand U19716 (N_19716,N_18065,N_18704);
or U19717 (N_19717,N_18529,N_18760);
and U19718 (N_19718,N_18672,N_18374);
xnor U19719 (N_19719,N_18529,N_18228);
nor U19720 (N_19720,N_18521,N_18048);
and U19721 (N_19721,N_18547,N_18551);
or U19722 (N_19722,N_18649,N_18919);
xnor U19723 (N_19723,N_18734,N_18951);
nand U19724 (N_19724,N_18182,N_18620);
nand U19725 (N_19725,N_18539,N_18969);
or U19726 (N_19726,N_18576,N_18065);
xor U19727 (N_19727,N_18719,N_18511);
xor U19728 (N_19728,N_18286,N_18363);
xor U19729 (N_19729,N_18706,N_18967);
nor U19730 (N_19730,N_18253,N_18733);
nor U19731 (N_19731,N_18023,N_18245);
nand U19732 (N_19732,N_18965,N_18214);
nor U19733 (N_19733,N_18957,N_18557);
or U19734 (N_19734,N_18859,N_18224);
or U19735 (N_19735,N_18427,N_18922);
xor U19736 (N_19736,N_18502,N_18358);
nor U19737 (N_19737,N_18318,N_18116);
and U19738 (N_19738,N_18536,N_18050);
nor U19739 (N_19739,N_18791,N_18358);
nand U19740 (N_19740,N_18035,N_18789);
or U19741 (N_19741,N_18471,N_18399);
or U19742 (N_19742,N_18931,N_18587);
nor U19743 (N_19743,N_18944,N_18512);
and U19744 (N_19744,N_18702,N_18980);
or U19745 (N_19745,N_18113,N_18089);
nor U19746 (N_19746,N_18492,N_18716);
nor U19747 (N_19747,N_18439,N_18567);
and U19748 (N_19748,N_18174,N_18017);
and U19749 (N_19749,N_18407,N_18479);
nand U19750 (N_19750,N_18849,N_18903);
or U19751 (N_19751,N_18655,N_18406);
xnor U19752 (N_19752,N_18864,N_18925);
xnor U19753 (N_19753,N_18120,N_18384);
and U19754 (N_19754,N_18889,N_18240);
or U19755 (N_19755,N_18392,N_18972);
and U19756 (N_19756,N_18043,N_18533);
or U19757 (N_19757,N_18391,N_18359);
xor U19758 (N_19758,N_18065,N_18809);
xnor U19759 (N_19759,N_18222,N_18662);
and U19760 (N_19760,N_18859,N_18757);
nand U19761 (N_19761,N_18811,N_18252);
xnor U19762 (N_19762,N_18608,N_18152);
xnor U19763 (N_19763,N_18273,N_18807);
xor U19764 (N_19764,N_18154,N_18343);
nand U19765 (N_19765,N_18724,N_18363);
or U19766 (N_19766,N_18032,N_18159);
nand U19767 (N_19767,N_18963,N_18258);
nand U19768 (N_19768,N_18873,N_18638);
nor U19769 (N_19769,N_18068,N_18114);
or U19770 (N_19770,N_18951,N_18242);
nand U19771 (N_19771,N_18689,N_18858);
or U19772 (N_19772,N_18938,N_18108);
nand U19773 (N_19773,N_18223,N_18091);
nand U19774 (N_19774,N_18286,N_18470);
nand U19775 (N_19775,N_18404,N_18711);
or U19776 (N_19776,N_18556,N_18902);
xor U19777 (N_19777,N_18891,N_18747);
xor U19778 (N_19778,N_18890,N_18518);
xnor U19779 (N_19779,N_18254,N_18734);
nor U19780 (N_19780,N_18713,N_18432);
nand U19781 (N_19781,N_18227,N_18902);
nand U19782 (N_19782,N_18119,N_18271);
xnor U19783 (N_19783,N_18390,N_18912);
nor U19784 (N_19784,N_18680,N_18586);
or U19785 (N_19785,N_18264,N_18031);
xor U19786 (N_19786,N_18438,N_18218);
nand U19787 (N_19787,N_18203,N_18670);
or U19788 (N_19788,N_18252,N_18040);
nor U19789 (N_19789,N_18944,N_18743);
nor U19790 (N_19790,N_18149,N_18270);
nor U19791 (N_19791,N_18073,N_18871);
xor U19792 (N_19792,N_18497,N_18980);
or U19793 (N_19793,N_18618,N_18469);
and U19794 (N_19794,N_18002,N_18395);
xnor U19795 (N_19795,N_18955,N_18546);
nor U19796 (N_19796,N_18405,N_18533);
nor U19797 (N_19797,N_18107,N_18498);
or U19798 (N_19798,N_18248,N_18747);
nand U19799 (N_19799,N_18087,N_18223);
nand U19800 (N_19800,N_18046,N_18941);
or U19801 (N_19801,N_18423,N_18118);
and U19802 (N_19802,N_18183,N_18398);
or U19803 (N_19803,N_18213,N_18337);
nor U19804 (N_19804,N_18212,N_18501);
nand U19805 (N_19805,N_18089,N_18385);
and U19806 (N_19806,N_18003,N_18839);
or U19807 (N_19807,N_18277,N_18231);
xor U19808 (N_19808,N_18604,N_18983);
nor U19809 (N_19809,N_18683,N_18713);
or U19810 (N_19810,N_18146,N_18748);
nor U19811 (N_19811,N_18184,N_18853);
nand U19812 (N_19812,N_18215,N_18039);
nor U19813 (N_19813,N_18984,N_18606);
xor U19814 (N_19814,N_18836,N_18430);
and U19815 (N_19815,N_18410,N_18435);
or U19816 (N_19816,N_18536,N_18233);
and U19817 (N_19817,N_18744,N_18531);
nor U19818 (N_19818,N_18101,N_18368);
and U19819 (N_19819,N_18685,N_18459);
xnor U19820 (N_19820,N_18935,N_18290);
or U19821 (N_19821,N_18069,N_18673);
or U19822 (N_19822,N_18793,N_18273);
nor U19823 (N_19823,N_18952,N_18647);
nand U19824 (N_19824,N_18608,N_18549);
and U19825 (N_19825,N_18151,N_18886);
nor U19826 (N_19826,N_18377,N_18626);
nand U19827 (N_19827,N_18888,N_18196);
or U19828 (N_19828,N_18102,N_18044);
or U19829 (N_19829,N_18835,N_18509);
nand U19830 (N_19830,N_18117,N_18715);
or U19831 (N_19831,N_18012,N_18437);
xnor U19832 (N_19832,N_18072,N_18789);
nor U19833 (N_19833,N_18058,N_18338);
or U19834 (N_19834,N_18729,N_18455);
nand U19835 (N_19835,N_18121,N_18507);
nor U19836 (N_19836,N_18673,N_18732);
nand U19837 (N_19837,N_18864,N_18027);
xor U19838 (N_19838,N_18531,N_18899);
nor U19839 (N_19839,N_18666,N_18160);
nand U19840 (N_19840,N_18036,N_18214);
nor U19841 (N_19841,N_18007,N_18291);
and U19842 (N_19842,N_18415,N_18953);
and U19843 (N_19843,N_18579,N_18352);
xor U19844 (N_19844,N_18874,N_18093);
or U19845 (N_19845,N_18256,N_18799);
and U19846 (N_19846,N_18558,N_18108);
and U19847 (N_19847,N_18025,N_18752);
nor U19848 (N_19848,N_18116,N_18587);
or U19849 (N_19849,N_18817,N_18204);
or U19850 (N_19850,N_18977,N_18676);
nand U19851 (N_19851,N_18890,N_18892);
xor U19852 (N_19852,N_18858,N_18315);
nand U19853 (N_19853,N_18455,N_18618);
nor U19854 (N_19854,N_18144,N_18696);
and U19855 (N_19855,N_18699,N_18250);
or U19856 (N_19856,N_18265,N_18543);
nand U19857 (N_19857,N_18027,N_18015);
nor U19858 (N_19858,N_18856,N_18007);
nand U19859 (N_19859,N_18519,N_18628);
and U19860 (N_19860,N_18835,N_18189);
or U19861 (N_19861,N_18670,N_18773);
nand U19862 (N_19862,N_18013,N_18238);
and U19863 (N_19863,N_18392,N_18127);
and U19864 (N_19864,N_18392,N_18064);
nor U19865 (N_19865,N_18120,N_18043);
or U19866 (N_19866,N_18347,N_18382);
or U19867 (N_19867,N_18771,N_18802);
nand U19868 (N_19868,N_18663,N_18656);
xor U19869 (N_19869,N_18366,N_18421);
nand U19870 (N_19870,N_18779,N_18633);
nand U19871 (N_19871,N_18534,N_18466);
nand U19872 (N_19872,N_18843,N_18707);
or U19873 (N_19873,N_18120,N_18988);
nor U19874 (N_19874,N_18642,N_18943);
and U19875 (N_19875,N_18788,N_18965);
or U19876 (N_19876,N_18793,N_18987);
xnor U19877 (N_19877,N_18956,N_18447);
nand U19878 (N_19878,N_18649,N_18754);
or U19879 (N_19879,N_18292,N_18595);
nor U19880 (N_19880,N_18028,N_18699);
and U19881 (N_19881,N_18087,N_18394);
nor U19882 (N_19882,N_18651,N_18477);
nand U19883 (N_19883,N_18705,N_18447);
nand U19884 (N_19884,N_18058,N_18766);
or U19885 (N_19885,N_18985,N_18867);
and U19886 (N_19886,N_18196,N_18862);
and U19887 (N_19887,N_18145,N_18208);
xor U19888 (N_19888,N_18442,N_18951);
and U19889 (N_19889,N_18517,N_18833);
nor U19890 (N_19890,N_18672,N_18091);
and U19891 (N_19891,N_18447,N_18344);
nor U19892 (N_19892,N_18933,N_18980);
nor U19893 (N_19893,N_18120,N_18109);
and U19894 (N_19894,N_18988,N_18486);
nand U19895 (N_19895,N_18137,N_18422);
nor U19896 (N_19896,N_18185,N_18012);
nor U19897 (N_19897,N_18632,N_18339);
xnor U19898 (N_19898,N_18306,N_18887);
and U19899 (N_19899,N_18535,N_18699);
xor U19900 (N_19900,N_18089,N_18721);
nor U19901 (N_19901,N_18784,N_18970);
and U19902 (N_19902,N_18325,N_18227);
nor U19903 (N_19903,N_18368,N_18518);
xor U19904 (N_19904,N_18753,N_18008);
nor U19905 (N_19905,N_18679,N_18934);
and U19906 (N_19906,N_18666,N_18952);
and U19907 (N_19907,N_18289,N_18018);
nand U19908 (N_19908,N_18157,N_18986);
and U19909 (N_19909,N_18755,N_18518);
nand U19910 (N_19910,N_18907,N_18918);
and U19911 (N_19911,N_18169,N_18394);
xor U19912 (N_19912,N_18840,N_18564);
or U19913 (N_19913,N_18957,N_18198);
nand U19914 (N_19914,N_18481,N_18347);
xnor U19915 (N_19915,N_18057,N_18309);
nand U19916 (N_19916,N_18396,N_18454);
or U19917 (N_19917,N_18785,N_18379);
or U19918 (N_19918,N_18521,N_18530);
nor U19919 (N_19919,N_18432,N_18624);
nor U19920 (N_19920,N_18476,N_18473);
nand U19921 (N_19921,N_18418,N_18530);
and U19922 (N_19922,N_18393,N_18023);
xor U19923 (N_19923,N_18887,N_18689);
xor U19924 (N_19924,N_18060,N_18891);
nand U19925 (N_19925,N_18049,N_18513);
or U19926 (N_19926,N_18552,N_18853);
nand U19927 (N_19927,N_18509,N_18786);
or U19928 (N_19928,N_18796,N_18503);
nor U19929 (N_19929,N_18020,N_18750);
nand U19930 (N_19930,N_18181,N_18089);
nand U19931 (N_19931,N_18277,N_18934);
nor U19932 (N_19932,N_18859,N_18849);
or U19933 (N_19933,N_18664,N_18681);
nand U19934 (N_19934,N_18054,N_18777);
or U19935 (N_19935,N_18866,N_18005);
and U19936 (N_19936,N_18932,N_18118);
or U19937 (N_19937,N_18065,N_18078);
and U19938 (N_19938,N_18666,N_18793);
and U19939 (N_19939,N_18386,N_18421);
and U19940 (N_19940,N_18525,N_18523);
nor U19941 (N_19941,N_18492,N_18991);
nor U19942 (N_19942,N_18802,N_18515);
xnor U19943 (N_19943,N_18749,N_18824);
xor U19944 (N_19944,N_18453,N_18821);
nor U19945 (N_19945,N_18649,N_18314);
nand U19946 (N_19946,N_18573,N_18315);
and U19947 (N_19947,N_18678,N_18194);
nand U19948 (N_19948,N_18060,N_18319);
nor U19949 (N_19949,N_18244,N_18226);
xnor U19950 (N_19950,N_18910,N_18727);
nand U19951 (N_19951,N_18322,N_18104);
nor U19952 (N_19952,N_18946,N_18618);
xor U19953 (N_19953,N_18558,N_18093);
xor U19954 (N_19954,N_18354,N_18636);
and U19955 (N_19955,N_18077,N_18236);
or U19956 (N_19956,N_18949,N_18147);
nor U19957 (N_19957,N_18412,N_18213);
and U19958 (N_19958,N_18187,N_18215);
and U19959 (N_19959,N_18801,N_18116);
xnor U19960 (N_19960,N_18849,N_18496);
xnor U19961 (N_19961,N_18458,N_18833);
or U19962 (N_19962,N_18910,N_18591);
nand U19963 (N_19963,N_18390,N_18383);
and U19964 (N_19964,N_18297,N_18362);
xnor U19965 (N_19965,N_18611,N_18554);
nor U19966 (N_19966,N_18054,N_18003);
and U19967 (N_19967,N_18832,N_18339);
nor U19968 (N_19968,N_18836,N_18422);
nor U19969 (N_19969,N_18515,N_18167);
or U19970 (N_19970,N_18203,N_18472);
xor U19971 (N_19971,N_18415,N_18128);
and U19972 (N_19972,N_18701,N_18366);
nor U19973 (N_19973,N_18118,N_18154);
nand U19974 (N_19974,N_18917,N_18993);
and U19975 (N_19975,N_18820,N_18165);
and U19976 (N_19976,N_18833,N_18799);
xnor U19977 (N_19977,N_18876,N_18800);
nor U19978 (N_19978,N_18737,N_18506);
xnor U19979 (N_19979,N_18585,N_18173);
xor U19980 (N_19980,N_18926,N_18925);
nor U19981 (N_19981,N_18795,N_18374);
nor U19982 (N_19982,N_18223,N_18615);
and U19983 (N_19983,N_18601,N_18918);
xor U19984 (N_19984,N_18630,N_18373);
or U19985 (N_19985,N_18848,N_18116);
xnor U19986 (N_19986,N_18738,N_18485);
nand U19987 (N_19987,N_18208,N_18204);
and U19988 (N_19988,N_18774,N_18849);
and U19989 (N_19989,N_18959,N_18279);
and U19990 (N_19990,N_18802,N_18005);
nand U19991 (N_19991,N_18083,N_18601);
nand U19992 (N_19992,N_18087,N_18190);
or U19993 (N_19993,N_18234,N_18770);
nor U19994 (N_19994,N_18228,N_18896);
nor U19995 (N_19995,N_18636,N_18213);
xor U19996 (N_19996,N_18626,N_18643);
nand U19997 (N_19997,N_18110,N_18517);
or U19998 (N_19998,N_18052,N_18248);
xor U19999 (N_19999,N_18243,N_18766);
nor U20000 (N_20000,N_19993,N_19388);
xor U20001 (N_20001,N_19689,N_19159);
nand U20002 (N_20002,N_19705,N_19646);
nand U20003 (N_20003,N_19264,N_19868);
nor U20004 (N_20004,N_19593,N_19673);
nand U20005 (N_20005,N_19751,N_19873);
nor U20006 (N_20006,N_19354,N_19639);
nor U20007 (N_20007,N_19475,N_19203);
xnor U20008 (N_20008,N_19502,N_19206);
or U20009 (N_20009,N_19349,N_19329);
and U20010 (N_20010,N_19557,N_19843);
nor U20011 (N_20011,N_19890,N_19205);
nand U20012 (N_20012,N_19902,N_19411);
xor U20013 (N_20013,N_19005,N_19066);
and U20014 (N_20014,N_19883,N_19587);
and U20015 (N_20015,N_19169,N_19439);
or U20016 (N_20016,N_19261,N_19103);
nor U20017 (N_20017,N_19207,N_19848);
nor U20018 (N_20018,N_19758,N_19013);
nor U20019 (N_20019,N_19684,N_19432);
xor U20020 (N_20020,N_19394,N_19938);
xor U20021 (N_20021,N_19399,N_19567);
nor U20022 (N_20022,N_19006,N_19841);
and U20023 (N_20023,N_19197,N_19281);
or U20024 (N_20024,N_19359,N_19213);
xnor U20025 (N_20025,N_19139,N_19970);
and U20026 (N_20026,N_19348,N_19721);
nand U20027 (N_20027,N_19484,N_19398);
xnor U20028 (N_20028,N_19680,N_19371);
nand U20029 (N_20029,N_19230,N_19645);
and U20030 (N_20030,N_19161,N_19940);
xnor U20031 (N_20031,N_19373,N_19086);
xor U20032 (N_20032,N_19518,N_19154);
or U20033 (N_20033,N_19947,N_19494);
nor U20034 (N_20034,N_19421,N_19919);
or U20035 (N_20035,N_19107,N_19943);
xor U20036 (N_20036,N_19468,N_19910);
xor U20037 (N_20037,N_19333,N_19315);
xor U20038 (N_20038,N_19761,N_19956);
xnor U20039 (N_20039,N_19276,N_19483);
and U20040 (N_20040,N_19142,N_19922);
and U20041 (N_20041,N_19621,N_19093);
xnor U20042 (N_20042,N_19355,N_19460);
nand U20043 (N_20043,N_19814,N_19457);
xor U20044 (N_20044,N_19434,N_19323);
nand U20045 (N_20045,N_19630,N_19260);
or U20046 (N_20046,N_19897,N_19955);
and U20047 (N_20047,N_19099,N_19743);
xor U20048 (N_20048,N_19528,N_19782);
xor U20049 (N_20049,N_19941,N_19072);
nand U20050 (N_20050,N_19239,N_19974);
xor U20051 (N_20051,N_19458,N_19643);
xnor U20052 (N_20052,N_19773,N_19456);
nor U20053 (N_20053,N_19280,N_19998);
and U20054 (N_20054,N_19662,N_19225);
nand U20055 (N_20055,N_19004,N_19561);
xor U20056 (N_20056,N_19619,N_19585);
or U20057 (N_20057,N_19384,N_19414);
or U20058 (N_20058,N_19083,N_19760);
nor U20059 (N_20059,N_19454,N_19248);
or U20060 (N_20060,N_19081,N_19061);
and U20061 (N_20061,N_19918,N_19606);
and U20062 (N_20062,N_19803,N_19003);
xnor U20063 (N_20063,N_19025,N_19641);
or U20064 (N_20064,N_19604,N_19199);
or U20065 (N_20065,N_19889,N_19599);
and U20066 (N_20066,N_19701,N_19982);
nand U20067 (N_20067,N_19032,N_19617);
xnor U20068 (N_20068,N_19298,N_19827);
xnor U20069 (N_20069,N_19470,N_19235);
and U20070 (N_20070,N_19908,N_19163);
and U20071 (N_20071,N_19968,N_19234);
xnor U20072 (N_20072,N_19117,N_19926);
nor U20073 (N_20073,N_19609,N_19045);
or U20074 (N_20074,N_19605,N_19710);
nor U20075 (N_20075,N_19148,N_19815);
nor U20076 (N_20076,N_19226,N_19444);
or U20077 (N_20077,N_19435,N_19440);
nand U20078 (N_20078,N_19591,N_19211);
nor U20079 (N_20079,N_19765,N_19912);
or U20080 (N_20080,N_19129,N_19736);
xor U20081 (N_20081,N_19627,N_19964);
nor U20082 (N_20082,N_19876,N_19101);
and U20083 (N_20083,N_19907,N_19364);
xor U20084 (N_20084,N_19324,N_19675);
nor U20085 (N_20085,N_19429,N_19186);
or U20086 (N_20086,N_19629,N_19582);
and U20087 (N_20087,N_19789,N_19709);
or U20088 (N_20088,N_19951,N_19997);
nor U20089 (N_20089,N_19408,N_19790);
and U20090 (N_20090,N_19492,N_19122);
or U20091 (N_20091,N_19866,N_19877);
and U20092 (N_20092,N_19430,N_19506);
or U20093 (N_20093,N_19427,N_19724);
or U20094 (N_20094,N_19375,N_19043);
xor U20095 (N_20095,N_19389,N_19610);
and U20096 (N_20096,N_19425,N_19836);
or U20097 (N_20097,N_19089,N_19450);
xnor U20098 (N_20098,N_19929,N_19923);
and U20099 (N_20099,N_19381,N_19644);
nor U20100 (N_20100,N_19949,N_19720);
or U20101 (N_20101,N_19719,N_19742);
nand U20102 (N_20102,N_19880,N_19633);
nand U20103 (N_20103,N_19774,N_19026);
nor U20104 (N_20104,N_19672,N_19537);
nor U20105 (N_20105,N_19763,N_19040);
and U20106 (N_20106,N_19337,N_19366);
nor U20107 (N_20107,N_19553,N_19330);
or U20108 (N_20108,N_19068,N_19054);
nand U20109 (N_20109,N_19698,N_19124);
nand U20110 (N_20110,N_19303,N_19471);
xor U20111 (N_20111,N_19541,N_19138);
xor U20112 (N_20112,N_19438,N_19077);
nand U20113 (N_20113,N_19634,N_19856);
nor U20114 (N_20114,N_19747,N_19130);
or U20115 (N_20115,N_19070,N_19224);
nand U20116 (N_20116,N_19284,N_19635);
nor U20117 (N_20117,N_19175,N_19624);
nor U20118 (N_20118,N_19022,N_19740);
or U20119 (N_20119,N_19344,N_19573);
and U20120 (N_20120,N_19016,N_19608);
or U20121 (N_20121,N_19356,N_19534);
xnor U20122 (N_20122,N_19150,N_19896);
nor U20123 (N_20123,N_19063,N_19002);
and U20124 (N_20124,N_19125,N_19056);
nand U20125 (N_20125,N_19691,N_19478);
nand U20126 (N_20126,N_19447,N_19249);
and U20127 (N_20127,N_19479,N_19113);
nand U20128 (N_20128,N_19404,N_19813);
nand U20129 (N_20129,N_19808,N_19036);
or U20130 (N_20130,N_19166,N_19283);
nor U20131 (N_20131,N_19328,N_19946);
nand U20132 (N_20132,N_19227,N_19852);
and U20133 (N_20133,N_19788,N_19273);
nor U20134 (N_20134,N_19603,N_19526);
xnor U20135 (N_20135,N_19115,N_19589);
or U20136 (N_20136,N_19892,N_19800);
or U20137 (N_20137,N_19011,N_19271);
or U20138 (N_20138,N_19551,N_19885);
or U20139 (N_20139,N_19702,N_19165);
xor U20140 (N_20140,N_19326,N_19776);
and U20141 (N_20141,N_19795,N_19485);
or U20142 (N_20142,N_19441,N_19893);
xor U20143 (N_20143,N_19809,N_19141);
and U20144 (N_20144,N_19764,N_19727);
nor U20145 (N_20145,N_19669,N_19676);
xnor U20146 (N_20146,N_19677,N_19382);
xnor U20147 (N_20147,N_19204,N_19697);
or U20148 (N_20148,N_19527,N_19029);
nand U20149 (N_20149,N_19516,N_19924);
or U20150 (N_20150,N_19978,N_19168);
nand U20151 (N_20151,N_19110,N_19493);
and U20152 (N_20152,N_19623,N_19647);
nor U20153 (N_20153,N_19810,N_19772);
nand U20154 (N_20154,N_19167,N_19096);
xnor U20155 (N_20155,N_19078,N_19508);
xnor U20156 (N_20156,N_19878,N_19732);
or U20157 (N_20157,N_19863,N_19402);
and U20158 (N_20158,N_19396,N_19542);
or U20159 (N_20159,N_19729,N_19085);
or U20160 (N_20160,N_19855,N_19419);
and U20161 (N_20161,N_19445,N_19500);
nand U20162 (N_20162,N_19285,N_19833);
or U20163 (N_20163,N_19847,N_19395);
or U20164 (N_20164,N_19505,N_19074);
nand U20165 (N_20165,N_19321,N_19681);
xnor U20166 (N_20166,N_19958,N_19174);
nand U20167 (N_20167,N_19361,N_19256);
and U20168 (N_20168,N_19839,N_19812);
nand U20169 (N_20169,N_19584,N_19400);
xor U20170 (N_20170,N_19980,N_19509);
or U20171 (N_20171,N_19291,N_19640);
nand U20172 (N_20172,N_19874,N_19424);
nand U20173 (N_20173,N_19659,N_19648);
nand U20174 (N_20174,N_19631,N_19496);
xor U20175 (N_20175,N_19318,N_19614);
nor U20176 (N_20176,N_19601,N_19416);
and U20177 (N_20177,N_19871,N_19247);
nand U20178 (N_20178,N_19210,N_19936);
or U20179 (N_20179,N_19901,N_19904);
and U20180 (N_20180,N_19133,N_19297);
nor U20181 (N_20181,N_19854,N_19305);
nand U20182 (N_20182,N_19486,N_19274);
and U20183 (N_20183,N_19977,N_19934);
xnor U20184 (N_20184,N_19804,N_19383);
xnor U20185 (N_20185,N_19781,N_19965);
or U20186 (N_20186,N_19762,N_19718);
or U20187 (N_20187,N_19825,N_19626);
nor U20188 (N_20188,N_19988,N_19132);
xnor U20189 (N_20189,N_19925,N_19933);
nand U20190 (N_20190,N_19898,N_19149);
and U20191 (N_20191,N_19018,N_19872);
nand U20192 (N_20192,N_19030,N_19531);
xor U20193 (N_20193,N_19302,N_19869);
xnor U20194 (N_20194,N_19008,N_19620);
nand U20195 (N_20195,N_19467,N_19272);
and U20196 (N_20196,N_19953,N_19538);
nor U20197 (N_20197,N_19688,N_19309);
nor U20198 (N_20198,N_19222,N_19613);
and U20199 (N_20199,N_19819,N_19463);
nor U20200 (N_20200,N_19187,N_19637);
or U20201 (N_20201,N_19112,N_19816);
xnor U20202 (N_20202,N_19410,N_19237);
or U20203 (N_20203,N_19409,N_19906);
or U20204 (N_20204,N_19325,N_19192);
and U20205 (N_20205,N_19094,N_19595);
nor U20206 (N_20206,N_19015,N_19491);
xnor U20207 (N_20207,N_19654,N_19202);
and U20208 (N_20208,N_19277,N_19306);
xor U20209 (N_20209,N_19164,N_19838);
and U20210 (N_20210,N_19658,N_19525);
and U20211 (N_20211,N_19236,N_19657);
or U20212 (N_20212,N_19307,N_19067);
nand U20213 (N_20213,N_19785,N_19973);
nor U20214 (N_20214,N_19162,N_19504);
and U20215 (N_20215,N_19991,N_19488);
nand U20216 (N_20216,N_19048,N_19310);
xor U20217 (N_20217,N_19944,N_19377);
and U20218 (N_20218,N_19487,N_19461);
nor U20219 (N_20219,N_19822,N_19905);
nor U20220 (N_20220,N_19135,N_19232);
and U20221 (N_20221,N_19752,N_19423);
nand U20222 (N_20222,N_19278,N_19250);
or U20223 (N_20223,N_19353,N_19246);
and U20224 (N_20224,N_19136,N_19108);
xnor U20225 (N_20225,N_19615,N_19792);
xor U20226 (N_20226,N_19095,N_19313);
and U20227 (N_20227,N_19652,N_19731);
xor U20228 (N_20228,N_19805,N_19547);
nand U20229 (N_20229,N_19798,N_19565);
or U20230 (N_20230,N_19577,N_19569);
xnor U20231 (N_20231,N_19268,N_19472);
nor U20232 (N_20232,N_19343,N_19228);
nand U20233 (N_20233,N_19661,N_19055);
xor U20234 (N_20234,N_19365,N_19442);
and U20235 (N_20235,N_19000,N_19049);
and U20236 (N_20236,N_19734,N_19220);
xor U20237 (N_20237,N_19091,N_19368);
or U20238 (N_20238,N_19759,N_19052);
and U20239 (N_20239,N_19594,N_19288);
and U20240 (N_20240,N_19571,N_19564);
and U20241 (N_20241,N_19830,N_19338);
xnor U20242 (N_20242,N_19510,N_19104);
nand U20243 (N_20243,N_19862,N_19127);
nand U20244 (N_20244,N_19304,N_19495);
and U20245 (N_20245,N_19548,N_19158);
or U20246 (N_20246,N_19448,N_19826);
or U20247 (N_20247,N_19481,N_19215);
xnor U20248 (N_20248,N_19179,N_19153);
nand U20249 (N_20249,N_19121,N_19791);
xor U20250 (N_20250,N_19722,N_19357);
xnor U20251 (N_20251,N_19392,N_19331);
or U20252 (N_20252,N_19476,N_19524);
or U20253 (N_20253,N_19437,N_19563);
nor U20254 (N_20254,N_19556,N_19027);
nand U20255 (N_20255,N_19433,N_19144);
or U20256 (N_20256,N_19327,N_19196);
nand U20257 (N_20257,N_19935,N_19738);
xor U20258 (N_20258,N_19649,N_19317);
xor U20259 (N_20259,N_19831,N_19216);
and U20260 (N_20260,N_19775,N_19928);
nor U20261 (N_20261,N_19820,N_19363);
or U20262 (N_20262,N_19231,N_19021);
or U20263 (N_20263,N_19536,N_19540);
and U20264 (N_20264,N_19378,N_19058);
xnor U20265 (N_20265,N_19581,N_19976);
or U20266 (N_20266,N_19501,N_19984);
and U20267 (N_20267,N_19693,N_19844);
xnor U20268 (N_20268,N_19916,N_19969);
nor U20269 (N_20269,N_19320,N_19017);
nand U20270 (N_20270,N_19157,N_19807);
xnor U20271 (N_20271,N_19939,N_19031);
or U20272 (N_20272,N_19257,N_19300);
nand U20273 (N_20273,N_19181,N_19683);
nor U20274 (N_20274,N_19019,N_19670);
or U20275 (N_20275,N_19687,N_19219);
or U20276 (N_20276,N_19996,N_19900);
or U20277 (N_20277,N_19459,N_19466);
xor U20278 (N_20278,N_19369,N_19778);
and U20279 (N_20279,N_19725,N_19097);
nor U20280 (N_20280,N_19682,N_19728);
nor U20281 (N_20281,N_19137,N_19412);
nand U20282 (N_20282,N_19241,N_19704);
and U20283 (N_20283,N_19694,N_19299);
nand U20284 (N_20284,N_19490,N_19663);
nand U20285 (N_20285,N_19927,N_19037);
xnor U20286 (N_20286,N_19262,N_19376);
or U20287 (N_20287,N_19265,N_19979);
xor U20288 (N_20288,N_19064,N_19543);
or U20289 (N_20289,N_19692,N_19514);
and U20290 (N_20290,N_19263,N_19134);
xor U20291 (N_20291,N_19178,N_19428);
nor U20292 (N_20292,N_19678,N_19143);
and U20293 (N_20293,N_19746,N_19797);
nand U20294 (N_20294,N_19963,N_19931);
nand U20295 (N_20295,N_19651,N_19082);
and U20296 (N_20296,N_19990,N_19886);
nor U20297 (N_20297,N_19799,N_19832);
xnor U20298 (N_20298,N_19041,N_19566);
and U20299 (N_20299,N_19749,N_19850);
nand U20300 (N_20300,N_19279,N_19884);
xor U20301 (N_20301,N_19152,N_19867);
and U20302 (N_20302,N_19674,N_19576);
nor U20303 (N_20303,N_19989,N_19242);
nand U20304 (N_20304,N_19699,N_19555);
or U20305 (N_20305,N_19287,N_19301);
nor U20306 (N_20306,N_19560,N_19597);
or U20307 (N_20307,N_19726,N_19986);
and U20308 (N_20308,N_19828,N_19332);
nand U20309 (N_20309,N_19190,N_19861);
xnor U20310 (N_20310,N_19511,N_19628);
and U20311 (N_20311,N_19817,N_19123);
xnor U20312 (N_20312,N_19787,N_19497);
or U20313 (N_20313,N_19942,N_19069);
and U20314 (N_20314,N_19367,N_19253);
and U20315 (N_20315,N_19917,N_19853);
xor U20316 (N_20316,N_19572,N_19347);
nand U20317 (N_20317,N_19351,N_19529);
or U20318 (N_20318,N_19223,N_19849);
nor U20319 (N_20319,N_19530,N_19611);
xnor U20320 (N_20320,N_19712,N_19308);
or U20321 (N_20321,N_19888,N_19258);
xor U20322 (N_20322,N_19735,N_19962);
nor U20323 (N_20323,N_19930,N_19730);
and U20324 (N_20324,N_19360,N_19858);
or U20325 (N_20325,N_19600,N_19811);
or U20326 (N_20326,N_19171,N_19744);
and U20327 (N_20327,N_19446,N_19464);
xnor U20328 (N_20328,N_19784,N_19051);
and U20329 (N_20329,N_19960,N_19859);
nand U20330 (N_20330,N_19075,N_19345);
nand U20331 (N_20331,N_19499,N_19715);
xnor U20332 (N_20332,N_19950,N_19339);
and U20333 (N_20333,N_19616,N_19894);
nor U20334 (N_20334,N_19767,N_19293);
and U20335 (N_20335,N_19887,N_19296);
or U20336 (N_20336,N_19046,N_19334);
nand U20337 (N_20337,N_19212,N_19106);
nor U20338 (N_20338,N_19275,N_19546);
nor U20339 (N_20339,N_19198,N_19975);
nor U20340 (N_20340,N_19050,N_19602);
or U20341 (N_20341,N_19452,N_19145);
nand U20342 (N_20342,N_19568,N_19266);
xnor U20343 (N_20343,N_19469,N_19177);
xnor U20344 (N_20344,N_19578,N_19292);
or U20345 (N_20345,N_19407,N_19370);
and U20346 (N_20346,N_19882,N_19057);
and U20347 (N_20347,N_19182,N_19282);
nor U20348 (N_20348,N_19455,N_19387);
nand U20349 (N_20349,N_19380,N_19655);
nand U20350 (N_20350,N_19985,N_19480);
nand U20351 (N_20351,N_19717,N_19632);
xnor U20352 (N_20352,N_19519,N_19155);
xnor U20353 (N_20353,N_19131,N_19286);
nand U20354 (N_20354,N_19522,N_19422);
nor U20355 (N_20355,N_19176,N_19405);
nand U20356 (N_20356,N_19482,N_19341);
xor U20357 (N_20357,N_19753,N_19267);
or U20358 (N_20358,N_19214,N_19544);
nand U20359 (N_20359,N_19517,N_19120);
and U20360 (N_20360,N_19802,N_19417);
nor U20361 (N_20361,N_19583,N_19660);
nand U20362 (N_20362,N_19851,N_19834);
nor U20363 (N_20363,N_19769,N_19243);
or U20364 (N_20364,N_19562,N_19636);
xor U20365 (N_20365,N_19653,N_19350);
nand U20366 (N_20366,N_19770,N_19346);
nor U20367 (N_20367,N_19044,N_19754);
xnor U20368 (N_20368,N_19590,N_19579);
xnor U20369 (N_20369,N_19489,N_19570);
nor U20370 (N_20370,N_19116,N_19290);
xor U20371 (N_20371,N_19756,N_19172);
nor U20372 (N_20372,N_19695,N_19513);
or U20373 (N_20373,N_19671,N_19431);
nand U20374 (N_20374,N_19014,N_19160);
nor U20375 (N_20375,N_19462,N_19845);
nor U20376 (N_20376,N_19385,N_19532);
nor U20377 (N_20377,N_19667,N_19098);
nand U20378 (N_20378,N_19716,N_19118);
nor U20379 (N_20379,N_19294,N_19793);
xnor U20380 (N_20380,N_19474,N_19959);
nor U20381 (N_20381,N_19062,N_19737);
and U20382 (N_20382,N_19588,N_19685);
nor U20383 (N_20383,N_19386,N_19195);
and U20384 (N_20384,N_19316,N_19857);
or U20385 (N_20385,N_19146,N_19105);
or U20386 (N_20386,N_19102,N_19352);
or U20387 (N_20387,N_19038,N_19768);
xnor U20388 (N_20388,N_19393,N_19358);
xor U20389 (N_20389,N_19552,N_19750);
nand U20390 (N_20390,N_19700,N_19766);
and U20391 (N_20391,N_19690,N_19270);
nor U20392 (N_20392,N_19259,N_19783);
xor U20393 (N_20393,N_19507,N_19042);
nor U20394 (N_20394,N_19140,N_19967);
nand U20395 (N_20395,N_19913,N_19390);
nor U20396 (N_20396,N_19100,N_19686);
or U20397 (N_20397,N_19846,N_19379);
xor U20398 (N_20398,N_19001,N_19992);
nand U20399 (N_20399,N_19840,N_19209);
nor U20400 (N_20400,N_19995,N_19443);
xnor U20401 (N_20401,N_19703,N_19771);
or U20402 (N_20402,N_19708,N_19920);
nand U20403 (N_20403,N_19777,N_19033);
xor U20404 (N_20404,N_19954,N_19948);
or U20405 (N_20405,N_19665,N_19295);
nor U20406 (N_20406,N_19696,N_19932);
and U20407 (N_20407,N_19679,N_19073);
nand U20408 (N_20408,N_19666,N_19523);
and U20409 (N_20409,N_19521,N_19244);
nand U20410 (N_20410,N_19245,N_19255);
xnor U20411 (N_20411,N_19047,N_19193);
and U20412 (N_20412,N_19739,N_19945);
nand U20413 (N_20413,N_19084,N_19558);
nand U20414 (N_20414,N_19554,N_19007);
or U20415 (N_20415,N_19983,N_19028);
nor U20416 (N_20416,N_19269,N_19184);
nand U20417 (N_20417,N_19335,N_19966);
nand U20418 (N_20418,N_19312,N_19533);
nor U20419 (N_20419,N_19638,N_19080);
or U20420 (N_20420,N_19012,N_19994);
and U20421 (N_20421,N_19860,N_19706);
and U20422 (N_20422,N_19053,N_19575);
nor U20423 (N_20423,N_19217,N_19961);
or U20424 (N_20424,N_19451,N_19559);
nand U20425 (N_20425,N_19915,N_19806);
or U20426 (N_20426,N_19034,N_19612);
nand U20427 (N_20427,N_19188,N_19909);
nor U20428 (N_20428,N_19233,N_19254);
and U20429 (N_20429,N_19823,N_19596);
and U20430 (N_20430,N_19707,N_19126);
and U20431 (N_20431,N_19401,N_19170);
xnor U20432 (N_20432,N_19023,N_19189);
xnor U20433 (N_20433,N_19650,N_19515);
or U20434 (N_20434,N_19342,N_19173);
nor U20435 (N_20435,N_19914,N_19201);
xnor U20436 (N_20436,N_19087,N_19111);
nand U20437 (N_20437,N_19088,N_19837);
xor U20438 (N_20438,N_19218,N_19473);
and U20439 (N_20439,N_19336,N_19039);
nand U20440 (N_20440,N_19311,N_19420);
and U20441 (N_20441,N_19981,N_19714);
or U20442 (N_20442,N_19194,N_19539);
xor U20443 (N_20443,N_19374,N_19545);
and U20444 (N_20444,N_19314,N_19128);
nand U20445 (N_20445,N_19911,N_19745);
xor U20446 (N_20446,N_19971,N_19191);
and U20447 (N_20447,N_19957,N_19656);
and U20448 (N_20448,N_19065,N_19748);
or U20449 (N_20449,N_19875,N_19151);
or U20450 (N_20450,N_19397,N_19801);
xnor U20451 (N_20451,N_19972,N_19780);
or U20452 (N_20452,N_19208,N_19415);
nor U20453 (N_20453,N_19535,N_19477);
xnor U20454 (N_20454,N_19937,N_19520);
xnor U20455 (N_20455,N_19625,N_19436);
nand U20456 (N_20456,N_19622,N_19009);
nand U20457 (N_20457,N_19921,N_19406);
nand U20458 (N_20458,N_19618,N_19586);
xnor U20459 (N_20459,N_19842,N_19999);
xnor U20460 (N_20460,N_19449,N_19418);
nor U20461 (N_20461,N_19010,N_19741);
nand U20462 (N_20462,N_19060,N_19092);
or U20463 (N_20463,N_19664,N_19723);
nand U20464 (N_20464,N_19079,N_19835);
or U20465 (N_20465,N_19200,N_19322);
nand U20466 (N_20466,N_19607,N_19183);
nand U20467 (N_20467,N_19829,N_19512);
or U20468 (N_20468,N_19498,N_19818);
or U20469 (N_20469,N_19870,N_19879);
xnor U20470 (N_20470,N_19574,N_19865);
nor U20471 (N_20471,N_19550,N_19549);
and U20472 (N_20472,N_19426,N_19413);
nand U20473 (N_20473,N_19952,N_19711);
or U20474 (N_20474,N_19403,N_19733);
nand U20475 (N_20475,N_19180,N_19071);
and U20476 (N_20476,N_19895,N_19668);
xnor U20477 (N_20477,N_19903,N_19340);
nand U20478 (N_20478,N_19251,N_19864);
and U20479 (N_20479,N_19642,N_19119);
and U20480 (N_20480,N_19114,N_19156);
or U20481 (N_20481,N_19592,N_19289);
or U20482 (N_20482,N_19881,N_19757);
and U20483 (N_20483,N_19024,N_19362);
or U20484 (N_20484,N_19391,N_19824);
xnor U20485 (N_20485,N_19147,N_19372);
or U20486 (N_20486,N_19035,N_19453);
xor U20487 (N_20487,N_19794,N_19185);
nor U20488 (N_20488,N_19779,N_19821);
nor U20489 (N_20489,N_19076,N_19598);
or U20490 (N_20490,N_19755,N_19713);
xnor U20491 (N_20491,N_19252,N_19786);
nor U20492 (N_20492,N_19899,N_19240);
nor U20493 (N_20493,N_19319,N_19109);
or U20494 (N_20494,N_19238,N_19059);
xnor U20495 (N_20495,N_19987,N_19229);
nand U20496 (N_20496,N_19020,N_19221);
and U20497 (N_20497,N_19090,N_19580);
or U20498 (N_20498,N_19465,N_19891);
and U20499 (N_20499,N_19503,N_19796);
and U20500 (N_20500,N_19493,N_19111);
nor U20501 (N_20501,N_19198,N_19175);
or U20502 (N_20502,N_19962,N_19744);
and U20503 (N_20503,N_19125,N_19449);
nand U20504 (N_20504,N_19689,N_19979);
or U20505 (N_20505,N_19789,N_19019);
nand U20506 (N_20506,N_19120,N_19888);
xor U20507 (N_20507,N_19921,N_19070);
nand U20508 (N_20508,N_19057,N_19277);
and U20509 (N_20509,N_19468,N_19311);
or U20510 (N_20510,N_19429,N_19565);
and U20511 (N_20511,N_19496,N_19125);
and U20512 (N_20512,N_19252,N_19654);
nand U20513 (N_20513,N_19121,N_19249);
xnor U20514 (N_20514,N_19595,N_19877);
xor U20515 (N_20515,N_19430,N_19551);
and U20516 (N_20516,N_19793,N_19000);
nor U20517 (N_20517,N_19732,N_19577);
nor U20518 (N_20518,N_19862,N_19564);
nand U20519 (N_20519,N_19987,N_19363);
nor U20520 (N_20520,N_19994,N_19689);
xnor U20521 (N_20521,N_19175,N_19336);
nor U20522 (N_20522,N_19420,N_19794);
xnor U20523 (N_20523,N_19060,N_19465);
or U20524 (N_20524,N_19397,N_19367);
and U20525 (N_20525,N_19751,N_19551);
nor U20526 (N_20526,N_19383,N_19955);
and U20527 (N_20527,N_19476,N_19420);
and U20528 (N_20528,N_19382,N_19205);
and U20529 (N_20529,N_19884,N_19769);
or U20530 (N_20530,N_19903,N_19095);
and U20531 (N_20531,N_19018,N_19506);
xor U20532 (N_20532,N_19866,N_19606);
nor U20533 (N_20533,N_19650,N_19924);
nor U20534 (N_20534,N_19831,N_19278);
nor U20535 (N_20535,N_19423,N_19998);
and U20536 (N_20536,N_19352,N_19973);
or U20537 (N_20537,N_19484,N_19516);
or U20538 (N_20538,N_19437,N_19446);
or U20539 (N_20539,N_19405,N_19442);
or U20540 (N_20540,N_19664,N_19536);
nor U20541 (N_20541,N_19174,N_19182);
xor U20542 (N_20542,N_19333,N_19977);
and U20543 (N_20543,N_19460,N_19889);
or U20544 (N_20544,N_19461,N_19733);
and U20545 (N_20545,N_19266,N_19928);
xnor U20546 (N_20546,N_19902,N_19246);
or U20547 (N_20547,N_19784,N_19308);
nor U20548 (N_20548,N_19189,N_19320);
nor U20549 (N_20549,N_19984,N_19936);
nor U20550 (N_20550,N_19609,N_19533);
and U20551 (N_20551,N_19285,N_19147);
and U20552 (N_20552,N_19069,N_19183);
nand U20553 (N_20553,N_19136,N_19572);
or U20554 (N_20554,N_19878,N_19979);
and U20555 (N_20555,N_19234,N_19514);
and U20556 (N_20556,N_19573,N_19225);
nor U20557 (N_20557,N_19637,N_19424);
xor U20558 (N_20558,N_19443,N_19347);
or U20559 (N_20559,N_19519,N_19724);
xor U20560 (N_20560,N_19511,N_19449);
or U20561 (N_20561,N_19047,N_19201);
or U20562 (N_20562,N_19193,N_19783);
or U20563 (N_20563,N_19183,N_19014);
and U20564 (N_20564,N_19523,N_19150);
nor U20565 (N_20565,N_19686,N_19715);
xnor U20566 (N_20566,N_19404,N_19720);
xor U20567 (N_20567,N_19648,N_19354);
nor U20568 (N_20568,N_19013,N_19162);
nor U20569 (N_20569,N_19539,N_19035);
and U20570 (N_20570,N_19464,N_19570);
xor U20571 (N_20571,N_19481,N_19240);
nand U20572 (N_20572,N_19560,N_19924);
nor U20573 (N_20573,N_19323,N_19280);
xnor U20574 (N_20574,N_19894,N_19896);
nand U20575 (N_20575,N_19450,N_19716);
xor U20576 (N_20576,N_19176,N_19751);
and U20577 (N_20577,N_19944,N_19452);
nand U20578 (N_20578,N_19644,N_19921);
and U20579 (N_20579,N_19928,N_19028);
nand U20580 (N_20580,N_19682,N_19019);
nor U20581 (N_20581,N_19827,N_19048);
nand U20582 (N_20582,N_19937,N_19039);
xnor U20583 (N_20583,N_19270,N_19042);
xor U20584 (N_20584,N_19698,N_19318);
xnor U20585 (N_20585,N_19616,N_19989);
nor U20586 (N_20586,N_19189,N_19462);
xnor U20587 (N_20587,N_19370,N_19945);
nor U20588 (N_20588,N_19057,N_19649);
xor U20589 (N_20589,N_19517,N_19831);
nor U20590 (N_20590,N_19927,N_19928);
xor U20591 (N_20591,N_19790,N_19002);
xnor U20592 (N_20592,N_19704,N_19637);
or U20593 (N_20593,N_19348,N_19906);
xor U20594 (N_20594,N_19512,N_19385);
and U20595 (N_20595,N_19890,N_19858);
xor U20596 (N_20596,N_19410,N_19506);
and U20597 (N_20597,N_19889,N_19289);
nand U20598 (N_20598,N_19934,N_19011);
nor U20599 (N_20599,N_19404,N_19671);
and U20600 (N_20600,N_19921,N_19525);
xnor U20601 (N_20601,N_19726,N_19423);
and U20602 (N_20602,N_19232,N_19831);
nor U20603 (N_20603,N_19682,N_19037);
nand U20604 (N_20604,N_19523,N_19963);
and U20605 (N_20605,N_19307,N_19923);
xnor U20606 (N_20606,N_19557,N_19380);
nor U20607 (N_20607,N_19057,N_19672);
xor U20608 (N_20608,N_19045,N_19647);
nand U20609 (N_20609,N_19282,N_19590);
or U20610 (N_20610,N_19647,N_19520);
or U20611 (N_20611,N_19287,N_19027);
xnor U20612 (N_20612,N_19814,N_19460);
nand U20613 (N_20613,N_19238,N_19751);
nor U20614 (N_20614,N_19003,N_19751);
nand U20615 (N_20615,N_19665,N_19711);
nor U20616 (N_20616,N_19626,N_19238);
nand U20617 (N_20617,N_19532,N_19489);
nor U20618 (N_20618,N_19432,N_19299);
xnor U20619 (N_20619,N_19913,N_19312);
or U20620 (N_20620,N_19731,N_19949);
or U20621 (N_20621,N_19989,N_19202);
and U20622 (N_20622,N_19885,N_19287);
nor U20623 (N_20623,N_19658,N_19994);
xor U20624 (N_20624,N_19956,N_19752);
nor U20625 (N_20625,N_19900,N_19601);
and U20626 (N_20626,N_19247,N_19740);
xor U20627 (N_20627,N_19193,N_19627);
or U20628 (N_20628,N_19123,N_19490);
xnor U20629 (N_20629,N_19116,N_19453);
nand U20630 (N_20630,N_19836,N_19283);
xor U20631 (N_20631,N_19226,N_19276);
nand U20632 (N_20632,N_19327,N_19080);
nand U20633 (N_20633,N_19209,N_19123);
nor U20634 (N_20634,N_19765,N_19641);
xnor U20635 (N_20635,N_19200,N_19924);
or U20636 (N_20636,N_19514,N_19080);
nor U20637 (N_20637,N_19712,N_19027);
xnor U20638 (N_20638,N_19908,N_19600);
and U20639 (N_20639,N_19401,N_19399);
and U20640 (N_20640,N_19358,N_19269);
or U20641 (N_20641,N_19630,N_19067);
nor U20642 (N_20642,N_19191,N_19464);
and U20643 (N_20643,N_19809,N_19618);
or U20644 (N_20644,N_19612,N_19114);
xor U20645 (N_20645,N_19909,N_19213);
or U20646 (N_20646,N_19614,N_19899);
nor U20647 (N_20647,N_19212,N_19909);
xnor U20648 (N_20648,N_19758,N_19386);
or U20649 (N_20649,N_19434,N_19092);
xor U20650 (N_20650,N_19099,N_19387);
and U20651 (N_20651,N_19701,N_19237);
or U20652 (N_20652,N_19261,N_19418);
nor U20653 (N_20653,N_19164,N_19491);
nor U20654 (N_20654,N_19419,N_19034);
or U20655 (N_20655,N_19871,N_19286);
xor U20656 (N_20656,N_19396,N_19207);
xnor U20657 (N_20657,N_19473,N_19687);
and U20658 (N_20658,N_19695,N_19634);
nand U20659 (N_20659,N_19137,N_19551);
xor U20660 (N_20660,N_19226,N_19866);
and U20661 (N_20661,N_19516,N_19683);
nor U20662 (N_20662,N_19210,N_19359);
and U20663 (N_20663,N_19061,N_19374);
nand U20664 (N_20664,N_19617,N_19035);
and U20665 (N_20665,N_19726,N_19081);
nor U20666 (N_20666,N_19075,N_19299);
or U20667 (N_20667,N_19138,N_19196);
xor U20668 (N_20668,N_19672,N_19080);
nor U20669 (N_20669,N_19765,N_19983);
xor U20670 (N_20670,N_19053,N_19460);
xor U20671 (N_20671,N_19704,N_19063);
or U20672 (N_20672,N_19696,N_19095);
xnor U20673 (N_20673,N_19533,N_19483);
nor U20674 (N_20674,N_19262,N_19118);
and U20675 (N_20675,N_19451,N_19885);
nand U20676 (N_20676,N_19629,N_19043);
or U20677 (N_20677,N_19218,N_19576);
or U20678 (N_20678,N_19919,N_19731);
nand U20679 (N_20679,N_19491,N_19874);
nand U20680 (N_20680,N_19050,N_19866);
nor U20681 (N_20681,N_19934,N_19110);
xor U20682 (N_20682,N_19181,N_19517);
nor U20683 (N_20683,N_19072,N_19661);
or U20684 (N_20684,N_19458,N_19764);
and U20685 (N_20685,N_19858,N_19609);
and U20686 (N_20686,N_19461,N_19337);
xor U20687 (N_20687,N_19098,N_19573);
and U20688 (N_20688,N_19125,N_19083);
xnor U20689 (N_20689,N_19124,N_19128);
nand U20690 (N_20690,N_19401,N_19410);
nor U20691 (N_20691,N_19340,N_19821);
nor U20692 (N_20692,N_19403,N_19686);
nor U20693 (N_20693,N_19466,N_19533);
nand U20694 (N_20694,N_19134,N_19452);
xor U20695 (N_20695,N_19178,N_19219);
and U20696 (N_20696,N_19355,N_19326);
xnor U20697 (N_20697,N_19856,N_19140);
xnor U20698 (N_20698,N_19385,N_19567);
and U20699 (N_20699,N_19603,N_19572);
and U20700 (N_20700,N_19915,N_19450);
xnor U20701 (N_20701,N_19600,N_19756);
xor U20702 (N_20702,N_19967,N_19698);
and U20703 (N_20703,N_19963,N_19258);
nand U20704 (N_20704,N_19483,N_19485);
or U20705 (N_20705,N_19934,N_19281);
nor U20706 (N_20706,N_19117,N_19302);
nor U20707 (N_20707,N_19642,N_19095);
xor U20708 (N_20708,N_19057,N_19713);
and U20709 (N_20709,N_19914,N_19523);
nand U20710 (N_20710,N_19090,N_19877);
and U20711 (N_20711,N_19407,N_19644);
nor U20712 (N_20712,N_19272,N_19523);
xor U20713 (N_20713,N_19816,N_19316);
xnor U20714 (N_20714,N_19098,N_19623);
xnor U20715 (N_20715,N_19225,N_19392);
nand U20716 (N_20716,N_19239,N_19364);
nor U20717 (N_20717,N_19516,N_19804);
and U20718 (N_20718,N_19482,N_19683);
or U20719 (N_20719,N_19926,N_19821);
nor U20720 (N_20720,N_19820,N_19951);
or U20721 (N_20721,N_19381,N_19210);
nor U20722 (N_20722,N_19210,N_19025);
and U20723 (N_20723,N_19554,N_19012);
xor U20724 (N_20724,N_19508,N_19230);
or U20725 (N_20725,N_19541,N_19502);
nor U20726 (N_20726,N_19989,N_19015);
or U20727 (N_20727,N_19399,N_19975);
or U20728 (N_20728,N_19723,N_19878);
and U20729 (N_20729,N_19762,N_19074);
and U20730 (N_20730,N_19330,N_19353);
xor U20731 (N_20731,N_19751,N_19175);
nand U20732 (N_20732,N_19887,N_19758);
and U20733 (N_20733,N_19471,N_19106);
or U20734 (N_20734,N_19817,N_19581);
nand U20735 (N_20735,N_19081,N_19426);
nor U20736 (N_20736,N_19793,N_19193);
xnor U20737 (N_20737,N_19596,N_19549);
xor U20738 (N_20738,N_19121,N_19083);
xnor U20739 (N_20739,N_19414,N_19609);
nor U20740 (N_20740,N_19389,N_19805);
xnor U20741 (N_20741,N_19449,N_19049);
xnor U20742 (N_20742,N_19624,N_19677);
xnor U20743 (N_20743,N_19202,N_19114);
and U20744 (N_20744,N_19725,N_19136);
xnor U20745 (N_20745,N_19070,N_19575);
nor U20746 (N_20746,N_19491,N_19708);
and U20747 (N_20747,N_19978,N_19040);
nor U20748 (N_20748,N_19586,N_19175);
nand U20749 (N_20749,N_19018,N_19692);
or U20750 (N_20750,N_19642,N_19351);
and U20751 (N_20751,N_19746,N_19869);
xor U20752 (N_20752,N_19840,N_19256);
nor U20753 (N_20753,N_19118,N_19510);
and U20754 (N_20754,N_19242,N_19739);
and U20755 (N_20755,N_19987,N_19755);
nor U20756 (N_20756,N_19078,N_19915);
xor U20757 (N_20757,N_19306,N_19766);
nand U20758 (N_20758,N_19654,N_19456);
xor U20759 (N_20759,N_19948,N_19416);
or U20760 (N_20760,N_19160,N_19065);
nand U20761 (N_20761,N_19422,N_19110);
nand U20762 (N_20762,N_19005,N_19940);
or U20763 (N_20763,N_19410,N_19748);
nand U20764 (N_20764,N_19844,N_19948);
nor U20765 (N_20765,N_19966,N_19883);
nor U20766 (N_20766,N_19579,N_19396);
nor U20767 (N_20767,N_19927,N_19439);
xnor U20768 (N_20768,N_19418,N_19891);
and U20769 (N_20769,N_19292,N_19430);
nand U20770 (N_20770,N_19274,N_19602);
and U20771 (N_20771,N_19766,N_19384);
and U20772 (N_20772,N_19370,N_19069);
or U20773 (N_20773,N_19048,N_19955);
or U20774 (N_20774,N_19653,N_19779);
xnor U20775 (N_20775,N_19605,N_19914);
or U20776 (N_20776,N_19107,N_19053);
and U20777 (N_20777,N_19024,N_19777);
nor U20778 (N_20778,N_19241,N_19116);
nand U20779 (N_20779,N_19407,N_19650);
xnor U20780 (N_20780,N_19481,N_19056);
nand U20781 (N_20781,N_19767,N_19427);
and U20782 (N_20782,N_19474,N_19147);
or U20783 (N_20783,N_19874,N_19213);
nand U20784 (N_20784,N_19063,N_19032);
nand U20785 (N_20785,N_19393,N_19198);
nor U20786 (N_20786,N_19559,N_19648);
nor U20787 (N_20787,N_19022,N_19850);
and U20788 (N_20788,N_19613,N_19292);
and U20789 (N_20789,N_19996,N_19374);
xor U20790 (N_20790,N_19275,N_19021);
nor U20791 (N_20791,N_19882,N_19690);
or U20792 (N_20792,N_19684,N_19054);
nand U20793 (N_20793,N_19367,N_19787);
and U20794 (N_20794,N_19384,N_19907);
nor U20795 (N_20795,N_19438,N_19556);
and U20796 (N_20796,N_19265,N_19440);
xnor U20797 (N_20797,N_19344,N_19796);
nor U20798 (N_20798,N_19100,N_19527);
or U20799 (N_20799,N_19726,N_19775);
or U20800 (N_20800,N_19017,N_19199);
and U20801 (N_20801,N_19508,N_19935);
nand U20802 (N_20802,N_19997,N_19112);
or U20803 (N_20803,N_19422,N_19338);
xor U20804 (N_20804,N_19253,N_19624);
xor U20805 (N_20805,N_19687,N_19284);
nand U20806 (N_20806,N_19940,N_19289);
xor U20807 (N_20807,N_19499,N_19599);
and U20808 (N_20808,N_19728,N_19773);
or U20809 (N_20809,N_19968,N_19621);
or U20810 (N_20810,N_19369,N_19735);
xor U20811 (N_20811,N_19309,N_19322);
and U20812 (N_20812,N_19882,N_19407);
nor U20813 (N_20813,N_19995,N_19330);
xor U20814 (N_20814,N_19777,N_19571);
or U20815 (N_20815,N_19093,N_19278);
nor U20816 (N_20816,N_19520,N_19446);
xor U20817 (N_20817,N_19086,N_19208);
xor U20818 (N_20818,N_19815,N_19569);
and U20819 (N_20819,N_19898,N_19048);
nand U20820 (N_20820,N_19504,N_19989);
and U20821 (N_20821,N_19953,N_19389);
and U20822 (N_20822,N_19981,N_19475);
or U20823 (N_20823,N_19205,N_19629);
and U20824 (N_20824,N_19124,N_19948);
nor U20825 (N_20825,N_19901,N_19807);
and U20826 (N_20826,N_19517,N_19040);
nand U20827 (N_20827,N_19668,N_19971);
nand U20828 (N_20828,N_19542,N_19234);
xor U20829 (N_20829,N_19118,N_19237);
or U20830 (N_20830,N_19044,N_19864);
xnor U20831 (N_20831,N_19424,N_19763);
nand U20832 (N_20832,N_19213,N_19068);
xor U20833 (N_20833,N_19833,N_19842);
xor U20834 (N_20834,N_19613,N_19960);
or U20835 (N_20835,N_19474,N_19749);
nand U20836 (N_20836,N_19236,N_19350);
xnor U20837 (N_20837,N_19799,N_19476);
nor U20838 (N_20838,N_19441,N_19211);
nand U20839 (N_20839,N_19298,N_19645);
or U20840 (N_20840,N_19888,N_19827);
xnor U20841 (N_20841,N_19486,N_19073);
or U20842 (N_20842,N_19101,N_19912);
nand U20843 (N_20843,N_19882,N_19646);
or U20844 (N_20844,N_19640,N_19143);
xnor U20845 (N_20845,N_19548,N_19524);
and U20846 (N_20846,N_19039,N_19237);
and U20847 (N_20847,N_19363,N_19493);
and U20848 (N_20848,N_19899,N_19101);
nor U20849 (N_20849,N_19999,N_19007);
or U20850 (N_20850,N_19240,N_19122);
nor U20851 (N_20851,N_19093,N_19318);
xor U20852 (N_20852,N_19625,N_19852);
and U20853 (N_20853,N_19152,N_19417);
nand U20854 (N_20854,N_19333,N_19193);
nor U20855 (N_20855,N_19254,N_19303);
xnor U20856 (N_20856,N_19131,N_19514);
xor U20857 (N_20857,N_19252,N_19829);
nor U20858 (N_20858,N_19442,N_19253);
nand U20859 (N_20859,N_19381,N_19447);
or U20860 (N_20860,N_19760,N_19197);
and U20861 (N_20861,N_19740,N_19951);
nor U20862 (N_20862,N_19910,N_19255);
xor U20863 (N_20863,N_19006,N_19844);
xor U20864 (N_20864,N_19262,N_19178);
nor U20865 (N_20865,N_19793,N_19773);
nand U20866 (N_20866,N_19600,N_19029);
or U20867 (N_20867,N_19058,N_19157);
or U20868 (N_20868,N_19921,N_19414);
nor U20869 (N_20869,N_19250,N_19285);
or U20870 (N_20870,N_19904,N_19715);
xnor U20871 (N_20871,N_19618,N_19482);
xnor U20872 (N_20872,N_19982,N_19586);
nand U20873 (N_20873,N_19333,N_19526);
and U20874 (N_20874,N_19734,N_19601);
xnor U20875 (N_20875,N_19826,N_19289);
xor U20876 (N_20876,N_19860,N_19069);
nand U20877 (N_20877,N_19623,N_19995);
xor U20878 (N_20878,N_19979,N_19371);
nand U20879 (N_20879,N_19838,N_19577);
xor U20880 (N_20880,N_19252,N_19335);
or U20881 (N_20881,N_19796,N_19008);
nand U20882 (N_20882,N_19827,N_19427);
and U20883 (N_20883,N_19775,N_19331);
nor U20884 (N_20884,N_19830,N_19871);
nand U20885 (N_20885,N_19374,N_19249);
xor U20886 (N_20886,N_19782,N_19526);
nand U20887 (N_20887,N_19145,N_19901);
nor U20888 (N_20888,N_19603,N_19077);
and U20889 (N_20889,N_19934,N_19103);
or U20890 (N_20890,N_19693,N_19344);
and U20891 (N_20891,N_19839,N_19032);
and U20892 (N_20892,N_19064,N_19029);
and U20893 (N_20893,N_19813,N_19844);
or U20894 (N_20894,N_19068,N_19288);
nor U20895 (N_20895,N_19406,N_19589);
nor U20896 (N_20896,N_19395,N_19116);
and U20897 (N_20897,N_19423,N_19646);
xnor U20898 (N_20898,N_19020,N_19820);
nor U20899 (N_20899,N_19980,N_19439);
nor U20900 (N_20900,N_19328,N_19455);
nand U20901 (N_20901,N_19361,N_19850);
nand U20902 (N_20902,N_19147,N_19963);
nor U20903 (N_20903,N_19036,N_19613);
and U20904 (N_20904,N_19164,N_19023);
nand U20905 (N_20905,N_19321,N_19548);
and U20906 (N_20906,N_19205,N_19291);
xor U20907 (N_20907,N_19294,N_19628);
xnor U20908 (N_20908,N_19215,N_19097);
nand U20909 (N_20909,N_19289,N_19681);
or U20910 (N_20910,N_19291,N_19383);
or U20911 (N_20911,N_19462,N_19994);
and U20912 (N_20912,N_19430,N_19997);
and U20913 (N_20913,N_19242,N_19346);
nor U20914 (N_20914,N_19797,N_19325);
and U20915 (N_20915,N_19682,N_19457);
nand U20916 (N_20916,N_19593,N_19987);
xor U20917 (N_20917,N_19732,N_19674);
or U20918 (N_20918,N_19348,N_19967);
or U20919 (N_20919,N_19048,N_19223);
nor U20920 (N_20920,N_19317,N_19621);
and U20921 (N_20921,N_19424,N_19457);
nor U20922 (N_20922,N_19541,N_19771);
and U20923 (N_20923,N_19048,N_19909);
and U20924 (N_20924,N_19276,N_19392);
or U20925 (N_20925,N_19091,N_19440);
xnor U20926 (N_20926,N_19051,N_19763);
xnor U20927 (N_20927,N_19588,N_19362);
or U20928 (N_20928,N_19195,N_19850);
and U20929 (N_20929,N_19104,N_19509);
xor U20930 (N_20930,N_19479,N_19714);
and U20931 (N_20931,N_19351,N_19161);
nand U20932 (N_20932,N_19465,N_19335);
nor U20933 (N_20933,N_19115,N_19172);
and U20934 (N_20934,N_19953,N_19322);
xnor U20935 (N_20935,N_19237,N_19245);
xnor U20936 (N_20936,N_19834,N_19539);
or U20937 (N_20937,N_19552,N_19330);
xor U20938 (N_20938,N_19359,N_19069);
and U20939 (N_20939,N_19097,N_19232);
xnor U20940 (N_20940,N_19976,N_19907);
nand U20941 (N_20941,N_19138,N_19677);
and U20942 (N_20942,N_19667,N_19461);
xnor U20943 (N_20943,N_19924,N_19591);
nand U20944 (N_20944,N_19187,N_19529);
xnor U20945 (N_20945,N_19170,N_19407);
or U20946 (N_20946,N_19589,N_19563);
nor U20947 (N_20947,N_19747,N_19144);
nor U20948 (N_20948,N_19464,N_19619);
and U20949 (N_20949,N_19629,N_19266);
and U20950 (N_20950,N_19213,N_19742);
nand U20951 (N_20951,N_19673,N_19787);
nand U20952 (N_20952,N_19509,N_19758);
nor U20953 (N_20953,N_19248,N_19980);
and U20954 (N_20954,N_19202,N_19200);
nand U20955 (N_20955,N_19996,N_19313);
nor U20956 (N_20956,N_19978,N_19506);
xor U20957 (N_20957,N_19384,N_19036);
nand U20958 (N_20958,N_19395,N_19413);
xnor U20959 (N_20959,N_19554,N_19577);
xnor U20960 (N_20960,N_19649,N_19223);
nand U20961 (N_20961,N_19590,N_19770);
xnor U20962 (N_20962,N_19003,N_19067);
xnor U20963 (N_20963,N_19022,N_19766);
nor U20964 (N_20964,N_19385,N_19117);
nand U20965 (N_20965,N_19127,N_19665);
or U20966 (N_20966,N_19854,N_19513);
nor U20967 (N_20967,N_19615,N_19251);
and U20968 (N_20968,N_19024,N_19421);
nor U20969 (N_20969,N_19028,N_19698);
xor U20970 (N_20970,N_19161,N_19384);
xnor U20971 (N_20971,N_19090,N_19202);
xor U20972 (N_20972,N_19669,N_19196);
nand U20973 (N_20973,N_19277,N_19341);
xnor U20974 (N_20974,N_19516,N_19944);
xor U20975 (N_20975,N_19331,N_19350);
and U20976 (N_20976,N_19221,N_19572);
nor U20977 (N_20977,N_19125,N_19286);
or U20978 (N_20978,N_19749,N_19152);
or U20979 (N_20979,N_19757,N_19850);
or U20980 (N_20980,N_19435,N_19569);
xor U20981 (N_20981,N_19172,N_19060);
nor U20982 (N_20982,N_19315,N_19995);
nor U20983 (N_20983,N_19669,N_19796);
nand U20984 (N_20984,N_19892,N_19743);
and U20985 (N_20985,N_19850,N_19742);
nand U20986 (N_20986,N_19497,N_19966);
nand U20987 (N_20987,N_19177,N_19873);
nor U20988 (N_20988,N_19277,N_19622);
and U20989 (N_20989,N_19391,N_19666);
nand U20990 (N_20990,N_19966,N_19991);
nor U20991 (N_20991,N_19696,N_19351);
or U20992 (N_20992,N_19755,N_19941);
nor U20993 (N_20993,N_19333,N_19257);
xor U20994 (N_20994,N_19888,N_19643);
xnor U20995 (N_20995,N_19167,N_19975);
nand U20996 (N_20996,N_19112,N_19146);
xor U20997 (N_20997,N_19711,N_19568);
and U20998 (N_20998,N_19158,N_19497);
xnor U20999 (N_20999,N_19458,N_19145);
or U21000 (N_21000,N_20402,N_20597);
or U21001 (N_21001,N_20080,N_20638);
nand U21002 (N_21002,N_20579,N_20957);
and U21003 (N_21003,N_20216,N_20200);
or U21004 (N_21004,N_20149,N_20030);
and U21005 (N_21005,N_20570,N_20115);
or U21006 (N_21006,N_20013,N_20501);
or U21007 (N_21007,N_20525,N_20762);
xnor U21008 (N_21008,N_20511,N_20314);
or U21009 (N_21009,N_20681,N_20686);
xnor U21010 (N_21010,N_20932,N_20333);
nand U21011 (N_21011,N_20476,N_20391);
nor U21012 (N_21012,N_20411,N_20769);
xor U21013 (N_21013,N_20680,N_20857);
and U21014 (N_21014,N_20089,N_20838);
nand U21015 (N_21015,N_20822,N_20003);
nor U21016 (N_21016,N_20405,N_20202);
nor U21017 (N_21017,N_20169,N_20166);
nand U21018 (N_21018,N_20771,N_20455);
xnor U21019 (N_21019,N_20557,N_20327);
or U21020 (N_21020,N_20925,N_20374);
or U21021 (N_21021,N_20528,N_20183);
xor U21022 (N_21022,N_20279,N_20052);
nor U21023 (N_21023,N_20161,N_20793);
and U21024 (N_21024,N_20531,N_20599);
nor U21025 (N_21025,N_20732,N_20099);
and U21026 (N_21026,N_20361,N_20340);
nand U21027 (N_21027,N_20434,N_20380);
or U21028 (N_21028,N_20929,N_20900);
xnor U21029 (N_21029,N_20672,N_20723);
nand U21030 (N_21030,N_20009,N_20109);
and U21031 (N_21031,N_20590,N_20260);
or U21032 (N_21032,N_20170,N_20817);
xor U21033 (N_21033,N_20312,N_20317);
nor U21034 (N_21034,N_20945,N_20265);
nor U21035 (N_21035,N_20076,N_20687);
xnor U21036 (N_21036,N_20592,N_20330);
or U21037 (N_21037,N_20020,N_20372);
nor U21038 (N_21038,N_20022,N_20187);
or U21039 (N_21039,N_20882,N_20060);
nand U21040 (N_21040,N_20948,N_20286);
xor U21041 (N_21041,N_20228,N_20494);
nor U21042 (N_21042,N_20600,N_20789);
nor U21043 (N_21043,N_20868,N_20474);
nor U21044 (N_21044,N_20475,N_20015);
or U21045 (N_21045,N_20065,N_20255);
nand U21046 (N_21046,N_20223,N_20603);
or U21047 (N_21047,N_20140,N_20843);
and U21048 (N_21048,N_20119,N_20173);
or U21049 (N_21049,N_20496,N_20852);
nor U21050 (N_21050,N_20881,N_20921);
or U21051 (N_21051,N_20385,N_20826);
nor U21052 (N_21052,N_20427,N_20536);
xor U21053 (N_21053,N_20270,N_20870);
nor U21054 (N_21054,N_20561,N_20650);
and U21055 (N_21055,N_20998,N_20114);
xnor U21056 (N_21056,N_20025,N_20103);
nor U21057 (N_21057,N_20970,N_20155);
nand U21058 (N_21058,N_20923,N_20702);
xnor U21059 (N_21059,N_20079,N_20378);
or U21060 (N_21060,N_20985,N_20643);
nor U21061 (N_21061,N_20437,N_20211);
nor U21062 (N_21062,N_20731,N_20457);
nand U21063 (N_21063,N_20224,N_20440);
nand U21064 (N_21064,N_20084,N_20087);
xnor U21065 (N_21065,N_20163,N_20978);
and U21066 (N_21066,N_20352,N_20398);
and U21067 (N_21067,N_20553,N_20575);
nand U21068 (N_21068,N_20741,N_20546);
and U21069 (N_21069,N_20645,N_20990);
or U21070 (N_21070,N_20979,N_20240);
or U21071 (N_21071,N_20653,N_20168);
xor U21072 (N_21072,N_20282,N_20021);
or U21073 (N_21073,N_20300,N_20469);
nand U21074 (N_21074,N_20757,N_20273);
xor U21075 (N_21075,N_20112,N_20639);
or U21076 (N_21076,N_20151,N_20285);
and U21077 (N_21077,N_20134,N_20542);
or U21078 (N_21078,N_20544,N_20002);
nor U21079 (N_21079,N_20413,N_20956);
or U21080 (N_21080,N_20520,N_20477);
and U21081 (N_21081,N_20001,N_20675);
and U21082 (N_21082,N_20818,N_20866);
xor U21083 (N_21083,N_20752,N_20038);
or U21084 (N_21084,N_20696,N_20659);
xor U21085 (N_21085,N_20246,N_20484);
xor U21086 (N_21086,N_20035,N_20693);
or U21087 (N_21087,N_20037,N_20063);
xnor U21088 (N_21088,N_20941,N_20069);
nand U21089 (N_21089,N_20298,N_20690);
or U21090 (N_21090,N_20143,N_20368);
or U21091 (N_21091,N_20988,N_20887);
xor U21092 (N_21092,N_20966,N_20664);
xor U21093 (N_21093,N_20295,N_20628);
or U21094 (N_21094,N_20431,N_20328);
or U21095 (N_21095,N_20589,N_20231);
or U21096 (N_21096,N_20267,N_20635);
xor U21097 (N_21097,N_20976,N_20299);
or U21098 (N_21098,N_20981,N_20392);
nor U21099 (N_21099,N_20316,N_20624);
nor U21100 (N_21100,N_20626,N_20896);
nand U21101 (N_21101,N_20806,N_20666);
xor U21102 (N_21102,N_20417,N_20902);
nand U21103 (N_21103,N_20796,N_20182);
or U21104 (N_21104,N_20185,N_20699);
xor U21105 (N_21105,N_20620,N_20930);
or U21106 (N_21106,N_20602,N_20082);
nand U21107 (N_21107,N_20172,N_20801);
and U21108 (N_21108,N_20668,N_20233);
or U21109 (N_21109,N_20506,N_20607);
and U21110 (N_21110,N_20266,N_20623);
nand U21111 (N_21111,N_20019,N_20967);
and U21112 (N_21112,N_20220,N_20420);
xor U21113 (N_21113,N_20613,N_20236);
nor U21114 (N_21114,N_20920,N_20781);
or U21115 (N_21115,N_20113,N_20492);
or U21116 (N_21116,N_20294,N_20346);
and U21117 (N_21117,N_20018,N_20767);
or U21118 (N_21118,N_20011,N_20891);
xnor U21119 (N_21119,N_20379,N_20345);
xor U21120 (N_21120,N_20257,N_20101);
or U21121 (N_21121,N_20839,N_20414);
nand U21122 (N_21122,N_20780,N_20308);
nor U21123 (N_21123,N_20387,N_20051);
xnor U21124 (N_21124,N_20856,N_20844);
nand U21125 (N_21125,N_20463,N_20439);
nand U21126 (N_21126,N_20679,N_20263);
nand U21127 (N_21127,N_20321,N_20125);
or U21128 (N_21128,N_20232,N_20832);
nor U21129 (N_21129,N_20522,N_20548);
nor U21130 (N_21130,N_20962,N_20895);
nor U21131 (N_21131,N_20786,N_20987);
nor U21132 (N_21132,N_20869,N_20809);
nand U21133 (N_21133,N_20291,N_20351);
nand U21134 (N_21134,N_20132,N_20629);
xnor U21135 (N_21135,N_20523,N_20999);
or U21136 (N_21136,N_20761,N_20212);
and U21137 (N_21137,N_20918,N_20106);
nand U21138 (N_21138,N_20622,N_20448);
or U21139 (N_21139,N_20341,N_20239);
and U21140 (N_21140,N_20715,N_20581);
xor U21141 (N_21141,N_20192,N_20139);
and U21142 (N_21142,N_20652,N_20532);
nand U21143 (N_21143,N_20176,N_20738);
and U21144 (N_21144,N_20326,N_20563);
nor U21145 (N_21145,N_20794,N_20100);
or U21146 (N_21146,N_20334,N_20540);
nand U21147 (N_21147,N_20608,N_20452);
or U21148 (N_21148,N_20824,N_20517);
and U21149 (N_21149,N_20876,N_20621);
nand U21150 (N_21150,N_20423,N_20828);
and U21151 (N_21151,N_20377,N_20678);
or U21152 (N_21152,N_20245,N_20836);
nor U21153 (N_21153,N_20807,N_20552);
nor U21154 (N_21154,N_20443,N_20671);
or U21155 (N_21155,N_20823,N_20012);
xnor U21156 (N_21156,N_20545,N_20847);
nand U21157 (N_21157,N_20403,N_20584);
nand U21158 (N_21158,N_20797,N_20924);
xor U21159 (N_21159,N_20425,N_20127);
nand U21160 (N_21160,N_20248,N_20028);
or U21161 (N_21161,N_20062,N_20432);
or U21162 (N_21162,N_20649,N_20049);
or U21163 (N_21163,N_20859,N_20772);
nand U21164 (N_21164,N_20210,N_20335);
nor U21165 (N_21165,N_20081,N_20473);
nand U21166 (N_21166,N_20310,N_20467);
nor U21167 (N_21167,N_20568,N_20512);
or U21168 (N_21168,N_20651,N_20997);
xor U21169 (N_21169,N_20877,N_20784);
or U21170 (N_21170,N_20449,N_20039);
nand U21171 (N_21171,N_20208,N_20193);
nand U21172 (N_21172,N_20805,N_20878);
nor U21173 (N_21173,N_20207,N_20369);
nand U21174 (N_21174,N_20505,N_20913);
xor U21175 (N_21175,N_20903,N_20479);
and U21176 (N_21176,N_20861,N_20096);
nand U21177 (N_21177,N_20331,N_20213);
nor U21178 (N_21178,N_20630,N_20661);
nand U21179 (N_21179,N_20831,N_20008);
and U21180 (N_21180,N_20992,N_20787);
or U21181 (N_21181,N_20122,N_20515);
or U21182 (N_21182,N_20795,N_20243);
or U21183 (N_21183,N_20670,N_20935);
nand U21184 (N_21184,N_20167,N_20555);
nor U21185 (N_21185,N_20097,N_20683);
xor U21186 (N_21186,N_20980,N_20899);
and U21187 (N_21187,N_20936,N_20908);
and U21188 (N_21188,N_20130,N_20851);
and U21189 (N_21189,N_20296,N_20461);
and U21190 (N_21190,N_20524,N_20788);
nand U21191 (N_21191,N_20890,N_20964);
or U21192 (N_21192,N_20489,N_20318);
nor U21193 (N_21193,N_20107,N_20578);
and U21194 (N_21194,N_20867,N_20588);
and U21195 (N_21195,N_20137,N_20458);
or U21196 (N_21196,N_20803,N_20293);
or U21197 (N_21197,N_20014,N_20395);
nor U21198 (N_21198,N_20560,N_20388);
nor U21199 (N_21199,N_20819,N_20749);
and U21200 (N_21200,N_20961,N_20480);
nand U21201 (N_21201,N_20865,N_20031);
nor U21202 (N_21202,N_20066,N_20829);
and U21203 (N_21203,N_20586,N_20808);
nand U21204 (N_21204,N_20901,N_20487);
and U21205 (N_21205,N_20004,N_20526);
and U21206 (N_21206,N_20005,N_20641);
nand U21207 (N_21207,N_20539,N_20888);
or U21208 (N_21208,N_20533,N_20971);
xnor U21209 (N_21209,N_20104,N_20691);
and U21210 (N_21210,N_20313,N_20493);
xnor U21211 (N_21211,N_20569,N_20284);
nand U21212 (N_21212,N_20883,N_20689);
nor U21213 (N_21213,N_20952,N_20827);
nand U21214 (N_21214,N_20916,N_20339);
or U21215 (N_21215,N_20792,N_20124);
and U21216 (N_21216,N_20986,N_20301);
xnor U21217 (N_21217,N_20148,N_20841);
or U21218 (N_21218,N_20892,N_20186);
or U21219 (N_21219,N_20509,N_20644);
or U21220 (N_21220,N_20872,N_20059);
xor U21221 (N_21221,N_20583,N_20943);
nor U21222 (N_21222,N_20070,N_20604);
xor U21223 (N_21223,N_20311,N_20057);
or U21224 (N_21224,N_20230,N_20911);
nor U21225 (N_21225,N_20105,N_20048);
xor U21226 (N_21226,N_20766,N_20303);
or U21227 (N_21227,N_20329,N_20776);
and U21228 (N_21228,N_20085,N_20768);
or U21229 (N_21229,N_20904,N_20835);
and U21230 (N_21230,N_20550,N_20221);
nor U21231 (N_21231,N_20381,N_20409);
nor U21232 (N_21232,N_20047,N_20848);
and U21233 (N_21233,N_20529,N_20500);
or U21234 (N_21234,N_20587,N_20110);
nor U21235 (N_21235,N_20102,N_20343);
nand U21236 (N_21236,N_20142,N_20753);
and U21237 (N_21237,N_20460,N_20919);
nand U21238 (N_21238,N_20810,N_20042);
nand U21239 (N_21239,N_20276,N_20968);
xnor U21240 (N_21240,N_20421,N_20034);
nand U21241 (N_21241,N_20556,N_20033);
or U21242 (N_21242,N_20386,N_20363);
nor U21243 (N_21243,N_20779,N_20078);
or U21244 (N_21244,N_20754,N_20595);
nor U21245 (N_21245,N_20910,N_20247);
and U21246 (N_21246,N_20725,N_20485);
or U21247 (N_21247,N_20946,N_20072);
and U21248 (N_21248,N_20609,N_20171);
nand U21249 (N_21249,N_20174,N_20642);
nor U21250 (N_21250,N_20252,N_20949);
nor U21251 (N_21251,N_20275,N_20707);
and U21252 (N_21252,N_20601,N_20775);
or U21253 (N_21253,N_20799,N_20618);
nand U21254 (N_21254,N_20222,N_20942);
nand U21255 (N_21255,N_20740,N_20075);
nand U21256 (N_21256,N_20704,N_20237);
nor U21257 (N_21257,N_20855,N_20503);
or U21258 (N_21258,N_20906,N_20886);
and U21259 (N_21259,N_20606,N_20399);
nand U21260 (N_21260,N_20325,N_20108);
nand U21261 (N_21261,N_20697,N_20927);
or U21262 (N_21262,N_20154,N_20567);
nor U21263 (N_21263,N_20880,N_20393);
or U21264 (N_21264,N_20656,N_20464);
and U21265 (N_21265,N_20046,N_20763);
nand U21266 (N_21266,N_20574,N_20206);
or U21267 (N_21267,N_20041,N_20858);
xnor U21268 (N_21268,N_20073,N_20996);
nor U21269 (N_21269,N_20518,N_20415);
nor U21270 (N_21270,N_20993,N_20714);
nor U21271 (N_21271,N_20010,N_20319);
xnor U21272 (N_21272,N_20488,N_20180);
nor U21273 (N_21273,N_20241,N_20783);
or U21274 (N_21274,N_20138,N_20281);
nand U21275 (N_21275,N_20663,N_20879);
nand U21276 (N_21276,N_20147,N_20674);
xor U21277 (N_21277,N_20288,N_20396);
nand U21278 (N_21278,N_20144,N_20422);
nor U21279 (N_21279,N_20055,N_20893);
or U21280 (N_21280,N_20898,N_20268);
xor U21281 (N_21281,N_20324,N_20156);
xnor U21282 (N_21282,N_20755,N_20750);
and U21283 (N_21283,N_20131,N_20937);
and U21284 (N_21284,N_20874,N_20287);
or U21285 (N_21285,N_20371,N_20864);
and U21286 (N_21286,N_20989,N_20482);
and U21287 (N_21287,N_20933,N_20745);
xor U21288 (N_21288,N_20214,N_20748);
xor U21289 (N_21289,N_20472,N_20453);
nand U21290 (N_21290,N_20362,N_20922);
nand U21291 (N_21291,N_20323,N_20834);
xnor U21292 (N_21292,N_20721,N_20056);
or U21293 (N_21293,N_20706,N_20000);
nand U21294 (N_21294,N_20953,N_20969);
nor U21295 (N_21295,N_20277,N_20365);
xnor U21296 (N_21296,N_20845,N_20129);
or U21297 (N_21297,N_20160,N_20820);
or U21298 (N_21298,N_20181,N_20007);
or U21299 (N_21299,N_20777,N_20456);
nand U21300 (N_21300,N_20145,N_20627);
xor U21301 (N_21301,N_20465,N_20636);
and U21302 (N_21302,N_20963,N_20433);
or U21303 (N_21303,N_20735,N_20006);
nor U21304 (N_21304,N_20594,N_20029);
and U21305 (N_21305,N_20338,N_20337);
or U21306 (N_21306,N_20198,N_20537);
xnor U21307 (N_21307,N_20778,N_20812);
or U21308 (N_21308,N_20430,N_20435);
nand U21309 (N_21309,N_20673,N_20184);
xor U21310 (N_21310,N_20682,N_20242);
xor U21311 (N_21311,N_20747,N_20153);
nand U21312 (N_21312,N_20490,N_20800);
xnor U21313 (N_21313,N_20593,N_20495);
and U21314 (N_21314,N_20716,N_20229);
nor U21315 (N_21315,N_20278,N_20840);
xor U21316 (N_21316,N_20302,N_20734);
or U21317 (N_21317,N_20743,N_20905);
nand U21318 (N_21318,N_20585,N_20032);
nand U21319 (N_21319,N_20177,N_20632);
and U21320 (N_21320,N_20357,N_20894);
nor U21321 (N_21321,N_20068,N_20133);
xor U21322 (N_21322,N_20370,N_20092);
or U21323 (N_21323,N_20067,N_20217);
or U21324 (N_21324,N_20191,N_20928);
xor U21325 (N_21325,N_20884,N_20804);
and U21326 (N_21326,N_20195,N_20717);
nor U21327 (N_21327,N_20849,N_20416);
or U21328 (N_21328,N_20640,N_20373);
xor U21329 (N_21329,N_20907,N_20677);
and U21330 (N_21330,N_20519,N_20053);
xnor U21331 (N_21331,N_20662,N_20758);
nor U21332 (N_21332,N_20446,N_20660);
and U21333 (N_21333,N_20815,N_20135);
nor U21334 (N_21334,N_20259,N_20685);
xor U21335 (N_21335,N_20401,N_20159);
nor U21336 (N_21336,N_20535,N_20215);
nor U21337 (N_21337,N_20157,N_20562);
and U21338 (N_21338,N_20554,N_20499);
and U21339 (N_21339,N_20050,N_20853);
or U21340 (N_21340,N_20158,N_20564);
nand U21341 (N_21341,N_20814,N_20665);
or U21342 (N_21342,N_20975,N_20647);
nand U21343 (N_21343,N_20045,N_20023);
or U21344 (N_21344,N_20530,N_20719);
xnor U21345 (N_21345,N_20366,N_20534);
nor U21346 (N_21346,N_20958,N_20447);
and U21347 (N_21347,N_20790,N_20646);
nand U21348 (N_21348,N_20591,N_20269);
and U21349 (N_21349,N_20514,N_20359);
or U21350 (N_21350,N_20513,N_20304);
nor U21351 (N_21351,N_20091,N_20605);
nor U21352 (N_21352,N_20253,N_20558);
and U21353 (N_21353,N_20309,N_20912);
and U21354 (N_21354,N_20703,N_20959);
and U21355 (N_21355,N_20305,N_20272);
or U21356 (N_21356,N_20724,N_20141);
nor U21357 (N_21357,N_20718,N_20262);
and U21358 (N_21358,N_20218,N_20336);
nand U21359 (N_21359,N_20454,N_20965);
and U21360 (N_21360,N_20175,N_20244);
and U21361 (N_21361,N_20737,N_20438);
nand U21362 (N_21362,N_20376,N_20058);
nor U21363 (N_21363,N_20367,N_20667);
or U21364 (N_21364,N_20297,N_20654);
or U21365 (N_21365,N_20322,N_20315);
nand U21366 (N_21366,N_20390,N_20254);
and U21367 (N_21367,N_20611,N_20375);
nand U21368 (N_21368,N_20917,N_20655);
nand U21369 (N_21369,N_20850,N_20126);
nor U21370 (N_21370,N_20445,N_20356);
xor U21371 (N_21371,N_20727,N_20016);
nor U21372 (N_21372,N_20984,N_20705);
or U21373 (N_21373,N_20394,N_20692);
nand U21374 (N_21374,N_20350,N_20098);
nand U21375 (N_21375,N_20994,N_20711);
or U21376 (N_21376,N_20760,N_20821);
or U21377 (N_21377,N_20939,N_20813);
nor U21378 (N_21378,N_20701,N_20698);
xnor U21379 (N_21379,N_20353,N_20428);
xor U21380 (N_21380,N_20885,N_20842);
nand U21381 (N_21381,N_20344,N_20944);
or U21382 (N_21382,N_20770,N_20165);
nor U21383 (N_21383,N_20364,N_20450);
xnor U21384 (N_21384,N_20973,N_20547);
xor U21385 (N_21385,N_20064,N_20196);
and U21386 (N_21386,N_20742,N_20982);
or U21387 (N_21387,N_20773,N_20116);
or U21388 (N_21388,N_20798,N_20614);
xor U21389 (N_21389,N_20190,N_20090);
nor U21390 (N_21390,N_20938,N_20444);
or U21391 (N_21391,N_20283,N_20201);
nor U21392 (N_21392,N_20619,N_20830);
nand U21393 (N_21393,N_20261,N_20914);
or U21394 (N_21394,N_20451,N_20470);
nor U21395 (N_21395,N_20383,N_20384);
xnor U21396 (N_21396,N_20825,N_20347);
and U21397 (N_21397,N_20095,N_20249);
and U21398 (N_21398,N_20120,N_20093);
nand U21399 (N_21399,N_20871,N_20708);
or U21400 (N_21400,N_20764,N_20408);
nand U21401 (N_21401,N_20676,N_20576);
and U21402 (N_21402,N_20354,N_20227);
and U21403 (N_21403,N_20342,N_20136);
or U21404 (N_21404,N_20459,N_20991);
xor U21405 (N_21405,N_20150,N_20657);
xor U21406 (N_21406,N_20977,N_20290);
or U21407 (N_21407,N_20024,N_20419);
nor U21408 (N_21408,N_20926,N_20862);
xnor U21409 (N_21409,N_20205,N_20483);
nand U21410 (N_21410,N_20118,N_20785);
nor U21411 (N_21411,N_20695,N_20950);
or U21412 (N_21412,N_20036,N_20765);
and U21413 (N_21413,N_20209,N_20983);
and U21414 (N_21414,N_20027,N_20404);
nor U21415 (N_21415,N_20947,N_20722);
nand U21416 (N_21416,N_20225,N_20580);
nor U21417 (N_21417,N_20258,N_20292);
nor U21418 (N_21418,N_20559,N_20617);
or U21419 (N_21419,N_20498,N_20688);
and U21420 (N_21420,N_20960,N_20094);
nand U21421 (N_21421,N_20955,N_20468);
nor U21422 (N_21422,N_20406,N_20486);
and U21423 (N_21423,N_20410,N_20128);
nand U21424 (N_21424,N_20234,N_20759);
and U21425 (N_21425,N_20694,N_20863);
nand U21426 (N_21426,N_20730,N_20194);
or U21427 (N_21427,N_20264,N_20426);
nor U21428 (N_21428,N_20951,N_20407);
nor U21429 (N_21429,N_20846,N_20728);
nor U21430 (N_21430,N_20710,N_20199);
xor U21431 (N_21431,N_20491,N_20634);
nand U21432 (N_21432,N_20582,N_20429);
xor U21433 (N_21433,N_20700,N_20811);
nor U21434 (N_21434,N_20572,N_20397);
and U21435 (N_21435,N_20507,N_20179);
nor U21436 (N_21436,N_20162,N_20400);
or U21437 (N_21437,N_20543,N_20510);
nor U21438 (N_21438,N_20478,N_20729);
or U21439 (N_21439,N_20088,N_20791);
or U21440 (N_21440,N_20637,N_20615);
nor U21441 (N_21441,N_20565,N_20044);
nand U21442 (N_21442,N_20756,N_20238);
nor U21443 (N_21443,N_20713,N_20086);
xor U21444 (N_21444,N_20389,N_20197);
xor U21445 (N_21445,N_20837,N_20164);
nand U21446 (N_21446,N_20860,N_20504);
xor U21447 (N_21447,N_20521,N_20471);
nand U21448 (N_21448,N_20424,N_20442);
xor U21449 (N_21449,N_20875,N_20625);
nor U21450 (N_21450,N_20616,N_20077);
or U21451 (N_21451,N_20436,N_20497);
nand U21452 (N_21452,N_20481,N_20320);
or U21453 (N_21453,N_20782,N_20873);
and U21454 (N_21454,N_20571,N_20071);
nand U21455 (N_21455,N_20382,N_20631);
or U21456 (N_21456,N_20934,N_20751);
nor U21457 (N_21457,N_20658,N_20188);
nor U21458 (N_21458,N_20203,N_20121);
xnor U21459 (N_21459,N_20909,N_20502);
xor U21460 (N_21460,N_20974,N_20358);
nor U21461 (N_21461,N_20736,N_20566);
or U21462 (N_21462,N_20466,N_20348);
and U21463 (N_21463,N_20307,N_20720);
nor U21464 (N_21464,N_20083,N_20204);
nand U21465 (N_21465,N_20219,N_20854);
xor U21466 (N_21466,N_20889,N_20816);
or U21467 (N_21467,N_20355,N_20931);
nor U21468 (N_21468,N_20418,N_20774);
nand U21469 (N_21469,N_20360,N_20538);
nor U21470 (N_21470,N_20256,N_20669);
nor U21471 (N_21471,N_20648,N_20043);
xor U21472 (N_21472,N_20235,N_20915);
nor U21473 (N_21473,N_20280,N_20633);
and U21474 (N_21474,N_20972,N_20516);
and U21475 (N_21475,N_20226,N_20802);
or U21476 (N_21476,N_20733,N_20061);
or U21477 (N_21477,N_20527,N_20349);
or U21478 (N_21478,N_20712,N_20598);
nand U21479 (N_21479,N_20746,N_20612);
or U21480 (N_21480,N_20954,N_20251);
xor U21481 (N_21481,N_20897,N_20117);
or U21482 (N_21482,N_20332,N_20040);
and U21483 (N_21483,N_20271,N_20549);
nor U21484 (N_21484,N_20744,N_20026);
nand U21485 (N_21485,N_20189,N_20709);
xor U21486 (N_21486,N_20178,N_20573);
nand U21487 (N_21487,N_20508,N_20017);
or U21488 (N_21488,N_20441,N_20940);
nor U21489 (N_21489,N_20306,N_20833);
or U21490 (N_21490,N_20412,N_20111);
nor U21491 (N_21491,N_20289,N_20726);
nor U21492 (N_21492,N_20577,N_20684);
xor U21493 (N_21493,N_20739,N_20146);
nand U21494 (N_21494,N_20995,N_20551);
nor U21495 (N_21495,N_20596,N_20274);
nand U21496 (N_21496,N_20152,N_20462);
and U21497 (N_21497,N_20054,N_20074);
or U21498 (N_21498,N_20610,N_20541);
nand U21499 (N_21499,N_20250,N_20123);
nor U21500 (N_21500,N_20188,N_20546);
nand U21501 (N_21501,N_20482,N_20029);
nand U21502 (N_21502,N_20171,N_20524);
nor U21503 (N_21503,N_20807,N_20477);
or U21504 (N_21504,N_20976,N_20317);
and U21505 (N_21505,N_20696,N_20604);
xnor U21506 (N_21506,N_20537,N_20442);
and U21507 (N_21507,N_20819,N_20575);
nor U21508 (N_21508,N_20298,N_20797);
nor U21509 (N_21509,N_20215,N_20496);
xor U21510 (N_21510,N_20886,N_20482);
nor U21511 (N_21511,N_20636,N_20996);
or U21512 (N_21512,N_20705,N_20536);
or U21513 (N_21513,N_20606,N_20800);
nand U21514 (N_21514,N_20103,N_20612);
nor U21515 (N_21515,N_20144,N_20523);
nor U21516 (N_21516,N_20173,N_20950);
and U21517 (N_21517,N_20517,N_20224);
or U21518 (N_21518,N_20137,N_20477);
nand U21519 (N_21519,N_20563,N_20504);
or U21520 (N_21520,N_20797,N_20180);
and U21521 (N_21521,N_20120,N_20000);
or U21522 (N_21522,N_20654,N_20871);
xor U21523 (N_21523,N_20296,N_20453);
nand U21524 (N_21524,N_20832,N_20680);
nand U21525 (N_21525,N_20306,N_20593);
nor U21526 (N_21526,N_20341,N_20708);
nor U21527 (N_21527,N_20756,N_20918);
xnor U21528 (N_21528,N_20287,N_20666);
xor U21529 (N_21529,N_20840,N_20660);
and U21530 (N_21530,N_20319,N_20451);
nand U21531 (N_21531,N_20251,N_20851);
nand U21532 (N_21532,N_20635,N_20302);
xor U21533 (N_21533,N_20827,N_20107);
or U21534 (N_21534,N_20663,N_20806);
nor U21535 (N_21535,N_20430,N_20717);
nor U21536 (N_21536,N_20601,N_20254);
xnor U21537 (N_21537,N_20263,N_20943);
xnor U21538 (N_21538,N_20010,N_20162);
and U21539 (N_21539,N_20132,N_20319);
xor U21540 (N_21540,N_20431,N_20934);
nor U21541 (N_21541,N_20376,N_20450);
and U21542 (N_21542,N_20508,N_20126);
and U21543 (N_21543,N_20827,N_20595);
and U21544 (N_21544,N_20792,N_20613);
xnor U21545 (N_21545,N_20906,N_20237);
xor U21546 (N_21546,N_20328,N_20964);
and U21547 (N_21547,N_20704,N_20642);
nand U21548 (N_21548,N_20216,N_20538);
nor U21549 (N_21549,N_20316,N_20163);
xor U21550 (N_21550,N_20633,N_20835);
nor U21551 (N_21551,N_20379,N_20597);
xnor U21552 (N_21552,N_20297,N_20429);
xor U21553 (N_21553,N_20312,N_20198);
nor U21554 (N_21554,N_20597,N_20436);
nand U21555 (N_21555,N_20874,N_20705);
xor U21556 (N_21556,N_20687,N_20429);
nand U21557 (N_21557,N_20660,N_20640);
or U21558 (N_21558,N_20896,N_20430);
or U21559 (N_21559,N_20715,N_20700);
or U21560 (N_21560,N_20130,N_20768);
or U21561 (N_21561,N_20535,N_20428);
or U21562 (N_21562,N_20657,N_20179);
and U21563 (N_21563,N_20929,N_20705);
xor U21564 (N_21564,N_20084,N_20123);
nor U21565 (N_21565,N_20609,N_20844);
and U21566 (N_21566,N_20184,N_20036);
and U21567 (N_21567,N_20753,N_20093);
nand U21568 (N_21568,N_20328,N_20362);
or U21569 (N_21569,N_20605,N_20012);
and U21570 (N_21570,N_20015,N_20445);
and U21571 (N_21571,N_20776,N_20440);
nand U21572 (N_21572,N_20865,N_20563);
nor U21573 (N_21573,N_20769,N_20862);
nand U21574 (N_21574,N_20352,N_20437);
nor U21575 (N_21575,N_20663,N_20579);
xnor U21576 (N_21576,N_20597,N_20270);
xnor U21577 (N_21577,N_20343,N_20442);
nand U21578 (N_21578,N_20809,N_20855);
nand U21579 (N_21579,N_20799,N_20414);
or U21580 (N_21580,N_20655,N_20275);
xor U21581 (N_21581,N_20349,N_20645);
and U21582 (N_21582,N_20832,N_20956);
xor U21583 (N_21583,N_20167,N_20006);
nand U21584 (N_21584,N_20246,N_20654);
and U21585 (N_21585,N_20578,N_20638);
nand U21586 (N_21586,N_20511,N_20708);
or U21587 (N_21587,N_20080,N_20164);
nand U21588 (N_21588,N_20946,N_20897);
nand U21589 (N_21589,N_20336,N_20764);
or U21590 (N_21590,N_20730,N_20891);
nor U21591 (N_21591,N_20251,N_20849);
and U21592 (N_21592,N_20556,N_20255);
nor U21593 (N_21593,N_20200,N_20564);
and U21594 (N_21594,N_20018,N_20043);
nor U21595 (N_21595,N_20783,N_20442);
nor U21596 (N_21596,N_20341,N_20901);
nor U21597 (N_21597,N_20542,N_20328);
or U21598 (N_21598,N_20927,N_20679);
nor U21599 (N_21599,N_20755,N_20354);
nand U21600 (N_21600,N_20860,N_20621);
xnor U21601 (N_21601,N_20247,N_20379);
nor U21602 (N_21602,N_20005,N_20520);
or U21603 (N_21603,N_20659,N_20677);
xor U21604 (N_21604,N_20095,N_20251);
xnor U21605 (N_21605,N_20929,N_20334);
xor U21606 (N_21606,N_20922,N_20829);
nand U21607 (N_21607,N_20265,N_20806);
nand U21608 (N_21608,N_20587,N_20241);
and U21609 (N_21609,N_20110,N_20537);
nor U21610 (N_21610,N_20312,N_20651);
nor U21611 (N_21611,N_20901,N_20362);
and U21612 (N_21612,N_20222,N_20121);
nand U21613 (N_21613,N_20474,N_20103);
and U21614 (N_21614,N_20644,N_20146);
or U21615 (N_21615,N_20997,N_20933);
and U21616 (N_21616,N_20666,N_20961);
xor U21617 (N_21617,N_20189,N_20221);
xnor U21618 (N_21618,N_20790,N_20283);
or U21619 (N_21619,N_20023,N_20470);
nand U21620 (N_21620,N_20439,N_20138);
xnor U21621 (N_21621,N_20275,N_20825);
nor U21622 (N_21622,N_20211,N_20103);
or U21623 (N_21623,N_20707,N_20510);
or U21624 (N_21624,N_20022,N_20690);
nand U21625 (N_21625,N_20359,N_20865);
nor U21626 (N_21626,N_20186,N_20398);
or U21627 (N_21627,N_20507,N_20857);
or U21628 (N_21628,N_20266,N_20512);
and U21629 (N_21629,N_20083,N_20741);
nor U21630 (N_21630,N_20072,N_20629);
or U21631 (N_21631,N_20245,N_20930);
xor U21632 (N_21632,N_20090,N_20752);
nor U21633 (N_21633,N_20464,N_20994);
nand U21634 (N_21634,N_20459,N_20614);
nor U21635 (N_21635,N_20433,N_20728);
nor U21636 (N_21636,N_20640,N_20483);
nor U21637 (N_21637,N_20139,N_20722);
nand U21638 (N_21638,N_20272,N_20341);
and U21639 (N_21639,N_20528,N_20429);
xnor U21640 (N_21640,N_20429,N_20878);
or U21641 (N_21641,N_20435,N_20357);
or U21642 (N_21642,N_20140,N_20658);
nand U21643 (N_21643,N_20866,N_20997);
nor U21644 (N_21644,N_20816,N_20181);
nand U21645 (N_21645,N_20762,N_20518);
or U21646 (N_21646,N_20798,N_20985);
or U21647 (N_21647,N_20715,N_20558);
or U21648 (N_21648,N_20504,N_20715);
xnor U21649 (N_21649,N_20088,N_20401);
and U21650 (N_21650,N_20535,N_20976);
nor U21651 (N_21651,N_20592,N_20301);
and U21652 (N_21652,N_20668,N_20166);
and U21653 (N_21653,N_20268,N_20558);
and U21654 (N_21654,N_20045,N_20311);
or U21655 (N_21655,N_20337,N_20418);
nand U21656 (N_21656,N_20714,N_20681);
and U21657 (N_21657,N_20998,N_20480);
and U21658 (N_21658,N_20367,N_20765);
xnor U21659 (N_21659,N_20781,N_20089);
or U21660 (N_21660,N_20055,N_20619);
or U21661 (N_21661,N_20840,N_20464);
nand U21662 (N_21662,N_20791,N_20136);
xnor U21663 (N_21663,N_20718,N_20658);
or U21664 (N_21664,N_20190,N_20778);
nand U21665 (N_21665,N_20259,N_20369);
nor U21666 (N_21666,N_20141,N_20727);
and U21667 (N_21667,N_20452,N_20821);
nand U21668 (N_21668,N_20889,N_20248);
or U21669 (N_21669,N_20458,N_20069);
xnor U21670 (N_21670,N_20193,N_20851);
nand U21671 (N_21671,N_20156,N_20012);
nor U21672 (N_21672,N_20475,N_20692);
and U21673 (N_21673,N_20078,N_20373);
or U21674 (N_21674,N_20419,N_20770);
xnor U21675 (N_21675,N_20036,N_20346);
xnor U21676 (N_21676,N_20811,N_20361);
xor U21677 (N_21677,N_20827,N_20346);
and U21678 (N_21678,N_20562,N_20227);
nand U21679 (N_21679,N_20190,N_20989);
and U21680 (N_21680,N_20869,N_20747);
or U21681 (N_21681,N_20689,N_20017);
or U21682 (N_21682,N_20738,N_20229);
and U21683 (N_21683,N_20875,N_20819);
nor U21684 (N_21684,N_20252,N_20245);
nand U21685 (N_21685,N_20483,N_20463);
nand U21686 (N_21686,N_20801,N_20716);
and U21687 (N_21687,N_20986,N_20837);
or U21688 (N_21688,N_20283,N_20461);
xor U21689 (N_21689,N_20261,N_20333);
and U21690 (N_21690,N_20397,N_20985);
nor U21691 (N_21691,N_20215,N_20760);
nand U21692 (N_21692,N_20620,N_20108);
xnor U21693 (N_21693,N_20442,N_20666);
nand U21694 (N_21694,N_20821,N_20626);
or U21695 (N_21695,N_20780,N_20051);
nor U21696 (N_21696,N_20568,N_20653);
nand U21697 (N_21697,N_20200,N_20105);
nand U21698 (N_21698,N_20269,N_20131);
xor U21699 (N_21699,N_20514,N_20115);
nor U21700 (N_21700,N_20757,N_20857);
or U21701 (N_21701,N_20316,N_20382);
or U21702 (N_21702,N_20140,N_20364);
nand U21703 (N_21703,N_20409,N_20982);
nor U21704 (N_21704,N_20002,N_20473);
nor U21705 (N_21705,N_20119,N_20192);
and U21706 (N_21706,N_20008,N_20609);
xor U21707 (N_21707,N_20096,N_20284);
and U21708 (N_21708,N_20072,N_20525);
or U21709 (N_21709,N_20487,N_20494);
xor U21710 (N_21710,N_20625,N_20029);
nor U21711 (N_21711,N_20488,N_20371);
nand U21712 (N_21712,N_20129,N_20827);
or U21713 (N_21713,N_20557,N_20480);
nand U21714 (N_21714,N_20091,N_20745);
nor U21715 (N_21715,N_20891,N_20977);
or U21716 (N_21716,N_20372,N_20458);
or U21717 (N_21717,N_20418,N_20742);
and U21718 (N_21718,N_20598,N_20457);
nand U21719 (N_21719,N_20061,N_20991);
nand U21720 (N_21720,N_20530,N_20624);
xnor U21721 (N_21721,N_20092,N_20928);
nor U21722 (N_21722,N_20242,N_20254);
and U21723 (N_21723,N_20308,N_20162);
and U21724 (N_21724,N_20508,N_20801);
and U21725 (N_21725,N_20726,N_20327);
and U21726 (N_21726,N_20075,N_20272);
and U21727 (N_21727,N_20626,N_20047);
or U21728 (N_21728,N_20091,N_20694);
nor U21729 (N_21729,N_20193,N_20005);
nor U21730 (N_21730,N_20576,N_20337);
xnor U21731 (N_21731,N_20585,N_20593);
nor U21732 (N_21732,N_20844,N_20278);
nor U21733 (N_21733,N_20282,N_20307);
xor U21734 (N_21734,N_20638,N_20503);
nand U21735 (N_21735,N_20781,N_20434);
or U21736 (N_21736,N_20603,N_20659);
and U21737 (N_21737,N_20746,N_20387);
xor U21738 (N_21738,N_20048,N_20298);
xnor U21739 (N_21739,N_20117,N_20303);
and U21740 (N_21740,N_20019,N_20893);
and U21741 (N_21741,N_20244,N_20281);
xor U21742 (N_21742,N_20482,N_20672);
nand U21743 (N_21743,N_20205,N_20695);
xnor U21744 (N_21744,N_20520,N_20725);
xnor U21745 (N_21745,N_20473,N_20815);
xnor U21746 (N_21746,N_20064,N_20211);
and U21747 (N_21747,N_20303,N_20667);
or U21748 (N_21748,N_20247,N_20824);
nand U21749 (N_21749,N_20507,N_20341);
nand U21750 (N_21750,N_20699,N_20752);
or U21751 (N_21751,N_20608,N_20669);
nor U21752 (N_21752,N_20650,N_20830);
and U21753 (N_21753,N_20324,N_20146);
nor U21754 (N_21754,N_20660,N_20148);
nand U21755 (N_21755,N_20981,N_20849);
nand U21756 (N_21756,N_20834,N_20110);
and U21757 (N_21757,N_20939,N_20849);
and U21758 (N_21758,N_20005,N_20565);
and U21759 (N_21759,N_20302,N_20241);
and U21760 (N_21760,N_20003,N_20958);
and U21761 (N_21761,N_20258,N_20078);
or U21762 (N_21762,N_20337,N_20096);
or U21763 (N_21763,N_20513,N_20005);
xor U21764 (N_21764,N_20507,N_20283);
nand U21765 (N_21765,N_20322,N_20943);
nand U21766 (N_21766,N_20676,N_20812);
or U21767 (N_21767,N_20031,N_20930);
nor U21768 (N_21768,N_20516,N_20926);
xor U21769 (N_21769,N_20047,N_20368);
xnor U21770 (N_21770,N_20384,N_20375);
or U21771 (N_21771,N_20828,N_20270);
or U21772 (N_21772,N_20562,N_20256);
xnor U21773 (N_21773,N_20367,N_20143);
nand U21774 (N_21774,N_20681,N_20906);
nor U21775 (N_21775,N_20919,N_20255);
or U21776 (N_21776,N_20602,N_20375);
and U21777 (N_21777,N_20448,N_20222);
and U21778 (N_21778,N_20073,N_20329);
nand U21779 (N_21779,N_20573,N_20175);
nor U21780 (N_21780,N_20089,N_20430);
xor U21781 (N_21781,N_20408,N_20151);
and U21782 (N_21782,N_20551,N_20904);
xor U21783 (N_21783,N_20342,N_20885);
nor U21784 (N_21784,N_20172,N_20312);
nand U21785 (N_21785,N_20110,N_20694);
xor U21786 (N_21786,N_20979,N_20447);
nand U21787 (N_21787,N_20832,N_20260);
xnor U21788 (N_21788,N_20607,N_20092);
xnor U21789 (N_21789,N_20358,N_20539);
nor U21790 (N_21790,N_20453,N_20320);
xor U21791 (N_21791,N_20756,N_20285);
xnor U21792 (N_21792,N_20685,N_20197);
and U21793 (N_21793,N_20699,N_20112);
and U21794 (N_21794,N_20646,N_20916);
nor U21795 (N_21795,N_20993,N_20579);
xor U21796 (N_21796,N_20688,N_20481);
and U21797 (N_21797,N_20453,N_20483);
and U21798 (N_21798,N_20349,N_20830);
or U21799 (N_21799,N_20531,N_20485);
nor U21800 (N_21800,N_20751,N_20722);
nor U21801 (N_21801,N_20523,N_20637);
nand U21802 (N_21802,N_20128,N_20028);
nand U21803 (N_21803,N_20368,N_20703);
xnor U21804 (N_21804,N_20864,N_20967);
nand U21805 (N_21805,N_20083,N_20724);
or U21806 (N_21806,N_20379,N_20918);
and U21807 (N_21807,N_20298,N_20658);
or U21808 (N_21808,N_20175,N_20999);
nand U21809 (N_21809,N_20745,N_20326);
and U21810 (N_21810,N_20246,N_20044);
xor U21811 (N_21811,N_20543,N_20741);
nor U21812 (N_21812,N_20604,N_20859);
xor U21813 (N_21813,N_20786,N_20037);
or U21814 (N_21814,N_20643,N_20652);
nand U21815 (N_21815,N_20585,N_20276);
or U21816 (N_21816,N_20620,N_20857);
nor U21817 (N_21817,N_20325,N_20948);
and U21818 (N_21818,N_20937,N_20824);
nand U21819 (N_21819,N_20196,N_20396);
and U21820 (N_21820,N_20240,N_20506);
and U21821 (N_21821,N_20088,N_20083);
nand U21822 (N_21822,N_20671,N_20263);
nor U21823 (N_21823,N_20063,N_20113);
and U21824 (N_21824,N_20007,N_20361);
nand U21825 (N_21825,N_20894,N_20186);
nand U21826 (N_21826,N_20462,N_20650);
nand U21827 (N_21827,N_20448,N_20331);
and U21828 (N_21828,N_20478,N_20655);
nand U21829 (N_21829,N_20773,N_20186);
nand U21830 (N_21830,N_20642,N_20995);
xnor U21831 (N_21831,N_20782,N_20551);
and U21832 (N_21832,N_20490,N_20005);
nor U21833 (N_21833,N_20057,N_20184);
or U21834 (N_21834,N_20812,N_20660);
and U21835 (N_21835,N_20934,N_20540);
xnor U21836 (N_21836,N_20017,N_20577);
nand U21837 (N_21837,N_20977,N_20878);
nor U21838 (N_21838,N_20010,N_20473);
and U21839 (N_21839,N_20133,N_20924);
nand U21840 (N_21840,N_20067,N_20415);
nand U21841 (N_21841,N_20293,N_20241);
xnor U21842 (N_21842,N_20341,N_20088);
nor U21843 (N_21843,N_20452,N_20029);
nor U21844 (N_21844,N_20790,N_20393);
or U21845 (N_21845,N_20527,N_20577);
nand U21846 (N_21846,N_20927,N_20442);
and U21847 (N_21847,N_20724,N_20275);
nor U21848 (N_21848,N_20864,N_20568);
xor U21849 (N_21849,N_20145,N_20577);
nand U21850 (N_21850,N_20557,N_20838);
nor U21851 (N_21851,N_20605,N_20049);
nor U21852 (N_21852,N_20289,N_20382);
nor U21853 (N_21853,N_20890,N_20799);
nor U21854 (N_21854,N_20114,N_20904);
and U21855 (N_21855,N_20933,N_20587);
nand U21856 (N_21856,N_20493,N_20882);
or U21857 (N_21857,N_20966,N_20804);
nand U21858 (N_21858,N_20913,N_20887);
nand U21859 (N_21859,N_20872,N_20322);
nand U21860 (N_21860,N_20531,N_20035);
nand U21861 (N_21861,N_20593,N_20974);
or U21862 (N_21862,N_20546,N_20184);
nor U21863 (N_21863,N_20286,N_20944);
or U21864 (N_21864,N_20303,N_20803);
or U21865 (N_21865,N_20584,N_20086);
and U21866 (N_21866,N_20248,N_20533);
xor U21867 (N_21867,N_20380,N_20521);
xnor U21868 (N_21868,N_20322,N_20460);
nand U21869 (N_21869,N_20870,N_20330);
xor U21870 (N_21870,N_20717,N_20894);
xor U21871 (N_21871,N_20904,N_20459);
or U21872 (N_21872,N_20820,N_20302);
and U21873 (N_21873,N_20747,N_20284);
nor U21874 (N_21874,N_20327,N_20420);
nand U21875 (N_21875,N_20924,N_20572);
or U21876 (N_21876,N_20203,N_20304);
xor U21877 (N_21877,N_20767,N_20658);
nor U21878 (N_21878,N_20778,N_20404);
and U21879 (N_21879,N_20771,N_20177);
or U21880 (N_21880,N_20980,N_20090);
and U21881 (N_21881,N_20633,N_20760);
xor U21882 (N_21882,N_20083,N_20647);
xnor U21883 (N_21883,N_20338,N_20433);
nand U21884 (N_21884,N_20193,N_20945);
nand U21885 (N_21885,N_20873,N_20249);
and U21886 (N_21886,N_20983,N_20560);
xor U21887 (N_21887,N_20735,N_20869);
xnor U21888 (N_21888,N_20252,N_20383);
nor U21889 (N_21889,N_20657,N_20624);
and U21890 (N_21890,N_20932,N_20893);
or U21891 (N_21891,N_20222,N_20614);
nand U21892 (N_21892,N_20805,N_20239);
nand U21893 (N_21893,N_20938,N_20394);
nand U21894 (N_21894,N_20900,N_20061);
or U21895 (N_21895,N_20494,N_20148);
and U21896 (N_21896,N_20482,N_20307);
nor U21897 (N_21897,N_20101,N_20522);
nor U21898 (N_21898,N_20705,N_20470);
nor U21899 (N_21899,N_20268,N_20242);
nand U21900 (N_21900,N_20315,N_20526);
and U21901 (N_21901,N_20689,N_20842);
xnor U21902 (N_21902,N_20505,N_20726);
nand U21903 (N_21903,N_20378,N_20590);
or U21904 (N_21904,N_20003,N_20353);
nand U21905 (N_21905,N_20881,N_20750);
xor U21906 (N_21906,N_20963,N_20720);
xnor U21907 (N_21907,N_20419,N_20960);
or U21908 (N_21908,N_20959,N_20084);
or U21909 (N_21909,N_20697,N_20071);
nor U21910 (N_21910,N_20848,N_20246);
or U21911 (N_21911,N_20703,N_20972);
nand U21912 (N_21912,N_20583,N_20053);
and U21913 (N_21913,N_20088,N_20058);
xor U21914 (N_21914,N_20114,N_20716);
nor U21915 (N_21915,N_20857,N_20298);
or U21916 (N_21916,N_20685,N_20826);
and U21917 (N_21917,N_20025,N_20894);
xor U21918 (N_21918,N_20956,N_20858);
or U21919 (N_21919,N_20323,N_20583);
xnor U21920 (N_21920,N_20409,N_20324);
xnor U21921 (N_21921,N_20266,N_20579);
xor U21922 (N_21922,N_20361,N_20162);
or U21923 (N_21923,N_20401,N_20355);
or U21924 (N_21924,N_20372,N_20690);
or U21925 (N_21925,N_20419,N_20741);
xnor U21926 (N_21926,N_20638,N_20442);
xnor U21927 (N_21927,N_20983,N_20598);
or U21928 (N_21928,N_20157,N_20722);
or U21929 (N_21929,N_20844,N_20311);
or U21930 (N_21930,N_20027,N_20830);
nand U21931 (N_21931,N_20352,N_20073);
nor U21932 (N_21932,N_20460,N_20723);
and U21933 (N_21933,N_20169,N_20862);
nor U21934 (N_21934,N_20246,N_20884);
nor U21935 (N_21935,N_20010,N_20537);
or U21936 (N_21936,N_20634,N_20106);
nor U21937 (N_21937,N_20058,N_20502);
nor U21938 (N_21938,N_20356,N_20950);
and U21939 (N_21939,N_20566,N_20909);
and U21940 (N_21940,N_20568,N_20767);
nor U21941 (N_21941,N_20069,N_20963);
or U21942 (N_21942,N_20336,N_20726);
or U21943 (N_21943,N_20496,N_20506);
xor U21944 (N_21944,N_20221,N_20478);
xnor U21945 (N_21945,N_20182,N_20430);
and U21946 (N_21946,N_20787,N_20284);
nor U21947 (N_21947,N_20464,N_20417);
and U21948 (N_21948,N_20517,N_20923);
xnor U21949 (N_21949,N_20282,N_20934);
and U21950 (N_21950,N_20937,N_20507);
nand U21951 (N_21951,N_20925,N_20169);
nor U21952 (N_21952,N_20890,N_20869);
nor U21953 (N_21953,N_20045,N_20790);
or U21954 (N_21954,N_20879,N_20520);
nand U21955 (N_21955,N_20388,N_20845);
xnor U21956 (N_21956,N_20837,N_20780);
or U21957 (N_21957,N_20266,N_20775);
nand U21958 (N_21958,N_20669,N_20695);
nand U21959 (N_21959,N_20031,N_20877);
or U21960 (N_21960,N_20417,N_20612);
or U21961 (N_21961,N_20122,N_20031);
and U21962 (N_21962,N_20727,N_20817);
or U21963 (N_21963,N_20372,N_20452);
or U21964 (N_21964,N_20041,N_20373);
xor U21965 (N_21965,N_20186,N_20646);
xnor U21966 (N_21966,N_20446,N_20088);
xor U21967 (N_21967,N_20739,N_20766);
nor U21968 (N_21968,N_20654,N_20728);
nor U21969 (N_21969,N_20257,N_20053);
or U21970 (N_21970,N_20892,N_20503);
or U21971 (N_21971,N_20257,N_20408);
xor U21972 (N_21972,N_20906,N_20725);
or U21973 (N_21973,N_20771,N_20024);
and U21974 (N_21974,N_20345,N_20033);
nand U21975 (N_21975,N_20696,N_20473);
and U21976 (N_21976,N_20352,N_20017);
xor U21977 (N_21977,N_20357,N_20702);
or U21978 (N_21978,N_20521,N_20455);
nor U21979 (N_21979,N_20440,N_20482);
nand U21980 (N_21980,N_20940,N_20192);
nand U21981 (N_21981,N_20376,N_20344);
nor U21982 (N_21982,N_20529,N_20858);
nand U21983 (N_21983,N_20819,N_20189);
or U21984 (N_21984,N_20497,N_20152);
nor U21985 (N_21985,N_20259,N_20562);
or U21986 (N_21986,N_20047,N_20898);
nand U21987 (N_21987,N_20035,N_20343);
or U21988 (N_21988,N_20966,N_20473);
nand U21989 (N_21989,N_20949,N_20495);
xor U21990 (N_21990,N_20091,N_20623);
or U21991 (N_21991,N_20416,N_20238);
nand U21992 (N_21992,N_20639,N_20988);
nor U21993 (N_21993,N_20098,N_20742);
xnor U21994 (N_21994,N_20282,N_20077);
or U21995 (N_21995,N_20331,N_20208);
nand U21996 (N_21996,N_20300,N_20879);
nand U21997 (N_21997,N_20415,N_20349);
or U21998 (N_21998,N_20487,N_20042);
and U21999 (N_21999,N_20072,N_20788);
nand U22000 (N_22000,N_21981,N_21826);
nand U22001 (N_22001,N_21166,N_21637);
or U22002 (N_22002,N_21967,N_21906);
nor U22003 (N_22003,N_21953,N_21174);
or U22004 (N_22004,N_21626,N_21223);
and U22005 (N_22005,N_21351,N_21197);
nor U22006 (N_22006,N_21383,N_21522);
or U22007 (N_22007,N_21893,N_21369);
or U22008 (N_22008,N_21877,N_21433);
nor U22009 (N_22009,N_21661,N_21738);
nor U22010 (N_22010,N_21611,N_21085);
nand U22011 (N_22011,N_21175,N_21810);
nor U22012 (N_22012,N_21071,N_21663);
xor U22013 (N_22013,N_21016,N_21007);
nand U22014 (N_22014,N_21603,N_21377);
and U22015 (N_22015,N_21599,N_21779);
and U22016 (N_22016,N_21443,N_21279);
nor U22017 (N_22017,N_21534,N_21116);
nor U22018 (N_22018,N_21922,N_21628);
or U22019 (N_22019,N_21356,N_21364);
and U22020 (N_22020,N_21004,N_21244);
and U22021 (N_22021,N_21644,N_21501);
nand U22022 (N_22022,N_21586,N_21406);
or U22023 (N_22023,N_21718,N_21510);
nand U22024 (N_22024,N_21793,N_21683);
nor U22025 (N_22025,N_21427,N_21263);
nand U22026 (N_22026,N_21054,N_21104);
nor U22027 (N_22027,N_21574,N_21361);
xor U22028 (N_22028,N_21362,N_21024);
xnor U22029 (N_22029,N_21341,N_21310);
or U22030 (N_22030,N_21062,N_21014);
and U22031 (N_22031,N_21230,N_21401);
or U22032 (N_22032,N_21802,N_21192);
and U22033 (N_22033,N_21431,N_21493);
or U22034 (N_22034,N_21910,N_21524);
or U22035 (N_22035,N_21163,N_21667);
nand U22036 (N_22036,N_21971,N_21529);
xnor U22037 (N_22037,N_21641,N_21449);
or U22038 (N_22038,N_21213,N_21190);
nor U22039 (N_22039,N_21528,N_21010);
and U22040 (N_22040,N_21198,N_21972);
nor U22041 (N_22041,N_21030,N_21115);
nor U22042 (N_22042,N_21161,N_21656);
nor U22043 (N_22043,N_21622,N_21289);
nor U22044 (N_22044,N_21086,N_21479);
and U22045 (N_22045,N_21069,N_21535);
xor U22046 (N_22046,N_21357,N_21927);
and U22047 (N_22047,N_21410,N_21789);
nor U22048 (N_22048,N_21128,N_21896);
nor U22049 (N_22049,N_21933,N_21143);
nor U22050 (N_22050,N_21748,N_21499);
nand U22051 (N_22051,N_21009,N_21011);
or U22052 (N_22052,N_21977,N_21869);
nand U22053 (N_22053,N_21079,N_21898);
and U22054 (N_22054,N_21508,N_21891);
or U22055 (N_22055,N_21248,N_21767);
or U22056 (N_22056,N_21480,N_21582);
and U22057 (N_22057,N_21468,N_21117);
nor U22058 (N_22058,N_21160,N_21777);
xnor U22059 (N_22059,N_21956,N_21668);
xor U22060 (N_22060,N_21900,N_21658);
nor U22061 (N_22061,N_21268,N_21019);
or U22062 (N_22062,N_21285,N_21465);
xnor U22063 (N_22063,N_21220,N_21428);
and U22064 (N_22064,N_21476,N_21037);
and U22065 (N_22065,N_21039,N_21945);
xnor U22066 (N_22066,N_21478,N_21875);
xnor U22067 (N_22067,N_21243,N_21858);
nor U22068 (N_22068,N_21863,N_21634);
and U22069 (N_22069,N_21507,N_21295);
and U22070 (N_22070,N_21890,N_21380);
xor U22071 (N_22071,N_21600,N_21850);
xnor U22072 (N_22072,N_21338,N_21643);
nand U22073 (N_22073,N_21808,N_21191);
nand U22074 (N_22074,N_21090,N_21114);
xnor U22075 (N_22075,N_21936,N_21202);
nand U22076 (N_22076,N_21672,N_21650);
and U22077 (N_22077,N_21843,N_21354);
or U22078 (N_22078,N_21536,N_21318);
and U22079 (N_22079,N_21473,N_21477);
nor U22080 (N_22080,N_21515,N_21787);
or U22081 (N_22081,N_21761,N_21888);
nor U22082 (N_22082,N_21878,N_21939);
nor U22083 (N_22083,N_21017,N_21076);
nand U22084 (N_22084,N_21892,N_21099);
nor U22085 (N_22085,N_21615,N_21408);
and U22086 (N_22086,N_21821,N_21734);
xor U22087 (N_22087,N_21975,N_21050);
xor U22088 (N_22088,N_21188,N_21796);
nand U22089 (N_22089,N_21141,N_21924);
or U22090 (N_22090,N_21760,N_21901);
and U22091 (N_22091,N_21199,N_21332);
xnor U22092 (N_22092,N_21862,N_21331);
or U22093 (N_22093,N_21766,N_21563);
nor U22094 (N_22094,N_21602,N_21625);
nand U22095 (N_22095,N_21610,N_21883);
nand U22096 (N_22096,N_21570,N_21897);
nand U22097 (N_22097,N_21944,N_21684);
nand U22098 (N_22098,N_21105,N_21549);
and U22099 (N_22099,N_21502,N_21275);
xnor U22100 (N_22100,N_21206,N_21585);
or U22101 (N_22101,N_21077,N_21072);
nor U22102 (N_22102,N_21110,N_21540);
nand U22103 (N_22103,N_21947,N_21389);
or U22104 (N_22104,N_21474,N_21339);
or U22105 (N_22105,N_21904,N_21228);
nand U22106 (N_22106,N_21358,N_21287);
nand U22107 (N_22107,N_21520,N_21012);
nor U22108 (N_22108,N_21726,N_21677);
and U22109 (N_22109,N_21035,N_21930);
xnor U22110 (N_22110,N_21708,N_21227);
xnor U22111 (N_22111,N_21960,N_21542);
nand U22112 (N_22112,N_21621,N_21973);
xnor U22113 (N_22113,N_21184,N_21132);
nor U22114 (N_22114,N_21412,N_21470);
or U22115 (N_22115,N_21784,N_21309);
nor U22116 (N_22116,N_21703,N_21692);
nand U22117 (N_22117,N_21997,N_21544);
nand U22118 (N_22118,N_21998,N_21759);
nand U22119 (N_22119,N_21136,N_21416);
nor U22120 (N_22120,N_21229,N_21269);
or U22121 (N_22121,N_21879,N_21438);
nor U22122 (N_22122,N_21475,N_21154);
nor U22123 (N_22123,N_21903,N_21329);
nand U22124 (N_22124,N_21913,N_21375);
or U22125 (N_22125,N_21120,N_21179);
nand U22126 (N_22126,N_21770,N_21003);
xor U22127 (N_22127,N_21064,N_21834);
nor U22128 (N_22128,N_21592,N_21509);
or U22129 (N_22129,N_21264,N_21532);
or U22130 (N_22130,N_21245,N_21253);
nand U22131 (N_22131,N_21647,N_21974);
or U22132 (N_22132,N_21125,N_21583);
nor U22133 (N_22133,N_21815,N_21818);
or U22134 (N_22134,N_21950,N_21340);
xnor U22135 (N_22135,N_21089,N_21735);
nor U22136 (N_22136,N_21550,N_21022);
xnor U22137 (N_22137,N_21941,N_21838);
or U22138 (N_22138,N_21320,N_21813);
xor U22139 (N_22139,N_21378,N_21660);
and U22140 (N_22140,N_21776,N_21741);
or U22141 (N_22141,N_21249,N_21178);
nor U22142 (N_22142,N_21607,N_21046);
xnor U22143 (N_22143,N_21601,N_21402);
xor U22144 (N_22144,N_21538,N_21589);
or U22145 (N_22145,N_21926,N_21494);
and U22146 (N_22146,N_21982,N_21284);
nor U22147 (N_22147,N_21758,N_21307);
or U22148 (N_22148,N_21173,N_21094);
xor U22149 (N_22149,N_21492,N_21659);
or U22150 (N_22150,N_21261,N_21469);
or U22151 (N_22151,N_21788,N_21382);
and U22152 (N_22152,N_21780,N_21068);
nor U22153 (N_22153,N_21856,N_21194);
nand U22154 (N_22154,N_21561,N_21551);
or U22155 (N_22155,N_21485,N_21032);
and U22156 (N_22156,N_21066,N_21384);
nor U22157 (N_22157,N_21809,N_21078);
or U22158 (N_22158,N_21347,N_21140);
nor U22159 (N_22159,N_21365,N_21543);
nor U22160 (N_22160,N_21440,N_21744);
xnor U22161 (N_22161,N_21291,N_21546);
nor U22162 (N_22162,N_21451,N_21719);
xnor U22163 (N_22163,N_21326,N_21405);
nand U22164 (N_22164,N_21573,N_21966);
nand U22165 (N_22165,N_21633,N_21624);
xor U22166 (N_22166,N_21915,N_21595);
xor U22167 (N_22167,N_21505,N_21642);
xnor U22168 (N_22168,N_21733,N_21588);
xnor U22169 (N_22169,N_21021,N_21652);
nor U22170 (N_22170,N_21225,N_21409);
nand U22171 (N_22171,N_21335,N_21999);
and U22172 (N_22172,N_21518,N_21434);
nand U22173 (N_22173,N_21149,N_21424);
nand U22174 (N_22174,N_21895,N_21655);
xnor U22175 (N_22175,N_21547,N_21609);
and U22176 (N_22176,N_21096,N_21806);
nor U22177 (N_22177,N_21993,N_21101);
nand U22178 (N_22178,N_21819,N_21247);
nor U22179 (N_22179,N_21262,N_21860);
nand U22180 (N_22180,N_21321,N_21047);
and U22181 (N_22181,N_21627,N_21539);
xnor U22182 (N_22182,N_21209,N_21506);
or U22183 (N_22183,N_21432,N_21687);
xnor U22184 (N_22184,N_21436,N_21290);
nor U22185 (N_22185,N_21832,N_21422);
and U22186 (N_22186,N_21949,N_21980);
or U22187 (N_22187,N_21623,N_21311);
or U22188 (N_22188,N_21569,N_21131);
nor U22189 (N_22189,N_21466,N_21205);
and U22190 (N_22190,N_21374,N_21593);
and U22191 (N_22191,N_21155,N_21292);
nor U22192 (N_22192,N_21376,N_21908);
xnor U22193 (N_22193,N_21800,N_21619);
or U22194 (N_22194,N_21948,N_21403);
or U22195 (N_22195,N_21581,N_21545);
or U22196 (N_22196,N_21969,N_21560);
nor U22197 (N_22197,N_21246,N_21496);
or U22198 (N_22198,N_21727,N_21387);
and U22199 (N_22199,N_21350,N_21804);
xor U22200 (N_22200,N_21137,N_21454);
and U22201 (N_22201,N_21725,N_21854);
nor U22202 (N_22202,N_21273,N_21087);
xor U22203 (N_22203,N_21839,N_21256);
nand U22204 (N_22204,N_21598,N_21183);
and U22205 (N_22205,N_21270,N_21053);
nand U22206 (N_22206,N_21885,N_21482);
nand U22207 (N_22207,N_21305,N_21559);
xnor U22208 (N_22208,N_21337,N_21394);
or U22209 (N_22209,N_21989,N_21257);
nor U22210 (N_22210,N_21168,N_21083);
xnor U22211 (N_22211,N_21330,N_21323);
or U22212 (N_22212,N_21371,N_21210);
or U22213 (N_22213,N_21799,N_21812);
and U22214 (N_22214,N_21527,N_21461);
and U22215 (N_22215,N_21689,N_21940);
nor U22216 (N_22216,N_21366,N_21430);
or U22217 (N_22217,N_21180,N_21504);
or U22218 (N_22218,N_21754,N_21001);
and U22219 (N_22219,N_21840,N_21992);
or U22220 (N_22220,N_21251,N_21126);
or U22221 (N_22221,N_21828,N_21768);
or U22222 (N_22222,N_21979,N_21937);
and U22223 (N_22223,N_21919,N_21029);
and U22224 (N_22224,N_21724,N_21233);
xor U22225 (N_22225,N_21639,N_21413);
and U22226 (N_22226,N_21058,N_21669);
and U22227 (N_22227,N_21189,N_21781);
nand U22228 (N_22228,N_21617,N_21782);
nand U22229 (N_22229,N_21630,N_21678);
and U22230 (N_22230,N_21907,N_21632);
or U22231 (N_22231,N_21497,N_21605);
and U22232 (N_22232,N_21437,N_21055);
or U22233 (N_22233,N_21204,N_21283);
xor U22234 (N_22234,N_21674,N_21203);
and U22235 (N_22235,N_21103,N_21124);
nor U22236 (N_22236,N_21577,N_21170);
and U22237 (N_22237,N_21300,N_21235);
xor U22238 (N_22238,N_21359,N_21201);
or U22239 (N_22239,N_21801,N_21743);
nand U22240 (N_22240,N_21541,N_21565);
or U22241 (N_22241,N_21397,N_21272);
or U22242 (N_22242,N_21372,N_21399);
nor U22243 (N_22243,N_21830,N_21106);
nor U22244 (N_22244,N_21604,N_21267);
or U22245 (N_22245,N_21629,N_21938);
and U22246 (N_22246,N_21928,N_21763);
and U22247 (N_22247,N_21098,N_21691);
xnor U22248 (N_22248,N_21914,N_21961);
or U22249 (N_22249,N_21277,N_21680);
nor U22250 (N_22250,N_21729,N_21219);
nand U22251 (N_22251,N_21348,N_21135);
nand U22252 (N_22252,N_21934,N_21709);
or U22253 (N_22253,N_21837,N_21827);
or U22254 (N_22254,N_21968,N_21921);
xnor U22255 (N_22255,N_21108,N_21212);
or U22256 (N_22256,N_21278,N_21404);
nand U22257 (N_22257,N_21336,N_21312);
nand U22258 (N_22258,N_21833,N_21552);
nor U22259 (N_22259,N_21558,N_21556);
xor U22260 (N_22260,N_21195,N_21730);
nor U22261 (N_22261,N_21322,N_21048);
xor U22262 (N_22262,N_21060,N_21463);
and U22263 (N_22263,N_21297,N_21005);
xnor U22264 (N_22264,N_21844,N_21696);
nand U22265 (N_22265,N_21705,N_21442);
nand U22266 (N_22266,N_21360,N_21852);
nand U22267 (N_22267,N_21905,N_21835);
or U22268 (N_22268,N_21831,N_21435);
xnor U22269 (N_22269,N_21177,N_21157);
or U22270 (N_22270,N_21635,N_21158);
nor U22271 (N_22271,N_21608,N_21697);
nand U22272 (N_22272,N_21462,N_21008);
nand U22273 (N_22273,N_21122,N_21418);
nand U22274 (N_22274,N_21861,N_21313);
nor U22275 (N_22275,N_21649,N_21281);
or U22276 (N_22276,N_21486,N_21028);
and U22277 (N_22277,N_21067,N_21638);
nor U22278 (N_22278,N_21031,N_21484);
nand U22279 (N_22279,N_21749,N_21495);
nand U22280 (N_22280,N_21458,N_21093);
xor U22281 (N_22281,N_21015,N_21805);
nand U22282 (N_22282,N_21693,N_21241);
and U22283 (N_22283,N_21316,N_21407);
or U22284 (N_22284,N_21685,N_21386);
nand U22285 (N_22285,N_21823,N_21144);
nand U22286 (N_22286,N_21757,N_21590);
nor U22287 (N_22287,N_21186,N_21457);
and U22288 (N_22288,N_21453,N_21196);
xnor U22289 (N_22289,N_21258,N_21074);
nand U22290 (N_22290,N_21917,N_21620);
nand U22291 (N_22291,N_21824,N_21242);
or U22292 (N_22292,N_21185,N_21483);
and U22293 (N_22293,N_21503,N_21343);
nand U22294 (N_22294,N_21034,N_21769);
or U22295 (N_22295,N_21742,N_21065);
and U22296 (N_22296,N_21816,N_21234);
xor U22297 (N_22297,N_21952,N_21786);
nand U22298 (N_22298,N_21591,N_21159);
nand U22299 (N_22299,N_21481,N_21792);
nor U22300 (N_22300,N_21848,N_21712);
nor U22301 (N_22301,N_21841,N_21931);
and U22302 (N_22302,N_21798,N_21794);
nor U22303 (N_22303,N_21095,N_21498);
xor U22304 (N_22304,N_21344,N_21571);
nand U22305 (N_22305,N_21723,N_21148);
xor U22306 (N_22306,N_21452,N_21537);
and U22307 (N_22307,N_21765,N_21020);
nand U22308 (N_22308,N_21446,N_21584);
nand U22309 (N_22309,N_21164,N_21847);
nand U22310 (N_22310,N_21215,N_21075);
nor U22311 (N_22311,N_21162,N_21613);
or U22312 (N_22312,N_21679,N_21704);
nor U22313 (N_22313,N_21150,N_21328);
xor U22314 (N_22314,N_21829,N_21579);
or U22315 (N_22315,N_21699,N_21390);
and U22316 (N_22316,N_21027,N_21640);
or U22317 (N_22317,N_21460,N_21119);
nand U22318 (N_22318,N_21274,N_21773);
or U22319 (N_22319,N_21013,N_21129);
or U22320 (N_22320,N_21923,N_21167);
and U22321 (N_22321,N_21471,N_21807);
or U22322 (N_22322,N_21222,N_21063);
nand U22323 (N_22323,N_21260,N_21111);
or U22324 (N_22324,N_21884,N_21994);
xnor U22325 (N_22325,N_21675,N_21746);
or U22326 (N_22326,N_21052,N_21511);
or U22327 (N_22327,N_21049,N_21084);
nor U22328 (N_22328,N_21018,N_21271);
or U22329 (N_22329,N_21224,N_21207);
and U22330 (N_22330,N_21865,N_21200);
and U22331 (N_22331,N_21447,N_21282);
and U22332 (N_22332,N_21690,N_21785);
and U22333 (N_22333,N_21464,N_21123);
xnor U22334 (N_22334,N_21385,N_21134);
or U22335 (N_22335,N_21169,N_21526);
nand U22336 (N_22336,N_21088,N_21707);
and U22337 (N_22337,N_21706,N_21415);
nor U22338 (N_22338,N_21346,N_21868);
nand U22339 (N_22339,N_21426,N_21396);
xor U22340 (N_22340,N_21646,N_21102);
xnor U22341 (N_22341,N_21946,N_21889);
xnor U22342 (N_22342,N_21750,N_21513);
xnor U22343 (N_22343,N_21702,N_21756);
nand U22344 (N_22344,N_21880,N_21845);
nand U22345 (N_22345,N_21575,N_21391);
nor U22346 (N_22346,N_21059,N_21252);
xor U22347 (N_22347,N_21716,N_21298);
xnor U22348 (N_22348,N_21962,N_21739);
nand U22349 (N_22349,N_21817,N_21182);
nand U22350 (N_22350,N_21181,N_21500);
and U22351 (N_22351,N_21942,N_21152);
xnor U22352 (N_22352,N_21187,N_21671);
nor U22353 (N_22353,N_21286,N_21172);
or U22354 (N_22354,N_21487,N_21894);
nor U22355 (N_22355,N_21682,N_21315);
or U22356 (N_22356,N_21045,N_21755);
nand U22357 (N_22357,N_21606,N_21459);
or U22358 (N_22358,N_21752,N_21700);
and U22359 (N_22359,N_21963,N_21395);
nand U22360 (N_22360,N_21873,N_21231);
nand U22361 (N_22361,N_21214,N_21218);
xnor U22362 (N_22362,N_21398,N_21349);
xnor U22363 (N_22363,N_21491,N_21523);
and U22364 (N_22364,N_21056,N_21911);
and U22365 (N_22365,N_21073,N_21236);
or U22366 (N_22366,N_21618,N_21568);
xnor U22367 (N_22367,N_21925,N_21368);
or U22368 (N_22368,N_21280,N_21803);
nor U22369 (N_22369,N_21751,N_21996);
nand U22370 (N_22370,N_21811,N_21855);
or U22371 (N_22371,N_21717,N_21964);
xor U22372 (N_22372,N_21293,N_21455);
and U22373 (N_22373,N_21142,N_21043);
nand U22374 (N_22374,N_21145,N_21825);
or U22375 (N_22375,N_21519,N_21775);
and U22376 (N_22376,N_21317,N_21955);
and U22377 (N_22377,N_21853,N_21871);
xor U22378 (N_22378,N_21648,N_21732);
xnor U22379 (N_22379,N_21866,N_21562);
nand U22380 (N_22380,N_21334,N_21753);
nand U22381 (N_22381,N_21651,N_21082);
or U22382 (N_22382,N_21423,N_21736);
nand U22383 (N_22383,N_21208,N_21092);
nor U22384 (N_22384,N_21567,N_21450);
nand U22385 (N_22385,N_21701,N_21918);
or U22386 (N_22386,N_21920,N_21299);
and U22387 (N_22387,N_21533,N_21238);
or U22388 (N_22388,N_21276,N_21211);
xor U22389 (N_22389,N_21747,N_21294);
nor U22390 (N_22390,N_21514,N_21899);
nand U22391 (N_22391,N_21932,N_21239);
xor U22392 (N_22392,N_21070,N_21327);
nand U22393 (N_22393,N_21265,N_21421);
or U22394 (N_22394,N_21370,N_21051);
or U22395 (N_22395,N_21985,N_21681);
and U22396 (N_22396,N_21025,N_21314);
nor U22397 (N_22397,N_21731,N_21176);
and U22398 (N_22398,N_21587,N_21666);
and U22399 (N_22399,N_21373,N_21118);
nor U22400 (N_22400,N_21886,N_21393);
and U22401 (N_22401,N_21417,N_21130);
and U22402 (N_22402,N_21572,N_21887);
nor U22403 (N_22403,N_21851,N_21429);
and U22404 (N_22404,N_21490,N_21363);
or U22405 (N_22405,N_21456,N_21042);
nor U22406 (N_22406,N_21302,N_21156);
and U22407 (N_22407,N_21044,N_21984);
or U22408 (N_22408,N_21916,N_21420);
nand U22409 (N_22409,N_21566,N_21288);
and U22410 (N_22410,N_21367,N_21721);
nor U22411 (N_22411,N_21138,N_21772);
or U22412 (N_22412,N_21983,N_21472);
xor U22413 (N_22413,N_21594,N_21943);
xor U22414 (N_22414,N_21673,N_21745);
xor U22415 (N_22415,N_21867,N_21531);
or U22416 (N_22416,N_21870,N_21151);
and U22417 (N_22417,N_21995,N_21990);
or U22418 (N_22418,N_21388,N_21872);
nand U22419 (N_22419,N_21411,N_21146);
xor U22420 (N_22420,N_21597,N_21100);
and U22421 (N_22421,N_21445,N_21790);
or U22422 (N_22422,N_21728,N_21392);
or U22423 (N_22423,N_21217,N_21714);
nor U22424 (N_22424,N_21576,N_21849);
nand U22425 (N_22425,N_21970,N_21778);
nand U22426 (N_22426,N_21061,N_21147);
xor U22427 (N_22427,N_21171,N_21836);
nand U22428 (N_22428,N_21006,N_21112);
and U22429 (N_22429,N_21722,N_21250);
nand U22430 (N_22430,N_21842,N_21308);
or U22431 (N_22431,N_21516,N_21857);
nor U22432 (N_22432,N_21023,N_21814);
and U22433 (N_22433,N_21616,N_21319);
nand U22434 (N_22434,N_21081,N_21226);
nand U22435 (N_22435,N_21791,N_21564);
xor U22436 (N_22436,N_21554,N_21991);
nand U22437 (N_22437,N_21439,N_21555);
and U22438 (N_22438,N_21694,N_21797);
and U22439 (N_22439,N_21662,N_21153);
or U22440 (N_22440,N_21381,N_21107);
xnor U22441 (N_22441,N_21688,N_21109);
and U22442 (N_22442,N_21113,N_21425);
and U22443 (N_22443,N_21036,N_21342);
and U22444 (N_22444,N_21986,N_21240);
or U22445 (N_22445,N_21165,N_21400);
nand U22446 (N_22446,N_21266,N_21127);
nand U22447 (N_22447,N_21737,N_21959);
and U22448 (N_22448,N_21876,N_21657);
and U22449 (N_22449,N_21000,N_21715);
and U22450 (N_22450,N_21139,N_21232);
and U22451 (N_22451,N_21216,N_21121);
xnor U22452 (N_22452,N_21133,N_21912);
or U22453 (N_22453,N_21612,N_21002);
nor U22454 (N_22454,N_21951,N_21987);
xor U22455 (N_22455,N_21353,N_21237);
nor U22456 (N_22456,N_21301,N_21676);
xnor U22457 (N_22457,N_21414,N_21448);
xnor U22458 (N_22458,N_21653,N_21324);
or U22459 (N_22459,N_21352,N_21864);
nand U22460 (N_22460,N_21713,N_21379);
xor U22461 (N_22461,N_21881,N_21345);
nand U22462 (N_22462,N_21026,N_21419);
nor U22463 (N_22463,N_21664,N_21521);
nor U22464 (N_22464,N_21710,N_21553);
xor U22465 (N_22465,N_21304,N_21467);
xnor U22466 (N_22466,N_21902,N_21444);
and U22467 (N_22467,N_21525,N_21488);
nor U22468 (N_22468,N_21614,N_21774);
nor U22469 (N_22469,N_21040,N_21255);
or U22470 (N_22470,N_21846,N_21686);
nand U22471 (N_22471,N_21631,N_21333);
and U22472 (N_22472,N_21057,N_21254);
and U22473 (N_22473,N_21740,N_21874);
and U22474 (N_22474,N_21935,N_21965);
xnor U22475 (N_22475,N_21193,N_21771);
and U22476 (N_22476,N_21303,N_21698);
nor U22477 (N_22477,N_21654,N_21548);
xor U22478 (N_22478,N_21978,N_21441);
or U22479 (N_22479,N_21306,N_21822);
xnor U22480 (N_22480,N_21762,N_21695);
and U22481 (N_22481,N_21221,N_21041);
and U22482 (N_22482,N_21530,N_21882);
xnor U22483 (N_22483,N_21097,N_21033);
nor U22484 (N_22484,N_21080,N_21557);
and U22485 (N_22485,N_21958,N_21296);
nor U22486 (N_22486,N_21783,N_21859);
nand U22487 (N_22487,N_21512,N_21795);
nand U22488 (N_22488,N_21711,N_21580);
xnor U22489 (N_22489,N_21489,N_21355);
xor U22490 (N_22490,N_21645,N_21578);
nor U22491 (N_22491,N_21720,N_21636);
nand U22492 (N_22492,N_21259,N_21957);
and U22493 (N_22493,N_21976,N_21764);
nor U22494 (N_22494,N_21909,N_21517);
nor U22495 (N_22495,N_21665,N_21038);
nor U22496 (N_22496,N_21091,N_21596);
nand U22497 (N_22497,N_21954,N_21820);
nor U22498 (N_22498,N_21670,N_21325);
nor U22499 (N_22499,N_21988,N_21929);
nor U22500 (N_22500,N_21732,N_21214);
and U22501 (N_22501,N_21333,N_21256);
or U22502 (N_22502,N_21612,N_21842);
nand U22503 (N_22503,N_21855,N_21183);
or U22504 (N_22504,N_21876,N_21252);
or U22505 (N_22505,N_21682,N_21485);
and U22506 (N_22506,N_21521,N_21950);
nor U22507 (N_22507,N_21519,N_21157);
nand U22508 (N_22508,N_21017,N_21850);
or U22509 (N_22509,N_21492,N_21543);
nand U22510 (N_22510,N_21423,N_21921);
xnor U22511 (N_22511,N_21387,N_21771);
and U22512 (N_22512,N_21313,N_21807);
nand U22513 (N_22513,N_21295,N_21818);
or U22514 (N_22514,N_21572,N_21351);
and U22515 (N_22515,N_21423,N_21494);
and U22516 (N_22516,N_21470,N_21924);
xnor U22517 (N_22517,N_21035,N_21875);
and U22518 (N_22518,N_21090,N_21578);
nand U22519 (N_22519,N_21949,N_21266);
nor U22520 (N_22520,N_21254,N_21509);
nor U22521 (N_22521,N_21573,N_21451);
and U22522 (N_22522,N_21189,N_21289);
xor U22523 (N_22523,N_21266,N_21003);
nand U22524 (N_22524,N_21684,N_21965);
xnor U22525 (N_22525,N_21637,N_21597);
nand U22526 (N_22526,N_21069,N_21963);
nor U22527 (N_22527,N_21707,N_21668);
and U22528 (N_22528,N_21296,N_21175);
nand U22529 (N_22529,N_21868,N_21729);
and U22530 (N_22530,N_21399,N_21247);
or U22531 (N_22531,N_21511,N_21492);
nor U22532 (N_22532,N_21512,N_21308);
nor U22533 (N_22533,N_21403,N_21681);
xor U22534 (N_22534,N_21082,N_21847);
and U22535 (N_22535,N_21484,N_21680);
or U22536 (N_22536,N_21192,N_21934);
nand U22537 (N_22537,N_21446,N_21865);
or U22538 (N_22538,N_21824,N_21473);
nand U22539 (N_22539,N_21923,N_21404);
or U22540 (N_22540,N_21513,N_21517);
and U22541 (N_22541,N_21565,N_21672);
or U22542 (N_22542,N_21224,N_21717);
or U22543 (N_22543,N_21748,N_21569);
or U22544 (N_22544,N_21122,N_21788);
nand U22545 (N_22545,N_21412,N_21430);
nor U22546 (N_22546,N_21295,N_21577);
and U22547 (N_22547,N_21983,N_21466);
or U22548 (N_22548,N_21000,N_21344);
xnor U22549 (N_22549,N_21817,N_21013);
or U22550 (N_22550,N_21803,N_21057);
and U22551 (N_22551,N_21831,N_21811);
nand U22552 (N_22552,N_21096,N_21148);
and U22553 (N_22553,N_21483,N_21793);
or U22554 (N_22554,N_21740,N_21003);
nor U22555 (N_22555,N_21392,N_21282);
nor U22556 (N_22556,N_21639,N_21551);
or U22557 (N_22557,N_21202,N_21960);
xor U22558 (N_22558,N_21936,N_21331);
and U22559 (N_22559,N_21487,N_21723);
xor U22560 (N_22560,N_21909,N_21991);
nor U22561 (N_22561,N_21317,N_21899);
nand U22562 (N_22562,N_21303,N_21480);
nor U22563 (N_22563,N_21709,N_21813);
nand U22564 (N_22564,N_21257,N_21649);
nand U22565 (N_22565,N_21194,N_21263);
and U22566 (N_22566,N_21621,N_21145);
nand U22567 (N_22567,N_21644,N_21065);
nand U22568 (N_22568,N_21860,N_21505);
or U22569 (N_22569,N_21032,N_21082);
nor U22570 (N_22570,N_21383,N_21048);
or U22571 (N_22571,N_21538,N_21077);
and U22572 (N_22572,N_21261,N_21209);
nand U22573 (N_22573,N_21698,N_21064);
xnor U22574 (N_22574,N_21258,N_21029);
xnor U22575 (N_22575,N_21581,N_21009);
or U22576 (N_22576,N_21603,N_21529);
or U22577 (N_22577,N_21880,N_21553);
nor U22578 (N_22578,N_21286,N_21136);
or U22579 (N_22579,N_21064,N_21606);
xor U22580 (N_22580,N_21915,N_21738);
nor U22581 (N_22581,N_21627,N_21507);
and U22582 (N_22582,N_21318,N_21158);
or U22583 (N_22583,N_21500,N_21705);
nor U22584 (N_22584,N_21456,N_21537);
nand U22585 (N_22585,N_21874,N_21295);
nand U22586 (N_22586,N_21942,N_21696);
nor U22587 (N_22587,N_21077,N_21644);
nand U22588 (N_22588,N_21502,N_21196);
nor U22589 (N_22589,N_21206,N_21235);
and U22590 (N_22590,N_21176,N_21813);
nand U22591 (N_22591,N_21664,N_21044);
nand U22592 (N_22592,N_21158,N_21319);
nand U22593 (N_22593,N_21194,N_21232);
or U22594 (N_22594,N_21325,N_21203);
or U22595 (N_22595,N_21615,N_21860);
or U22596 (N_22596,N_21990,N_21832);
nand U22597 (N_22597,N_21734,N_21429);
xnor U22598 (N_22598,N_21317,N_21793);
nand U22599 (N_22599,N_21019,N_21739);
nor U22600 (N_22600,N_21567,N_21654);
nand U22601 (N_22601,N_21280,N_21370);
nand U22602 (N_22602,N_21485,N_21873);
nor U22603 (N_22603,N_21715,N_21279);
nor U22604 (N_22604,N_21298,N_21502);
nor U22605 (N_22605,N_21956,N_21358);
and U22606 (N_22606,N_21765,N_21589);
and U22607 (N_22607,N_21004,N_21692);
nor U22608 (N_22608,N_21298,N_21781);
nand U22609 (N_22609,N_21174,N_21007);
and U22610 (N_22610,N_21884,N_21347);
and U22611 (N_22611,N_21733,N_21060);
or U22612 (N_22612,N_21830,N_21187);
nor U22613 (N_22613,N_21621,N_21611);
and U22614 (N_22614,N_21902,N_21399);
nand U22615 (N_22615,N_21270,N_21518);
xor U22616 (N_22616,N_21457,N_21615);
xor U22617 (N_22617,N_21279,N_21194);
or U22618 (N_22618,N_21694,N_21061);
nand U22619 (N_22619,N_21611,N_21517);
or U22620 (N_22620,N_21996,N_21529);
xnor U22621 (N_22621,N_21700,N_21745);
xnor U22622 (N_22622,N_21121,N_21700);
or U22623 (N_22623,N_21000,N_21890);
nand U22624 (N_22624,N_21921,N_21960);
xor U22625 (N_22625,N_21341,N_21421);
xor U22626 (N_22626,N_21361,N_21753);
xnor U22627 (N_22627,N_21079,N_21674);
nand U22628 (N_22628,N_21989,N_21399);
xnor U22629 (N_22629,N_21057,N_21996);
or U22630 (N_22630,N_21361,N_21812);
nand U22631 (N_22631,N_21103,N_21479);
nand U22632 (N_22632,N_21459,N_21350);
xnor U22633 (N_22633,N_21797,N_21300);
and U22634 (N_22634,N_21661,N_21452);
and U22635 (N_22635,N_21943,N_21964);
nor U22636 (N_22636,N_21245,N_21104);
and U22637 (N_22637,N_21638,N_21920);
nand U22638 (N_22638,N_21798,N_21510);
and U22639 (N_22639,N_21419,N_21933);
xor U22640 (N_22640,N_21196,N_21697);
xnor U22641 (N_22641,N_21520,N_21699);
and U22642 (N_22642,N_21915,N_21837);
nor U22643 (N_22643,N_21335,N_21294);
nand U22644 (N_22644,N_21751,N_21522);
nor U22645 (N_22645,N_21440,N_21587);
or U22646 (N_22646,N_21913,N_21058);
and U22647 (N_22647,N_21209,N_21802);
nand U22648 (N_22648,N_21502,N_21699);
or U22649 (N_22649,N_21829,N_21904);
nand U22650 (N_22650,N_21755,N_21528);
or U22651 (N_22651,N_21095,N_21816);
or U22652 (N_22652,N_21784,N_21196);
nand U22653 (N_22653,N_21161,N_21671);
nand U22654 (N_22654,N_21403,N_21409);
nor U22655 (N_22655,N_21208,N_21096);
and U22656 (N_22656,N_21147,N_21644);
or U22657 (N_22657,N_21477,N_21214);
xor U22658 (N_22658,N_21741,N_21711);
nand U22659 (N_22659,N_21200,N_21613);
nand U22660 (N_22660,N_21739,N_21313);
nor U22661 (N_22661,N_21587,N_21352);
nand U22662 (N_22662,N_21944,N_21188);
and U22663 (N_22663,N_21641,N_21334);
nand U22664 (N_22664,N_21424,N_21952);
and U22665 (N_22665,N_21461,N_21690);
nor U22666 (N_22666,N_21154,N_21695);
nor U22667 (N_22667,N_21978,N_21428);
nor U22668 (N_22668,N_21900,N_21619);
or U22669 (N_22669,N_21372,N_21003);
nor U22670 (N_22670,N_21986,N_21270);
xor U22671 (N_22671,N_21228,N_21708);
xor U22672 (N_22672,N_21821,N_21724);
and U22673 (N_22673,N_21534,N_21151);
or U22674 (N_22674,N_21477,N_21273);
or U22675 (N_22675,N_21890,N_21912);
or U22676 (N_22676,N_21460,N_21199);
or U22677 (N_22677,N_21006,N_21294);
nor U22678 (N_22678,N_21901,N_21664);
nor U22679 (N_22679,N_21550,N_21539);
or U22680 (N_22680,N_21800,N_21563);
or U22681 (N_22681,N_21180,N_21134);
or U22682 (N_22682,N_21858,N_21947);
nand U22683 (N_22683,N_21545,N_21307);
xor U22684 (N_22684,N_21564,N_21152);
xnor U22685 (N_22685,N_21072,N_21850);
nand U22686 (N_22686,N_21284,N_21413);
nand U22687 (N_22687,N_21336,N_21500);
and U22688 (N_22688,N_21877,N_21693);
xnor U22689 (N_22689,N_21632,N_21765);
nor U22690 (N_22690,N_21719,N_21717);
or U22691 (N_22691,N_21826,N_21843);
and U22692 (N_22692,N_21767,N_21427);
and U22693 (N_22693,N_21593,N_21487);
nand U22694 (N_22694,N_21626,N_21868);
and U22695 (N_22695,N_21565,N_21217);
and U22696 (N_22696,N_21494,N_21615);
or U22697 (N_22697,N_21163,N_21882);
xnor U22698 (N_22698,N_21618,N_21600);
xor U22699 (N_22699,N_21919,N_21954);
or U22700 (N_22700,N_21684,N_21184);
nor U22701 (N_22701,N_21696,N_21760);
and U22702 (N_22702,N_21608,N_21808);
nand U22703 (N_22703,N_21251,N_21230);
xor U22704 (N_22704,N_21369,N_21480);
nand U22705 (N_22705,N_21255,N_21337);
nand U22706 (N_22706,N_21845,N_21625);
and U22707 (N_22707,N_21059,N_21558);
nor U22708 (N_22708,N_21973,N_21855);
or U22709 (N_22709,N_21225,N_21060);
nor U22710 (N_22710,N_21079,N_21403);
nor U22711 (N_22711,N_21922,N_21130);
nor U22712 (N_22712,N_21583,N_21820);
xnor U22713 (N_22713,N_21550,N_21810);
or U22714 (N_22714,N_21247,N_21317);
nor U22715 (N_22715,N_21509,N_21024);
xnor U22716 (N_22716,N_21858,N_21227);
xor U22717 (N_22717,N_21455,N_21506);
xor U22718 (N_22718,N_21893,N_21630);
nor U22719 (N_22719,N_21105,N_21930);
nand U22720 (N_22720,N_21003,N_21575);
nor U22721 (N_22721,N_21520,N_21500);
nor U22722 (N_22722,N_21758,N_21131);
xor U22723 (N_22723,N_21199,N_21515);
nand U22724 (N_22724,N_21842,N_21633);
nor U22725 (N_22725,N_21883,N_21260);
xnor U22726 (N_22726,N_21175,N_21047);
or U22727 (N_22727,N_21823,N_21994);
xor U22728 (N_22728,N_21129,N_21904);
xnor U22729 (N_22729,N_21355,N_21923);
and U22730 (N_22730,N_21844,N_21950);
nand U22731 (N_22731,N_21657,N_21965);
nand U22732 (N_22732,N_21453,N_21677);
xor U22733 (N_22733,N_21689,N_21601);
or U22734 (N_22734,N_21891,N_21832);
nor U22735 (N_22735,N_21981,N_21417);
nor U22736 (N_22736,N_21802,N_21594);
or U22737 (N_22737,N_21024,N_21448);
nand U22738 (N_22738,N_21887,N_21047);
xor U22739 (N_22739,N_21305,N_21591);
or U22740 (N_22740,N_21860,N_21409);
xnor U22741 (N_22741,N_21934,N_21632);
and U22742 (N_22742,N_21702,N_21076);
nor U22743 (N_22743,N_21953,N_21743);
or U22744 (N_22744,N_21797,N_21698);
and U22745 (N_22745,N_21894,N_21759);
nand U22746 (N_22746,N_21044,N_21748);
nand U22747 (N_22747,N_21193,N_21427);
and U22748 (N_22748,N_21319,N_21735);
and U22749 (N_22749,N_21431,N_21880);
and U22750 (N_22750,N_21069,N_21734);
nor U22751 (N_22751,N_21053,N_21907);
and U22752 (N_22752,N_21547,N_21409);
xnor U22753 (N_22753,N_21978,N_21214);
or U22754 (N_22754,N_21206,N_21937);
nor U22755 (N_22755,N_21986,N_21326);
xor U22756 (N_22756,N_21558,N_21147);
nor U22757 (N_22757,N_21123,N_21615);
or U22758 (N_22758,N_21118,N_21274);
xnor U22759 (N_22759,N_21546,N_21302);
nor U22760 (N_22760,N_21473,N_21384);
nand U22761 (N_22761,N_21104,N_21102);
xor U22762 (N_22762,N_21086,N_21445);
or U22763 (N_22763,N_21217,N_21155);
xnor U22764 (N_22764,N_21500,N_21145);
xnor U22765 (N_22765,N_21512,N_21143);
xnor U22766 (N_22766,N_21861,N_21824);
nand U22767 (N_22767,N_21816,N_21140);
or U22768 (N_22768,N_21262,N_21187);
nand U22769 (N_22769,N_21894,N_21383);
xnor U22770 (N_22770,N_21738,N_21778);
xnor U22771 (N_22771,N_21532,N_21948);
nor U22772 (N_22772,N_21348,N_21532);
xor U22773 (N_22773,N_21109,N_21346);
and U22774 (N_22774,N_21063,N_21711);
and U22775 (N_22775,N_21598,N_21746);
nand U22776 (N_22776,N_21204,N_21310);
nand U22777 (N_22777,N_21366,N_21473);
nor U22778 (N_22778,N_21155,N_21460);
or U22779 (N_22779,N_21918,N_21157);
nand U22780 (N_22780,N_21740,N_21242);
or U22781 (N_22781,N_21446,N_21229);
nand U22782 (N_22782,N_21591,N_21728);
xor U22783 (N_22783,N_21460,N_21364);
xor U22784 (N_22784,N_21476,N_21500);
nand U22785 (N_22785,N_21893,N_21602);
xnor U22786 (N_22786,N_21277,N_21240);
nor U22787 (N_22787,N_21397,N_21908);
nor U22788 (N_22788,N_21088,N_21038);
xnor U22789 (N_22789,N_21860,N_21395);
xor U22790 (N_22790,N_21189,N_21447);
or U22791 (N_22791,N_21082,N_21684);
or U22792 (N_22792,N_21827,N_21025);
and U22793 (N_22793,N_21276,N_21969);
nand U22794 (N_22794,N_21174,N_21277);
nand U22795 (N_22795,N_21045,N_21441);
nand U22796 (N_22796,N_21320,N_21118);
and U22797 (N_22797,N_21369,N_21610);
nor U22798 (N_22798,N_21240,N_21668);
xnor U22799 (N_22799,N_21169,N_21155);
nor U22800 (N_22800,N_21635,N_21529);
nand U22801 (N_22801,N_21149,N_21385);
nor U22802 (N_22802,N_21303,N_21611);
nand U22803 (N_22803,N_21370,N_21235);
and U22804 (N_22804,N_21867,N_21118);
xnor U22805 (N_22805,N_21509,N_21433);
nor U22806 (N_22806,N_21510,N_21758);
nor U22807 (N_22807,N_21987,N_21649);
xor U22808 (N_22808,N_21124,N_21134);
nor U22809 (N_22809,N_21795,N_21045);
nand U22810 (N_22810,N_21913,N_21554);
xnor U22811 (N_22811,N_21966,N_21412);
xnor U22812 (N_22812,N_21849,N_21518);
nor U22813 (N_22813,N_21181,N_21378);
nor U22814 (N_22814,N_21351,N_21988);
or U22815 (N_22815,N_21723,N_21535);
nand U22816 (N_22816,N_21733,N_21093);
or U22817 (N_22817,N_21612,N_21145);
nor U22818 (N_22818,N_21911,N_21712);
xor U22819 (N_22819,N_21265,N_21950);
nand U22820 (N_22820,N_21493,N_21211);
and U22821 (N_22821,N_21211,N_21786);
xnor U22822 (N_22822,N_21442,N_21563);
or U22823 (N_22823,N_21615,N_21689);
nor U22824 (N_22824,N_21406,N_21346);
and U22825 (N_22825,N_21277,N_21178);
and U22826 (N_22826,N_21373,N_21722);
nor U22827 (N_22827,N_21670,N_21480);
or U22828 (N_22828,N_21598,N_21467);
nand U22829 (N_22829,N_21689,N_21490);
and U22830 (N_22830,N_21024,N_21695);
or U22831 (N_22831,N_21257,N_21055);
or U22832 (N_22832,N_21082,N_21361);
and U22833 (N_22833,N_21592,N_21276);
and U22834 (N_22834,N_21220,N_21069);
xor U22835 (N_22835,N_21542,N_21365);
and U22836 (N_22836,N_21837,N_21736);
nand U22837 (N_22837,N_21295,N_21967);
nor U22838 (N_22838,N_21370,N_21293);
nand U22839 (N_22839,N_21225,N_21312);
nand U22840 (N_22840,N_21793,N_21637);
xnor U22841 (N_22841,N_21740,N_21577);
nand U22842 (N_22842,N_21276,N_21682);
nor U22843 (N_22843,N_21266,N_21992);
or U22844 (N_22844,N_21280,N_21830);
nand U22845 (N_22845,N_21614,N_21802);
nor U22846 (N_22846,N_21999,N_21124);
or U22847 (N_22847,N_21040,N_21106);
nor U22848 (N_22848,N_21789,N_21122);
xnor U22849 (N_22849,N_21721,N_21660);
xnor U22850 (N_22850,N_21750,N_21054);
xor U22851 (N_22851,N_21973,N_21328);
and U22852 (N_22852,N_21270,N_21108);
nor U22853 (N_22853,N_21836,N_21647);
nor U22854 (N_22854,N_21943,N_21156);
and U22855 (N_22855,N_21092,N_21214);
or U22856 (N_22856,N_21858,N_21926);
nand U22857 (N_22857,N_21465,N_21318);
xnor U22858 (N_22858,N_21625,N_21174);
nand U22859 (N_22859,N_21287,N_21991);
nand U22860 (N_22860,N_21220,N_21593);
xor U22861 (N_22861,N_21399,N_21167);
xnor U22862 (N_22862,N_21722,N_21650);
xnor U22863 (N_22863,N_21627,N_21656);
nand U22864 (N_22864,N_21859,N_21276);
nand U22865 (N_22865,N_21109,N_21464);
xor U22866 (N_22866,N_21709,N_21694);
nand U22867 (N_22867,N_21267,N_21154);
xor U22868 (N_22868,N_21187,N_21217);
nor U22869 (N_22869,N_21178,N_21241);
and U22870 (N_22870,N_21631,N_21299);
and U22871 (N_22871,N_21192,N_21614);
or U22872 (N_22872,N_21196,N_21799);
nor U22873 (N_22873,N_21378,N_21914);
xnor U22874 (N_22874,N_21264,N_21936);
or U22875 (N_22875,N_21915,N_21071);
and U22876 (N_22876,N_21589,N_21568);
or U22877 (N_22877,N_21068,N_21893);
and U22878 (N_22878,N_21290,N_21872);
or U22879 (N_22879,N_21049,N_21609);
nand U22880 (N_22880,N_21484,N_21280);
xor U22881 (N_22881,N_21811,N_21853);
and U22882 (N_22882,N_21761,N_21880);
or U22883 (N_22883,N_21922,N_21903);
or U22884 (N_22884,N_21568,N_21895);
or U22885 (N_22885,N_21119,N_21354);
or U22886 (N_22886,N_21933,N_21798);
nor U22887 (N_22887,N_21646,N_21327);
xor U22888 (N_22888,N_21387,N_21826);
or U22889 (N_22889,N_21873,N_21160);
and U22890 (N_22890,N_21268,N_21761);
xnor U22891 (N_22891,N_21435,N_21059);
and U22892 (N_22892,N_21924,N_21143);
xnor U22893 (N_22893,N_21943,N_21314);
xnor U22894 (N_22894,N_21526,N_21881);
nor U22895 (N_22895,N_21617,N_21042);
and U22896 (N_22896,N_21412,N_21382);
nor U22897 (N_22897,N_21853,N_21172);
nand U22898 (N_22898,N_21807,N_21339);
or U22899 (N_22899,N_21349,N_21918);
xor U22900 (N_22900,N_21510,N_21685);
nand U22901 (N_22901,N_21195,N_21525);
or U22902 (N_22902,N_21812,N_21892);
or U22903 (N_22903,N_21673,N_21403);
or U22904 (N_22904,N_21566,N_21035);
nor U22905 (N_22905,N_21531,N_21860);
or U22906 (N_22906,N_21666,N_21918);
or U22907 (N_22907,N_21525,N_21957);
and U22908 (N_22908,N_21300,N_21573);
nor U22909 (N_22909,N_21328,N_21376);
nor U22910 (N_22910,N_21360,N_21516);
xnor U22911 (N_22911,N_21213,N_21718);
nor U22912 (N_22912,N_21152,N_21914);
or U22913 (N_22913,N_21826,N_21259);
xnor U22914 (N_22914,N_21104,N_21522);
nor U22915 (N_22915,N_21118,N_21292);
and U22916 (N_22916,N_21851,N_21607);
or U22917 (N_22917,N_21354,N_21884);
nor U22918 (N_22918,N_21894,N_21549);
or U22919 (N_22919,N_21195,N_21350);
xnor U22920 (N_22920,N_21114,N_21785);
or U22921 (N_22921,N_21455,N_21320);
xnor U22922 (N_22922,N_21864,N_21291);
or U22923 (N_22923,N_21717,N_21864);
nor U22924 (N_22924,N_21448,N_21570);
and U22925 (N_22925,N_21283,N_21060);
nor U22926 (N_22926,N_21840,N_21448);
nand U22927 (N_22927,N_21649,N_21886);
xnor U22928 (N_22928,N_21004,N_21851);
and U22929 (N_22929,N_21534,N_21161);
or U22930 (N_22930,N_21496,N_21037);
or U22931 (N_22931,N_21393,N_21883);
or U22932 (N_22932,N_21084,N_21006);
or U22933 (N_22933,N_21286,N_21348);
and U22934 (N_22934,N_21485,N_21724);
and U22935 (N_22935,N_21410,N_21137);
and U22936 (N_22936,N_21090,N_21974);
nor U22937 (N_22937,N_21919,N_21253);
or U22938 (N_22938,N_21405,N_21368);
nand U22939 (N_22939,N_21938,N_21028);
and U22940 (N_22940,N_21576,N_21133);
xnor U22941 (N_22941,N_21295,N_21786);
xor U22942 (N_22942,N_21261,N_21802);
nor U22943 (N_22943,N_21426,N_21916);
xor U22944 (N_22944,N_21118,N_21960);
xor U22945 (N_22945,N_21658,N_21815);
xnor U22946 (N_22946,N_21791,N_21452);
nor U22947 (N_22947,N_21993,N_21706);
xor U22948 (N_22948,N_21600,N_21575);
nor U22949 (N_22949,N_21283,N_21030);
xnor U22950 (N_22950,N_21249,N_21609);
or U22951 (N_22951,N_21159,N_21264);
or U22952 (N_22952,N_21624,N_21049);
xor U22953 (N_22953,N_21091,N_21353);
and U22954 (N_22954,N_21927,N_21989);
nand U22955 (N_22955,N_21470,N_21203);
and U22956 (N_22956,N_21991,N_21502);
or U22957 (N_22957,N_21399,N_21448);
xor U22958 (N_22958,N_21805,N_21556);
or U22959 (N_22959,N_21476,N_21967);
or U22960 (N_22960,N_21595,N_21376);
or U22961 (N_22961,N_21666,N_21638);
and U22962 (N_22962,N_21151,N_21545);
or U22963 (N_22963,N_21383,N_21025);
nand U22964 (N_22964,N_21911,N_21311);
nand U22965 (N_22965,N_21527,N_21376);
or U22966 (N_22966,N_21090,N_21943);
nand U22967 (N_22967,N_21757,N_21181);
or U22968 (N_22968,N_21827,N_21011);
nor U22969 (N_22969,N_21439,N_21591);
xor U22970 (N_22970,N_21207,N_21663);
or U22971 (N_22971,N_21012,N_21891);
or U22972 (N_22972,N_21208,N_21730);
or U22973 (N_22973,N_21704,N_21683);
nor U22974 (N_22974,N_21433,N_21967);
or U22975 (N_22975,N_21862,N_21797);
nand U22976 (N_22976,N_21919,N_21220);
and U22977 (N_22977,N_21460,N_21501);
nor U22978 (N_22978,N_21118,N_21849);
xor U22979 (N_22979,N_21567,N_21833);
xor U22980 (N_22980,N_21643,N_21665);
nand U22981 (N_22981,N_21327,N_21914);
and U22982 (N_22982,N_21639,N_21458);
or U22983 (N_22983,N_21452,N_21511);
and U22984 (N_22984,N_21018,N_21725);
xnor U22985 (N_22985,N_21912,N_21042);
and U22986 (N_22986,N_21749,N_21038);
and U22987 (N_22987,N_21897,N_21620);
nand U22988 (N_22988,N_21663,N_21370);
nor U22989 (N_22989,N_21756,N_21959);
xor U22990 (N_22990,N_21362,N_21792);
or U22991 (N_22991,N_21982,N_21693);
or U22992 (N_22992,N_21552,N_21013);
and U22993 (N_22993,N_21991,N_21096);
xor U22994 (N_22994,N_21664,N_21698);
nand U22995 (N_22995,N_21850,N_21695);
or U22996 (N_22996,N_21723,N_21503);
and U22997 (N_22997,N_21391,N_21990);
nor U22998 (N_22998,N_21052,N_21687);
nor U22999 (N_22999,N_21353,N_21990);
nor U23000 (N_23000,N_22023,N_22408);
nand U23001 (N_23001,N_22340,N_22143);
and U23002 (N_23002,N_22650,N_22256);
or U23003 (N_23003,N_22603,N_22560);
nor U23004 (N_23004,N_22027,N_22971);
and U23005 (N_23005,N_22025,N_22814);
or U23006 (N_23006,N_22329,N_22757);
and U23007 (N_23007,N_22267,N_22706);
nor U23008 (N_23008,N_22477,N_22754);
nor U23009 (N_23009,N_22456,N_22767);
nor U23010 (N_23010,N_22655,N_22834);
xor U23011 (N_23011,N_22326,N_22646);
xnor U23012 (N_23012,N_22682,N_22826);
nor U23013 (N_23013,N_22547,N_22186);
and U23014 (N_23014,N_22417,N_22697);
or U23015 (N_23015,N_22736,N_22428);
nand U23016 (N_23016,N_22606,N_22903);
and U23017 (N_23017,N_22298,N_22191);
nor U23018 (N_23018,N_22967,N_22555);
nor U23019 (N_23019,N_22483,N_22858);
xnor U23020 (N_23020,N_22578,N_22209);
xor U23021 (N_23021,N_22139,N_22470);
xor U23022 (N_23022,N_22899,N_22800);
and U23023 (N_23023,N_22149,N_22528);
or U23024 (N_23024,N_22792,N_22557);
and U23025 (N_23025,N_22914,N_22459);
and U23026 (N_23026,N_22839,N_22647);
nor U23027 (N_23027,N_22120,N_22553);
xor U23028 (N_23028,N_22011,N_22577);
nand U23029 (N_23029,N_22878,N_22857);
or U23030 (N_23030,N_22364,N_22531);
or U23031 (N_23031,N_22999,N_22929);
or U23032 (N_23032,N_22794,N_22702);
xnor U23033 (N_23033,N_22173,N_22179);
xor U23034 (N_23034,N_22146,N_22226);
or U23035 (N_23035,N_22112,N_22601);
nand U23036 (N_23036,N_22835,N_22550);
and U23037 (N_23037,N_22922,N_22439);
and U23038 (N_23038,N_22730,N_22221);
xnor U23039 (N_23039,N_22419,N_22368);
nand U23040 (N_23040,N_22691,N_22161);
xnor U23041 (N_23041,N_22561,N_22180);
nor U23042 (N_23042,N_22400,N_22463);
and U23043 (N_23043,N_22295,N_22866);
and U23044 (N_23044,N_22644,N_22401);
nand U23045 (N_23045,N_22748,N_22688);
nor U23046 (N_23046,N_22192,N_22067);
xor U23047 (N_23047,N_22225,N_22246);
xor U23048 (N_23048,N_22480,N_22404);
xnor U23049 (N_23049,N_22030,N_22896);
and U23050 (N_23050,N_22604,N_22167);
nor U23051 (N_23051,N_22862,N_22222);
and U23052 (N_23052,N_22559,N_22572);
nand U23053 (N_23053,N_22924,N_22598);
or U23054 (N_23054,N_22418,N_22659);
and U23055 (N_23055,N_22938,N_22307);
nand U23056 (N_23056,N_22345,N_22586);
and U23057 (N_23057,N_22770,N_22367);
nor U23058 (N_23058,N_22336,N_22305);
and U23059 (N_23059,N_22580,N_22460);
or U23060 (N_23060,N_22836,N_22570);
or U23061 (N_23061,N_22796,N_22930);
or U23062 (N_23062,N_22163,N_22510);
xnor U23063 (N_23063,N_22687,N_22521);
nand U23064 (N_23064,N_22845,N_22133);
xor U23065 (N_23065,N_22822,N_22735);
xor U23066 (N_23066,N_22506,N_22193);
nand U23067 (N_23067,N_22071,N_22979);
and U23068 (N_23068,N_22708,N_22332);
xor U23069 (N_23069,N_22338,N_22563);
nor U23070 (N_23070,N_22216,N_22339);
nor U23071 (N_23071,N_22158,N_22852);
nand U23072 (N_23072,N_22153,N_22512);
nor U23073 (N_23073,N_22874,N_22414);
and U23074 (N_23074,N_22271,N_22261);
nand U23075 (N_23075,N_22694,N_22156);
and U23076 (N_23076,N_22584,N_22362);
or U23077 (N_23077,N_22763,N_22849);
nand U23078 (N_23078,N_22063,N_22441);
xor U23079 (N_23079,N_22962,N_22094);
or U23080 (N_23080,N_22968,N_22692);
and U23081 (N_23081,N_22703,N_22619);
nor U23082 (N_23082,N_22473,N_22426);
nand U23083 (N_23083,N_22876,N_22709);
or U23084 (N_23084,N_22496,N_22765);
nor U23085 (N_23085,N_22723,N_22116);
and U23086 (N_23086,N_22396,N_22147);
xnor U23087 (N_23087,N_22928,N_22994);
and U23088 (N_23088,N_22840,N_22031);
nor U23089 (N_23089,N_22579,N_22233);
xor U23090 (N_23090,N_22085,N_22643);
nand U23091 (N_23091,N_22445,N_22091);
nand U23092 (N_23092,N_22049,N_22587);
or U23093 (N_23093,N_22070,N_22970);
xor U23094 (N_23094,N_22452,N_22328);
or U23095 (N_23095,N_22423,N_22170);
and U23096 (N_23096,N_22207,N_22466);
and U23097 (N_23097,N_22107,N_22389);
or U23098 (N_23098,N_22597,N_22178);
or U23099 (N_23099,N_22824,N_22039);
nand U23100 (N_23100,N_22168,N_22318);
xnor U23101 (N_23101,N_22213,N_22169);
and U23102 (N_23102,N_22361,N_22501);
xor U23103 (N_23103,N_22679,N_22782);
or U23104 (N_23104,N_22040,N_22020);
and U23105 (N_23105,N_22830,N_22160);
xor U23106 (N_23106,N_22548,N_22205);
or U23107 (N_23107,N_22371,N_22589);
nand U23108 (N_23108,N_22627,N_22095);
nand U23109 (N_23109,N_22821,N_22022);
nand U23110 (N_23110,N_22248,N_22253);
xnor U23111 (N_23111,N_22288,N_22969);
and U23112 (N_23112,N_22100,N_22433);
and U23113 (N_23113,N_22780,N_22720);
nor U23114 (N_23114,N_22744,N_22341);
or U23115 (N_23115,N_22282,N_22393);
and U23116 (N_23116,N_22327,N_22069);
nand U23117 (N_23117,N_22176,N_22135);
and U23118 (N_23118,N_22010,N_22721);
nand U23119 (N_23119,N_22718,N_22229);
and U23120 (N_23120,N_22319,N_22057);
and U23121 (N_23121,N_22019,N_22036);
xnor U23122 (N_23122,N_22403,N_22853);
nor U23123 (N_23123,N_22048,N_22901);
xnor U23124 (N_23124,N_22677,N_22435);
nand U23125 (N_23125,N_22942,N_22781);
and U23126 (N_23126,N_22861,N_22385);
and U23127 (N_23127,N_22908,N_22014);
or U23128 (N_23128,N_22114,N_22081);
nor U23129 (N_23129,N_22804,N_22947);
nor U23130 (N_23130,N_22130,N_22602);
nor U23131 (N_23131,N_22125,N_22753);
and U23132 (N_23132,N_22093,N_22725);
xor U23133 (N_23133,N_22497,N_22710);
xor U23134 (N_23134,N_22424,N_22645);
or U23135 (N_23135,N_22514,N_22458);
nor U23136 (N_23136,N_22972,N_22185);
or U23137 (N_23137,N_22883,N_22195);
nor U23138 (N_23138,N_22657,N_22281);
or U23139 (N_23139,N_22529,N_22372);
xor U23140 (N_23140,N_22806,N_22165);
nand U23141 (N_23141,N_22099,N_22076);
nand U23142 (N_23142,N_22653,N_22457);
or U23143 (N_23143,N_22632,N_22527);
nand U23144 (N_23144,N_22043,N_22363);
nor U23145 (N_23145,N_22787,N_22231);
xnor U23146 (N_23146,N_22144,N_22771);
nor U23147 (N_23147,N_22360,N_22008);
xnor U23148 (N_23148,N_22311,N_22427);
or U23149 (N_23149,N_22696,N_22541);
xnor U23150 (N_23150,N_22951,N_22569);
nand U23151 (N_23151,N_22097,N_22485);
or U23152 (N_23152,N_22838,N_22296);
and U23153 (N_23153,N_22775,N_22421);
nand U23154 (N_23154,N_22406,N_22912);
nor U23155 (N_23155,N_22953,N_22534);
or U23156 (N_23156,N_22941,N_22518);
nor U23157 (N_23157,N_22002,N_22592);
xnor U23158 (N_23158,N_22028,N_22998);
nor U23159 (N_23159,N_22240,N_22284);
xor U23160 (N_23160,N_22755,N_22618);
and U23161 (N_23161,N_22232,N_22910);
or U23162 (N_23162,N_22060,N_22954);
or U23163 (N_23163,N_22609,N_22795);
nand U23164 (N_23164,N_22275,N_22218);
nor U23165 (N_23165,N_22384,N_22825);
xnor U23166 (N_23166,N_22891,N_22162);
xnor U23167 (N_23167,N_22892,N_22286);
and U23168 (N_23168,N_22174,N_22481);
nor U23169 (N_23169,N_22032,N_22378);
and U23170 (N_23170,N_22668,N_22283);
or U23171 (N_23171,N_22773,N_22292);
and U23172 (N_23172,N_22948,N_22734);
xor U23173 (N_23173,N_22402,N_22933);
nand U23174 (N_23174,N_22551,N_22995);
and U23175 (N_23175,N_22515,N_22072);
nand U23176 (N_23176,N_22034,N_22376);
nor U23177 (N_23177,N_22488,N_22890);
nor U23178 (N_23178,N_22552,N_22467);
nand U23179 (N_23179,N_22616,N_22098);
and U23180 (N_23180,N_22390,N_22759);
nor U23181 (N_23181,N_22882,N_22513);
nand U23182 (N_23182,N_22184,N_22009);
and U23183 (N_23183,N_22793,N_22489);
or U23184 (N_23184,N_22898,N_22926);
and U23185 (N_23185,N_22410,N_22370);
and U23186 (N_23186,N_22096,N_22837);
nand U23187 (N_23187,N_22660,N_22206);
nand U23188 (N_23188,N_22591,N_22084);
and U23189 (N_23189,N_22394,N_22052);
nand U23190 (N_23190,N_22199,N_22608);
and U23191 (N_23191,N_22776,N_22752);
or U23192 (N_23192,N_22599,N_22260);
xor U23193 (N_23193,N_22511,N_22317);
nand U23194 (N_23194,N_22722,N_22092);
or U23195 (N_23195,N_22148,N_22202);
nand U23196 (N_23196,N_22425,N_22919);
xnor U23197 (N_23197,N_22409,N_22411);
nor U23198 (N_23198,N_22145,N_22904);
and U23199 (N_23199,N_22254,N_22651);
xnor U23200 (N_23200,N_22383,N_22422);
or U23201 (N_23201,N_22639,N_22065);
xnor U23202 (N_23202,N_22880,N_22662);
nor U23203 (N_23203,N_22881,N_22637);
nor U23204 (N_23204,N_22879,N_22301);
nor U23205 (N_23205,N_22415,N_22516);
nor U23206 (N_23206,N_22622,N_22211);
xnor U23207 (N_23207,N_22607,N_22965);
or U23208 (N_23208,N_22138,N_22519);
nor U23209 (N_23209,N_22568,N_22259);
nor U23210 (N_23210,N_22681,N_22988);
and U23211 (N_23211,N_22234,N_22728);
and U23212 (N_23212,N_22605,N_22869);
and U23213 (N_23213,N_22214,N_22851);
xor U23214 (N_23214,N_22333,N_22699);
xor U23215 (N_23215,N_22936,N_22877);
or U23216 (N_23216,N_22724,N_22287);
xnor U23217 (N_23217,N_22678,N_22508);
xnor U23218 (N_23218,N_22870,N_22129);
xor U23219 (N_23219,N_22064,N_22236);
xnor U23220 (N_23220,N_22935,N_22686);
or U23221 (N_23221,N_22056,N_22134);
nand U23222 (N_23222,N_22083,N_22676);
xnor U23223 (N_23223,N_22247,N_22986);
and U23224 (N_23224,N_22151,N_22102);
and U23225 (N_23225,N_22154,N_22983);
nor U23226 (N_23226,N_22255,N_22499);
xor U23227 (N_23227,N_22623,N_22732);
and U23228 (N_23228,N_22820,N_22429);
nor U23229 (N_23229,N_22007,N_22086);
and U23230 (N_23230,N_22331,N_22815);
nand U23231 (N_23231,N_22166,N_22630);
or U23232 (N_23232,N_22054,N_22062);
or U23233 (N_23233,N_22617,N_22119);
and U23234 (N_23234,N_22110,N_22871);
nand U23235 (N_23235,N_22888,N_22756);
nand U23236 (N_23236,N_22689,N_22540);
nand U23237 (N_23237,N_22729,N_22289);
and U23238 (N_23238,N_22377,N_22749);
nor U23239 (N_23239,N_22537,N_22194);
or U23240 (N_23240,N_22352,N_22012);
xor U23241 (N_23241,N_22320,N_22044);
nor U23242 (N_23242,N_22711,N_22073);
xnor U23243 (N_23243,N_22652,N_22810);
xor U23244 (N_23244,N_22268,N_22958);
xnor U23245 (N_23245,N_22693,N_22399);
or U23246 (N_23246,N_22374,N_22313);
nor U23247 (N_23247,N_22238,N_22157);
nand U23248 (N_23248,N_22128,N_22842);
xor U23249 (N_23249,N_22524,N_22981);
or U23250 (N_23250,N_22131,N_22306);
or U23251 (N_23251,N_22803,N_22545);
nor U23252 (N_23252,N_22172,N_22111);
xor U23253 (N_23253,N_22493,N_22159);
or U23254 (N_23254,N_22745,N_22931);
xor U23255 (N_23255,N_22454,N_22854);
or U23256 (N_23256,N_22113,N_22432);
nor U23257 (N_23257,N_22004,N_22818);
or U23258 (N_23258,N_22263,N_22142);
nor U23259 (N_23259,N_22035,N_22141);
or U23260 (N_23260,N_22127,N_22562);
nor U23261 (N_23261,N_22921,N_22358);
nor U23262 (N_23262,N_22766,N_22475);
xnor U23263 (N_23263,N_22886,N_22407);
nor U23264 (N_23264,N_22731,N_22916);
or U23265 (N_23265,N_22504,N_22611);
nand U23266 (N_23266,N_22164,N_22913);
xnor U23267 (N_23267,N_22900,N_22208);
nand U23268 (N_23268,N_22443,N_22526);
nand U23269 (N_23269,N_22554,N_22809);
nor U23270 (N_23270,N_22397,N_22576);
or U23271 (N_23271,N_22285,N_22638);
nor U23272 (N_23272,N_22380,N_22182);
nor U23273 (N_23273,N_22841,N_22798);
nor U23274 (N_23274,N_22906,N_22080);
nand U23275 (N_23275,N_22359,N_22717);
or U23276 (N_23276,N_22074,N_22183);
xor U23277 (N_23277,N_22405,N_22945);
nor U23278 (N_23278,N_22442,N_22447);
or U23279 (N_23279,N_22449,N_22391);
nor U23280 (N_23280,N_22784,N_22768);
nor U23281 (N_23281,N_22181,N_22859);
or U23282 (N_23282,N_22297,N_22046);
or U23283 (N_23283,N_22121,N_22889);
or U23284 (N_23284,N_22105,N_22117);
nor U23285 (N_23285,N_22024,N_22633);
or U23286 (N_23286,N_22189,N_22462);
or U23287 (N_23287,N_22530,N_22479);
nand U23288 (N_23288,N_22210,N_22799);
and U23289 (N_23289,N_22843,N_22266);
nor U23290 (N_23290,N_22103,N_22992);
xnor U23291 (N_23291,N_22029,N_22949);
xor U23292 (N_23292,N_22705,N_22438);
xor U23293 (N_23293,N_22520,N_22375);
nand U23294 (N_23294,N_22038,N_22716);
and U23295 (N_23295,N_22349,N_22507);
xnor U23296 (N_23296,N_22386,N_22982);
nand U23297 (N_23297,N_22590,N_22201);
nor U23298 (N_23298,N_22270,N_22430);
nand U23299 (N_23299,N_22783,N_22819);
and U23300 (N_23300,N_22543,N_22902);
nand U23301 (N_23301,N_22635,N_22525);
or U23302 (N_23302,N_22293,N_22269);
xnor U23303 (N_23303,N_22244,N_22667);
or U23304 (N_23304,N_22715,N_22943);
xnor U23305 (N_23305,N_22621,N_22087);
and U23306 (N_23306,N_22868,N_22614);
nand U23307 (N_23307,N_22549,N_22785);
nor U23308 (N_23308,N_22055,N_22321);
xnor U23309 (N_23309,N_22495,N_22015);
xor U23310 (N_23310,N_22956,N_22037);
xor U23311 (N_23311,N_22198,N_22137);
or U23312 (N_23312,N_22001,N_22847);
nor U23313 (N_23313,N_22991,N_22101);
nor U23314 (N_23314,N_22726,N_22050);
xor U23315 (N_23315,N_22684,N_22152);
xor U23316 (N_23316,N_22701,N_22434);
and U23317 (N_23317,N_22536,N_22873);
nand U23318 (N_23318,N_22769,N_22132);
nand U23319 (N_23319,N_22021,N_22813);
and U23320 (N_23320,N_22346,N_22583);
nand U23321 (N_23321,N_22713,N_22104);
xor U23322 (N_23322,N_22556,N_22350);
or U23323 (N_23323,N_22887,N_22140);
xor U23324 (N_23324,N_22649,N_22079);
and U23325 (N_23325,N_22600,N_22228);
nor U23326 (N_23326,N_22844,N_22567);
nand U23327 (N_23327,N_22227,N_22582);
xor U23328 (N_23328,N_22016,N_22685);
nand U23329 (N_23329,N_22628,N_22864);
and U23330 (N_23330,N_22944,N_22314);
or U23331 (N_23331,N_22907,N_22648);
xnor U23332 (N_23332,N_22344,N_22656);
and U23333 (N_23333,N_22950,N_22805);
nand U23334 (N_23334,N_22276,N_22666);
and U23335 (N_23335,N_22575,N_22751);
and U23336 (N_23336,N_22077,N_22190);
nor U23337 (N_23337,N_22237,N_22779);
and U23338 (N_23338,N_22934,N_22239);
xor U23339 (N_23339,N_22373,N_22278);
and U23340 (N_23340,N_22817,N_22932);
nor U23341 (N_23341,N_22355,N_22764);
or U23342 (N_23342,N_22505,N_22875);
nand U23343 (N_23343,N_22727,N_22279);
xor U23344 (N_23344,N_22961,N_22829);
nand U23345 (N_23345,N_22446,N_22823);
or U23346 (N_23346,N_22960,N_22867);
nor U23347 (N_23347,N_22658,N_22343);
nor U23348 (N_23348,N_22303,N_22465);
nor U23349 (N_23349,N_22224,N_22624);
or U23350 (N_23350,N_22946,N_22017);
nand U23351 (N_23351,N_22005,N_22000);
nor U23352 (N_23352,N_22532,N_22641);
and U23353 (N_23353,N_22833,N_22626);
nand U23354 (N_23354,N_22444,N_22850);
xor U23355 (N_23355,N_22539,N_22801);
and U23356 (N_23356,N_22420,N_22090);
or U23357 (N_23357,N_22760,N_22546);
and U23358 (N_23358,N_22917,N_22468);
and U23359 (N_23359,N_22330,N_22106);
nor U23360 (N_23360,N_22342,N_22574);
xnor U23361 (N_23361,N_22976,N_22354);
or U23362 (N_23362,N_22348,N_22300);
xor U23363 (N_23363,N_22894,N_22963);
and U23364 (N_23364,N_22089,N_22761);
nor U23365 (N_23365,N_22985,N_22750);
or U23366 (N_23366,N_22033,N_22461);
nor U23367 (N_23367,N_22381,N_22957);
xor U23368 (N_23368,N_22778,N_22669);
nand U23369 (N_23369,N_22013,N_22788);
nand U23370 (N_23370,N_22041,N_22250);
nor U23371 (N_23371,N_22920,N_22905);
or U23372 (N_23372,N_22966,N_22634);
or U23373 (N_23373,N_22440,N_22264);
xor U23374 (N_23374,N_22596,N_22828);
nor U23375 (N_23375,N_22392,N_22413);
xnor U23376 (N_23376,N_22451,N_22595);
and U23377 (N_23377,N_22797,N_22290);
or U23378 (N_23378,N_22334,N_22455);
or U23379 (N_23379,N_22118,N_22996);
nor U23380 (N_23380,N_22993,N_22789);
nor U23381 (N_23381,N_22664,N_22807);
and U23382 (N_23382,N_22500,N_22827);
nor U23383 (N_23383,N_22066,N_22498);
nor U23384 (N_23384,N_22448,N_22472);
and U23385 (N_23385,N_22059,N_22078);
xnor U23386 (N_23386,N_22631,N_22245);
nand U23387 (N_23387,N_22661,N_22122);
nor U23388 (N_23388,N_22310,N_22704);
nand U23389 (N_23389,N_22517,N_22989);
and U23390 (N_23390,N_22431,N_22047);
nand U23391 (N_23391,N_22739,N_22816);
xnor U23392 (N_23392,N_22223,N_22042);
and U23393 (N_23393,N_22812,N_22774);
or U23394 (N_23394,N_22923,N_22885);
xor U23395 (N_23395,N_22476,N_22758);
nor U23396 (N_23396,N_22337,N_22200);
nand U23397 (N_23397,N_22594,N_22610);
or U23398 (N_23398,N_22915,N_22719);
nand U23399 (N_23399,N_22625,N_22535);
or U23400 (N_23400,N_22277,N_22503);
and U23401 (N_23401,N_22573,N_22353);
xor U23402 (N_23402,N_22509,N_22808);
and U23403 (N_23403,N_22243,N_22058);
nor U23404 (N_23404,N_22698,N_22217);
nand U23405 (N_23405,N_22856,N_22252);
and U23406 (N_23406,N_22395,N_22683);
nor U23407 (N_23407,N_22642,N_22502);
and U23408 (N_23408,N_22474,N_22884);
nor U23409 (N_23409,N_22109,N_22155);
xor U23410 (N_23410,N_22990,N_22241);
nand U23411 (N_23411,N_22357,N_22469);
or U23412 (N_23412,N_22257,N_22762);
nand U23413 (N_23413,N_22280,N_22964);
xor U23414 (N_23414,N_22309,N_22663);
or U23415 (N_23415,N_22335,N_22187);
nor U23416 (N_23416,N_22737,N_22203);
and U23417 (N_23417,N_22219,N_22262);
or U23418 (N_23418,N_22484,N_22542);
nor U23419 (N_23419,N_22196,N_22487);
and U23420 (N_23420,N_22249,N_22068);
nor U23421 (N_23421,N_22136,N_22860);
or U23422 (N_23422,N_22984,N_22108);
nand U23423 (N_23423,N_22675,N_22802);
nor U23424 (N_23424,N_22347,N_22061);
and U23425 (N_23425,N_22436,N_22671);
or U23426 (N_23426,N_22003,N_22733);
xnor U23427 (N_23427,N_22695,N_22053);
xor U23428 (N_23428,N_22482,N_22453);
or U23429 (N_23429,N_22450,N_22558);
nand U23430 (N_23430,N_22620,N_22365);
nand U23431 (N_23431,N_22872,N_22315);
xor U23432 (N_23432,N_22416,N_22670);
and U23433 (N_23433,N_22251,N_22322);
and U23434 (N_23434,N_22743,N_22124);
xor U23435 (N_23435,N_22323,N_22690);
or U23436 (N_23436,N_22777,N_22351);
and U23437 (N_23437,N_22294,N_22564);
or U23438 (N_23438,N_22673,N_22379);
nor U23439 (N_23439,N_22265,N_22665);
nor U23440 (N_23440,N_22940,N_22171);
and U23441 (N_23441,N_22123,N_22486);
and U23442 (N_23442,N_22846,N_22491);
nand U23443 (N_23443,N_22316,N_22088);
or U23444 (N_23444,N_22366,N_22654);
xor U23445 (N_23445,N_22565,N_22045);
or U23446 (N_23446,N_22707,N_22175);
xnor U23447 (N_23447,N_22273,N_22700);
and U23448 (N_23448,N_22291,N_22018);
nand U23449 (N_23449,N_22714,N_22955);
xnor U23450 (N_23450,N_22790,N_22082);
xnor U23451 (N_23451,N_22494,N_22230);
or U23452 (N_23452,N_22272,N_22831);
nor U23453 (N_23453,N_22593,N_22911);
nand U23454 (N_23454,N_22308,N_22324);
nor U23455 (N_23455,N_22412,N_22974);
nor U23456 (N_23456,N_22987,N_22612);
nand U23457 (N_23457,N_22978,N_22588);
nand U23458 (N_23458,N_22026,N_22977);
nor U23459 (N_23459,N_22464,N_22613);
nor U23460 (N_23460,N_22126,N_22188);
xor U23461 (N_23461,N_22636,N_22672);
xor U23462 (N_23462,N_22522,N_22544);
or U23463 (N_23463,N_22242,N_22772);
nand U23464 (N_23464,N_22523,N_22571);
xor U23465 (N_23465,N_22235,N_22738);
nand U23466 (N_23466,N_22712,N_22492);
or U23467 (N_23467,N_22855,N_22674);
nand U23468 (N_23468,N_22791,N_22478);
nor U23469 (N_23469,N_22897,N_22746);
nor U23470 (N_23470,N_22927,N_22177);
xor U23471 (N_23471,N_22212,N_22051);
nand U23472 (N_23472,N_22369,N_22197);
and U23473 (N_23473,N_22388,N_22848);
nand U23474 (N_23474,N_22865,N_22382);
xnor U23475 (N_23475,N_22959,N_22680);
nand U23476 (N_23476,N_22615,N_22863);
and U23477 (N_23477,N_22585,N_22918);
and U23478 (N_23478,N_22538,N_22811);
nand U23479 (N_23479,N_22302,N_22937);
nand U23480 (N_23480,N_22566,N_22925);
nand U23481 (N_23481,N_22832,N_22997);
and U23482 (N_23482,N_22356,N_22893);
nor U23483 (N_23483,N_22312,N_22490);
nand U23484 (N_23484,N_22398,N_22973);
nor U23485 (N_23485,N_22741,N_22115);
nor U23486 (N_23486,N_22640,N_22215);
or U23487 (N_23487,N_22075,N_22980);
nand U23488 (N_23488,N_22006,N_22975);
nor U23489 (N_23489,N_22325,N_22629);
nand U23490 (N_23490,N_22471,N_22939);
nor U23491 (N_23491,N_22895,N_22740);
or U23492 (N_23492,N_22204,N_22304);
nor U23493 (N_23493,N_22387,N_22258);
nor U23494 (N_23494,N_22220,N_22274);
nor U23495 (N_23495,N_22150,N_22742);
or U23496 (N_23496,N_22437,N_22299);
nor U23497 (N_23497,N_22581,N_22909);
nor U23498 (N_23498,N_22747,N_22786);
or U23499 (N_23499,N_22533,N_22952);
nand U23500 (N_23500,N_22459,N_22763);
nor U23501 (N_23501,N_22957,N_22651);
nor U23502 (N_23502,N_22527,N_22100);
xor U23503 (N_23503,N_22397,N_22943);
nand U23504 (N_23504,N_22652,N_22534);
nor U23505 (N_23505,N_22385,N_22638);
nand U23506 (N_23506,N_22946,N_22316);
nand U23507 (N_23507,N_22672,N_22995);
xnor U23508 (N_23508,N_22880,N_22916);
or U23509 (N_23509,N_22577,N_22509);
xor U23510 (N_23510,N_22725,N_22251);
nor U23511 (N_23511,N_22245,N_22416);
and U23512 (N_23512,N_22791,N_22168);
and U23513 (N_23513,N_22590,N_22263);
and U23514 (N_23514,N_22670,N_22576);
nor U23515 (N_23515,N_22020,N_22300);
or U23516 (N_23516,N_22459,N_22129);
nand U23517 (N_23517,N_22473,N_22406);
or U23518 (N_23518,N_22683,N_22996);
or U23519 (N_23519,N_22358,N_22041);
and U23520 (N_23520,N_22965,N_22145);
and U23521 (N_23521,N_22123,N_22144);
nand U23522 (N_23522,N_22467,N_22426);
or U23523 (N_23523,N_22839,N_22736);
and U23524 (N_23524,N_22840,N_22939);
xor U23525 (N_23525,N_22311,N_22401);
nand U23526 (N_23526,N_22007,N_22974);
and U23527 (N_23527,N_22363,N_22437);
and U23528 (N_23528,N_22820,N_22258);
nor U23529 (N_23529,N_22389,N_22651);
nor U23530 (N_23530,N_22445,N_22318);
nor U23531 (N_23531,N_22796,N_22439);
nand U23532 (N_23532,N_22481,N_22024);
nand U23533 (N_23533,N_22820,N_22347);
or U23534 (N_23534,N_22761,N_22781);
xor U23535 (N_23535,N_22668,N_22046);
or U23536 (N_23536,N_22424,N_22613);
and U23537 (N_23537,N_22839,N_22955);
nor U23538 (N_23538,N_22919,N_22029);
nor U23539 (N_23539,N_22204,N_22070);
xor U23540 (N_23540,N_22796,N_22980);
and U23541 (N_23541,N_22982,N_22306);
and U23542 (N_23542,N_22808,N_22632);
or U23543 (N_23543,N_22903,N_22997);
and U23544 (N_23544,N_22863,N_22072);
nor U23545 (N_23545,N_22220,N_22320);
or U23546 (N_23546,N_22910,N_22896);
nand U23547 (N_23547,N_22748,N_22874);
nand U23548 (N_23548,N_22522,N_22683);
and U23549 (N_23549,N_22459,N_22430);
and U23550 (N_23550,N_22265,N_22588);
or U23551 (N_23551,N_22846,N_22713);
or U23552 (N_23552,N_22735,N_22464);
and U23553 (N_23553,N_22860,N_22538);
and U23554 (N_23554,N_22537,N_22462);
xnor U23555 (N_23555,N_22042,N_22316);
xor U23556 (N_23556,N_22572,N_22577);
nand U23557 (N_23557,N_22248,N_22577);
nand U23558 (N_23558,N_22189,N_22635);
nor U23559 (N_23559,N_22110,N_22994);
xor U23560 (N_23560,N_22538,N_22692);
nand U23561 (N_23561,N_22900,N_22409);
nor U23562 (N_23562,N_22749,N_22145);
xnor U23563 (N_23563,N_22339,N_22347);
and U23564 (N_23564,N_22896,N_22364);
nor U23565 (N_23565,N_22321,N_22997);
and U23566 (N_23566,N_22551,N_22644);
or U23567 (N_23567,N_22530,N_22831);
or U23568 (N_23568,N_22370,N_22124);
or U23569 (N_23569,N_22551,N_22788);
nand U23570 (N_23570,N_22145,N_22861);
and U23571 (N_23571,N_22267,N_22412);
or U23572 (N_23572,N_22507,N_22177);
nand U23573 (N_23573,N_22682,N_22770);
or U23574 (N_23574,N_22043,N_22978);
nor U23575 (N_23575,N_22472,N_22267);
or U23576 (N_23576,N_22160,N_22812);
xor U23577 (N_23577,N_22657,N_22502);
nor U23578 (N_23578,N_22840,N_22932);
xor U23579 (N_23579,N_22430,N_22558);
and U23580 (N_23580,N_22811,N_22762);
nand U23581 (N_23581,N_22035,N_22301);
nand U23582 (N_23582,N_22458,N_22709);
nand U23583 (N_23583,N_22209,N_22754);
and U23584 (N_23584,N_22999,N_22894);
nor U23585 (N_23585,N_22723,N_22304);
nand U23586 (N_23586,N_22068,N_22864);
and U23587 (N_23587,N_22359,N_22586);
and U23588 (N_23588,N_22702,N_22919);
or U23589 (N_23589,N_22880,N_22644);
or U23590 (N_23590,N_22913,N_22521);
nor U23591 (N_23591,N_22750,N_22417);
xnor U23592 (N_23592,N_22925,N_22647);
nand U23593 (N_23593,N_22294,N_22830);
or U23594 (N_23594,N_22979,N_22752);
nand U23595 (N_23595,N_22366,N_22800);
nor U23596 (N_23596,N_22268,N_22819);
nor U23597 (N_23597,N_22836,N_22926);
xor U23598 (N_23598,N_22444,N_22692);
nor U23599 (N_23599,N_22298,N_22579);
or U23600 (N_23600,N_22771,N_22320);
nor U23601 (N_23601,N_22381,N_22567);
or U23602 (N_23602,N_22931,N_22506);
nor U23603 (N_23603,N_22529,N_22896);
nor U23604 (N_23604,N_22636,N_22664);
and U23605 (N_23605,N_22667,N_22105);
and U23606 (N_23606,N_22979,N_22850);
or U23607 (N_23607,N_22973,N_22687);
or U23608 (N_23608,N_22725,N_22135);
and U23609 (N_23609,N_22360,N_22561);
and U23610 (N_23610,N_22469,N_22687);
and U23611 (N_23611,N_22455,N_22975);
nor U23612 (N_23612,N_22853,N_22758);
nand U23613 (N_23613,N_22770,N_22086);
nor U23614 (N_23614,N_22720,N_22705);
or U23615 (N_23615,N_22717,N_22512);
nand U23616 (N_23616,N_22233,N_22414);
xnor U23617 (N_23617,N_22917,N_22101);
nor U23618 (N_23618,N_22135,N_22551);
nand U23619 (N_23619,N_22727,N_22988);
and U23620 (N_23620,N_22528,N_22094);
or U23621 (N_23621,N_22205,N_22249);
nor U23622 (N_23622,N_22748,N_22137);
and U23623 (N_23623,N_22225,N_22881);
nor U23624 (N_23624,N_22707,N_22281);
xor U23625 (N_23625,N_22803,N_22705);
xnor U23626 (N_23626,N_22751,N_22509);
nand U23627 (N_23627,N_22789,N_22159);
or U23628 (N_23628,N_22670,N_22138);
nor U23629 (N_23629,N_22869,N_22514);
nand U23630 (N_23630,N_22274,N_22015);
nand U23631 (N_23631,N_22032,N_22545);
or U23632 (N_23632,N_22201,N_22402);
and U23633 (N_23633,N_22710,N_22069);
xor U23634 (N_23634,N_22557,N_22380);
nand U23635 (N_23635,N_22282,N_22227);
nand U23636 (N_23636,N_22406,N_22606);
or U23637 (N_23637,N_22847,N_22667);
nand U23638 (N_23638,N_22474,N_22014);
nand U23639 (N_23639,N_22495,N_22081);
nand U23640 (N_23640,N_22152,N_22803);
nor U23641 (N_23641,N_22625,N_22123);
nor U23642 (N_23642,N_22792,N_22219);
nor U23643 (N_23643,N_22924,N_22788);
or U23644 (N_23644,N_22748,N_22539);
or U23645 (N_23645,N_22479,N_22422);
nor U23646 (N_23646,N_22039,N_22674);
and U23647 (N_23647,N_22813,N_22497);
xnor U23648 (N_23648,N_22797,N_22455);
xor U23649 (N_23649,N_22785,N_22993);
xor U23650 (N_23650,N_22077,N_22964);
xnor U23651 (N_23651,N_22679,N_22093);
xor U23652 (N_23652,N_22624,N_22264);
nand U23653 (N_23653,N_22264,N_22724);
xnor U23654 (N_23654,N_22618,N_22151);
nand U23655 (N_23655,N_22558,N_22343);
nand U23656 (N_23656,N_22357,N_22573);
nor U23657 (N_23657,N_22201,N_22480);
xor U23658 (N_23658,N_22528,N_22107);
xor U23659 (N_23659,N_22541,N_22892);
or U23660 (N_23660,N_22481,N_22042);
nand U23661 (N_23661,N_22089,N_22229);
or U23662 (N_23662,N_22873,N_22360);
and U23663 (N_23663,N_22357,N_22840);
nor U23664 (N_23664,N_22497,N_22430);
or U23665 (N_23665,N_22683,N_22114);
xnor U23666 (N_23666,N_22795,N_22559);
xor U23667 (N_23667,N_22252,N_22240);
and U23668 (N_23668,N_22430,N_22166);
nand U23669 (N_23669,N_22957,N_22785);
xor U23670 (N_23670,N_22266,N_22097);
or U23671 (N_23671,N_22987,N_22647);
or U23672 (N_23672,N_22354,N_22483);
and U23673 (N_23673,N_22756,N_22735);
or U23674 (N_23674,N_22738,N_22519);
and U23675 (N_23675,N_22329,N_22377);
nand U23676 (N_23676,N_22791,N_22140);
nor U23677 (N_23677,N_22167,N_22860);
nor U23678 (N_23678,N_22415,N_22635);
xor U23679 (N_23679,N_22804,N_22667);
nand U23680 (N_23680,N_22016,N_22748);
xnor U23681 (N_23681,N_22573,N_22254);
nand U23682 (N_23682,N_22783,N_22807);
nand U23683 (N_23683,N_22769,N_22939);
nor U23684 (N_23684,N_22545,N_22060);
nor U23685 (N_23685,N_22823,N_22657);
and U23686 (N_23686,N_22922,N_22248);
xor U23687 (N_23687,N_22634,N_22248);
and U23688 (N_23688,N_22509,N_22071);
and U23689 (N_23689,N_22556,N_22056);
or U23690 (N_23690,N_22936,N_22730);
xor U23691 (N_23691,N_22211,N_22278);
and U23692 (N_23692,N_22797,N_22583);
or U23693 (N_23693,N_22393,N_22880);
nor U23694 (N_23694,N_22799,N_22207);
nor U23695 (N_23695,N_22269,N_22403);
xor U23696 (N_23696,N_22048,N_22026);
nor U23697 (N_23697,N_22551,N_22182);
xnor U23698 (N_23698,N_22471,N_22565);
or U23699 (N_23699,N_22006,N_22426);
nor U23700 (N_23700,N_22187,N_22243);
nor U23701 (N_23701,N_22967,N_22216);
or U23702 (N_23702,N_22536,N_22898);
and U23703 (N_23703,N_22341,N_22794);
nand U23704 (N_23704,N_22239,N_22381);
or U23705 (N_23705,N_22276,N_22189);
and U23706 (N_23706,N_22332,N_22366);
and U23707 (N_23707,N_22974,N_22797);
xnor U23708 (N_23708,N_22147,N_22287);
nor U23709 (N_23709,N_22570,N_22526);
and U23710 (N_23710,N_22618,N_22602);
or U23711 (N_23711,N_22832,N_22730);
or U23712 (N_23712,N_22345,N_22392);
nand U23713 (N_23713,N_22784,N_22278);
and U23714 (N_23714,N_22169,N_22921);
or U23715 (N_23715,N_22753,N_22628);
nand U23716 (N_23716,N_22281,N_22922);
or U23717 (N_23717,N_22360,N_22186);
nor U23718 (N_23718,N_22537,N_22214);
nand U23719 (N_23719,N_22381,N_22102);
nor U23720 (N_23720,N_22113,N_22490);
xnor U23721 (N_23721,N_22514,N_22748);
and U23722 (N_23722,N_22423,N_22562);
nor U23723 (N_23723,N_22407,N_22439);
or U23724 (N_23724,N_22218,N_22842);
or U23725 (N_23725,N_22317,N_22831);
nand U23726 (N_23726,N_22915,N_22224);
nand U23727 (N_23727,N_22402,N_22560);
xor U23728 (N_23728,N_22058,N_22547);
nor U23729 (N_23729,N_22357,N_22158);
xnor U23730 (N_23730,N_22639,N_22832);
xor U23731 (N_23731,N_22890,N_22318);
nand U23732 (N_23732,N_22882,N_22846);
and U23733 (N_23733,N_22047,N_22698);
nor U23734 (N_23734,N_22832,N_22235);
and U23735 (N_23735,N_22901,N_22236);
or U23736 (N_23736,N_22703,N_22103);
xnor U23737 (N_23737,N_22932,N_22108);
and U23738 (N_23738,N_22518,N_22053);
nand U23739 (N_23739,N_22293,N_22900);
nand U23740 (N_23740,N_22883,N_22707);
nor U23741 (N_23741,N_22693,N_22079);
nor U23742 (N_23742,N_22878,N_22017);
nand U23743 (N_23743,N_22841,N_22777);
xnor U23744 (N_23744,N_22340,N_22297);
and U23745 (N_23745,N_22185,N_22683);
and U23746 (N_23746,N_22172,N_22259);
nor U23747 (N_23747,N_22764,N_22806);
nor U23748 (N_23748,N_22209,N_22832);
nor U23749 (N_23749,N_22854,N_22736);
nand U23750 (N_23750,N_22812,N_22026);
or U23751 (N_23751,N_22449,N_22533);
nand U23752 (N_23752,N_22976,N_22446);
nand U23753 (N_23753,N_22488,N_22471);
and U23754 (N_23754,N_22053,N_22531);
nor U23755 (N_23755,N_22894,N_22822);
nand U23756 (N_23756,N_22252,N_22595);
nand U23757 (N_23757,N_22981,N_22925);
or U23758 (N_23758,N_22175,N_22264);
or U23759 (N_23759,N_22494,N_22796);
nand U23760 (N_23760,N_22990,N_22102);
xor U23761 (N_23761,N_22666,N_22884);
and U23762 (N_23762,N_22239,N_22251);
xnor U23763 (N_23763,N_22623,N_22823);
or U23764 (N_23764,N_22014,N_22755);
and U23765 (N_23765,N_22452,N_22016);
or U23766 (N_23766,N_22743,N_22530);
xor U23767 (N_23767,N_22545,N_22750);
xnor U23768 (N_23768,N_22896,N_22454);
xnor U23769 (N_23769,N_22499,N_22850);
xnor U23770 (N_23770,N_22106,N_22617);
xor U23771 (N_23771,N_22032,N_22494);
and U23772 (N_23772,N_22733,N_22701);
or U23773 (N_23773,N_22058,N_22505);
or U23774 (N_23774,N_22026,N_22509);
and U23775 (N_23775,N_22388,N_22405);
xnor U23776 (N_23776,N_22397,N_22552);
nor U23777 (N_23777,N_22875,N_22694);
xnor U23778 (N_23778,N_22005,N_22169);
or U23779 (N_23779,N_22544,N_22481);
or U23780 (N_23780,N_22634,N_22616);
nand U23781 (N_23781,N_22277,N_22325);
nor U23782 (N_23782,N_22565,N_22001);
nor U23783 (N_23783,N_22766,N_22850);
nor U23784 (N_23784,N_22388,N_22211);
and U23785 (N_23785,N_22947,N_22089);
or U23786 (N_23786,N_22870,N_22639);
nand U23787 (N_23787,N_22444,N_22521);
nand U23788 (N_23788,N_22130,N_22278);
nand U23789 (N_23789,N_22658,N_22462);
or U23790 (N_23790,N_22592,N_22273);
xnor U23791 (N_23791,N_22926,N_22478);
and U23792 (N_23792,N_22503,N_22312);
nor U23793 (N_23793,N_22968,N_22884);
nand U23794 (N_23794,N_22534,N_22751);
nand U23795 (N_23795,N_22746,N_22714);
nand U23796 (N_23796,N_22555,N_22773);
and U23797 (N_23797,N_22786,N_22907);
nand U23798 (N_23798,N_22250,N_22771);
xor U23799 (N_23799,N_22296,N_22376);
xor U23800 (N_23800,N_22931,N_22360);
nand U23801 (N_23801,N_22080,N_22913);
or U23802 (N_23802,N_22878,N_22941);
and U23803 (N_23803,N_22113,N_22579);
nand U23804 (N_23804,N_22199,N_22770);
or U23805 (N_23805,N_22932,N_22763);
or U23806 (N_23806,N_22137,N_22927);
or U23807 (N_23807,N_22033,N_22933);
xnor U23808 (N_23808,N_22609,N_22800);
nand U23809 (N_23809,N_22900,N_22713);
xnor U23810 (N_23810,N_22575,N_22400);
xor U23811 (N_23811,N_22655,N_22432);
and U23812 (N_23812,N_22668,N_22885);
and U23813 (N_23813,N_22117,N_22606);
and U23814 (N_23814,N_22387,N_22400);
xor U23815 (N_23815,N_22396,N_22383);
nand U23816 (N_23816,N_22704,N_22862);
nor U23817 (N_23817,N_22473,N_22348);
nor U23818 (N_23818,N_22919,N_22868);
xor U23819 (N_23819,N_22097,N_22935);
nand U23820 (N_23820,N_22674,N_22709);
nand U23821 (N_23821,N_22713,N_22621);
and U23822 (N_23822,N_22203,N_22287);
nand U23823 (N_23823,N_22078,N_22254);
xor U23824 (N_23824,N_22771,N_22204);
nor U23825 (N_23825,N_22419,N_22268);
xnor U23826 (N_23826,N_22425,N_22960);
and U23827 (N_23827,N_22311,N_22329);
and U23828 (N_23828,N_22100,N_22007);
and U23829 (N_23829,N_22036,N_22180);
xnor U23830 (N_23830,N_22626,N_22105);
and U23831 (N_23831,N_22879,N_22923);
or U23832 (N_23832,N_22860,N_22601);
nand U23833 (N_23833,N_22334,N_22336);
or U23834 (N_23834,N_22279,N_22340);
or U23835 (N_23835,N_22451,N_22327);
xnor U23836 (N_23836,N_22742,N_22698);
nor U23837 (N_23837,N_22485,N_22107);
nor U23838 (N_23838,N_22369,N_22263);
nor U23839 (N_23839,N_22800,N_22383);
nand U23840 (N_23840,N_22019,N_22552);
xor U23841 (N_23841,N_22633,N_22897);
or U23842 (N_23842,N_22722,N_22138);
nor U23843 (N_23843,N_22485,N_22930);
nor U23844 (N_23844,N_22709,N_22657);
and U23845 (N_23845,N_22458,N_22188);
nand U23846 (N_23846,N_22839,N_22638);
nor U23847 (N_23847,N_22365,N_22276);
and U23848 (N_23848,N_22424,N_22854);
or U23849 (N_23849,N_22982,N_22717);
or U23850 (N_23850,N_22935,N_22841);
xnor U23851 (N_23851,N_22581,N_22763);
xnor U23852 (N_23852,N_22776,N_22890);
or U23853 (N_23853,N_22116,N_22083);
or U23854 (N_23854,N_22430,N_22196);
and U23855 (N_23855,N_22983,N_22792);
nand U23856 (N_23856,N_22407,N_22046);
xnor U23857 (N_23857,N_22557,N_22948);
xnor U23858 (N_23858,N_22157,N_22328);
and U23859 (N_23859,N_22256,N_22829);
and U23860 (N_23860,N_22303,N_22699);
nand U23861 (N_23861,N_22748,N_22793);
nor U23862 (N_23862,N_22111,N_22189);
xor U23863 (N_23863,N_22714,N_22601);
xor U23864 (N_23864,N_22096,N_22901);
xor U23865 (N_23865,N_22533,N_22809);
xnor U23866 (N_23866,N_22184,N_22286);
or U23867 (N_23867,N_22978,N_22241);
or U23868 (N_23868,N_22681,N_22924);
xnor U23869 (N_23869,N_22436,N_22642);
xnor U23870 (N_23870,N_22234,N_22313);
nand U23871 (N_23871,N_22035,N_22041);
or U23872 (N_23872,N_22271,N_22092);
and U23873 (N_23873,N_22744,N_22880);
and U23874 (N_23874,N_22875,N_22842);
or U23875 (N_23875,N_22299,N_22245);
nor U23876 (N_23876,N_22602,N_22616);
nand U23877 (N_23877,N_22824,N_22863);
nor U23878 (N_23878,N_22690,N_22227);
nor U23879 (N_23879,N_22044,N_22689);
nand U23880 (N_23880,N_22718,N_22967);
xor U23881 (N_23881,N_22287,N_22180);
nor U23882 (N_23882,N_22267,N_22771);
xor U23883 (N_23883,N_22060,N_22126);
nor U23884 (N_23884,N_22273,N_22544);
nor U23885 (N_23885,N_22171,N_22908);
or U23886 (N_23886,N_22596,N_22357);
or U23887 (N_23887,N_22453,N_22486);
nand U23888 (N_23888,N_22101,N_22236);
or U23889 (N_23889,N_22597,N_22485);
nor U23890 (N_23890,N_22566,N_22038);
and U23891 (N_23891,N_22645,N_22721);
xnor U23892 (N_23892,N_22956,N_22475);
or U23893 (N_23893,N_22653,N_22223);
and U23894 (N_23894,N_22675,N_22390);
and U23895 (N_23895,N_22162,N_22704);
nor U23896 (N_23896,N_22585,N_22643);
nand U23897 (N_23897,N_22164,N_22440);
and U23898 (N_23898,N_22811,N_22334);
nand U23899 (N_23899,N_22738,N_22305);
and U23900 (N_23900,N_22628,N_22030);
xnor U23901 (N_23901,N_22250,N_22756);
nor U23902 (N_23902,N_22660,N_22305);
nand U23903 (N_23903,N_22191,N_22272);
nand U23904 (N_23904,N_22895,N_22163);
nor U23905 (N_23905,N_22554,N_22224);
and U23906 (N_23906,N_22533,N_22913);
or U23907 (N_23907,N_22186,N_22893);
nand U23908 (N_23908,N_22738,N_22505);
nor U23909 (N_23909,N_22855,N_22305);
or U23910 (N_23910,N_22383,N_22510);
and U23911 (N_23911,N_22844,N_22525);
xor U23912 (N_23912,N_22791,N_22136);
nand U23913 (N_23913,N_22587,N_22654);
and U23914 (N_23914,N_22290,N_22528);
nand U23915 (N_23915,N_22321,N_22667);
nand U23916 (N_23916,N_22587,N_22383);
nand U23917 (N_23917,N_22627,N_22398);
and U23918 (N_23918,N_22008,N_22843);
or U23919 (N_23919,N_22805,N_22669);
and U23920 (N_23920,N_22343,N_22526);
and U23921 (N_23921,N_22180,N_22541);
and U23922 (N_23922,N_22137,N_22997);
and U23923 (N_23923,N_22854,N_22991);
xnor U23924 (N_23924,N_22847,N_22275);
or U23925 (N_23925,N_22213,N_22469);
nand U23926 (N_23926,N_22333,N_22621);
nand U23927 (N_23927,N_22552,N_22437);
or U23928 (N_23928,N_22037,N_22493);
xnor U23929 (N_23929,N_22627,N_22676);
nor U23930 (N_23930,N_22213,N_22700);
nor U23931 (N_23931,N_22300,N_22240);
nor U23932 (N_23932,N_22328,N_22834);
or U23933 (N_23933,N_22103,N_22295);
xnor U23934 (N_23934,N_22862,N_22229);
xor U23935 (N_23935,N_22451,N_22817);
xnor U23936 (N_23936,N_22478,N_22579);
nand U23937 (N_23937,N_22790,N_22992);
xor U23938 (N_23938,N_22566,N_22030);
or U23939 (N_23939,N_22207,N_22983);
xnor U23940 (N_23940,N_22895,N_22734);
nand U23941 (N_23941,N_22169,N_22075);
or U23942 (N_23942,N_22948,N_22387);
nor U23943 (N_23943,N_22066,N_22137);
and U23944 (N_23944,N_22059,N_22785);
nand U23945 (N_23945,N_22005,N_22520);
or U23946 (N_23946,N_22314,N_22067);
or U23947 (N_23947,N_22588,N_22508);
xor U23948 (N_23948,N_22331,N_22507);
nor U23949 (N_23949,N_22734,N_22779);
nand U23950 (N_23950,N_22031,N_22872);
nor U23951 (N_23951,N_22424,N_22003);
nand U23952 (N_23952,N_22548,N_22644);
xor U23953 (N_23953,N_22785,N_22130);
or U23954 (N_23954,N_22461,N_22801);
xor U23955 (N_23955,N_22158,N_22570);
and U23956 (N_23956,N_22049,N_22179);
xor U23957 (N_23957,N_22927,N_22116);
xnor U23958 (N_23958,N_22982,N_22403);
and U23959 (N_23959,N_22378,N_22727);
xnor U23960 (N_23960,N_22692,N_22661);
nor U23961 (N_23961,N_22269,N_22901);
or U23962 (N_23962,N_22739,N_22975);
nor U23963 (N_23963,N_22457,N_22129);
and U23964 (N_23964,N_22304,N_22951);
nand U23965 (N_23965,N_22265,N_22436);
xor U23966 (N_23966,N_22012,N_22626);
or U23967 (N_23967,N_22055,N_22501);
and U23968 (N_23968,N_22593,N_22698);
nand U23969 (N_23969,N_22057,N_22928);
xor U23970 (N_23970,N_22798,N_22726);
nor U23971 (N_23971,N_22465,N_22822);
nor U23972 (N_23972,N_22848,N_22429);
and U23973 (N_23973,N_22219,N_22471);
or U23974 (N_23974,N_22275,N_22251);
nand U23975 (N_23975,N_22724,N_22321);
nand U23976 (N_23976,N_22274,N_22639);
nor U23977 (N_23977,N_22470,N_22355);
or U23978 (N_23978,N_22394,N_22346);
nor U23979 (N_23979,N_22092,N_22054);
nor U23980 (N_23980,N_22715,N_22288);
or U23981 (N_23981,N_22014,N_22941);
and U23982 (N_23982,N_22872,N_22651);
or U23983 (N_23983,N_22931,N_22876);
nand U23984 (N_23984,N_22565,N_22486);
or U23985 (N_23985,N_22239,N_22447);
nor U23986 (N_23986,N_22439,N_22867);
nor U23987 (N_23987,N_22681,N_22618);
nor U23988 (N_23988,N_22784,N_22939);
xor U23989 (N_23989,N_22007,N_22899);
and U23990 (N_23990,N_22345,N_22441);
xnor U23991 (N_23991,N_22367,N_22508);
and U23992 (N_23992,N_22193,N_22164);
nand U23993 (N_23993,N_22032,N_22655);
or U23994 (N_23994,N_22369,N_22698);
xnor U23995 (N_23995,N_22913,N_22418);
or U23996 (N_23996,N_22808,N_22381);
nand U23997 (N_23997,N_22381,N_22903);
or U23998 (N_23998,N_22009,N_22144);
nand U23999 (N_23999,N_22382,N_22572);
nand U24000 (N_24000,N_23582,N_23956);
and U24001 (N_24001,N_23487,N_23482);
nor U24002 (N_24002,N_23721,N_23287);
or U24003 (N_24003,N_23369,N_23569);
nand U24004 (N_24004,N_23943,N_23379);
nor U24005 (N_24005,N_23208,N_23404);
and U24006 (N_24006,N_23797,N_23921);
xor U24007 (N_24007,N_23823,N_23019);
nand U24008 (N_24008,N_23554,N_23636);
nand U24009 (N_24009,N_23145,N_23543);
xor U24010 (N_24010,N_23705,N_23164);
nand U24011 (N_24011,N_23461,N_23066);
or U24012 (N_24012,N_23957,N_23684);
or U24013 (N_24013,N_23455,N_23516);
nor U24014 (N_24014,N_23193,N_23565);
or U24015 (N_24015,N_23784,N_23967);
xnor U24016 (N_24016,N_23899,N_23133);
xnor U24017 (N_24017,N_23631,N_23934);
xnor U24018 (N_24018,N_23002,N_23526);
nor U24019 (N_24019,N_23170,N_23521);
and U24020 (N_24020,N_23809,N_23655);
nor U24021 (N_24021,N_23345,N_23220);
nor U24022 (N_24022,N_23732,N_23428);
nand U24023 (N_24023,N_23770,N_23948);
xor U24024 (N_24024,N_23283,N_23387);
nand U24025 (N_24025,N_23878,N_23323);
or U24026 (N_24026,N_23710,N_23058);
nand U24027 (N_24027,N_23557,N_23095);
xor U24028 (N_24028,N_23465,N_23927);
or U24029 (N_24029,N_23272,N_23984);
or U24030 (N_24030,N_23480,N_23911);
or U24031 (N_24031,N_23155,N_23234);
and U24032 (N_24032,N_23832,N_23143);
xor U24033 (N_24033,N_23575,N_23626);
and U24034 (N_24034,N_23925,N_23816);
nand U24035 (N_24035,N_23898,N_23433);
or U24036 (N_24036,N_23835,N_23200);
nor U24037 (N_24037,N_23510,N_23184);
or U24038 (N_24038,N_23817,N_23976);
nor U24039 (N_24039,N_23402,N_23787);
xor U24040 (N_24040,N_23445,N_23698);
or U24041 (N_24041,N_23910,N_23980);
and U24042 (N_24042,N_23897,N_23974);
nand U24043 (N_24043,N_23198,N_23011);
nand U24044 (N_24044,N_23488,N_23504);
and U24045 (N_24045,N_23194,N_23420);
nor U24046 (N_24046,N_23701,N_23879);
nand U24047 (N_24047,N_23667,N_23235);
nand U24048 (N_24048,N_23139,N_23001);
nand U24049 (N_24049,N_23337,N_23138);
and U24050 (N_24050,N_23175,N_23546);
and U24051 (N_24051,N_23434,N_23312);
nor U24052 (N_24052,N_23935,N_23845);
xor U24053 (N_24053,N_23038,N_23328);
xor U24054 (N_24054,N_23396,N_23747);
and U24055 (N_24055,N_23630,N_23755);
and U24056 (N_24056,N_23661,N_23275);
nor U24057 (N_24057,N_23609,N_23243);
xnor U24058 (N_24058,N_23733,N_23665);
xor U24059 (N_24059,N_23421,N_23891);
nand U24060 (N_24060,N_23130,N_23860);
and U24061 (N_24061,N_23375,N_23707);
nor U24062 (N_24062,N_23473,N_23205);
nor U24063 (N_24063,N_23195,N_23033);
nand U24064 (N_24064,N_23830,N_23185);
and U24065 (N_24065,N_23416,N_23996);
or U24066 (N_24066,N_23658,N_23656);
and U24067 (N_24067,N_23127,N_23269);
nor U24068 (N_24068,N_23744,N_23573);
nor U24069 (N_24069,N_23777,N_23886);
or U24070 (N_24070,N_23848,N_23827);
and U24071 (N_24071,N_23334,N_23091);
and U24072 (N_24072,N_23442,N_23076);
nand U24073 (N_24073,N_23893,N_23551);
nand U24074 (N_24074,N_23302,N_23940);
xor U24075 (N_24075,N_23726,N_23637);
nand U24076 (N_24076,N_23278,N_23116);
nor U24077 (N_24077,N_23794,N_23960);
nor U24078 (N_24078,N_23137,N_23591);
nand U24079 (N_24079,N_23715,N_23505);
or U24080 (N_24080,N_23887,N_23883);
or U24081 (N_24081,N_23782,N_23494);
nand U24082 (N_24082,N_23862,N_23840);
nand U24083 (N_24083,N_23238,N_23515);
or U24084 (N_24084,N_23263,N_23252);
and U24085 (N_24085,N_23606,N_23950);
nor U24086 (N_24086,N_23617,N_23540);
nor U24087 (N_24087,N_23563,N_23621);
nand U24088 (N_24088,N_23714,N_23348);
and U24089 (N_24089,N_23588,N_23204);
nor U24090 (N_24090,N_23536,N_23666);
or U24091 (N_24091,N_23178,N_23959);
or U24092 (N_24092,N_23767,N_23431);
or U24093 (N_24093,N_23758,N_23281);
xor U24094 (N_24094,N_23248,N_23983);
or U24095 (N_24095,N_23136,N_23368);
nor U24096 (N_24096,N_23413,N_23232);
or U24097 (N_24097,N_23367,N_23821);
nand U24098 (N_24098,N_23014,N_23293);
nand U24099 (N_24099,N_23214,N_23930);
xnor U24100 (N_24100,N_23928,N_23042);
or U24101 (N_24101,N_23780,N_23620);
nand U24102 (N_24102,N_23037,N_23713);
and U24103 (N_24103,N_23599,N_23892);
xor U24104 (N_24104,N_23868,N_23447);
xor U24105 (N_24105,N_23353,N_23171);
nand U24106 (N_24106,N_23100,N_23507);
xor U24107 (N_24107,N_23598,N_23069);
nor U24108 (N_24108,N_23962,N_23354);
and U24109 (N_24109,N_23295,N_23394);
nand U24110 (N_24110,N_23438,N_23471);
nor U24111 (N_24111,N_23633,N_23933);
and U24112 (N_24112,N_23972,N_23785);
nand U24113 (N_24113,N_23815,N_23305);
nand U24114 (N_24114,N_23687,N_23904);
xnor U24115 (N_24115,N_23228,N_23535);
or U24116 (N_24116,N_23871,N_23056);
nand U24117 (N_24117,N_23239,N_23452);
and U24118 (N_24118,N_23762,N_23463);
nor U24119 (N_24119,N_23577,N_23645);
nand U24120 (N_24120,N_23070,N_23528);
nor U24121 (N_24121,N_23722,N_23788);
nand U24122 (N_24122,N_23912,N_23282);
or U24123 (N_24123,N_23253,N_23285);
nand U24124 (N_24124,N_23458,N_23873);
or U24125 (N_24125,N_23855,N_23724);
xor U24126 (N_24126,N_23059,N_23124);
xor U24127 (N_24127,N_23046,N_23663);
xor U24128 (N_24128,N_23680,N_23807);
or U24129 (N_24129,N_23118,N_23121);
xor U24130 (N_24130,N_23660,N_23920);
nand U24131 (N_24131,N_23783,N_23727);
and U24132 (N_24132,N_23843,N_23558);
nand U24133 (N_24133,N_23335,N_23246);
xor U24134 (N_24134,N_23363,N_23905);
xor U24135 (N_24135,N_23362,N_23392);
nand U24136 (N_24136,N_23849,N_23825);
nor U24137 (N_24137,N_23189,N_23651);
and U24138 (N_24138,N_23530,N_23989);
or U24139 (N_24139,N_23853,N_23015);
xor U24140 (N_24140,N_23219,N_23477);
and U24141 (N_24141,N_23319,N_23481);
and U24142 (N_24142,N_23614,N_23115);
nor U24143 (N_24143,N_23561,N_23939);
nand U24144 (N_24144,N_23364,N_23958);
nand U24145 (N_24145,N_23129,N_23432);
nand U24146 (N_24146,N_23074,N_23737);
nand U24147 (N_24147,N_23225,N_23542);
or U24148 (N_24148,N_23509,N_23885);
and U24149 (N_24149,N_23310,N_23222);
nor U24150 (N_24150,N_23642,N_23766);
nor U24151 (N_24151,N_23229,N_23119);
nand U24152 (N_24152,N_23775,N_23212);
and U24153 (N_24153,N_23901,N_23942);
or U24154 (N_24154,N_23403,N_23632);
nor U24155 (N_24155,N_23114,N_23992);
and U24156 (N_24156,N_23538,N_23023);
nand U24157 (N_24157,N_23771,N_23067);
nor U24158 (N_24158,N_23479,N_23694);
or U24159 (N_24159,N_23411,N_23035);
and U24160 (N_24160,N_23993,N_23531);
or U24161 (N_24161,N_23099,N_23051);
or U24162 (N_24162,N_23102,N_23435);
or U24163 (N_24163,N_23690,N_23215);
and U24164 (N_24164,N_23749,N_23007);
nand U24165 (N_24165,N_23547,N_23358);
nand U24166 (N_24166,N_23670,N_23768);
and U24167 (N_24167,N_23450,N_23408);
nand U24168 (N_24168,N_23604,N_23679);
and U24169 (N_24169,N_23997,N_23415);
nor U24170 (N_24170,N_23708,N_23826);
nor U24171 (N_24171,N_23031,N_23339);
nand U24172 (N_24172,N_23559,N_23789);
xnor U24173 (N_24173,N_23859,N_23361);
xor U24174 (N_24174,N_23365,N_23329);
or U24175 (N_24175,N_23806,N_23401);
or U24176 (N_24176,N_23009,N_23987);
or U24177 (N_24177,N_23090,N_23266);
or U24178 (N_24178,N_23330,N_23915);
or U24179 (N_24179,N_23810,N_23233);
nand U24180 (N_24180,N_23366,N_23196);
nor U24181 (N_24181,N_23357,N_23792);
and U24182 (N_24182,N_23944,N_23791);
nor U24183 (N_24183,N_23192,N_23795);
and U24184 (N_24184,N_23981,N_23340);
and U24185 (N_24185,N_23664,N_23341);
or U24186 (N_24186,N_23439,N_23390);
xor U24187 (N_24187,N_23267,N_23616);
nor U24188 (N_24188,N_23371,N_23103);
nand U24189 (N_24189,N_23055,N_23227);
nand U24190 (N_24190,N_23486,N_23751);
xnor U24191 (N_24191,N_23608,N_23838);
xor U24192 (N_24192,N_23533,N_23648);
nand U24193 (N_24193,N_23050,N_23571);
nand U24194 (N_24194,N_23167,N_23472);
and U24195 (N_24195,N_23088,N_23240);
xnor U24196 (N_24196,N_23894,N_23493);
nor U24197 (N_24197,N_23678,N_23740);
and U24198 (N_24198,N_23796,N_23441);
and U24199 (N_24199,N_23596,N_23382);
nor U24200 (N_24200,N_23414,N_23866);
or U24201 (N_24201,N_23818,N_23120);
nor U24202 (N_24202,N_23029,N_23291);
or U24203 (N_24203,N_23875,N_23147);
and U24204 (N_24204,N_23083,N_23057);
nor U24205 (N_24205,N_23410,N_23326);
and U24206 (N_24206,N_23929,N_23292);
xor U24207 (N_24207,N_23581,N_23372);
nand U24208 (N_24208,N_23534,N_23675);
or U24209 (N_24209,N_23047,N_23824);
xnor U24210 (N_24210,N_23869,N_23462);
and U24211 (N_24211,N_23496,N_23627);
and U24212 (N_24212,N_23995,N_23677);
and U24213 (N_24213,N_23322,N_23761);
xor U24214 (N_24214,N_23146,N_23580);
nand U24215 (N_24215,N_23622,N_23584);
or U24216 (N_24216,N_23065,N_23045);
nor U24217 (N_24217,N_23373,N_23804);
nor U24218 (N_24218,N_23748,N_23464);
nor U24219 (N_24219,N_23643,N_23113);
nand U24220 (N_24220,N_23590,N_23570);
and U24221 (N_24221,N_23021,N_23026);
and U24222 (N_24222,N_23044,N_23881);
nor U24223 (N_24223,N_23603,N_23209);
nor U24224 (N_24224,N_23393,N_23491);
nand U24225 (N_24225,N_23437,N_23468);
nand U24226 (N_24226,N_23978,N_23126);
nor U24227 (N_24227,N_23641,N_23560);
nor U24228 (N_24228,N_23895,N_23772);
or U24229 (N_24229,N_23311,N_23903);
and U24230 (N_24230,N_23865,N_23159);
xnor U24231 (N_24231,N_23638,N_23412);
and U24232 (N_24232,N_23982,N_23218);
nor U24233 (N_24233,N_23512,N_23877);
xor U24234 (N_24234,N_23304,N_23717);
nand U24235 (N_24235,N_23738,N_23852);
xor U24236 (N_24236,N_23634,N_23841);
nand U24237 (N_24237,N_23320,N_23203);
nor U24238 (N_24238,N_23757,N_23681);
or U24239 (N_24239,N_23025,N_23084);
and U24240 (N_24240,N_23592,N_23990);
nand U24241 (N_24241,N_23562,N_23237);
or U24242 (N_24242,N_23858,N_23216);
or U24243 (N_24243,N_23250,N_23276);
nor U24244 (N_24244,N_23446,N_23896);
or U24245 (N_24245,N_23629,N_23331);
nor U24246 (N_24246,N_23712,N_23469);
nor U24247 (N_24247,N_23376,N_23112);
or U24248 (N_24248,N_23064,N_23254);
xor U24249 (N_24249,N_23075,N_23579);
nand U24250 (N_24250,N_23107,N_23359);
and U24251 (N_24251,N_23600,N_23842);
and U24252 (N_24252,N_23188,N_23979);
xnor U24253 (N_24253,N_23585,N_23476);
nand U24254 (N_24254,N_23650,N_23077);
or U24255 (N_24255,N_23160,N_23425);
nand U24256 (N_24256,N_23882,N_23153);
nand U24257 (N_24257,N_23436,N_23131);
xnor U24258 (N_24258,N_23524,N_23583);
and U24259 (N_24259,N_23743,N_23764);
xor U24260 (N_24260,N_23729,N_23702);
nor U24261 (N_24261,N_23773,N_23094);
nor U24262 (N_24262,N_23296,N_23259);
and U24263 (N_24263,N_23264,N_23224);
nand U24264 (N_24264,N_23079,N_23087);
and U24265 (N_24265,N_23819,N_23041);
nor U24266 (N_24266,N_23669,N_23833);
nand U24267 (N_24267,N_23300,N_23048);
nand U24268 (N_24268,N_23696,N_23072);
or U24269 (N_24269,N_23970,N_23578);
nand U24270 (N_24270,N_23166,N_23625);
nor U24271 (N_24271,N_23697,N_23514);
or U24272 (N_24272,N_23662,N_23973);
and U24273 (N_24273,N_23676,N_23036);
nor U24274 (N_24274,N_23602,N_23231);
nand U24275 (N_24275,N_23333,N_23242);
nand U24276 (N_24276,N_23187,N_23975);
nand U24277 (N_24277,N_23098,N_23135);
and U24278 (N_24278,N_23279,N_23385);
nand U24279 (N_24279,N_23556,N_23741);
or U24280 (N_24280,N_23502,N_23418);
xor U24281 (N_24281,N_23836,N_23965);
and U24282 (N_24282,N_23256,N_23105);
or U24283 (N_24283,N_23101,N_23900);
nand U24284 (N_24284,N_23478,N_23406);
nand U24285 (N_24285,N_23321,N_23870);
and U24286 (N_24286,N_23597,N_23117);
and U24287 (N_24287,N_23255,N_23844);
and U24288 (N_24288,N_23356,N_23917);
and U24289 (N_24289,N_23988,N_23347);
nor U24290 (N_24290,N_23889,N_23317);
or U24291 (N_24291,N_23244,N_23265);
nor U24292 (N_24292,N_23013,N_23409);
nor U24293 (N_24293,N_23539,N_23020);
xnor U24294 (N_24294,N_23258,N_23888);
and U24295 (N_24295,N_23230,N_23467);
and U24296 (N_24296,N_23709,N_23168);
nor U24297 (N_24297,N_23008,N_23398);
xnor U24298 (N_24298,N_23776,N_23532);
and U24299 (N_24299,N_23805,N_23052);
xnor U24300 (N_24300,N_23649,N_23210);
and U24301 (N_24301,N_23183,N_23874);
nor U24302 (N_24302,N_23123,N_23395);
nand U24303 (N_24303,N_23426,N_23864);
nor U24304 (N_24304,N_23288,N_23190);
nand U24305 (N_24305,N_23032,N_23611);
nand U24306 (N_24306,N_23191,N_23812);
nor U24307 (N_24307,N_23271,N_23399);
nor U24308 (N_24308,N_23097,N_23765);
or U24309 (N_24309,N_23994,N_23861);
nand U24310 (N_24310,N_23682,N_23977);
nand U24311 (N_24311,N_23144,N_23344);
nand U24312 (N_24312,N_23377,N_23017);
or U24313 (N_24313,N_23711,N_23954);
or U24314 (N_24314,N_23572,N_23683);
and U24315 (N_24315,N_23104,N_23180);
or U24316 (N_24316,N_23890,N_23407);
nor U24317 (N_24317,N_23484,N_23417);
xor U24318 (N_24318,N_23273,N_23553);
nor U24319 (N_24319,N_23595,N_23061);
nor U24320 (N_24320,N_23027,N_23644);
xnor U24321 (N_24321,N_23054,N_23063);
xnor U24322 (N_24322,N_23245,N_23525);
xnor U24323 (N_24323,N_23610,N_23814);
xor U24324 (N_24324,N_23945,N_23924);
nor U24325 (N_24325,N_23423,N_23280);
or U24326 (N_24326,N_23400,N_23004);
xnor U24327 (N_24327,N_23820,N_23798);
nand U24328 (N_24328,N_23086,N_23926);
and U24329 (N_24329,N_23759,N_23342);
xnor U24330 (N_24330,N_23274,N_23251);
nand U24331 (N_24331,N_23549,N_23257);
xor U24332 (N_24332,N_23918,N_23781);
or U24333 (N_24333,N_23746,N_23386);
nor U24334 (N_24334,N_23492,N_23763);
nand U24335 (N_24335,N_23217,N_23449);
xnor U24336 (N_24336,N_23700,N_23932);
nor U24337 (N_24337,N_23654,N_23081);
or U24338 (N_24338,N_23018,N_23298);
and U24339 (N_24339,N_23919,N_23022);
nand U24340 (N_24340,N_23652,N_23774);
nor U24341 (N_24341,N_23173,N_23628);
nor U24342 (N_24342,N_23005,N_23564);
nand U24343 (N_24343,N_23270,N_23043);
nand U24344 (N_24344,N_23779,N_23503);
nor U24345 (N_24345,N_23040,N_23750);
nor U24346 (N_24346,N_23914,N_23586);
nand U24347 (N_24347,N_23306,N_23589);
or U24348 (N_24348,N_23688,N_23163);
or U24349 (N_24349,N_23725,N_23080);
or U24350 (N_24350,N_23092,N_23388);
and U24351 (N_24351,N_23073,N_23938);
nor U24352 (N_24352,N_23448,N_23529);
nand U24353 (N_24353,N_23686,N_23734);
nor U24354 (N_24354,N_23947,N_23140);
nor U24355 (N_24355,N_23062,N_23111);
or U24356 (N_24356,N_23955,N_23391);
nor U24357 (N_24357,N_23157,N_23381);
or U24358 (N_24358,N_23325,N_23501);
xnor U24359 (N_24359,N_23207,N_23152);
nand U24360 (N_24360,N_23703,N_23016);
and U24361 (N_24361,N_23850,N_23922);
nand U24362 (N_24362,N_23953,N_23324);
xor U24363 (N_24363,N_23837,N_23618);
xnor U24364 (N_24364,N_23012,N_23695);
or U24365 (N_24365,N_23769,N_23498);
xor U24366 (N_24366,N_23752,N_23223);
and U24367 (N_24367,N_23566,N_23182);
nor U24368 (N_24368,N_23659,N_23673);
nand U24369 (N_24369,N_23527,N_23440);
and U24370 (N_24370,N_23277,N_23884);
nand U24371 (N_24371,N_23568,N_23247);
xor U24372 (N_24372,N_23813,N_23704);
and U24373 (N_24373,N_23459,N_23500);
and U24374 (N_24374,N_23110,N_23172);
or U24375 (N_24375,N_23262,N_23151);
and U24376 (N_24376,N_23613,N_23719);
xor U24377 (N_24377,N_23671,N_23149);
nand U24378 (N_24378,N_23349,N_23511);
nand U24379 (N_24379,N_23906,N_23537);
and U24380 (N_24380,N_23174,N_23158);
xor U24381 (N_24381,N_23261,N_23854);
nor U24382 (N_24382,N_23313,N_23847);
and U24383 (N_24383,N_23093,N_23483);
xnor U24384 (N_24384,N_23457,N_23699);
or U24385 (N_24385,N_23552,N_23615);
xor U24386 (N_24386,N_23177,N_23451);
or U24387 (N_24387,N_23730,N_23010);
xor U24388 (N_24388,N_23513,N_23307);
xnor U24389 (N_24389,N_23653,N_23343);
or U24390 (N_24390,N_23474,N_23199);
xnor U24391 (N_24391,N_23460,N_23692);
and U24392 (N_24392,N_23808,N_23786);
nand U24393 (N_24393,N_23268,N_23221);
nand U24394 (N_24394,N_23165,N_23141);
or U24395 (N_24395,N_23060,N_23723);
nand U24396 (N_24396,N_23108,N_23518);
or U24397 (N_24397,N_23249,N_23134);
nand U24398 (N_24398,N_23085,N_23360);
xor U24399 (N_24399,N_23444,N_23986);
nor U24400 (N_24400,N_23380,N_23639);
nor U24401 (N_24401,N_23370,N_23148);
nand U24402 (N_24402,N_23132,N_23475);
xor U24403 (N_24403,N_23049,N_23497);
xnor U24404 (N_24404,N_23422,N_23756);
or U24405 (N_24405,N_23213,N_23355);
nor U24406 (N_24406,N_23966,N_23156);
or U24407 (N_24407,N_23576,N_23424);
and U24408 (N_24408,N_23499,N_23693);
and U24409 (N_24409,N_23941,N_23829);
xor U24410 (N_24410,N_23674,N_23623);
or U24411 (N_24411,N_23969,N_23383);
and U24412 (N_24412,N_23397,N_23857);
nor U24413 (N_24413,N_23211,N_23946);
nand U24414 (N_24414,N_23053,N_23068);
nor U24415 (N_24415,N_23574,N_23071);
xnor U24416 (N_24416,N_23519,N_23952);
or U24417 (N_24417,N_23991,N_23754);
nand U24418 (N_24418,N_23856,N_23909);
and U24419 (N_24419,N_23142,N_23739);
xor U24420 (N_24420,N_23485,N_23949);
nor U24421 (N_24421,N_23640,N_23802);
nand U24422 (N_24422,N_23299,N_23799);
nand U24423 (N_24423,N_23389,N_23454);
and U24424 (N_24424,N_23161,N_23689);
and U24425 (N_24425,N_23872,N_23619);
nor U24426 (N_24426,N_23520,N_23150);
or U24427 (N_24427,N_23290,N_23508);
or U24428 (N_24428,N_23587,N_23309);
or U24429 (N_24429,N_23913,N_23332);
nor U24430 (N_24430,N_23506,N_23206);
nor U24431 (N_24431,N_23202,N_23923);
xor U24432 (N_24432,N_23828,N_23753);
nor U24433 (N_24433,N_23624,N_23003);
xnor U24434 (N_24434,N_23303,N_23024);
xor U24435 (N_24435,N_23880,N_23963);
xor U24436 (N_24436,N_23286,N_23831);
or U24437 (N_24437,N_23668,N_23490);
or U24438 (N_24438,N_23594,N_23778);
xnor U24439 (N_24439,N_23811,N_23998);
nand U24440 (N_24440,N_23236,N_23327);
nand U24441 (N_24441,N_23907,N_23523);
nand U24442 (N_24442,N_23284,N_23541);
and U24443 (N_24443,N_23039,N_23720);
and U24444 (N_24444,N_23028,N_23226);
xor U24445 (N_24445,N_23834,N_23089);
nor U24446 (N_24446,N_23078,N_23867);
and U24447 (N_24447,N_23308,N_23034);
nand U24448 (N_24448,N_23352,N_23672);
nor U24449 (N_24449,N_23745,N_23790);
or U24450 (N_24450,N_23154,N_23593);
nor U24451 (N_24451,N_23961,N_23801);
and U24452 (N_24452,N_23106,N_23489);
nand U24453 (N_24453,N_23350,N_23082);
xnor U24454 (N_24454,N_23470,N_23122);
xor U24455 (N_24455,N_23346,N_23742);
xnor U24456 (N_24456,N_23916,N_23931);
nor U24457 (N_24457,N_23793,N_23241);
xor U24458 (N_24458,N_23125,N_23294);
and U24459 (N_24459,N_23181,N_23384);
and U24460 (N_24460,N_23453,N_23456);
and U24461 (N_24461,N_23544,N_23443);
nand U24462 (N_24462,N_23006,N_23876);
nor U24463 (N_24463,N_23545,N_23260);
nor U24464 (N_24464,N_23657,N_23378);
nand U24465 (N_24465,N_23405,N_23601);
xor U24466 (N_24466,N_23419,N_23128);
xor U24467 (N_24467,N_23316,N_23522);
nand U24468 (N_24468,N_23176,N_23338);
or U24469 (N_24469,N_23646,N_23550);
or U24470 (N_24470,N_23186,N_23803);
nand U24471 (N_24471,N_23736,N_23548);
or U24472 (N_24472,N_23691,N_23968);
or U24473 (N_24473,N_23297,N_23985);
xor U24474 (N_24474,N_23517,N_23971);
or U24475 (N_24475,N_23902,N_23863);
and U24476 (N_24476,N_23951,N_23466);
xor U24477 (N_24477,N_23685,N_23201);
xnor U24478 (N_24478,N_23999,N_23289);
or U24479 (N_24479,N_23937,N_23567);
and U24480 (N_24480,N_23555,N_23495);
nand U24481 (N_24481,N_23336,N_23318);
nand U24482 (N_24482,N_23612,N_23030);
or U24483 (N_24483,N_23429,N_23374);
nor U24484 (N_24484,N_23822,N_23908);
or U24485 (N_24485,N_23846,N_23000);
or U24486 (N_24486,N_23800,N_23301);
or U24487 (N_24487,N_23315,N_23635);
and U24488 (N_24488,N_23430,N_23197);
nor U24489 (N_24489,N_23427,N_23731);
xnor U24490 (N_24490,N_23936,N_23728);
and U24491 (N_24491,N_23647,N_23839);
and U24492 (N_24492,N_23605,N_23179);
and U24493 (N_24493,N_23162,N_23851);
and U24494 (N_24494,N_23706,N_23109);
nor U24495 (N_24495,N_23964,N_23096);
nor U24496 (N_24496,N_23718,N_23735);
xnor U24497 (N_24497,N_23607,N_23760);
xnor U24498 (N_24498,N_23314,N_23169);
and U24499 (N_24499,N_23716,N_23351);
and U24500 (N_24500,N_23044,N_23280);
xnor U24501 (N_24501,N_23498,N_23181);
xor U24502 (N_24502,N_23790,N_23170);
xnor U24503 (N_24503,N_23928,N_23662);
xnor U24504 (N_24504,N_23003,N_23554);
nor U24505 (N_24505,N_23237,N_23586);
nor U24506 (N_24506,N_23060,N_23941);
xor U24507 (N_24507,N_23854,N_23522);
and U24508 (N_24508,N_23197,N_23427);
nor U24509 (N_24509,N_23295,N_23813);
nor U24510 (N_24510,N_23175,N_23021);
nor U24511 (N_24511,N_23759,N_23034);
or U24512 (N_24512,N_23858,N_23961);
and U24513 (N_24513,N_23038,N_23464);
or U24514 (N_24514,N_23783,N_23018);
and U24515 (N_24515,N_23669,N_23845);
or U24516 (N_24516,N_23269,N_23068);
xor U24517 (N_24517,N_23177,N_23701);
and U24518 (N_24518,N_23211,N_23856);
or U24519 (N_24519,N_23287,N_23267);
nor U24520 (N_24520,N_23490,N_23818);
nand U24521 (N_24521,N_23465,N_23540);
nor U24522 (N_24522,N_23400,N_23755);
and U24523 (N_24523,N_23969,N_23883);
and U24524 (N_24524,N_23225,N_23432);
xor U24525 (N_24525,N_23105,N_23418);
xor U24526 (N_24526,N_23906,N_23217);
and U24527 (N_24527,N_23957,N_23479);
nor U24528 (N_24528,N_23557,N_23498);
or U24529 (N_24529,N_23501,N_23965);
xor U24530 (N_24530,N_23345,N_23493);
or U24531 (N_24531,N_23280,N_23272);
or U24532 (N_24532,N_23199,N_23560);
nand U24533 (N_24533,N_23118,N_23706);
nand U24534 (N_24534,N_23404,N_23660);
nor U24535 (N_24535,N_23848,N_23335);
xnor U24536 (N_24536,N_23052,N_23295);
or U24537 (N_24537,N_23974,N_23015);
nor U24538 (N_24538,N_23689,N_23870);
or U24539 (N_24539,N_23036,N_23512);
and U24540 (N_24540,N_23620,N_23064);
nor U24541 (N_24541,N_23771,N_23206);
nand U24542 (N_24542,N_23234,N_23671);
xor U24543 (N_24543,N_23505,N_23128);
or U24544 (N_24544,N_23221,N_23312);
or U24545 (N_24545,N_23458,N_23060);
nor U24546 (N_24546,N_23303,N_23154);
xor U24547 (N_24547,N_23301,N_23599);
or U24548 (N_24548,N_23045,N_23620);
xor U24549 (N_24549,N_23290,N_23123);
nand U24550 (N_24550,N_23429,N_23233);
and U24551 (N_24551,N_23875,N_23702);
nand U24552 (N_24552,N_23115,N_23028);
and U24553 (N_24553,N_23216,N_23879);
nor U24554 (N_24554,N_23362,N_23460);
nor U24555 (N_24555,N_23412,N_23985);
or U24556 (N_24556,N_23238,N_23835);
nor U24557 (N_24557,N_23895,N_23418);
nor U24558 (N_24558,N_23978,N_23330);
xnor U24559 (N_24559,N_23401,N_23767);
and U24560 (N_24560,N_23435,N_23000);
and U24561 (N_24561,N_23969,N_23530);
xor U24562 (N_24562,N_23616,N_23525);
xor U24563 (N_24563,N_23373,N_23324);
nand U24564 (N_24564,N_23940,N_23387);
nand U24565 (N_24565,N_23306,N_23025);
or U24566 (N_24566,N_23740,N_23040);
nand U24567 (N_24567,N_23629,N_23991);
or U24568 (N_24568,N_23267,N_23187);
or U24569 (N_24569,N_23713,N_23884);
and U24570 (N_24570,N_23677,N_23854);
or U24571 (N_24571,N_23397,N_23153);
xor U24572 (N_24572,N_23518,N_23753);
xnor U24573 (N_24573,N_23589,N_23506);
or U24574 (N_24574,N_23160,N_23421);
and U24575 (N_24575,N_23663,N_23840);
or U24576 (N_24576,N_23481,N_23842);
nand U24577 (N_24577,N_23543,N_23165);
or U24578 (N_24578,N_23336,N_23688);
xnor U24579 (N_24579,N_23726,N_23227);
or U24580 (N_24580,N_23306,N_23640);
or U24581 (N_24581,N_23026,N_23834);
or U24582 (N_24582,N_23324,N_23530);
or U24583 (N_24583,N_23659,N_23283);
xor U24584 (N_24584,N_23773,N_23724);
nor U24585 (N_24585,N_23318,N_23482);
and U24586 (N_24586,N_23158,N_23709);
nand U24587 (N_24587,N_23165,N_23527);
nand U24588 (N_24588,N_23194,N_23604);
nand U24589 (N_24589,N_23319,N_23742);
xor U24590 (N_24590,N_23406,N_23759);
nor U24591 (N_24591,N_23137,N_23413);
or U24592 (N_24592,N_23577,N_23186);
nand U24593 (N_24593,N_23204,N_23262);
xor U24594 (N_24594,N_23007,N_23155);
or U24595 (N_24595,N_23907,N_23088);
nor U24596 (N_24596,N_23233,N_23608);
nand U24597 (N_24597,N_23104,N_23846);
and U24598 (N_24598,N_23445,N_23819);
and U24599 (N_24599,N_23530,N_23598);
and U24600 (N_24600,N_23843,N_23281);
and U24601 (N_24601,N_23419,N_23054);
nand U24602 (N_24602,N_23696,N_23901);
xnor U24603 (N_24603,N_23644,N_23744);
nor U24604 (N_24604,N_23527,N_23092);
nor U24605 (N_24605,N_23403,N_23866);
xor U24606 (N_24606,N_23788,N_23441);
and U24607 (N_24607,N_23300,N_23705);
or U24608 (N_24608,N_23841,N_23198);
xnor U24609 (N_24609,N_23853,N_23326);
nor U24610 (N_24610,N_23508,N_23293);
xnor U24611 (N_24611,N_23056,N_23810);
or U24612 (N_24612,N_23258,N_23615);
nor U24613 (N_24613,N_23775,N_23080);
nor U24614 (N_24614,N_23521,N_23740);
or U24615 (N_24615,N_23907,N_23272);
nand U24616 (N_24616,N_23698,N_23796);
nand U24617 (N_24617,N_23022,N_23920);
xor U24618 (N_24618,N_23172,N_23313);
nand U24619 (N_24619,N_23319,N_23927);
nor U24620 (N_24620,N_23988,N_23572);
nand U24621 (N_24621,N_23642,N_23536);
nand U24622 (N_24622,N_23482,N_23833);
and U24623 (N_24623,N_23157,N_23318);
and U24624 (N_24624,N_23122,N_23461);
nand U24625 (N_24625,N_23714,N_23831);
xor U24626 (N_24626,N_23389,N_23381);
nor U24627 (N_24627,N_23164,N_23263);
nand U24628 (N_24628,N_23875,N_23965);
and U24629 (N_24629,N_23208,N_23901);
xnor U24630 (N_24630,N_23204,N_23957);
nor U24631 (N_24631,N_23356,N_23161);
xnor U24632 (N_24632,N_23632,N_23404);
xnor U24633 (N_24633,N_23658,N_23366);
nand U24634 (N_24634,N_23710,N_23844);
or U24635 (N_24635,N_23389,N_23990);
xor U24636 (N_24636,N_23211,N_23894);
or U24637 (N_24637,N_23090,N_23239);
nor U24638 (N_24638,N_23166,N_23754);
nand U24639 (N_24639,N_23544,N_23382);
and U24640 (N_24640,N_23607,N_23595);
and U24641 (N_24641,N_23295,N_23678);
and U24642 (N_24642,N_23650,N_23073);
and U24643 (N_24643,N_23486,N_23948);
and U24644 (N_24644,N_23190,N_23036);
nor U24645 (N_24645,N_23353,N_23339);
or U24646 (N_24646,N_23697,N_23523);
or U24647 (N_24647,N_23418,N_23055);
nand U24648 (N_24648,N_23594,N_23222);
nor U24649 (N_24649,N_23674,N_23888);
xor U24650 (N_24650,N_23753,N_23461);
and U24651 (N_24651,N_23379,N_23589);
nand U24652 (N_24652,N_23178,N_23824);
and U24653 (N_24653,N_23568,N_23467);
nand U24654 (N_24654,N_23645,N_23740);
and U24655 (N_24655,N_23250,N_23347);
nand U24656 (N_24656,N_23849,N_23268);
nand U24657 (N_24657,N_23910,N_23425);
nand U24658 (N_24658,N_23499,N_23161);
nand U24659 (N_24659,N_23951,N_23624);
nand U24660 (N_24660,N_23141,N_23795);
nand U24661 (N_24661,N_23865,N_23995);
and U24662 (N_24662,N_23921,N_23347);
and U24663 (N_24663,N_23963,N_23102);
and U24664 (N_24664,N_23969,N_23354);
or U24665 (N_24665,N_23358,N_23415);
or U24666 (N_24666,N_23979,N_23444);
nor U24667 (N_24667,N_23871,N_23023);
or U24668 (N_24668,N_23027,N_23928);
and U24669 (N_24669,N_23337,N_23802);
nor U24670 (N_24670,N_23347,N_23941);
or U24671 (N_24671,N_23467,N_23087);
nor U24672 (N_24672,N_23501,N_23366);
or U24673 (N_24673,N_23636,N_23638);
or U24674 (N_24674,N_23062,N_23904);
nand U24675 (N_24675,N_23138,N_23942);
and U24676 (N_24676,N_23819,N_23388);
nor U24677 (N_24677,N_23066,N_23925);
xnor U24678 (N_24678,N_23828,N_23936);
xor U24679 (N_24679,N_23496,N_23876);
and U24680 (N_24680,N_23244,N_23401);
or U24681 (N_24681,N_23413,N_23224);
and U24682 (N_24682,N_23413,N_23029);
and U24683 (N_24683,N_23419,N_23160);
nand U24684 (N_24684,N_23057,N_23609);
nor U24685 (N_24685,N_23506,N_23200);
and U24686 (N_24686,N_23750,N_23905);
xor U24687 (N_24687,N_23098,N_23363);
nor U24688 (N_24688,N_23923,N_23119);
nand U24689 (N_24689,N_23310,N_23739);
nor U24690 (N_24690,N_23770,N_23698);
xor U24691 (N_24691,N_23642,N_23545);
and U24692 (N_24692,N_23339,N_23721);
or U24693 (N_24693,N_23559,N_23134);
nor U24694 (N_24694,N_23336,N_23271);
or U24695 (N_24695,N_23624,N_23373);
or U24696 (N_24696,N_23896,N_23701);
nand U24697 (N_24697,N_23809,N_23883);
nor U24698 (N_24698,N_23373,N_23226);
and U24699 (N_24699,N_23978,N_23908);
and U24700 (N_24700,N_23761,N_23654);
or U24701 (N_24701,N_23315,N_23902);
and U24702 (N_24702,N_23223,N_23638);
nand U24703 (N_24703,N_23978,N_23828);
or U24704 (N_24704,N_23391,N_23962);
and U24705 (N_24705,N_23535,N_23651);
nor U24706 (N_24706,N_23965,N_23227);
nand U24707 (N_24707,N_23775,N_23710);
xor U24708 (N_24708,N_23898,N_23142);
and U24709 (N_24709,N_23276,N_23695);
or U24710 (N_24710,N_23323,N_23228);
or U24711 (N_24711,N_23339,N_23263);
nor U24712 (N_24712,N_23109,N_23990);
and U24713 (N_24713,N_23428,N_23519);
nand U24714 (N_24714,N_23361,N_23528);
nand U24715 (N_24715,N_23815,N_23803);
and U24716 (N_24716,N_23197,N_23105);
nor U24717 (N_24717,N_23836,N_23675);
nor U24718 (N_24718,N_23134,N_23737);
nand U24719 (N_24719,N_23446,N_23514);
nand U24720 (N_24720,N_23834,N_23594);
xnor U24721 (N_24721,N_23558,N_23421);
xor U24722 (N_24722,N_23682,N_23497);
or U24723 (N_24723,N_23422,N_23221);
or U24724 (N_24724,N_23717,N_23834);
nor U24725 (N_24725,N_23334,N_23399);
and U24726 (N_24726,N_23731,N_23690);
nor U24727 (N_24727,N_23064,N_23380);
xnor U24728 (N_24728,N_23904,N_23582);
or U24729 (N_24729,N_23964,N_23127);
xor U24730 (N_24730,N_23711,N_23765);
or U24731 (N_24731,N_23367,N_23055);
xnor U24732 (N_24732,N_23896,N_23192);
xor U24733 (N_24733,N_23684,N_23936);
nand U24734 (N_24734,N_23248,N_23021);
and U24735 (N_24735,N_23415,N_23648);
xor U24736 (N_24736,N_23947,N_23116);
xnor U24737 (N_24737,N_23251,N_23690);
nand U24738 (N_24738,N_23903,N_23488);
or U24739 (N_24739,N_23062,N_23245);
nand U24740 (N_24740,N_23340,N_23284);
and U24741 (N_24741,N_23032,N_23599);
or U24742 (N_24742,N_23988,N_23410);
and U24743 (N_24743,N_23461,N_23258);
xor U24744 (N_24744,N_23792,N_23124);
or U24745 (N_24745,N_23827,N_23330);
and U24746 (N_24746,N_23859,N_23123);
or U24747 (N_24747,N_23644,N_23211);
and U24748 (N_24748,N_23792,N_23906);
nor U24749 (N_24749,N_23233,N_23297);
or U24750 (N_24750,N_23526,N_23421);
nand U24751 (N_24751,N_23020,N_23596);
and U24752 (N_24752,N_23545,N_23372);
and U24753 (N_24753,N_23459,N_23725);
nor U24754 (N_24754,N_23953,N_23913);
xor U24755 (N_24755,N_23045,N_23673);
xnor U24756 (N_24756,N_23142,N_23568);
xnor U24757 (N_24757,N_23890,N_23815);
xor U24758 (N_24758,N_23845,N_23325);
nand U24759 (N_24759,N_23253,N_23556);
nand U24760 (N_24760,N_23472,N_23524);
xor U24761 (N_24761,N_23761,N_23403);
nand U24762 (N_24762,N_23321,N_23565);
or U24763 (N_24763,N_23226,N_23811);
nor U24764 (N_24764,N_23617,N_23942);
nand U24765 (N_24765,N_23065,N_23213);
nand U24766 (N_24766,N_23371,N_23129);
and U24767 (N_24767,N_23529,N_23095);
or U24768 (N_24768,N_23636,N_23291);
nand U24769 (N_24769,N_23759,N_23372);
xnor U24770 (N_24770,N_23490,N_23369);
nor U24771 (N_24771,N_23964,N_23419);
nor U24772 (N_24772,N_23718,N_23839);
xor U24773 (N_24773,N_23775,N_23564);
and U24774 (N_24774,N_23533,N_23562);
or U24775 (N_24775,N_23499,N_23728);
or U24776 (N_24776,N_23528,N_23957);
or U24777 (N_24777,N_23830,N_23439);
nand U24778 (N_24778,N_23916,N_23255);
nor U24779 (N_24779,N_23494,N_23215);
nand U24780 (N_24780,N_23852,N_23222);
and U24781 (N_24781,N_23680,N_23746);
and U24782 (N_24782,N_23873,N_23861);
and U24783 (N_24783,N_23904,N_23996);
nand U24784 (N_24784,N_23816,N_23489);
nor U24785 (N_24785,N_23790,N_23558);
or U24786 (N_24786,N_23138,N_23318);
or U24787 (N_24787,N_23396,N_23278);
or U24788 (N_24788,N_23181,N_23945);
nand U24789 (N_24789,N_23649,N_23809);
or U24790 (N_24790,N_23826,N_23536);
or U24791 (N_24791,N_23317,N_23897);
nor U24792 (N_24792,N_23824,N_23624);
xnor U24793 (N_24793,N_23161,N_23424);
nor U24794 (N_24794,N_23115,N_23168);
or U24795 (N_24795,N_23070,N_23127);
nor U24796 (N_24796,N_23793,N_23975);
xor U24797 (N_24797,N_23203,N_23928);
or U24798 (N_24798,N_23338,N_23737);
nor U24799 (N_24799,N_23855,N_23861);
nor U24800 (N_24800,N_23791,N_23288);
or U24801 (N_24801,N_23724,N_23952);
or U24802 (N_24802,N_23546,N_23213);
nand U24803 (N_24803,N_23856,N_23496);
or U24804 (N_24804,N_23994,N_23605);
or U24805 (N_24805,N_23335,N_23153);
nor U24806 (N_24806,N_23592,N_23784);
nor U24807 (N_24807,N_23221,N_23953);
nand U24808 (N_24808,N_23534,N_23321);
and U24809 (N_24809,N_23069,N_23442);
nand U24810 (N_24810,N_23332,N_23717);
and U24811 (N_24811,N_23901,N_23131);
and U24812 (N_24812,N_23936,N_23352);
or U24813 (N_24813,N_23138,N_23243);
or U24814 (N_24814,N_23658,N_23377);
nor U24815 (N_24815,N_23058,N_23872);
xor U24816 (N_24816,N_23174,N_23854);
nand U24817 (N_24817,N_23943,N_23625);
or U24818 (N_24818,N_23206,N_23134);
and U24819 (N_24819,N_23087,N_23488);
or U24820 (N_24820,N_23685,N_23375);
or U24821 (N_24821,N_23929,N_23443);
and U24822 (N_24822,N_23144,N_23014);
and U24823 (N_24823,N_23852,N_23618);
or U24824 (N_24824,N_23290,N_23942);
nor U24825 (N_24825,N_23989,N_23555);
and U24826 (N_24826,N_23111,N_23651);
and U24827 (N_24827,N_23603,N_23543);
nand U24828 (N_24828,N_23463,N_23528);
xor U24829 (N_24829,N_23395,N_23755);
xor U24830 (N_24830,N_23312,N_23907);
xor U24831 (N_24831,N_23400,N_23589);
and U24832 (N_24832,N_23302,N_23799);
or U24833 (N_24833,N_23847,N_23830);
nand U24834 (N_24834,N_23602,N_23046);
or U24835 (N_24835,N_23217,N_23862);
nor U24836 (N_24836,N_23942,N_23482);
xor U24837 (N_24837,N_23351,N_23483);
nand U24838 (N_24838,N_23524,N_23550);
xor U24839 (N_24839,N_23230,N_23083);
or U24840 (N_24840,N_23545,N_23800);
nor U24841 (N_24841,N_23875,N_23327);
and U24842 (N_24842,N_23240,N_23260);
and U24843 (N_24843,N_23003,N_23270);
or U24844 (N_24844,N_23975,N_23212);
or U24845 (N_24845,N_23789,N_23643);
xor U24846 (N_24846,N_23007,N_23012);
nand U24847 (N_24847,N_23664,N_23921);
and U24848 (N_24848,N_23867,N_23588);
xor U24849 (N_24849,N_23718,N_23240);
xnor U24850 (N_24850,N_23955,N_23536);
and U24851 (N_24851,N_23002,N_23946);
and U24852 (N_24852,N_23522,N_23210);
nand U24853 (N_24853,N_23847,N_23553);
and U24854 (N_24854,N_23087,N_23503);
nor U24855 (N_24855,N_23121,N_23533);
xnor U24856 (N_24856,N_23068,N_23944);
or U24857 (N_24857,N_23647,N_23210);
or U24858 (N_24858,N_23639,N_23793);
xnor U24859 (N_24859,N_23563,N_23236);
or U24860 (N_24860,N_23993,N_23306);
and U24861 (N_24861,N_23527,N_23613);
nand U24862 (N_24862,N_23136,N_23906);
xor U24863 (N_24863,N_23101,N_23450);
or U24864 (N_24864,N_23816,N_23271);
nor U24865 (N_24865,N_23469,N_23350);
nand U24866 (N_24866,N_23609,N_23944);
xor U24867 (N_24867,N_23064,N_23584);
xor U24868 (N_24868,N_23904,N_23511);
or U24869 (N_24869,N_23497,N_23097);
or U24870 (N_24870,N_23245,N_23564);
nor U24871 (N_24871,N_23035,N_23807);
nor U24872 (N_24872,N_23658,N_23051);
nand U24873 (N_24873,N_23906,N_23712);
nor U24874 (N_24874,N_23707,N_23185);
nor U24875 (N_24875,N_23182,N_23345);
nand U24876 (N_24876,N_23822,N_23625);
nor U24877 (N_24877,N_23275,N_23562);
xnor U24878 (N_24878,N_23819,N_23881);
or U24879 (N_24879,N_23535,N_23987);
or U24880 (N_24880,N_23617,N_23348);
and U24881 (N_24881,N_23194,N_23953);
and U24882 (N_24882,N_23820,N_23089);
or U24883 (N_24883,N_23752,N_23083);
nand U24884 (N_24884,N_23031,N_23049);
and U24885 (N_24885,N_23517,N_23321);
nor U24886 (N_24886,N_23935,N_23075);
or U24887 (N_24887,N_23988,N_23357);
and U24888 (N_24888,N_23180,N_23981);
and U24889 (N_24889,N_23147,N_23261);
and U24890 (N_24890,N_23846,N_23970);
or U24891 (N_24891,N_23196,N_23298);
xnor U24892 (N_24892,N_23410,N_23603);
nand U24893 (N_24893,N_23809,N_23142);
or U24894 (N_24894,N_23573,N_23178);
or U24895 (N_24895,N_23636,N_23829);
and U24896 (N_24896,N_23811,N_23878);
nand U24897 (N_24897,N_23008,N_23687);
and U24898 (N_24898,N_23818,N_23727);
and U24899 (N_24899,N_23371,N_23153);
and U24900 (N_24900,N_23624,N_23992);
nor U24901 (N_24901,N_23813,N_23399);
xor U24902 (N_24902,N_23296,N_23873);
nor U24903 (N_24903,N_23022,N_23549);
and U24904 (N_24904,N_23078,N_23863);
or U24905 (N_24905,N_23371,N_23981);
nor U24906 (N_24906,N_23152,N_23953);
or U24907 (N_24907,N_23832,N_23493);
xnor U24908 (N_24908,N_23013,N_23769);
nand U24909 (N_24909,N_23052,N_23259);
and U24910 (N_24910,N_23086,N_23271);
and U24911 (N_24911,N_23744,N_23443);
and U24912 (N_24912,N_23303,N_23709);
xnor U24913 (N_24913,N_23669,N_23842);
and U24914 (N_24914,N_23015,N_23768);
and U24915 (N_24915,N_23620,N_23198);
nor U24916 (N_24916,N_23262,N_23056);
xnor U24917 (N_24917,N_23612,N_23456);
nand U24918 (N_24918,N_23144,N_23875);
nor U24919 (N_24919,N_23832,N_23776);
or U24920 (N_24920,N_23402,N_23245);
nand U24921 (N_24921,N_23531,N_23928);
nand U24922 (N_24922,N_23579,N_23201);
nand U24923 (N_24923,N_23522,N_23022);
xor U24924 (N_24924,N_23365,N_23780);
xor U24925 (N_24925,N_23842,N_23292);
nor U24926 (N_24926,N_23280,N_23507);
nor U24927 (N_24927,N_23443,N_23235);
and U24928 (N_24928,N_23612,N_23044);
nand U24929 (N_24929,N_23240,N_23046);
nand U24930 (N_24930,N_23354,N_23461);
and U24931 (N_24931,N_23546,N_23255);
xnor U24932 (N_24932,N_23398,N_23671);
nand U24933 (N_24933,N_23390,N_23132);
xnor U24934 (N_24934,N_23395,N_23502);
or U24935 (N_24935,N_23150,N_23886);
or U24936 (N_24936,N_23936,N_23154);
and U24937 (N_24937,N_23811,N_23853);
or U24938 (N_24938,N_23362,N_23077);
or U24939 (N_24939,N_23099,N_23075);
and U24940 (N_24940,N_23953,N_23907);
nand U24941 (N_24941,N_23036,N_23293);
or U24942 (N_24942,N_23089,N_23393);
xnor U24943 (N_24943,N_23578,N_23992);
xnor U24944 (N_24944,N_23478,N_23643);
nand U24945 (N_24945,N_23324,N_23046);
xnor U24946 (N_24946,N_23537,N_23923);
xor U24947 (N_24947,N_23002,N_23561);
xor U24948 (N_24948,N_23387,N_23655);
nor U24949 (N_24949,N_23802,N_23283);
and U24950 (N_24950,N_23180,N_23006);
nand U24951 (N_24951,N_23423,N_23027);
or U24952 (N_24952,N_23502,N_23802);
xor U24953 (N_24953,N_23434,N_23106);
and U24954 (N_24954,N_23473,N_23189);
xnor U24955 (N_24955,N_23087,N_23114);
xor U24956 (N_24956,N_23553,N_23818);
and U24957 (N_24957,N_23375,N_23110);
or U24958 (N_24958,N_23366,N_23195);
nor U24959 (N_24959,N_23682,N_23609);
and U24960 (N_24960,N_23992,N_23302);
or U24961 (N_24961,N_23626,N_23263);
or U24962 (N_24962,N_23937,N_23244);
and U24963 (N_24963,N_23814,N_23308);
nand U24964 (N_24964,N_23208,N_23998);
nor U24965 (N_24965,N_23703,N_23406);
nand U24966 (N_24966,N_23510,N_23189);
and U24967 (N_24967,N_23613,N_23008);
nand U24968 (N_24968,N_23671,N_23445);
xor U24969 (N_24969,N_23871,N_23735);
and U24970 (N_24970,N_23986,N_23159);
or U24971 (N_24971,N_23466,N_23856);
xnor U24972 (N_24972,N_23384,N_23575);
or U24973 (N_24973,N_23107,N_23592);
nor U24974 (N_24974,N_23529,N_23611);
nor U24975 (N_24975,N_23437,N_23251);
nand U24976 (N_24976,N_23564,N_23652);
nand U24977 (N_24977,N_23573,N_23504);
nor U24978 (N_24978,N_23763,N_23195);
xnor U24979 (N_24979,N_23573,N_23929);
xor U24980 (N_24980,N_23560,N_23555);
xor U24981 (N_24981,N_23582,N_23291);
or U24982 (N_24982,N_23491,N_23814);
nand U24983 (N_24983,N_23536,N_23046);
xor U24984 (N_24984,N_23611,N_23704);
and U24985 (N_24985,N_23404,N_23184);
xnor U24986 (N_24986,N_23730,N_23151);
nor U24987 (N_24987,N_23714,N_23401);
nor U24988 (N_24988,N_23248,N_23240);
nor U24989 (N_24989,N_23587,N_23936);
xnor U24990 (N_24990,N_23179,N_23368);
and U24991 (N_24991,N_23221,N_23536);
or U24992 (N_24992,N_23687,N_23402);
xnor U24993 (N_24993,N_23791,N_23084);
nor U24994 (N_24994,N_23306,N_23538);
and U24995 (N_24995,N_23069,N_23456);
and U24996 (N_24996,N_23844,N_23695);
or U24997 (N_24997,N_23646,N_23466);
nand U24998 (N_24998,N_23440,N_23707);
or U24999 (N_24999,N_23174,N_23121);
and U25000 (N_25000,N_24410,N_24748);
and U25001 (N_25001,N_24957,N_24980);
and U25002 (N_25002,N_24134,N_24981);
xnor U25003 (N_25003,N_24488,N_24452);
and U25004 (N_25004,N_24683,N_24232);
and U25005 (N_25005,N_24689,N_24933);
xnor U25006 (N_25006,N_24456,N_24361);
nand U25007 (N_25007,N_24270,N_24719);
xor U25008 (N_25008,N_24946,N_24570);
xor U25009 (N_25009,N_24593,N_24994);
xor U25010 (N_25010,N_24846,N_24224);
nand U25011 (N_25011,N_24960,N_24945);
nor U25012 (N_25012,N_24419,N_24122);
nor U25013 (N_25013,N_24659,N_24422);
nor U25014 (N_25014,N_24901,N_24679);
or U25015 (N_25015,N_24813,N_24167);
and U25016 (N_25016,N_24790,N_24226);
xor U25017 (N_25017,N_24789,N_24268);
or U25018 (N_25018,N_24185,N_24557);
xor U25019 (N_25019,N_24269,N_24080);
nand U25020 (N_25020,N_24553,N_24250);
nor U25021 (N_25021,N_24105,N_24999);
nand U25022 (N_25022,N_24832,N_24070);
nand U25023 (N_25023,N_24707,N_24225);
or U25024 (N_25024,N_24931,N_24428);
nand U25025 (N_25025,N_24483,N_24735);
or U25026 (N_25026,N_24806,N_24145);
or U25027 (N_25027,N_24868,N_24401);
xor U25028 (N_25028,N_24702,N_24919);
xnor U25029 (N_25029,N_24510,N_24616);
and U25030 (N_25030,N_24026,N_24814);
nand U25031 (N_25031,N_24545,N_24035);
and U25032 (N_25032,N_24258,N_24711);
or U25033 (N_25033,N_24115,N_24217);
nand U25034 (N_25034,N_24387,N_24759);
xnor U25035 (N_25035,N_24163,N_24306);
or U25036 (N_25036,N_24620,N_24494);
or U25037 (N_25037,N_24643,N_24180);
and U25038 (N_25038,N_24514,N_24742);
nand U25039 (N_25039,N_24328,N_24988);
nand U25040 (N_25040,N_24463,N_24117);
or U25041 (N_25041,N_24773,N_24447);
or U25042 (N_25042,N_24388,N_24495);
nor U25043 (N_25043,N_24534,N_24146);
nand U25044 (N_25044,N_24920,N_24772);
and U25045 (N_25045,N_24639,N_24302);
and U25046 (N_25046,N_24943,N_24233);
and U25047 (N_25047,N_24331,N_24758);
xnor U25048 (N_25048,N_24648,N_24379);
nand U25049 (N_25049,N_24694,N_24985);
nand U25050 (N_25050,N_24755,N_24717);
and U25051 (N_25051,N_24910,N_24047);
and U25052 (N_25052,N_24631,N_24136);
nor U25053 (N_25053,N_24100,N_24952);
nand U25054 (N_25054,N_24573,N_24987);
nor U25055 (N_25055,N_24461,N_24768);
nand U25056 (N_25056,N_24611,N_24090);
nand U25057 (N_25057,N_24157,N_24671);
xnor U25058 (N_25058,N_24529,N_24692);
nand U25059 (N_25059,N_24609,N_24210);
or U25060 (N_25060,N_24374,N_24405);
and U25061 (N_25061,N_24155,N_24108);
xor U25062 (N_25062,N_24727,N_24237);
and U25063 (N_25063,N_24103,N_24182);
and U25064 (N_25064,N_24354,N_24785);
xor U25065 (N_25065,N_24754,N_24974);
nor U25066 (N_25066,N_24950,N_24552);
xor U25067 (N_25067,N_24441,N_24372);
nor U25068 (N_25068,N_24876,N_24211);
and U25069 (N_25069,N_24138,N_24203);
and U25070 (N_25070,N_24130,N_24420);
nand U25071 (N_25071,N_24497,N_24840);
or U25072 (N_25072,N_24932,N_24236);
or U25073 (N_25073,N_24997,N_24575);
xnor U25074 (N_25074,N_24953,N_24560);
xor U25075 (N_25075,N_24338,N_24290);
or U25076 (N_25076,N_24862,N_24831);
and U25077 (N_25077,N_24364,N_24585);
and U25078 (N_25078,N_24949,N_24436);
nand U25079 (N_25079,N_24907,N_24536);
and U25080 (N_25080,N_24209,N_24688);
or U25081 (N_25081,N_24594,N_24438);
xor U25082 (N_25082,N_24468,N_24809);
nor U25083 (N_25083,N_24606,N_24148);
nor U25084 (N_25084,N_24651,N_24263);
or U25085 (N_25085,N_24431,N_24549);
nand U25086 (N_25086,N_24044,N_24712);
and U25087 (N_25087,N_24822,N_24349);
and U25088 (N_25088,N_24486,N_24774);
nor U25089 (N_25089,N_24027,N_24474);
and U25090 (N_25090,N_24398,N_24296);
and U25091 (N_25091,N_24556,N_24693);
xnor U25092 (N_25092,N_24872,N_24308);
nor U25093 (N_25093,N_24903,N_24650);
xnor U25094 (N_25094,N_24778,N_24260);
or U25095 (N_25095,N_24409,N_24499);
and U25096 (N_25096,N_24665,N_24332);
xnor U25097 (N_25097,N_24445,N_24954);
or U25098 (N_25098,N_24111,N_24287);
or U25099 (N_25099,N_24925,N_24179);
nand U25100 (N_25100,N_24547,N_24595);
xor U25101 (N_25101,N_24627,N_24662);
and U25102 (N_25102,N_24731,N_24887);
xnor U25103 (N_25103,N_24640,N_24206);
xnor U25104 (N_25104,N_24292,N_24603);
or U25105 (N_25105,N_24764,N_24819);
or U25106 (N_25106,N_24176,N_24200);
and U25107 (N_25107,N_24393,N_24928);
xnor U25108 (N_25108,N_24187,N_24617);
xnor U25109 (N_25109,N_24976,N_24830);
xor U25110 (N_25110,N_24709,N_24346);
and U25111 (N_25111,N_24747,N_24125);
or U25112 (N_25112,N_24208,N_24112);
and U25113 (N_25113,N_24473,N_24891);
nor U25114 (N_25114,N_24934,N_24285);
xor U25115 (N_25115,N_24038,N_24500);
xor U25116 (N_25116,N_24291,N_24675);
xor U25117 (N_25117,N_24610,N_24921);
or U25118 (N_25118,N_24028,N_24131);
nor U25119 (N_25119,N_24343,N_24571);
and U25120 (N_25120,N_24626,N_24437);
nor U25121 (N_25121,N_24649,N_24561);
and U25122 (N_25122,N_24221,N_24266);
nor U25123 (N_25123,N_24995,N_24658);
nand U25124 (N_25124,N_24516,N_24905);
nor U25125 (N_25125,N_24858,N_24255);
and U25126 (N_25126,N_24466,N_24721);
nor U25127 (N_25127,N_24188,N_24339);
nor U25128 (N_25128,N_24760,N_24827);
or U25129 (N_25129,N_24215,N_24894);
or U25130 (N_25130,N_24723,N_24607);
nand U25131 (N_25131,N_24818,N_24798);
and U25132 (N_25132,N_24867,N_24329);
and U25133 (N_25133,N_24817,N_24579);
or U25134 (N_25134,N_24863,N_24548);
xnor U25135 (N_25135,N_24301,N_24893);
and U25136 (N_25136,N_24701,N_24158);
or U25137 (N_25137,N_24067,N_24278);
and U25138 (N_25138,N_24162,N_24964);
or U25139 (N_25139,N_24892,N_24020);
nor U25140 (N_25140,N_24257,N_24192);
or U25141 (N_25141,N_24634,N_24885);
or U25142 (N_25142,N_24961,N_24883);
and U25143 (N_25143,N_24000,N_24722);
or U25144 (N_25144,N_24505,N_24168);
xor U25145 (N_25145,N_24655,N_24150);
nand U25146 (N_25146,N_24889,N_24811);
xnor U25147 (N_25147,N_24312,N_24147);
nand U25148 (N_25148,N_24710,N_24776);
and U25149 (N_25149,N_24589,N_24929);
and U25150 (N_25150,N_24184,N_24309);
or U25151 (N_25151,N_24274,N_24788);
and U25152 (N_25152,N_24057,N_24775);
nand U25153 (N_25153,N_24771,N_24159);
nand U25154 (N_25154,N_24761,N_24153);
or U25155 (N_25155,N_24969,N_24890);
or U25156 (N_25156,N_24213,N_24056);
and U25157 (N_25157,N_24698,N_24395);
and U25158 (N_25158,N_24578,N_24060);
and U25159 (N_25159,N_24807,N_24016);
xor U25160 (N_25160,N_24491,N_24124);
xnor U25161 (N_25161,N_24815,N_24475);
and U25162 (N_25162,N_24795,N_24632);
and U25163 (N_25163,N_24726,N_24879);
nor U25164 (N_25164,N_24947,N_24356);
nor U25165 (N_25165,N_24657,N_24520);
and U25166 (N_25166,N_24336,N_24295);
and U25167 (N_25167,N_24528,N_24251);
and U25168 (N_25168,N_24597,N_24604);
and U25169 (N_25169,N_24962,N_24697);
nand U25170 (N_25170,N_24462,N_24245);
and U25171 (N_25171,N_24990,N_24622);
and U25172 (N_25172,N_24537,N_24254);
xor U25173 (N_25173,N_24527,N_24078);
or U25174 (N_25174,N_24927,N_24873);
and U25175 (N_25175,N_24440,N_24457);
nand U25176 (N_25176,N_24460,N_24975);
xor U25177 (N_25177,N_24915,N_24390);
nor U25178 (N_25178,N_24277,N_24635);
nor U25179 (N_25179,N_24851,N_24040);
nand U25180 (N_25180,N_24008,N_24244);
xnor U25181 (N_25181,N_24874,N_24479);
nor U25182 (N_25182,N_24212,N_24864);
nor U25183 (N_25183,N_24860,N_24304);
nand U25184 (N_25184,N_24142,N_24839);
and U25185 (N_25185,N_24967,N_24956);
and U25186 (N_25186,N_24050,N_24271);
nor U25187 (N_25187,N_24025,N_24470);
nand U25188 (N_25188,N_24471,N_24484);
and U25189 (N_25189,N_24538,N_24133);
and U25190 (N_25190,N_24317,N_24565);
or U25191 (N_25191,N_24123,N_24991);
nor U25192 (N_25192,N_24318,N_24355);
or U25193 (N_25193,N_24143,N_24544);
xnor U25194 (N_25194,N_24766,N_24160);
nor U25195 (N_25195,N_24299,N_24310);
xnor U25196 (N_25196,N_24704,N_24024);
nand U25197 (N_25197,N_24902,N_24888);
nand U25198 (N_25198,N_24046,N_24077);
xor U25199 (N_25199,N_24417,N_24496);
nor U25200 (N_25200,N_24850,N_24684);
and U25201 (N_25201,N_24191,N_24881);
or U25202 (N_25202,N_24998,N_24079);
nand U25203 (N_25203,N_24403,N_24577);
and U25204 (N_25204,N_24321,N_24563);
nand U25205 (N_25205,N_24786,N_24204);
nor U25206 (N_25206,N_24909,N_24531);
xor U25207 (N_25207,N_24175,N_24453);
nand U25208 (N_25208,N_24653,N_24939);
nand U25209 (N_25209,N_24829,N_24968);
or U25210 (N_25210,N_24645,N_24414);
nand U25211 (N_25211,N_24068,N_24564);
or U25212 (N_25212,N_24367,N_24061);
xor U25213 (N_25213,N_24094,N_24502);
and U25214 (N_25214,N_24524,N_24242);
or U25215 (N_25215,N_24661,N_24847);
nand U25216 (N_25216,N_24912,N_24582);
or U25217 (N_25217,N_24033,N_24246);
or U25218 (N_25218,N_24663,N_24938);
or U25219 (N_25219,N_24132,N_24039);
nor U25220 (N_25220,N_24983,N_24518);
or U25221 (N_25221,N_24107,N_24218);
xnor U25222 (N_25222,N_24015,N_24848);
xor U25223 (N_25223,N_24880,N_24247);
xor U25224 (N_25224,N_24982,N_24335);
nor U25225 (N_25225,N_24127,N_24114);
xnor U25226 (N_25226,N_24362,N_24637);
nor U25227 (N_25227,N_24451,N_24342);
nor U25228 (N_25228,N_24053,N_24030);
nor U25229 (N_25229,N_24161,N_24439);
nor U25230 (N_25230,N_24426,N_24333);
or U25231 (N_25231,N_24828,N_24793);
or U25232 (N_25232,N_24316,N_24170);
xor U25233 (N_25233,N_24716,N_24120);
nand U25234 (N_25234,N_24618,N_24383);
and U25235 (N_25235,N_24699,N_24836);
nor U25236 (N_25236,N_24678,N_24360);
nand U25237 (N_25237,N_24849,N_24190);
nor U25238 (N_25238,N_24703,N_24546);
nand U25239 (N_25239,N_24743,N_24313);
nor U25240 (N_25240,N_24326,N_24744);
xnor U25241 (N_25241,N_24104,N_24235);
and U25242 (N_25242,N_24402,N_24581);
xnor U25243 (N_25243,N_24444,N_24216);
or U25244 (N_25244,N_24081,N_24871);
or U25245 (N_25245,N_24116,N_24930);
or U25246 (N_25246,N_24171,N_24083);
xnor U25247 (N_25247,N_24085,N_24695);
and U25248 (N_25248,N_24427,N_24799);
or U25249 (N_25249,N_24911,N_24823);
and U25250 (N_25250,N_24002,N_24353);
xnor U25251 (N_25251,N_24740,N_24532);
nor U25252 (N_25252,N_24430,N_24064);
nand U25253 (N_25253,N_24913,N_24877);
xor U25254 (N_25254,N_24381,N_24051);
and U25255 (N_25255,N_24262,N_24177);
xor U25256 (N_25256,N_24400,N_24164);
xnor U25257 (N_25257,N_24222,N_24530);
xor U25258 (N_25258,N_24992,N_24612);
xnor U25259 (N_25259,N_24614,N_24073);
and U25260 (N_25260,N_24673,N_24899);
and U25261 (N_25261,N_24917,N_24680);
or U25262 (N_25262,N_24037,N_24259);
or U25263 (N_25263,N_24782,N_24023);
or U25264 (N_25264,N_24455,N_24842);
xnor U25265 (N_25265,N_24566,N_24895);
xor U25266 (N_25266,N_24487,N_24587);
and U25267 (N_25267,N_24567,N_24307);
or U25268 (N_25268,N_24202,N_24784);
nand U25269 (N_25269,N_24368,N_24825);
or U25270 (N_25270,N_24623,N_24800);
xor U25271 (N_25271,N_24063,N_24031);
xor U25272 (N_25272,N_24109,N_24667);
nor U25273 (N_25273,N_24739,N_24730);
xor U25274 (N_25274,N_24074,N_24359);
and U25275 (N_25275,N_24629,N_24865);
and U25276 (N_25276,N_24265,N_24979);
and U25277 (N_25277,N_24152,N_24756);
nand U25278 (N_25278,N_24093,N_24059);
and U25279 (N_25279,N_24151,N_24713);
nor U25280 (N_25280,N_24465,N_24344);
and U25281 (N_25281,N_24696,N_24173);
and U25282 (N_25282,N_24660,N_24904);
nand U25283 (N_25283,N_24805,N_24686);
nand U25284 (N_25284,N_24812,N_24166);
nor U25285 (N_25285,N_24273,N_24036);
or U25286 (N_25286,N_24382,N_24554);
nor U25287 (N_25287,N_24485,N_24195);
nor U25288 (N_25288,N_24870,N_24392);
nand U25289 (N_25289,N_24602,N_24559);
or U25290 (N_25290,N_24320,N_24019);
xor U25291 (N_25291,N_24220,N_24408);
nand U25292 (N_25292,N_24972,N_24196);
nand U25293 (N_25293,N_24097,N_24810);
nor U25294 (N_25294,N_24407,N_24646);
xor U25295 (N_25295,N_24178,N_24095);
or U25296 (N_25296,N_24522,N_24376);
xnor U25297 (N_25297,N_24551,N_24797);
nor U25298 (N_25298,N_24685,N_24238);
nand U25299 (N_25299,N_24241,N_24069);
or U25300 (N_25300,N_24370,N_24350);
or U25301 (N_25301,N_24275,N_24165);
nor U25302 (N_25302,N_24239,N_24540);
and U25303 (N_25303,N_24248,N_24323);
nand U25304 (N_25304,N_24749,N_24838);
or U25305 (N_25305,N_24855,N_24896);
xnor U25306 (N_25306,N_24391,N_24866);
xnor U25307 (N_25307,N_24448,N_24550);
xor U25308 (N_25308,N_24796,N_24129);
or U25309 (N_25309,N_24140,N_24777);
nand U25310 (N_25310,N_24543,N_24613);
nor U25311 (N_25311,N_24319,N_24062);
or U25312 (N_25312,N_24358,N_24802);
nand U25313 (N_25313,N_24459,N_24449);
nor U25314 (N_25314,N_24337,N_24942);
nor U25315 (N_25315,N_24517,N_24853);
xnor U25316 (N_25316,N_24845,N_24854);
xnor U25317 (N_25317,N_24615,N_24936);
and U25318 (N_25318,N_24377,N_24276);
nand U25319 (N_25319,N_24197,N_24415);
nor U25320 (N_25320,N_24482,N_24480);
xor U25321 (N_25321,N_24837,N_24986);
xnor U25322 (N_25322,N_24397,N_24674);
nand U25323 (N_25323,N_24590,N_24334);
nor U25324 (N_25324,N_24186,N_24608);
nor U25325 (N_25325,N_24619,N_24508);
xnor U25326 (N_25326,N_24965,N_24113);
and U25327 (N_25327,N_24708,N_24562);
or U25328 (N_25328,N_24154,N_24670);
xnor U25329 (N_25329,N_24071,N_24458);
nor U25330 (N_25330,N_24843,N_24194);
or U25331 (N_25331,N_24808,N_24207);
nor U25332 (N_25332,N_24264,N_24737);
or U25333 (N_25333,N_24384,N_24054);
nand U25334 (N_25334,N_24523,N_24385);
and U25335 (N_25335,N_24283,N_24511);
nor U25336 (N_25336,N_24017,N_24325);
or U25337 (N_25337,N_24820,N_24745);
or U25338 (N_25338,N_24007,N_24753);
xor U25339 (N_25339,N_24884,N_24642);
or U25340 (N_25340,N_24021,N_24803);
nor U25341 (N_25341,N_24924,N_24230);
nor U25342 (N_25342,N_24507,N_24014);
and U25343 (N_25343,N_24380,N_24013);
or U25344 (N_25344,N_24375,N_24289);
and U25345 (N_25345,N_24418,N_24664);
nor U25346 (N_25346,N_24844,N_24412);
or U25347 (N_25347,N_24741,N_24984);
nand U25348 (N_25348,N_24135,N_24914);
or U25349 (N_25349,N_24009,N_24141);
or U25350 (N_25350,N_24003,N_24169);
and U25351 (N_25351,N_24625,N_24916);
nor U25352 (N_25352,N_24783,N_24801);
nand U25353 (N_25353,N_24413,N_24373);
nand U25354 (N_25354,N_24096,N_24584);
nor U25355 (N_25355,N_24322,N_24092);
xnor U25356 (N_25356,N_24004,N_24751);
and U25357 (N_25357,N_24477,N_24476);
and U25358 (N_25358,N_24857,N_24729);
or U25359 (N_25359,N_24029,N_24227);
nor U25360 (N_25360,N_24298,N_24311);
or U25361 (N_25361,N_24791,N_24824);
nor U25362 (N_25362,N_24034,N_24351);
nand U25363 (N_25363,N_24001,N_24330);
or U25364 (N_25364,N_24011,N_24205);
nand U25365 (N_25365,N_24706,N_24432);
or U25366 (N_25366,N_24416,N_24568);
xnor U25367 (N_25367,N_24596,N_24324);
or U25368 (N_25368,N_24705,N_24633);
or U25369 (N_25369,N_24055,N_24253);
and U25370 (N_25370,N_24315,N_24087);
nor U25371 (N_25371,N_24971,N_24586);
nand U25372 (N_25372,N_24293,N_24628);
or U25373 (N_25373,N_24442,N_24279);
nor U25374 (N_25374,N_24424,N_24781);
or U25375 (N_25375,N_24940,N_24724);
xor U25376 (N_25376,N_24833,N_24792);
xnor U25377 (N_25377,N_24601,N_24119);
nor U25378 (N_25378,N_24834,N_24411);
nor U25379 (N_25379,N_24365,N_24763);
or U25380 (N_25380,N_24089,N_24045);
nor U25381 (N_25381,N_24647,N_24010);
or U25382 (N_25382,N_24533,N_24826);
and U25383 (N_25383,N_24509,N_24937);
nand U25384 (N_25384,N_24583,N_24005);
nor U25385 (N_25385,N_24535,N_24728);
xnor U25386 (N_25386,N_24340,N_24048);
nor U25387 (N_25387,N_24977,N_24072);
xor U25388 (N_25388,N_24435,N_24454);
or U25389 (N_25389,N_24525,N_24174);
or U25390 (N_25390,N_24765,N_24720);
xor U25391 (N_25391,N_24908,N_24327);
or U25392 (N_25392,N_24715,N_24128);
nor U25393 (N_25393,N_24082,N_24654);
nor U25394 (N_25394,N_24841,N_24926);
nor U25395 (N_25395,N_24521,N_24746);
xor U25396 (N_25396,N_24032,N_24006);
nand U25397 (N_25397,N_24139,N_24280);
and U25398 (N_25398,N_24288,N_24624);
xnor U25399 (N_25399,N_24598,N_24922);
and U25400 (N_25400,N_24856,N_24600);
and U25401 (N_25401,N_24102,N_24861);
nand U25402 (N_25402,N_24043,N_24366);
or U25403 (N_25403,N_24869,N_24098);
and U25404 (N_25404,N_24446,N_24515);
nor U25405 (N_25405,N_24252,N_24691);
nand U25406 (N_25406,N_24978,N_24429);
nand U25407 (N_25407,N_24574,N_24588);
nor U25408 (N_25408,N_24106,N_24406);
and U25409 (N_25409,N_24101,N_24681);
nand U25410 (N_25410,N_24677,N_24394);
and U25411 (N_25411,N_24404,N_24223);
nand U25412 (N_25412,N_24668,N_24580);
and U25413 (N_25413,N_24638,N_24464);
and U25414 (N_25414,N_24666,N_24732);
nand U25415 (N_25415,N_24725,N_24513);
nand U25416 (N_25416,N_24541,N_24989);
nor U25417 (N_25417,N_24240,N_24300);
or U25418 (N_25418,N_24519,N_24878);
nand U25419 (N_25419,N_24490,N_24423);
and U25420 (N_25420,N_24183,N_24886);
nor U25421 (N_25421,N_24088,N_24099);
nand U25422 (N_25422,N_24970,N_24075);
nor U25423 (N_25423,N_24882,N_24201);
nand U25424 (N_25424,N_24700,N_24126);
or U25425 (N_25425,N_24012,N_24229);
xor U25426 (N_25426,N_24630,N_24555);
nand U25427 (N_25427,N_24172,N_24363);
nand U25428 (N_25428,N_24121,N_24501);
nand U25429 (N_25429,N_24231,N_24804);
nor U25430 (N_25430,N_24018,N_24752);
nor U25431 (N_25431,N_24303,N_24656);
and U25432 (N_25432,N_24219,N_24421);
nor U25433 (N_25433,N_24049,N_24714);
nor U25434 (N_25434,N_24558,N_24503);
xnor U25435 (N_25435,N_24996,N_24498);
nor U25436 (N_25436,N_24993,N_24973);
and U25437 (N_25437,N_24935,N_24314);
or U25438 (N_25438,N_24347,N_24644);
and U25439 (N_25439,N_24542,N_24757);
or U25440 (N_25440,N_24481,N_24425);
or U25441 (N_25441,N_24676,N_24592);
nor U25442 (N_25442,N_24512,N_24348);
and U25443 (N_25443,N_24572,N_24794);
nor U25444 (N_25444,N_24076,N_24493);
nand U25445 (N_25445,N_24690,N_24652);
xnor U25446 (N_25446,N_24599,N_24767);
or U25447 (N_25447,N_24282,N_24469);
and U25448 (N_25448,N_24389,N_24816);
nand U25449 (N_25449,N_24506,N_24958);
xnor U25450 (N_25450,N_24305,N_24399);
nand U25451 (N_25451,N_24450,N_24770);
nand U25452 (N_25452,N_24576,N_24504);
xnor U25453 (N_25453,N_24762,N_24284);
xor U25454 (N_25454,N_24966,N_24738);
nand U25455 (N_25455,N_24897,N_24058);
nand U25456 (N_25456,N_24687,N_24272);
xnor U25457 (N_25457,N_24489,N_24636);
or U25458 (N_25458,N_24341,N_24234);
and U25459 (N_25459,N_24137,N_24780);
nor U25460 (N_25460,N_24352,N_24526);
or U25461 (N_25461,N_24492,N_24900);
xnor U25462 (N_25462,N_24569,N_24261);
xor U25463 (N_25463,N_24951,N_24297);
or U25464 (N_25464,N_24199,N_24941);
or U25465 (N_25465,N_24256,N_24906);
and U25466 (N_25466,N_24682,N_24859);
or U25467 (N_25467,N_24243,N_24378);
nor U25468 (N_25468,N_24286,N_24472);
nand U25469 (N_25469,N_24065,N_24787);
xnor U25470 (N_25470,N_24267,N_24641);
nand U25471 (N_25471,N_24091,N_24779);
nand U25472 (N_25472,N_24669,N_24734);
nor U25473 (N_25473,N_24443,N_24041);
and U25474 (N_25474,N_24852,N_24156);
nor U25475 (N_25475,N_24959,N_24345);
nand U25476 (N_25476,N_24621,N_24042);
nor U25477 (N_25477,N_24249,N_24718);
xnor U25478 (N_25478,N_24066,N_24821);
nor U25479 (N_25479,N_24022,N_24478);
xor U25480 (N_25480,N_24371,N_24433);
nor U25481 (N_25481,N_24434,N_24357);
nand U25482 (N_25482,N_24605,N_24144);
nand U25483 (N_25483,N_24294,N_24052);
nand U25484 (N_25484,N_24948,N_24228);
nor U25485 (N_25485,N_24149,N_24539);
and U25486 (N_25486,N_24963,N_24118);
and U25487 (N_25487,N_24955,N_24591);
or U25488 (N_25488,N_24110,N_24875);
nor U25489 (N_25489,N_24084,N_24750);
or U25490 (N_25490,N_24672,N_24898);
or U25491 (N_25491,N_24369,N_24733);
xor U25492 (N_25492,N_24193,N_24467);
and U25493 (N_25493,N_24214,N_24736);
and U25494 (N_25494,N_24086,N_24769);
or U25495 (N_25495,N_24944,N_24189);
or U25496 (N_25496,N_24181,N_24923);
xnor U25497 (N_25497,N_24835,N_24918);
nand U25498 (N_25498,N_24396,N_24386);
or U25499 (N_25499,N_24281,N_24198);
xnor U25500 (N_25500,N_24961,N_24420);
xor U25501 (N_25501,N_24767,N_24131);
xor U25502 (N_25502,N_24030,N_24556);
nor U25503 (N_25503,N_24808,N_24463);
nand U25504 (N_25504,N_24693,N_24284);
nor U25505 (N_25505,N_24938,N_24011);
nand U25506 (N_25506,N_24577,N_24534);
and U25507 (N_25507,N_24084,N_24949);
or U25508 (N_25508,N_24046,N_24114);
and U25509 (N_25509,N_24311,N_24494);
or U25510 (N_25510,N_24335,N_24886);
nor U25511 (N_25511,N_24565,N_24361);
nand U25512 (N_25512,N_24008,N_24510);
and U25513 (N_25513,N_24339,N_24553);
nand U25514 (N_25514,N_24004,N_24834);
or U25515 (N_25515,N_24177,N_24203);
nand U25516 (N_25516,N_24338,N_24208);
or U25517 (N_25517,N_24369,N_24855);
nand U25518 (N_25518,N_24333,N_24462);
and U25519 (N_25519,N_24800,N_24685);
and U25520 (N_25520,N_24655,N_24260);
xnor U25521 (N_25521,N_24827,N_24415);
and U25522 (N_25522,N_24908,N_24637);
or U25523 (N_25523,N_24715,N_24042);
or U25524 (N_25524,N_24251,N_24006);
and U25525 (N_25525,N_24442,N_24718);
xor U25526 (N_25526,N_24722,N_24570);
or U25527 (N_25527,N_24574,N_24110);
nor U25528 (N_25528,N_24839,N_24118);
or U25529 (N_25529,N_24028,N_24467);
nor U25530 (N_25530,N_24731,N_24236);
xor U25531 (N_25531,N_24609,N_24930);
xnor U25532 (N_25532,N_24478,N_24832);
or U25533 (N_25533,N_24528,N_24797);
nand U25534 (N_25534,N_24364,N_24420);
and U25535 (N_25535,N_24565,N_24991);
xor U25536 (N_25536,N_24752,N_24755);
nand U25537 (N_25537,N_24193,N_24659);
and U25538 (N_25538,N_24663,N_24847);
nor U25539 (N_25539,N_24459,N_24794);
nand U25540 (N_25540,N_24061,N_24809);
xor U25541 (N_25541,N_24873,N_24662);
and U25542 (N_25542,N_24664,N_24872);
and U25543 (N_25543,N_24135,N_24318);
nor U25544 (N_25544,N_24791,N_24997);
or U25545 (N_25545,N_24666,N_24328);
or U25546 (N_25546,N_24341,N_24285);
xnor U25547 (N_25547,N_24102,N_24209);
xor U25548 (N_25548,N_24252,N_24626);
nor U25549 (N_25549,N_24737,N_24405);
or U25550 (N_25550,N_24811,N_24980);
nor U25551 (N_25551,N_24653,N_24193);
and U25552 (N_25552,N_24638,N_24811);
or U25553 (N_25553,N_24232,N_24541);
nor U25554 (N_25554,N_24838,N_24348);
nor U25555 (N_25555,N_24359,N_24796);
and U25556 (N_25556,N_24975,N_24448);
or U25557 (N_25557,N_24665,N_24888);
xnor U25558 (N_25558,N_24795,N_24749);
or U25559 (N_25559,N_24101,N_24910);
and U25560 (N_25560,N_24604,N_24504);
nand U25561 (N_25561,N_24189,N_24415);
and U25562 (N_25562,N_24361,N_24161);
nor U25563 (N_25563,N_24434,N_24539);
nand U25564 (N_25564,N_24709,N_24843);
nor U25565 (N_25565,N_24074,N_24621);
and U25566 (N_25566,N_24068,N_24205);
nand U25567 (N_25567,N_24207,N_24270);
and U25568 (N_25568,N_24551,N_24341);
nor U25569 (N_25569,N_24583,N_24007);
or U25570 (N_25570,N_24093,N_24096);
nor U25571 (N_25571,N_24033,N_24105);
or U25572 (N_25572,N_24271,N_24013);
nand U25573 (N_25573,N_24155,N_24017);
xnor U25574 (N_25574,N_24426,N_24607);
xor U25575 (N_25575,N_24267,N_24753);
nand U25576 (N_25576,N_24239,N_24476);
xnor U25577 (N_25577,N_24856,N_24830);
or U25578 (N_25578,N_24001,N_24663);
nand U25579 (N_25579,N_24290,N_24981);
xor U25580 (N_25580,N_24853,N_24297);
xnor U25581 (N_25581,N_24503,N_24921);
xnor U25582 (N_25582,N_24991,N_24828);
nand U25583 (N_25583,N_24416,N_24399);
nand U25584 (N_25584,N_24388,N_24329);
xor U25585 (N_25585,N_24475,N_24643);
or U25586 (N_25586,N_24437,N_24623);
nor U25587 (N_25587,N_24944,N_24793);
or U25588 (N_25588,N_24345,N_24428);
or U25589 (N_25589,N_24364,N_24306);
and U25590 (N_25590,N_24069,N_24838);
nor U25591 (N_25591,N_24576,N_24573);
nand U25592 (N_25592,N_24723,N_24411);
or U25593 (N_25593,N_24619,N_24615);
and U25594 (N_25594,N_24004,N_24316);
nand U25595 (N_25595,N_24089,N_24821);
or U25596 (N_25596,N_24312,N_24943);
xor U25597 (N_25597,N_24025,N_24244);
nor U25598 (N_25598,N_24523,N_24205);
xor U25599 (N_25599,N_24788,N_24618);
xnor U25600 (N_25600,N_24954,N_24828);
and U25601 (N_25601,N_24454,N_24548);
xnor U25602 (N_25602,N_24151,N_24351);
and U25603 (N_25603,N_24377,N_24037);
or U25604 (N_25604,N_24362,N_24872);
or U25605 (N_25605,N_24521,N_24563);
and U25606 (N_25606,N_24385,N_24666);
or U25607 (N_25607,N_24669,N_24525);
xor U25608 (N_25608,N_24445,N_24057);
nand U25609 (N_25609,N_24219,N_24593);
or U25610 (N_25610,N_24969,N_24796);
xor U25611 (N_25611,N_24936,N_24748);
or U25612 (N_25612,N_24218,N_24321);
nand U25613 (N_25613,N_24261,N_24637);
or U25614 (N_25614,N_24362,N_24656);
and U25615 (N_25615,N_24330,N_24129);
or U25616 (N_25616,N_24222,N_24433);
and U25617 (N_25617,N_24756,N_24029);
xnor U25618 (N_25618,N_24815,N_24891);
or U25619 (N_25619,N_24620,N_24562);
xor U25620 (N_25620,N_24924,N_24455);
xnor U25621 (N_25621,N_24109,N_24039);
and U25622 (N_25622,N_24827,N_24704);
or U25623 (N_25623,N_24488,N_24214);
or U25624 (N_25624,N_24713,N_24426);
or U25625 (N_25625,N_24133,N_24686);
nor U25626 (N_25626,N_24280,N_24608);
and U25627 (N_25627,N_24473,N_24985);
xor U25628 (N_25628,N_24744,N_24880);
or U25629 (N_25629,N_24978,N_24500);
xor U25630 (N_25630,N_24298,N_24554);
xnor U25631 (N_25631,N_24855,N_24337);
nand U25632 (N_25632,N_24110,N_24254);
nor U25633 (N_25633,N_24897,N_24274);
and U25634 (N_25634,N_24929,N_24012);
and U25635 (N_25635,N_24640,N_24290);
nand U25636 (N_25636,N_24944,N_24429);
nand U25637 (N_25637,N_24750,N_24814);
or U25638 (N_25638,N_24239,N_24454);
nor U25639 (N_25639,N_24497,N_24338);
nand U25640 (N_25640,N_24971,N_24413);
nand U25641 (N_25641,N_24944,N_24250);
nor U25642 (N_25642,N_24035,N_24832);
nand U25643 (N_25643,N_24824,N_24596);
xnor U25644 (N_25644,N_24965,N_24976);
nand U25645 (N_25645,N_24324,N_24858);
xnor U25646 (N_25646,N_24309,N_24316);
xnor U25647 (N_25647,N_24472,N_24966);
xor U25648 (N_25648,N_24321,N_24969);
and U25649 (N_25649,N_24638,N_24788);
xnor U25650 (N_25650,N_24661,N_24698);
and U25651 (N_25651,N_24667,N_24657);
nor U25652 (N_25652,N_24725,N_24585);
nor U25653 (N_25653,N_24386,N_24125);
nand U25654 (N_25654,N_24562,N_24062);
nand U25655 (N_25655,N_24226,N_24762);
or U25656 (N_25656,N_24235,N_24971);
nor U25657 (N_25657,N_24019,N_24041);
and U25658 (N_25658,N_24802,N_24246);
nand U25659 (N_25659,N_24782,N_24804);
and U25660 (N_25660,N_24362,N_24897);
xor U25661 (N_25661,N_24108,N_24096);
nand U25662 (N_25662,N_24449,N_24856);
nand U25663 (N_25663,N_24694,N_24117);
nor U25664 (N_25664,N_24901,N_24975);
and U25665 (N_25665,N_24367,N_24910);
nand U25666 (N_25666,N_24025,N_24727);
or U25667 (N_25667,N_24469,N_24742);
and U25668 (N_25668,N_24638,N_24872);
xnor U25669 (N_25669,N_24186,N_24431);
xor U25670 (N_25670,N_24232,N_24441);
nor U25671 (N_25671,N_24004,N_24781);
or U25672 (N_25672,N_24713,N_24201);
xnor U25673 (N_25673,N_24855,N_24404);
xor U25674 (N_25674,N_24424,N_24120);
and U25675 (N_25675,N_24596,N_24162);
and U25676 (N_25676,N_24471,N_24669);
xnor U25677 (N_25677,N_24353,N_24695);
or U25678 (N_25678,N_24234,N_24546);
nor U25679 (N_25679,N_24899,N_24997);
or U25680 (N_25680,N_24206,N_24334);
nor U25681 (N_25681,N_24112,N_24430);
nor U25682 (N_25682,N_24884,N_24741);
nor U25683 (N_25683,N_24624,N_24332);
nand U25684 (N_25684,N_24284,N_24273);
nand U25685 (N_25685,N_24332,N_24364);
xnor U25686 (N_25686,N_24043,N_24515);
nand U25687 (N_25687,N_24124,N_24817);
nor U25688 (N_25688,N_24185,N_24478);
xor U25689 (N_25689,N_24254,N_24932);
xnor U25690 (N_25690,N_24191,N_24219);
nor U25691 (N_25691,N_24495,N_24556);
or U25692 (N_25692,N_24951,N_24254);
or U25693 (N_25693,N_24467,N_24685);
nor U25694 (N_25694,N_24281,N_24894);
nand U25695 (N_25695,N_24307,N_24152);
nand U25696 (N_25696,N_24530,N_24425);
and U25697 (N_25697,N_24279,N_24609);
xor U25698 (N_25698,N_24793,N_24015);
or U25699 (N_25699,N_24068,N_24256);
or U25700 (N_25700,N_24095,N_24511);
or U25701 (N_25701,N_24250,N_24924);
nand U25702 (N_25702,N_24271,N_24798);
xor U25703 (N_25703,N_24220,N_24913);
and U25704 (N_25704,N_24226,N_24701);
nor U25705 (N_25705,N_24948,N_24784);
xor U25706 (N_25706,N_24642,N_24790);
xor U25707 (N_25707,N_24849,N_24214);
xor U25708 (N_25708,N_24015,N_24218);
nor U25709 (N_25709,N_24521,N_24904);
nand U25710 (N_25710,N_24069,N_24763);
nand U25711 (N_25711,N_24839,N_24691);
nor U25712 (N_25712,N_24543,N_24366);
or U25713 (N_25713,N_24475,N_24692);
xnor U25714 (N_25714,N_24649,N_24311);
or U25715 (N_25715,N_24664,N_24796);
xor U25716 (N_25716,N_24779,N_24848);
nor U25717 (N_25717,N_24247,N_24930);
nor U25718 (N_25718,N_24501,N_24747);
nand U25719 (N_25719,N_24196,N_24347);
nor U25720 (N_25720,N_24070,N_24114);
and U25721 (N_25721,N_24304,N_24873);
and U25722 (N_25722,N_24428,N_24794);
nand U25723 (N_25723,N_24358,N_24795);
or U25724 (N_25724,N_24629,N_24610);
and U25725 (N_25725,N_24976,N_24714);
xnor U25726 (N_25726,N_24293,N_24567);
nand U25727 (N_25727,N_24085,N_24070);
nand U25728 (N_25728,N_24030,N_24698);
nand U25729 (N_25729,N_24819,N_24265);
nor U25730 (N_25730,N_24117,N_24809);
or U25731 (N_25731,N_24322,N_24467);
nor U25732 (N_25732,N_24611,N_24935);
or U25733 (N_25733,N_24575,N_24872);
or U25734 (N_25734,N_24832,N_24334);
nor U25735 (N_25735,N_24493,N_24548);
or U25736 (N_25736,N_24219,N_24962);
nor U25737 (N_25737,N_24438,N_24504);
nor U25738 (N_25738,N_24523,N_24952);
and U25739 (N_25739,N_24741,N_24090);
nand U25740 (N_25740,N_24556,N_24161);
and U25741 (N_25741,N_24332,N_24940);
nor U25742 (N_25742,N_24401,N_24727);
or U25743 (N_25743,N_24665,N_24477);
and U25744 (N_25744,N_24250,N_24479);
nand U25745 (N_25745,N_24509,N_24600);
xnor U25746 (N_25746,N_24710,N_24972);
nand U25747 (N_25747,N_24253,N_24960);
and U25748 (N_25748,N_24478,N_24647);
nand U25749 (N_25749,N_24325,N_24158);
nor U25750 (N_25750,N_24861,N_24849);
xor U25751 (N_25751,N_24643,N_24121);
nor U25752 (N_25752,N_24161,N_24055);
or U25753 (N_25753,N_24501,N_24114);
nor U25754 (N_25754,N_24727,N_24815);
and U25755 (N_25755,N_24256,N_24742);
and U25756 (N_25756,N_24434,N_24611);
nand U25757 (N_25757,N_24346,N_24356);
xor U25758 (N_25758,N_24182,N_24010);
nand U25759 (N_25759,N_24015,N_24201);
nor U25760 (N_25760,N_24869,N_24873);
or U25761 (N_25761,N_24757,N_24986);
nor U25762 (N_25762,N_24414,N_24663);
or U25763 (N_25763,N_24197,N_24800);
nand U25764 (N_25764,N_24162,N_24986);
nand U25765 (N_25765,N_24195,N_24331);
and U25766 (N_25766,N_24103,N_24377);
nand U25767 (N_25767,N_24192,N_24073);
nor U25768 (N_25768,N_24716,N_24202);
and U25769 (N_25769,N_24738,N_24817);
nor U25770 (N_25770,N_24630,N_24997);
or U25771 (N_25771,N_24240,N_24457);
xor U25772 (N_25772,N_24627,N_24262);
and U25773 (N_25773,N_24916,N_24859);
nor U25774 (N_25774,N_24653,N_24801);
xnor U25775 (N_25775,N_24079,N_24646);
and U25776 (N_25776,N_24949,N_24237);
nor U25777 (N_25777,N_24410,N_24458);
nand U25778 (N_25778,N_24336,N_24025);
nor U25779 (N_25779,N_24820,N_24972);
xor U25780 (N_25780,N_24273,N_24304);
nand U25781 (N_25781,N_24934,N_24831);
nor U25782 (N_25782,N_24081,N_24763);
nor U25783 (N_25783,N_24115,N_24041);
and U25784 (N_25784,N_24979,N_24021);
nor U25785 (N_25785,N_24998,N_24464);
nor U25786 (N_25786,N_24160,N_24427);
and U25787 (N_25787,N_24911,N_24182);
or U25788 (N_25788,N_24743,N_24208);
nor U25789 (N_25789,N_24970,N_24137);
and U25790 (N_25790,N_24527,N_24576);
nand U25791 (N_25791,N_24049,N_24942);
and U25792 (N_25792,N_24147,N_24887);
xnor U25793 (N_25793,N_24078,N_24571);
xor U25794 (N_25794,N_24459,N_24792);
or U25795 (N_25795,N_24449,N_24987);
or U25796 (N_25796,N_24620,N_24356);
nor U25797 (N_25797,N_24345,N_24065);
nand U25798 (N_25798,N_24033,N_24560);
nand U25799 (N_25799,N_24005,N_24353);
xor U25800 (N_25800,N_24515,N_24881);
and U25801 (N_25801,N_24279,N_24942);
nand U25802 (N_25802,N_24089,N_24327);
and U25803 (N_25803,N_24070,N_24947);
nand U25804 (N_25804,N_24511,N_24518);
nor U25805 (N_25805,N_24699,N_24667);
or U25806 (N_25806,N_24538,N_24563);
nand U25807 (N_25807,N_24170,N_24761);
and U25808 (N_25808,N_24297,N_24516);
nor U25809 (N_25809,N_24364,N_24500);
or U25810 (N_25810,N_24604,N_24755);
or U25811 (N_25811,N_24473,N_24509);
nor U25812 (N_25812,N_24047,N_24280);
or U25813 (N_25813,N_24822,N_24962);
or U25814 (N_25814,N_24993,N_24365);
xnor U25815 (N_25815,N_24854,N_24490);
nor U25816 (N_25816,N_24314,N_24005);
and U25817 (N_25817,N_24523,N_24927);
nand U25818 (N_25818,N_24461,N_24247);
nor U25819 (N_25819,N_24691,N_24433);
or U25820 (N_25820,N_24177,N_24619);
nand U25821 (N_25821,N_24911,N_24249);
and U25822 (N_25822,N_24304,N_24926);
or U25823 (N_25823,N_24115,N_24564);
nand U25824 (N_25824,N_24832,N_24275);
nand U25825 (N_25825,N_24170,N_24860);
nor U25826 (N_25826,N_24018,N_24379);
and U25827 (N_25827,N_24546,N_24938);
nand U25828 (N_25828,N_24491,N_24628);
xor U25829 (N_25829,N_24609,N_24415);
nand U25830 (N_25830,N_24200,N_24007);
nand U25831 (N_25831,N_24210,N_24227);
nand U25832 (N_25832,N_24402,N_24239);
and U25833 (N_25833,N_24486,N_24056);
and U25834 (N_25834,N_24037,N_24594);
nand U25835 (N_25835,N_24097,N_24748);
nand U25836 (N_25836,N_24859,N_24020);
or U25837 (N_25837,N_24534,N_24177);
or U25838 (N_25838,N_24534,N_24341);
and U25839 (N_25839,N_24024,N_24806);
nand U25840 (N_25840,N_24501,N_24921);
nor U25841 (N_25841,N_24551,N_24911);
xnor U25842 (N_25842,N_24043,N_24079);
and U25843 (N_25843,N_24912,N_24661);
nor U25844 (N_25844,N_24053,N_24505);
xor U25845 (N_25845,N_24840,N_24531);
xnor U25846 (N_25846,N_24158,N_24733);
nand U25847 (N_25847,N_24283,N_24991);
xnor U25848 (N_25848,N_24023,N_24767);
or U25849 (N_25849,N_24926,N_24903);
and U25850 (N_25850,N_24768,N_24827);
or U25851 (N_25851,N_24200,N_24621);
and U25852 (N_25852,N_24373,N_24190);
nor U25853 (N_25853,N_24909,N_24587);
xor U25854 (N_25854,N_24988,N_24877);
nor U25855 (N_25855,N_24666,N_24906);
nand U25856 (N_25856,N_24460,N_24263);
nor U25857 (N_25857,N_24817,N_24534);
nor U25858 (N_25858,N_24320,N_24376);
and U25859 (N_25859,N_24675,N_24140);
xor U25860 (N_25860,N_24232,N_24417);
and U25861 (N_25861,N_24953,N_24874);
nand U25862 (N_25862,N_24017,N_24538);
nor U25863 (N_25863,N_24665,N_24561);
and U25864 (N_25864,N_24565,N_24619);
nor U25865 (N_25865,N_24757,N_24341);
xor U25866 (N_25866,N_24395,N_24096);
and U25867 (N_25867,N_24799,N_24179);
xor U25868 (N_25868,N_24491,N_24958);
nor U25869 (N_25869,N_24909,N_24550);
nand U25870 (N_25870,N_24835,N_24757);
nand U25871 (N_25871,N_24649,N_24771);
nor U25872 (N_25872,N_24172,N_24139);
xnor U25873 (N_25873,N_24748,N_24893);
xor U25874 (N_25874,N_24255,N_24517);
nor U25875 (N_25875,N_24926,N_24914);
and U25876 (N_25876,N_24754,N_24593);
and U25877 (N_25877,N_24497,N_24584);
nor U25878 (N_25878,N_24807,N_24948);
nand U25879 (N_25879,N_24311,N_24028);
or U25880 (N_25880,N_24845,N_24983);
or U25881 (N_25881,N_24790,N_24161);
and U25882 (N_25882,N_24770,N_24822);
nand U25883 (N_25883,N_24167,N_24874);
nor U25884 (N_25884,N_24128,N_24358);
or U25885 (N_25885,N_24012,N_24840);
xor U25886 (N_25886,N_24107,N_24611);
xnor U25887 (N_25887,N_24005,N_24059);
xnor U25888 (N_25888,N_24948,N_24352);
nor U25889 (N_25889,N_24922,N_24062);
or U25890 (N_25890,N_24727,N_24525);
nor U25891 (N_25891,N_24106,N_24142);
nor U25892 (N_25892,N_24606,N_24994);
xnor U25893 (N_25893,N_24253,N_24726);
nand U25894 (N_25894,N_24528,N_24488);
nand U25895 (N_25895,N_24777,N_24948);
xnor U25896 (N_25896,N_24344,N_24959);
and U25897 (N_25897,N_24291,N_24740);
and U25898 (N_25898,N_24139,N_24157);
and U25899 (N_25899,N_24171,N_24267);
nand U25900 (N_25900,N_24682,N_24908);
and U25901 (N_25901,N_24354,N_24416);
xnor U25902 (N_25902,N_24759,N_24715);
nor U25903 (N_25903,N_24701,N_24752);
or U25904 (N_25904,N_24620,N_24800);
xnor U25905 (N_25905,N_24933,N_24403);
xnor U25906 (N_25906,N_24409,N_24936);
and U25907 (N_25907,N_24040,N_24013);
or U25908 (N_25908,N_24178,N_24007);
and U25909 (N_25909,N_24315,N_24907);
nand U25910 (N_25910,N_24594,N_24803);
or U25911 (N_25911,N_24346,N_24158);
nand U25912 (N_25912,N_24009,N_24971);
xor U25913 (N_25913,N_24262,N_24396);
nand U25914 (N_25914,N_24671,N_24660);
and U25915 (N_25915,N_24257,N_24079);
or U25916 (N_25916,N_24615,N_24654);
or U25917 (N_25917,N_24212,N_24638);
nor U25918 (N_25918,N_24239,N_24799);
or U25919 (N_25919,N_24018,N_24847);
nand U25920 (N_25920,N_24249,N_24023);
nand U25921 (N_25921,N_24923,N_24469);
nand U25922 (N_25922,N_24363,N_24453);
nor U25923 (N_25923,N_24158,N_24255);
or U25924 (N_25924,N_24300,N_24931);
and U25925 (N_25925,N_24866,N_24863);
nand U25926 (N_25926,N_24978,N_24507);
nor U25927 (N_25927,N_24031,N_24731);
and U25928 (N_25928,N_24116,N_24971);
nand U25929 (N_25929,N_24474,N_24211);
nand U25930 (N_25930,N_24455,N_24200);
nand U25931 (N_25931,N_24239,N_24038);
xor U25932 (N_25932,N_24768,N_24902);
xnor U25933 (N_25933,N_24174,N_24882);
nor U25934 (N_25934,N_24075,N_24273);
and U25935 (N_25935,N_24388,N_24170);
nor U25936 (N_25936,N_24453,N_24213);
and U25937 (N_25937,N_24399,N_24005);
xnor U25938 (N_25938,N_24869,N_24868);
xnor U25939 (N_25939,N_24378,N_24415);
or U25940 (N_25940,N_24771,N_24572);
nor U25941 (N_25941,N_24943,N_24507);
or U25942 (N_25942,N_24035,N_24528);
nand U25943 (N_25943,N_24091,N_24905);
nand U25944 (N_25944,N_24070,N_24900);
or U25945 (N_25945,N_24796,N_24866);
xor U25946 (N_25946,N_24800,N_24237);
nor U25947 (N_25947,N_24448,N_24281);
or U25948 (N_25948,N_24856,N_24198);
nor U25949 (N_25949,N_24113,N_24380);
nor U25950 (N_25950,N_24510,N_24270);
nand U25951 (N_25951,N_24928,N_24723);
or U25952 (N_25952,N_24542,N_24905);
nand U25953 (N_25953,N_24640,N_24427);
xnor U25954 (N_25954,N_24613,N_24418);
or U25955 (N_25955,N_24932,N_24710);
xnor U25956 (N_25956,N_24475,N_24219);
or U25957 (N_25957,N_24063,N_24809);
nor U25958 (N_25958,N_24964,N_24268);
nor U25959 (N_25959,N_24056,N_24177);
and U25960 (N_25960,N_24553,N_24893);
nand U25961 (N_25961,N_24132,N_24378);
nand U25962 (N_25962,N_24072,N_24479);
nor U25963 (N_25963,N_24992,N_24395);
and U25964 (N_25964,N_24196,N_24214);
nand U25965 (N_25965,N_24975,N_24806);
and U25966 (N_25966,N_24093,N_24954);
nor U25967 (N_25967,N_24522,N_24581);
nand U25968 (N_25968,N_24701,N_24317);
and U25969 (N_25969,N_24776,N_24540);
nor U25970 (N_25970,N_24917,N_24320);
nand U25971 (N_25971,N_24028,N_24358);
nand U25972 (N_25972,N_24909,N_24288);
and U25973 (N_25973,N_24681,N_24938);
xor U25974 (N_25974,N_24264,N_24768);
xnor U25975 (N_25975,N_24616,N_24219);
nand U25976 (N_25976,N_24629,N_24220);
nor U25977 (N_25977,N_24572,N_24787);
or U25978 (N_25978,N_24854,N_24453);
or U25979 (N_25979,N_24583,N_24266);
and U25980 (N_25980,N_24154,N_24536);
xor U25981 (N_25981,N_24838,N_24686);
and U25982 (N_25982,N_24148,N_24700);
nor U25983 (N_25983,N_24927,N_24752);
or U25984 (N_25984,N_24221,N_24319);
or U25985 (N_25985,N_24348,N_24902);
or U25986 (N_25986,N_24382,N_24952);
and U25987 (N_25987,N_24437,N_24533);
and U25988 (N_25988,N_24854,N_24645);
nor U25989 (N_25989,N_24342,N_24530);
and U25990 (N_25990,N_24349,N_24404);
nor U25991 (N_25991,N_24785,N_24692);
and U25992 (N_25992,N_24036,N_24507);
nor U25993 (N_25993,N_24745,N_24995);
nand U25994 (N_25994,N_24859,N_24371);
or U25995 (N_25995,N_24523,N_24716);
and U25996 (N_25996,N_24802,N_24794);
nand U25997 (N_25997,N_24059,N_24284);
and U25998 (N_25998,N_24926,N_24964);
and U25999 (N_25999,N_24642,N_24814);
or U26000 (N_26000,N_25229,N_25144);
and U26001 (N_26001,N_25692,N_25726);
or U26002 (N_26002,N_25690,N_25629);
nor U26003 (N_26003,N_25363,N_25032);
nand U26004 (N_26004,N_25920,N_25109);
nand U26005 (N_26005,N_25068,N_25395);
and U26006 (N_26006,N_25438,N_25227);
or U26007 (N_26007,N_25168,N_25867);
xor U26008 (N_26008,N_25236,N_25556);
or U26009 (N_26009,N_25527,N_25804);
xor U26010 (N_26010,N_25073,N_25078);
nand U26011 (N_26011,N_25082,N_25150);
and U26012 (N_26012,N_25178,N_25321);
nor U26013 (N_26013,N_25206,N_25512);
or U26014 (N_26014,N_25297,N_25449);
or U26015 (N_26015,N_25169,N_25094);
nand U26016 (N_26016,N_25593,N_25662);
nor U26017 (N_26017,N_25407,N_25376);
and U26018 (N_26018,N_25429,N_25898);
nand U26019 (N_26019,N_25614,N_25682);
nor U26020 (N_26020,N_25295,N_25261);
nor U26021 (N_26021,N_25319,N_25218);
xnor U26022 (N_26022,N_25877,N_25696);
nand U26023 (N_26023,N_25093,N_25419);
and U26024 (N_26024,N_25632,N_25160);
xor U26025 (N_26025,N_25208,N_25003);
nor U26026 (N_26026,N_25984,N_25318);
xor U26027 (N_26027,N_25286,N_25561);
and U26028 (N_26028,N_25903,N_25356);
or U26029 (N_26029,N_25374,N_25240);
nand U26030 (N_26030,N_25535,N_25572);
nand U26031 (N_26031,N_25377,N_25263);
xor U26032 (N_26032,N_25901,N_25567);
or U26033 (N_26033,N_25031,N_25767);
nor U26034 (N_26034,N_25313,N_25891);
xnor U26035 (N_26035,N_25355,N_25796);
or U26036 (N_26036,N_25345,N_25679);
xor U26037 (N_26037,N_25445,N_25409);
or U26038 (N_26038,N_25481,N_25484);
nand U26039 (N_26039,N_25272,N_25882);
or U26040 (N_26040,N_25279,N_25669);
and U26041 (N_26041,N_25963,N_25067);
nand U26042 (N_26042,N_25809,N_25241);
and U26043 (N_26043,N_25581,N_25305);
or U26044 (N_26044,N_25618,N_25952);
xor U26045 (N_26045,N_25475,N_25372);
xor U26046 (N_26046,N_25118,N_25414);
nor U26047 (N_26047,N_25412,N_25846);
and U26048 (N_26048,N_25428,N_25045);
xor U26049 (N_26049,N_25025,N_25883);
and U26050 (N_26050,N_25871,N_25986);
nand U26051 (N_26051,N_25075,N_25502);
xor U26052 (N_26052,N_25860,N_25728);
nand U26053 (N_26053,N_25341,N_25401);
xor U26054 (N_26054,N_25411,N_25661);
and U26055 (N_26055,N_25199,N_25390);
nand U26056 (N_26056,N_25887,N_25080);
nand U26057 (N_26057,N_25365,N_25184);
xor U26058 (N_26058,N_25322,N_25708);
nor U26059 (N_26059,N_25856,N_25258);
xnor U26060 (N_26060,N_25852,N_25774);
nor U26061 (N_26061,N_25251,N_25756);
xor U26062 (N_26062,N_25837,N_25918);
or U26063 (N_26063,N_25293,N_25672);
and U26064 (N_26064,N_25522,N_25501);
nand U26065 (N_26065,N_25105,N_25284);
and U26066 (N_26066,N_25091,N_25344);
and U26067 (N_26067,N_25613,N_25235);
nand U26068 (N_26068,N_25802,N_25248);
or U26069 (N_26069,N_25748,N_25291);
nand U26070 (N_26070,N_25530,N_25717);
and U26071 (N_26071,N_25173,N_25975);
nor U26072 (N_26072,N_25283,N_25273);
nand U26073 (N_26073,N_25420,N_25571);
nand U26074 (N_26074,N_25495,N_25418);
nand U26075 (N_26075,N_25554,N_25113);
and U26076 (N_26076,N_25114,N_25050);
xor U26077 (N_26077,N_25587,N_25465);
nand U26078 (N_26078,N_25904,N_25044);
nand U26079 (N_26079,N_25924,N_25642);
nand U26080 (N_26080,N_25453,N_25680);
xor U26081 (N_26081,N_25673,N_25749);
nand U26082 (N_26082,N_25203,N_25541);
nand U26083 (N_26083,N_25597,N_25892);
or U26084 (N_26084,N_25562,N_25899);
or U26085 (N_26085,N_25187,N_25165);
nor U26086 (N_26086,N_25383,N_25134);
nand U26087 (N_26087,N_25239,N_25219);
nand U26088 (N_26088,N_25553,N_25474);
nor U26089 (N_26089,N_25166,N_25398);
xnor U26090 (N_26090,N_25463,N_25569);
nor U26091 (N_26091,N_25129,N_25012);
and U26092 (N_26092,N_25700,N_25685);
nor U26093 (N_26093,N_25909,N_25471);
or U26094 (N_26094,N_25879,N_25213);
xnor U26095 (N_26095,N_25639,N_25062);
nor U26096 (N_26096,N_25095,N_25624);
xnor U26097 (N_26097,N_25699,N_25037);
xor U26098 (N_26098,N_25835,N_25081);
xnor U26099 (N_26099,N_25009,N_25958);
nor U26100 (N_26100,N_25029,N_25244);
nand U26101 (N_26101,N_25935,N_25353);
or U26102 (N_26102,N_25996,N_25740);
nor U26103 (N_26103,N_25531,N_25011);
or U26104 (N_26104,N_25087,N_25149);
and U26105 (N_26105,N_25505,N_25352);
or U26106 (N_26106,N_25954,N_25308);
nand U26107 (N_26107,N_25539,N_25196);
xor U26108 (N_26108,N_25874,N_25112);
nor U26109 (N_26109,N_25072,N_25070);
nor U26110 (N_26110,N_25342,N_25022);
xnor U26111 (N_26111,N_25040,N_25575);
and U26112 (N_26112,N_25974,N_25999);
and U26113 (N_26113,N_25643,N_25450);
or U26114 (N_26114,N_25434,N_25048);
and U26115 (N_26115,N_25066,N_25697);
or U26116 (N_26116,N_25724,N_25551);
or U26117 (N_26117,N_25183,N_25282);
xor U26118 (N_26118,N_25052,N_25979);
xnor U26119 (N_26119,N_25900,N_25202);
or U26120 (N_26120,N_25266,N_25497);
nor U26121 (N_26121,N_25425,N_25090);
nor U26122 (N_26122,N_25224,N_25253);
and U26123 (N_26123,N_25274,N_25223);
nor U26124 (N_26124,N_25755,N_25443);
nand U26125 (N_26125,N_25875,N_25432);
nand U26126 (N_26126,N_25010,N_25312);
or U26127 (N_26127,N_25674,N_25705);
nand U26128 (N_26128,N_25464,N_25711);
nand U26129 (N_26129,N_25651,N_25890);
nand U26130 (N_26130,N_25143,N_25819);
and U26131 (N_26131,N_25611,N_25015);
xnor U26132 (N_26132,N_25084,N_25691);
nand U26133 (N_26133,N_25734,N_25628);
nand U26134 (N_26134,N_25098,N_25806);
and U26135 (N_26135,N_25681,N_25369);
nand U26136 (N_26136,N_25446,N_25167);
and U26137 (N_26137,N_25406,N_25217);
nor U26138 (N_26138,N_25041,N_25665);
xor U26139 (N_26139,N_25177,N_25185);
and U26140 (N_26140,N_25099,N_25402);
and U26141 (N_26141,N_25439,N_25600);
and U26142 (N_26142,N_25759,N_25013);
and U26143 (N_26143,N_25146,N_25831);
xnor U26144 (N_26144,N_25659,N_25907);
xor U26145 (N_26145,N_25941,N_25454);
xnor U26146 (N_26146,N_25155,N_25287);
and U26147 (N_26147,N_25710,N_25405);
xor U26148 (N_26148,N_25544,N_25153);
and U26149 (N_26149,N_25536,N_25018);
nor U26150 (N_26150,N_25195,N_25054);
xnor U26151 (N_26151,N_25957,N_25592);
xnor U26152 (N_26152,N_25116,N_25334);
nand U26153 (N_26153,N_25413,N_25268);
or U26154 (N_26154,N_25815,N_25220);
xnor U26155 (N_26155,N_25936,N_25051);
and U26156 (N_26156,N_25653,N_25579);
and U26157 (N_26157,N_25917,N_25715);
nand U26158 (N_26158,N_25230,N_25427);
or U26159 (N_26159,N_25237,N_25107);
and U26160 (N_26160,N_25750,N_25778);
nand U26161 (N_26161,N_25706,N_25945);
nor U26162 (N_26162,N_25069,N_25033);
and U26163 (N_26163,N_25126,N_25462);
nor U26164 (N_26164,N_25059,N_25676);
and U26165 (N_26165,N_25612,N_25049);
or U26166 (N_26166,N_25915,N_25793);
nor U26167 (N_26167,N_25647,N_25442);
and U26168 (N_26168,N_25626,N_25346);
xnor U26169 (N_26169,N_25136,N_25872);
and U26170 (N_26170,N_25096,N_25212);
nor U26171 (N_26171,N_25311,N_25128);
nand U26172 (N_26172,N_25232,N_25088);
nand U26173 (N_26173,N_25876,N_25922);
and U26174 (N_26174,N_25255,N_25437);
or U26175 (N_26175,N_25826,N_25790);
or U26176 (N_26176,N_25939,N_25119);
and U26177 (N_26177,N_25937,N_25323);
nand U26178 (N_26178,N_25703,N_25042);
xnor U26179 (N_26179,N_25823,N_25847);
or U26180 (N_26180,N_25730,N_25364);
nand U26181 (N_26181,N_25304,N_25504);
nor U26182 (N_26182,N_25381,N_25855);
nand U26183 (N_26183,N_25300,N_25543);
nand U26184 (N_26184,N_25786,N_25038);
and U26185 (N_26185,N_25275,N_25280);
and U26186 (N_26186,N_25214,N_25158);
or U26187 (N_26187,N_25947,N_25995);
nand U26188 (N_26188,N_25367,N_25714);
or U26189 (N_26189,N_25912,N_25865);
nor U26190 (N_26190,N_25154,N_25635);
and U26191 (N_26191,N_25063,N_25789);
or U26192 (N_26192,N_25511,N_25760);
or U26193 (N_26193,N_25967,N_25870);
xor U26194 (N_26194,N_25079,N_25638);
and U26195 (N_26195,N_25076,N_25186);
and U26196 (N_26196,N_25943,N_25188);
or U26197 (N_26197,N_25940,N_25962);
xnor U26198 (N_26198,N_25435,N_25812);
nor U26199 (N_26199,N_25523,N_25982);
nand U26200 (N_26200,N_25634,N_25529);
and U26201 (N_26201,N_25197,N_25176);
nand U26202 (N_26202,N_25932,N_25808);
nor U26203 (N_26203,N_25725,N_25399);
or U26204 (N_26204,N_25654,N_25889);
xor U26205 (N_26205,N_25580,N_25452);
nand U26206 (N_26206,N_25884,N_25306);
nand U26207 (N_26207,N_25397,N_25633);
xnor U26208 (N_26208,N_25245,N_25392);
nand U26209 (N_26209,N_25097,N_25469);
or U26210 (N_26210,N_25542,N_25247);
nor U26211 (N_26211,N_25631,N_25960);
nor U26212 (N_26212,N_25441,N_25668);
and U26213 (N_26213,N_25997,N_25732);
nand U26214 (N_26214,N_25189,N_25086);
or U26215 (N_26215,N_25822,N_25309);
nand U26216 (N_26216,N_25228,N_25617);
xor U26217 (N_26217,N_25520,N_25650);
nand U26218 (N_26218,N_25162,N_25499);
or U26219 (N_26219,N_25458,N_25844);
and U26220 (N_26220,N_25034,N_25824);
xor U26221 (N_26221,N_25148,N_25115);
nor U26222 (N_26222,N_25752,N_25254);
and U26223 (N_26223,N_25636,N_25138);
nor U26224 (N_26224,N_25704,N_25301);
nand U26225 (N_26225,N_25416,N_25316);
xnor U26226 (N_26226,N_25869,N_25565);
or U26227 (N_26227,N_25472,N_25001);
nand U26228 (N_26228,N_25741,N_25104);
and U26229 (N_26229,N_25071,N_25781);
xnor U26230 (N_26230,N_25378,N_25548);
nand U26231 (N_26231,N_25145,N_25393);
xnor U26232 (N_26232,N_25832,N_25246);
and U26233 (N_26233,N_25314,N_25956);
and U26234 (N_26234,N_25276,N_25267);
xnor U26235 (N_26235,N_25191,N_25850);
xor U26236 (N_26236,N_25426,N_25757);
and U26237 (N_26237,N_25482,N_25403);
nand U26238 (N_26238,N_25905,N_25307);
nor U26239 (N_26239,N_25787,N_25335);
nor U26240 (N_26240,N_25055,N_25330);
nor U26241 (N_26241,N_25948,N_25720);
or U26242 (N_26242,N_25836,N_25568);
nor U26243 (N_26243,N_25422,N_25599);
and U26244 (N_26244,N_25842,N_25607);
nor U26245 (N_26245,N_25332,N_25921);
nand U26246 (N_26246,N_25016,N_25961);
xor U26247 (N_26247,N_25667,N_25289);
xor U26248 (N_26248,N_25983,N_25598);
xnor U26249 (N_26249,N_25368,N_25616);
nand U26250 (N_26250,N_25340,N_25135);
xnor U26251 (N_26251,N_25886,N_25798);
xor U26252 (N_26252,N_25591,N_25739);
xor U26253 (N_26253,N_25210,N_25596);
nor U26254 (N_26254,N_25359,N_25843);
xor U26255 (N_26255,N_25573,N_25758);
and U26256 (N_26256,N_25394,N_25215);
nor U26257 (N_26257,N_25973,N_25468);
nor U26258 (N_26258,N_25821,N_25585);
xnor U26259 (N_26259,N_25451,N_25868);
nor U26260 (N_26260,N_25737,N_25777);
and U26261 (N_26261,N_25343,N_25566);
and U26262 (N_26262,N_25396,N_25582);
or U26263 (N_26263,N_25026,N_25648);
nand U26264 (N_26264,N_25866,N_25124);
or U26265 (N_26265,N_25658,N_25926);
and U26266 (N_26266,N_25222,N_25689);
nor U26267 (N_26267,N_25117,N_25294);
and U26268 (N_26268,N_25198,N_25841);
nor U26269 (N_26269,N_25019,N_25814);
or U26270 (N_26270,N_25959,N_25719);
or U26271 (N_26271,N_25382,N_25200);
nor U26272 (N_26272,N_25557,N_25234);
nand U26273 (N_26273,N_25564,N_25763);
xor U26274 (N_26274,N_25992,N_25404);
nor U26275 (N_26275,N_25400,N_25545);
or U26276 (N_26276,N_25942,N_25339);
xor U26277 (N_26277,N_25328,N_25361);
nand U26278 (N_26278,N_25640,N_25857);
nand U26279 (N_26279,N_25265,N_25455);
nand U26280 (N_26280,N_25457,N_25385);
nand U26281 (N_26281,N_25863,N_25209);
nor U26282 (N_26282,N_25838,N_25830);
nand U26283 (N_26283,N_25485,N_25510);
xor U26284 (N_26284,N_25964,N_25036);
nor U26285 (N_26285,N_25546,N_25873);
nand U26286 (N_26286,N_25174,N_25745);
nand U26287 (N_26287,N_25586,N_25500);
nor U26288 (N_26288,N_25743,N_25965);
nand U26289 (N_26289,N_25270,N_25221);
xnor U26290 (N_26290,N_25906,N_25298);
xnor U26291 (N_26291,N_25656,N_25448);
and U26292 (N_26292,N_25480,N_25718);
nand U26293 (N_26293,N_25675,N_25461);
nand U26294 (N_26294,N_25595,N_25043);
nand U26295 (N_26295,N_25494,N_25285);
nand U26296 (N_26296,N_25688,N_25989);
and U26297 (N_26297,N_25046,N_25483);
or U26298 (N_26298,N_25845,N_25834);
nand U26299 (N_26299,N_25619,N_25243);
nor U26300 (N_26300,N_25366,N_25594);
nor U26301 (N_26301,N_25201,N_25147);
xor U26302 (N_26302,N_25506,N_25327);
nor U26303 (N_26303,N_25417,N_25137);
nor U26304 (N_26304,N_25408,N_25584);
and U26305 (N_26305,N_25558,N_25861);
xnor U26306 (N_26306,N_25934,N_25017);
or U26307 (N_26307,N_25157,N_25609);
and U26308 (N_26308,N_25881,N_25813);
xnor U26309 (N_26309,N_25005,N_25620);
or U26310 (N_26310,N_25955,N_25440);
nand U26311 (N_26311,N_25083,N_25902);
xnor U26312 (N_26312,N_25061,N_25772);
xnor U26313 (N_26313,N_25103,N_25047);
and U26314 (N_26314,N_25123,N_25858);
or U26315 (N_26315,N_25570,N_25583);
nand U26316 (N_26316,N_25931,N_25456);
xnor U26317 (N_26317,N_25677,N_25803);
xor U26318 (N_26318,N_25770,N_25436);
and U26319 (N_26319,N_25721,N_25788);
nand U26320 (N_26320,N_25514,N_25671);
nand U26321 (N_26321,N_25389,N_25998);
or U26322 (N_26322,N_25827,N_25338);
xnor U26323 (N_26323,N_25373,N_25193);
nand U26324 (N_26324,N_25775,N_25292);
nor U26325 (N_26325,N_25120,N_25459);
and U26326 (N_26326,N_25768,N_25664);
xor U26327 (N_26327,N_25204,N_25492);
nor U26328 (N_26328,N_25028,N_25919);
and U26329 (N_26329,N_25938,N_25387);
or U26330 (N_26330,N_25779,N_25362);
nor U26331 (N_26331,N_25498,N_25625);
and U26332 (N_26332,N_25713,N_25683);
and U26333 (N_26333,N_25916,N_25657);
or U26334 (N_26334,N_25466,N_25131);
nor U26335 (N_26335,N_25944,N_25560);
nand U26336 (N_26336,N_25516,N_25762);
nand U26337 (N_26337,N_25862,N_25142);
nand U26338 (N_26338,N_25641,N_25507);
and U26339 (N_26339,N_25260,N_25946);
and U26340 (N_26340,N_25994,N_25347);
nor U26341 (N_26341,N_25290,N_25526);
xor U26342 (N_26342,N_25655,N_25649);
nand U26343 (N_26343,N_25773,N_25388);
xnor U26344 (N_26344,N_25172,N_25085);
nand U26345 (N_26345,N_25735,N_25666);
xnor U26346 (N_26346,N_25460,N_25329);
nor U26347 (N_26347,N_25302,N_25859);
and U26348 (N_26348,N_25532,N_25547);
xor U26349 (N_26349,N_25895,N_25360);
or U26350 (N_26350,N_25391,N_25577);
nor U26351 (N_26351,N_25927,N_25252);
nand U26352 (N_26352,N_25077,N_25800);
and U26353 (N_26353,N_25893,N_25693);
xnor U26354 (N_26354,N_25180,N_25980);
xnor U26355 (N_26355,N_25431,N_25503);
nand U26356 (N_26356,N_25550,N_25021);
nand U26357 (N_26357,N_25008,N_25035);
xor U26358 (N_26358,N_25277,N_25249);
nor U26359 (N_26359,N_25132,N_25722);
nor U26360 (N_26360,N_25825,N_25194);
nor U26361 (N_26361,N_25479,N_25473);
xnor U26362 (N_26362,N_25805,N_25623);
xnor U26363 (N_26363,N_25100,N_25549);
and U26364 (N_26364,N_25039,N_25170);
nand U26365 (N_26365,N_25242,N_25761);
and U26366 (N_26366,N_25589,N_25751);
nor U26367 (N_26367,N_25508,N_25652);
or U26368 (N_26368,N_25766,N_25559);
xor U26369 (N_26369,N_25348,N_25192);
nand U26370 (N_26370,N_25660,N_25092);
nand U26371 (N_26371,N_25007,N_25140);
and U26372 (N_26372,N_25910,N_25002);
nor U26373 (N_26373,N_25264,N_25971);
and U26374 (N_26374,N_25027,N_25020);
and U26375 (N_26375,N_25970,N_25602);
nor U26376 (N_26376,N_25089,N_25430);
or U26377 (N_26377,N_25784,N_25226);
xnor U26378 (N_26378,N_25753,N_25238);
nand U26379 (N_26379,N_25256,N_25175);
nor U26380 (N_26380,N_25911,N_25349);
or U26381 (N_26381,N_25953,N_25179);
nand U26382 (N_26382,N_25670,N_25969);
xnor U26383 (N_26383,N_25731,N_25818);
or U26384 (N_26384,N_25949,N_25331);
or U26385 (N_26385,N_25744,N_25701);
and U26386 (N_26386,N_25684,N_25888);
nand U26387 (N_26387,N_25929,N_25278);
or U26388 (N_26388,N_25791,N_25151);
and U26389 (N_26389,N_25608,N_25820);
or U26390 (N_26390,N_25490,N_25106);
or U26391 (N_26391,N_25326,N_25783);
and U26392 (N_26392,N_25152,N_25156);
and U26393 (N_26393,N_25742,N_25782);
xor U26394 (N_26394,N_25030,N_25207);
or U26395 (N_26395,N_25769,N_25707);
nand U26396 (N_26396,N_25840,N_25590);
nand U26397 (N_26397,N_25977,N_25424);
or U26398 (N_26398,N_25771,N_25491);
and U26399 (N_26399,N_25627,N_25060);
and U26400 (N_26400,N_25563,N_25317);
nand U26401 (N_26401,N_25333,N_25914);
and U26402 (N_26402,N_25375,N_25923);
xnor U26403 (N_26403,N_25896,N_25880);
or U26404 (N_26404,N_25733,N_25644);
and U26405 (N_26405,N_25518,N_25930);
and U26406 (N_26406,N_25004,N_25878);
xor U26407 (N_26407,N_25476,N_25555);
nor U26408 (N_26408,N_25006,N_25130);
or U26409 (N_26409,N_25190,N_25588);
and U26410 (N_26410,N_25271,N_25951);
nand U26411 (N_26411,N_25358,N_25574);
or U26412 (N_26412,N_25534,N_25161);
or U26413 (N_26413,N_25678,N_25351);
nor U26414 (N_26414,N_25509,N_25380);
nand U26415 (N_26415,N_25801,N_25829);
nor U26416 (N_26416,N_25621,N_25848);
and U26417 (N_26417,N_25606,N_25727);
nand U26418 (N_26418,N_25601,N_25467);
or U26419 (N_26419,N_25849,N_25533);
nor U26420 (N_26420,N_25864,N_25171);
xor U26421 (N_26421,N_25310,N_25288);
nor U26422 (N_26422,N_25540,N_25746);
and U26423 (N_26423,N_25552,N_25121);
nor U26424 (N_26424,N_25250,N_25064);
nand U26425 (N_26425,N_25433,N_25630);
xnor U26426 (N_26426,N_25164,N_25410);
nand U26427 (N_26427,N_25976,N_25933);
nor U26428 (N_26428,N_25993,N_25139);
and U26429 (N_26429,N_25111,N_25159);
xor U26430 (N_26430,N_25127,N_25637);
xnor U26431 (N_26431,N_25981,N_25698);
nor U26432 (N_26432,N_25797,N_25421);
xnor U26433 (N_26433,N_25325,N_25663);
nand U26434 (N_26434,N_25894,N_25470);
nand U26435 (N_26435,N_25315,N_25320);
and U26436 (N_26436,N_25776,N_25000);
nor U26437 (N_26437,N_25102,N_25972);
xnor U26438 (N_26438,N_25141,N_25521);
and U26439 (N_26439,N_25794,N_25799);
nand U26440 (N_26440,N_25122,N_25816);
nand U26441 (N_26441,N_25053,N_25747);
nor U26442 (N_26442,N_25925,N_25477);
and U26443 (N_26443,N_25354,N_25828);
xnor U26444 (N_26444,N_25754,N_25336);
xor U26445 (N_26445,N_25576,N_25444);
and U26446 (N_26446,N_25513,N_25324);
and U26447 (N_26447,N_25181,N_25269);
xor U26448 (N_26448,N_25058,N_25785);
or U26449 (N_26449,N_25225,N_25296);
nand U26450 (N_26450,N_25604,N_25610);
xnor U26451 (N_26451,N_25985,N_25489);
nand U26452 (N_26452,N_25057,N_25065);
or U26453 (N_26453,N_25885,N_25615);
or U26454 (N_26454,N_25163,N_25478);
xor U26455 (N_26455,N_25795,N_25056);
and U26456 (N_26456,N_25908,N_25839);
nand U26457 (N_26457,N_25496,N_25024);
nor U26458 (N_26458,N_25231,N_25108);
xor U26459 (N_26459,N_25528,N_25897);
nor U26460 (N_26460,N_25233,N_25738);
nor U26461 (N_26461,N_25350,N_25303);
nand U26462 (N_26462,N_25493,N_25990);
nor U26463 (N_26463,N_25695,N_25694);
xor U26464 (N_26464,N_25991,N_25780);
or U26465 (N_26465,N_25537,N_25423);
or U26466 (N_26466,N_25687,N_25357);
and U26467 (N_26467,N_25764,N_25259);
or U26468 (N_26468,N_25216,N_25205);
nand U26469 (N_26469,N_25023,N_25101);
xnor U26470 (N_26470,N_25281,N_25519);
xor U26471 (N_26471,N_25686,N_25928);
nor U26472 (N_26472,N_25125,N_25645);
or U26473 (N_26473,N_25736,N_25578);
nor U26474 (N_26474,N_25370,N_25833);
xor U26475 (N_26475,N_25133,N_25712);
and U26476 (N_26476,N_25913,N_25810);
nor U26477 (N_26477,N_25646,N_25447);
nand U26478 (N_26478,N_25262,N_25807);
and U26479 (N_26479,N_25978,N_25379);
xnor U26480 (N_26480,N_25014,N_25603);
nor U26481 (N_26481,N_25386,N_25486);
nand U26482 (N_26482,N_25182,N_25709);
nand U26483 (N_26483,N_25622,N_25966);
or U26484 (N_26484,N_25487,N_25723);
or U26485 (N_26485,N_25987,N_25817);
xor U26486 (N_26486,N_25525,N_25371);
xor U26487 (N_26487,N_25257,N_25488);
and U26488 (N_26488,N_25716,N_25299);
and U26489 (N_26489,N_25074,N_25524);
xnor U26490 (N_26490,N_25792,N_25517);
nor U26491 (N_26491,N_25702,N_25988);
nand U26492 (N_26492,N_25515,N_25811);
xor U26493 (N_26493,N_25211,N_25765);
and U26494 (N_26494,N_25384,N_25538);
xnor U26495 (N_26495,N_25968,N_25851);
or U26496 (N_26496,N_25415,N_25110);
and U26497 (N_26497,N_25854,N_25605);
xnor U26498 (N_26498,N_25337,N_25950);
nor U26499 (N_26499,N_25853,N_25729);
nand U26500 (N_26500,N_25618,N_25846);
or U26501 (N_26501,N_25300,N_25431);
or U26502 (N_26502,N_25771,N_25122);
nand U26503 (N_26503,N_25590,N_25103);
or U26504 (N_26504,N_25607,N_25451);
nand U26505 (N_26505,N_25883,N_25650);
nand U26506 (N_26506,N_25352,N_25576);
nand U26507 (N_26507,N_25308,N_25832);
nand U26508 (N_26508,N_25938,N_25585);
and U26509 (N_26509,N_25565,N_25945);
nand U26510 (N_26510,N_25114,N_25873);
and U26511 (N_26511,N_25821,N_25001);
and U26512 (N_26512,N_25718,N_25468);
xor U26513 (N_26513,N_25133,N_25040);
or U26514 (N_26514,N_25448,N_25545);
and U26515 (N_26515,N_25947,N_25073);
xor U26516 (N_26516,N_25998,N_25463);
or U26517 (N_26517,N_25826,N_25234);
xor U26518 (N_26518,N_25174,N_25545);
and U26519 (N_26519,N_25516,N_25143);
nor U26520 (N_26520,N_25636,N_25225);
or U26521 (N_26521,N_25599,N_25995);
nand U26522 (N_26522,N_25217,N_25474);
or U26523 (N_26523,N_25180,N_25211);
xnor U26524 (N_26524,N_25892,N_25762);
xnor U26525 (N_26525,N_25288,N_25906);
xnor U26526 (N_26526,N_25472,N_25417);
or U26527 (N_26527,N_25395,N_25329);
or U26528 (N_26528,N_25603,N_25621);
xor U26529 (N_26529,N_25021,N_25826);
or U26530 (N_26530,N_25267,N_25735);
or U26531 (N_26531,N_25987,N_25437);
xor U26532 (N_26532,N_25673,N_25775);
xnor U26533 (N_26533,N_25135,N_25725);
or U26534 (N_26534,N_25869,N_25751);
nand U26535 (N_26535,N_25869,N_25572);
and U26536 (N_26536,N_25137,N_25891);
or U26537 (N_26537,N_25557,N_25191);
or U26538 (N_26538,N_25582,N_25547);
nor U26539 (N_26539,N_25109,N_25095);
and U26540 (N_26540,N_25192,N_25851);
and U26541 (N_26541,N_25558,N_25067);
or U26542 (N_26542,N_25124,N_25074);
and U26543 (N_26543,N_25606,N_25654);
nand U26544 (N_26544,N_25399,N_25770);
or U26545 (N_26545,N_25633,N_25359);
and U26546 (N_26546,N_25292,N_25960);
and U26547 (N_26547,N_25290,N_25143);
nor U26548 (N_26548,N_25402,N_25326);
nand U26549 (N_26549,N_25569,N_25616);
nand U26550 (N_26550,N_25141,N_25169);
nor U26551 (N_26551,N_25167,N_25018);
xor U26552 (N_26552,N_25869,N_25138);
or U26553 (N_26553,N_25709,N_25756);
xnor U26554 (N_26554,N_25138,N_25335);
xor U26555 (N_26555,N_25650,N_25536);
or U26556 (N_26556,N_25318,N_25515);
and U26557 (N_26557,N_25381,N_25556);
xnor U26558 (N_26558,N_25927,N_25635);
nand U26559 (N_26559,N_25340,N_25381);
nor U26560 (N_26560,N_25375,N_25127);
nand U26561 (N_26561,N_25192,N_25610);
nor U26562 (N_26562,N_25276,N_25808);
and U26563 (N_26563,N_25556,N_25036);
nand U26564 (N_26564,N_25260,N_25770);
nor U26565 (N_26565,N_25704,N_25062);
nor U26566 (N_26566,N_25508,N_25631);
nor U26567 (N_26567,N_25473,N_25441);
or U26568 (N_26568,N_25229,N_25570);
nor U26569 (N_26569,N_25357,N_25066);
nor U26570 (N_26570,N_25157,N_25207);
nor U26571 (N_26571,N_25595,N_25360);
or U26572 (N_26572,N_25791,N_25163);
or U26573 (N_26573,N_25523,N_25698);
or U26574 (N_26574,N_25033,N_25559);
xor U26575 (N_26575,N_25485,N_25569);
xor U26576 (N_26576,N_25087,N_25731);
and U26577 (N_26577,N_25423,N_25592);
xor U26578 (N_26578,N_25839,N_25092);
or U26579 (N_26579,N_25083,N_25360);
nor U26580 (N_26580,N_25525,N_25351);
xor U26581 (N_26581,N_25784,N_25826);
nand U26582 (N_26582,N_25822,N_25518);
or U26583 (N_26583,N_25686,N_25775);
nand U26584 (N_26584,N_25162,N_25285);
or U26585 (N_26585,N_25175,N_25961);
nand U26586 (N_26586,N_25055,N_25253);
nand U26587 (N_26587,N_25921,N_25368);
and U26588 (N_26588,N_25936,N_25742);
nor U26589 (N_26589,N_25117,N_25483);
and U26590 (N_26590,N_25511,N_25534);
or U26591 (N_26591,N_25118,N_25811);
and U26592 (N_26592,N_25554,N_25413);
nand U26593 (N_26593,N_25174,N_25601);
nor U26594 (N_26594,N_25779,N_25515);
xnor U26595 (N_26595,N_25289,N_25336);
xor U26596 (N_26596,N_25961,N_25813);
and U26597 (N_26597,N_25177,N_25058);
nor U26598 (N_26598,N_25226,N_25805);
xor U26599 (N_26599,N_25196,N_25536);
nor U26600 (N_26600,N_25542,N_25481);
nand U26601 (N_26601,N_25263,N_25328);
xnor U26602 (N_26602,N_25825,N_25988);
xor U26603 (N_26603,N_25616,N_25048);
nor U26604 (N_26604,N_25255,N_25529);
nor U26605 (N_26605,N_25309,N_25712);
nand U26606 (N_26606,N_25859,N_25795);
nor U26607 (N_26607,N_25256,N_25000);
and U26608 (N_26608,N_25160,N_25363);
xor U26609 (N_26609,N_25806,N_25132);
nand U26610 (N_26610,N_25857,N_25886);
nor U26611 (N_26611,N_25099,N_25256);
nand U26612 (N_26612,N_25498,N_25393);
or U26613 (N_26613,N_25662,N_25894);
xor U26614 (N_26614,N_25626,N_25919);
xor U26615 (N_26615,N_25204,N_25431);
nand U26616 (N_26616,N_25376,N_25399);
or U26617 (N_26617,N_25796,N_25162);
or U26618 (N_26618,N_25470,N_25080);
and U26619 (N_26619,N_25805,N_25508);
nand U26620 (N_26620,N_25991,N_25777);
and U26621 (N_26621,N_25917,N_25617);
xor U26622 (N_26622,N_25918,N_25893);
and U26623 (N_26623,N_25712,N_25694);
nor U26624 (N_26624,N_25151,N_25110);
nand U26625 (N_26625,N_25050,N_25958);
nor U26626 (N_26626,N_25141,N_25335);
nand U26627 (N_26627,N_25352,N_25625);
nor U26628 (N_26628,N_25062,N_25243);
xor U26629 (N_26629,N_25149,N_25738);
or U26630 (N_26630,N_25725,N_25535);
nor U26631 (N_26631,N_25246,N_25149);
xor U26632 (N_26632,N_25774,N_25953);
nor U26633 (N_26633,N_25590,N_25983);
nand U26634 (N_26634,N_25739,N_25362);
xor U26635 (N_26635,N_25990,N_25774);
nand U26636 (N_26636,N_25835,N_25945);
or U26637 (N_26637,N_25125,N_25654);
or U26638 (N_26638,N_25767,N_25533);
nand U26639 (N_26639,N_25429,N_25622);
or U26640 (N_26640,N_25512,N_25657);
or U26641 (N_26641,N_25992,N_25186);
nand U26642 (N_26642,N_25192,N_25966);
nor U26643 (N_26643,N_25897,N_25029);
and U26644 (N_26644,N_25259,N_25804);
xnor U26645 (N_26645,N_25186,N_25424);
nand U26646 (N_26646,N_25941,N_25561);
or U26647 (N_26647,N_25838,N_25672);
nor U26648 (N_26648,N_25006,N_25508);
nand U26649 (N_26649,N_25928,N_25003);
and U26650 (N_26650,N_25949,N_25533);
or U26651 (N_26651,N_25864,N_25873);
xnor U26652 (N_26652,N_25613,N_25780);
xnor U26653 (N_26653,N_25256,N_25249);
nand U26654 (N_26654,N_25320,N_25510);
and U26655 (N_26655,N_25476,N_25988);
and U26656 (N_26656,N_25282,N_25602);
nor U26657 (N_26657,N_25125,N_25525);
or U26658 (N_26658,N_25151,N_25730);
nand U26659 (N_26659,N_25785,N_25679);
nor U26660 (N_26660,N_25479,N_25586);
xnor U26661 (N_26661,N_25293,N_25765);
or U26662 (N_26662,N_25205,N_25169);
xor U26663 (N_26663,N_25637,N_25893);
and U26664 (N_26664,N_25392,N_25499);
xnor U26665 (N_26665,N_25491,N_25726);
xnor U26666 (N_26666,N_25180,N_25155);
xor U26667 (N_26667,N_25943,N_25668);
or U26668 (N_26668,N_25927,N_25587);
xor U26669 (N_26669,N_25717,N_25869);
nor U26670 (N_26670,N_25331,N_25442);
xor U26671 (N_26671,N_25616,N_25767);
and U26672 (N_26672,N_25182,N_25474);
or U26673 (N_26673,N_25895,N_25668);
or U26674 (N_26674,N_25976,N_25074);
or U26675 (N_26675,N_25249,N_25519);
or U26676 (N_26676,N_25020,N_25448);
and U26677 (N_26677,N_25250,N_25368);
xor U26678 (N_26678,N_25349,N_25860);
or U26679 (N_26679,N_25594,N_25489);
nor U26680 (N_26680,N_25182,N_25744);
nor U26681 (N_26681,N_25267,N_25333);
nor U26682 (N_26682,N_25185,N_25465);
nor U26683 (N_26683,N_25204,N_25689);
or U26684 (N_26684,N_25911,N_25429);
nand U26685 (N_26685,N_25649,N_25195);
nand U26686 (N_26686,N_25452,N_25951);
xnor U26687 (N_26687,N_25757,N_25824);
nor U26688 (N_26688,N_25847,N_25998);
and U26689 (N_26689,N_25650,N_25091);
nor U26690 (N_26690,N_25984,N_25841);
and U26691 (N_26691,N_25203,N_25194);
nor U26692 (N_26692,N_25430,N_25545);
nand U26693 (N_26693,N_25510,N_25884);
and U26694 (N_26694,N_25090,N_25153);
xnor U26695 (N_26695,N_25114,N_25831);
nor U26696 (N_26696,N_25920,N_25587);
nand U26697 (N_26697,N_25167,N_25683);
xor U26698 (N_26698,N_25828,N_25266);
and U26699 (N_26699,N_25949,N_25472);
and U26700 (N_26700,N_25575,N_25012);
or U26701 (N_26701,N_25305,N_25800);
and U26702 (N_26702,N_25081,N_25448);
or U26703 (N_26703,N_25848,N_25209);
xor U26704 (N_26704,N_25088,N_25509);
or U26705 (N_26705,N_25136,N_25800);
nor U26706 (N_26706,N_25299,N_25723);
or U26707 (N_26707,N_25556,N_25577);
nand U26708 (N_26708,N_25947,N_25094);
nand U26709 (N_26709,N_25955,N_25844);
or U26710 (N_26710,N_25739,N_25610);
nand U26711 (N_26711,N_25452,N_25093);
or U26712 (N_26712,N_25301,N_25863);
nand U26713 (N_26713,N_25771,N_25364);
nor U26714 (N_26714,N_25651,N_25250);
nor U26715 (N_26715,N_25409,N_25544);
and U26716 (N_26716,N_25989,N_25459);
and U26717 (N_26717,N_25969,N_25638);
and U26718 (N_26718,N_25787,N_25305);
nor U26719 (N_26719,N_25250,N_25159);
nor U26720 (N_26720,N_25994,N_25634);
and U26721 (N_26721,N_25260,N_25408);
or U26722 (N_26722,N_25285,N_25740);
and U26723 (N_26723,N_25771,N_25159);
and U26724 (N_26724,N_25641,N_25568);
nor U26725 (N_26725,N_25478,N_25337);
nor U26726 (N_26726,N_25913,N_25439);
or U26727 (N_26727,N_25058,N_25403);
or U26728 (N_26728,N_25667,N_25182);
and U26729 (N_26729,N_25214,N_25603);
xor U26730 (N_26730,N_25020,N_25772);
or U26731 (N_26731,N_25107,N_25152);
nor U26732 (N_26732,N_25945,N_25184);
nand U26733 (N_26733,N_25584,N_25075);
xor U26734 (N_26734,N_25194,N_25062);
and U26735 (N_26735,N_25146,N_25753);
and U26736 (N_26736,N_25370,N_25250);
and U26737 (N_26737,N_25527,N_25360);
xnor U26738 (N_26738,N_25374,N_25077);
nor U26739 (N_26739,N_25020,N_25503);
nor U26740 (N_26740,N_25698,N_25065);
nor U26741 (N_26741,N_25115,N_25415);
and U26742 (N_26742,N_25319,N_25012);
nor U26743 (N_26743,N_25625,N_25025);
nand U26744 (N_26744,N_25202,N_25930);
or U26745 (N_26745,N_25341,N_25536);
or U26746 (N_26746,N_25705,N_25546);
nand U26747 (N_26747,N_25836,N_25153);
nor U26748 (N_26748,N_25645,N_25863);
or U26749 (N_26749,N_25822,N_25421);
or U26750 (N_26750,N_25409,N_25222);
or U26751 (N_26751,N_25166,N_25541);
nor U26752 (N_26752,N_25800,N_25259);
nand U26753 (N_26753,N_25124,N_25777);
and U26754 (N_26754,N_25019,N_25885);
or U26755 (N_26755,N_25399,N_25920);
or U26756 (N_26756,N_25851,N_25843);
and U26757 (N_26757,N_25570,N_25916);
and U26758 (N_26758,N_25152,N_25669);
xnor U26759 (N_26759,N_25801,N_25568);
nand U26760 (N_26760,N_25318,N_25092);
nor U26761 (N_26761,N_25751,N_25239);
xnor U26762 (N_26762,N_25063,N_25906);
nand U26763 (N_26763,N_25660,N_25102);
or U26764 (N_26764,N_25978,N_25717);
and U26765 (N_26765,N_25654,N_25361);
and U26766 (N_26766,N_25587,N_25608);
nand U26767 (N_26767,N_25487,N_25456);
xor U26768 (N_26768,N_25844,N_25757);
xnor U26769 (N_26769,N_25872,N_25182);
nand U26770 (N_26770,N_25110,N_25761);
and U26771 (N_26771,N_25993,N_25826);
nand U26772 (N_26772,N_25416,N_25032);
nor U26773 (N_26773,N_25704,N_25474);
xnor U26774 (N_26774,N_25799,N_25447);
or U26775 (N_26775,N_25262,N_25573);
nor U26776 (N_26776,N_25406,N_25088);
xnor U26777 (N_26777,N_25186,N_25461);
nor U26778 (N_26778,N_25987,N_25062);
or U26779 (N_26779,N_25289,N_25481);
nor U26780 (N_26780,N_25574,N_25761);
and U26781 (N_26781,N_25377,N_25458);
xor U26782 (N_26782,N_25422,N_25793);
nor U26783 (N_26783,N_25952,N_25569);
nor U26784 (N_26784,N_25431,N_25125);
nand U26785 (N_26785,N_25084,N_25119);
or U26786 (N_26786,N_25618,N_25459);
nor U26787 (N_26787,N_25773,N_25271);
or U26788 (N_26788,N_25197,N_25968);
xor U26789 (N_26789,N_25570,N_25601);
xnor U26790 (N_26790,N_25053,N_25083);
or U26791 (N_26791,N_25861,N_25989);
and U26792 (N_26792,N_25511,N_25989);
and U26793 (N_26793,N_25584,N_25386);
nand U26794 (N_26794,N_25244,N_25697);
and U26795 (N_26795,N_25428,N_25246);
or U26796 (N_26796,N_25755,N_25916);
nor U26797 (N_26797,N_25325,N_25642);
nand U26798 (N_26798,N_25225,N_25157);
xor U26799 (N_26799,N_25755,N_25900);
and U26800 (N_26800,N_25299,N_25322);
and U26801 (N_26801,N_25547,N_25736);
and U26802 (N_26802,N_25853,N_25337);
nand U26803 (N_26803,N_25264,N_25130);
xnor U26804 (N_26804,N_25692,N_25032);
xor U26805 (N_26805,N_25462,N_25133);
nand U26806 (N_26806,N_25186,N_25325);
nand U26807 (N_26807,N_25717,N_25107);
or U26808 (N_26808,N_25944,N_25620);
nor U26809 (N_26809,N_25427,N_25340);
nor U26810 (N_26810,N_25774,N_25996);
or U26811 (N_26811,N_25996,N_25350);
xor U26812 (N_26812,N_25357,N_25824);
nand U26813 (N_26813,N_25762,N_25683);
nor U26814 (N_26814,N_25936,N_25221);
xor U26815 (N_26815,N_25407,N_25972);
nor U26816 (N_26816,N_25287,N_25879);
xor U26817 (N_26817,N_25332,N_25547);
nor U26818 (N_26818,N_25514,N_25204);
or U26819 (N_26819,N_25985,N_25794);
xor U26820 (N_26820,N_25293,N_25736);
xor U26821 (N_26821,N_25313,N_25430);
and U26822 (N_26822,N_25961,N_25525);
or U26823 (N_26823,N_25913,N_25325);
and U26824 (N_26824,N_25608,N_25370);
or U26825 (N_26825,N_25541,N_25211);
xnor U26826 (N_26826,N_25012,N_25046);
nor U26827 (N_26827,N_25336,N_25148);
nor U26828 (N_26828,N_25531,N_25169);
xor U26829 (N_26829,N_25916,N_25806);
xnor U26830 (N_26830,N_25997,N_25576);
nand U26831 (N_26831,N_25799,N_25365);
and U26832 (N_26832,N_25291,N_25141);
and U26833 (N_26833,N_25470,N_25739);
nand U26834 (N_26834,N_25711,N_25828);
or U26835 (N_26835,N_25598,N_25374);
nor U26836 (N_26836,N_25759,N_25055);
xor U26837 (N_26837,N_25429,N_25204);
nand U26838 (N_26838,N_25171,N_25521);
nor U26839 (N_26839,N_25156,N_25096);
or U26840 (N_26840,N_25506,N_25244);
and U26841 (N_26841,N_25319,N_25264);
and U26842 (N_26842,N_25865,N_25479);
xnor U26843 (N_26843,N_25952,N_25342);
or U26844 (N_26844,N_25804,N_25242);
nor U26845 (N_26845,N_25554,N_25181);
xnor U26846 (N_26846,N_25220,N_25789);
nor U26847 (N_26847,N_25173,N_25476);
xor U26848 (N_26848,N_25991,N_25342);
nor U26849 (N_26849,N_25454,N_25198);
and U26850 (N_26850,N_25790,N_25289);
xnor U26851 (N_26851,N_25767,N_25140);
nand U26852 (N_26852,N_25888,N_25165);
nand U26853 (N_26853,N_25318,N_25661);
nand U26854 (N_26854,N_25604,N_25188);
or U26855 (N_26855,N_25048,N_25807);
nor U26856 (N_26856,N_25011,N_25604);
nor U26857 (N_26857,N_25845,N_25289);
xor U26858 (N_26858,N_25330,N_25974);
xnor U26859 (N_26859,N_25666,N_25423);
xor U26860 (N_26860,N_25996,N_25091);
nand U26861 (N_26861,N_25933,N_25123);
xor U26862 (N_26862,N_25136,N_25446);
or U26863 (N_26863,N_25886,N_25078);
or U26864 (N_26864,N_25495,N_25399);
and U26865 (N_26865,N_25418,N_25215);
nor U26866 (N_26866,N_25502,N_25863);
and U26867 (N_26867,N_25783,N_25503);
xnor U26868 (N_26868,N_25706,N_25459);
nor U26869 (N_26869,N_25537,N_25002);
and U26870 (N_26870,N_25767,N_25947);
nor U26871 (N_26871,N_25468,N_25797);
nor U26872 (N_26872,N_25721,N_25445);
or U26873 (N_26873,N_25954,N_25185);
and U26874 (N_26874,N_25402,N_25785);
and U26875 (N_26875,N_25139,N_25955);
nor U26876 (N_26876,N_25104,N_25433);
xnor U26877 (N_26877,N_25448,N_25153);
nand U26878 (N_26878,N_25928,N_25403);
and U26879 (N_26879,N_25586,N_25937);
xnor U26880 (N_26880,N_25123,N_25342);
nor U26881 (N_26881,N_25453,N_25184);
nand U26882 (N_26882,N_25563,N_25204);
and U26883 (N_26883,N_25573,N_25002);
nand U26884 (N_26884,N_25904,N_25022);
or U26885 (N_26885,N_25435,N_25190);
xor U26886 (N_26886,N_25954,N_25742);
or U26887 (N_26887,N_25224,N_25102);
xnor U26888 (N_26888,N_25549,N_25979);
and U26889 (N_26889,N_25579,N_25621);
or U26890 (N_26890,N_25418,N_25006);
xor U26891 (N_26891,N_25688,N_25516);
or U26892 (N_26892,N_25541,N_25335);
and U26893 (N_26893,N_25848,N_25159);
xor U26894 (N_26894,N_25207,N_25036);
and U26895 (N_26895,N_25002,N_25487);
nand U26896 (N_26896,N_25255,N_25265);
xnor U26897 (N_26897,N_25220,N_25681);
nor U26898 (N_26898,N_25176,N_25862);
xnor U26899 (N_26899,N_25170,N_25509);
or U26900 (N_26900,N_25229,N_25619);
or U26901 (N_26901,N_25529,N_25441);
xnor U26902 (N_26902,N_25383,N_25787);
nand U26903 (N_26903,N_25004,N_25229);
nand U26904 (N_26904,N_25905,N_25853);
nor U26905 (N_26905,N_25949,N_25998);
and U26906 (N_26906,N_25628,N_25848);
or U26907 (N_26907,N_25621,N_25607);
and U26908 (N_26908,N_25630,N_25092);
and U26909 (N_26909,N_25290,N_25068);
or U26910 (N_26910,N_25388,N_25928);
nor U26911 (N_26911,N_25425,N_25104);
or U26912 (N_26912,N_25404,N_25387);
nor U26913 (N_26913,N_25108,N_25742);
or U26914 (N_26914,N_25875,N_25290);
nand U26915 (N_26915,N_25965,N_25348);
or U26916 (N_26916,N_25980,N_25050);
and U26917 (N_26917,N_25110,N_25316);
or U26918 (N_26918,N_25965,N_25783);
or U26919 (N_26919,N_25444,N_25796);
xnor U26920 (N_26920,N_25803,N_25317);
nand U26921 (N_26921,N_25803,N_25632);
nor U26922 (N_26922,N_25217,N_25595);
nor U26923 (N_26923,N_25614,N_25347);
or U26924 (N_26924,N_25855,N_25882);
nor U26925 (N_26925,N_25477,N_25311);
nand U26926 (N_26926,N_25108,N_25787);
nor U26927 (N_26927,N_25464,N_25708);
and U26928 (N_26928,N_25076,N_25340);
and U26929 (N_26929,N_25919,N_25279);
and U26930 (N_26930,N_25087,N_25025);
and U26931 (N_26931,N_25771,N_25972);
nor U26932 (N_26932,N_25709,N_25773);
nand U26933 (N_26933,N_25332,N_25933);
nand U26934 (N_26934,N_25116,N_25345);
and U26935 (N_26935,N_25449,N_25346);
or U26936 (N_26936,N_25708,N_25427);
and U26937 (N_26937,N_25564,N_25402);
xor U26938 (N_26938,N_25287,N_25753);
nor U26939 (N_26939,N_25597,N_25791);
nand U26940 (N_26940,N_25695,N_25497);
or U26941 (N_26941,N_25694,N_25302);
or U26942 (N_26942,N_25435,N_25189);
nand U26943 (N_26943,N_25543,N_25583);
or U26944 (N_26944,N_25793,N_25760);
nor U26945 (N_26945,N_25646,N_25012);
xnor U26946 (N_26946,N_25996,N_25588);
nor U26947 (N_26947,N_25802,N_25006);
nor U26948 (N_26948,N_25570,N_25083);
xor U26949 (N_26949,N_25929,N_25180);
or U26950 (N_26950,N_25478,N_25415);
nor U26951 (N_26951,N_25220,N_25319);
nand U26952 (N_26952,N_25434,N_25124);
and U26953 (N_26953,N_25849,N_25652);
or U26954 (N_26954,N_25795,N_25158);
nor U26955 (N_26955,N_25682,N_25243);
and U26956 (N_26956,N_25950,N_25025);
and U26957 (N_26957,N_25860,N_25025);
nand U26958 (N_26958,N_25045,N_25892);
nor U26959 (N_26959,N_25968,N_25928);
nand U26960 (N_26960,N_25022,N_25866);
and U26961 (N_26961,N_25790,N_25478);
and U26962 (N_26962,N_25009,N_25250);
nor U26963 (N_26963,N_25345,N_25512);
or U26964 (N_26964,N_25720,N_25616);
and U26965 (N_26965,N_25935,N_25178);
nand U26966 (N_26966,N_25158,N_25130);
and U26967 (N_26967,N_25836,N_25767);
and U26968 (N_26968,N_25322,N_25488);
nand U26969 (N_26969,N_25962,N_25810);
nand U26970 (N_26970,N_25876,N_25380);
nand U26971 (N_26971,N_25208,N_25706);
or U26972 (N_26972,N_25096,N_25725);
and U26973 (N_26973,N_25166,N_25523);
and U26974 (N_26974,N_25906,N_25061);
xor U26975 (N_26975,N_25756,N_25176);
nand U26976 (N_26976,N_25159,N_25504);
nand U26977 (N_26977,N_25807,N_25458);
xnor U26978 (N_26978,N_25990,N_25210);
nor U26979 (N_26979,N_25643,N_25264);
xor U26980 (N_26980,N_25627,N_25085);
nand U26981 (N_26981,N_25060,N_25571);
or U26982 (N_26982,N_25944,N_25617);
nor U26983 (N_26983,N_25739,N_25854);
and U26984 (N_26984,N_25168,N_25292);
or U26985 (N_26985,N_25356,N_25968);
nor U26986 (N_26986,N_25382,N_25232);
nor U26987 (N_26987,N_25383,N_25489);
nor U26988 (N_26988,N_25249,N_25355);
nand U26989 (N_26989,N_25318,N_25822);
and U26990 (N_26990,N_25072,N_25809);
or U26991 (N_26991,N_25343,N_25152);
and U26992 (N_26992,N_25389,N_25767);
nor U26993 (N_26993,N_25714,N_25650);
nor U26994 (N_26994,N_25382,N_25845);
nand U26995 (N_26995,N_25853,N_25626);
and U26996 (N_26996,N_25432,N_25990);
or U26997 (N_26997,N_25474,N_25326);
nand U26998 (N_26998,N_25890,N_25373);
and U26999 (N_26999,N_25037,N_25127);
nand U27000 (N_27000,N_26988,N_26501);
and U27001 (N_27001,N_26483,N_26980);
nand U27002 (N_27002,N_26920,N_26470);
nor U27003 (N_27003,N_26826,N_26599);
xnor U27004 (N_27004,N_26236,N_26156);
and U27005 (N_27005,N_26247,N_26185);
nand U27006 (N_27006,N_26541,N_26543);
or U27007 (N_27007,N_26564,N_26100);
nand U27008 (N_27008,N_26024,N_26155);
and U27009 (N_27009,N_26556,N_26021);
xnor U27010 (N_27010,N_26636,N_26510);
nor U27011 (N_27011,N_26002,N_26647);
nand U27012 (N_27012,N_26915,N_26336);
nand U27013 (N_27013,N_26232,N_26057);
and U27014 (N_27014,N_26911,N_26596);
and U27015 (N_27015,N_26567,N_26088);
nand U27016 (N_27016,N_26951,N_26216);
or U27017 (N_27017,N_26699,N_26745);
or U27018 (N_27018,N_26984,N_26262);
nor U27019 (N_27019,N_26866,N_26391);
or U27020 (N_27020,N_26311,N_26707);
nand U27021 (N_27021,N_26508,N_26622);
nand U27022 (N_27022,N_26509,N_26977);
xnor U27023 (N_27023,N_26926,N_26670);
nand U27024 (N_27024,N_26740,N_26825);
and U27025 (N_27025,N_26069,N_26097);
xnor U27026 (N_27026,N_26293,N_26288);
and U27027 (N_27027,N_26186,N_26080);
and U27028 (N_27028,N_26929,N_26179);
or U27029 (N_27029,N_26150,N_26368);
xor U27030 (N_27030,N_26018,N_26862);
or U27031 (N_27031,N_26865,N_26890);
or U27032 (N_27032,N_26772,N_26015);
xor U27033 (N_27033,N_26377,N_26595);
nand U27034 (N_27034,N_26456,N_26779);
xor U27035 (N_27035,N_26671,N_26655);
or U27036 (N_27036,N_26346,N_26974);
nand U27037 (N_27037,N_26691,N_26847);
nand U27038 (N_27038,N_26507,N_26545);
nor U27039 (N_27039,N_26152,N_26652);
nor U27040 (N_27040,N_26738,N_26721);
nand U27041 (N_27041,N_26889,N_26759);
and U27042 (N_27042,N_26003,N_26171);
xor U27043 (N_27043,N_26276,N_26560);
or U27044 (N_27044,N_26375,N_26489);
xnor U27045 (N_27045,N_26552,N_26601);
nor U27046 (N_27046,N_26522,N_26815);
and U27047 (N_27047,N_26408,N_26918);
nand U27048 (N_27048,N_26258,N_26220);
xnor U27049 (N_27049,N_26893,N_26341);
or U27050 (N_27050,N_26925,N_26625);
and U27051 (N_27051,N_26923,N_26876);
nand U27052 (N_27052,N_26644,N_26400);
nor U27053 (N_27053,N_26267,N_26513);
xnor U27054 (N_27054,N_26874,N_26036);
xnor U27055 (N_27055,N_26044,N_26598);
and U27056 (N_27056,N_26557,N_26591);
xnor U27057 (N_27057,N_26761,N_26909);
nor U27058 (N_27058,N_26942,N_26366);
and U27059 (N_27059,N_26307,N_26189);
or U27060 (N_27060,N_26586,N_26621);
nor U27061 (N_27061,N_26175,N_26032);
nor U27062 (N_27062,N_26529,N_26861);
nand U27063 (N_27063,N_26637,N_26853);
nand U27064 (N_27064,N_26047,N_26756);
nand U27065 (N_27065,N_26705,N_26284);
xnor U27066 (N_27066,N_26187,N_26758);
xor U27067 (N_27067,N_26025,N_26246);
or U27068 (N_27068,N_26558,N_26157);
or U27069 (N_27069,N_26813,N_26023);
and U27070 (N_27070,N_26308,N_26103);
nand U27071 (N_27071,N_26950,N_26627);
nand U27072 (N_27072,N_26544,N_26206);
or U27073 (N_27073,N_26662,N_26766);
nand U27074 (N_27074,N_26070,N_26616);
xnor U27075 (N_27075,N_26362,N_26213);
xor U27076 (N_27076,N_26335,N_26374);
xnor U27077 (N_27077,N_26703,N_26131);
xor U27078 (N_27078,N_26450,N_26797);
nand U27079 (N_27079,N_26860,N_26342);
and U27080 (N_27080,N_26357,N_26237);
or U27081 (N_27081,N_26729,N_26141);
and U27082 (N_27082,N_26697,N_26611);
or U27083 (N_27083,N_26981,N_26111);
xor U27084 (N_27084,N_26623,N_26325);
nand U27085 (N_27085,N_26498,N_26146);
and U27086 (N_27086,N_26294,N_26251);
xnor U27087 (N_27087,N_26676,N_26050);
and U27088 (N_27088,N_26843,N_26663);
and U27089 (N_27089,N_26201,N_26245);
and U27090 (N_27090,N_26573,N_26228);
and U27091 (N_27091,N_26653,N_26741);
and U27092 (N_27092,N_26323,N_26020);
and U27093 (N_27093,N_26686,N_26566);
nor U27094 (N_27094,N_26300,N_26226);
nand U27095 (N_27095,N_26109,N_26240);
and U27096 (N_27096,N_26776,N_26736);
and U27097 (N_27097,N_26737,N_26711);
nor U27098 (N_27098,N_26429,N_26099);
xnor U27099 (N_27099,N_26638,N_26927);
nor U27100 (N_27100,N_26762,N_26607);
xor U27101 (N_27101,N_26409,N_26278);
or U27102 (N_27102,N_26993,N_26079);
nand U27103 (N_27103,N_26718,N_26301);
nand U27104 (N_27104,N_26775,N_26931);
xnor U27105 (N_27105,N_26561,N_26954);
and U27106 (N_27106,N_26190,N_26854);
or U27107 (N_27107,N_26844,N_26334);
nand U27108 (N_27108,N_26913,N_26401);
and U27109 (N_27109,N_26272,N_26493);
nor U27110 (N_27110,N_26807,N_26613);
or U27111 (N_27111,N_26863,N_26143);
or U27112 (N_27112,N_26778,N_26525);
xor U27113 (N_27113,N_26244,N_26932);
xnor U27114 (N_27114,N_26581,N_26518);
or U27115 (N_27115,N_26387,N_26753);
xor U27116 (N_27116,N_26577,N_26667);
nor U27117 (N_27117,N_26310,N_26597);
or U27118 (N_27118,N_26348,N_26687);
and U27119 (N_27119,N_26063,N_26678);
or U27120 (N_27120,N_26534,N_26484);
or U27121 (N_27121,N_26469,N_26081);
or U27122 (N_27122,N_26857,N_26649);
nand U27123 (N_27123,N_26682,N_26809);
or U27124 (N_27124,N_26971,N_26114);
xor U27125 (N_27125,N_26196,N_26041);
nor U27126 (N_27126,N_26646,N_26167);
xor U27127 (N_27127,N_26757,N_26821);
xor U27128 (N_27128,N_26702,N_26879);
nor U27129 (N_27129,N_26433,N_26046);
nor U27130 (N_27130,N_26065,N_26116);
or U27131 (N_27131,N_26316,N_26264);
nand U27132 (N_27132,N_26356,N_26282);
xor U27133 (N_27133,N_26716,N_26012);
and U27134 (N_27134,N_26209,N_26136);
or U27135 (N_27135,N_26767,N_26856);
xor U27136 (N_27136,N_26125,N_26651);
and U27137 (N_27137,N_26976,N_26940);
or U27138 (N_27138,N_26416,N_26239);
and U27139 (N_27139,N_26811,N_26227);
xnor U27140 (N_27140,N_26569,N_26936);
and U27141 (N_27141,N_26692,N_26679);
or U27142 (N_27142,N_26871,N_26841);
nand U27143 (N_27143,N_26121,N_26720);
nor U27144 (N_27144,N_26268,N_26314);
nand U27145 (N_27145,N_26881,N_26445);
and U27146 (N_27146,N_26796,N_26690);
or U27147 (N_27147,N_26004,N_26326);
nand U27148 (N_27148,N_26838,N_26331);
xor U27149 (N_27149,N_26748,N_26882);
xnor U27150 (N_27150,N_26091,N_26726);
xnor U27151 (N_27151,N_26304,N_26398);
or U27152 (N_27152,N_26798,N_26168);
xnor U27153 (N_27153,N_26299,N_26605);
or U27154 (N_27154,N_26447,N_26941);
nand U27155 (N_27155,N_26760,N_26263);
xnor U27156 (N_27156,N_26033,N_26176);
and U27157 (N_27157,N_26804,N_26805);
and U27158 (N_27158,N_26768,N_26831);
or U27159 (N_27159,N_26568,N_26207);
nor U27160 (N_27160,N_26743,N_26092);
nand U27161 (N_27161,N_26312,N_26824);
and U27162 (N_27162,N_26291,N_26473);
or U27163 (N_27163,N_26137,N_26793);
xnor U27164 (N_27164,N_26640,N_26438);
and U27165 (N_27165,N_26947,N_26580);
nand U27166 (N_27166,N_26269,N_26823);
nor U27167 (N_27167,N_26719,N_26480);
or U27168 (N_27168,N_26204,N_26203);
and U27169 (N_27169,N_26419,N_26275);
xnor U27170 (N_27170,N_26995,N_26769);
nor U27171 (N_27171,N_26631,N_26231);
xor U27172 (N_27172,N_26223,N_26487);
or U27173 (N_27173,N_26446,N_26290);
or U27174 (N_27174,N_26837,N_26836);
and U27175 (N_27175,N_26351,N_26074);
or U27176 (N_27176,N_26472,N_26297);
nand U27177 (N_27177,N_26818,N_26695);
nor U27178 (N_27178,N_26389,N_26814);
xor U27179 (N_27179,N_26358,N_26076);
and U27180 (N_27180,N_26192,N_26392);
nor U27181 (N_27181,N_26867,N_26332);
nand U27182 (N_27182,N_26765,N_26619);
nor U27183 (N_27183,N_26735,N_26642);
xnor U27184 (N_27184,N_26089,N_26124);
nor U27185 (N_27185,N_26829,N_26585);
and U27186 (N_27186,N_26043,N_26313);
nand U27187 (N_27187,N_26465,N_26259);
nor U27188 (N_27188,N_26490,N_26485);
and U27189 (N_27189,N_26017,N_26248);
and U27190 (N_27190,N_26296,N_26547);
or U27191 (N_27191,N_26364,N_26958);
or U27192 (N_27192,N_26660,N_26181);
nand U27193 (N_27193,N_26848,N_26395);
xnor U27194 (N_27194,N_26164,N_26031);
nor U27195 (N_27195,N_26051,N_26714);
and U27196 (N_27196,N_26126,N_26462);
or U27197 (N_27197,N_26086,N_26318);
xnor U27198 (N_27198,N_26333,N_26969);
and U27199 (N_27199,N_26302,N_26008);
nor U27200 (N_27200,N_26900,N_26777);
xor U27201 (N_27201,N_26540,N_26306);
xor U27202 (N_27202,N_26992,N_26799);
nand U27203 (N_27203,N_26424,N_26466);
xor U27204 (N_27204,N_26693,N_26014);
xnor U27205 (N_27205,N_26180,N_26576);
xor U27206 (N_27206,N_26688,N_26503);
xnor U27207 (N_27207,N_26412,N_26098);
or U27208 (N_27208,N_26430,N_26083);
nor U27209 (N_27209,N_26666,N_26790);
nor U27210 (N_27210,N_26355,N_26471);
or U27211 (N_27211,N_26635,N_26755);
nor U27212 (N_27212,N_26872,N_26914);
nor U27213 (N_27213,N_26037,N_26094);
or U27214 (N_27214,N_26795,N_26511);
or U27215 (N_27215,N_26764,N_26905);
nor U27216 (N_27216,N_26674,N_26460);
or U27217 (N_27217,N_26329,N_26855);
or U27218 (N_27218,N_26968,N_26040);
nor U27219 (N_27219,N_26614,N_26440);
xor U27220 (N_27220,N_26153,N_26084);
nand U27221 (N_27221,N_26917,N_26172);
nand U27222 (N_27222,N_26801,N_26096);
nand U27223 (N_27223,N_26641,N_26535);
nor U27224 (N_27224,N_26139,N_26000);
and U27225 (N_27225,N_26413,N_26059);
nor U27226 (N_27226,N_26110,N_26191);
xnor U27227 (N_27227,N_26056,N_26594);
and U27228 (N_27228,N_26461,N_26868);
and U27229 (N_27229,N_26160,N_26448);
nand U27230 (N_27230,N_26533,N_26378);
nor U27231 (N_27231,N_26255,N_26746);
and U27232 (N_27232,N_26235,N_26588);
and U27233 (N_27233,N_26376,N_26903);
nand U27234 (N_27234,N_26145,N_26944);
xor U27235 (N_27235,N_26928,N_26028);
nor U27236 (N_27236,N_26022,N_26620);
xnor U27237 (N_27237,N_26733,N_26270);
or U27238 (N_27238,N_26612,N_26706);
nor U27239 (N_27239,N_26698,N_26986);
or U27240 (N_27240,N_26794,N_26933);
nor U27241 (N_27241,N_26658,N_26385);
xnor U27242 (N_27242,N_26962,N_26921);
xor U27243 (N_27243,N_26787,N_26846);
nand U27244 (N_27244,N_26132,N_26873);
nand U27245 (N_27245,N_26791,N_26849);
nor U27246 (N_27246,N_26967,N_26442);
and U27247 (N_27247,N_26060,N_26820);
nor U27248 (N_27248,N_26633,N_26402);
and U27249 (N_27249,N_26935,N_26118);
and U27250 (N_27250,N_26709,N_26839);
nor U27251 (N_27251,N_26987,N_26407);
and U27252 (N_27252,N_26781,N_26500);
nor U27253 (N_27253,N_26423,N_26379);
and U27254 (N_27254,N_26006,N_26959);
nand U27255 (N_27255,N_26208,N_26979);
nand U27256 (N_27256,N_26783,N_26317);
xor U27257 (N_27257,N_26673,N_26369);
nor U27258 (N_27258,N_26010,N_26390);
and U27259 (N_27259,N_26732,N_26531);
or U27260 (N_27260,N_26583,N_26072);
or U27261 (N_27261,N_26277,N_26634);
and U27262 (N_27262,N_26327,N_26380);
xor U27263 (N_27263,N_26650,N_26193);
and U27264 (N_27264,N_26221,N_26101);
and U27265 (N_27265,N_26578,N_26039);
xnor U27266 (N_27266,N_26961,N_26481);
nor U27267 (N_27267,N_26506,N_26038);
xnor U27268 (N_27268,N_26054,N_26253);
or U27269 (N_27269,N_26906,N_26808);
xnor U27270 (N_27270,N_26883,N_26725);
nand U27271 (N_27271,N_26754,N_26800);
or U27272 (N_27272,N_26960,N_26710);
nor U27273 (N_27273,N_26451,N_26242);
nand U27274 (N_27274,N_26212,N_26123);
nand U27275 (N_27275,N_26701,N_26013);
xor U27276 (N_27276,N_26449,N_26426);
or U27277 (N_27277,N_26249,N_26455);
nand U27278 (N_27278,N_26624,N_26712);
or U27279 (N_27279,N_26989,N_26052);
nand U27280 (N_27280,N_26514,N_26045);
nand U27281 (N_27281,N_26049,N_26908);
nor U27282 (N_27282,N_26144,N_26538);
and U27283 (N_27283,N_26422,N_26488);
nor U27284 (N_27284,N_26352,N_26222);
or U27285 (N_27285,N_26108,N_26298);
xor U27286 (N_27286,N_26532,N_26238);
or U27287 (N_27287,N_26105,N_26322);
or U27288 (N_27288,N_26421,N_26388);
and U27289 (N_27289,N_26990,N_26668);
nand U27290 (N_27290,N_26496,N_26007);
xnor U27291 (N_27291,N_26945,N_26563);
or U27292 (N_27292,N_26998,N_26361);
nand U27293 (N_27293,N_26792,N_26806);
nand U27294 (N_27294,N_26632,N_26555);
or U27295 (N_27295,N_26648,N_26340);
xor U27296 (N_27296,N_26420,N_26656);
xor U27297 (N_27297,N_26425,N_26183);
and U27298 (N_27298,N_26159,N_26486);
xnor U27299 (N_27299,N_26482,N_26360);
and U27300 (N_27300,N_26075,N_26305);
nor U27301 (N_27301,N_26696,N_26082);
nand U27302 (N_27302,N_26770,N_26205);
nand U27303 (N_27303,N_26494,N_26924);
or U27304 (N_27304,N_26292,N_26188);
nand U27305 (N_27305,N_26224,N_26888);
or U27306 (N_27306,N_26816,N_26537);
nor U27307 (N_27307,N_26898,N_26948);
xnor U27308 (N_27308,N_26734,N_26521);
nor U27309 (N_27309,N_26571,N_26093);
xnor U27310 (N_27310,N_26752,N_26835);
and U27311 (N_27311,N_26279,N_26523);
and U27312 (N_27312,N_26274,N_26606);
and U27313 (N_27313,N_26468,N_26102);
or U27314 (N_27314,N_26542,N_26479);
nor U27315 (N_27315,N_26463,N_26672);
nor U27316 (N_27316,N_26475,N_26151);
or U27317 (N_27317,N_26464,N_26694);
nor U27318 (N_27318,N_26880,N_26243);
and U27319 (N_27319,N_26704,N_26418);
and U27320 (N_27320,N_26902,N_26178);
nand U27321 (N_27321,N_26444,N_26830);
nand U27322 (N_27322,N_26546,N_26684);
and U27323 (N_27323,N_26347,N_26283);
nor U27324 (N_27324,N_26127,N_26428);
nand U27325 (N_27325,N_26603,N_26727);
or U27326 (N_27326,N_26982,N_26700);
nand U27327 (N_27327,N_26436,N_26587);
nand U27328 (N_27328,N_26628,N_26104);
nor U27329 (N_27329,N_26949,N_26901);
xor U27330 (N_27330,N_26604,N_26415);
xnor U27331 (N_27331,N_26128,N_26570);
or U27332 (N_27332,N_26536,N_26345);
nand U27333 (N_27333,N_26367,N_26885);
and U27334 (N_27334,N_26910,N_26878);
and U27335 (N_27335,N_26439,N_26774);
xor U27336 (N_27336,N_26520,N_26359);
xnor U27337 (N_27337,N_26530,N_26952);
nand U27338 (N_27338,N_26399,N_26955);
and U27339 (N_27339,N_26802,N_26973);
xor U27340 (N_27340,N_26256,N_26930);
and U27341 (N_27341,N_26747,N_26182);
or U27342 (N_27342,N_26851,N_26551);
and U27343 (N_27343,N_26233,N_26845);
nor U27344 (N_27344,N_26659,N_26053);
xor U27345 (N_27345,N_26163,N_26285);
nand U27346 (N_27346,N_26202,N_26579);
nor U27347 (N_27347,N_26115,N_26840);
nand U27348 (N_27348,N_26966,N_26061);
nor U27349 (N_27349,N_26281,N_26991);
or U27350 (N_27350,N_26617,N_26645);
nor U27351 (N_27351,N_26295,N_26739);
nand U27352 (N_27352,N_26922,N_26750);
and U27353 (N_27353,N_26372,N_26934);
and U27354 (N_27354,N_26731,N_26884);
or U27355 (N_27355,N_26225,N_26610);
nor U27356 (N_27356,N_26199,N_26161);
or U27357 (N_27357,N_26230,N_26997);
nor U27358 (N_27358,N_26904,N_26504);
or U27359 (N_27359,N_26963,N_26441);
nor U27360 (N_27360,N_26215,N_26943);
and U27361 (N_27361,N_26035,N_26273);
or U27362 (N_27362,N_26027,N_26505);
and U27363 (N_27363,N_26058,N_26713);
or U27364 (N_27364,N_26894,N_26034);
xnor U27365 (N_27365,N_26639,N_26589);
xor U27366 (N_27366,N_26497,N_26026);
and U27367 (N_27367,N_26454,N_26550);
nor U27368 (N_27368,N_26875,N_26217);
nor U27369 (N_27369,N_26174,N_26383);
xnor U27370 (N_27370,N_26452,N_26728);
or U27371 (N_27371,N_26817,N_26887);
nor U27372 (N_27372,N_26122,N_26066);
nand U27373 (N_27373,N_26763,N_26320);
xnor U27374 (N_27374,N_26062,N_26938);
nor U27375 (N_27375,N_26474,N_26194);
or U27376 (N_27376,N_26397,N_26528);
and U27377 (N_27377,N_26953,N_26129);
and U27378 (N_27378,N_26675,N_26477);
xnor U27379 (N_27379,N_26077,N_26009);
nor U27380 (N_27380,N_26499,N_26553);
or U27381 (N_27381,N_26458,N_26029);
xor U27382 (N_27382,N_26615,N_26590);
xor U27383 (N_27383,N_26211,N_26661);
nand U27384 (N_27384,N_26437,N_26715);
or U27385 (N_27385,N_26166,N_26373);
nor U27386 (N_27386,N_26434,N_26120);
xor U27387 (N_27387,N_26257,N_26751);
nor U27388 (N_27388,N_26669,N_26095);
nor U27389 (N_27389,N_26722,N_26549);
xnor U27390 (N_27390,N_26173,N_26749);
xor U27391 (N_27391,N_26148,N_26218);
nand U27392 (N_27392,N_26177,N_26978);
nand U27393 (N_27393,N_26337,N_26386);
nand U27394 (N_27394,N_26353,N_26832);
or U27395 (N_27395,N_26384,N_26067);
and U27396 (N_27396,N_26459,N_26999);
nand U27397 (N_27397,N_26030,N_26453);
xor U27398 (N_27398,N_26019,N_26572);
nor U27399 (N_27399,N_26287,N_26261);
or U27400 (N_27400,N_26309,N_26524);
and U27401 (N_27401,N_26005,N_26833);
or U27402 (N_27402,N_26562,N_26254);
xnor U27403 (N_27403,N_26085,N_26071);
xnor U27404 (N_27404,N_26575,N_26939);
or U27405 (N_27405,N_26492,N_26803);
nor U27406 (N_27406,N_26162,N_26229);
nor U27407 (N_27407,N_26609,N_26600);
and U27408 (N_27408,N_26957,N_26970);
nor U27409 (N_27409,N_26068,N_26677);
nor U27410 (N_27410,N_26548,N_26565);
or U27411 (N_27411,N_26554,N_26516);
and U27412 (N_27412,N_26393,N_26476);
xor U27413 (N_27413,N_26512,N_26330);
nand U27414 (N_27414,N_26519,N_26850);
or U27415 (N_27415,N_26365,N_26912);
nand U27416 (N_27416,N_26324,N_26996);
nor U27417 (N_27417,N_26349,N_26048);
or U27418 (N_27418,N_26877,N_26994);
or U27419 (N_27419,N_26983,N_26394);
or U27420 (N_27420,N_26789,N_26526);
and U27421 (N_27421,N_26819,N_26895);
and U27422 (N_27422,N_26133,N_26574);
and U27423 (N_27423,N_26252,N_26234);
or U27424 (N_27424,N_26630,N_26657);
nor U27425 (N_27425,N_26897,N_26319);
or U27426 (N_27426,N_26812,N_26042);
and U27427 (N_27427,N_26689,N_26404);
nand U27428 (N_27428,N_26681,N_26055);
nand U27429 (N_27429,N_26654,N_26073);
or U27430 (N_27430,N_26250,N_26643);
xor U27431 (N_27431,N_26016,N_26158);
and U27432 (N_27432,N_26381,N_26142);
and U27433 (N_27433,N_26064,N_26289);
and U27434 (N_27434,N_26834,N_26457);
nor U27435 (N_27435,N_26328,N_26169);
nor U27436 (N_27436,N_26892,N_26975);
nand U27437 (N_27437,N_26350,N_26896);
xnor U27438 (N_27438,N_26785,N_26478);
xor U27439 (N_27439,N_26708,N_26828);
nor U27440 (N_27440,N_26937,N_26406);
nand U27441 (N_27441,N_26559,N_26403);
nor U27442 (N_27442,N_26431,N_26371);
or U27443 (N_27443,N_26899,N_26343);
and U27444 (N_27444,N_26265,N_26112);
or U27445 (N_27445,N_26810,N_26827);
xor U27446 (N_27446,N_26730,N_26214);
xor U27447 (N_27447,N_26724,N_26864);
nor U27448 (N_27448,N_26539,N_26138);
and U27449 (N_27449,N_26411,N_26443);
xor U27450 (N_27450,N_26629,N_26417);
nand U27451 (N_27451,N_26134,N_26321);
or U27452 (N_27452,N_26985,N_26087);
nor U27453 (N_27453,N_26717,N_26593);
and U27454 (N_27454,N_26260,N_26200);
nand U27455 (N_27455,N_26135,N_26432);
nand U27456 (N_27456,N_26130,N_26410);
xor U27457 (N_27457,N_26964,N_26241);
nor U27458 (N_27458,N_26107,N_26842);
and U27459 (N_27459,N_26266,N_26147);
and U27460 (N_27460,N_26370,N_26382);
xor U27461 (N_27461,N_26584,N_26723);
or U27462 (N_27462,N_26315,N_26858);
nand U27463 (N_27463,N_26685,N_26197);
xnor U27464 (N_27464,N_26665,N_26618);
and U27465 (N_27465,N_26435,N_26001);
xnor U27466 (N_27466,N_26149,N_26592);
and U27467 (N_27467,N_26582,N_26916);
xnor U27468 (N_27468,N_26427,N_26919);
nor U27469 (N_27469,N_26680,N_26602);
and U27470 (N_27470,N_26852,N_26744);
or U27471 (N_27471,N_26011,N_26782);
and U27472 (N_27472,N_26788,N_26414);
nand U27473 (N_27473,N_26078,N_26405);
or U27474 (N_27474,N_26467,N_26219);
or U27475 (N_27475,N_26396,N_26784);
nand U27476 (N_27476,N_26338,N_26527);
nand U27477 (N_27477,N_26113,N_26170);
or U27478 (N_27478,N_26870,N_26117);
nand U27479 (N_27479,N_26491,N_26742);
nor U27480 (N_27480,N_26090,N_26140);
or U27481 (N_27481,N_26515,N_26869);
nand U27482 (N_27482,N_26859,N_26303);
nor U27483 (N_27483,N_26198,N_26956);
xnor U27484 (N_27484,N_26354,N_26771);
xor U27485 (N_27485,N_26683,N_26271);
and U27486 (N_27486,N_26786,N_26626);
xnor U27487 (N_27487,N_26154,N_26195);
nand U27488 (N_27488,N_26119,N_26946);
xor U27489 (N_27489,N_26907,N_26608);
nor U27490 (N_27490,N_26773,N_26184);
nand U27491 (N_27491,N_26822,N_26363);
and U27492 (N_27492,N_26210,N_26517);
or U27493 (N_27493,N_26339,N_26664);
and U27494 (N_27494,N_26344,N_26972);
and U27495 (N_27495,N_26965,N_26502);
and U27496 (N_27496,N_26780,N_26891);
nor U27497 (N_27497,N_26165,N_26886);
nand U27498 (N_27498,N_26286,N_26280);
xor U27499 (N_27499,N_26106,N_26495);
nor U27500 (N_27500,N_26522,N_26833);
and U27501 (N_27501,N_26851,N_26946);
xor U27502 (N_27502,N_26896,N_26765);
nor U27503 (N_27503,N_26476,N_26412);
and U27504 (N_27504,N_26942,N_26855);
and U27505 (N_27505,N_26699,N_26320);
or U27506 (N_27506,N_26791,N_26271);
and U27507 (N_27507,N_26514,N_26220);
nor U27508 (N_27508,N_26739,N_26595);
xor U27509 (N_27509,N_26661,N_26672);
nand U27510 (N_27510,N_26587,N_26482);
nand U27511 (N_27511,N_26413,N_26942);
and U27512 (N_27512,N_26557,N_26577);
or U27513 (N_27513,N_26262,N_26300);
xor U27514 (N_27514,N_26338,N_26271);
and U27515 (N_27515,N_26070,N_26453);
nand U27516 (N_27516,N_26645,N_26584);
nand U27517 (N_27517,N_26020,N_26699);
xor U27518 (N_27518,N_26898,N_26498);
nor U27519 (N_27519,N_26801,N_26020);
or U27520 (N_27520,N_26864,N_26157);
and U27521 (N_27521,N_26333,N_26122);
or U27522 (N_27522,N_26847,N_26032);
xnor U27523 (N_27523,N_26816,N_26572);
xor U27524 (N_27524,N_26501,N_26945);
nor U27525 (N_27525,N_26114,N_26186);
and U27526 (N_27526,N_26443,N_26740);
nor U27527 (N_27527,N_26825,N_26332);
or U27528 (N_27528,N_26187,N_26042);
nand U27529 (N_27529,N_26804,N_26083);
xor U27530 (N_27530,N_26622,N_26954);
xor U27531 (N_27531,N_26283,N_26052);
or U27532 (N_27532,N_26759,N_26832);
and U27533 (N_27533,N_26981,N_26939);
nand U27534 (N_27534,N_26739,N_26320);
nand U27535 (N_27535,N_26723,N_26265);
and U27536 (N_27536,N_26791,N_26759);
and U27537 (N_27537,N_26493,N_26461);
xor U27538 (N_27538,N_26615,N_26394);
nor U27539 (N_27539,N_26913,N_26091);
or U27540 (N_27540,N_26093,N_26190);
or U27541 (N_27541,N_26648,N_26239);
and U27542 (N_27542,N_26639,N_26823);
or U27543 (N_27543,N_26633,N_26488);
and U27544 (N_27544,N_26853,N_26105);
nand U27545 (N_27545,N_26017,N_26007);
and U27546 (N_27546,N_26233,N_26839);
nand U27547 (N_27547,N_26639,N_26213);
and U27548 (N_27548,N_26503,N_26145);
or U27549 (N_27549,N_26659,N_26327);
or U27550 (N_27550,N_26057,N_26952);
or U27551 (N_27551,N_26785,N_26763);
and U27552 (N_27552,N_26193,N_26146);
and U27553 (N_27553,N_26152,N_26499);
nand U27554 (N_27554,N_26775,N_26739);
xnor U27555 (N_27555,N_26874,N_26117);
and U27556 (N_27556,N_26132,N_26994);
and U27557 (N_27557,N_26382,N_26158);
or U27558 (N_27558,N_26189,N_26553);
nor U27559 (N_27559,N_26530,N_26584);
and U27560 (N_27560,N_26740,N_26078);
nor U27561 (N_27561,N_26065,N_26689);
nand U27562 (N_27562,N_26707,N_26988);
nor U27563 (N_27563,N_26559,N_26175);
or U27564 (N_27564,N_26952,N_26892);
or U27565 (N_27565,N_26826,N_26255);
xnor U27566 (N_27566,N_26405,N_26963);
or U27567 (N_27567,N_26179,N_26977);
xor U27568 (N_27568,N_26778,N_26749);
xnor U27569 (N_27569,N_26301,N_26062);
and U27570 (N_27570,N_26481,N_26789);
nand U27571 (N_27571,N_26901,N_26096);
nand U27572 (N_27572,N_26529,N_26203);
and U27573 (N_27573,N_26176,N_26334);
nand U27574 (N_27574,N_26583,N_26887);
nor U27575 (N_27575,N_26538,N_26160);
xnor U27576 (N_27576,N_26771,N_26074);
and U27577 (N_27577,N_26229,N_26242);
and U27578 (N_27578,N_26270,N_26902);
nor U27579 (N_27579,N_26825,N_26209);
nor U27580 (N_27580,N_26845,N_26459);
nor U27581 (N_27581,N_26547,N_26233);
nand U27582 (N_27582,N_26214,N_26086);
and U27583 (N_27583,N_26608,N_26103);
or U27584 (N_27584,N_26695,N_26899);
nand U27585 (N_27585,N_26485,N_26314);
xor U27586 (N_27586,N_26052,N_26273);
or U27587 (N_27587,N_26286,N_26363);
nor U27588 (N_27588,N_26118,N_26087);
nand U27589 (N_27589,N_26502,N_26058);
xnor U27590 (N_27590,N_26662,N_26191);
xor U27591 (N_27591,N_26882,N_26518);
nand U27592 (N_27592,N_26828,N_26148);
nand U27593 (N_27593,N_26573,N_26999);
nand U27594 (N_27594,N_26649,N_26219);
or U27595 (N_27595,N_26776,N_26519);
or U27596 (N_27596,N_26343,N_26336);
and U27597 (N_27597,N_26727,N_26378);
nand U27598 (N_27598,N_26102,N_26611);
nor U27599 (N_27599,N_26697,N_26111);
and U27600 (N_27600,N_26193,N_26758);
xnor U27601 (N_27601,N_26477,N_26108);
or U27602 (N_27602,N_26254,N_26946);
nand U27603 (N_27603,N_26150,N_26389);
or U27604 (N_27604,N_26492,N_26822);
and U27605 (N_27605,N_26145,N_26459);
or U27606 (N_27606,N_26726,N_26071);
or U27607 (N_27607,N_26245,N_26569);
and U27608 (N_27608,N_26847,N_26089);
xnor U27609 (N_27609,N_26272,N_26037);
xor U27610 (N_27610,N_26957,N_26611);
nand U27611 (N_27611,N_26726,N_26834);
and U27612 (N_27612,N_26559,N_26005);
nor U27613 (N_27613,N_26513,N_26617);
or U27614 (N_27614,N_26653,N_26605);
nand U27615 (N_27615,N_26312,N_26639);
or U27616 (N_27616,N_26583,N_26559);
nand U27617 (N_27617,N_26421,N_26987);
nor U27618 (N_27618,N_26777,N_26562);
xnor U27619 (N_27619,N_26668,N_26969);
xor U27620 (N_27620,N_26205,N_26915);
nand U27621 (N_27621,N_26215,N_26419);
nand U27622 (N_27622,N_26453,N_26671);
nand U27623 (N_27623,N_26462,N_26509);
xnor U27624 (N_27624,N_26611,N_26765);
nor U27625 (N_27625,N_26731,N_26624);
nor U27626 (N_27626,N_26935,N_26305);
nand U27627 (N_27627,N_26520,N_26208);
xor U27628 (N_27628,N_26392,N_26855);
nand U27629 (N_27629,N_26417,N_26594);
nand U27630 (N_27630,N_26060,N_26761);
or U27631 (N_27631,N_26123,N_26188);
nand U27632 (N_27632,N_26168,N_26109);
and U27633 (N_27633,N_26952,N_26040);
and U27634 (N_27634,N_26081,N_26345);
xnor U27635 (N_27635,N_26535,N_26755);
and U27636 (N_27636,N_26392,N_26275);
nand U27637 (N_27637,N_26997,N_26028);
nor U27638 (N_27638,N_26191,N_26164);
or U27639 (N_27639,N_26400,N_26072);
nor U27640 (N_27640,N_26324,N_26651);
nor U27641 (N_27641,N_26035,N_26480);
nand U27642 (N_27642,N_26296,N_26074);
nor U27643 (N_27643,N_26693,N_26607);
and U27644 (N_27644,N_26557,N_26649);
and U27645 (N_27645,N_26436,N_26591);
nand U27646 (N_27646,N_26386,N_26654);
xnor U27647 (N_27647,N_26029,N_26666);
or U27648 (N_27648,N_26592,N_26103);
and U27649 (N_27649,N_26207,N_26832);
or U27650 (N_27650,N_26857,N_26275);
and U27651 (N_27651,N_26757,N_26855);
nor U27652 (N_27652,N_26786,N_26286);
and U27653 (N_27653,N_26471,N_26561);
and U27654 (N_27654,N_26196,N_26231);
nand U27655 (N_27655,N_26512,N_26439);
and U27656 (N_27656,N_26830,N_26188);
and U27657 (N_27657,N_26498,N_26921);
or U27658 (N_27658,N_26222,N_26202);
nor U27659 (N_27659,N_26613,N_26437);
nand U27660 (N_27660,N_26591,N_26029);
and U27661 (N_27661,N_26878,N_26323);
nand U27662 (N_27662,N_26154,N_26639);
nand U27663 (N_27663,N_26241,N_26978);
nor U27664 (N_27664,N_26371,N_26959);
nor U27665 (N_27665,N_26926,N_26826);
xnor U27666 (N_27666,N_26242,N_26886);
or U27667 (N_27667,N_26956,N_26324);
and U27668 (N_27668,N_26312,N_26557);
and U27669 (N_27669,N_26878,N_26908);
nand U27670 (N_27670,N_26923,N_26976);
and U27671 (N_27671,N_26068,N_26313);
nand U27672 (N_27672,N_26406,N_26886);
and U27673 (N_27673,N_26606,N_26837);
and U27674 (N_27674,N_26151,N_26764);
and U27675 (N_27675,N_26411,N_26018);
or U27676 (N_27676,N_26443,N_26886);
nor U27677 (N_27677,N_26236,N_26288);
and U27678 (N_27678,N_26727,N_26837);
and U27679 (N_27679,N_26991,N_26633);
nor U27680 (N_27680,N_26542,N_26414);
xnor U27681 (N_27681,N_26716,N_26841);
and U27682 (N_27682,N_26525,N_26463);
nor U27683 (N_27683,N_26586,N_26394);
xor U27684 (N_27684,N_26236,N_26611);
nor U27685 (N_27685,N_26226,N_26235);
nand U27686 (N_27686,N_26465,N_26422);
and U27687 (N_27687,N_26649,N_26759);
nand U27688 (N_27688,N_26035,N_26503);
xor U27689 (N_27689,N_26442,N_26899);
nor U27690 (N_27690,N_26741,N_26809);
or U27691 (N_27691,N_26046,N_26863);
nand U27692 (N_27692,N_26965,N_26074);
nor U27693 (N_27693,N_26013,N_26754);
nand U27694 (N_27694,N_26984,N_26655);
and U27695 (N_27695,N_26059,N_26048);
nor U27696 (N_27696,N_26207,N_26868);
nand U27697 (N_27697,N_26091,N_26775);
xor U27698 (N_27698,N_26322,N_26990);
or U27699 (N_27699,N_26540,N_26546);
and U27700 (N_27700,N_26976,N_26699);
or U27701 (N_27701,N_26374,N_26422);
nor U27702 (N_27702,N_26295,N_26995);
or U27703 (N_27703,N_26102,N_26885);
and U27704 (N_27704,N_26631,N_26237);
nand U27705 (N_27705,N_26806,N_26443);
and U27706 (N_27706,N_26803,N_26414);
nor U27707 (N_27707,N_26299,N_26931);
xor U27708 (N_27708,N_26335,N_26006);
and U27709 (N_27709,N_26579,N_26783);
or U27710 (N_27710,N_26492,N_26165);
nand U27711 (N_27711,N_26012,N_26678);
xnor U27712 (N_27712,N_26315,N_26937);
or U27713 (N_27713,N_26224,N_26428);
nor U27714 (N_27714,N_26443,N_26711);
nand U27715 (N_27715,N_26428,N_26676);
or U27716 (N_27716,N_26064,N_26059);
nand U27717 (N_27717,N_26492,N_26824);
nand U27718 (N_27718,N_26344,N_26613);
or U27719 (N_27719,N_26640,N_26943);
or U27720 (N_27720,N_26587,N_26832);
nand U27721 (N_27721,N_26301,N_26439);
and U27722 (N_27722,N_26570,N_26729);
nor U27723 (N_27723,N_26022,N_26023);
or U27724 (N_27724,N_26291,N_26239);
nand U27725 (N_27725,N_26879,N_26315);
xor U27726 (N_27726,N_26674,N_26908);
or U27727 (N_27727,N_26875,N_26735);
and U27728 (N_27728,N_26101,N_26807);
or U27729 (N_27729,N_26469,N_26434);
nand U27730 (N_27730,N_26999,N_26522);
nand U27731 (N_27731,N_26263,N_26969);
nor U27732 (N_27732,N_26820,N_26068);
or U27733 (N_27733,N_26572,N_26385);
and U27734 (N_27734,N_26860,N_26982);
nand U27735 (N_27735,N_26756,N_26267);
and U27736 (N_27736,N_26063,N_26517);
or U27737 (N_27737,N_26079,N_26789);
nand U27738 (N_27738,N_26643,N_26310);
and U27739 (N_27739,N_26436,N_26291);
nor U27740 (N_27740,N_26914,N_26173);
xor U27741 (N_27741,N_26329,N_26423);
nor U27742 (N_27742,N_26401,N_26567);
or U27743 (N_27743,N_26708,N_26789);
nor U27744 (N_27744,N_26628,N_26378);
xnor U27745 (N_27745,N_26388,N_26051);
and U27746 (N_27746,N_26438,N_26460);
and U27747 (N_27747,N_26515,N_26163);
and U27748 (N_27748,N_26798,N_26306);
nor U27749 (N_27749,N_26495,N_26492);
nor U27750 (N_27750,N_26172,N_26199);
or U27751 (N_27751,N_26664,N_26748);
or U27752 (N_27752,N_26363,N_26103);
and U27753 (N_27753,N_26056,N_26783);
nand U27754 (N_27754,N_26134,N_26653);
nand U27755 (N_27755,N_26834,N_26003);
or U27756 (N_27756,N_26419,N_26703);
nor U27757 (N_27757,N_26738,N_26676);
nor U27758 (N_27758,N_26279,N_26722);
nand U27759 (N_27759,N_26174,N_26338);
and U27760 (N_27760,N_26569,N_26325);
or U27761 (N_27761,N_26417,N_26895);
xor U27762 (N_27762,N_26064,N_26080);
or U27763 (N_27763,N_26137,N_26518);
nor U27764 (N_27764,N_26248,N_26094);
nand U27765 (N_27765,N_26880,N_26595);
nor U27766 (N_27766,N_26990,N_26745);
nor U27767 (N_27767,N_26710,N_26013);
xnor U27768 (N_27768,N_26020,N_26057);
nand U27769 (N_27769,N_26115,N_26985);
nand U27770 (N_27770,N_26728,N_26474);
nor U27771 (N_27771,N_26730,N_26857);
nand U27772 (N_27772,N_26673,N_26385);
or U27773 (N_27773,N_26260,N_26342);
nor U27774 (N_27774,N_26180,N_26678);
or U27775 (N_27775,N_26682,N_26287);
or U27776 (N_27776,N_26801,N_26873);
xor U27777 (N_27777,N_26573,N_26254);
xnor U27778 (N_27778,N_26354,N_26353);
xnor U27779 (N_27779,N_26593,N_26287);
nand U27780 (N_27780,N_26047,N_26860);
nand U27781 (N_27781,N_26983,N_26845);
nor U27782 (N_27782,N_26059,N_26719);
or U27783 (N_27783,N_26806,N_26441);
xor U27784 (N_27784,N_26376,N_26601);
nor U27785 (N_27785,N_26341,N_26361);
and U27786 (N_27786,N_26024,N_26079);
xnor U27787 (N_27787,N_26943,N_26961);
nand U27788 (N_27788,N_26205,N_26737);
and U27789 (N_27789,N_26711,N_26706);
or U27790 (N_27790,N_26944,N_26485);
xnor U27791 (N_27791,N_26545,N_26795);
nand U27792 (N_27792,N_26529,N_26076);
nand U27793 (N_27793,N_26675,N_26240);
nor U27794 (N_27794,N_26014,N_26913);
nor U27795 (N_27795,N_26513,N_26695);
and U27796 (N_27796,N_26032,N_26448);
or U27797 (N_27797,N_26185,N_26275);
and U27798 (N_27798,N_26486,N_26307);
nand U27799 (N_27799,N_26010,N_26387);
and U27800 (N_27800,N_26390,N_26962);
xnor U27801 (N_27801,N_26309,N_26445);
nand U27802 (N_27802,N_26446,N_26495);
and U27803 (N_27803,N_26010,N_26029);
nor U27804 (N_27804,N_26632,N_26219);
xnor U27805 (N_27805,N_26050,N_26140);
nor U27806 (N_27806,N_26700,N_26862);
and U27807 (N_27807,N_26010,N_26208);
nor U27808 (N_27808,N_26228,N_26876);
and U27809 (N_27809,N_26759,N_26119);
xnor U27810 (N_27810,N_26521,N_26940);
nand U27811 (N_27811,N_26153,N_26210);
and U27812 (N_27812,N_26842,N_26325);
nand U27813 (N_27813,N_26542,N_26361);
and U27814 (N_27814,N_26816,N_26057);
nor U27815 (N_27815,N_26342,N_26432);
xnor U27816 (N_27816,N_26903,N_26353);
nand U27817 (N_27817,N_26084,N_26711);
nand U27818 (N_27818,N_26449,N_26605);
and U27819 (N_27819,N_26614,N_26651);
nor U27820 (N_27820,N_26729,N_26105);
nor U27821 (N_27821,N_26103,N_26974);
or U27822 (N_27822,N_26726,N_26933);
and U27823 (N_27823,N_26560,N_26518);
and U27824 (N_27824,N_26601,N_26670);
nor U27825 (N_27825,N_26373,N_26274);
and U27826 (N_27826,N_26975,N_26845);
nor U27827 (N_27827,N_26391,N_26717);
nand U27828 (N_27828,N_26126,N_26192);
and U27829 (N_27829,N_26877,N_26556);
and U27830 (N_27830,N_26637,N_26398);
xnor U27831 (N_27831,N_26591,N_26736);
and U27832 (N_27832,N_26073,N_26243);
or U27833 (N_27833,N_26246,N_26520);
xnor U27834 (N_27834,N_26828,N_26996);
nand U27835 (N_27835,N_26896,N_26667);
nor U27836 (N_27836,N_26903,N_26190);
nor U27837 (N_27837,N_26490,N_26045);
nand U27838 (N_27838,N_26369,N_26516);
or U27839 (N_27839,N_26785,N_26576);
nor U27840 (N_27840,N_26276,N_26700);
and U27841 (N_27841,N_26419,N_26834);
xnor U27842 (N_27842,N_26953,N_26062);
nand U27843 (N_27843,N_26839,N_26910);
and U27844 (N_27844,N_26491,N_26561);
nor U27845 (N_27845,N_26709,N_26061);
nand U27846 (N_27846,N_26973,N_26565);
nor U27847 (N_27847,N_26782,N_26297);
or U27848 (N_27848,N_26158,N_26470);
nand U27849 (N_27849,N_26542,N_26840);
and U27850 (N_27850,N_26315,N_26312);
nand U27851 (N_27851,N_26254,N_26302);
nand U27852 (N_27852,N_26417,N_26982);
or U27853 (N_27853,N_26844,N_26184);
and U27854 (N_27854,N_26225,N_26024);
xnor U27855 (N_27855,N_26466,N_26909);
or U27856 (N_27856,N_26468,N_26594);
nor U27857 (N_27857,N_26196,N_26429);
and U27858 (N_27858,N_26234,N_26603);
nor U27859 (N_27859,N_26028,N_26340);
or U27860 (N_27860,N_26318,N_26803);
nor U27861 (N_27861,N_26237,N_26059);
and U27862 (N_27862,N_26600,N_26514);
nand U27863 (N_27863,N_26319,N_26881);
and U27864 (N_27864,N_26245,N_26947);
and U27865 (N_27865,N_26003,N_26435);
and U27866 (N_27866,N_26776,N_26374);
or U27867 (N_27867,N_26911,N_26811);
and U27868 (N_27868,N_26967,N_26316);
nor U27869 (N_27869,N_26858,N_26331);
nand U27870 (N_27870,N_26017,N_26811);
or U27871 (N_27871,N_26263,N_26576);
or U27872 (N_27872,N_26631,N_26822);
nand U27873 (N_27873,N_26104,N_26085);
or U27874 (N_27874,N_26397,N_26023);
and U27875 (N_27875,N_26168,N_26847);
or U27876 (N_27876,N_26131,N_26732);
nand U27877 (N_27877,N_26801,N_26927);
nor U27878 (N_27878,N_26251,N_26681);
and U27879 (N_27879,N_26598,N_26814);
nand U27880 (N_27880,N_26455,N_26884);
nor U27881 (N_27881,N_26240,N_26900);
xor U27882 (N_27882,N_26378,N_26928);
nor U27883 (N_27883,N_26023,N_26156);
nor U27884 (N_27884,N_26753,N_26659);
nor U27885 (N_27885,N_26200,N_26262);
nor U27886 (N_27886,N_26151,N_26759);
or U27887 (N_27887,N_26560,N_26132);
xor U27888 (N_27888,N_26157,N_26469);
xor U27889 (N_27889,N_26124,N_26275);
nand U27890 (N_27890,N_26111,N_26480);
and U27891 (N_27891,N_26017,N_26603);
nand U27892 (N_27892,N_26974,N_26866);
nor U27893 (N_27893,N_26190,N_26863);
nand U27894 (N_27894,N_26608,N_26138);
xnor U27895 (N_27895,N_26642,N_26224);
and U27896 (N_27896,N_26475,N_26124);
and U27897 (N_27897,N_26192,N_26782);
xnor U27898 (N_27898,N_26116,N_26890);
nor U27899 (N_27899,N_26735,N_26249);
and U27900 (N_27900,N_26224,N_26325);
xnor U27901 (N_27901,N_26185,N_26714);
nor U27902 (N_27902,N_26118,N_26917);
xor U27903 (N_27903,N_26391,N_26515);
xnor U27904 (N_27904,N_26590,N_26577);
xor U27905 (N_27905,N_26546,N_26873);
and U27906 (N_27906,N_26383,N_26354);
and U27907 (N_27907,N_26711,N_26992);
xnor U27908 (N_27908,N_26637,N_26114);
nor U27909 (N_27909,N_26063,N_26543);
and U27910 (N_27910,N_26323,N_26487);
xnor U27911 (N_27911,N_26299,N_26262);
and U27912 (N_27912,N_26491,N_26588);
nand U27913 (N_27913,N_26547,N_26792);
nor U27914 (N_27914,N_26042,N_26465);
xor U27915 (N_27915,N_26955,N_26925);
xor U27916 (N_27916,N_26232,N_26417);
and U27917 (N_27917,N_26145,N_26307);
or U27918 (N_27918,N_26709,N_26520);
nor U27919 (N_27919,N_26693,N_26435);
and U27920 (N_27920,N_26344,N_26600);
or U27921 (N_27921,N_26711,N_26057);
and U27922 (N_27922,N_26954,N_26907);
xnor U27923 (N_27923,N_26321,N_26433);
xor U27924 (N_27924,N_26437,N_26219);
or U27925 (N_27925,N_26142,N_26925);
nor U27926 (N_27926,N_26715,N_26327);
nor U27927 (N_27927,N_26348,N_26312);
and U27928 (N_27928,N_26582,N_26271);
nand U27929 (N_27929,N_26576,N_26332);
nor U27930 (N_27930,N_26090,N_26564);
and U27931 (N_27931,N_26682,N_26594);
and U27932 (N_27932,N_26998,N_26575);
and U27933 (N_27933,N_26459,N_26128);
nand U27934 (N_27934,N_26548,N_26478);
xor U27935 (N_27935,N_26724,N_26941);
or U27936 (N_27936,N_26435,N_26507);
nor U27937 (N_27937,N_26518,N_26936);
nand U27938 (N_27938,N_26304,N_26482);
or U27939 (N_27939,N_26711,N_26355);
nand U27940 (N_27940,N_26918,N_26081);
xor U27941 (N_27941,N_26216,N_26436);
or U27942 (N_27942,N_26097,N_26713);
nor U27943 (N_27943,N_26542,N_26946);
xnor U27944 (N_27944,N_26384,N_26581);
nand U27945 (N_27945,N_26295,N_26498);
nand U27946 (N_27946,N_26454,N_26774);
and U27947 (N_27947,N_26973,N_26545);
or U27948 (N_27948,N_26056,N_26800);
nand U27949 (N_27949,N_26346,N_26299);
nor U27950 (N_27950,N_26953,N_26663);
xor U27951 (N_27951,N_26654,N_26886);
nor U27952 (N_27952,N_26531,N_26703);
or U27953 (N_27953,N_26507,N_26745);
xnor U27954 (N_27954,N_26565,N_26230);
or U27955 (N_27955,N_26500,N_26120);
nor U27956 (N_27956,N_26186,N_26813);
xnor U27957 (N_27957,N_26785,N_26416);
and U27958 (N_27958,N_26286,N_26122);
nor U27959 (N_27959,N_26953,N_26440);
nor U27960 (N_27960,N_26792,N_26278);
nand U27961 (N_27961,N_26264,N_26192);
and U27962 (N_27962,N_26550,N_26325);
nor U27963 (N_27963,N_26395,N_26561);
or U27964 (N_27964,N_26096,N_26390);
and U27965 (N_27965,N_26334,N_26050);
nor U27966 (N_27966,N_26892,N_26288);
nand U27967 (N_27967,N_26837,N_26838);
xnor U27968 (N_27968,N_26012,N_26327);
nand U27969 (N_27969,N_26515,N_26695);
and U27970 (N_27970,N_26659,N_26824);
and U27971 (N_27971,N_26628,N_26201);
xor U27972 (N_27972,N_26943,N_26419);
nand U27973 (N_27973,N_26313,N_26197);
nor U27974 (N_27974,N_26941,N_26413);
nor U27975 (N_27975,N_26451,N_26476);
nor U27976 (N_27976,N_26798,N_26315);
nand U27977 (N_27977,N_26333,N_26847);
xor U27978 (N_27978,N_26817,N_26138);
and U27979 (N_27979,N_26627,N_26030);
xnor U27980 (N_27980,N_26054,N_26582);
xnor U27981 (N_27981,N_26705,N_26922);
and U27982 (N_27982,N_26339,N_26349);
or U27983 (N_27983,N_26075,N_26524);
or U27984 (N_27984,N_26417,N_26471);
xor U27985 (N_27985,N_26656,N_26431);
nand U27986 (N_27986,N_26129,N_26313);
xnor U27987 (N_27987,N_26251,N_26710);
nor U27988 (N_27988,N_26849,N_26568);
and U27989 (N_27989,N_26515,N_26614);
nor U27990 (N_27990,N_26248,N_26357);
or U27991 (N_27991,N_26511,N_26180);
and U27992 (N_27992,N_26801,N_26080);
nand U27993 (N_27993,N_26130,N_26201);
nand U27994 (N_27994,N_26169,N_26758);
xor U27995 (N_27995,N_26861,N_26552);
and U27996 (N_27996,N_26538,N_26823);
nand U27997 (N_27997,N_26680,N_26102);
and U27998 (N_27998,N_26092,N_26319);
and U27999 (N_27999,N_26016,N_26120);
xor U28000 (N_28000,N_27643,N_27215);
nand U28001 (N_28001,N_27512,N_27622);
xor U28002 (N_28002,N_27167,N_27415);
nor U28003 (N_28003,N_27555,N_27154);
xnor U28004 (N_28004,N_27232,N_27039);
xnor U28005 (N_28005,N_27141,N_27911);
and U28006 (N_28006,N_27488,N_27564);
xor U28007 (N_28007,N_27427,N_27260);
nand U28008 (N_28008,N_27537,N_27716);
and U28009 (N_28009,N_27422,N_27290);
nor U28010 (N_28010,N_27848,N_27379);
or U28011 (N_28011,N_27582,N_27693);
nand U28012 (N_28012,N_27075,N_27481);
nand U28013 (N_28013,N_27866,N_27019);
xnor U28014 (N_28014,N_27103,N_27806);
xnor U28015 (N_28015,N_27910,N_27960);
nand U28016 (N_28016,N_27558,N_27183);
nor U28017 (N_28017,N_27925,N_27596);
nand U28018 (N_28018,N_27822,N_27767);
xnor U28019 (N_28019,N_27938,N_27185);
nand U28020 (N_28020,N_27626,N_27340);
nor U28021 (N_28021,N_27342,N_27414);
nor U28022 (N_28022,N_27800,N_27688);
and U28023 (N_28023,N_27906,N_27684);
and U28024 (N_28024,N_27660,N_27839);
or U28025 (N_28025,N_27847,N_27599);
nor U28026 (N_28026,N_27190,N_27631);
nand U28027 (N_28027,N_27413,N_27197);
or U28028 (N_28028,N_27172,N_27506);
xor U28029 (N_28029,N_27874,N_27179);
nand U28030 (N_28030,N_27694,N_27174);
nand U28031 (N_28031,N_27679,N_27971);
or U28032 (N_28032,N_27177,N_27907);
nor U28033 (N_28033,N_27020,N_27160);
nor U28034 (N_28034,N_27431,N_27901);
and U28035 (N_28035,N_27089,N_27478);
nor U28036 (N_28036,N_27888,N_27718);
and U28037 (N_28037,N_27311,N_27871);
nand U28038 (N_28038,N_27516,N_27509);
nor U28039 (N_28039,N_27662,N_27271);
nand U28040 (N_28040,N_27743,N_27973);
nor U28041 (N_28041,N_27374,N_27578);
or U28042 (N_28042,N_27817,N_27323);
xor U28043 (N_28043,N_27850,N_27354);
nand U28044 (N_28044,N_27956,N_27893);
xor U28045 (N_28045,N_27265,N_27169);
nand U28046 (N_28046,N_27088,N_27915);
nor U28047 (N_28047,N_27671,N_27708);
or U28048 (N_28048,N_27119,N_27037);
or U28049 (N_28049,N_27081,N_27436);
nand U28050 (N_28050,N_27491,N_27018);
xor U28051 (N_28051,N_27859,N_27793);
or U28052 (N_28052,N_27341,N_27730);
nand U28053 (N_28053,N_27394,N_27362);
nor U28054 (N_28054,N_27916,N_27992);
xnor U28055 (N_28055,N_27247,N_27411);
nand U28056 (N_28056,N_27844,N_27476);
xor U28057 (N_28057,N_27490,N_27745);
and U28058 (N_28058,N_27444,N_27281);
and U28059 (N_28059,N_27267,N_27051);
nand U28060 (N_28060,N_27155,N_27189);
nand U28061 (N_28061,N_27496,N_27303);
nor U28062 (N_28062,N_27222,N_27041);
and U28063 (N_28063,N_27331,N_27269);
nor U28064 (N_28064,N_27410,N_27950);
nand U28065 (N_28065,N_27968,N_27614);
or U28066 (N_28066,N_27810,N_27263);
nand U28067 (N_28067,N_27315,N_27601);
nand U28068 (N_28068,N_27854,N_27638);
and U28069 (N_28069,N_27367,N_27941);
or U28070 (N_28070,N_27001,N_27337);
and U28071 (N_28071,N_27248,N_27762);
nor U28072 (N_28072,N_27188,N_27869);
or U28073 (N_28073,N_27515,N_27784);
and U28074 (N_28074,N_27621,N_27291);
nand U28075 (N_28075,N_27139,N_27565);
xnor U28076 (N_28076,N_27369,N_27698);
xnor U28077 (N_28077,N_27495,N_27937);
nand U28078 (N_28078,N_27192,N_27191);
nand U28079 (N_28079,N_27732,N_27405);
xor U28080 (N_28080,N_27213,N_27021);
nor U28081 (N_28081,N_27585,N_27385);
or U28082 (N_28082,N_27485,N_27140);
xor U28083 (N_28083,N_27097,N_27908);
xor U28084 (N_28084,N_27113,N_27744);
and U28085 (N_28085,N_27138,N_27957);
nor U28086 (N_28086,N_27691,N_27640);
xnor U28087 (N_28087,N_27737,N_27975);
nand U28088 (N_28088,N_27771,N_27508);
nor U28089 (N_28089,N_27759,N_27980);
nor U28090 (N_28090,N_27650,N_27796);
xnor U28091 (N_28091,N_27469,N_27005);
or U28092 (N_28092,N_27628,N_27392);
nand U28093 (N_28093,N_27579,N_27867);
nand U28094 (N_28094,N_27896,N_27373);
and U28095 (N_28095,N_27753,N_27317);
or U28096 (N_28096,N_27209,N_27674);
or U28097 (N_28097,N_27296,N_27324);
xnor U28098 (N_28098,N_27282,N_27297);
xor U28099 (N_28099,N_27636,N_27335);
nor U28100 (N_28100,N_27078,N_27522);
or U28101 (N_28101,N_27846,N_27002);
or U28102 (N_28102,N_27059,N_27196);
xor U28103 (N_28103,N_27229,N_27024);
or U28104 (N_28104,N_27498,N_27243);
xor U28105 (N_28105,N_27013,N_27775);
and U28106 (N_28106,N_27251,N_27382);
and U28107 (N_28107,N_27993,N_27548);
xnor U28108 (N_28108,N_27991,N_27393);
xnor U28109 (N_28109,N_27518,N_27715);
or U28110 (N_28110,N_27738,N_27357);
and U28111 (N_28111,N_27349,N_27946);
nand U28112 (N_28112,N_27388,N_27090);
xor U28113 (N_28113,N_27895,N_27409);
nand U28114 (N_28114,N_27722,N_27124);
nor U28115 (N_28115,N_27602,N_27117);
nand U28116 (N_28116,N_27023,N_27010);
nor U28117 (N_28117,N_27658,N_27418);
and U28118 (N_28118,N_27524,N_27554);
nor U28119 (N_28119,N_27381,N_27986);
nor U28120 (N_28120,N_27507,N_27562);
or U28121 (N_28121,N_27539,N_27497);
or U28122 (N_28122,N_27456,N_27985);
nor U28123 (N_28123,N_27742,N_27584);
nor U28124 (N_28124,N_27559,N_27840);
and U28125 (N_28125,N_27761,N_27987);
nand U28126 (N_28126,N_27990,N_27092);
or U28127 (N_28127,N_27923,N_27459);
nor U28128 (N_28128,N_27821,N_27580);
nor U28129 (N_28129,N_27238,N_27082);
nand U28130 (N_28130,N_27783,N_27003);
nand U28131 (N_28131,N_27791,N_27187);
nor U28132 (N_28132,N_27173,N_27466);
or U28133 (N_28133,N_27300,N_27032);
and U28134 (N_28134,N_27913,N_27760);
nor U28135 (N_28135,N_27406,N_27079);
nor U28136 (N_28136,N_27242,N_27890);
nor U28137 (N_28137,N_27057,N_27995);
nand U28138 (N_28138,N_27472,N_27450);
nor U28139 (N_28139,N_27408,N_27989);
nor U28140 (N_28140,N_27186,N_27678);
or U28141 (N_28141,N_27503,N_27811);
nor U28142 (N_28142,N_27273,N_27130);
or U28143 (N_28143,N_27820,N_27223);
and U28144 (N_28144,N_27677,N_27065);
nor U28145 (N_28145,N_27216,N_27587);
and U28146 (N_28146,N_27787,N_27948);
and U28147 (N_28147,N_27504,N_27977);
xor U28148 (N_28148,N_27107,N_27752);
nor U28149 (N_28149,N_27253,N_27400);
nand U28150 (N_28150,N_27045,N_27055);
xnor U28151 (N_28151,N_27484,N_27513);
and U28152 (N_28152,N_27531,N_27511);
xor U28153 (N_28153,N_27148,N_27774);
and U28154 (N_28154,N_27280,N_27012);
xor U28155 (N_28155,N_27729,N_27348);
and U28156 (N_28156,N_27339,N_27115);
and U28157 (N_28157,N_27210,N_27104);
and U28158 (N_28158,N_27552,N_27686);
and U28159 (N_28159,N_27245,N_27390);
nor U28160 (N_28160,N_27309,N_27900);
nor U28161 (N_28161,N_27723,N_27590);
or U28162 (N_28162,N_27573,N_27050);
nor U28163 (N_28163,N_27345,N_27486);
or U28164 (N_28164,N_27212,N_27788);
nand U28165 (N_28165,N_27884,N_27049);
nand U28166 (N_28166,N_27852,N_27963);
xor U28167 (N_28167,N_27417,N_27195);
nand U28168 (N_28168,N_27231,N_27804);
and U28169 (N_28169,N_27270,N_27670);
nand U28170 (N_28170,N_27333,N_27036);
nand U28171 (N_28171,N_27028,N_27689);
and U28172 (N_28172,N_27945,N_27276);
nor U28173 (N_28173,N_27605,N_27816);
nand U28174 (N_28174,N_27813,N_27721);
nor U28175 (N_28175,N_27122,N_27735);
or U28176 (N_28176,N_27812,N_27208);
and U28177 (N_28177,N_27114,N_27446);
xor U28178 (N_28178,N_27668,N_27627);
nand U28179 (N_28179,N_27700,N_27007);
xnor U28180 (N_28180,N_27619,N_27087);
or U28181 (N_28181,N_27842,N_27483);
xnor U28182 (N_28182,N_27157,N_27110);
nor U28183 (N_28183,N_27933,N_27171);
nand U28184 (N_28184,N_27040,N_27862);
nor U28185 (N_28185,N_27940,N_27182);
nand U28186 (N_28186,N_27268,N_27334);
nand U28187 (N_28187,N_27633,N_27125);
and U28188 (N_28188,N_27778,N_27999);
xor U28189 (N_28189,N_27288,N_27560);
nor U28190 (N_28190,N_27831,N_27672);
nand U28191 (N_28191,N_27731,N_27246);
or U28192 (N_28192,N_27758,N_27876);
nand U28193 (N_28193,N_27184,N_27814);
and U28194 (N_28194,N_27434,N_27329);
or U28195 (N_28195,N_27170,N_27285);
xor U28196 (N_28196,N_27266,N_27914);
nand U28197 (N_28197,N_27561,N_27378);
xnor U28198 (N_28198,N_27261,N_27889);
xor U28199 (N_28199,N_27287,N_27519);
nand U28200 (N_28200,N_27361,N_27624);
xnor U28201 (N_28201,N_27494,N_27949);
nor U28202 (N_28202,N_27194,N_27607);
xnor U28203 (N_28203,N_27733,N_27589);
or U28204 (N_28204,N_27604,N_27623);
nor U28205 (N_28205,N_27147,N_27967);
or U28206 (N_28206,N_27663,N_27625);
and U28207 (N_28207,N_27074,N_27353);
or U28208 (N_28208,N_27085,N_27551);
and U28209 (N_28209,N_27838,N_27048);
nor U28210 (N_28210,N_27439,N_27064);
or U28211 (N_28211,N_27568,N_27894);
nor U28212 (N_28212,N_27666,N_27827);
xnor U28213 (N_28213,N_27371,N_27538);
and U28214 (N_28214,N_27756,N_27609);
or U28215 (N_28215,N_27868,N_27637);
nor U28216 (N_28216,N_27520,N_27563);
nor U28217 (N_28217,N_27424,N_27720);
nand U28218 (N_28218,N_27416,N_27805);
nand U28219 (N_28219,N_27274,N_27219);
xor U28220 (N_28220,N_27873,N_27134);
or U28221 (N_28221,N_27314,N_27221);
and U28222 (N_28222,N_27951,N_27440);
and U28223 (N_28223,N_27086,N_27642);
and U28224 (N_28224,N_27084,N_27308);
xnor U28225 (N_28225,N_27815,N_27566);
nand U28226 (N_28226,N_27206,N_27632);
and U28227 (N_28227,N_27754,N_27403);
or U28228 (N_28228,N_27818,N_27043);
nand U28229 (N_28229,N_27437,N_27033);
nor U28230 (N_28230,N_27717,N_27819);
xor U28231 (N_28231,N_27256,N_27930);
xor U28232 (N_28232,N_27830,N_27961);
nand U28233 (N_28233,N_27461,N_27380);
xnor U28234 (N_28234,N_27465,N_27404);
nor U28235 (N_28235,N_27644,N_27105);
and U28236 (N_28236,N_27149,N_27284);
nand U28237 (N_28237,N_27741,N_27098);
nand U28238 (N_28238,N_27430,N_27858);
xor U28239 (N_28239,N_27740,N_27006);
or U28240 (N_28240,N_27029,N_27581);
xnor U28241 (N_28241,N_27947,N_27710);
nand U28242 (N_28242,N_27824,N_27054);
or U28243 (N_28243,N_27060,N_27545);
xnor U28244 (N_28244,N_27667,N_27225);
and U28245 (N_28245,N_27880,N_27591);
and U28246 (N_28246,N_27843,N_27499);
nand U28247 (N_28247,N_27473,N_27258);
or U28248 (N_28248,N_27978,N_27398);
xnor U28249 (N_28249,N_27794,N_27988);
and U28250 (N_28250,N_27161,N_27226);
xor U28251 (N_28251,N_27919,N_27726);
or U28252 (N_28252,N_27257,N_27533);
nand U28253 (N_28253,N_27798,N_27709);
xnor U28254 (N_28254,N_27047,N_27457);
or U28255 (N_28255,N_27143,N_27096);
xor U28256 (N_28256,N_27254,N_27034);
xor U28257 (N_28257,N_27181,N_27200);
and U28258 (N_28258,N_27872,N_27176);
xor U28259 (N_28259,N_27252,N_27351);
xor U28260 (N_28260,N_27121,N_27505);
and U28261 (N_28261,N_27825,N_27077);
or U28262 (N_28262,N_27364,N_27395);
nand U28263 (N_28263,N_27714,N_27707);
xor U28264 (N_28264,N_27111,N_27305);
and U28265 (N_28265,N_27904,N_27801);
or U28266 (N_28266,N_27629,N_27675);
nor U28267 (N_28267,N_27336,N_27454);
nand U28268 (N_28268,N_27468,N_27014);
xnor U28269 (N_28269,N_27926,N_27412);
nor U28270 (N_28270,N_27249,N_27031);
or U28271 (N_28271,N_27312,N_27489);
nand U28272 (N_28272,N_27201,N_27493);
xnor U28273 (N_28273,N_27523,N_27135);
xnor U28274 (N_28274,N_27396,N_27487);
xor U28275 (N_28275,N_27535,N_27687);
xnor U28276 (N_28276,N_27885,N_27569);
nor U28277 (N_28277,N_27779,N_27883);
or U28278 (N_28278,N_27510,N_27166);
xnor U28279 (N_28279,N_27441,N_27851);
nand U28280 (N_28280,N_27199,N_27841);
or U28281 (N_28281,N_27118,N_27865);
nand U28282 (N_28282,N_27294,N_27870);
xor U28283 (N_28283,N_27630,N_27724);
or U28284 (N_28284,N_27272,N_27165);
or U28285 (N_28285,N_27091,N_27070);
xnor U28286 (N_28286,N_27375,N_27072);
and U28287 (N_28287,N_27429,N_27463);
and U28288 (N_28288,N_27931,N_27255);
nor U28289 (N_28289,N_27344,N_27703);
nor U28290 (N_28290,N_27328,N_27244);
and U28291 (N_28291,N_27583,N_27586);
and U28292 (N_28292,N_27681,N_27377);
or U28293 (N_28293,N_27570,N_27879);
xor U28294 (N_28294,N_27015,N_27860);
nand U28295 (N_28295,N_27777,N_27616);
nor U28296 (N_28296,N_27202,N_27474);
xor U28297 (N_28297,N_27891,N_27056);
nor U28298 (N_28298,N_27809,N_27776);
nor U28299 (N_28299,N_27802,N_27592);
nand U28300 (N_28300,N_27479,N_27435);
nor U28301 (N_28301,N_27112,N_27000);
nor U28302 (N_28302,N_27211,N_27952);
and U28303 (N_28303,N_27711,N_27534);
nor U28304 (N_28304,N_27932,N_27797);
xnor U28305 (N_28305,N_27180,N_27445);
xnor U28306 (N_28306,N_27557,N_27144);
and U28307 (N_28307,N_27407,N_27358);
and U28308 (N_28308,N_27017,N_27123);
nor U28309 (N_28309,N_27598,N_27239);
or U28310 (N_28310,N_27690,N_27327);
or U28311 (N_28311,N_27250,N_27136);
or U28312 (N_28312,N_27608,N_27347);
or U28313 (N_28313,N_27620,N_27939);
nor U28314 (N_28314,N_27163,N_27647);
xnor U28315 (N_28315,N_27443,N_27073);
xnor U28316 (N_28316,N_27882,N_27203);
nor U28317 (N_28317,N_27067,N_27321);
nand U28318 (N_28318,N_27706,N_27764);
or U28319 (N_28319,N_27521,N_27542);
nand U28320 (N_28320,N_27976,N_27655);
nand U28321 (N_28321,N_27235,N_27918);
and U28322 (N_28322,N_27669,N_27318);
nand U28323 (N_28323,N_27420,N_27464);
and U28324 (N_28324,N_27799,N_27363);
or U28325 (N_28325,N_27228,N_27026);
and U28326 (N_28326,N_27343,N_27419);
nor U28327 (N_28327,N_27008,N_27790);
and U28328 (N_28328,N_27823,N_27536);
and U28329 (N_28329,N_27304,N_27127);
and U28330 (N_28330,N_27836,N_27207);
xor U28331 (N_28331,N_27289,N_27530);
xnor U28332 (N_28332,N_27834,N_27702);
and U28333 (N_28333,N_27350,N_27151);
or U28334 (N_28334,N_27603,N_27102);
and U28335 (N_28335,N_27205,N_27142);
nand U28336 (N_28336,N_27984,N_27829);
or U28337 (N_28337,N_27052,N_27974);
xnor U28338 (N_28338,N_27982,N_27046);
and U28339 (N_28339,N_27025,N_27164);
nand U28340 (N_28340,N_27983,N_27673);
nand U28341 (N_28341,N_27279,N_27359);
or U28342 (N_28342,N_27168,N_27158);
nand U28343 (N_28343,N_27612,N_27338);
nand U28344 (N_28344,N_27728,N_27757);
nor U28345 (N_28345,N_27071,N_27746);
xnor U28346 (N_28346,N_27397,N_27692);
nor U28347 (N_28347,N_27944,N_27540);
or U28348 (N_28348,N_27654,N_27386);
xnor U28349 (N_28349,N_27099,N_27917);
nor U28350 (N_28350,N_27966,N_27264);
or U28351 (N_28351,N_27763,N_27998);
nor U28352 (N_28352,N_27769,N_27480);
and U28353 (N_28353,N_27886,N_27795);
xnor U28354 (N_28354,N_27068,N_27204);
xor U28355 (N_28355,N_27645,N_27855);
nor U28356 (N_28356,N_27832,N_27193);
or U28357 (N_28357,N_27042,N_27828);
and U28358 (N_28358,N_27748,N_27278);
or U28359 (N_28359,N_27845,N_27175);
nor U28360 (N_28360,N_27458,N_27150);
nor U28361 (N_28361,N_27922,N_27368);
xor U28362 (N_28362,N_27061,N_27792);
and U28363 (N_28363,N_27835,N_27109);
or U28364 (N_28364,N_27330,N_27384);
and U28365 (N_28365,N_27705,N_27100);
and U28366 (N_28366,N_27234,N_27864);
and U28367 (N_28367,N_27313,N_27546);
and U28368 (N_28368,N_27528,N_27525);
nand U28369 (N_28369,N_27970,N_27389);
and U28370 (N_28370,N_27549,N_27979);
xnor U28371 (N_28371,N_27929,N_27106);
xnor U28372 (N_28372,N_27310,N_27962);
nand U28373 (N_28373,N_27943,N_27217);
or U28374 (N_28374,N_27902,N_27502);
nand U28375 (N_28375,N_27685,N_27853);
xnor U28376 (N_28376,N_27030,N_27126);
nor U28377 (N_28377,N_27652,N_27571);
and U28378 (N_28378,N_27892,N_27402);
and U28379 (N_28379,N_27004,N_27550);
xor U28380 (N_28380,N_27713,N_27076);
xor U28381 (N_28381,N_27969,N_27661);
nand U28382 (N_28382,N_27897,N_27936);
or U28383 (N_28383,N_27083,N_27162);
nand U28384 (N_28384,N_27768,N_27606);
or U28385 (N_28385,N_27553,N_27611);
xor U28386 (N_28386,N_27286,N_27452);
and U28387 (N_28387,N_27651,N_27133);
or U28388 (N_28388,N_27449,N_27292);
or U28389 (N_28389,N_27575,N_27712);
nor U28390 (N_28390,N_27682,N_27218);
and U28391 (N_28391,N_27996,N_27588);
nor U28392 (N_28392,N_27198,N_27942);
nor U28393 (N_28393,N_27275,N_27066);
and U28394 (N_28394,N_27322,N_27556);
or U28395 (N_28395,N_27293,N_27877);
or U28396 (N_28396,N_27927,N_27346);
nor U28397 (N_28397,N_27016,N_27898);
or U28398 (N_28398,N_27826,N_27069);
nor U28399 (N_28399,N_27924,N_27965);
nor U28400 (N_28400,N_27649,N_27120);
xor U28401 (N_28401,N_27696,N_27541);
and U28402 (N_28402,N_27352,N_27356);
or U28403 (N_28403,N_27697,N_27594);
or U28404 (N_28404,N_27425,N_27749);
and U28405 (N_28405,N_27383,N_27921);
or U28406 (N_28406,N_27856,N_27467);
nand U28407 (N_28407,N_27224,N_27448);
or U28408 (N_28408,N_27803,N_27526);
or U28409 (N_28409,N_27220,N_27500);
and U28410 (N_28410,N_27447,N_27302);
and U28411 (N_28411,N_27230,N_27887);
xnor U28412 (N_28412,N_27233,N_27751);
nand U28413 (N_28413,N_27909,N_27849);
nor U28414 (N_28414,N_27475,N_27320);
xor U28415 (N_28415,N_27146,N_27426);
nand U28416 (N_28416,N_27755,N_27736);
nor U28417 (N_28417,N_27460,N_27517);
xor U28418 (N_28418,N_27132,N_27316);
xor U28419 (N_28419,N_27899,N_27656);
xor U28420 (N_28420,N_27837,N_27453);
xnor U28421 (N_28421,N_27372,N_27782);
xnor U28422 (N_28422,N_27298,N_27326);
or U28423 (N_28423,N_27063,N_27237);
xor U28424 (N_28424,N_27227,N_27370);
nand U28425 (N_28425,N_27492,N_27038);
and U28426 (N_28426,N_27438,N_27325);
xor U28427 (N_28427,N_27959,N_27617);
nand U28428 (N_28428,N_27332,N_27833);
nor U28429 (N_28429,N_27955,N_27905);
or U28430 (N_28430,N_27241,N_27391);
nand U28431 (N_28431,N_27131,N_27366);
nor U28432 (N_28432,N_27972,N_27739);
or U28433 (N_28433,N_27595,N_27773);
nand U28434 (N_28434,N_27306,N_27572);
and U28435 (N_28435,N_27470,N_27683);
nor U28436 (N_28436,N_27301,N_27547);
xor U28437 (N_28437,N_27451,N_27145);
xor U28438 (N_28438,N_27455,N_27719);
or U28439 (N_28439,N_27615,N_27080);
or U28440 (N_28440,N_27781,N_27665);
or U28441 (N_28441,N_27657,N_27259);
xnor U28442 (N_28442,N_27994,N_27981);
xnor U28443 (N_28443,N_27577,N_27646);
and U28444 (N_28444,N_27432,N_27861);
nand U28445 (N_28445,N_27421,N_27808);
nand U28446 (N_28446,N_27863,N_27664);
and U28447 (N_28447,N_27178,N_27307);
nand U28448 (N_28448,N_27035,N_27574);
nor U28449 (N_28449,N_27128,N_27704);
or U28450 (N_28450,N_27482,N_27727);
xor U28451 (N_28451,N_27094,N_27928);
nand U28452 (N_28452,N_27011,N_27428);
nand U28453 (N_28453,N_27648,N_27399);
and U28454 (N_28454,N_27964,N_27527);
and U28455 (N_28455,N_27116,N_27734);
nand U28456 (N_28456,N_27789,N_27462);
nand U28457 (N_28457,N_27857,N_27600);
nand U28458 (N_28458,N_27283,N_27997);
nand U28459 (N_28459,N_27567,N_27137);
and U28460 (N_28460,N_27360,N_27695);
xnor U28461 (N_28461,N_27770,N_27634);
or U28462 (N_28462,N_27214,N_27954);
xor U28463 (N_28463,N_27699,N_27780);
xnor U28464 (N_28464,N_27613,N_27639);
and U28465 (N_28465,N_27920,N_27772);
xnor U28466 (N_28466,N_27058,N_27543);
xnor U28467 (N_28467,N_27477,N_27442);
nand U28468 (N_28468,N_27355,N_27610);
nand U28469 (N_28469,N_27532,N_27875);
xnor U28470 (N_28470,N_27701,N_27953);
nor U28471 (N_28471,N_27299,N_27401);
or U28472 (N_28472,N_27062,N_27912);
and U28473 (N_28473,N_27881,N_27022);
nor U28474 (N_28474,N_27544,N_27152);
and U28475 (N_28475,N_27501,N_27765);
or U28476 (N_28476,N_27053,N_27725);
or U28477 (N_28477,N_27277,N_27514);
and U28478 (N_28478,N_27576,N_27095);
xnor U28479 (N_28479,N_27676,N_27156);
nand U28480 (N_28480,N_27618,N_27433);
nor U28481 (N_28481,N_27786,N_27159);
or U28482 (N_28482,N_27807,N_27747);
nand U28483 (N_28483,N_27766,N_27240);
or U28484 (N_28484,N_27659,N_27423);
or U28485 (N_28485,N_27044,N_27934);
nor U28486 (N_28486,N_27365,N_27236);
xnor U28487 (N_28487,N_27376,N_27295);
nor U28488 (N_28488,N_27878,N_27597);
nor U28489 (N_28489,N_27027,N_27785);
or U28490 (N_28490,N_27108,N_27129);
and U28491 (N_28491,N_27680,N_27635);
and U28492 (N_28492,N_27471,N_27935);
and U28493 (N_28493,N_27529,N_27093);
and U28494 (N_28494,N_27653,N_27262);
or U28495 (N_28495,N_27750,N_27903);
or U28496 (N_28496,N_27153,N_27009);
nand U28497 (N_28497,N_27101,N_27593);
nand U28498 (N_28498,N_27387,N_27641);
or U28499 (N_28499,N_27958,N_27319);
nor U28500 (N_28500,N_27568,N_27089);
xor U28501 (N_28501,N_27523,N_27871);
xor U28502 (N_28502,N_27206,N_27776);
nand U28503 (N_28503,N_27169,N_27419);
nand U28504 (N_28504,N_27516,N_27531);
or U28505 (N_28505,N_27810,N_27350);
xnor U28506 (N_28506,N_27092,N_27846);
and U28507 (N_28507,N_27783,N_27518);
nand U28508 (N_28508,N_27671,N_27467);
and U28509 (N_28509,N_27039,N_27951);
nor U28510 (N_28510,N_27546,N_27164);
nor U28511 (N_28511,N_27651,N_27927);
xnor U28512 (N_28512,N_27425,N_27395);
and U28513 (N_28513,N_27461,N_27252);
and U28514 (N_28514,N_27388,N_27710);
or U28515 (N_28515,N_27369,N_27417);
nor U28516 (N_28516,N_27405,N_27613);
xnor U28517 (N_28517,N_27464,N_27086);
nor U28518 (N_28518,N_27034,N_27905);
nor U28519 (N_28519,N_27308,N_27784);
nor U28520 (N_28520,N_27428,N_27797);
xnor U28521 (N_28521,N_27358,N_27929);
or U28522 (N_28522,N_27898,N_27941);
and U28523 (N_28523,N_27655,N_27564);
and U28524 (N_28524,N_27403,N_27098);
or U28525 (N_28525,N_27462,N_27619);
nand U28526 (N_28526,N_27564,N_27520);
or U28527 (N_28527,N_27582,N_27392);
nor U28528 (N_28528,N_27840,N_27001);
or U28529 (N_28529,N_27573,N_27574);
nand U28530 (N_28530,N_27032,N_27008);
nor U28531 (N_28531,N_27202,N_27400);
and U28532 (N_28532,N_27124,N_27906);
or U28533 (N_28533,N_27208,N_27253);
nor U28534 (N_28534,N_27015,N_27638);
or U28535 (N_28535,N_27528,N_27899);
nor U28536 (N_28536,N_27976,N_27792);
or U28537 (N_28537,N_27407,N_27018);
and U28538 (N_28538,N_27632,N_27545);
and U28539 (N_28539,N_27985,N_27113);
xor U28540 (N_28540,N_27225,N_27650);
or U28541 (N_28541,N_27759,N_27734);
nor U28542 (N_28542,N_27446,N_27175);
or U28543 (N_28543,N_27861,N_27668);
and U28544 (N_28544,N_27290,N_27711);
xor U28545 (N_28545,N_27928,N_27098);
nand U28546 (N_28546,N_27687,N_27753);
and U28547 (N_28547,N_27011,N_27137);
nand U28548 (N_28548,N_27566,N_27874);
and U28549 (N_28549,N_27584,N_27297);
nand U28550 (N_28550,N_27450,N_27886);
nor U28551 (N_28551,N_27198,N_27468);
and U28552 (N_28552,N_27512,N_27410);
nor U28553 (N_28553,N_27784,N_27856);
and U28554 (N_28554,N_27480,N_27661);
or U28555 (N_28555,N_27143,N_27208);
or U28556 (N_28556,N_27020,N_27567);
xor U28557 (N_28557,N_27253,N_27120);
nor U28558 (N_28558,N_27296,N_27003);
nand U28559 (N_28559,N_27077,N_27266);
or U28560 (N_28560,N_27698,N_27610);
nor U28561 (N_28561,N_27434,N_27390);
or U28562 (N_28562,N_27490,N_27549);
xnor U28563 (N_28563,N_27760,N_27258);
nand U28564 (N_28564,N_27270,N_27696);
xnor U28565 (N_28565,N_27501,N_27154);
or U28566 (N_28566,N_27295,N_27474);
nand U28567 (N_28567,N_27736,N_27090);
and U28568 (N_28568,N_27820,N_27897);
xnor U28569 (N_28569,N_27406,N_27080);
nand U28570 (N_28570,N_27240,N_27499);
or U28571 (N_28571,N_27099,N_27356);
nand U28572 (N_28572,N_27522,N_27926);
or U28573 (N_28573,N_27555,N_27971);
xor U28574 (N_28574,N_27794,N_27224);
and U28575 (N_28575,N_27651,N_27066);
xor U28576 (N_28576,N_27552,N_27927);
nor U28577 (N_28577,N_27149,N_27066);
nand U28578 (N_28578,N_27112,N_27751);
nor U28579 (N_28579,N_27570,N_27166);
nor U28580 (N_28580,N_27852,N_27359);
or U28581 (N_28581,N_27753,N_27995);
nor U28582 (N_28582,N_27524,N_27113);
nor U28583 (N_28583,N_27192,N_27147);
or U28584 (N_28584,N_27825,N_27421);
xnor U28585 (N_28585,N_27701,N_27708);
nor U28586 (N_28586,N_27649,N_27680);
nand U28587 (N_28587,N_27605,N_27455);
nand U28588 (N_28588,N_27032,N_27368);
nand U28589 (N_28589,N_27618,N_27813);
and U28590 (N_28590,N_27809,N_27982);
and U28591 (N_28591,N_27028,N_27696);
nor U28592 (N_28592,N_27400,N_27298);
or U28593 (N_28593,N_27831,N_27362);
xor U28594 (N_28594,N_27619,N_27333);
nor U28595 (N_28595,N_27793,N_27885);
and U28596 (N_28596,N_27388,N_27438);
and U28597 (N_28597,N_27924,N_27181);
and U28598 (N_28598,N_27333,N_27859);
and U28599 (N_28599,N_27866,N_27951);
and U28600 (N_28600,N_27085,N_27305);
and U28601 (N_28601,N_27680,N_27235);
and U28602 (N_28602,N_27447,N_27931);
or U28603 (N_28603,N_27335,N_27621);
nand U28604 (N_28604,N_27696,N_27427);
nand U28605 (N_28605,N_27285,N_27741);
or U28606 (N_28606,N_27866,N_27229);
nor U28607 (N_28607,N_27635,N_27135);
xnor U28608 (N_28608,N_27175,N_27289);
nand U28609 (N_28609,N_27677,N_27861);
nand U28610 (N_28610,N_27304,N_27323);
xor U28611 (N_28611,N_27270,N_27258);
nand U28612 (N_28612,N_27268,N_27633);
and U28613 (N_28613,N_27078,N_27705);
or U28614 (N_28614,N_27079,N_27271);
xor U28615 (N_28615,N_27264,N_27462);
or U28616 (N_28616,N_27666,N_27710);
nor U28617 (N_28617,N_27847,N_27772);
or U28618 (N_28618,N_27388,N_27960);
or U28619 (N_28619,N_27869,N_27640);
and U28620 (N_28620,N_27177,N_27608);
nand U28621 (N_28621,N_27614,N_27249);
nand U28622 (N_28622,N_27326,N_27880);
or U28623 (N_28623,N_27114,N_27048);
or U28624 (N_28624,N_27541,N_27025);
and U28625 (N_28625,N_27901,N_27132);
and U28626 (N_28626,N_27575,N_27755);
and U28627 (N_28627,N_27759,N_27901);
nor U28628 (N_28628,N_27375,N_27674);
or U28629 (N_28629,N_27922,N_27612);
nand U28630 (N_28630,N_27870,N_27721);
or U28631 (N_28631,N_27620,N_27543);
and U28632 (N_28632,N_27953,N_27621);
xnor U28633 (N_28633,N_27493,N_27390);
nand U28634 (N_28634,N_27860,N_27947);
or U28635 (N_28635,N_27562,N_27497);
nor U28636 (N_28636,N_27822,N_27381);
nand U28637 (N_28637,N_27600,N_27261);
or U28638 (N_28638,N_27296,N_27861);
nand U28639 (N_28639,N_27944,N_27698);
or U28640 (N_28640,N_27901,N_27299);
nand U28641 (N_28641,N_27536,N_27100);
nor U28642 (N_28642,N_27690,N_27442);
and U28643 (N_28643,N_27952,N_27558);
or U28644 (N_28644,N_27320,N_27705);
nand U28645 (N_28645,N_27550,N_27557);
nor U28646 (N_28646,N_27925,N_27300);
nand U28647 (N_28647,N_27301,N_27764);
xor U28648 (N_28648,N_27870,N_27729);
nor U28649 (N_28649,N_27014,N_27493);
nor U28650 (N_28650,N_27212,N_27123);
xor U28651 (N_28651,N_27653,N_27781);
nor U28652 (N_28652,N_27064,N_27028);
nand U28653 (N_28653,N_27986,N_27671);
nand U28654 (N_28654,N_27040,N_27402);
xnor U28655 (N_28655,N_27655,N_27774);
nand U28656 (N_28656,N_27306,N_27486);
nand U28657 (N_28657,N_27152,N_27777);
nor U28658 (N_28658,N_27166,N_27805);
nor U28659 (N_28659,N_27254,N_27836);
nand U28660 (N_28660,N_27830,N_27693);
nor U28661 (N_28661,N_27132,N_27450);
xor U28662 (N_28662,N_27728,N_27672);
and U28663 (N_28663,N_27197,N_27142);
xnor U28664 (N_28664,N_27201,N_27306);
and U28665 (N_28665,N_27626,N_27046);
or U28666 (N_28666,N_27564,N_27835);
xnor U28667 (N_28667,N_27663,N_27746);
and U28668 (N_28668,N_27166,N_27780);
and U28669 (N_28669,N_27214,N_27835);
xor U28670 (N_28670,N_27598,N_27276);
nand U28671 (N_28671,N_27369,N_27535);
nor U28672 (N_28672,N_27938,N_27560);
and U28673 (N_28673,N_27810,N_27257);
nand U28674 (N_28674,N_27972,N_27159);
xnor U28675 (N_28675,N_27400,N_27346);
or U28676 (N_28676,N_27713,N_27820);
nor U28677 (N_28677,N_27206,N_27787);
or U28678 (N_28678,N_27564,N_27436);
and U28679 (N_28679,N_27106,N_27902);
xnor U28680 (N_28680,N_27497,N_27424);
and U28681 (N_28681,N_27358,N_27714);
nand U28682 (N_28682,N_27866,N_27631);
and U28683 (N_28683,N_27503,N_27038);
xnor U28684 (N_28684,N_27481,N_27299);
and U28685 (N_28685,N_27514,N_27211);
nand U28686 (N_28686,N_27565,N_27760);
xor U28687 (N_28687,N_27370,N_27778);
xnor U28688 (N_28688,N_27364,N_27840);
or U28689 (N_28689,N_27720,N_27632);
nor U28690 (N_28690,N_27149,N_27495);
and U28691 (N_28691,N_27032,N_27351);
nor U28692 (N_28692,N_27048,N_27088);
xor U28693 (N_28693,N_27638,N_27349);
and U28694 (N_28694,N_27312,N_27170);
and U28695 (N_28695,N_27147,N_27166);
nand U28696 (N_28696,N_27435,N_27990);
xnor U28697 (N_28697,N_27839,N_27738);
and U28698 (N_28698,N_27519,N_27192);
and U28699 (N_28699,N_27960,N_27373);
or U28700 (N_28700,N_27344,N_27594);
xnor U28701 (N_28701,N_27617,N_27802);
and U28702 (N_28702,N_27764,N_27782);
xor U28703 (N_28703,N_27755,N_27277);
and U28704 (N_28704,N_27828,N_27814);
or U28705 (N_28705,N_27751,N_27975);
nand U28706 (N_28706,N_27633,N_27689);
and U28707 (N_28707,N_27672,N_27267);
xnor U28708 (N_28708,N_27233,N_27675);
xnor U28709 (N_28709,N_27315,N_27502);
and U28710 (N_28710,N_27837,N_27239);
nand U28711 (N_28711,N_27041,N_27254);
nor U28712 (N_28712,N_27301,N_27593);
or U28713 (N_28713,N_27446,N_27632);
xnor U28714 (N_28714,N_27116,N_27063);
and U28715 (N_28715,N_27372,N_27998);
xnor U28716 (N_28716,N_27362,N_27971);
or U28717 (N_28717,N_27379,N_27252);
and U28718 (N_28718,N_27615,N_27431);
and U28719 (N_28719,N_27870,N_27467);
nor U28720 (N_28720,N_27578,N_27287);
xor U28721 (N_28721,N_27135,N_27997);
xnor U28722 (N_28722,N_27761,N_27248);
nor U28723 (N_28723,N_27805,N_27128);
nand U28724 (N_28724,N_27499,N_27874);
nor U28725 (N_28725,N_27172,N_27456);
and U28726 (N_28726,N_27196,N_27109);
xor U28727 (N_28727,N_27342,N_27801);
and U28728 (N_28728,N_27236,N_27380);
nand U28729 (N_28729,N_27423,N_27506);
nor U28730 (N_28730,N_27426,N_27065);
xor U28731 (N_28731,N_27373,N_27995);
xor U28732 (N_28732,N_27051,N_27397);
or U28733 (N_28733,N_27950,N_27285);
nor U28734 (N_28734,N_27786,N_27979);
or U28735 (N_28735,N_27597,N_27973);
nand U28736 (N_28736,N_27900,N_27822);
nand U28737 (N_28737,N_27923,N_27740);
nand U28738 (N_28738,N_27800,N_27973);
xor U28739 (N_28739,N_27185,N_27562);
nor U28740 (N_28740,N_27546,N_27925);
xnor U28741 (N_28741,N_27415,N_27904);
nand U28742 (N_28742,N_27242,N_27616);
nor U28743 (N_28743,N_27943,N_27513);
and U28744 (N_28744,N_27898,N_27481);
nor U28745 (N_28745,N_27826,N_27485);
or U28746 (N_28746,N_27944,N_27358);
nor U28747 (N_28747,N_27654,N_27445);
nor U28748 (N_28748,N_27206,N_27517);
nor U28749 (N_28749,N_27160,N_27819);
nand U28750 (N_28750,N_27208,N_27433);
and U28751 (N_28751,N_27778,N_27024);
or U28752 (N_28752,N_27042,N_27636);
nand U28753 (N_28753,N_27910,N_27441);
xor U28754 (N_28754,N_27377,N_27645);
and U28755 (N_28755,N_27971,N_27031);
or U28756 (N_28756,N_27937,N_27046);
or U28757 (N_28757,N_27950,N_27997);
xnor U28758 (N_28758,N_27899,N_27526);
and U28759 (N_28759,N_27950,N_27488);
nor U28760 (N_28760,N_27649,N_27117);
nor U28761 (N_28761,N_27455,N_27202);
xor U28762 (N_28762,N_27041,N_27384);
and U28763 (N_28763,N_27015,N_27071);
or U28764 (N_28764,N_27981,N_27597);
and U28765 (N_28765,N_27628,N_27943);
nor U28766 (N_28766,N_27178,N_27328);
nand U28767 (N_28767,N_27644,N_27692);
nand U28768 (N_28768,N_27634,N_27670);
nand U28769 (N_28769,N_27722,N_27821);
xor U28770 (N_28770,N_27101,N_27538);
nand U28771 (N_28771,N_27050,N_27520);
xnor U28772 (N_28772,N_27663,N_27510);
and U28773 (N_28773,N_27799,N_27581);
and U28774 (N_28774,N_27073,N_27980);
xnor U28775 (N_28775,N_27180,N_27496);
nor U28776 (N_28776,N_27985,N_27651);
and U28777 (N_28777,N_27200,N_27109);
nor U28778 (N_28778,N_27683,N_27001);
nand U28779 (N_28779,N_27739,N_27153);
nor U28780 (N_28780,N_27541,N_27698);
xnor U28781 (N_28781,N_27037,N_27445);
or U28782 (N_28782,N_27476,N_27632);
nand U28783 (N_28783,N_27074,N_27994);
or U28784 (N_28784,N_27969,N_27049);
xor U28785 (N_28785,N_27073,N_27261);
or U28786 (N_28786,N_27060,N_27047);
or U28787 (N_28787,N_27310,N_27461);
or U28788 (N_28788,N_27454,N_27561);
nor U28789 (N_28789,N_27810,N_27655);
and U28790 (N_28790,N_27455,N_27035);
xor U28791 (N_28791,N_27541,N_27234);
nor U28792 (N_28792,N_27758,N_27355);
nor U28793 (N_28793,N_27785,N_27381);
and U28794 (N_28794,N_27887,N_27706);
nor U28795 (N_28795,N_27797,N_27641);
or U28796 (N_28796,N_27781,N_27909);
and U28797 (N_28797,N_27960,N_27503);
nor U28798 (N_28798,N_27854,N_27485);
and U28799 (N_28799,N_27646,N_27379);
xnor U28800 (N_28800,N_27300,N_27840);
nor U28801 (N_28801,N_27407,N_27606);
nand U28802 (N_28802,N_27050,N_27826);
xnor U28803 (N_28803,N_27889,N_27614);
xor U28804 (N_28804,N_27197,N_27071);
nor U28805 (N_28805,N_27953,N_27033);
or U28806 (N_28806,N_27058,N_27048);
xor U28807 (N_28807,N_27623,N_27009);
nand U28808 (N_28808,N_27590,N_27802);
or U28809 (N_28809,N_27520,N_27744);
and U28810 (N_28810,N_27168,N_27945);
nand U28811 (N_28811,N_27068,N_27541);
xor U28812 (N_28812,N_27524,N_27254);
and U28813 (N_28813,N_27972,N_27195);
nor U28814 (N_28814,N_27428,N_27201);
xor U28815 (N_28815,N_27724,N_27762);
nand U28816 (N_28816,N_27416,N_27457);
nor U28817 (N_28817,N_27723,N_27234);
or U28818 (N_28818,N_27740,N_27677);
or U28819 (N_28819,N_27211,N_27471);
xnor U28820 (N_28820,N_27664,N_27058);
and U28821 (N_28821,N_27163,N_27439);
nand U28822 (N_28822,N_27770,N_27152);
and U28823 (N_28823,N_27024,N_27655);
nor U28824 (N_28824,N_27791,N_27565);
nor U28825 (N_28825,N_27230,N_27851);
nand U28826 (N_28826,N_27419,N_27159);
xnor U28827 (N_28827,N_27987,N_27851);
and U28828 (N_28828,N_27855,N_27981);
or U28829 (N_28829,N_27444,N_27572);
or U28830 (N_28830,N_27637,N_27790);
nand U28831 (N_28831,N_27404,N_27284);
nor U28832 (N_28832,N_27438,N_27663);
and U28833 (N_28833,N_27271,N_27798);
and U28834 (N_28834,N_27505,N_27709);
nand U28835 (N_28835,N_27968,N_27829);
and U28836 (N_28836,N_27985,N_27457);
nand U28837 (N_28837,N_27375,N_27266);
nor U28838 (N_28838,N_27330,N_27197);
nand U28839 (N_28839,N_27157,N_27160);
nor U28840 (N_28840,N_27877,N_27577);
or U28841 (N_28841,N_27603,N_27924);
nor U28842 (N_28842,N_27210,N_27751);
nand U28843 (N_28843,N_27190,N_27095);
and U28844 (N_28844,N_27545,N_27562);
nand U28845 (N_28845,N_27369,N_27738);
and U28846 (N_28846,N_27138,N_27400);
and U28847 (N_28847,N_27436,N_27423);
or U28848 (N_28848,N_27195,N_27492);
nand U28849 (N_28849,N_27959,N_27023);
or U28850 (N_28850,N_27495,N_27227);
nor U28851 (N_28851,N_27723,N_27258);
or U28852 (N_28852,N_27790,N_27420);
xnor U28853 (N_28853,N_27337,N_27223);
and U28854 (N_28854,N_27421,N_27921);
and U28855 (N_28855,N_27420,N_27810);
xor U28856 (N_28856,N_27836,N_27963);
and U28857 (N_28857,N_27515,N_27319);
nor U28858 (N_28858,N_27102,N_27132);
and U28859 (N_28859,N_27273,N_27025);
xor U28860 (N_28860,N_27031,N_27982);
or U28861 (N_28861,N_27660,N_27673);
xor U28862 (N_28862,N_27713,N_27743);
nor U28863 (N_28863,N_27354,N_27445);
nand U28864 (N_28864,N_27519,N_27071);
nand U28865 (N_28865,N_27572,N_27813);
nor U28866 (N_28866,N_27016,N_27963);
nand U28867 (N_28867,N_27133,N_27178);
xnor U28868 (N_28868,N_27435,N_27392);
xor U28869 (N_28869,N_27204,N_27711);
or U28870 (N_28870,N_27793,N_27726);
xor U28871 (N_28871,N_27193,N_27557);
nor U28872 (N_28872,N_27872,N_27643);
nand U28873 (N_28873,N_27443,N_27205);
or U28874 (N_28874,N_27610,N_27514);
nand U28875 (N_28875,N_27799,N_27838);
or U28876 (N_28876,N_27948,N_27375);
nor U28877 (N_28877,N_27985,N_27100);
or U28878 (N_28878,N_27995,N_27930);
nand U28879 (N_28879,N_27007,N_27226);
xor U28880 (N_28880,N_27600,N_27765);
and U28881 (N_28881,N_27525,N_27886);
nand U28882 (N_28882,N_27222,N_27847);
xnor U28883 (N_28883,N_27711,N_27361);
nand U28884 (N_28884,N_27471,N_27407);
or U28885 (N_28885,N_27669,N_27280);
xor U28886 (N_28886,N_27993,N_27624);
nor U28887 (N_28887,N_27089,N_27102);
and U28888 (N_28888,N_27253,N_27499);
xnor U28889 (N_28889,N_27933,N_27842);
or U28890 (N_28890,N_27101,N_27678);
nand U28891 (N_28891,N_27902,N_27886);
or U28892 (N_28892,N_27891,N_27524);
xor U28893 (N_28893,N_27162,N_27323);
xor U28894 (N_28894,N_27100,N_27995);
xnor U28895 (N_28895,N_27652,N_27879);
or U28896 (N_28896,N_27888,N_27892);
nor U28897 (N_28897,N_27817,N_27229);
or U28898 (N_28898,N_27983,N_27055);
nor U28899 (N_28899,N_27016,N_27686);
nand U28900 (N_28900,N_27792,N_27208);
and U28901 (N_28901,N_27654,N_27280);
nand U28902 (N_28902,N_27023,N_27510);
or U28903 (N_28903,N_27654,N_27293);
or U28904 (N_28904,N_27541,N_27980);
and U28905 (N_28905,N_27006,N_27124);
or U28906 (N_28906,N_27435,N_27933);
and U28907 (N_28907,N_27008,N_27410);
nor U28908 (N_28908,N_27216,N_27858);
nand U28909 (N_28909,N_27082,N_27007);
xnor U28910 (N_28910,N_27259,N_27019);
nand U28911 (N_28911,N_27770,N_27978);
nand U28912 (N_28912,N_27253,N_27985);
nor U28913 (N_28913,N_27667,N_27785);
xnor U28914 (N_28914,N_27191,N_27454);
and U28915 (N_28915,N_27576,N_27889);
and U28916 (N_28916,N_27092,N_27726);
nand U28917 (N_28917,N_27324,N_27920);
or U28918 (N_28918,N_27415,N_27756);
nor U28919 (N_28919,N_27581,N_27779);
and U28920 (N_28920,N_27215,N_27707);
nand U28921 (N_28921,N_27474,N_27371);
nand U28922 (N_28922,N_27188,N_27949);
or U28923 (N_28923,N_27016,N_27395);
or U28924 (N_28924,N_27101,N_27132);
nor U28925 (N_28925,N_27793,N_27239);
and U28926 (N_28926,N_27612,N_27324);
and U28927 (N_28927,N_27676,N_27558);
xnor U28928 (N_28928,N_27147,N_27280);
nand U28929 (N_28929,N_27096,N_27224);
and U28930 (N_28930,N_27672,N_27586);
or U28931 (N_28931,N_27293,N_27520);
nor U28932 (N_28932,N_27348,N_27790);
nand U28933 (N_28933,N_27604,N_27110);
or U28934 (N_28934,N_27770,N_27187);
or U28935 (N_28935,N_27534,N_27060);
and U28936 (N_28936,N_27437,N_27018);
nand U28937 (N_28937,N_27980,N_27187);
and U28938 (N_28938,N_27852,N_27459);
nand U28939 (N_28939,N_27814,N_27287);
or U28940 (N_28940,N_27483,N_27042);
and U28941 (N_28941,N_27787,N_27007);
and U28942 (N_28942,N_27845,N_27136);
xnor U28943 (N_28943,N_27893,N_27001);
nor U28944 (N_28944,N_27452,N_27901);
xor U28945 (N_28945,N_27954,N_27177);
and U28946 (N_28946,N_27319,N_27358);
or U28947 (N_28947,N_27264,N_27423);
xnor U28948 (N_28948,N_27786,N_27745);
nand U28949 (N_28949,N_27043,N_27928);
xor U28950 (N_28950,N_27847,N_27788);
nand U28951 (N_28951,N_27564,N_27929);
or U28952 (N_28952,N_27149,N_27115);
xnor U28953 (N_28953,N_27938,N_27218);
nor U28954 (N_28954,N_27116,N_27226);
or U28955 (N_28955,N_27691,N_27494);
nor U28956 (N_28956,N_27373,N_27157);
nand U28957 (N_28957,N_27754,N_27640);
nor U28958 (N_28958,N_27551,N_27266);
and U28959 (N_28959,N_27331,N_27610);
nor U28960 (N_28960,N_27679,N_27417);
nor U28961 (N_28961,N_27035,N_27235);
xnor U28962 (N_28962,N_27075,N_27330);
or U28963 (N_28963,N_27919,N_27119);
xor U28964 (N_28964,N_27651,N_27543);
and U28965 (N_28965,N_27656,N_27952);
or U28966 (N_28966,N_27057,N_27745);
nand U28967 (N_28967,N_27729,N_27071);
nand U28968 (N_28968,N_27149,N_27948);
and U28969 (N_28969,N_27891,N_27039);
and U28970 (N_28970,N_27160,N_27734);
or U28971 (N_28971,N_27614,N_27549);
or U28972 (N_28972,N_27327,N_27574);
xnor U28973 (N_28973,N_27036,N_27037);
xor U28974 (N_28974,N_27790,N_27991);
nor U28975 (N_28975,N_27922,N_27740);
xnor U28976 (N_28976,N_27291,N_27770);
or U28977 (N_28977,N_27247,N_27774);
nor U28978 (N_28978,N_27458,N_27952);
nor U28979 (N_28979,N_27008,N_27266);
and U28980 (N_28980,N_27369,N_27095);
or U28981 (N_28981,N_27465,N_27370);
nor U28982 (N_28982,N_27251,N_27265);
xnor U28983 (N_28983,N_27241,N_27646);
or U28984 (N_28984,N_27579,N_27934);
xor U28985 (N_28985,N_27718,N_27629);
or U28986 (N_28986,N_27351,N_27835);
nor U28987 (N_28987,N_27317,N_27335);
xnor U28988 (N_28988,N_27363,N_27160);
or U28989 (N_28989,N_27915,N_27532);
or U28990 (N_28990,N_27313,N_27849);
nand U28991 (N_28991,N_27685,N_27473);
or U28992 (N_28992,N_27552,N_27057);
xor U28993 (N_28993,N_27342,N_27364);
xnor U28994 (N_28994,N_27327,N_27426);
or U28995 (N_28995,N_27212,N_27527);
nand U28996 (N_28996,N_27067,N_27548);
nor U28997 (N_28997,N_27039,N_27657);
nor U28998 (N_28998,N_27595,N_27038);
or U28999 (N_28999,N_27814,N_27583);
or U29000 (N_29000,N_28621,N_28305);
nand U29001 (N_29001,N_28989,N_28120);
or U29002 (N_29002,N_28761,N_28662);
or U29003 (N_29003,N_28463,N_28406);
and U29004 (N_29004,N_28117,N_28724);
nor U29005 (N_29005,N_28018,N_28592);
and U29006 (N_29006,N_28212,N_28778);
or U29007 (N_29007,N_28666,N_28611);
xnor U29008 (N_29008,N_28960,N_28736);
nor U29009 (N_29009,N_28694,N_28471);
and U29010 (N_29010,N_28162,N_28325);
nand U29011 (N_29011,N_28988,N_28822);
or U29012 (N_29012,N_28740,N_28278);
xnor U29013 (N_29013,N_28226,N_28073);
or U29014 (N_29014,N_28535,N_28399);
and U29015 (N_29015,N_28557,N_28546);
nor U29016 (N_29016,N_28910,N_28404);
or U29017 (N_29017,N_28444,N_28007);
or U29018 (N_29018,N_28764,N_28905);
nor U29019 (N_29019,N_28633,N_28802);
nand U29020 (N_29020,N_28563,N_28532);
nand U29021 (N_29021,N_28958,N_28808);
nand U29022 (N_29022,N_28234,N_28787);
nor U29023 (N_29023,N_28722,N_28575);
nor U29024 (N_29024,N_28338,N_28015);
and U29025 (N_29025,N_28704,N_28883);
xnor U29026 (N_29026,N_28052,N_28811);
nor U29027 (N_29027,N_28119,N_28980);
nor U29028 (N_29028,N_28213,N_28771);
nand U29029 (N_29029,N_28098,N_28997);
nand U29030 (N_29030,N_28555,N_28357);
nand U29031 (N_29031,N_28340,N_28070);
or U29032 (N_29032,N_28919,N_28579);
or U29033 (N_29033,N_28693,N_28613);
or U29034 (N_29034,N_28277,N_28675);
and U29035 (N_29035,N_28914,N_28819);
or U29036 (N_29036,N_28328,N_28653);
nand U29037 (N_29037,N_28135,N_28799);
nor U29038 (N_29038,N_28847,N_28063);
and U29039 (N_29039,N_28986,N_28922);
xnor U29040 (N_29040,N_28195,N_28640);
and U29041 (N_29041,N_28189,N_28295);
or U29042 (N_29042,N_28924,N_28155);
nand U29043 (N_29043,N_28908,N_28042);
or U29044 (N_29044,N_28779,N_28496);
nor U29045 (N_29045,N_28795,N_28522);
or U29046 (N_29046,N_28425,N_28728);
nand U29047 (N_29047,N_28465,N_28450);
nor U29048 (N_29048,N_28279,N_28370);
nor U29049 (N_29049,N_28389,N_28788);
nor U29050 (N_29050,N_28159,N_28805);
nand U29051 (N_29051,N_28210,N_28040);
nand U29052 (N_29052,N_28829,N_28921);
nand U29053 (N_29053,N_28687,N_28826);
nand U29054 (N_29054,N_28060,N_28225);
xor U29055 (N_29055,N_28252,N_28456);
nor U29056 (N_29056,N_28203,N_28747);
nand U29057 (N_29057,N_28880,N_28918);
nor U29058 (N_29058,N_28689,N_28710);
or U29059 (N_29059,N_28056,N_28840);
and U29060 (N_29060,N_28428,N_28623);
or U29061 (N_29061,N_28545,N_28996);
xnor U29062 (N_29062,N_28182,N_28083);
xnor U29063 (N_29063,N_28447,N_28881);
nand U29064 (N_29064,N_28620,N_28390);
nor U29065 (N_29065,N_28319,N_28221);
nand U29066 (N_29066,N_28269,N_28267);
nand U29067 (N_29067,N_28096,N_28616);
nand U29068 (N_29068,N_28048,N_28601);
or U29069 (N_29069,N_28000,N_28153);
nor U29070 (N_29070,N_28172,N_28499);
nand U29071 (N_29071,N_28851,N_28925);
and U29072 (N_29072,N_28928,N_28359);
and U29073 (N_29073,N_28625,N_28410);
xnor U29074 (N_29074,N_28296,N_28538);
and U29075 (N_29075,N_28072,N_28598);
nor U29076 (N_29076,N_28187,N_28849);
and U29077 (N_29077,N_28080,N_28767);
and U29078 (N_29078,N_28109,N_28004);
and U29079 (N_29079,N_28681,N_28092);
nor U29080 (N_29080,N_28594,N_28976);
or U29081 (N_29081,N_28223,N_28937);
xor U29082 (N_29082,N_28176,N_28630);
and U29083 (N_29083,N_28642,N_28421);
nor U29084 (N_29084,N_28917,N_28173);
nand U29085 (N_29085,N_28100,N_28457);
nor U29086 (N_29086,N_28256,N_28397);
nand U29087 (N_29087,N_28049,N_28301);
or U29088 (N_29088,N_28373,N_28418);
or U29089 (N_29089,N_28186,N_28250);
xor U29090 (N_29090,N_28896,N_28263);
and U29091 (N_29091,N_28029,N_28597);
and U29092 (N_29092,N_28346,N_28932);
or U29093 (N_29093,N_28244,N_28130);
nand U29094 (N_29094,N_28141,N_28061);
or U29095 (N_29095,N_28419,N_28243);
nand U29096 (N_29096,N_28344,N_28430);
and U29097 (N_29097,N_28360,N_28230);
nand U29098 (N_29098,N_28035,N_28859);
or U29099 (N_29099,N_28038,N_28401);
and U29100 (N_29100,N_28409,N_28755);
xnor U29101 (N_29101,N_28549,N_28103);
nor U29102 (N_29102,N_28750,N_28132);
nor U29103 (N_29103,N_28490,N_28517);
and U29104 (N_29104,N_28426,N_28364);
or U29105 (N_29105,N_28206,N_28509);
xor U29106 (N_29106,N_28032,N_28909);
nor U29107 (N_29107,N_28864,N_28715);
and U29108 (N_29108,N_28797,N_28125);
nor U29109 (N_29109,N_28468,N_28129);
xor U29110 (N_29110,N_28139,N_28233);
or U29111 (N_29111,N_28031,N_28235);
or U29112 (N_29112,N_28671,N_28887);
nor U29113 (N_29113,N_28588,N_28743);
xnor U29114 (N_29114,N_28804,N_28238);
xnor U29115 (N_29115,N_28494,N_28054);
or U29116 (N_29116,N_28564,N_28984);
or U29117 (N_29117,N_28962,N_28565);
nand U29118 (N_29118,N_28712,N_28383);
or U29119 (N_29119,N_28758,N_28116);
xor U29120 (N_29120,N_28923,N_28765);
xor U29121 (N_29121,N_28991,N_28264);
xor U29122 (N_29122,N_28998,N_28138);
xor U29123 (N_29123,N_28122,N_28615);
or U29124 (N_29124,N_28580,N_28348);
and U29125 (N_29125,N_28491,N_28034);
and U29126 (N_29126,N_28593,N_28515);
nand U29127 (N_29127,N_28003,N_28508);
xor U29128 (N_29128,N_28570,N_28807);
and U29129 (N_29129,N_28610,N_28907);
nor U29130 (N_29130,N_28144,N_28773);
nor U29131 (N_29131,N_28014,N_28474);
nor U29132 (N_29132,N_28201,N_28574);
or U29133 (N_29133,N_28664,N_28302);
nand U29134 (N_29134,N_28553,N_28744);
or U29135 (N_29135,N_28059,N_28420);
or U29136 (N_29136,N_28703,N_28618);
or U29137 (N_29137,N_28500,N_28275);
xor U29138 (N_29138,N_28151,N_28794);
nand U29139 (N_29139,N_28867,N_28118);
xnor U29140 (N_29140,N_28249,N_28013);
or U29141 (N_29141,N_28875,N_28803);
nor U29142 (N_29142,N_28090,N_28957);
nand U29143 (N_29143,N_28432,N_28916);
and U29144 (N_29144,N_28483,N_28165);
nand U29145 (N_29145,N_28951,N_28197);
nor U29146 (N_29146,N_28403,N_28241);
nor U29147 (N_29147,N_28478,N_28486);
nor U29148 (N_29148,N_28770,N_28314);
nor U29149 (N_29149,N_28208,N_28429);
nor U29150 (N_29150,N_28273,N_28502);
and U29151 (N_29151,N_28837,N_28475);
nor U29152 (N_29152,N_28583,N_28652);
or U29153 (N_29153,N_28733,N_28774);
nand U29154 (N_29154,N_28326,N_28115);
nand U29155 (N_29155,N_28303,N_28461);
nor U29156 (N_29156,N_28091,N_28068);
and U29157 (N_29157,N_28408,N_28436);
and U29158 (N_29158,N_28940,N_28530);
and U29159 (N_29159,N_28431,N_28622);
and U29160 (N_29160,N_28396,N_28683);
nand U29161 (N_29161,N_28738,N_28350);
xnor U29162 (N_29162,N_28441,N_28608);
nor U29163 (N_29163,N_28796,N_28493);
nor U29164 (N_29164,N_28965,N_28516);
or U29165 (N_29165,N_28691,N_28595);
nor U29166 (N_29166,N_28892,N_28634);
xnor U29167 (N_29167,N_28832,N_28933);
nand U29168 (N_29168,N_28413,N_28284);
and U29169 (N_29169,N_28143,N_28523);
nand U29170 (N_29170,N_28395,N_28462);
nand U29171 (N_29171,N_28150,N_28414);
nor U29172 (N_29172,N_28894,N_28087);
and U29173 (N_29173,N_28518,N_28198);
and U29174 (N_29174,N_28558,N_28596);
or U29175 (N_29175,N_28676,N_28639);
nor U29176 (N_29176,N_28424,N_28873);
nor U29177 (N_29177,N_28775,N_28946);
or U29178 (N_29178,N_28351,N_28028);
nand U29179 (N_29179,N_28655,N_28154);
nor U29180 (N_29180,N_28607,N_28262);
and U29181 (N_29181,N_28020,N_28635);
or U29182 (N_29182,N_28086,N_28260);
xnor U29183 (N_29183,N_28169,N_28503);
and U29184 (N_29184,N_28245,N_28714);
xor U29185 (N_29185,N_28854,N_28551);
and U29186 (N_29186,N_28720,N_28813);
nor U29187 (N_29187,N_28547,N_28355);
nand U29188 (N_29188,N_28349,N_28372);
xnor U29189 (N_29189,N_28524,N_28816);
or U29190 (N_29190,N_28079,N_28232);
or U29191 (N_29191,N_28320,N_28985);
xnor U29192 (N_29192,N_28137,N_28205);
nor U29193 (N_29193,N_28757,N_28104);
nor U29194 (N_29194,N_28239,N_28845);
nand U29195 (N_29195,N_28037,N_28077);
nor U29196 (N_29196,N_28412,N_28973);
nor U29197 (N_29197,N_28809,N_28696);
xnor U29198 (N_29198,N_28217,N_28181);
nor U29199 (N_29199,N_28011,N_28046);
and U29200 (N_29200,N_28812,N_28300);
nand U29201 (N_29201,N_28053,N_28285);
or U29202 (N_29202,N_28888,N_28171);
or U29203 (N_29203,N_28573,N_28862);
xnor U29204 (N_29204,N_28097,N_28879);
xnor U29205 (N_29205,N_28900,N_28204);
and U29206 (N_29206,N_28170,N_28484);
nor U29207 (N_29207,N_28392,N_28834);
xor U29208 (N_29208,N_28184,N_28654);
nor U29209 (N_29209,N_28307,N_28646);
nor U29210 (N_29210,N_28990,N_28836);
xor U29211 (N_29211,N_28352,N_28612);
or U29212 (N_29212,N_28339,N_28790);
and U29213 (N_29213,N_28776,N_28663);
or U29214 (N_29214,N_28378,N_28711);
xnor U29215 (N_29215,N_28669,N_28271);
or U29216 (N_29216,N_28216,N_28734);
nor U29217 (N_29217,N_28614,N_28163);
and U29218 (N_29218,N_28566,N_28741);
xor U29219 (N_29219,N_28199,N_28058);
or U29220 (N_29220,N_28148,N_28308);
nand U29221 (N_29221,N_28999,N_28342);
nand U29222 (N_29222,N_28178,N_28248);
xnor U29223 (N_29223,N_28036,N_28876);
xnor U29224 (N_29224,N_28030,N_28679);
nor U29225 (N_29225,N_28543,N_28247);
xnor U29226 (N_29226,N_28433,N_28619);
xnor U29227 (N_29227,N_28820,N_28541);
nor U29228 (N_29228,N_28912,N_28697);
nor U29229 (N_29229,N_28071,N_28394);
nor U29230 (N_29230,N_28719,N_28763);
nand U29231 (N_29231,N_28782,N_28064);
or U29232 (N_29232,N_28857,N_28361);
or U29233 (N_29233,N_28180,N_28974);
nor U29234 (N_29234,N_28707,N_28648);
or U29235 (N_29235,N_28033,N_28511);
and U29236 (N_29236,N_28993,N_28982);
nor U29237 (N_29237,N_28971,N_28236);
xnor U29238 (N_29238,N_28047,N_28514);
nand U29239 (N_29239,N_28131,N_28582);
and U29240 (N_29240,N_28823,N_28938);
and U29241 (N_29241,N_28731,N_28067);
nor U29242 (N_29242,N_28581,N_28629);
xnor U29243 (N_29243,N_28402,N_28016);
and U29244 (N_29244,N_28477,N_28057);
and U29245 (N_29245,N_28435,N_28688);
nor U29246 (N_29246,N_28954,N_28334);
and U29247 (N_29247,N_28886,N_28878);
nand U29248 (N_29248,N_28605,N_28085);
nor U29249 (N_29249,N_28602,N_28786);
or U29250 (N_29250,N_28560,N_28229);
or U29251 (N_29251,N_28228,N_28705);
nand U29252 (N_29252,N_28529,N_28631);
nor U29253 (N_29253,N_28175,N_28944);
or U29254 (N_29254,N_28684,N_28084);
xnor U29255 (N_29255,N_28737,N_28762);
and U29256 (N_29256,N_28202,N_28112);
xor U29257 (N_29257,N_28113,N_28959);
xor U29258 (N_29258,N_28008,N_28191);
or U29259 (N_29259,N_28994,N_28536);
nor U29260 (N_29260,N_28146,N_28968);
nand U29261 (N_29261,N_28472,N_28088);
xnor U29262 (N_29262,N_28211,N_28473);
nand U29263 (N_29263,N_28017,N_28855);
and U29264 (N_29264,N_28495,N_28480);
or U29265 (N_29265,N_28453,N_28214);
xor U29266 (N_29266,N_28281,N_28405);
or U29267 (N_29267,N_28953,N_28901);
or U29268 (N_29268,N_28665,N_28293);
or U29269 (N_29269,N_28780,N_28254);
xor U29270 (N_29270,N_28843,N_28542);
xnor U29271 (N_29271,N_28891,N_28386);
or U29272 (N_29272,N_28824,N_28074);
nor U29273 (N_29273,N_28082,N_28865);
xnor U29274 (N_29274,N_28931,N_28266);
xnor U29275 (N_29275,N_28445,N_28835);
nand U29276 (N_29276,N_28161,N_28200);
nor U29277 (N_29277,N_28667,N_28895);
nor U29278 (N_29278,N_28945,N_28527);
nand U29279 (N_29279,N_28259,N_28488);
xor U29280 (N_29280,N_28627,N_28603);
nor U29281 (N_29281,N_28709,N_28019);
or U29282 (N_29282,N_28680,N_28793);
and U29283 (N_29283,N_28967,N_28391);
xnor U29284 (N_29284,N_28045,N_28806);
nor U29285 (N_29285,N_28830,N_28505);
xor U29286 (N_29286,N_28833,N_28587);
or U29287 (N_29287,N_28686,N_28479);
nor U29288 (N_29288,N_28699,N_28858);
or U29289 (N_29289,N_28449,N_28481);
nor U29290 (N_29290,N_28814,N_28026);
and U29291 (N_29291,N_28730,N_28860);
nor U29292 (N_29292,N_28193,N_28578);
or U29293 (N_29293,N_28321,N_28981);
nand U29294 (N_29294,N_28800,N_28632);
and U29295 (N_29295,N_28539,N_28044);
nand U29296 (N_29296,N_28489,N_28550);
nand U29297 (N_29297,N_28911,N_28651);
nor U29298 (N_29298,N_28739,N_28643);
xnor U29299 (N_29299,N_28673,N_28287);
nor U29300 (N_29300,N_28451,N_28852);
nand U29301 (N_29301,N_28388,N_28936);
and U29302 (N_29302,N_28220,N_28685);
or U29303 (N_29303,N_28955,N_28427);
xnor U29304 (N_29304,N_28745,N_28102);
nand U29305 (N_29305,N_28218,N_28291);
or U29306 (N_29306,N_28561,N_28963);
nor U29307 (N_29307,N_28567,N_28136);
nand U29308 (N_29308,N_28889,N_28751);
xor U29309 (N_29309,N_28604,N_28158);
and U29310 (N_29310,N_28591,N_28874);
nor U29311 (N_29311,N_28368,N_28363);
xnor U29312 (N_29312,N_28012,N_28906);
or U29313 (N_29313,N_28825,N_28975);
or U29314 (N_29314,N_28487,N_28310);
xor U29315 (N_29315,N_28341,N_28298);
nand U29316 (N_29316,N_28838,N_28345);
and U29317 (N_29317,N_28915,N_28358);
nand U29318 (N_29318,N_28682,N_28149);
nand U29319 (N_29319,N_28979,N_28124);
or U29320 (N_29320,N_28853,N_28898);
nor U29321 (N_29321,N_28306,N_28177);
nor U29322 (N_29322,N_28785,N_28466);
xor U29323 (N_29323,N_28939,N_28526);
xnor U29324 (N_29324,N_28600,N_28270);
and U29325 (N_29325,N_28385,N_28884);
and U29326 (N_29326,N_28970,N_28010);
xor U29327 (N_29327,N_28768,N_28777);
or U29328 (N_29328,N_28987,N_28374);
nor U29329 (N_29329,N_28972,N_28265);
nand U29330 (N_29330,N_28766,N_28842);
and U29331 (N_29331,N_28961,N_28152);
nand U29332 (N_29332,N_28941,N_28400);
nor U29333 (N_29333,N_28382,N_28448);
xor U29334 (N_29334,N_28258,N_28369);
or U29335 (N_29335,N_28817,N_28659);
nor U29336 (N_29336,N_28644,N_28164);
nor U29337 (N_29337,N_28443,N_28268);
nand U29338 (N_29338,N_28661,N_28492);
xor U29339 (N_29339,N_28280,N_28668);
or U29340 (N_29340,N_28167,N_28950);
nand U29341 (N_29341,N_28274,N_28781);
nand U29342 (N_29342,N_28706,N_28868);
or U29343 (N_29343,N_28726,N_28095);
and U29344 (N_29344,N_28123,N_28160);
or U29345 (N_29345,N_28882,N_28393);
and U29346 (N_29346,N_28801,N_28670);
or U29347 (N_29347,N_28528,N_28869);
xor U29348 (N_29348,N_28927,N_28188);
xnor U29349 (N_29349,N_28147,N_28498);
nor U29350 (N_29350,N_28460,N_28798);
xnor U29351 (N_29351,N_28562,N_28043);
or U29352 (N_29352,N_28890,N_28365);
and U29353 (N_29353,N_28041,N_28930);
nand U29354 (N_29354,N_28647,N_28772);
nand U29355 (N_29355,N_28168,N_28025);
nor U29356 (N_29356,N_28183,N_28324);
nor U29357 (N_29357,N_28556,N_28069);
xor U29358 (N_29358,N_28128,N_28005);
or U29359 (N_29359,N_28075,N_28437);
and U29360 (N_29360,N_28754,N_28501);
and U29361 (N_29361,N_28039,N_28133);
nand U29362 (N_29362,N_28827,N_28375);
nand U29363 (N_29363,N_28134,N_28947);
xor U29364 (N_29364,N_28948,N_28081);
xor U29365 (N_29365,N_28343,N_28729);
or U29366 (N_29366,N_28742,N_28335);
nor U29367 (N_29367,N_28455,N_28089);
nand U29368 (N_29368,N_28126,N_28789);
xor U29369 (N_29369,N_28690,N_28354);
xnor U29370 (N_29370,N_28554,N_28617);
or U29371 (N_29371,N_28966,N_28559);
nand U29372 (N_29372,N_28657,N_28194);
and U29373 (N_29373,N_28283,N_28815);
and U29374 (N_29374,N_28899,N_28288);
nor U29375 (N_29375,N_28756,N_28952);
nand U29376 (N_29376,N_28590,N_28784);
xor U29377 (N_29377,N_28377,N_28387);
or U29378 (N_29378,N_28844,N_28371);
nand U29379 (N_29379,N_28099,N_28330);
nor U29380 (N_29380,N_28871,N_28848);
xnor U29381 (N_29381,N_28577,N_28272);
xor U29382 (N_29382,N_28695,N_28992);
and U29383 (N_29383,N_28407,N_28367);
or U29384 (N_29384,N_28841,N_28534);
xnor U29385 (N_29385,N_28913,N_28105);
xnor U29386 (N_29386,N_28521,N_28347);
nand U29387 (N_29387,N_28943,N_28190);
nand U29388 (N_29388,N_28094,N_28692);
xor U29389 (N_29389,N_28196,N_28312);
or U29390 (N_29390,N_28585,N_28628);
and U29391 (N_29391,N_28818,N_28584);
nand U29392 (N_29392,N_28791,N_28513);
nor U29393 (N_29393,N_28902,N_28166);
nor U29394 (N_29394,N_28251,N_28318);
xnor U29395 (N_29395,N_28519,N_28304);
nor U29396 (N_29396,N_28062,N_28626);
or U29397 (N_29397,N_28353,N_28856);
nor U29398 (N_29398,N_28893,N_28609);
nand U29399 (N_29399,N_28411,N_28897);
or U29400 (N_29400,N_28446,N_28356);
xor U29401 (N_29401,N_28309,N_28713);
and U29402 (N_29402,N_28219,N_28145);
nor U29403 (N_29403,N_28290,N_28066);
nand U29404 (N_29404,N_28641,N_28009);
xnor U29405 (N_29405,N_28255,N_28716);
nor U29406 (N_29406,N_28006,N_28322);
nand U29407 (N_29407,N_28110,N_28942);
or U29408 (N_29408,N_28485,N_28674);
xnor U29409 (N_29409,N_28650,N_28442);
xor U29410 (N_29410,N_28752,N_28289);
nand U29411 (N_29411,N_28828,N_28022);
and U29412 (N_29412,N_28531,N_28636);
xor U29413 (N_29413,N_28544,N_28076);
nor U29414 (N_29414,N_28440,N_28415);
xnor U29415 (N_29415,N_28101,N_28949);
xnor U29416 (N_29416,N_28329,N_28292);
nor U29417 (N_29417,N_28174,N_28156);
nor U29418 (N_29418,N_28246,N_28111);
xnor U29419 (N_29419,N_28956,N_28157);
or U29420 (N_29420,N_28261,N_28753);
nand U29421 (N_29421,N_28540,N_28434);
nand U29422 (N_29422,N_28732,N_28336);
nand U29423 (N_29423,N_28525,N_28242);
or U29424 (N_29424,N_28055,N_28331);
nand U29425 (N_29425,N_28381,N_28380);
and U29426 (N_29426,N_28571,N_28315);
and U29427 (N_29427,N_28850,N_28866);
nand U29428 (N_29428,N_28759,N_28439);
nor U29429 (N_29429,N_28746,N_28257);
or U29430 (N_29430,N_28727,N_28332);
xor U29431 (N_29431,N_28645,N_28995);
nand U29432 (N_29432,N_28701,N_28660);
or U29433 (N_29433,N_28964,N_28452);
or U29434 (N_29434,N_28376,N_28969);
nor U29435 (N_29435,N_28422,N_28839);
nand U29436 (N_29436,N_28885,N_28209);
and U29437 (N_29437,N_28237,N_28192);
or U29438 (N_29438,N_28624,N_28783);
nand U29439 (N_29439,N_28537,N_28467);
and U29440 (N_29440,N_28977,N_28438);
or U29441 (N_29441,N_28586,N_28311);
or U29442 (N_29442,N_28276,N_28333);
nand U29443 (N_29443,N_28735,N_28224);
xor U29444 (N_29444,N_28398,N_28337);
xor U29445 (N_29445,N_28708,N_28978);
nor U29446 (N_29446,N_28464,N_28846);
nor U29447 (N_29447,N_28533,N_28677);
nand U29448 (N_29448,N_28903,N_28106);
nor U29449 (N_29449,N_28114,N_28215);
nand U29450 (N_29450,N_28904,N_28185);
and U29451 (N_29451,N_28725,N_28821);
nor U29452 (N_29452,N_28286,N_28861);
and U29453 (N_29453,N_28327,N_28497);
nor U29454 (N_29454,N_28506,N_28127);
and U29455 (N_29455,N_28142,N_28638);
and U29456 (N_29456,N_28459,N_28379);
nor U29457 (N_29457,N_28872,N_28576);
xnor U29458 (N_29458,N_28929,N_28934);
nor U29459 (N_29459,N_28672,N_28294);
xor U29460 (N_29460,N_28323,N_28027);
or U29461 (N_29461,N_28760,N_28926);
xor U29462 (N_29462,N_28606,N_28108);
xnor U29463 (N_29463,N_28983,N_28749);
nand U29464 (N_29464,N_28316,N_28482);
or U29465 (N_29465,N_28282,N_28678);
xor U29466 (N_29466,N_28810,N_28572);
and U29467 (N_29467,N_28510,N_28416);
xor U29468 (N_29468,N_28227,N_28568);
xnor U29469 (N_29469,N_28179,N_28051);
nand U29470 (N_29470,N_28222,N_28792);
xor U29471 (N_29471,N_28458,N_28240);
or U29472 (N_29472,N_28050,N_28920);
and U29473 (N_29473,N_28935,N_28384);
nand U29474 (N_29474,N_28702,N_28552);
or U29475 (N_29475,N_28065,N_28093);
or U29476 (N_29476,N_28718,N_28721);
and U29477 (N_29477,N_28024,N_28121);
xor U29478 (N_29478,N_28504,N_28313);
nor U29479 (N_29479,N_28548,N_28417);
and U29480 (N_29480,N_28512,N_28021);
nand U29481 (N_29481,N_28317,N_28078);
nand U29482 (N_29482,N_28297,N_28454);
xnor U29483 (N_29483,N_28231,N_28362);
and U29484 (N_29484,N_28207,N_28423);
and U29485 (N_29485,N_28470,N_28700);
and U29486 (N_29486,N_28658,N_28520);
xor U29487 (N_29487,N_28717,N_28507);
xor U29488 (N_29488,N_28476,N_28637);
xor U29489 (N_29489,N_28140,N_28569);
nand U29490 (N_29490,N_28366,N_28002);
or U29491 (N_29491,N_28107,N_28723);
nand U29492 (N_29492,N_28870,N_28649);
xnor U29493 (N_29493,N_28253,N_28299);
and U29494 (N_29494,N_28656,N_28589);
nor U29495 (N_29495,N_28023,N_28599);
and U29496 (N_29496,N_28698,N_28831);
xor U29497 (N_29497,N_28863,N_28769);
nor U29498 (N_29498,N_28748,N_28469);
xor U29499 (N_29499,N_28001,N_28877);
or U29500 (N_29500,N_28424,N_28117);
or U29501 (N_29501,N_28742,N_28399);
xor U29502 (N_29502,N_28072,N_28231);
or U29503 (N_29503,N_28977,N_28499);
or U29504 (N_29504,N_28658,N_28170);
nor U29505 (N_29505,N_28932,N_28317);
or U29506 (N_29506,N_28788,N_28170);
nand U29507 (N_29507,N_28267,N_28970);
nand U29508 (N_29508,N_28250,N_28607);
xor U29509 (N_29509,N_28626,N_28094);
or U29510 (N_29510,N_28434,N_28513);
or U29511 (N_29511,N_28343,N_28227);
and U29512 (N_29512,N_28248,N_28914);
nor U29513 (N_29513,N_28241,N_28901);
nor U29514 (N_29514,N_28351,N_28084);
and U29515 (N_29515,N_28011,N_28352);
nor U29516 (N_29516,N_28179,N_28824);
nor U29517 (N_29517,N_28619,N_28046);
nand U29518 (N_29518,N_28395,N_28243);
xor U29519 (N_29519,N_28456,N_28212);
xor U29520 (N_29520,N_28760,N_28092);
nand U29521 (N_29521,N_28324,N_28157);
nor U29522 (N_29522,N_28374,N_28501);
and U29523 (N_29523,N_28118,N_28290);
nor U29524 (N_29524,N_28238,N_28833);
or U29525 (N_29525,N_28525,N_28715);
and U29526 (N_29526,N_28715,N_28340);
nor U29527 (N_29527,N_28039,N_28905);
and U29528 (N_29528,N_28430,N_28529);
nor U29529 (N_29529,N_28089,N_28879);
nor U29530 (N_29530,N_28127,N_28349);
nor U29531 (N_29531,N_28715,N_28862);
nand U29532 (N_29532,N_28462,N_28229);
nand U29533 (N_29533,N_28732,N_28369);
xor U29534 (N_29534,N_28174,N_28175);
nor U29535 (N_29535,N_28306,N_28160);
nor U29536 (N_29536,N_28773,N_28091);
xor U29537 (N_29537,N_28862,N_28433);
nor U29538 (N_29538,N_28122,N_28528);
nand U29539 (N_29539,N_28395,N_28314);
nand U29540 (N_29540,N_28338,N_28098);
and U29541 (N_29541,N_28397,N_28533);
nor U29542 (N_29542,N_28516,N_28710);
xor U29543 (N_29543,N_28552,N_28109);
xnor U29544 (N_29544,N_28279,N_28707);
nand U29545 (N_29545,N_28806,N_28222);
nand U29546 (N_29546,N_28024,N_28955);
nor U29547 (N_29547,N_28489,N_28461);
nor U29548 (N_29548,N_28631,N_28316);
and U29549 (N_29549,N_28723,N_28444);
and U29550 (N_29550,N_28480,N_28966);
or U29551 (N_29551,N_28427,N_28872);
and U29552 (N_29552,N_28761,N_28136);
nor U29553 (N_29553,N_28185,N_28210);
nor U29554 (N_29554,N_28980,N_28293);
xor U29555 (N_29555,N_28469,N_28312);
nand U29556 (N_29556,N_28863,N_28464);
and U29557 (N_29557,N_28963,N_28294);
and U29558 (N_29558,N_28303,N_28049);
xnor U29559 (N_29559,N_28406,N_28212);
xor U29560 (N_29560,N_28539,N_28058);
xor U29561 (N_29561,N_28746,N_28605);
nor U29562 (N_29562,N_28948,N_28623);
nand U29563 (N_29563,N_28617,N_28173);
nor U29564 (N_29564,N_28685,N_28500);
xor U29565 (N_29565,N_28373,N_28302);
nor U29566 (N_29566,N_28423,N_28568);
nand U29567 (N_29567,N_28820,N_28825);
nor U29568 (N_29568,N_28498,N_28395);
and U29569 (N_29569,N_28030,N_28032);
nand U29570 (N_29570,N_28870,N_28134);
nand U29571 (N_29571,N_28364,N_28510);
xnor U29572 (N_29572,N_28034,N_28650);
or U29573 (N_29573,N_28827,N_28486);
or U29574 (N_29574,N_28163,N_28378);
xnor U29575 (N_29575,N_28811,N_28943);
nand U29576 (N_29576,N_28359,N_28696);
xnor U29577 (N_29577,N_28132,N_28481);
nor U29578 (N_29578,N_28089,N_28447);
or U29579 (N_29579,N_28799,N_28569);
xor U29580 (N_29580,N_28607,N_28898);
and U29581 (N_29581,N_28330,N_28350);
and U29582 (N_29582,N_28317,N_28356);
and U29583 (N_29583,N_28862,N_28955);
xnor U29584 (N_29584,N_28914,N_28789);
xnor U29585 (N_29585,N_28076,N_28912);
xnor U29586 (N_29586,N_28482,N_28936);
xnor U29587 (N_29587,N_28857,N_28861);
nand U29588 (N_29588,N_28982,N_28505);
xnor U29589 (N_29589,N_28248,N_28039);
or U29590 (N_29590,N_28329,N_28771);
or U29591 (N_29591,N_28202,N_28927);
xnor U29592 (N_29592,N_28317,N_28793);
nand U29593 (N_29593,N_28868,N_28536);
xor U29594 (N_29594,N_28706,N_28884);
or U29595 (N_29595,N_28831,N_28887);
and U29596 (N_29596,N_28969,N_28943);
and U29597 (N_29597,N_28318,N_28494);
nor U29598 (N_29598,N_28625,N_28445);
xnor U29599 (N_29599,N_28949,N_28627);
nand U29600 (N_29600,N_28301,N_28226);
or U29601 (N_29601,N_28983,N_28176);
xnor U29602 (N_29602,N_28245,N_28984);
and U29603 (N_29603,N_28382,N_28948);
nor U29604 (N_29604,N_28135,N_28127);
and U29605 (N_29605,N_28186,N_28060);
xor U29606 (N_29606,N_28251,N_28369);
xor U29607 (N_29607,N_28268,N_28294);
nor U29608 (N_29608,N_28582,N_28016);
xor U29609 (N_29609,N_28934,N_28347);
xor U29610 (N_29610,N_28457,N_28372);
xnor U29611 (N_29611,N_28100,N_28691);
and U29612 (N_29612,N_28428,N_28494);
nor U29613 (N_29613,N_28712,N_28231);
xnor U29614 (N_29614,N_28687,N_28843);
nor U29615 (N_29615,N_28430,N_28912);
and U29616 (N_29616,N_28408,N_28578);
and U29617 (N_29617,N_28598,N_28419);
nand U29618 (N_29618,N_28402,N_28650);
nand U29619 (N_29619,N_28543,N_28280);
and U29620 (N_29620,N_28662,N_28312);
and U29621 (N_29621,N_28937,N_28262);
and U29622 (N_29622,N_28246,N_28478);
or U29623 (N_29623,N_28775,N_28479);
or U29624 (N_29624,N_28333,N_28979);
or U29625 (N_29625,N_28320,N_28091);
or U29626 (N_29626,N_28388,N_28420);
xor U29627 (N_29627,N_28117,N_28191);
xnor U29628 (N_29628,N_28966,N_28744);
and U29629 (N_29629,N_28469,N_28108);
xnor U29630 (N_29630,N_28194,N_28101);
or U29631 (N_29631,N_28003,N_28614);
nor U29632 (N_29632,N_28062,N_28686);
nor U29633 (N_29633,N_28810,N_28709);
and U29634 (N_29634,N_28811,N_28412);
and U29635 (N_29635,N_28596,N_28217);
nand U29636 (N_29636,N_28978,N_28539);
and U29637 (N_29637,N_28920,N_28253);
nand U29638 (N_29638,N_28602,N_28446);
and U29639 (N_29639,N_28304,N_28373);
xor U29640 (N_29640,N_28111,N_28349);
nand U29641 (N_29641,N_28445,N_28410);
nand U29642 (N_29642,N_28011,N_28447);
nand U29643 (N_29643,N_28790,N_28847);
or U29644 (N_29644,N_28079,N_28938);
xnor U29645 (N_29645,N_28195,N_28926);
and U29646 (N_29646,N_28835,N_28230);
or U29647 (N_29647,N_28516,N_28283);
xor U29648 (N_29648,N_28270,N_28584);
nor U29649 (N_29649,N_28294,N_28813);
and U29650 (N_29650,N_28001,N_28755);
nand U29651 (N_29651,N_28361,N_28218);
nand U29652 (N_29652,N_28368,N_28921);
nor U29653 (N_29653,N_28601,N_28169);
and U29654 (N_29654,N_28989,N_28767);
or U29655 (N_29655,N_28247,N_28660);
xnor U29656 (N_29656,N_28138,N_28184);
or U29657 (N_29657,N_28492,N_28234);
or U29658 (N_29658,N_28774,N_28782);
xor U29659 (N_29659,N_28414,N_28494);
xnor U29660 (N_29660,N_28157,N_28264);
and U29661 (N_29661,N_28499,N_28640);
nand U29662 (N_29662,N_28809,N_28256);
nor U29663 (N_29663,N_28589,N_28343);
nor U29664 (N_29664,N_28728,N_28459);
xnor U29665 (N_29665,N_28542,N_28886);
or U29666 (N_29666,N_28679,N_28182);
nand U29667 (N_29667,N_28133,N_28286);
and U29668 (N_29668,N_28821,N_28779);
nand U29669 (N_29669,N_28556,N_28316);
and U29670 (N_29670,N_28151,N_28496);
xor U29671 (N_29671,N_28747,N_28310);
or U29672 (N_29672,N_28363,N_28749);
nor U29673 (N_29673,N_28721,N_28412);
xor U29674 (N_29674,N_28746,N_28522);
nor U29675 (N_29675,N_28517,N_28336);
and U29676 (N_29676,N_28912,N_28259);
and U29677 (N_29677,N_28756,N_28796);
and U29678 (N_29678,N_28663,N_28933);
nor U29679 (N_29679,N_28915,N_28419);
or U29680 (N_29680,N_28463,N_28531);
nor U29681 (N_29681,N_28011,N_28947);
or U29682 (N_29682,N_28928,N_28627);
nand U29683 (N_29683,N_28537,N_28239);
xor U29684 (N_29684,N_28175,N_28598);
nor U29685 (N_29685,N_28274,N_28579);
and U29686 (N_29686,N_28709,N_28585);
nor U29687 (N_29687,N_28250,N_28145);
and U29688 (N_29688,N_28792,N_28764);
and U29689 (N_29689,N_28944,N_28154);
nor U29690 (N_29690,N_28342,N_28573);
nor U29691 (N_29691,N_28142,N_28160);
nor U29692 (N_29692,N_28477,N_28926);
xnor U29693 (N_29693,N_28046,N_28188);
or U29694 (N_29694,N_28758,N_28620);
and U29695 (N_29695,N_28358,N_28037);
or U29696 (N_29696,N_28624,N_28248);
nor U29697 (N_29697,N_28812,N_28323);
xnor U29698 (N_29698,N_28308,N_28698);
nor U29699 (N_29699,N_28518,N_28572);
nor U29700 (N_29700,N_28480,N_28680);
nand U29701 (N_29701,N_28650,N_28817);
or U29702 (N_29702,N_28692,N_28409);
or U29703 (N_29703,N_28501,N_28197);
xor U29704 (N_29704,N_28038,N_28977);
nand U29705 (N_29705,N_28935,N_28477);
or U29706 (N_29706,N_28933,N_28794);
nand U29707 (N_29707,N_28760,N_28073);
and U29708 (N_29708,N_28549,N_28943);
and U29709 (N_29709,N_28164,N_28790);
xor U29710 (N_29710,N_28589,N_28417);
nand U29711 (N_29711,N_28749,N_28147);
xnor U29712 (N_29712,N_28178,N_28724);
xnor U29713 (N_29713,N_28259,N_28224);
nand U29714 (N_29714,N_28293,N_28620);
or U29715 (N_29715,N_28061,N_28176);
or U29716 (N_29716,N_28443,N_28524);
nor U29717 (N_29717,N_28177,N_28168);
or U29718 (N_29718,N_28158,N_28179);
xnor U29719 (N_29719,N_28449,N_28134);
or U29720 (N_29720,N_28634,N_28697);
or U29721 (N_29721,N_28444,N_28008);
and U29722 (N_29722,N_28119,N_28048);
xnor U29723 (N_29723,N_28814,N_28479);
or U29724 (N_29724,N_28585,N_28795);
nand U29725 (N_29725,N_28893,N_28067);
or U29726 (N_29726,N_28321,N_28496);
nand U29727 (N_29727,N_28062,N_28835);
or U29728 (N_29728,N_28798,N_28658);
and U29729 (N_29729,N_28234,N_28238);
nand U29730 (N_29730,N_28832,N_28938);
nor U29731 (N_29731,N_28981,N_28980);
or U29732 (N_29732,N_28718,N_28681);
nor U29733 (N_29733,N_28065,N_28156);
nor U29734 (N_29734,N_28475,N_28031);
nand U29735 (N_29735,N_28673,N_28992);
xnor U29736 (N_29736,N_28187,N_28049);
nor U29737 (N_29737,N_28365,N_28096);
nand U29738 (N_29738,N_28806,N_28125);
and U29739 (N_29739,N_28260,N_28661);
xor U29740 (N_29740,N_28799,N_28186);
nand U29741 (N_29741,N_28928,N_28516);
or U29742 (N_29742,N_28023,N_28447);
and U29743 (N_29743,N_28524,N_28517);
xor U29744 (N_29744,N_28198,N_28546);
nand U29745 (N_29745,N_28387,N_28547);
nor U29746 (N_29746,N_28054,N_28134);
nand U29747 (N_29747,N_28467,N_28162);
xor U29748 (N_29748,N_28754,N_28877);
nand U29749 (N_29749,N_28996,N_28566);
or U29750 (N_29750,N_28914,N_28374);
and U29751 (N_29751,N_28947,N_28629);
or U29752 (N_29752,N_28308,N_28828);
nand U29753 (N_29753,N_28767,N_28639);
nor U29754 (N_29754,N_28916,N_28192);
or U29755 (N_29755,N_28674,N_28707);
or U29756 (N_29756,N_28158,N_28620);
nand U29757 (N_29757,N_28818,N_28364);
nand U29758 (N_29758,N_28988,N_28294);
and U29759 (N_29759,N_28005,N_28439);
or U29760 (N_29760,N_28141,N_28343);
xor U29761 (N_29761,N_28413,N_28041);
xnor U29762 (N_29762,N_28695,N_28107);
nor U29763 (N_29763,N_28722,N_28001);
and U29764 (N_29764,N_28161,N_28328);
nor U29765 (N_29765,N_28308,N_28797);
and U29766 (N_29766,N_28090,N_28467);
and U29767 (N_29767,N_28295,N_28499);
nor U29768 (N_29768,N_28765,N_28140);
and U29769 (N_29769,N_28746,N_28188);
or U29770 (N_29770,N_28303,N_28171);
xor U29771 (N_29771,N_28046,N_28525);
xor U29772 (N_29772,N_28013,N_28651);
nand U29773 (N_29773,N_28994,N_28927);
nand U29774 (N_29774,N_28889,N_28709);
and U29775 (N_29775,N_28422,N_28571);
nand U29776 (N_29776,N_28645,N_28938);
nand U29777 (N_29777,N_28859,N_28703);
or U29778 (N_29778,N_28196,N_28502);
xnor U29779 (N_29779,N_28504,N_28501);
nand U29780 (N_29780,N_28879,N_28717);
nor U29781 (N_29781,N_28887,N_28465);
nor U29782 (N_29782,N_28138,N_28312);
xnor U29783 (N_29783,N_28555,N_28012);
nor U29784 (N_29784,N_28147,N_28217);
or U29785 (N_29785,N_28214,N_28572);
nand U29786 (N_29786,N_28346,N_28098);
xnor U29787 (N_29787,N_28642,N_28801);
xnor U29788 (N_29788,N_28195,N_28571);
nand U29789 (N_29789,N_28483,N_28781);
xor U29790 (N_29790,N_28992,N_28399);
nor U29791 (N_29791,N_28567,N_28911);
or U29792 (N_29792,N_28024,N_28619);
xnor U29793 (N_29793,N_28435,N_28320);
nand U29794 (N_29794,N_28575,N_28285);
xnor U29795 (N_29795,N_28802,N_28752);
and U29796 (N_29796,N_28485,N_28254);
nor U29797 (N_29797,N_28070,N_28579);
nor U29798 (N_29798,N_28828,N_28458);
or U29799 (N_29799,N_28233,N_28282);
nor U29800 (N_29800,N_28690,N_28641);
xor U29801 (N_29801,N_28151,N_28076);
and U29802 (N_29802,N_28803,N_28549);
xor U29803 (N_29803,N_28529,N_28227);
or U29804 (N_29804,N_28652,N_28554);
nor U29805 (N_29805,N_28250,N_28284);
nand U29806 (N_29806,N_28205,N_28139);
xnor U29807 (N_29807,N_28804,N_28101);
nand U29808 (N_29808,N_28195,N_28938);
nand U29809 (N_29809,N_28050,N_28992);
nor U29810 (N_29810,N_28373,N_28826);
nand U29811 (N_29811,N_28630,N_28328);
xor U29812 (N_29812,N_28428,N_28963);
or U29813 (N_29813,N_28834,N_28055);
nor U29814 (N_29814,N_28015,N_28507);
xnor U29815 (N_29815,N_28175,N_28714);
or U29816 (N_29816,N_28202,N_28978);
and U29817 (N_29817,N_28958,N_28910);
nand U29818 (N_29818,N_28698,N_28074);
and U29819 (N_29819,N_28997,N_28198);
xnor U29820 (N_29820,N_28590,N_28106);
nand U29821 (N_29821,N_28551,N_28995);
and U29822 (N_29822,N_28657,N_28636);
nor U29823 (N_29823,N_28613,N_28633);
xnor U29824 (N_29824,N_28134,N_28487);
nor U29825 (N_29825,N_28990,N_28842);
nand U29826 (N_29826,N_28939,N_28620);
nor U29827 (N_29827,N_28764,N_28050);
or U29828 (N_29828,N_28226,N_28214);
xnor U29829 (N_29829,N_28721,N_28545);
nand U29830 (N_29830,N_28444,N_28728);
nor U29831 (N_29831,N_28053,N_28493);
and U29832 (N_29832,N_28312,N_28086);
nor U29833 (N_29833,N_28182,N_28017);
nand U29834 (N_29834,N_28849,N_28491);
nand U29835 (N_29835,N_28743,N_28470);
and U29836 (N_29836,N_28004,N_28108);
nand U29837 (N_29837,N_28687,N_28152);
xnor U29838 (N_29838,N_28288,N_28584);
or U29839 (N_29839,N_28019,N_28002);
xnor U29840 (N_29840,N_28442,N_28734);
and U29841 (N_29841,N_28570,N_28166);
or U29842 (N_29842,N_28069,N_28301);
nor U29843 (N_29843,N_28950,N_28394);
and U29844 (N_29844,N_28328,N_28675);
nand U29845 (N_29845,N_28866,N_28054);
nor U29846 (N_29846,N_28484,N_28769);
and U29847 (N_29847,N_28175,N_28036);
xnor U29848 (N_29848,N_28135,N_28130);
nor U29849 (N_29849,N_28827,N_28952);
xnor U29850 (N_29850,N_28580,N_28939);
xor U29851 (N_29851,N_28722,N_28655);
and U29852 (N_29852,N_28487,N_28207);
or U29853 (N_29853,N_28887,N_28648);
nand U29854 (N_29854,N_28672,N_28512);
nand U29855 (N_29855,N_28936,N_28985);
nor U29856 (N_29856,N_28507,N_28464);
and U29857 (N_29857,N_28471,N_28774);
or U29858 (N_29858,N_28196,N_28011);
xnor U29859 (N_29859,N_28390,N_28247);
and U29860 (N_29860,N_28258,N_28462);
and U29861 (N_29861,N_28343,N_28816);
xnor U29862 (N_29862,N_28467,N_28805);
nand U29863 (N_29863,N_28158,N_28922);
nand U29864 (N_29864,N_28397,N_28289);
and U29865 (N_29865,N_28688,N_28091);
xnor U29866 (N_29866,N_28512,N_28059);
xor U29867 (N_29867,N_28001,N_28977);
nand U29868 (N_29868,N_28199,N_28589);
nor U29869 (N_29869,N_28733,N_28465);
or U29870 (N_29870,N_28261,N_28704);
nand U29871 (N_29871,N_28255,N_28607);
nand U29872 (N_29872,N_28446,N_28913);
nor U29873 (N_29873,N_28860,N_28964);
nor U29874 (N_29874,N_28748,N_28580);
or U29875 (N_29875,N_28195,N_28587);
or U29876 (N_29876,N_28663,N_28596);
nand U29877 (N_29877,N_28181,N_28241);
or U29878 (N_29878,N_28948,N_28616);
or U29879 (N_29879,N_28035,N_28212);
nor U29880 (N_29880,N_28608,N_28863);
or U29881 (N_29881,N_28000,N_28399);
and U29882 (N_29882,N_28839,N_28362);
xor U29883 (N_29883,N_28184,N_28371);
or U29884 (N_29884,N_28757,N_28524);
and U29885 (N_29885,N_28962,N_28739);
xor U29886 (N_29886,N_28047,N_28181);
nor U29887 (N_29887,N_28752,N_28268);
or U29888 (N_29888,N_28836,N_28589);
nor U29889 (N_29889,N_28445,N_28221);
or U29890 (N_29890,N_28522,N_28062);
nor U29891 (N_29891,N_28026,N_28318);
nor U29892 (N_29892,N_28760,N_28982);
nor U29893 (N_29893,N_28277,N_28241);
nand U29894 (N_29894,N_28678,N_28863);
or U29895 (N_29895,N_28952,N_28157);
nor U29896 (N_29896,N_28766,N_28921);
and U29897 (N_29897,N_28371,N_28558);
or U29898 (N_29898,N_28580,N_28856);
or U29899 (N_29899,N_28138,N_28992);
nor U29900 (N_29900,N_28247,N_28118);
nor U29901 (N_29901,N_28619,N_28348);
nor U29902 (N_29902,N_28873,N_28247);
nand U29903 (N_29903,N_28048,N_28023);
nand U29904 (N_29904,N_28984,N_28074);
nor U29905 (N_29905,N_28560,N_28697);
nor U29906 (N_29906,N_28324,N_28979);
and U29907 (N_29907,N_28592,N_28929);
nor U29908 (N_29908,N_28946,N_28972);
and U29909 (N_29909,N_28057,N_28460);
xnor U29910 (N_29910,N_28684,N_28483);
nor U29911 (N_29911,N_28212,N_28643);
nor U29912 (N_29912,N_28566,N_28435);
xor U29913 (N_29913,N_28603,N_28717);
and U29914 (N_29914,N_28314,N_28107);
and U29915 (N_29915,N_28905,N_28566);
and U29916 (N_29916,N_28663,N_28579);
and U29917 (N_29917,N_28396,N_28757);
or U29918 (N_29918,N_28575,N_28717);
nand U29919 (N_29919,N_28858,N_28621);
and U29920 (N_29920,N_28876,N_28613);
and U29921 (N_29921,N_28931,N_28836);
xnor U29922 (N_29922,N_28994,N_28508);
nand U29923 (N_29923,N_28450,N_28179);
nor U29924 (N_29924,N_28113,N_28268);
xor U29925 (N_29925,N_28088,N_28464);
nand U29926 (N_29926,N_28949,N_28485);
nand U29927 (N_29927,N_28944,N_28655);
nand U29928 (N_29928,N_28983,N_28526);
xnor U29929 (N_29929,N_28076,N_28475);
or U29930 (N_29930,N_28768,N_28649);
nand U29931 (N_29931,N_28989,N_28091);
xor U29932 (N_29932,N_28038,N_28544);
or U29933 (N_29933,N_28109,N_28199);
and U29934 (N_29934,N_28543,N_28161);
nor U29935 (N_29935,N_28796,N_28861);
and U29936 (N_29936,N_28351,N_28750);
or U29937 (N_29937,N_28016,N_28349);
xor U29938 (N_29938,N_28655,N_28219);
xor U29939 (N_29939,N_28713,N_28097);
or U29940 (N_29940,N_28396,N_28719);
or U29941 (N_29941,N_28784,N_28152);
nor U29942 (N_29942,N_28680,N_28046);
or U29943 (N_29943,N_28022,N_28125);
nor U29944 (N_29944,N_28799,N_28949);
nor U29945 (N_29945,N_28717,N_28196);
xnor U29946 (N_29946,N_28739,N_28945);
or U29947 (N_29947,N_28902,N_28686);
nand U29948 (N_29948,N_28637,N_28129);
and U29949 (N_29949,N_28500,N_28663);
nand U29950 (N_29950,N_28013,N_28600);
xnor U29951 (N_29951,N_28185,N_28620);
nor U29952 (N_29952,N_28372,N_28949);
xor U29953 (N_29953,N_28754,N_28410);
nand U29954 (N_29954,N_28633,N_28865);
and U29955 (N_29955,N_28952,N_28019);
xnor U29956 (N_29956,N_28382,N_28544);
nand U29957 (N_29957,N_28921,N_28964);
xor U29958 (N_29958,N_28835,N_28989);
and U29959 (N_29959,N_28823,N_28757);
and U29960 (N_29960,N_28812,N_28449);
xnor U29961 (N_29961,N_28602,N_28428);
xor U29962 (N_29962,N_28799,N_28143);
xor U29963 (N_29963,N_28684,N_28184);
or U29964 (N_29964,N_28654,N_28936);
or U29965 (N_29965,N_28253,N_28759);
nand U29966 (N_29966,N_28116,N_28724);
or U29967 (N_29967,N_28727,N_28556);
and U29968 (N_29968,N_28108,N_28663);
and U29969 (N_29969,N_28349,N_28552);
and U29970 (N_29970,N_28303,N_28211);
or U29971 (N_29971,N_28399,N_28406);
xnor U29972 (N_29972,N_28036,N_28736);
or U29973 (N_29973,N_28081,N_28085);
nor U29974 (N_29974,N_28265,N_28790);
or U29975 (N_29975,N_28478,N_28394);
nor U29976 (N_29976,N_28367,N_28341);
or U29977 (N_29977,N_28079,N_28781);
or U29978 (N_29978,N_28682,N_28359);
or U29979 (N_29979,N_28580,N_28647);
or U29980 (N_29980,N_28340,N_28357);
or U29981 (N_29981,N_28388,N_28577);
nor U29982 (N_29982,N_28023,N_28807);
xnor U29983 (N_29983,N_28549,N_28458);
and U29984 (N_29984,N_28626,N_28356);
nor U29985 (N_29985,N_28975,N_28183);
or U29986 (N_29986,N_28932,N_28644);
xor U29987 (N_29987,N_28900,N_28574);
or U29988 (N_29988,N_28078,N_28681);
nand U29989 (N_29989,N_28751,N_28865);
nor U29990 (N_29990,N_28378,N_28815);
xor U29991 (N_29991,N_28647,N_28361);
or U29992 (N_29992,N_28591,N_28020);
or U29993 (N_29993,N_28240,N_28788);
and U29994 (N_29994,N_28676,N_28151);
nor U29995 (N_29995,N_28294,N_28337);
nand U29996 (N_29996,N_28160,N_28828);
nand U29997 (N_29997,N_28525,N_28852);
nand U29998 (N_29998,N_28963,N_28880);
nor U29999 (N_29999,N_28215,N_28996);
and U30000 (N_30000,N_29778,N_29724);
xor U30001 (N_30001,N_29087,N_29994);
xnor U30002 (N_30002,N_29225,N_29424);
xor U30003 (N_30003,N_29849,N_29137);
nand U30004 (N_30004,N_29649,N_29246);
nand U30005 (N_30005,N_29310,N_29083);
or U30006 (N_30006,N_29272,N_29103);
and U30007 (N_30007,N_29909,N_29675);
and U30008 (N_30008,N_29925,N_29893);
and U30009 (N_30009,N_29253,N_29062);
nor U30010 (N_30010,N_29433,N_29385);
or U30011 (N_30011,N_29088,N_29125);
nand U30012 (N_30012,N_29284,N_29290);
nand U30013 (N_30013,N_29219,N_29606);
nor U30014 (N_30014,N_29034,N_29511);
xnor U30015 (N_30015,N_29391,N_29589);
xnor U30016 (N_30016,N_29816,N_29817);
nand U30017 (N_30017,N_29264,N_29944);
nand U30018 (N_30018,N_29677,N_29612);
nand U30019 (N_30019,N_29962,N_29400);
or U30020 (N_30020,N_29469,N_29767);
nor U30021 (N_30021,N_29099,N_29494);
nor U30022 (N_30022,N_29930,N_29269);
nand U30023 (N_30023,N_29401,N_29493);
and U30024 (N_30024,N_29529,N_29305);
nand U30025 (N_30025,N_29259,N_29879);
nor U30026 (N_30026,N_29690,N_29389);
and U30027 (N_30027,N_29108,N_29254);
or U30028 (N_30028,N_29781,N_29757);
and U30029 (N_30029,N_29093,N_29460);
nand U30030 (N_30030,N_29251,N_29159);
nor U30031 (N_30031,N_29474,N_29814);
or U30032 (N_30032,N_29797,N_29117);
xor U30033 (N_30033,N_29359,N_29411);
nor U30034 (N_30034,N_29111,N_29971);
xor U30035 (N_30035,N_29704,N_29322);
xnor U30036 (N_30036,N_29847,N_29840);
and U30037 (N_30037,N_29277,N_29209);
xor U30038 (N_30038,N_29397,N_29100);
nor U30039 (N_30039,N_29366,N_29697);
nand U30040 (N_30040,N_29886,N_29967);
nand U30041 (N_30041,N_29887,N_29488);
or U30042 (N_30042,N_29454,N_29740);
nand U30043 (N_30043,N_29946,N_29725);
xnor U30044 (N_30044,N_29819,N_29321);
xor U30045 (N_30045,N_29075,N_29216);
or U30046 (N_30046,N_29676,N_29278);
and U30047 (N_30047,N_29168,N_29098);
nand U30048 (N_30048,N_29863,N_29080);
and U30049 (N_30049,N_29593,N_29170);
xnor U30050 (N_30050,N_29453,N_29599);
xor U30051 (N_30051,N_29796,N_29794);
nand U30052 (N_30052,N_29459,N_29245);
or U30053 (N_30053,N_29714,N_29053);
or U30054 (N_30054,N_29989,N_29236);
nor U30055 (N_30055,N_29215,N_29515);
xor U30056 (N_30056,N_29086,N_29996);
nand U30057 (N_30057,N_29294,N_29597);
nand U30058 (N_30058,N_29727,N_29659);
or U30059 (N_30059,N_29622,N_29779);
nor U30060 (N_30060,N_29519,N_29713);
or U30061 (N_30061,N_29067,N_29340);
nand U30062 (N_30062,N_29949,N_29233);
and U30063 (N_30063,N_29422,N_29073);
nor U30064 (N_30064,N_29789,N_29506);
and U30065 (N_30065,N_29437,N_29534);
nor U30066 (N_30066,N_29785,N_29427);
nand U30067 (N_30067,N_29995,N_29641);
nor U30068 (N_30068,N_29326,N_29113);
nor U30069 (N_30069,N_29364,N_29047);
xor U30070 (N_30070,N_29404,N_29694);
nor U30071 (N_30071,N_29361,N_29350);
or U30072 (N_30072,N_29749,N_29820);
nor U30073 (N_30073,N_29861,N_29221);
xnor U30074 (N_30074,N_29162,N_29402);
nor U30075 (N_30075,N_29540,N_29271);
and U30076 (N_30076,N_29716,N_29191);
xnor U30077 (N_30077,N_29561,N_29434);
and U30078 (N_30078,N_29743,N_29299);
nand U30079 (N_30079,N_29395,N_29337);
nor U30080 (N_30080,N_29639,N_29920);
nor U30081 (N_30081,N_29268,N_29393);
xnor U30082 (N_30082,N_29405,N_29806);
nand U30083 (N_30083,N_29478,N_29430);
nand U30084 (N_30084,N_29369,N_29428);
and U30085 (N_30085,N_29832,N_29448);
nor U30086 (N_30086,N_29429,N_29983);
nor U30087 (N_30087,N_29963,N_29208);
or U30088 (N_30088,N_29683,N_29482);
xor U30089 (N_30089,N_29856,N_29764);
nand U30090 (N_30090,N_29040,N_29241);
and U30091 (N_30091,N_29839,N_29009);
nand U30092 (N_30092,N_29383,N_29061);
nor U30093 (N_30093,N_29239,N_29423);
or U30094 (N_30094,N_29346,N_29250);
nand U30095 (N_30095,N_29917,N_29458);
and U30096 (N_30096,N_29986,N_29877);
nand U30097 (N_30097,N_29687,N_29288);
and U30098 (N_30098,N_29588,N_29844);
nor U30099 (N_30099,N_29370,N_29421);
nor U30100 (N_30100,N_29557,N_29384);
nor U30101 (N_30101,N_29595,N_29889);
xor U30102 (N_30102,N_29523,N_29637);
nor U30103 (N_30103,N_29633,N_29503);
nand U30104 (N_30104,N_29499,N_29664);
xor U30105 (N_30105,N_29997,N_29498);
and U30106 (N_30106,N_29267,N_29763);
nor U30107 (N_30107,N_29938,N_29851);
nor U30108 (N_30108,N_29896,N_29858);
and U30109 (N_30109,N_29201,N_29541);
nor U30110 (N_30110,N_29138,N_29901);
nand U30111 (N_30111,N_29802,N_29948);
nand U30112 (N_30112,N_29505,N_29578);
nand U30113 (N_30113,N_29336,N_29712);
or U30114 (N_30114,N_29536,N_29332);
nor U30115 (N_30115,N_29991,N_29771);
nor U30116 (N_30116,N_29569,N_29375);
xor U30117 (N_30117,N_29487,N_29984);
nor U30118 (N_30118,N_29450,N_29471);
or U30119 (N_30119,N_29243,N_29584);
nor U30120 (N_30120,N_29609,N_29618);
and U30121 (N_30121,N_29701,N_29335);
and U30122 (N_30122,N_29413,N_29957);
and U30123 (N_30123,N_29501,N_29163);
or U30124 (N_30124,N_29234,N_29377);
or U30125 (N_30125,N_29952,N_29547);
xnor U30126 (N_30126,N_29528,N_29263);
nand U30127 (N_30127,N_29635,N_29741);
nand U30128 (N_30128,N_29992,N_29733);
nand U30129 (N_30129,N_29753,N_29049);
or U30130 (N_30130,N_29857,N_29703);
or U30131 (N_30131,N_29171,N_29555);
nand U30132 (N_30132,N_29583,N_29031);
and U30133 (N_30133,N_29046,N_29530);
nor U30134 (N_30134,N_29248,N_29455);
or U30135 (N_30135,N_29329,N_29640);
nand U30136 (N_30136,N_29830,N_29442);
xor U30137 (N_30137,N_29751,N_29197);
and U30138 (N_30138,N_29222,N_29975);
nand U30139 (N_30139,N_29287,N_29959);
xor U30140 (N_30140,N_29072,N_29484);
nor U30141 (N_30141,N_29898,N_29688);
or U30142 (N_30142,N_29860,N_29682);
nor U30143 (N_30143,N_29205,N_29419);
xor U30144 (N_30144,N_29089,N_29656);
and U30145 (N_30145,N_29123,N_29153);
nor U30146 (N_30146,N_29064,N_29709);
or U30147 (N_30147,N_29672,N_29476);
nand U30148 (N_30148,N_29472,N_29373);
nor U30149 (N_30149,N_29642,N_29367);
xor U30150 (N_30150,N_29485,N_29852);
or U30151 (N_30151,N_29490,N_29821);
and U30152 (N_30152,N_29029,N_29550);
nand U30153 (N_30153,N_29296,N_29576);
or U30154 (N_30154,N_29002,N_29591);
nor U30155 (N_30155,N_29556,N_29431);
or U30156 (N_30156,N_29070,N_29926);
xnor U30157 (N_30157,N_29812,N_29152);
and U30158 (N_30158,N_29325,N_29463);
and U30159 (N_30159,N_29365,N_29068);
or U30160 (N_30160,N_29516,N_29653);
xor U30161 (N_30161,N_29360,N_29614);
and U30162 (N_30162,N_29766,N_29242);
nor U30163 (N_30163,N_29846,N_29607);
nand U30164 (N_30164,N_29227,N_29939);
or U30165 (N_30165,N_29600,N_29174);
nor U30166 (N_30166,N_29303,N_29041);
nand U30167 (N_30167,N_29900,N_29065);
or U30168 (N_30168,N_29924,N_29140);
nand U30169 (N_30169,N_29217,N_29931);
nand U30170 (N_30170,N_29543,N_29120);
or U30171 (N_30171,N_29803,N_29235);
nand U30172 (N_30172,N_29643,N_29730);
and U30173 (N_30173,N_29207,N_29085);
nand U30174 (N_30174,N_29573,N_29097);
nand U30175 (N_30175,N_29035,N_29507);
or U30176 (N_30176,N_29956,N_29565);
nand U30177 (N_30177,N_29107,N_29890);
and U30178 (N_30178,N_29416,N_29392);
xnor U30179 (N_30179,N_29842,N_29489);
and U30180 (N_30180,N_29344,N_29624);
nand U30181 (N_30181,N_29323,N_29621);
nand U30182 (N_30182,N_29927,N_29590);
or U30183 (N_30183,N_29461,N_29412);
nand U30184 (N_30184,N_29567,N_29409);
or U30185 (N_30185,N_29969,N_29603);
nor U30186 (N_30186,N_29330,N_29300);
nand U30187 (N_30187,N_29908,N_29261);
xnor U30188 (N_30188,N_29016,N_29403);
or U30189 (N_30189,N_29020,N_29980);
or U30190 (N_30190,N_29435,N_29647);
nor U30191 (N_30191,N_29045,N_29870);
nor U30192 (N_30192,N_29809,N_29723);
xor U30193 (N_30193,N_29203,N_29492);
nand U30194 (N_30194,N_29457,N_29014);
or U30195 (N_30195,N_29738,N_29554);
and U30196 (N_30196,N_29180,N_29148);
nand U30197 (N_30197,N_29575,N_29824);
and U30198 (N_30198,N_29028,N_29645);
and U30199 (N_30199,N_29151,N_29306);
xnor U30200 (N_30200,N_29545,N_29204);
xnor U30201 (N_30201,N_29169,N_29304);
nor U30202 (N_30202,N_29032,N_29702);
nand U30203 (N_30203,N_29388,N_29513);
or U30204 (N_30204,N_29281,N_29445);
or U30205 (N_30205,N_29313,N_29116);
nor U30206 (N_30206,N_29696,N_29297);
xor U30207 (N_30207,N_29732,N_29628);
and U30208 (N_30208,N_29291,N_29951);
or U30209 (N_30209,N_29240,N_29342);
nor U30210 (N_30210,N_29982,N_29255);
nand U30211 (N_30211,N_29610,N_29620);
nand U30212 (N_30212,N_29737,N_29906);
nor U30213 (N_30213,N_29750,N_29880);
nor U30214 (N_30214,N_29426,N_29521);
xor U30215 (N_30215,N_29021,N_29721);
nand U30216 (N_30216,N_29532,N_29178);
nand U30217 (N_30217,N_29700,N_29990);
xnor U30218 (N_30218,N_29408,N_29232);
nor U30219 (N_30219,N_29985,N_29841);
nand U30220 (N_30220,N_29497,N_29695);
and U30221 (N_30221,N_29155,N_29466);
xnor U30222 (N_30222,N_29976,N_29387);
nor U30223 (N_30223,N_29055,N_29648);
nand U30224 (N_30224,N_29773,N_29671);
and U30225 (N_30225,N_29228,N_29605);
xor U30226 (N_30226,N_29551,N_29285);
nand U30227 (N_30227,N_29810,N_29950);
nor U30228 (N_30228,N_29376,N_29167);
nor U30229 (N_30229,N_29128,N_29292);
nor U30230 (N_30230,N_29914,N_29586);
or U30231 (N_30231,N_29467,N_29566);
or U30232 (N_30232,N_29793,N_29772);
or U30233 (N_30233,N_29465,N_29092);
or U30234 (N_30234,N_29142,N_29827);
or U30235 (N_30235,N_29184,N_29504);
or U30236 (N_30236,N_29439,N_29007);
and U30237 (N_30237,N_29972,N_29934);
nor U30238 (N_30238,N_29722,N_29024);
nand U30239 (N_30239,N_29008,N_29182);
xor U30240 (N_30240,N_29496,N_29030);
xnor U30241 (N_30241,N_29734,N_29616);
nor U30242 (N_30242,N_29932,N_29850);
or U30243 (N_30243,N_29598,N_29273);
or U30244 (N_30244,N_29407,N_29899);
xnor U30245 (N_30245,N_29759,N_29728);
or U30246 (N_30246,N_29681,N_29374);
and U30247 (N_30247,N_29845,N_29059);
nor U30248 (N_30248,N_29394,N_29302);
or U30249 (N_30249,N_29692,N_29865);
xor U30250 (N_30250,N_29577,N_29755);
nand U30251 (N_30251,N_29940,N_29015);
xor U30252 (N_30252,N_29449,N_29632);
xor U30253 (N_30253,N_29145,N_29592);
nand U30254 (N_30254,N_29158,N_29351);
or U30255 (N_30255,N_29106,N_29022);
and U30256 (N_30256,N_29788,N_29762);
and U30257 (N_30257,N_29615,N_29480);
xnor U30258 (N_30258,N_29134,N_29126);
nand U30259 (N_30259,N_29136,N_29166);
nor U30260 (N_30260,N_29813,N_29071);
or U30261 (N_30261,N_29003,N_29043);
and U30262 (N_30262,N_29790,N_29838);
nand U30263 (N_30263,N_29756,N_29684);
nor U30264 (N_30264,N_29500,N_29579);
and U30265 (N_30265,N_29758,N_29110);
and U30266 (N_30266,N_29260,N_29320);
nand U30267 (N_30267,N_29122,N_29244);
and U30268 (N_30268,N_29052,N_29804);
xnor U30269 (N_30269,N_29538,N_29308);
or U30270 (N_30270,N_29188,N_29262);
nand U30271 (N_30271,N_29869,N_29999);
nor U30272 (N_30272,N_29746,N_29025);
or U30273 (N_30273,N_29096,N_29101);
nand U30274 (N_30274,N_29175,N_29345);
nor U30275 (N_30275,N_29440,N_29356);
nor U30276 (N_30276,N_29443,N_29878);
nor U30277 (N_30277,N_29033,N_29658);
nand U30278 (N_30278,N_29023,N_29587);
and U30279 (N_30279,N_29776,N_29911);
or U30280 (N_30280,N_29711,N_29456);
xnor U30281 (N_30281,N_29678,N_29707);
xnor U30282 (N_30282,N_29109,N_29141);
nor U30283 (N_30283,N_29314,N_29784);
and U30284 (N_30284,N_29646,N_29552);
and U30285 (N_30285,N_29754,N_29210);
nand U30286 (N_30286,N_29775,N_29509);
and U30287 (N_30287,N_29945,N_29298);
xor U30288 (N_30288,N_29194,N_29105);
or U30289 (N_30289,N_29828,N_29131);
or U30290 (N_30290,N_29179,N_29432);
or U30291 (N_30291,N_29143,N_29144);
nand U30292 (N_30292,N_29947,N_29673);
nand U30293 (N_30293,N_29582,N_29660);
or U30294 (N_30294,N_29293,N_29638);
nand U30295 (N_30295,N_29256,N_29922);
nor U30296 (N_30296,N_29871,N_29237);
nand U30297 (N_30297,N_29823,N_29317);
or U30298 (N_30298,N_29470,N_29399);
and U30299 (N_30299,N_29328,N_29602);
or U30300 (N_30300,N_29563,N_29661);
or U30301 (N_30301,N_29617,N_29249);
or U30302 (N_30302,N_29380,N_29124);
and U30303 (N_30303,N_29928,N_29627);
or U30304 (N_30304,N_29936,N_29218);
nand U30305 (N_30305,N_29955,N_29079);
xnor U30306 (N_30306,N_29973,N_29051);
or U30307 (N_30307,N_29252,N_29462);
or U30308 (N_30308,N_29885,N_29798);
and U30309 (N_30309,N_29542,N_29895);
nor U30310 (N_30310,N_29118,N_29836);
or U30311 (N_30311,N_29444,N_29199);
xor U30312 (N_30312,N_29524,N_29910);
and U30313 (N_30313,N_29919,N_29679);
or U30314 (N_30314,N_29343,N_29280);
and U30315 (N_30315,N_29729,N_29348);
xor U30316 (N_30316,N_29663,N_29368);
or U30317 (N_30317,N_29069,N_29902);
or U30318 (N_30318,N_29652,N_29146);
nor U30319 (N_30319,N_29058,N_29791);
or U30320 (N_30320,N_29196,N_29941);
xnor U30321 (N_30321,N_29974,N_29060);
nand U30322 (N_30322,N_29200,N_29888);
and U30323 (N_30323,N_29834,N_29198);
or U30324 (N_30324,N_29859,N_29913);
nor U30325 (N_30325,N_29825,N_29960);
nand U30326 (N_30326,N_29341,N_29266);
xnor U30327 (N_30327,N_29231,N_29881);
nor U30328 (N_30328,N_29691,N_29386);
nand U30329 (N_30329,N_29156,N_29708);
or U30330 (N_30330,N_29961,N_29082);
or U30331 (N_30331,N_29868,N_29044);
xor U30332 (N_30332,N_29212,N_29274);
nor U30333 (N_30333,N_29826,N_29347);
nand U30334 (N_30334,N_29537,N_29334);
nand U30335 (N_30335,N_29327,N_29993);
nand U30336 (N_30336,N_29855,N_29415);
nor U30337 (N_30337,N_29815,N_29650);
and U30338 (N_30338,N_29417,N_29634);
or U30339 (N_30339,N_29742,N_29414);
xor U30340 (N_30340,N_29301,N_29119);
and U30341 (N_30341,N_29017,N_29731);
nand U30342 (N_30342,N_29258,N_29929);
nand U30343 (N_30343,N_29211,N_29333);
or U30344 (N_30344,N_29001,N_29319);
xnor U30345 (N_30345,N_29866,N_29226);
or U30346 (N_30346,N_29363,N_29745);
xnor U30347 (N_30347,N_29981,N_29522);
nand U30348 (N_30348,N_29874,N_29229);
xor U30349 (N_30349,N_29872,N_29670);
xor U30350 (N_30350,N_29873,N_29176);
or U30351 (N_30351,N_29943,N_29279);
nand U30352 (N_30352,N_29854,N_29186);
xnor U30353 (N_30353,N_29693,N_29090);
and U30354 (N_30354,N_29553,N_29800);
or U30355 (N_30355,N_29420,N_29718);
nand U30356 (N_30356,N_29935,N_29719);
xor U30357 (N_30357,N_29165,N_29937);
or U30358 (N_30358,N_29121,N_29636);
xor U30359 (N_30359,N_29657,N_29183);
nand U30360 (N_30360,N_29782,N_29735);
xnor U30361 (N_30361,N_29894,N_29970);
nor U30362 (N_30362,N_29436,N_29526);
xor U30363 (N_30363,N_29953,N_29012);
or U30364 (N_30364,N_29883,N_29904);
and U30365 (N_30365,N_29195,N_29717);
nor U30366 (N_30366,N_29998,N_29942);
or U30367 (N_30367,N_29486,N_29964);
or U30368 (N_30368,N_29903,N_29132);
nor U30369 (N_30369,N_29843,N_29230);
nor U30370 (N_30370,N_29010,N_29127);
nand U30371 (N_30371,N_29094,N_29626);
nor U30372 (N_30372,N_29864,N_29081);
nand U30373 (N_30373,N_29568,N_29475);
or U30374 (N_30374,N_29315,N_29187);
nor U30375 (N_30375,N_29921,N_29780);
or U30376 (N_30376,N_29644,N_29238);
and U30377 (N_30377,N_29958,N_29477);
or U30378 (N_30378,N_29837,N_29418);
and U30379 (N_30379,N_29818,N_29202);
and U30380 (N_30380,N_29558,N_29206);
and U30381 (N_30381,N_29311,N_29792);
nor U30382 (N_30382,N_29744,N_29004);
nor U30383 (N_30383,N_29669,N_29307);
or U30384 (N_30384,N_29220,N_29161);
nand U30385 (N_30385,N_29479,N_29048);
xnor U30386 (N_30386,N_29581,N_29452);
nor U30387 (N_30387,N_29665,N_29446);
or U30388 (N_30388,N_29923,N_29706);
or U30389 (N_30389,N_29382,N_29608);
nor U30390 (N_30390,N_29979,N_29037);
nand U30391 (N_30391,N_29102,N_29654);
or U30392 (N_30392,N_29801,N_29698);
or U30393 (N_30393,N_29527,N_29104);
xor U30394 (N_30394,N_29726,N_29807);
nor U30395 (N_30395,N_29352,N_29130);
or U30396 (N_30396,N_29160,N_29822);
or U30397 (N_30397,N_29316,N_29077);
or U30398 (N_30398,N_29508,N_29966);
nor U30399 (N_30399,N_29564,N_29761);
nand U30400 (N_30400,N_29867,N_29036);
nor U30401 (N_30401,N_29685,N_29056);
xor U30402 (N_30402,N_29224,N_29585);
or U30403 (N_30403,N_29177,N_29154);
or U30404 (N_30404,N_29667,N_29084);
xnor U30405 (N_30405,N_29286,N_29774);
nor U30406 (N_30406,N_29912,N_29276);
nand U30407 (N_30407,N_29787,N_29398);
nor U30408 (N_30408,N_29447,N_29018);
nor U30409 (N_30409,N_29133,N_29027);
nand U30410 (N_30410,N_29918,N_29172);
or U30411 (N_30411,N_29662,N_29338);
nor U30412 (N_30412,N_29406,N_29987);
and U30413 (N_30413,N_29596,N_29265);
nand U30414 (N_30414,N_29808,N_29076);
and U30415 (N_30415,N_29915,N_29531);
nand U30416 (N_30416,N_29699,N_29190);
or U30417 (N_30417,N_29006,N_29517);
nor U30418 (N_30418,N_29349,N_29533);
nor U30419 (N_30419,N_29378,N_29038);
xor U30420 (N_30420,N_29988,N_29483);
nor U30421 (N_30421,N_29795,N_29559);
or U30422 (N_30422,N_29535,N_29760);
and U30423 (N_30423,N_29362,N_29026);
or U30424 (N_30424,N_29078,N_29495);
or U30425 (N_30425,N_29000,N_29897);
or U30426 (N_30426,N_29339,N_29135);
or U30427 (N_30427,N_29468,N_29147);
and U30428 (N_30428,N_29862,N_29115);
and U30429 (N_30429,N_29549,N_29655);
and U30430 (N_30430,N_29548,N_29525);
nand U30431 (N_30431,N_29765,N_29289);
xnor U30432 (N_30432,N_29481,N_29282);
or U30433 (N_30433,N_29625,N_29619);
nor U30434 (N_30434,N_29063,N_29112);
and U30435 (N_30435,N_29623,N_29114);
and U30436 (N_30436,N_29312,N_29129);
nand U30437 (N_30437,N_29371,N_29748);
or U30438 (N_30438,N_29213,N_29777);
or U30439 (N_30439,N_29630,N_29354);
and U30440 (N_30440,N_29013,N_29514);
nor U30441 (N_30441,N_29977,N_29283);
or U30442 (N_30442,N_29318,N_29933);
nor U30443 (N_30443,N_29150,N_29544);
nor U30444 (N_30444,N_29680,N_29629);
nand U30445 (N_30445,N_29054,N_29091);
nor U30446 (N_30446,N_29309,N_29066);
nor U30447 (N_30447,N_29876,N_29954);
or U30448 (N_30448,N_29752,N_29884);
xor U30449 (N_30449,N_29574,N_29425);
or U30450 (N_30450,N_29572,N_29185);
or U30451 (N_30451,N_29768,N_29686);
and U30452 (N_30452,N_29410,N_29848);
xnor U30453 (N_30453,N_29739,N_29057);
xor U30454 (N_30454,N_29358,N_29715);
nor U30455 (N_30455,N_29570,N_29441);
or U30456 (N_30456,N_29005,N_29042);
and U30457 (N_30457,N_29710,N_29562);
and U30458 (N_30458,N_29799,N_29512);
or U30459 (N_30459,N_29257,N_29668);
nand U30460 (N_30460,N_29074,N_29786);
or U30461 (N_30461,N_29580,N_29905);
and U30462 (N_30462,N_29631,N_29039);
nand U30463 (N_30463,N_29835,N_29811);
nor U30464 (N_30464,N_29892,N_29095);
and U30465 (N_30465,N_29571,N_29223);
nor U30466 (N_30466,N_29193,N_29747);
nor U30467 (N_30467,N_29907,N_29390);
nor U30468 (N_30468,N_29173,N_29502);
nand U30469 (N_30469,N_29968,N_29473);
nor U30470 (N_30470,N_29357,N_29396);
or U30471 (N_30471,N_29192,N_29666);
xnor U30472 (N_30472,N_29270,N_29783);
nand U30473 (N_30473,N_29978,N_29916);
nand U30474 (N_30474,N_29295,N_29247);
nor U30475 (N_30475,N_29601,N_29833);
or U30476 (N_30476,N_29189,N_29560);
nand U30477 (N_30477,N_29805,N_29736);
nor U30478 (N_30478,N_29769,N_29882);
and U30479 (N_30479,N_29451,N_29689);
and U30480 (N_30480,N_29875,N_29438);
or U30481 (N_30481,N_29604,N_29705);
nor U30482 (N_30482,N_29770,N_29149);
and U30483 (N_30483,N_29379,N_29720);
and U30484 (N_30484,N_29674,N_29831);
nand U30485 (N_30485,N_29353,N_29381);
or U30486 (N_30486,N_29520,N_29546);
nand U30487 (N_30487,N_29324,N_29181);
or U30488 (N_30488,N_29965,N_29518);
nand U30489 (N_30489,N_29611,N_29594);
or U30490 (N_30490,N_29853,N_29011);
nand U30491 (N_30491,N_29491,N_29891);
nand U30492 (N_30492,N_29355,N_29331);
nand U30493 (N_30493,N_29214,N_29275);
or U30494 (N_30494,N_29464,N_29539);
or U30495 (N_30495,N_29372,N_29157);
nor U30496 (N_30496,N_29019,N_29139);
xnor U30497 (N_30497,N_29510,N_29050);
or U30498 (N_30498,N_29164,N_29829);
xor U30499 (N_30499,N_29651,N_29613);
nor U30500 (N_30500,N_29938,N_29734);
nor U30501 (N_30501,N_29185,N_29661);
xor U30502 (N_30502,N_29385,N_29213);
nor U30503 (N_30503,N_29961,N_29049);
and U30504 (N_30504,N_29188,N_29040);
nor U30505 (N_30505,N_29475,N_29922);
and U30506 (N_30506,N_29950,N_29513);
nand U30507 (N_30507,N_29346,N_29932);
nor U30508 (N_30508,N_29879,N_29156);
xor U30509 (N_30509,N_29773,N_29242);
nand U30510 (N_30510,N_29785,N_29534);
nand U30511 (N_30511,N_29080,N_29004);
and U30512 (N_30512,N_29349,N_29298);
xnor U30513 (N_30513,N_29365,N_29059);
or U30514 (N_30514,N_29973,N_29114);
nand U30515 (N_30515,N_29052,N_29699);
or U30516 (N_30516,N_29953,N_29222);
or U30517 (N_30517,N_29221,N_29870);
xnor U30518 (N_30518,N_29243,N_29043);
and U30519 (N_30519,N_29368,N_29835);
or U30520 (N_30520,N_29580,N_29172);
nand U30521 (N_30521,N_29225,N_29625);
xor U30522 (N_30522,N_29188,N_29946);
nor U30523 (N_30523,N_29050,N_29955);
or U30524 (N_30524,N_29774,N_29897);
nand U30525 (N_30525,N_29027,N_29583);
xnor U30526 (N_30526,N_29364,N_29118);
nor U30527 (N_30527,N_29545,N_29161);
and U30528 (N_30528,N_29407,N_29731);
xnor U30529 (N_30529,N_29584,N_29625);
nor U30530 (N_30530,N_29604,N_29418);
xor U30531 (N_30531,N_29368,N_29396);
and U30532 (N_30532,N_29943,N_29289);
xor U30533 (N_30533,N_29405,N_29535);
nor U30534 (N_30534,N_29579,N_29237);
nand U30535 (N_30535,N_29493,N_29081);
or U30536 (N_30536,N_29532,N_29756);
or U30537 (N_30537,N_29092,N_29261);
nand U30538 (N_30538,N_29666,N_29019);
and U30539 (N_30539,N_29016,N_29896);
or U30540 (N_30540,N_29177,N_29174);
nand U30541 (N_30541,N_29397,N_29250);
xor U30542 (N_30542,N_29463,N_29944);
nor U30543 (N_30543,N_29750,N_29124);
nor U30544 (N_30544,N_29583,N_29936);
nand U30545 (N_30545,N_29462,N_29137);
xnor U30546 (N_30546,N_29085,N_29004);
and U30547 (N_30547,N_29171,N_29328);
nand U30548 (N_30548,N_29047,N_29419);
nand U30549 (N_30549,N_29751,N_29402);
nor U30550 (N_30550,N_29573,N_29020);
and U30551 (N_30551,N_29454,N_29448);
and U30552 (N_30552,N_29605,N_29371);
nand U30553 (N_30553,N_29113,N_29556);
nand U30554 (N_30554,N_29857,N_29534);
or U30555 (N_30555,N_29637,N_29173);
and U30556 (N_30556,N_29191,N_29241);
or U30557 (N_30557,N_29004,N_29670);
xor U30558 (N_30558,N_29923,N_29254);
xor U30559 (N_30559,N_29434,N_29433);
and U30560 (N_30560,N_29889,N_29877);
or U30561 (N_30561,N_29753,N_29294);
or U30562 (N_30562,N_29534,N_29423);
and U30563 (N_30563,N_29272,N_29160);
nor U30564 (N_30564,N_29151,N_29861);
and U30565 (N_30565,N_29656,N_29382);
nor U30566 (N_30566,N_29905,N_29872);
xnor U30567 (N_30567,N_29059,N_29199);
and U30568 (N_30568,N_29519,N_29412);
nand U30569 (N_30569,N_29811,N_29992);
nor U30570 (N_30570,N_29341,N_29957);
and U30571 (N_30571,N_29975,N_29579);
and U30572 (N_30572,N_29557,N_29222);
nor U30573 (N_30573,N_29444,N_29046);
nand U30574 (N_30574,N_29593,N_29990);
or U30575 (N_30575,N_29848,N_29849);
or U30576 (N_30576,N_29221,N_29183);
nor U30577 (N_30577,N_29548,N_29075);
or U30578 (N_30578,N_29832,N_29196);
or U30579 (N_30579,N_29344,N_29829);
xor U30580 (N_30580,N_29142,N_29759);
or U30581 (N_30581,N_29499,N_29365);
nor U30582 (N_30582,N_29132,N_29463);
or U30583 (N_30583,N_29711,N_29137);
and U30584 (N_30584,N_29132,N_29598);
or U30585 (N_30585,N_29116,N_29513);
nor U30586 (N_30586,N_29608,N_29663);
or U30587 (N_30587,N_29624,N_29398);
xor U30588 (N_30588,N_29563,N_29743);
and U30589 (N_30589,N_29430,N_29836);
and U30590 (N_30590,N_29756,N_29916);
nor U30591 (N_30591,N_29583,N_29062);
or U30592 (N_30592,N_29269,N_29020);
nor U30593 (N_30593,N_29782,N_29842);
xnor U30594 (N_30594,N_29463,N_29800);
or U30595 (N_30595,N_29076,N_29289);
or U30596 (N_30596,N_29579,N_29146);
nand U30597 (N_30597,N_29913,N_29007);
or U30598 (N_30598,N_29291,N_29689);
or U30599 (N_30599,N_29930,N_29560);
nand U30600 (N_30600,N_29727,N_29349);
and U30601 (N_30601,N_29425,N_29733);
nand U30602 (N_30602,N_29553,N_29081);
nand U30603 (N_30603,N_29110,N_29599);
nor U30604 (N_30604,N_29536,N_29893);
nand U30605 (N_30605,N_29254,N_29241);
or U30606 (N_30606,N_29955,N_29982);
xnor U30607 (N_30607,N_29324,N_29006);
nor U30608 (N_30608,N_29811,N_29729);
or U30609 (N_30609,N_29475,N_29594);
nor U30610 (N_30610,N_29606,N_29135);
nor U30611 (N_30611,N_29556,N_29622);
and U30612 (N_30612,N_29700,N_29429);
and U30613 (N_30613,N_29366,N_29216);
xor U30614 (N_30614,N_29170,N_29966);
nor U30615 (N_30615,N_29371,N_29514);
xor U30616 (N_30616,N_29257,N_29330);
or U30617 (N_30617,N_29155,N_29864);
nand U30618 (N_30618,N_29135,N_29604);
nand U30619 (N_30619,N_29539,N_29640);
xnor U30620 (N_30620,N_29255,N_29289);
nor U30621 (N_30621,N_29953,N_29864);
or U30622 (N_30622,N_29958,N_29497);
or U30623 (N_30623,N_29127,N_29519);
and U30624 (N_30624,N_29966,N_29770);
nor U30625 (N_30625,N_29579,N_29362);
nor U30626 (N_30626,N_29823,N_29393);
and U30627 (N_30627,N_29815,N_29786);
nor U30628 (N_30628,N_29155,N_29636);
xnor U30629 (N_30629,N_29412,N_29778);
and U30630 (N_30630,N_29196,N_29909);
nand U30631 (N_30631,N_29466,N_29205);
nand U30632 (N_30632,N_29294,N_29419);
xnor U30633 (N_30633,N_29686,N_29696);
nand U30634 (N_30634,N_29949,N_29904);
nor U30635 (N_30635,N_29320,N_29401);
xor U30636 (N_30636,N_29742,N_29085);
and U30637 (N_30637,N_29630,N_29785);
nor U30638 (N_30638,N_29290,N_29651);
and U30639 (N_30639,N_29685,N_29648);
and U30640 (N_30640,N_29564,N_29108);
nand U30641 (N_30641,N_29871,N_29591);
and U30642 (N_30642,N_29989,N_29959);
xnor U30643 (N_30643,N_29735,N_29825);
nor U30644 (N_30644,N_29955,N_29819);
or U30645 (N_30645,N_29828,N_29356);
xnor U30646 (N_30646,N_29324,N_29050);
nor U30647 (N_30647,N_29764,N_29512);
nor U30648 (N_30648,N_29275,N_29390);
nand U30649 (N_30649,N_29343,N_29479);
nor U30650 (N_30650,N_29561,N_29743);
xnor U30651 (N_30651,N_29968,N_29740);
and U30652 (N_30652,N_29190,N_29729);
nand U30653 (N_30653,N_29671,N_29215);
nor U30654 (N_30654,N_29429,N_29448);
xnor U30655 (N_30655,N_29541,N_29489);
and U30656 (N_30656,N_29986,N_29299);
nand U30657 (N_30657,N_29179,N_29834);
or U30658 (N_30658,N_29787,N_29813);
or U30659 (N_30659,N_29097,N_29583);
xor U30660 (N_30660,N_29715,N_29233);
nand U30661 (N_30661,N_29628,N_29416);
nor U30662 (N_30662,N_29815,N_29455);
xor U30663 (N_30663,N_29115,N_29889);
nand U30664 (N_30664,N_29955,N_29032);
nor U30665 (N_30665,N_29786,N_29211);
or U30666 (N_30666,N_29246,N_29826);
or U30667 (N_30667,N_29775,N_29556);
xor U30668 (N_30668,N_29203,N_29035);
or U30669 (N_30669,N_29148,N_29632);
xnor U30670 (N_30670,N_29704,N_29048);
or U30671 (N_30671,N_29176,N_29205);
and U30672 (N_30672,N_29307,N_29128);
or U30673 (N_30673,N_29616,N_29251);
or U30674 (N_30674,N_29292,N_29774);
nand U30675 (N_30675,N_29981,N_29075);
xor U30676 (N_30676,N_29468,N_29364);
nand U30677 (N_30677,N_29903,N_29375);
or U30678 (N_30678,N_29091,N_29537);
xor U30679 (N_30679,N_29886,N_29106);
or U30680 (N_30680,N_29795,N_29117);
nand U30681 (N_30681,N_29449,N_29868);
xor U30682 (N_30682,N_29403,N_29866);
xor U30683 (N_30683,N_29166,N_29114);
or U30684 (N_30684,N_29360,N_29093);
and U30685 (N_30685,N_29457,N_29709);
or U30686 (N_30686,N_29749,N_29552);
or U30687 (N_30687,N_29219,N_29491);
and U30688 (N_30688,N_29407,N_29796);
or U30689 (N_30689,N_29227,N_29716);
xnor U30690 (N_30690,N_29364,N_29401);
nor U30691 (N_30691,N_29417,N_29630);
or U30692 (N_30692,N_29402,N_29781);
nor U30693 (N_30693,N_29826,N_29451);
and U30694 (N_30694,N_29439,N_29817);
nand U30695 (N_30695,N_29866,N_29230);
nor U30696 (N_30696,N_29373,N_29388);
xor U30697 (N_30697,N_29395,N_29990);
or U30698 (N_30698,N_29627,N_29481);
nor U30699 (N_30699,N_29647,N_29808);
xor U30700 (N_30700,N_29972,N_29879);
xnor U30701 (N_30701,N_29989,N_29318);
or U30702 (N_30702,N_29824,N_29690);
nor U30703 (N_30703,N_29625,N_29400);
nand U30704 (N_30704,N_29268,N_29220);
nand U30705 (N_30705,N_29142,N_29435);
xor U30706 (N_30706,N_29920,N_29169);
or U30707 (N_30707,N_29404,N_29775);
nand U30708 (N_30708,N_29891,N_29285);
nand U30709 (N_30709,N_29200,N_29893);
nand U30710 (N_30710,N_29839,N_29795);
and U30711 (N_30711,N_29901,N_29251);
nor U30712 (N_30712,N_29824,N_29899);
nand U30713 (N_30713,N_29098,N_29441);
nor U30714 (N_30714,N_29769,N_29502);
and U30715 (N_30715,N_29418,N_29092);
nor U30716 (N_30716,N_29365,N_29482);
and U30717 (N_30717,N_29618,N_29239);
nor U30718 (N_30718,N_29793,N_29194);
and U30719 (N_30719,N_29002,N_29839);
nor U30720 (N_30720,N_29474,N_29209);
or U30721 (N_30721,N_29535,N_29318);
xnor U30722 (N_30722,N_29329,N_29069);
and U30723 (N_30723,N_29415,N_29576);
xor U30724 (N_30724,N_29969,N_29003);
or U30725 (N_30725,N_29184,N_29002);
or U30726 (N_30726,N_29729,N_29308);
and U30727 (N_30727,N_29495,N_29576);
xnor U30728 (N_30728,N_29708,N_29801);
nor U30729 (N_30729,N_29431,N_29913);
nor U30730 (N_30730,N_29589,N_29492);
and U30731 (N_30731,N_29094,N_29247);
nor U30732 (N_30732,N_29286,N_29815);
xnor U30733 (N_30733,N_29185,N_29213);
xor U30734 (N_30734,N_29163,N_29465);
nor U30735 (N_30735,N_29980,N_29022);
nand U30736 (N_30736,N_29509,N_29217);
nor U30737 (N_30737,N_29869,N_29718);
nand U30738 (N_30738,N_29991,N_29225);
or U30739 (N_30739,N_29883,N_29626);
nand U30740 (N_30740,N_29401,N_29095);
nand U30741 (N_30741,N_29980,N_29114);
nand U30742 (N_30742,N_29293,N_29893);
nor U30743 (N_30743,N_29339,N_29871);
nand U30744 (N_30744,N_29401,N_29188);
nand U30745 (N_30745,N_29146,N_29405);
and U30746 (N_30746,N_29201,N_29001);
and U30747 (N_30747,N_29422,N_29411);
and U30748 (N_30748,N_29550,N_29243);
or U30749 (N_30749,N_29462,N_29683);
xor U30750 (N_30750,N_29879,N_29053);
or U30751 (N_30751,N_29928,N_29669);
and U30752 (N_30752,N_29853,N_29789);
or U30753 (N_30753,N_29213,N_29378);
nand U30754 (N_30754,N_29878,N_29228);
and U30755 (N_30755,N_29169,N_29497);
or U30756 (N_30756,N_29060,N_29623);
or U30757 (N_30757,N_29555,N_29619);
and U30758 (N_30758,N_29316,N_29170);
xnor U30759 (N_30759,N_29574,N_29444);
xnor U30760 (N_30760,N_29963,N_29249);
nor U30761 (N_30761,N_29155,N_29390);
xnor U30762 (N_30762,N_29821,N_29353);
nor U30763 (N_30763,N_29352,N_29485);
and U30764 (N_30764,N_29828,N_29584);
nand U30765 (N_30765,N_29053,N_29456);
nor U30766 (N_30766,N_29193,N_29144);
nand U30767 (N_30767,N_29325,N_29104);
or U30768 (N_30768,N_29035,N_29851);
nor U30769 (N_30769,N_29350,N_29097);
and U30770 (N_30770,N_29280,N_29516);
nand U30771 (N_30771,N_29214,N_29499);
and U30772 (N_30772,N_29923,N_29632);
nor U30773 (N_30773,N_29232,N_29193);
or U30774 (N_30774,N_29736,N_29630);
xor U30775 (N_30775,N_29608,N_29973);
nor U30776 (N_30776,N_29083,N_29903);
nor U30777 (N_30777,N_29353,N_29525);
nand U30778 (N_30778,N_29262,N_29574);
and U30779 (N_30779,N_29886,N_29692);
xnor U30780 (N_30780,N_29370,N_29103);
nor U30781 (N_30781,N_29037,N_29897);
nor U30782 (N_30782,N_29073,N_29525);
nor U30783 (N_30783,N_29433,N_29889);
nand U30784 (N_30784,N_29128,N_29670);
or U30785 (N_30785,N_29920,N_29245);
or U30786 (N_30786,N_29737,N_29858);
nor U30787 (N_30787,N_29005,N_29978);
and U30788 (N_30788,N_29213,N_29289);
nor U30789 (N_30789,N_29459,N_29565);
xor U30790 (N_30790,N_29898,N_29809);
and U30791 (N_30791,N_29725,N_29072);
nor U30792 (N_30792,N_29636,N_29977);
xnor U30793 (N_30793,N_29411,N_29040);
nand U30794 (N_30794,N_29667,N_29799);
nand U30795 (N_30795,N_29879,N_29503);
nor U30796 (N_30796,N_29219,N_29057);
xor U30797 (N_30797,N_29621,N_29912);
nor U30798 (N_30798,N_29181,N_29230);
and U30799 (N_30799,N_29718,N_29081);
or U30800 (N_30800,N_29995,N_29952);
xor U30801 (N_30801,N_29662,N_29075);
and U30802 (N_30802,N_29694,N_29056);
nor U30803 (N_30803,N_29487,N_29970);
xnor U30804 (N_30804,N_29915,N_29030);
or U30805 (N_30805,N_29783,N_29049);
or U30806 (N_30806,N_29369,N_29088);
nand U30807 (N_30807,N_29304,N_29774);
nor U30808 (N_30808,N_29814,N_29629);
and U30809 (N_30809,N_29880,N_29364);
nand U30810 (N_30810,N_29665,N_29151);
nand U30811 (N_30811,N_29726,N_29076);
xnor U30812 (N_30812,N_29125,N_29319);
or U30813 (N_30813,N_29825,N_29108);
nor U30814 (N_30814,N_29553,N_29644);
nand U30815 (N_30815,N_29847,N_29175);
nor U30816 (N_30816,N_29413,N_29259);
or U30817 (N_30817,N_29725,N_29782);
or U30818 (N_30818,N_29635,N_29060);
xor U30819 (N_30819,N_29332,N_29766);
or U30820 (N_30820,N_29629,N_29277);
nand U30821 (N_30821,N_29998,N_29676);
nand U30822 (N_30822,N_29469,N_29481);
nand U30823 (N_30823,N_29518,N_29609);
xor U30824 (N_30824,N_29871,N_29415);
nand U30825 (N_30825,N_29368,N_29838);
xor U30826 (N_30826,N_29702,N_29761);
and U30827 (N_30827,N_29077,N_29955);
and U30828 (N_30828,N_29714,N_29730);
or U30829 (N_30829,N_29494,N_29979);
nand U30830 (N_30830,N_29992,N_29920);
or U30831 (N_30831,N_29984,N_29704);
and U30832 (N_30832,N_29662,N_29747);
or U30833 (N_30833,N_29166,N_29788);
or U30834 (N_30834,N_29365,N_29639);
nor U30835 (N_30835,N_29981,N_29300);
nand U30836 (N_30836,N_29662,N_29567);
or U30837 (N_30837,N_29562,N_29236);
xnor U30838 (N_30838,N_29027,N_29410);
and U30839 (N_30839,N_29280,N_29892);
nand U30840 (N_30840,N_29776,N_29949);
xnor U30841 (N_30841,N_29348,N_29352);
nand U30842 (N_30842,N_29848,N_29896);
xor U30843 (N_30843,N_29319,N_29547);
nor U30844 (N_30844,N_29468,N_29832);
xor U30845 (N_30845,N_29110,N_29959);
nand U30846 (N_30846,N_29350,N_29189);
nand U30847 (N_30847,N_29507,N_29508);
nand U30848 (N_30848,N_29752,N_29042);
xor U30849 (N_30849,N_29708,N_29462);
and U30850 (N_30850,N_29644,N_29775);
and U30851 (N_30851,N_29305,N_29919);
nand U30852 (N_30852,N_29287,N_29331);
xnor U30853 (N_30853,N_29386,N_29837);
nor U30854 (N_30854,N_29714,N_29634);
nor U30855 (N_30855,N_29920,N_29321);
nor U30856 (N_30856,N_29186,N_29670);
and U30857 (N_30857,N_29673,N_29514);
nand U30858 (N_30858,N_29717,N_29800);
xnor U30859 (N_30859,N_29098,N_29841);
nor U30860 (N_30860,N_29295,N_29871);
xor U30861 (N_30861,N_29269,N_29151);
nor U30862 (N_30862,N_29719,N_29531);
nor U30863 (N_30863,N_29788,N_29963);
xor U30864 (N_30864,N_29208,N_29671);
nor U30865 (N_30865,N_29197,N_29614);
nand U30866 (N_30866,N_29865,N_29058);
nor U30867 (N_30867,N_29593,N_29308);
and U30868 (N_30868,N_29163,N_29067);
and U30869 (N_30869,N_29358,N_29627);
nand U30870 (N_30870,N_29096,N_29293);
or U30871 (N_30871,N_29009,N_29863);
or U30872 (N_30872,N_29413,N_29647);
or U30873 (N_30873,N_29898,N_29786);
nor U30874 (N_30874,N_29252,N_29912);
or U30875 (N_30875,N_29875,N_29312);
xor U30876 (N_30876,N_29252,N_29458);
and U30877 (N_30877,N_29355,N_29986);
and U30878 (N_30878,N_29741,N_29582);
xor U30879 (N_30879,N_29813,N_29847);
xnor U30880 (N_30880,N_29514,N_29591);
and U30881 (N_30881,N_29991,N_29798);
or U30882 (N_30882,N_29709,N_29757);
nor U30883 (N_30883,N_29671,N_29998);
or U30884 (N_30884,N_29810,N_29173);
xor U30885 (N_30885,N_29459,N_29691);
and U30886 (N_30886,N_29822,N_29448);
nor U30887 (N_30887,N_29713,N_29726);
and U30888 (N_30888,N_29377,N_29403);
xor U30889 (N_30889,N_29444,N_29401);
nor U30890 (N_30890,N_29045,N_29305);
nand U30891 (N_30891,N_29219,N_29576);
or U30892 (N_30892,N_29969,N_29840);
xnor U30893 (N_30893,N_29635,N_29697);
and U30894 (N_30894,N_29818,N_29238);
nand U30895 (N_30895,N_29332,N_29130);
nor U30896 (N_30896,N_29227,N_29618);
xor U30897 (N_30897,N_29382,N_29357);
nand U30898 (N_30898,N_29276,N_29467);
nand U30899 (N_30899,N_29369,N_29208);
nand U30900 (N_30900,N_29488,N_29644);
and U30901 (N_30901,N_29855,N_29055);
nor U30902 (N_30902,N_29477,N_29014);
nor U30903 (N_30903,N_29609,N_29930);
and U30904 (N_30904,N_29665,N_29130);
or U30905 (N_30905,N_29567,N_29067);
nor U30906 (N_30906,N_29289,N_29679);
and U30907 (N_30907,N_29803,N_29868);
xor U30908 (N_30908,N_29652,N_29108);
xnor U30909 (N_30909,N_29429,N_29715);
and U30910 (N_30910,N_29356,N_29797);
nand U30911 (N_30911,N_29972,N_29695);
nor U30912 (N_30912,N_29469,N_29680);
xnor U30913 (N_30913,N_29194,N_29187);
nor U30914 (N_30914,N_29992,N_29269);
xor U30915 (N_30915,N_29414,N_29927);
and U30916 (N_30916,N_29514,N_29822);
nand U30917 (N_30917,N_29565,N_29102);
nor U30918 (N_30918,N_29413,N_29086);
xor U30919 (N_30919,N_29506,N_29697);
and U30920 (N_30920,N_29467,N_29745);
nand U30921 (N_30921,N_29089,N_29467);
or U30922 (N_30922,N_29297,N_29322);
and U30923 (N_30923,N_29195,N_29537);
and U30924 (N_30924,N_29707,N_29973);
or U30925 (N_30925,N_29279,N_29856);
or U30926 (N_30926,N_29601,N_29994);
nand U30927 (N_30927,N_29607,N_29577);
and U30928 (N_30928,N_29842,N_29726);
or U30929 (N_30929,N_29870,N_29349);
and U30930 (N_30930,N_29320,N_29409);
nor U30931 (N_30931,N_29267,N_29154);
nand U30932 (N_30932,N_29336,N_29428);
and U30933 (N_30933,N_29673,N_29106);
and U30934 (N_30934,N_29932,N_29784);
nor U30935 (N_30935,N_29290,N_29472);
and U30936 (N_30936,N_29073,N_29526);
nand U30937 (N_30937,N_29180,N_29984);
or U30938 (N_30938,N_29188,N_29120);
xor U30939 (N_30939,N_29770,N_29057);
nand U30940 (N_30940,N_29233,N_29662);
and U30941 (N_30941,N_29082,N_29786);
xnor U30942 (N_30942,N_29790,N_29510);
xor U30943 (N_30943,N_29206,N_29739);
nor U30944 (N_30944,N_29915,N_29653);
and U30945 (N_30945,N_29776,N_29244);
nor U30946 (N_30946,N_29645,N_29802);
and U30947 (N_30947,N_29533,N_29507);
xor U30948 (N_30948,N_29592,N_29292);
or U30949 (N_30949,N_29959,N_29847);
xor U30950 (N_30950,N_29484,N_29297);
nand U30951 (N_30951,N_29466,N_29012);
or U30952 (N_30952,N_29639,N_29655);
xnor U30953 (N_30953,N_29173,N_29616);
nand U30954 (N_30954,N_29587,N_29624);
nor U30955 (N_30955,N_29260,N_29906);
and U30956 (N_30956,N_29932,N_29769);
and U30957 (N_30957,N_29277,N_29602);
and U30958 (N_30958,N_29477,N_29110);
or U30959 (N_30959,N_29488,N_29341);
and U30960 (N_30960,N_29175,N_29996);
nor U30961 (N_30961,N_29567,N_29895);
xnor U30962 (N_30962,N_29948,N_29894);
or U30963 (N_30963,N_29246,N_29932);
xnor U30964 (N_30964,N_29425,N_29954);
and U30965 (N_30965,N_29309,N_29935);
nand U30966 (N_30966,N_29109,N_29812);
xor U30967 (N_30967,N_29212,N_29904);
or U30968 (N_30968,N_29811,N_29987);
or U30969 (N_30969,N_29083,N_29677);
nor U30970 (N_30970,N_29828,N_29385);
or U30971 (N_30971,N_29822,N_29812);
nor U30972 (N_30972,N_29845,N_29137);
and U30973 (N_30973,N_29225,N_29779);
and U30974 (N_30974,N_29180,N_29007);
and U30975 (N_30975,N_29247,N_29903);
nand U30976 (N_30976,N_29170,N_29524);
nor U30977 (N_30977,N_29069,N_29043);
xor U30978 (N_30978,N_29505,N_29457);
xor U30979 (N_30979,N_29910,N_29038);
nand U30980 (N_30980,N_29318,N_29456);
nor U30981 (N_30981,N_29725,N_29405);
or U30982 (N_30982,N_29236,N_29905);
xor U30983 (N_30983,N_29254,N_29053);
nor U30984 (N_30984,N_29341,N_29964);
nor U30985 (N_30985,N_29537,N_29220);
and U30986 (N_30986,N_29547,N_29236);
or U30987 (N_30987,N_29533,N_29489);
nor U30988 (N_30988,N_29297,N_29300);
nand U30989 (N_30989,N_29627,N_29382);
xnor U30990 (N_30990,N_29027,N_29547);
and U30991 (N_30991,N_29653,N_29283);
nand U30992 (N_30992,N_29429,N_29317);
and U30993 (N_30993,N_29178,N_29146);
xor U30994 (N_30994,N_29413,N_29370);
and U30995 (N_30995,N_29794,N_29436);
nand U30996 (N_30996,N_29902,N_29813);
xnor U30997 (N_30997,N_29124,N_29792);
and U30998 (N_30998,N_29217,N_29497);
xnor U30999 (N_30999,N_29354,N_29326);
and U31000 (N_31000,N_30509,N_30484);
xnor U31001 (N_31001,N_30421,N_30016);
and U31002 (N_31002,N_30606,N_30921);
xnor U31003 (N_31003,N_30204,N_30680);
or U31004 (N_31004,N_30405,N_30822);
nand U31005 (N_31005,N_30562,N_30592);
and U31006 (N_31006,N_30503,N_30635);
and U31007 (N_31007,N_30798,N_30220);
nand U31008 (N_31008,N_30830,N_30681);
nor U31009 (N_31009,N_30231,N_30664);
or U31010 (N_31010,N_30886,N_30683);
nand U31011 (N_31011,N_30194,N_30237);
nor U31012 (N_31012,N_30604,N_30410);
nor U31013 (N_31013,N_30071,N_30124);
nand U31014 (N_31014,N_30967,N_30435);
or U31015 (N_31015,N_30702,N_30618);
xor U31016 (N_31016,N_30156,N_30375);
nor U31017 (N_31017,N_30729,N_30443);
and U31018 (N_31018,N_30189,N_30235);
or U31019 (N_31019,N_30361,N_30153);
and U31020 (N_31020,N_30021,N_30179);
and U31021 (N_31021,N_30232,N_30873);
xnor U31022 (N_31022,N_30453,N_30505);
nor U31023 (N_31023,N_30811,N_30900);
nand U31024 (N_31024,N_30565,N_30837);
nor U31025 (N_31025,N_30667,N_30968);
xor U31026 (N_31026,N_30706,N_30715);
nor U31027 (N_31027,N_30936,N_30623);
or U31028 (N_31028,N_30521,N_30908);
and U31029 (N_31029,N_30969,N_30858);
nand U31030 (N_31030,N_30863,N_30791);
nor U31031 (N_31031,N_30613,N_30965);
nand U31032 (N_31032,N_30054,N_30763);
nor U31033 (N_31033,N_30458,N_30083);
and U31034 (N_31034,N_30317,N_30076);
and U31035 (N_31035,N_30332,N_30834);
nor U31036 (N_31036,N_30695,N_30622);
xor U31037 (N_31037,N_30499,N_30903);
or U31038 (N_31038,N_30414,N_30947);
xor U31039 (N_31039,N_30923,N_30734);
xor U31040 (N_31040,N_30784,N_30335);
xor U31041 (N_31041,N_30993,N_30496);
and U31042 (N_31042,N_30704,N_30452);
or U31043 (N_31043,N_30411,N_30052);
xnor U31044 (N_31044,N_30497,N_30018);
or U31045 (N_31045,N_30001,N_30190);
or U31046 (N_31046,N_30213,N_30493);
and U31047 (N_31047,N_30563,N_30673);
xor U31048 (N_31048,N_30044,N_30318);
nor U31049 (N_31049,N_30262,N_30730);
nor U31050 (N_31050,N_30924,N_30469);
nand U31051 (N_31051,N_30017,N_30531);
nor U31052 (N_31052,N_30420,N_30254);
or U31053 (N_31053,N_30196,N_30860);
and U31054 (N_31054,N_30275,N_30561);
nand U31055 (N_31055,N_30431,N_30226);
and U31056 (N_31056,N_30754,N_30333);
nor U31057 (N_31057,N_30627,N_30210);
nor U31058 (N_31058,N_30475,N_30963);
or U31059 (N_31059,N_30060,N_30841);
xnor U31060 (N_31060,N_30387,N_30856);
xor U31061 (N_31061,N_30670,N_30719);
xnor U31062 (N_31062,N_30535,N_30488);
and U31063 (N_31063,N_30518,N_30019);
nand U31064 (N_31064,N_30129,N_30632);
or U31065 (N_31065,N_30176,N_30109);
xor U31066 (N_31066,N_30705,N_30331);
nor U31067 (N_31067,N_30642,N_30624);
xnor U31068 (N_31068,N_30161,N_30160);
xnor U31069 (N_31069,N_30755,N_30185);
or U31070 (N_31070,N_30494,N_30649);
or U31071 (N_31071,N_30788,N_30316);
nor U31072 (N_31072,N_30504,N_30540);
or U31073 (N_31073,N_30888,N_30739);
nor U31074 (N_31074,N_30010,N_30417);
nand U31075 (N_31075,N_30820,N_30720);
and U31076 (N_31076,N_30412,N_30193);
and U31077 (N_31077,N_30108,N_30004);
nand U31078 (N_31078,N_30438,N_30802);
nor U31079 (N_31079,N_30195,N_30750);
xor U31080 (N_31080,N_30264,N_30177);
or U31081 (N_31081,N_30013,N_30512);
xnor U31082 (N_31082,N_30736,N_30214);
xor U31083 (N_31083,N_30997,N_30353);
and U31084 (N_31084,N_30343,N_30957);
or U31085 (N_31085,N_30815,N_30290);
nor U31086 (N_31086,N_30139,N_30660);
nand U31087 (N_31087,N_30869,N_30517);
and U31088 (N_31088,N_30534,N_30383);
nor U31089 (N_31089,N_30300,N_30693);
and U31090 (N_31090,N_30897,N_30182);
and U31091 (N_31091,N_30883,N_30146);
nor U31092 (N_31092,N_30910,N_30790);
or U31093 (N_31093,N_30772,N_30418);
nand U31094 (N_31094,N_30057,N_30898);
nand U31095 (N_31095,N_30575,N_30662);
nor U31096 (N_31096,N_30832,N_30793);
nor U31097 (N_31097,N_30106,N_30741);
nor U31098 (N_31098,N_30848,N_30944);
nor U31099 (N_31099,N_30892,N_30581);
or U31100 (N_31100,N_30197,N_30943);
and U31101 (N_31101,N_30015,N_30567);
and U31102 (N_31102,N_30777,N_30404);
nor U31103 (N_31103,N_30323,N_30771);
nor U31104 (N_31104,N_30979,N_30896);
xor U31105 (N_31105,N_30637,N_30255);
or U31106 (N_31106,N_30816,N_30389);
nor U31107 (N_31107,N_30654,N_30099);
xnor U31108 (N_31108,N_30895,N_30628);
nand U31109 (N_31109,N_30425,N_30966);
or U31110 (N_31110,N_30173,N_30625);
or U31111 (N_31111,N_30620,N_30442);
nor U31112 (N_31112,N_30906,N_30448);
or U31113 (N_31113,N_30158,N_30279);
and U31114 (N_31114,N_30629,N_30064);
xor U31115 (N_31115,N_30223,N_30587);
xor U31116 (N_31116,N_30296,N_30803);
nand U31117 (N_31117,N_30265,N_30258);
nor U31118 (N_31118,N_30133,N_30689);
nor U31119 (N_31119,N_30519,N_30167);
nand U31120 (N_31120,N_30073,N_30520);
nand U31121 (N_31121,N_30961,N_30838);
xnor U31122 (N_31122,N_30070,N_30962);
nor U31123 (N_31123,N_30263,N_30655);
or U31124 (N_31124,N_30676,N_30240);
nor U31125 (N_31125,N_30596,N_30269);
or U31126 (N_31126,N_30023,N_30684);
nand U31127 (N_31127,N_30590,N_30981);
and U31128 (N_31128,N_30477,N_30393);
and U31129 (N_31129,N_30674,N_30359);
xor U31130 (N_31130,N_30585,N_30381);
nor U31131 (N_31131,N_30239,N_30074);
nor U31132 (N_31132,N_30862,N_30697);
or U31133 (N_31133,N_30145,N_30956);
and U31134 (N_31134,N_30636,N_30914);
nand U31135 (N_31135,N_30125,N_30761);
or U31136 (N_31136,N_30261,N_30135);
xnor U31137 (N_31137,N_30857,N_30441);
xnor U31138 (N_31138,N_30349,N_30447);
and U31139 (N_31139,N_30002,N_30692);
or U31140 (N_31140,N_30882,N_30564);
or U31141 (N_31141,N_30992,N_30779);
and U31142 (N_31142,N_30360,N_30691);
and U31143 (N_31143,N_30374,N_30927);
nand U31144 (N_31144,N_30462,N_30933);
and U31145 (N_31145,N_30753,N_30200);
or U31146 (N_31146,N_30183,N_30707);
nor U31147 (N_31147,N_30097,N_30789);
or U31148 (N_31148,N_30492,N_30292);
and U31149 (N_31149,N_30334,N_30942);
xor U31150 (N_31150,N_30000,N_30994);
or U31151 (N_31151,N_30971,N_30209);
xor U31152 (N_31152,N_30887,N_30170);
and U31153 (N_31153,N_30029,N_30487);
nand U31154 (N_31154,N_30749,N_30319);
and U31155 (N_31155,N_30775,N_30650);
and U31156 (N_31156,N_30807,N_30571);
or U31157 (N_31157,N_30473,N_30868);
nand U31158 (N_31158,N_30014,N_30935);
xor U31159 (N_31159,N_30817,N_30075);
nor U31160 (N_31160,N_30552,N_30424);
or U31161 (N_31161,N_30368,N_30917);
xnor U31162 (N_31162,N_30941,N_30355);
and U31163 (N_31163,N_30039,N_30267);
nand U31164 (N_31164,N_30086,N_30364);
or U31165 (N_31165,N_30102,N_30234);
xor U31166 (N_31166,N_30370,N_30061);
and U31167 (N_31167,N_30049,N_30259);
or U31168 (N_31168,N_30459,N_30416);
nor U31169 (N_31169,N_30216,N_30247);
nor U31170 (N_31170,N_30825,N_30350);
xnor U31171 (N_31171,N_30938,N_30651);
and U31172 (N_31172,N_30806,N_30491);
xor U31173 (N_31173,N_30329,N_30630);
nor U31174 (N_31174,N_30640,N_30178);
nor U31175 (N_31175,N_30770,N_30143);
or U31176 (N_31176,N_30758,N_30767);
and U31177 (N_31177,N_30845,N_30105);
nor U31178 (N_31178,N_30808,N_30095);
or U31179 (N_31179,N_30212,N_30276);
or U31180 (N_31180,N_30025,N_30022);
xnor U31181 (N_31181,N_30043,N_30168);
xnor U31182 (N_31182,N_30399,N_30085);
nand U31183 (N_31183,N_30294,N_30050);
or U31184 (N_31184,N_30123,N_30644);
nand U31185 (N_31185,N_30877,N_30037);
nand U31186 (N_31186,N_30429,N_30909);
xnor U31187 (N_31187,N_30396,N_30946);
or U31188 (N_31188,N_30445,N_30768);
and U31189 (N_31189,N_30859,N_30465);
and U31190 (N_31190,N_30184,N_30550);
or U31191 (N_31191,N_30042,N_30568);
or U31192 (N_31192,N_30077,N_30867);
nand U31193 (N_31193,N_30631,N_30011);
nor U31194 (N_31194,N_30744,N_30723);
and U31195 (N_31195,N_30668,N_30919);
and U31196 (N_31196,N_30752,N_30608);
or U31197 (N_31197,N_30787,N_30082);
or U31198 (N_31198,N_30030,N_30257);
nand U31199 (N_31199,N_30566,N_30524);
xnor U31200 (N_31200,N_30471,N_30051);
nor U31201 (N_31201,N_30401,N_30577);
and U31202 (N_31202,N_30298,N_30849);
and U31203 (N_31203,N_30669,N_30155);
xor U31204 (N_31204,N_30395,N_30774);
nand U31205 (N_31205,N_30315,N_30485);
xor U31206 (N_31206,N_30498,N_30242);
or U31207 (N_31207,N_30324,N_30751);
nand U31208 (N_31208,N_30376,N_30615);
nand U31209 (N_31209,N_30081,N_30989);
nand U31210 (N_31210,N_30136,N_30764);
xor U31211 (N_31211,N_30999,N_30740);
or U31212 (N_31212,N_30152,N_30913);
and U31213 (N_31213,N_30973,N_30652);
xnor U31214 (N_31214,N_30326,N_30369);
nand U31215 (N_31215,N_30301,N_30172);
and U31216 (N_31216,N_30211,N_30960);
nor U31217 (N_31217,N_30871,N_30388);
or U31218 (N_31218,N_30525,N_30926);
and U31219 (N_31219,N_30078,N_30474);
nor U31220 (N_31220,N_30407,N_30809);
xnor U31221 (N_31221,N_30657,N_30422);
and U31222 (N_31222,N_30142,N_30058);
nor U31223 (N_31223,N_30544,N_30020);
nor U31224 (N_31224,N_30778,N_30948);
or U31225 (N_31225,N_30783,N_30773);
and U31226 (N_31226,N_30026,N_30826);
nand U31227 (N_31227,N_30786,N_30154);
nor U31228 (N_31228,N_30688,N_30502);
and U31229 (N_31229,N_30354,N_30894);
nor U31230 (N_31230,N_30527,N_30277);
nor U31231 (N_31231,N_30780,N_30582);
or U31232 (N_31232,N_30415,N_30975);
or U31233 (N_31233,N_30104,N_30716);
and U31234 (N_31234,N_30905,N_30330);
xnor U31235 (N_31235,N_30089,N_30548);
and U31236 (N_31236,N_30621,N_30677);
nand U31237 (N_31237,N_30922,N_30365);
and U31238 (N_31238,N_30874,N_30202);
and U31239 (N_31239,N_30814,N_30479);
nor U31240 (N_31240,N_30675,N_30286);
xor U31241 (N_31241,N_30358,N_30252);
xnor U31242 (N_31242,N_30157,N_30040);
and U31243 (N_31243,N_30273,N_30976);
nand U31244 (N_31244,N_30824,N_30311);
nand U31245 (N_31245,N_30547,N_30915);
nand U31246 (N_31246,N_30672,N_30150);
nor U31247 (N_31247,N_30983,N_30437);
nor U31248 (N_31248,N_30352,N_30542);
and U31249 (N_31249,N_30690,N_30970);
nor U31250 (N_31250,N_30743,N_30954);
xnor U31251 (N_31251,N_30470,N_30732);
nor U31252 (N_31252,N_30828,N_30737);
and U31253 (N_31253,N_30367,N_30612);
nor U31254 (N_31254,N_30593,N_30041);
nor U31255 (N_31255,N_30510,N_30466);
nor U31256 (N_31256,N_30686,N_30610);
nor U31257 (N_31257,N_30937,N_30557);
or U31258 (N_31258,N_30117,N_30794);
and U31259 (N_31259,N_30746,N_30248);
and U31260 (N_31260,N_30928,N_30047);
xor U31261 (N_31261,N_30038,N_30745);
nand U31262 (N_31262,N_30710,N_30634);
xnor U31263 (N_31263,N_30701,N_30907);
nor U31264 (N_31264,N_30765,N_30472);
nor U31265 (N_31265,N_30756,N_30080);
nor U31266 (N_31266,N_30322,N_30506);
nand U31267 (N_31267,N_30428,N_30112);
and U31268 (N_31268,N_30454,N_30536);
xnor U31269 (N_31269,N_30647,N_30884);
and U31270 (N_31270,N_30875,N_30034);
xor U31271 (N_31271,N_30804,N_30363);
nor U31272 (N_31272,N_30299,N_30511);
nand U31273 (N_31273,N_30096,N_30107);
and U31274 (N_31274,N_30529,N_30394);
and U31275 (N_31275,N_30222,N_30084);
nor U31276 (N_31276,N_30059,N_30293);
nand U31277 (N_31277,N_30995,N_30591);
and U31278 (N_31278,N_30379,N_30762);
and U31279 (N_31279,N_30617,N_30451);
nor U31280 (N_31280,N_30377,N_30988);
xor U31281 (N_31281,N_30588,N_30666);
xnor U31282 (N_31282,N_30633,N_30818);
nand U31283 (N_31283,N_30218,N_30539);
or U31284 (N_31284,N_30813,N_30118);
and U31285 (N_31285,N_30409,N_30574);
nor U31286 (N_31286,N_30166,N_30931);
nand U31287 (N_31287,N_30440,N_30310);
nand U31288 (N_31288,N_30855,N_30785);
nor U31289 (N_31289,N_30008,N_30847);
nand U31290 (N_31290,N_30031,N_30427);
xor U31291 (N_31291,N_30284,N_30062);
xor U31292 (N_31292,N_30821,N_30243);
nor U31293 (N_31293,N_30130,N_30313);
xor U31294 (N_31294,N_30805,N_30795);
nor U31295 (N_31295,N_30238,N_30162);
nand U31296 (N_31296,N_30092,N_30554);
xor U31297 (N_31297,N_30230,N_30700);
nor U31298 (N_31298,N_30920,N_30229);
and U31299 (N_31299,N_30221,N_30551);
and U31300 (N_31300,N_30345,N_30980);
nor U31301 (N_31301,N_30328,N_30602);
nand U31302 (N_31302,N_30866,N_30678);
or U31303 (N_31303,N_30726,N_30287);
nor U31304 (N_31304,N_30978,N_30297);
nor U31305 (N_31305,N_30757,N_30072);
nand U31306 (N_31306,N_30735,N_30147);
nand U31307 (N_31307,N_30712,N_30048);
xor U31308 (N_31308,N_30289,N_30100);
nand U31309 (N_31309,N_30308,N_30573);
nand U31310 (N_31310,N_30271,N_30281);
or U31311 (N_31311,N_30952,N_30274);
xor U31312 (N_31312,N_30653,N_30932);
and U31313 (N_31313,N_30836,N_30207);
nand U31314 (N_31314,N_30586,N_30638);
nor U31315 (N_31315,N_30346,N_30731);
nor U31316 (N_31316,N_30246,N_30904);
or U31317 (N_31317,N_30115,N_30314);
or U31318 (N_31318,N_30199,N_30439);
nand U31319 (N_31319,N_30164,N_30482);
nand U31320 (N_31320,N_30141,N_30413);
xor U31321 (N_31321,N_30005,N_30063);
xor U31322 (N_31322,N_30865,N_30645);
nor U31323 (N_31323,N_30486,N_30722);
or U31324 (N_31324,N_30801,N_30530);
and U31325 (N_31325,N_30351,N_30348);
and U31326 (N_31326,N_30419,N_30468);
xor U31327 (N_31327,N_30386,N_30120);
nand U31328 (N_31328,N_30027,N_30426);
and U31329 (N_31329,N_30347,N_30169);
and U31330 (N_31330,N_30341,N_30951);
and U31331 (N_31331,N_30569,N_30852);
and U31332 (N_31332,N_30984,N_30872);
or U31333 (N_31333,N_30955,N_30291);
xor U31334 (N_31334,N_30977,N_30879);
or U31335 (N_31335,N_30579,N_30727);
nor U31336 (N_31336,N_30366,N_30028);
nand U31337 (N_31337,N_30457,N_30890);
nand U31338 (N_31338,N_30748,N_30217);
nor U31339 (N_31339,N_30390,N_30843);
and U31340 (N_31340,N_30782,N_30225);
and U31341 (N_31341,N_30434,N_30609);
and U31342 (N_31342,N_30595,N_30703);
nor U31343 (N_31343,N_30219,N_30639);
nor U31344 (N_31344,N_30699,N_30528);
xor U31345 (N_31345,N_30066,N_30641);
nand U31346 (N_31346,N_30698,N_30507);
nor U31347 (N_31347,N_30304,N_30605);
nand U31348 (N_31348,N_30121,N_30449);
or U31349 (N_31349,N_30934,N_30228);
xnor U31350 (N_31350,N_30796,N_30823);
xnor U31351 (N_31351,N_30035,N_30171);
or U31352 (N_31352,N_30131,N_30972);
nand U31353 (N_31353,N_30456,N_30578);
or U31354 (N_31354,N_30854,N_30024);
nor U31355 (N_31355,N_30305,N_30088);
or U31356 (N_31356,N_30810,N_30893);
nor U31357 (N_31357,N_30831,N_30490);
xnor U31358 (N_31358,N_30087,N_30268);
or U31359 (N_31359,N_30839,N_30398);
nor U31360 (N_31360,N_30513,N_30881);
xor U31361 (N_31361,N_30522,N_30840);
xor U31362 (N_31362,N_30378,N_30256);
xor U31363 (N_31363,N_30583,N_30656);
nor U31364 (N_31364,N_30373,N_30385);
xor U31365 (N_31365,N_30400,N_30713);
nand U31366 (N_31366,N_30514,N_30009);
or U31367 (N_31367,N_30140,N_30306);
nor U31368 (N_31368,N_30889,N_30516);
and U31369 (N_31369,N_30844,N_30558);
nand U31370 (N_31370,N_30094,N_30260);
nor U31371 (N_31371,N_30175,N_30007);
xnor U31372 (N_31372,N_30853,N_30481);
nor U31373 (N_31373,N_30045,N_30250);
or U31374 (N_31374,N_30208,N_30188);
nor U31375 (N_31375,N_30283,N_30103);
and U31376 (N_31376,N_30101,N_30724);
nand U31377 (N_31377,N_30646,N_30114);
or U31378 (N_31378,N_30594,N_30584);
xor U31379 (N_31379,N_30959,N_30526);
and U31380 (N_31380,N_30733,N_30990);
xor U31381 (N_31381,N_30930,N_30278);
xor U31382 (N_31382,N_30601,N_30643);
and U31383 (N_31383,N_30397,N_30245);
and U31384 (N_31384,N_30191,N_30392);
nor U31385 (N_31385,N_30012,N_30149);
or U31386 (N_31386,N_30053,N_30382);
and U31387 (N_31387,N_30201,N_30861);
nand U31388 (N_31388,N_30537,N_30949);
and U31389 (N_31389,N_30891,N_30682);
nand U31390 (N_31390,N_30648,N_30307);
xor U31391 (N_31391,N_30523,N_30320);
and U31392 (N_31392,N_30126,N_30068);
and U31393 (N_31393,N_30899,N_30603);
and U31394 (N_31394,N_30549,N_30056);
or U31395 (N_31395,N_30340,N_30192);
nor U31396 (N_31396,N_30996,N_30998);
or U31397 (N_31397,N_30325,N_30950);
nor U31398 (N_31398,N_30819,N_30864);
and U31399 (N_31399,N_30272,N_30288);
nand U31400 (N_31400,N_30384,N_30541);
and U31401 (N_31401,N_30236,N_30455);
and U31402 (N_31402,N_30151,N_30885);
or U31403 (N_31403,N_30911,N_30708);
nand U31404 (N_31404,N_30543,N_30134);
and U31405 (N_31405,N_30444,N_30111);
nor U31406 (N_31406,N_30781,N_30402);
or U31407 (N_31407,N_30538,N_30128);
and U31408 (N_31408,N_30846,N_30776);
and U31409 (N_31409,N_30792,N_30501);
nand U31410 (N_31410,N_30233,N_30203);
nand U31411 (N_31411,N_30337,N_30186);
or U31412 (N_31412,N_30122,N_30312);
or U31413 (N_31413,N_30769,N_30835);
and U31414 (N_31414,N_30423,N_30721);
and U31415 (N_31415,N_30659,N_30067);
xnor U31416 (N_31416,N_30555,N_30616);
or U31417 (N_31417,N_30483,N_30093);
nand U31418 (N_31418,N_30215,N_30137);
xor U31419 (N_31419,N_30430,N_30282);
and U31420 (N_31420,N_30991,N_30597);
or U31421 (N_31421,N_30138,N_30295);
nor U31422 (N_31422,N_30032,N_30827);
nand U31423 (N_31423,N_30687,N_30180);
or U31424 (N_31424,N_30036,N_30945);
nor U31425 (N_31425,N_30940,N_30336);
nor U31426 (N_31426,N_30829,N_30205);
nor U31427 (N_31427,N_30033,N_30851);
nor U31428 (N_31428,N_30987,N_30850);
and U31429 (N_31429,N_30589,N_30572);
or U31430 (N_31430,N_30546,N_30685);
xor U31431 (N_31431,N_30266,N_30148);
and U31432 (N_31432,N_30939,N_30280);
nor U31433 (N_31433,N_30515,N_30356);
and U31434 (N_31434,N_30165,N_30742);
and U31435 (N_31435,N_30251,N_30461);
nor U31436 (N_31436,N_30738,N_30436);
nor U31437 (N_31437,N_30241,N_30302);
xor U31438 (N_31438,N_30450,N_30500);
nor U31439 (N_31439,N_30508,N_30912);
nand U31440 (N_31440,N_30974,N_30065);
xnor U31441 (N_31441,N_30559,N_30665);
and U31442 (N_31442,N_30694,N_30132);
and U31443 (N_31443,N_30362,N_30055);
or U31444 (N_31444,N_30460,N_30598);
or U31445 (N_31445,N_30728,N_30116);
and U31446 (N_31446,N_30342,N_30159);
and U31447 (N_31447,N_30476,N_30303);
nor U31448 (N_31448,N_30187,N_30925);
nor U31449 (N_31449,N_30480,N_30406);
and U31450 (N_31450,N_30321,N_30982);
nand U31451 (N_31451,N_30679,N_30463);
nand U31452 (N_31452,N_30986,N_30626);
nand U31453 (N_31453,N_30929,N_30098);
and U31454 (N_31454,N_30576,N_30339);
and U31455 (N_31455,N_30718,N_30725);
nor U31456 (N_31456,N_30580,N_30696);
xor U31457 (N_31457,N_30403,N_30599);
nand U31458 (N_31458,N_30113,N_30489);
or U31459 (N_31459,N_30357,N_30880);
nor U31460 (N_31460,N_30614,N_30953);
xnor U31461 (N_31461,N_30163,N_30532);
or U31462 (N_31462,N_30227,N_30711);
nor U31463 (N_31463,N_30717,N_30270);
xnor U31464 (N_31464,N_30478,N_30812);
or U31465 (N_31465,N_30760,N_30709);
and U31466 (N_31466,N_30570,N_30408);
nor U31467 (N_31467,N_30876,N_30800);
or U31468 (N_31468,N_30611,N_30842);
xor U31469 (N_31469,N_30174,N_30918);
or U31470 (N_31470,N_30901,N_30003);
xor U31471 (N_31471,N_30958,N_30338);
or U31472 (N_31472,N_30619,N_30467);
or U31473 (N_31473,N_30380,N_30079);
or U31474 (N_31474,N_30069,N_30902);
nand U31475 (N_31475,N_30556,N_30006);
xnor U31476 (N_31476,N_30607,N_30446);
nand U31477 (N_31477,N_30253,N_30495);
nor U31478 (N_31478,N_30371,N_30964);
and U31479 (N_31479,N_30119,N_30714);
or U31480 (N_31480,N_30249,N_30285);
or U31481 (N_31481,N_30110,N_30127);
xnor U31482 (N_31482,N_30799,N_30797);
xnor U31483 (N_31483,N_30464,N_30833);
nor U31484 (N_31484,N_30391,N_30747);
and U31485 (N_31485,N_30766,N_30878);
and U31486 (N_31486,N_30244,N_30916);
and U31487 (N_31487,N_30560,N_30658);
or U31488 (N_31488,N_30046,N_30870);
nand U31489 (N_31489,N_30327,N_30671);
nor U31490 (N_31490,N_30432,N_30181);
or U31491 (N_31491,N_30553,N_30663);
nand U31492 (N_31492,N_30545,N_30090);
nor U31493 (N_31493,N_30433,N_30985);
and U31494 (N_31494,N_30198,N_30372);
nand U31495 (N_31495,N_30661,N_30533);
nand U31496 (N_31496,N_30309,N_30344);
nor U31497 (N_31497,N_30759,N_30144);
xor U31498 (N_31498,N_30600,N_30091);
xnor U31499 (N_31499,N_30224,N_30206);
nand U31500 (N_31500,N_30483,N_30267);
xor U31501 (N_31501,N_30420,N_30403);
or U31502 (N_31502,N_30222,N_30396);
nor U31503 (N_31503,N_30559,N_30666);
or U31504 (N_31504,N_30943,N_30658);
or U31505 (N_31505,N_30276,N_30616);
and U31506 (N_31506,N_30125,N_30137);
and U31507 (N_31507,N_30077,N_30371);
nand U31508 (N_31508,N_30742,N_30133);
and U31509 (N_31509,N_30019,N_30453);
or U31510 (N_31510,N_30030,N_30310);
and U31511 (N_31511,N_30453,N_30585);
or U31512 (N_31512,N_30286,N_30905);
nor U31513 (N_31513,N_30971,N_30424);
and U31514 (N_31514,N_30184,N_30283);
nor U31515 (N_31515,N_30057,N_30225);
xnor U31516 (N_31516,N_30748,N_30607);
xnor U31517 (N_31517,N_30280,N_30974);
and U31518 (N_31518,N_30918,N_30580);
nor U31519 (N_31519,N_30082,N_30762);
nor U31520 (N_31520,N_30521,N_30158);
or U31521 (N_31521,N_30549,N_30544);
and U31522 (N_31522,N_30310,N_30113);
or U31523 (N_31523,N_30933,N_30908);
and U31524 (N_31524,N_30841,N_30888);
or U31525 (N_31525,N_30412,N_30656);
nand U31526 (N_31526,N_30968,N_30737);
and U31527 (N_31527,N_30438,N_30084);
and U31528 (N_31528,N_30985,N_30884);
nor U31529 (N_31529,N_30424,N_30054);
nand U31530 (N_31530,N_30813,N_30272);
or U31531 (N_31531,N_30807,N_30300);
and U31532 (N_31532,N_30441,N_30012);
xor U31533 (N_31533,N_30104,N_30912);
nand U31534 (N_31534,N_30933,N_30777);
and U31535 (N_31535,N_30082,N_30031);
or U31536 (N_31536,N_30326,N_30390);
xnor U31537 (N_31537,N_30274,N_30132);
or U31538 (N_31538,N_30998,N_30382);
nor U31539 (N_31539,N_30642,N_30117);
or U31540 (N_31540,N_30389,N_30480);
xnor U31541 (N_31541,N_30180,N_30453);
nor U31542 (N_31542,N_30011,N_30882);
nand U31543 (N_31543,N_30724,N_30161);
nor U31544 (N_31544,N_30864,N_30908);
or U31545 (N_31545,N_30145,N_30636);
nand U31546 (N_31546,N_30455,N_30485);
xnor U31547 (N_31547,N_30663,N_30574);
and U31548 (N_31548,N_30799,N_30623);
and U31549 (N_31549,N_30270,N_30825);
nor U31550 (N_31550,N_30136,N_30785);
or U31551 (N_31551,N_30586,N_30113);
and U31552 (N_31552,N_30381,N_30497);
or U31553 (N_31553,N_30808,N_30884);
xor U31554 (N_31554,N_30800,N_30178);
and U31555 (N_31555,N_30233,N_30079);
nor U31556 (N_31556,N_30512,N_30059);
nor U31557 (N_31557,N_30204,N_30800);
and U31558 (N_31558,N_30976,N_30129);
nor U31559 (N_31559,N_30379,N_30598);
nor U31560 (N_31560,N_30561,N_30493);
nand U31561 (N_31561,N_30278,N_30369);
nor U31562 (N_31562,N_30500,N_30280);
nor U31563 (N_31563,N_30659,N_30108);
and U31564 (N_31564,N_30734,N_30894);
nand U31565 (N_31565,N_30445,N_30139);
nand U31566 (N_31566,N_30255,N_30545);
or U31567 (N_31567,N_30149,N_30441);
and U31568 (N_31568,N_30245,N_30486);
nand U31569 (N_31569,N_30676,N_30000);
or U31570 (N_31570,N_30111,N_30980);
xor U31571 (N_31571,N_30497,N_30025);
nor U31572 (N_31572,N_30411,N_30329);
xnor U31573 (N_31573,N_30557,N_30652);
or U31574 (N_31574,N_30141,N_30885);
xnor U31575 (N_31575,N_30303,N_30179);
and U31576 (N_31576,N_30752,N_30997);
or U31577 (N_31577,N_30234,N_30008);
xnor U31578 (N_31578,N_30799,N_30458);
nand U31579 (N_31579,N_30547,N_30373);
nor U31580 (N_31580,N_30911,N_30482);
nor U31581 (N_31581,N_30671,N_30644);
or U31582 (N_31582,N_30221,N_30078);
and U31583 (N_31583,N_30766,N_30442);
or U31584 (N_31584,N_30859,N_30518);
and U31585 (N_31585,N_30498,N_30309);
nand U31586 (N_31586,N_30961,N_30414);
or U31587 (N_31587,N_30885,N_30389);
or U31588 (N_31588,N_30346,N_30142);
nand U31589 (N_31589,N_30722,N_30497);
or U31590 (N_31590,N_30719,N_30335);
xor U31591 (N_31591,N_30848,N_30667);
or U31592 (N_31592,N_30316,N_30913);
xnor U31593 (N_31593,N_30860,N_30723);
or U31594 (N_31594,N_30311,N_30158);
nand U31595 (N_31595,N_30441,N_30651);
or U31596 (N_31596,N_30842,N_30920);
nand U31597 (N_31597,N_30430,N_30835);
xnor U31598 (N_31598,N_30002,N_30598);
nor U31599 (N_31599,N_30533,N_30430);
nand U31600 (N_31600,N_30380,N_30623);
and U31601 (N_31601,N_30974,N_30251);
nand U31602 (N_31602,N_30452,N_30875);
and U31603 (N_31603,N_30346,N_30736);
and U31604 (N_31604,N_30853,N_30178);
or U31605 (N_31605,N_30918,N_30148);
nand U31606 (N_31606,N_30573,N_30170);
nand U31607 (N_31607,N_30501,N_30723);
nand U31608 (N_31608,N_30346,N_30893);
and U31609 (N_31609,N_30388,N_30532);
nor U31610 (N_31610,N_30006,N_30087);
or U31611 (N_31611,N_30986,N_30967);
xor U31612 (N_31612,N_30227,N_30681);
and U31613 (N_31613,N_30480,N_30796);
and U31614 (N_31614,N_30468,N_30393);
xnor U31615 (N_31615,N_30894,N_30557);
nand U31616 (N_31616,N_30690,N_30393);
nor U31617 (N_31617,N_30306,N_30564);
and U31618 (N_31618,N_30055,N_30743);
nand U31619 (N_31619,N_30203,N_30264);
nand U31620 (N_31620,N_30709,N_30312);
and U31621 (N_31621,N_30544,N_30244);
xor U31622 (N_31622,N_30298,N_30257);
and U31623 (N_31623,N_30850,N_30973);
nor U31624 (N_31624,N_30077,N_30917);
nand U31625 (N_31625,N_30166,N_30888);
or U31626 (N_31626,N_30687,N_30319);
or U31627 (N_31627,N_30832,N_30383);
xnor U31628 (N_31628,N_30180,N_30258);
nor U31629 (N_31629,N_30641,N_30340);
and U31630 (N_31630,N_30369,N_30161);
and U31631 (N_31631,N_30525,N_30204);
xor U31632 (N_31632,N_30439,N_30221);
nor U31633 (N_31633,N_30825,N_30748);
xnor U31634 (N_31634,N_30844,N_30436);
xor U31635 (N_31635,N_30727,N_30978);
nor U31636 (N_31636,N_30808,N_30079);
nor U31637 (N_31637,N_30882,N_30320);
nor U31638 (N_31638,N_30345,N_30243);
nor U31639 (N_31639,N_30370,N_30044);
xor U31640 (N_31640,N_30996,N_30641);
and U31641 (N_31641,N_30515,N_30552);
and U31642 (N_31642,N_30647,N_30866);
and U31643 (N_31643,N_30442,N_30656);
nor U31644 (N_31644,N_30328,N_30184);
xnor U31645 (N_31645,N_30993,N_30527);
and U31646 (N_31646,N_30394,N_30704);
nand U31647 (N_31647,N_30997,N_30671);
and U31648 (N_31648,N_30372,N_30158);
xor U31649 (N_31649,N_30315,N_30151);
xor U31650 (N_31650,N_30576,N_30713);
xnor U31651 (N_31651,N_30564,N_30446);
and U31652 (N_31652,N_30811,N_30749);
nor U31653 (N_31653,N_30637,N_30936);
and U31654 (N_31654,N_30118,N_30005);
xor U31655 (N_31655,N_30851,N_30801);
or U31656 (N_31656,N_30503,N_30281);
or U31657 (N_31657,N_30532,N_30412);
and U31658 (N_31658,N_30017,N_30053);
or U31659 (N_31659,N_30886,N_30408);
nor U31660 (N_31660,N_30963,N_30007);
or U31661 (N_31661,N_30369,N_30251);
xor U31662 (N_31662,N_30813,N_30799);
nor U31663 (N_31663,N_30703,N_30325);
xor U31664 (N_31664,N_30369,N_30379);
nor U31665 (N_31665,N_30036,N_30075);
xor U31666 (N_31666,N_30901,N_30532);
xnor U31667 (N_31667,N_30276,N_30866);
or U31668 (N_31668,N_30394,N_30789);
nor U31669 (N_31669,N_30719,N_30191);
or U31670 (N_31670,N_30715,N_30085);
nor U31671 (N_31671,N_30655,N_30601);
or U31672 (N_31672,N_30403,N_30366);
nor U31673 (N_31673,N_30903,N_30740);
xnor U31674 (N_31674,N_30903,N_30973);
nor U31675 (N_31675,N_30619,N_30859);
nor U31676 (N_31676,N_30424,N_30693);
xnor U31677 (N_31677,N_30373,N_30095);
or U31678 (N_31678,N_30372,N_30590);
and U31679 (N_31679,N_30051,N_30317);
nor U31680 (N_31680,N_30083,N_30919);
nor U31681 (N_31681,N_30815,N_30857);
xor U31682 (N_31682,N_30486,N_30530);
nand U31683 (N_31683,N_30954,N_30267);
xor U31684 (N_31684,N_30140,N_30353);
and U31685 (N_31685,N_30618,N_30486);
or U31686 (N_31686,N_30104,N_30621);
and U31687 (N_31687,N_30800,N_30151);
xnor U31688 (N_31688,N_30189,N_30083);
xor U31689 (N_31689,N_30922,N_30276);
or U31690 (N_31690,N_30998,N_30141);
xnor U31691 (N_31691,N_30115,N_30895);
and U31692 (N_31692,N_30888,N_30616);
and U31693 (N_31693,N_30305,N_30456);
nand U31694 (N_31694,N_30988,N_30706);
nand U31695 (N_31695,N_30742,N_30914);
nand U31696 (N_31696,N_30603,N_30308);
nor U31697 (N_31697,N_30490,N_30509);
xnor U31698 (N_31698,N_30214,N_30439);
and U31699 (N_31699,N_30318,N_30636);
xnor U31700 (N_31700,N_30193,N_30317);
nand U31701 (N_31701,N_30742,N_30583);
nor U31702 (N_31702,N_30295,N_30856);
or U31703 (N_31703,N_30435,N_30807);
xor U31704 (N_31704,N_30308,N_30001);
nand U31705 (N_31705,N_30476,N_30950);
nand U31706 (N_31706,N_30888,N_30086);
xnor U31707 (N_31707,N_30167,N_30418);
nand U31708 (N_31708,N_30403,N_30114);
or U31709 (N_31709,N_30704,N_30299);
nand U31710 (N_31710,N_30835,N_30946);
and U31711 (N_31711,N_30693,N_30210);
and U31712 (N_31712,N_30441,N_30862);
nand U31713 (N_31713,N_30114,N_30593);
xor U31714 (N_31714,N_30971,N_30054);
nand U31715 (N_31715,N_30128,N_30062);
nor U31716 (N_31716,N_30062,N_30945);
or U31717 (N_31717,N_30659,N_30691);
and U31718 (N_31718,N_30691,N_30437);
nor U31719 (N_31719,N_30400,N_30340);
and U31720 (N_31720,N_30575,N_30030);
nor U31721 (N_31721,N_30724,N_30903);
xor U31722 (N_31722,N_30117,N_30918);
nand U31723 (N_31723,N_30828,N_30921);
nor U31724 (N_31724,N_30379,N_30269);
nand U31725 (N_31725,N_30408,N_30918);
xnor U31726 (N_31726,N_30165,N_30361);
nand U31727 (N_31727,N_30759,N_30646);
nand U31728 (N_31728,N_30931,N_30971);
nand U31729 (N_31729,N_30245,N_30155);
and U31730 (N_31730,N_30515,N_30756);
or U31731 (N_31731,N_30892,N_30392);
or U31732 (N_31732,N_30031,N_30280);
nor U31733 (N_31733,N_30209,N_30359);
and U31734 (N_31734,N_30124,N_30735);
or U31735 (N_31735,N_30862,N_30692);
nor U31736 (N_31736,N_30363,N_30058);
or U31737 (N_31737,N_30854,N_30790);
nand U31738 (N_31738,N_30256,N_30056);
xnor U31739 (N_31739,N_30070,N_30205);
or U31740 (N_31740,N_30408,N_30922);
nand U31741 (N_31741,N_30076,N_30631);
xor U31742 (N_31742,N_30496,N_30600);
xnor U31743 (N_31743,N_30153,N_30767);
xnor U31744 (N_31744,N_30856,N_30098);
nor U31745 (N_31745,N_30745,N_30171);
or U31746 (N_31746,N_30731,N_30994);
nand U31747 (N_31747,N_30902,N_30678);
xnor U31748 (N_31748,N_30393,N_30787);
xnor U31749 (N_31749,N_30785,N_30023);
and U31750 (N_31750,N_30533,N_30471);
xor U31751 (N_31751,N_30370,N_30230);
nor U31752 (N_31752,N_30161,N_30119);
nand U31753 (N_31753,N_30817,N_30215);
nor U31754 (N_31754,N_30924,N_30562);
xnor U31755 (N_31755,N_30263,N_30040);
and U31756 (N_31756,N_30908,N_30744);
or U31757 (N_31757,N_30862,N_30949);
nor U31758 (N_31758,N_30209,N_30333);
nand U31759 (N_31759,N_30775,N_30065);
nand U31760 (N_31760,N_30084,N_30651);
xor U31761 (N_31761,N_30233,N_30505);
nor U31762 (N_31762,N_30639,N_30287);
and U31763 (N_31763,N_30399,N_30430);
xor U31764 (N_31764,N_30760,N_30005);
xnor U31765 (N_31765,N_30523,N_30073);
xnor U31766 (N_31766,N_30946,N_30832);
nand U31767 (N_31767,N_30133,N_30050);
nand U31768 (N_31768,N_30373,N_30799);
nor U31769 (N_31769,N_30047,N_30257);
nor U31770 (N_31770,N_30258,N_30419);
or U31771 (N_31771,N_30863,N_30669);
or U31772 (N_31772,N_30634,N_30037);
or U31773 (N_31773,N_30891,N_30657);
nor U31774 (N_31774,N_30326,N_30434);
nor U31775 (N_31775,N_30081,N_30494);
nor U31776 (N_31776,N_30925,N_30483);
or U31777 (N_31777,N_30869,N_30196);
nand U31778 (N_31778,N_30415,N_30234);
nor U31779 (N_31779,N_30399,N_30988);
nand U31780 (N_31780,N_30329,N_30299);
nor U31781 (N_31781,N_30034,N_30524);
xnor U31782 (N_31782,N_30474,N_30641);
nand U31783 (N_31783,N_30989,N_30410);
or U31784 (N_31784,N_30342,N_30754);
xor U31785 (N_31785,N_30459,N_30129);
and U31786 (N_31786,N_30393,N_30291);
or U31787 (N_31787,N_30854,N_30891);
nor U31788 (N_31788,N_30616,N_30401);
nor U31789 (N_31789,N_30060,N_30792);
nor U31790 (N_31790,N_30839,N_30043);
nor U31791 (N_31791,N_30631,N_30842);
nand U31792 (N_31792,N_30287,N_30199);
xor U31793 (N_31793,N_30215,N_30708);
and U31794 (N_31794,N_30701,N_30307);
nand U31795 (N_31795,N_30429,N_30942);
nand U31796 (N_31796,N_30956,N_30840);
and U31797 (N_31797,N_30076,N_30109);
nand U31798 (N_31798,N_30141,N_30876);
xnor U31799 (N_31799,N_30360,N_30180);
or U31800 (N_31800,N_30029,N_30706);
nor U31801 (N_31801,N_30499,N_30541);
nor U31802 (N_31802,N_30362,N_30335);
nor U31803 (N_31803,N_30853,N_30805);
or U31804 (N_31804,N_30987,N_30881);
nor U31805 (N_31805,N_30548,N_30034);
or U31806 (N_31806,N_30385,N_30486);
nor U31807 (N_31807,N_30082,N_30262);
and U31808 (N_31808,N_30940,N_30038);
or U31809 (N_31809,N_30569,N_30472);
and U31810 (N_31810,N_30062,N_30918);
nor U31811 (N_31811,N_30995,N_30060);
nor U31812 (N_31812,N_30809,N_30460);
nand U31813 (N_31813,N_30469,N_30605);
nor U31814 (N_31814,N_30037,N_30642);
nand U31815 (N_31815,N_30325,N_30981);
and U31816 (N_31816,N_30884,N_30420);
nand U31817 (N_31817,N_30181,N_30153);
xor U31818 (N_31818,N_30557,N_30028);
xnor U31819 (N_31819,N_30190,N_30284);
and U31820 (N_31820,N_30198,N_30036);
and U31821 (N_31821,N_30464,N_30245);
nor U31822 (N_31822,N_30051,N_30058);
nand U31823 (N_31823,N_30812,N_30154);
xnor U31824 (N_31824,N_30611,N_30360);
nor U31825 (N_31825,N_30454,N_30782);
or U31826 (N_31826,N_30996,N_30300);
nand U31827 (N_31827,N_30010,N_30480);
or U31828 (N_31828,N_30988,N_30822);
and U31829 (N_31829,N_30117,N_30661);
nor U31830 (N_31830,N_30382,N_30740);
xor U31831 (N_31831,N_30169,N_30081);
nor U31832 (N_31832,N_30946,N_30834);
nor U31833 (N_31833,N_30219,N_30387);
and U31834 (N_31834,N_30841,N_30491);
nand U31835 (N_31835,N_30276,N_30472);
or U31836 (N_31836,N_30474,N_30192);
xor U31837 (N_31837,N_30704,N_30490);
and U31838 (N_31838,N_30682,N_30175);
and U31839 (N_31839,N_30938,N_30355);
nor U31840 (N_31840,N_30306,N_30502);
xnor U31841 (N_31841,N_30010,N_30813);
and U31842 (N_31842,N_30601,N_30137);
or U31843 (N_31843,N_30170,N_30240);
nand U31844 (N_31844,N_30980,N_30263);
xor U31845 (N_31845,N_30679,N_30440);
and U31846 (N_31846,N_30758,N_30073);
xor U31847 (N_31847,N_30523,N_30810);
nand U31848 (N_31848,N_30776,N_30725);
xnor U31849 (N_31849,N_30561,N_30245);
nor U31850 (N_31850,N_30899,N_30999);
nand U31851 (N_31851,N_30784,N_30488);
and U31852 (N_31852,N_30567,N_30225);
xnor U31853 (N_31853,N_30251,N_30049);
xnor U31854 (N_31854,N_30527,N_30889);
and U31855 (N_31855,N_30494,N_30967);
and U31856 (N_31856,N_30526,N_30737);
nor U31857 (N_31857,N_30867,N_30687);
or U31858 (N_31858,N_30874,N_30268);
or U31859 (N_31859,N_30914,N_30631);
xor U31860 (N_31860,N_30959,N_30030);
nor U31861 (N_31861,N_30272,N_30796);
or U31862 (N_31862,N_30193,N_30705);
and U31863 (N_31863,N_30234,N_30012);
xnor U31864 (N_31864,N_30547,N_30346);
and U31865 (N_31865,N_30501,N_30751);
and U31866 (N_31866,N_30251,N_30288);
or U31867 (N_31867,N_30918,N_30277);
nand U31868 (N_31868,N_30923,N_30233);
and U31869 (N_31869,N_30089,N_30963);
and U31870 (N_31870,N_30581,N_30535);
nor U31871 (N_31871,N_30442,N_30593);
xnor U31872 (N_31872,N_30151,N_30616);
nor U31873 (N_31873,N_30479,N_30914);
xor U31874 (N_31874,N_30768,N_30573);
and U31875 (N_31875,N_30323,N_30325);
xnor U31876 (N_31876,N_30618,N_30883);
and U31877 (N_31877,N_30736,N_30261);
and U31878 (N_31878,N_30457,N_30374);
nor U31879 (N_31879,N_30414,N_30907);
nor U31880 (N_31880,N_30674,N_30350);
nor U31881 (N_31881,N_30660,N_30938);
or U31882 (N_31882,N_30638,N_30944);
xor U31883 (N_31883,N_30218,N_30787);
nor U31884 (N_31884,N_30015,N_30257);
and U31885 (N_31885,N_30638,N_30322);
nand U31886 (N_31886,N_30100,N_30582);
nor U31887 (N_31887,N_30640,N_30060);
and U31888 (N_31888,N_30121,N_30146);
and U31889 (N_31889,N_30634,N_30496);
and U31890 (N_31890,N_30701,N_30204);
nor U31891 (N_31891,N_30050,N_30209);
nor U31892 (N_31892,N_30416,N_30055);
xnor U31893 (N_31893,N_30441,N_30910);
xor U31894 (N_31894,N_30916,N_30021);
nor U31895 (N_31895,N_30490,N_30501);
or U31896 (N_31896,N_30126,N_30908);
xnor U31897 (N_31897,N_30084,N_30937);
and U31898 (N_31898,N_30447,N_30180);
xor U31899 (N_31899,N_30060,N_30018);
xnor U31900 (N_31900,N_30589,N_30445);
nand U31901 (N_31901,N_30146,N_30442);
nor U31902 (N_31902,N_30294,N_30052);
and U31903 (N_31903,N_30987,N_30527);
xor U31904 (N_31904,N_30974,N_30855);
nand U31905 (N_31905,N_30496,N_30068);
nand U31906 (N_31906,N_30242,N_30769);
nor U31907 (N_31907,N_30591,N_30794);
and U31908 (N_31908,N_30577,N_30184);
nand U31909 (N_31909,N_30846,N_30729);
xor U31910 (N_31910,N_30519,N_30336);
nand U31911 (N_31911,N_30142,N_30126);
xor U31912 (N_31912,N_30565,N_30314);
nand U31913 (N_31913,N_30920,N_30939);
or U31914 (N_31914,N_30430,N_30891);
and U31915 (N_31915,N_30998,N_30188);
and U31916 (N_31916,N_30679,N_30008);
and U31917 (N_31917,N_30781,N_30560);
nand U31918 (N_31918,N_30189,N_30951);
xor U31919 (N_31919,N_30302,N_30411);
xor U31920 (N_31920,N_30209,N_30835);
xnor U31921 (N_31921,N_30857,N_30192);
nand U31922 (N_31922,N_30699,N_30450);
xor U31923 (N_31923,N_30297,N_30303);
nor U31924 (N_31924,N_30027,N_30471);
xnor U31925 (N_31925,N_30608,N_30267);
xor U31926 (N_31926,N_30752,N_30517);
and U31927 (N_31927,N_30199,N_30782);
nor U31928 (N_31928,N_30273,N_30264);
xnor U31929 (N_31929,N_30580,N_30120);
and U31930 (N_31930,N_30271,N_30895);
and U31931 (N_31931,N_30953,N_30708);
nand U31932 (N_31932,N_30118,N_30229);
nor U31933 (N_31933,N_30781,N_30463);
nand U31934 (N_31934,N_30743,N_30592);
nor U31935 (N_31935,N_30196,N_30688);
nand U31936 (N_31936,N_30549,N_30444);
and U31937 (N_31937,N_30420,N_30301);
nor U31938 (N_31938,N_30137,N_30889);
xor U31939 (N_31939,N_30207,N_30887);
xor U31940 (N_31940,N_30768,N_30230);
nor U31941 (N_31941,N_30131,N_30960);
and U31942 (N_31942,N_30514,N_30658);
or U31943 (N_31943,N_30053,N_30778);
nand U31944 (N_31944,N_30062,N_30895);
and U31945 (N_31945,N_30810,N_30206);
or U31946 (N_31946,N_30142,N_30305);
nor U31947 (N_31947,N_30348,N_30906);
xor U31948 (N_31948,N_30225,N_30460);
and U31949 (N_31949,N_30767,N_30546);
and U31950 (N_31950,N_30009,N_30044);
and U31951 (N_31951,N_30202,N_30049);
nand U31952 (N_31952,N_30631,N_30708);
or U31953 (N_31953,N_30575,N_30206);
nor U31954 (N_31954,N_30611,N_30448);
xnor U31955 (N_31955,N_30427,N_30117);
and U31956 (N_31956,N_30436,N_30407);
nand U31957 (N_31957,N_30651,N_30955);
nand U31958 (N_31958,N_30779,N_30894);
or U31959 (N_31959,N_30619,N_30206);
nor U31960 (N_31960,N_30164,N_30735);
nor U31961 (N_31961,N_30010,N_30360);
xnor U31962 (N_31962,N_30877,N_30906);
nand U31963 (N_31963,N_30794,N_30238);
or U31964 (N_31964,N_30157,N_30907);
and U31965 (N_31965,N_30114,N_30389);
nor U31966 (N_31966,N_30276,N_30285);
or U31967 (N_31967,N_30925,N_30437);
nand U31968 (N_31968,N_30950,N_30003);
and U31969 (N_31969,N_30646,N_30318);
nor U31970 (N_31970,N_30598,N_30377);
and U31971 (N_31971,N_30435,N_30324);
nor U31972 (N_31972,N_30350,N_30528);
xnor U31973 (N_31973,N_30863,N_30856);
xnor U31974 (N_31974,N_30883,N_30367);
nor U31975 (N_31975,N_30186,N_30576);
or U31976 (N_31976,N_30930,N_30778);
and U31977 (N_31977,N_30501,N_30421);
nor U31978 (N_31978,N_30913,N_30888);
and U31979 (N_31979,N_30658,N_30524);
nand U31980 (N_31980,N_30602,N_30451);
xnor U31981 (N_31981,N_30577,N_30121);
nand U31982 (N_31982,N_30451,N_30685);
and U31983 (N_31983,N_30161,N_30429);
nand U31984 (N_31984,N_30675,N_30462);
nor U31985 (N_31985,N_30150,N_30374);
and U31986 (N_31986,N_30855,N_30636);
nor U31987 (N_31987,N_30520,N_30684);
nor U31988 (N_31988,N_30725,N_30964);
xor U31989 (N_31989,N_30800,N_30458);
xor U31990 (N_31990,N_30341,N_30272);
and U31991 (N_31991,N_30554,N_30968);
xnor U31992 (N_31992,N_30179,N_30047);
and U31993 (N_31993,N_30857,N_30172);
nor U31994 (N_31994,N_30618,N_30085);
or U31995 (N_31995,N_30971,N_30146);
nor U31996 (N_31996,N_30440,N_30960);
xnor U31997 (N_31997,N_30035,N_30180);
nor U31998 (N_31998,N_30420,N_30810);
nor U31999 (N_31999,N_30704,N_30831);
nor U32000 (N_32000,N_31554,N_31148);
xor U32001 (N_32001,N_31671,N_31439);
nor U32002 (N_32002,N_31212,N_31121);
or U32003 (N_32003,N_31060,N_31521);
and U32004 (N_32004,N_31483,N_31039);
or U32005 (N_32005,N_31442,N_31835);
or U32006 (N_32006,N_31926,N_31870);
xor U32007 (N_32007,N_31820,N_31793);
xnor U32008 (N_32008,N_31074,N_31110);
nand U32009 (N_32009,N_31508,N_31139);
and U32010 (N_32010,N_31706,N_31791);
xor U32011 (N_32011,N_31731,N_31070);
nor U32012 (N_32012,N_31654,N_31075);
nand U32013 (N_32013,N_31268,N_31659);
nand U32014 (N_32014,N_31510,N_31799);
or U32015 (N_32015,N_31974,N_31366);
or U32016 (N_32016,N_31548,N_31657);
nor U32017 (N_32017,N_31157,N_31445);
or U32018 (N_32018,N_31704,N_31381);
nand U32019 (N_32019,N_31936,N_31197);
nor U32020 (N_32020,N_31584,N_31296);
or U32021 (N_32021,N_31363,N_31574);
and U32022 (N_32022,N_31913,N_31173);
xnor U32023 (N_32023,N_31095,N_31355);
and U32024 (N_32024,N_31246,N_31801);
nor U32025 (N_32025,N_31899,N_31956);
nand U32026 (N_32026,N_31502,N_31608);
nor U32027 (N_32027,N_31871,N_31617);
or U32028 (N_32028,N_31973,N_31347);
or U32029 (N_32029,N_31580,N_31317);
or U32030 (N_32030,N_31934,N_31995);
xnor U32031 (N_32031,N_31542,N_31778);
or U32032 (N_32032,N_31632,N_31901);
nor U32033 (N_32033,N_31134,N_31307);
xor U32034 (N_32034,N_31045,N_31655);
nand U32035 (N_32035,N_31985,N_31408);
xnor U32036 (N_32036,N_31484,N_31619);
and U32037 (N_32037,N_31325,N_31822);
nor U32038 (N_32038,N_31456,N_31509);
nand U32039 (N_32039,N_31145,N_31981);
or U32040 (N_32040,N_31334,N_31297);
nor U32041 (N_32041,N_31749,N_31775);
nor U32042 (N_32042,N_31519,N_31006);
or U32043 (N_32043,N_31499,N_31993);
nor U32044 (N_32044,N_31462,N_31579);
nor U32045 (N_32045,N_31433,N_31191);
nor U32046 (N_32046,N_31876,N_31222);
nand U32047 (N_32047,N_31189,N_31768);
nand U32048 (N_32048,N_31021,N_31549);
and U32049 (N_32049,N_31674,N_31787);
nand U32050 (N_32050,N_31625,N_31373);
or U32051 (N_32051,N_31624,N_31398);
or U32052 (N_32052,N_31898,N_31160);
nor U32053 (N_32053,N_31961,N_31728);
or U32054 (N_32054,N_31477,N_31903);
and U32055 (N_32055,N_31798,N_31088);
nand U32056 (N_32056,N_31566,N_31261);
and U32057 (N_32057,N_31658,N_31496);
xnor U32058 (N_32058,N_31220,N_31991);
and U32059 (N_32059,N_31829,N_31165);
and U32060 (N_32060,N_31466,N_31938);
xnor U32061 (N_32061,N_31194,N_31323);
nor U32062 (N_32062,N_31602,N_31495);
nand U32063 (N_32063,N_31953,N_31567);
nor U32064 (N_32064,N_31747,N_31353);
and U32065 (N_32065,N_31278,N_31065);
xor U32066 (N_32066,N_31845,N_31356);
or U32067 (N_32067,N_31911,N_31879);
or U32068 (N_32068,N_31957,N_31281);
nor U32069 (N_32069,N_31622,N_31629);
xor U32070 (N_32070,N_31645,N_31885);
or U32071 (N_32071,N_31818,N_31744);
nand U32072 (N_32072,N_31977,N_31169);
nor U32073 (N_32073,N_31526,N_31666);
or U32074 (N_32074,N_31858,N_31722);
nand U32075 (N_32075,N_31630,N_31716);
nor U32076 (N_32076,N_31192,N_31767);
nand U32077 (N_32077,N_31950,N_31792);
xnor U32078 (N_32078,N_31403,N_31515);
xor U32079 (N_32079,N_31342,N_31422);
or U32080 (N_32080,N_31664,N_31505);
nand U32081 (N_32081,N_31853,N_31796);
and U32082 (N_32082,N_31201,N_31850);
nor U32083 (N_32083,N_31258,N_31400);
xnor U32084 (N_32084,N_31419,N_31746);
nand U32085 (N_32085,N_31489,N_31073);
xor U32086 (N_32086,N_31589,N_31770);
nand U32087 (N_32087,N_31545,N_31046);
xnor U32088 (N_32088,N_31223,N_31717);
xnor U32089 (N_32089,N_31676,N_31406);
and U32090 (N_32090,N_31457,N_31942);
xnor U32091 (N_32091,N_31507,N_31378);
nor U32092 (N_32092,N_31198,N_31030);
xnor U32093 (N_32093,N_31104,N_31399);
nor U32094 (N_32094,N_31735,N_31849);
or U32095 (N_32095,N_31014,N_31018);
or U32096 (N_32096,N_31841,N_31971);
nor U32097 (N_32097,N_31817,N_31960);
nand U32098 (N_32098,N_31809,N_31975);
nand U32099 (N_32099,N_31079,N_31581);
nand U32100 (N_32100,N_31464,N_31182);
and U32101 (N_32101,N_31232,N_31970);
or U32102 (N_32102,N_31937,N_31874);
or U32103 (N_32103,N_31183,N_31056);
and U32104 (N_32104,N_31748,N_31054);
nand U32105 (N_32105,N_31390,N_31168);
nand U32106 (N_32106,N_31072,N_31648);
nand U32107 (N_32107,N_31551,N_31776);
and U32108 (N_32108,N_31873,N_31636);
nor U32109 (N_32109,N_31618,N_31029);
and U32110 (N_32110,N_31115,N_31958);
or U32111 (N_32111,N_31783,N_31553);
nand U32112 (N_32112,N_31446,N_31328);
nor U32113 (N_32113,N_31651,N_31550);
or U32114 (N_32114,N_31641,N_31572);
and U32115 (N_32115,N_31158,N_31431);
nor U32116 (N_32116,N_31091,N_31867);
nor U32117 (N_32117,N_31569,N_31245);
and U32118 (N_32118,N_31781,N_31605);
xor U32119 (N_32119,N_31239,N_31837);
or U32120 (N_32120,N_31085,N_31314);
nand U32121 (N_32121,N_31467,N_31090);
nand U32122 (N_32122,N_31919,N_31335);
or U32123 (N_32123,N_31393,N_31276);
or U32124 (N_32124,N_31537,N_31935);
or U32125 (N_32125,N_31760,N_31807);
nand U32126 (N_32126,N_31059,N_31785);
nand U32127 (N_32127,N_31329,N_31238);
nor U32128 (N_32128,N_31080,N_31256);
and U32129 (N_32129,N_31391,N_31247);
or U32130 (N_32130,N_31711,N_31005);
nor U32131 (N_32131,N_31585,N_31897);
and U32132 (N_32132,N_31471,N_31894);
nand U32133 (N_32133,N_31772,N_31988);
or U32134 (N_32134,N_31282,N_31561);
and U32135 (N_32135,N_31862,N_31650);
nor U32136 (N_32136,N_31214,N_31343);
and U32137 (N_32137,N_31250,N_31371);
nand U32138 (N_32138,N_31848,N_31416);
and U32139 (N_32139,N_31494,N_31927);
nor U32140 (N_32140,N_31843,N_31933);
or U32141 (N_32141,N_31100,N_31774);
or U32142 (N_32142,N_31609,N_31719);
nor U32143 (N_32143,N_31293,N_31233);
nor U32144 (N_32144,N_31790,N_31939);
nor U32145 (N_32145,N_31610,N_31538);
nor U32146 (N_32146,N_31432,N_31915);
and U32147 (N_32147,N_31407,N_31291);
nor U32148 (N_32148,N_31252,N_31861);
xor U32149 (N_32149,N_31844,N_31362);
nand U32150 (N_32150,N_31628,N_31924);
xnor U32151 (N_32151,N_31725,N_31009);
or U32152 (N_32152,N_31751,N_31230);
and U32153 (N_32153,N_31583,N_31076);
or U32154 (N_32154,N_31642,N_31779);
nor U32155 (N_32155,N_31701,N_31083);
or U32156 (N_32156,N_31132,N_31156);
or U32157 (N_32157,N_31318,N_31374);
and U32158 (N_32158,N_31063,N_31591);
and U32159 (N_32159,N_31576,N_31922);
nor U32160 (N_32160,N_31965,N_31200);
nor U32161 (N_32161,N_31210,N_31405);
and U32162 (N_32162,N_31396,N_31249);
nor U32163 (N_32163,N_31154,N_31721);
nor U32164 (N_32164,N_31336,N_31368);
nor U32165 (N_32165,N_31708,N_31959);
nand U32166 (N_32166,N_31058,N_31892);
and U32167 (N_32167,N_31162,N_31627);
nand U32168 (N_32168,N_31951,N_31454);
nor U32169 (N_32169,N_31524,N_31102);
nor U32170 (N_32170,N_31663,N_31500);
nand U32171 (N_32171,N_31487,N_31773);
nand U32172 (N_32172,N_31043,N_31444);
nand U32173 (N_32173,N_31027,N_31479);
xor U32174 (N_32174,N_31308,N_31527);
or U32175 (N_32175,N_31022,N_31225);
and U32176 (N_32176,N_31730,N_31235);
and U32177 (N_32177,N_31350,N_31469);
or U32178 (N_32178,N_31380,N_31559);
and U32179 (N_32179,N_31228,N_31440);
xor U32180 (N_32180,N_31516,N_31705);
nor U32181 (N_32181,N_31434,N_31904);
or U32182 (N_32182,N_31920,N_31122);
or U32183 (N_32183,N_31601,N_31888);
and U32184 (N_32184,N_31383,N_31755);
xor U32185 (N_32185,N_31866,N_31679);
nand U32186 (N_32186,N_31036,N_31137);
xnor U32187 (N_32187,N_31007,N_31288);
nand U32188 (N_32188,N_31427,N_31682);
nand U32189 (N_32189,N_31259,N_31199);
nand U32190 (N_32190,N_31541,N_31805);
xor U32191 (N_32191,N_31757,N_31370);
nor U32192 (N_32192,N_31680,N_31195);
and U32193 (N_32193,N_31093,N_31397);
nor U32194 (N_32194,N_31204,N_31667);
xor U32195 (N_32195,N_31797,N_31944);
nand U32196 (N_32196,N_31086,N_31529);
nand U32197 (N_32197,N_31825,N_31114);
or U32198 (N_32198,N_31333,N_31734);
or U32199 (N_32199,N_31877,N_31826);
xor U32200 (N_32200,N_31236,N_31568);
nor U32201 (N_32201,N_31603,N_31864);
nor U32202 (N_32202,N_31759,N_31423);
xor U32203 (N_32203,N_31890,N_31522);
and U32204 (N_32204,N_31571,N_31340);
nand U32205 (N_32205,N_31119,N_31414);
nand U32206 (N_32206,N_31794,N_31896);
xor U32207 (N_32207,N_31038,N_31593);
nor U32208 (N_32208,N_31016,N_31337);
nand U32209 (N_32209,N_31980,N_31395);
and U32210 (N_32210,N_31543,N_31819);
and U32211 (N_32211,N_31780,N_31763);
and U32212 (N_32212,N_31756,N_31812);
and U32213 (N_32213,N_31109,N_31834);
nand U32214 (N_32214,N_31752,N_31740);
or U32215 (N_32215,N_31525,N_31348);
xnor U32216 (N_32216,N_31164,N_31042);
and U32217 (N_32217,N_31685,N_31856);
nor U32218 (N_32218,N_31695,N_31555);
nand U32219 (N_32219,N_31025,N_31983);
nor U32220 (N_32220,N_31053,N_31242);
nand U32221 (N_32221,N_31263,N_31590);
nand U32222 (N_32222,N_31923,N_31754);
nor U32223 (N_32223,N_31129,N_31905);
xnor U32224 (N_32224,N_31461,N_31426);
nand U32225 (N_32225,N_31670,N_31177);
xnor U32226 (N_32226,N_31392,N_31782);
nand U32227 (N_32227,N_31193,N_31311);
nor U32228 (N_32228,N_31178,N_31997);
nor U32229 (N_32229,N_31112,N_31428);
nand U32230 (N_32230,N_31000,N_31758);
xnor U32231 (N_32231,N_31539,N_31547);
nand U32232 (N_32232,N_31878,N_31324);
and U32233 (N_32233,N_31764,N_31465);
nor U32234 (N_32234,N_31635,N_31217);
nand U32235 (N_32235,N_31305,N_31604);
and U32236 (N_32236,N_31880,N_31170);
xor U32237 (N_32237,N_31240,N_31116);
nand U32238 (N_32238,N_31251,N_31714);
xnor U32239 (N_32239,N_31718,N_31300);
xnor U32240 (N_32240,N_31019,N_31094);
and U32241 (N_32241,N_31669,N_31954);
nand U32242 (N_32242,N_31034,N_31048);
xor U32243 (N_32243,N_31443,N_31715);
nand U32244 (N_32244,N_31587,N_31289);
or U32245 (N_32245,N_31410,N_31626);
xor U32246 (N_32246,N_31552,N_31101);
or U32247 (N_32247,N_31544,N_31498);
or U32248 (N_32248,N_31745,N_31049);
and U32249 (N_32249,N_31556,N_31097);
nand U32250 (N_32250,N_31883,N_31118);
nand U32251 (N_32251,N_31616,N_31430);
nor U32252 (N_32252,N_31710,N_31458);
and U32253 (N_32253,N_31451,N_31437);
or U32254 (N_32254,N_31203,N_31349);
or U32255 (N_32255,N_31441,N_31528);
and U32256 (N_32256,N_31044,N_31720);
or U32257 (N_32257,N_31827,N_31227);
and U32258 (N_32258,N_31033,N_31150);
nand U32259 (N_32259,N_31943,N_31409);
nand U32260 (N_32260,N_31921,N_31388);
and U32261 (N_32261,N_31436,N_31262);
and U32262 (N_32262,N_31788,N_31990);
xnor U32263 (N_32263,N_31292,N_31769);
xnor U32264 (N_32264,N_31023,N_31125);
and U32265 (N_32265,N_31486,N_31771);
and U32266 (N_32266,N_31570,N_31836);
nor U32267 (N_32267,N_31248,N_31175);
nor U32268 (N_32268,N_31514,N_31142);
and U32269 (N_32269,N_31267,N_31532);
nor U32270 (N_32270,N_31099,N_31662);
or U32271 (N_32271,N_31917,N_31703);
nand U32272 (N_32272,N_31215,N_31346);
or U32273 (N_32273,N_31476,N_31017);
or U32274 (N_32274,N_31123,N_31517);
nand U32275 (N_32275,N_31302,N_31345);
nand U32276 (N_32276,N_31481,N_31918);
or U32277 (N_32277,N_31989,N_31106);
nor U32278 (N_32278,N_31810,N_31639);
nor U32279 (N_32279,N_31186,N_31052);
or U32280 (N_32280,N_31316,N_31190);
and U32281 (N_32281,N_31611,N_31096);
and U32282 (N_32282,N_31724,N_31986);
xor U32283 (N_32283,N_31141,N_31916);
or U32284 (N_32284,N_31159,N_31683);
xor U32285 (N_32285,N_31449,N_31886);
or U32286 (N_32286,N_31815,N_31167);
nand U32287 (N_32287,N_31599,N_31932);
xor U32288 (N_32288,N_31146,N_31377);
or U32289 (N_32289,N_31062,N_31723);
or U32290 (N_32290,N_31153,N_31803);
and U32291 (N_32291,N_31729,N_31420);
xor U32292 (N_32292,N_31909,N_31697);
nor U32293 (N_32293,N_31762,N_31813);
or U32294 (N_32294,N_31174,N_31089);
or U32295 (N_32295,N_31415,N_31224);
nor U32296 (N_32296,N_31518,N_31575);
and U32297 (N_32297,N_31806,N_31925);
xnor U32298 (N_32298,N_31357,N_31172);
and U32299 (N_32299,N_31906,N_31784);
nand U32300 (N_32300,N_31875,N_31560);
xor U32301 (N_32301,N_31187,N_31425);
nor U32302 (N_32302,N_31531,N_31131);
nor U32303 (N_32303,N_31071,N_31497);
or U32304 (N_32304,N_31557,N_31107);
or U32305 (N_32305,N_31084,N_31105);
or U32306 (N_32306,N_31057,N_31530);
and U32307 (N_32307,N_31375,N_31802);
xnor U32308 (N_32308,N_31613,N_31741);
and U32309 (N_32309,N_31600,N_31050);
or U32310 (N_32310,N_31637,N_31143);
xor U32311 (N_32311,N_31621,N_31882);
nor U32312 (N_32312,N_31546,N_31984);
nor U32313 (N_32313,N_31020,N_31594);
xnor U32314 (N_32314,N_31087,N_31360);
xnor U32315 (N_32315,N_31313,N_31179);
or U32316 (N_32316,N_31713,N_31586);
nand U32317 (N_32317,N_31511,N_31234);
xor U32318 (N_32318,N_31066,N_31945);
and U32319 (N_32319,N_31631,N_31996);
xnor U32320 (N_32320,N_31155,N_31686);
or U32321 (N_32321,N_31035,N_31068);
nor U32322 (N_32322,N_31492,N_31176);
xnor U32323 (N_32323,N_31438,N_31821);
nand U32324 (N_32324,N_31520,N_31859);
nand U32325 (N_32325,N_31969,N_31298);
and U32326 (N_32326,N_31460,N_31633);
xor U32327 (N_32327,N_31257,N_31588);
nor U32328 (N_32328,N_31816,N_31067);
nand U32329 (N_32329,N_31208,N_31852);
and U32330 (N_32330,N_31237,N_31506);
xnor U32331 (N_32331,N_31144,N_31893);
and U32332 (N_32332,N_31681,N_31978);
or U32333 (N_32333,N_31900,N_31108);
or U32334 (N_32334,N_31055,N_31166);
nand U32335 (N_32335,N_31219,N_31929);
nand U32336 (N_32336,N_31795,N_31128);
and U32337 (N_32337,N_31949,N_31643);
xnor U32338 (N_32338,N_31301,N_31188);
nand U32339 (N_32339,N_31216,N_31254);
and U32340 (N_32340,N_31404,N_31709);
nand U32341 (N_32341,N_31279,N_31895);
xnor U32342 (N_32342,N_31394,N_31808);
nand U32343 (N_32343,N_31003,N_31351);
nand U32344 (N_32344,N_31914,N_31061);
xor U32345 (N_32345,N_31330,N_31478);
nor U32346 (N_32346,N_31450,N_31452);
and U32347 (N_32347,N_31361,N_31800);
or U32348 (N_32348,N_31275,N_31833);
and U32349 (N_32349,N_31868,N_31207);
and U32350 (N_32350,N_31742,N_31688);
nand U32351 (N_32351,N_31750,N_31504);
xor U32352 (N_32352,N_31647,N_31002);
nor U32353 (N_32353,N_31948,N_31766);
xnor U32354 (N_32354,N_31320,N_31967);
and U32355 (N_32355,N_31623,N_31928);
nor U32356 (N_32356,N_31202,N_31592);
nand U32357 (N_32357,N_31290,N_31952);
nor U32358 (N_32358,N_31184,N_31309);
and U32359 (N_32359,N_31832,N_31907);
and U32360 (N_32360,N_31678,N_31359);
nor U32361 (N_32361,N_31424,N_31732);
nor U32362 (N_32362,N_31272,N_31789);
or U32363 (N_32363,N_31999,N_31015);
nor U32364 (N_32364,N_31205,N_31577);
and U32365 (N_32365,N_31855,N_31133);
and U32366 (N_32366,N_31135,N_31596);
nor U32367 (N_32367,N_31041,N_31693);
xor U32368 (N_32368,N_31607,N_31998);
and U32369 (N_32369,N_31563,N_31372);
nand U32370 (N_32370,N_31321,N_31270);
nand U32371 (N_32371,N_31113,N_31653);
and U32372 (N_32372,N_31830,N_31684);
nand U32373 (N_32373,N_31804,N_31260);
xnor U32374 (N_32374,N_31031,N_31331);
nand U32375 (N_32375,N_31051,N_31738);
xor U32376 (N_32376,N_31299,N_31354);
or U32377 (N_32377,N_31266,N_31384);
nor U32378 (N_32378,N_31947,N_31699);
nand U32379 (N_32379,N_31908,N_31429);
and U32380 (N_32380,N_31614,N_31612);
nor U32381 (N_32381,N_31700,N_31672);
or U32382 (N_32382,N_31698,N_31660);
and U32383 (N_32383,N_31620,N_31493);
or U32384 (N_32384,N_31946,N_31727);
nor U32385 (N_32385,N_31872,N_31863);
xor U32386 (N_32386,N_31582,N_31448);
nor U32387 (N_32387,N_31402,N_31064);
and U32388 (N_32388,N_31823,N_31828);
xor U32389 (N_32389,N_31455,N_31306);
nor U32390 (N_32390,N_31136,N_31365);
nand U32391 (N_32391,N_31712,N_31312);
and U32392 (N_32392,N_31691,N_31902);
nand U32393 (N_32393,N_31972,N_31702);
nand U32394 (N_32394,N_31024,N_31344);
nor U32395 (N_32395,N_31512,N_31421);
and U32396 (N_32396,N_31675,N_31474);
xor U32397 (N_32397,N_31982,N_31130);
or U32398 (N_32398,N_31447,N_31338);
xor U32399 (N_32399,N_31111,N_31124);
xor U32400 (N_32400,N_31147,N_31941);
or U32401 (N_32401,N_31367,N_31847);
and U32402 (N_32402,N_31271,N_31860);
or U32403 (N_32403,N_31523,N_31322);
or U32404 (N_32404,N_31418,N_31595);
xnor U32405 (N_32405,N_31001,N_31689);
and U32406 (N_32406,N_31968,N_31814);
or U32407 (N_32407,N_31839,N_31824);
or U32408 (N_32408,N_31226,N_31533);
nand U32409 (N_32409,N_31707,N_31152);
nand U32410 (N_32410,N_31211,N_31196);
xnor U32411 (N_32411,N_31319,N_31930);
or U32412 (N_32412,N_31857,N_31846);
nand U32413 (N_32413,N_31010,N_31138);
xor U32414 (N_32414,N_31077,N_31218);
xor U32415 (N_32415,N_31501,N_31185);
xnor U32416 (N_32416,N_31206,N_31221);
xor U32417 (N_32417,N_31026,N_31241);
and U32418 (N_32418,N_31668,N_31181);
nand U32419 (N_32419,N_31475,N_31253);
nand U32420 (N_32420,N_31976,N_31482);
nand U32421 (N_32421,N_31283,N_31078);
xnor U32422 (N_32422,N_31120,N_31103);
nor U32423 (N_32423,N_31480,N_31535);
xor U32424 (N_32424,N_31327,N_31865);
nor U32425 (N_32425,N_31284,N_31578);
and U32426 (N_32426,N_31013,N_31274);
nor U32427 (N_32427,N_31032,N_31811);
nand U32428 (N_32428,N_31652,N_31485);
nand U32429 (N_32429,N_31411,N_31994);
and U32430 (N_32430,N_31412,N_31273);
nor U32431 (N_32431,N_31739,N_31040);
nor U32432 (N_32432,N_31352,N_31513);
xor U32433 (N_32433,N_31294,N_31286);
xnor U32434 (N_32434,N_31092,N_31687);
nor U32435 (N_32435,N_31149,N_31962);
or U32436 (N_32436,N_31401,N_31955);
nand U32437 (N_32437,N_31726,N_31161);
and U32438 (N_32438,N_31037,N_31615);
or U32439 (N_32439,N_31417,N_31231);
and U32440 (N_32440,N_31332,N_31376);
xnor U32441 (N_32441,N_31364,N_31851);
nor U32442 (N_32442,N_31656,N_31606);
or U32443 (N_32443,N_31004,N_31598);
xnor U32444 (N_32444,N_31468,N_31534);
or U32445 (N_32445,N_31761,N_31387);
and U32446 (N_32446,N_31536,N_31011);
nor U32447 (N_32447,N_31151,N_31126);
nor U32448 (N_32448,N_31069,N_31470);
xnor U32449 (N_32449,N_31127,N_31966);
nand U32450 (N_32450,N_31081,N_31047);
nand U32451 (N_32451,N_31646,N_31887);
nand U32452 (N_32452,N_31379,N_31082);
and U32453 (N_32453,N_31987,N_31884);
nand U32454 (N_32454,N_31008,N_31665);
xor U32455 (N_32455,N_31171,N_31453);
and U32456 (N_32456,N_31558,N_31640);
or U32457 (N_32457,N_31940,N_31389);
nor U32458 (N_32458,N_31565,N_31304);
and U32459 (N_32459,N_31473,N_31341);
nand U32460 (N_32460,N_31840,N_31597);
nand U32461 (N_32461,N_31677,N_31265);
nor U32462 (N_32462,N_31694,N_31491);
or U32463 (N_32463,N_31117,N_31315);
or U32464 (N_32464,N_31891,N_31280);
and U32465 (N_32465,N_31842,N_31910);
nand U32466 (N_32466,N_31562,N_31488);
nand U32467 (N_32467,N_31358,N_31326);
or U32468 (N_32468,N_31303,N_31255);
or U32469 (N_32469,N_31503,N_31564);
and U32470 (N_32470,N_31012,N_31382);
xnor U32471 (N_32471,N_31435,N_31765);
or U32472 (N_32472,N_31854,N_31733);
xor U32473 (N_32473,N_31912,N_31737);
nand U32474 (N_32474,N_31696,N_31209);
xor U32475 (N_32475,N_31869,N_31964);
nor U32476 (N_32476,N_31838,N_31992);
xor U32477 (N_32477,N_31786,N_31673);
nor U32478 (N_32478,N_31472,N_31889);
or U32479 (N_32479,N_31213,N_31269);
or U32480 (N_32480,N_31229,N_31459);
nor U32481 (N_32481,N_31413,N_31638);
xor U32482 (N_32482,N_31692,N_31634);
nor U32483 (N_32483,N_31277,N_31180);
nor U32484 (N_32484,N_31385,N_31963);
nor U32485 (N_32485,N_31386,N_31649);
nor U32486 (N_32486,N_31369,N_31573);
nor U32487 (N_32487,N_31244,N_31881);
and U32488 (N_32488,N_31661,N_31285);
nand U32489 (N_32489,N_31463,N_31295);
nand U32490 (N_32490,N_31979,N_31490);
and U32491 (N_32491,N_31140,N_31098);
and U32492 (N_32492,N_31690,N_31028);
nor U32493 (N_32493,N_31753,N_31264);
or U32494 (N_32494,N_31777,N_31831);
xnor U32495 (N_32495,N_31163,N_31339);
nand U32496 (N_32496,N_31310,N_31243);
and U32497 (N_32497,N_31644,N_31287);
or U32498 (N_32498,N_31736,N_31540);
xor U32499 (N_32499,N_31743,N_31931);
nand U32500 (N_32500,N_31851,N_31839);
xnor U32501 (N_32501,N_31237,N_31650);
nand U32502 (N_32502,N_31628,N_31563);
nor U32503 (N_32503,N_31709,N_31507);
or U32504 (N_32504,N_31711,N_31228);
nor U32505 (N_32505,N_31671,N_31229);
xnor U32506 (N_32506,N_31524,N_31527);
nand U32507 (N_32507,N_31211,N_31784);
or U32508 (N_32508,N_31854,N_31350);
nand U32509 (N_32509,N_31886,N_31551);
xor U32510 (N_32510,N_31954,N_31324);
xnor U32511 (N_32511,N_31686,N_31365);
nand U32512 (N_32512,N_31082,N_31182);
nor U32513 (N_32513,N_31074,N_31196);
or U32514 (N_32514,N_31520,N_31288);
and U32515 (N_32515,N_31716,N_31480);
and U32516 (N_32516,N_31067,N_31068);
and U32517 (N_32517,N_31768,N_31466);
or U32518 (N_32518,N_31889,N_31425);
nor U32519 (N_32519,N_31422,N_31839);
or U32520 (N_32520,N_31633,N_31628);
xor U32521 (N_32521,N_31374,N_31517);
or U32522 (N_32522,N_31486,N_31767);
and U32523 (N_32523,N_31333,N_31699);
nor U32524 (N_32524,N_31988,N_31285);
nand U32525 (N_32525,N_31943,N_31933);
nand U32526 (N_32526,N_31613,N_31965);
xnor U32527 (N_32527,N_31313,N_31443);
or U32528 (N_32528,N_31418,N_31727);
xnor U32529 (N_32529,N_31194,N_31341);
and U32530 (N_32530,N_31881,N_31488);
or U32531 (N_32531,N_31323,N_31006);
nand U32532 (N_32532,N_31139,N_31803);
xor U32533 (N_32533,N_31689,N_31987);
xor U32534 (N_32534,N_31870,N_31548);
nand U32535 (N_32535,N_31175,N_31445);
nor U32536 (N_32536,N_31676,N_31680);
and U32537 (N_32537,N_31356,N_31727);
nor U32538 (N_32538,N_31680,N_31233);
nor U32539 (N_32539,N_31244,N_31369);
nor U32540 (N_32540,N_31943,N_31771);
or U32541 (N_32541,N_31552,N_31933);
xor U32542 (N_32542,N_31085,N_31657);
nor U32543 (N_32543,N_31927,N_31072);
and U32544 (N_32544,N_31541,N_31316);
and U32545 (N_32545,N_31764,N_31538);
or U32546 (N_32546,N_31339,N_31138);
nand U32547 (N_32547,N_31926,N_31620);
and U32548 (N_32548,N_31415,N_31340);
or U32549 (N_32549,N_31075,N_31769);
and U32550 (N_32550,N_31299,N_31558);
nor U32551 (N_32551,N_31927,N_31002);
or U32552 (N_32552,N_31542,N_31674);
nor U32553 (N_32553,N_31750,N_31169);
and U32554 (N_32554,N_31314,N_31862);
xnor U32555 (N_32555,N_31536,N_31062);
or U32556 (N_32556,N_31124,N_31485);
and U32557 (N_32557,N_31336,N_31976);
nand U32558 (N_32558,N_31775,N_31289);
nand U32559 (N_32559,N_31534,N_31499);
and U32560 (N_32560,N_31080,N_31500);
nor U32561 (N_32561,N_31154,N_31507);
and U32562 (N_32562,N_31225,N_31984);
nor U32563 (N_32563,N_31245,N_31797);
or U32564 (N_32564,N_31316,N_31092);
or U32565 (N_32565,N_31570,N_31553);
or U32566 (N_32566,N_31988,N_31327);
nor U32567 (N_32567,N_31683,N_31235);
and U32568 (N_32568,N_31980,N_31463);
nand U32569 (N_32569,N_31769,N_31007);
and U32570 (N_32570,N_31708,N_31473);
and U32571 (N_32571,N_31425,N_31342);
nand U32572 (N_32572,N_31926,N_31764);
or U32573 (N_32573,N_31861,N_31391);
nor U32574 (N_32574,N_31847,N_31858);
nor U32575 (N_32575,N_31857,N_31576);
nor U32576 (N_32576,N_31219,N_31785);
xnor U32577 (N_32577,N_31216,N_31928);
nand U32578 (N_32578,N_31891,N_31819);
nand U32579 (N_32579,N_31649,N_31973);
xnor U32580 (N_32580,N_31273,N_31215);
nand U32581 (N_32581,N_31067,N_31420);
nor U32582 (N_32582,N_31486,N_31170);
and U32583 (N_32583,N_31378,N_31616);
nor U32584 (N_32584,N_31732,N_31952);
or U32585 (N_32585,N_31994,N_31613);
nor U32586 (N_32586,N_31395,N_31425);
and U32587 (N_32587,N_31985,N_31523);
xnor U32588 (N_32588,N_31147,N_31389);
nand U32589 (N_32589,N_31203,N_31828);
or U32590 (N_32590,N_31051,N_31670);
nor U32591 (N_32591,N_31302,N_31387);
nor U32592 (N_32592,N_31706,N_31426);
or U32593 (N_32593,N_31895,N_31304);
nor U32594 (N_32594,N_31017,N_31309);
xnor U32595 (N_32595,N_31728,N_31830);
and U32596 (N_32596,N_31240,N_31058);
xnor U32597 (N_32597,N_31720,N_31667);
nand U32598 (N_32598,N_31806,N_31629);
nor U32599 (N_32599,N_31427,N_31819);
and U32600 (N_32600,N_31452,N_31528);
nor U32601 (N_32601,N_31672,N_31727);
or U32602 (N_32602,N_31162,N_31036);
and U32603 (N_32603,N_31928,N_31213);
nor U32604 (N_32604,N_31704,N_31502);
or U32605 (N_32605,N_31347,N_31452);
and U32606 (N_32606,N_31932,N_31281);
or U32607 (N_32607,N_31161,N_31479);
nor U32608 (N_32608,N_31488,N_31097);
and U32609 (N_32609,N_31216,N_31643);
nand U32610 (N_32610,N_31462,N_31313);
or U32611 (N_32611,N_31917,N_31457);
nor U32612 (N_32612,N_31022,N_31426);
nor U32613 (N_32613,N_31074,N_31769);
xor U32614 (N_32614,N_31505,N_31550);
and U32615 (N_32615,N_31710,N_31638);
or U32616 (N_32616,N_31408,N_31478);
nand U32617 (N_32617,N_31672,N_31127);
xor U32618 (N_32618,N_31808,N_31442);
nor U32619 (N_32619,N_31802,N_31244);
and U32620 (N_32620,N_31465,N_31662);
nor U32621 (N_32621,N_31806,N_31899);
nand U32622 (N_32622,N_31285,N_31680);
xnor U32623 (N_32623,N_31236,N_31938);
or U32624 (N_32624,N_31524,N_31219);
nor U32625 (N_32625,N_31981,N_31385);
or U32626 (N_32626,N_31247,N_31160);
and U32627 (N_32627,N_31166,N_31518);
nor U32628 (N_32628,N_31087,N_31614);
nor U32629 (N_32629,N_31237,N_31258);
xnor U32630 (N_32630,N_31933,N_31400);
nand U32631 (N_32631,N_31507,N_31203);
xor U32632 (N_32632,N_31052,N_31714);
nand U32633 (N_32633,N_31637,N_31444);
nor U32634 (N_32634,N_31475,N_31189);
xor U32635 (N_32635,N_31385,N_31558);
xnor U32636 (N_32636,N_31063,N_31590);
nor U32637 (N_32637,N_31575,N_31500);
xnor U32638 (N_32638,N_31350,N_31571);
xor U32639 (N_32639,N_31644,N_31339);
and U32640 (N_32640,N_31518,N_31583);
nor U32641 (N_32641,N_31829,N_31332);
nand U32642 (N_32642,N_31362,N_31849);
nor U32643 (N_32643,N_31846,N_31002);
nor U32644 (N_32644,N_31980,N_31603);
or U32645 (N_32645,N_31275,N_31692);
or U32646 (N_32646,N_31352,N_31113);
xor U32647 (N_32647,N_31329,N_31855);
nor U32648 (N_32648,N_31335,N_31748);
and U32649 (N_32649,N_31893,N_31892);
xor U32650 (N_32650,N_31908,N_31857);
nor U32651 (N_32651,N_31301,N_31348);
nor U32652 (N_32652,N_31020,N_31139);
and U32653 (N_32653,N_31270,N_31280);
xnor U32654 (N_32654,N_31489,N_31178);
and U32655 (N_32655,N_31845,N_31584);
xnor U32656 (N_32656,N_31893,N_31926);
xnor U32657 (N_32657,N_31221,N_31935);
nor U32658 (N_32658,N_31659,N_31263);
xor U32659 (N_32659,N_31558,N_31450);
or U32660 (N_32660,N_31227,N_31888);
and U32661 (N_32661,N_31384,N_31041);
or U32662 (N_32662,N_31807,N_31224);
or U32663 (N_32663,N_31360,N_31159);
or U32664 (N_32664,N_31372,N_31623);
nor U32665 (N_32665,N_31689,N_31844);
or U32666 (N_32666,N_31093,N_31521);
or U32667 (N_32667,N_31578,N_31653);
xnor U32668 (N_32668,N_31623,N_31475);
and U32669 (N_32669,N_31324,N_31078);
or U32670 (N_32670,N_31308,N_31796);
xnor U32671 (N_32671,N_31475,N_31229);
xor U32672 (N_32672,N_31940,N_31153);
and U32673 (N_32673,N_31745,N_31128);
nand U32674 (N_32674,N_31938,N_31086);
nor U32675 (N_32675,N_31450,N_31944);
or U32676 (N_32676,N_31509,N_31529);
or U32677 (N_32677,N_31533,N_31655);
and U32678 (N_32678,N_31707,N_31533);
xnor U32679 (N_32679,N_31758,N_31434);
nand U32680 (N_32680,N_31647,N_31926);
nor U32681 (N_32681,N_31517,N_31504);
or U32682 (N_32682,N_31764,N_31428);
or U32683 (N_32683,N_31050,N_31687);
nand U32684 (N_32684,N_31093,N_31769);
nand U32685 (N_32685,N_31769,N_31632);
and U32686 (N_32686,N_31465,N_31881);
or U32687 (N_32687,N_31978,N_31114);
nor U32688 (N_32688,N_31771,N_31408);
or U32689 (N_32689,N_31168,N_31631);
or U32690 (N_32690,N_31432,N_31317);
and U32691 (N_32691,N_31712,N_31163);
or U32692 (N_32692,N_31008,N_31761);
xor U32693 (N_32693,N_31675,N_31674);
or U32694 (N_32694,N_31787,N_31007);
nand U32695 (N_32695,N_31529,N_31896);
xor U32696 (N_32696,N_31876,N_31598);
or U32697 (N_32697,N_31084,N_31643);
nand U32698 (N_32698,N_31821,N_31726);
nand U32699 (N_32699,N_31147,N_31411);
nor U32700 (N_32700,N_31251,N_31603);
nand U32701 (N_32701,N_31565,N_31459);
or U32702 (N_32702,N_31276,N_31623);
xor U32703 (N_32703,N_31703,N_31968);
or U32704 (N_32704,N_31403,N_31728);
xor U32705 (N_32705,N_31930,N_31804);
xnor U32706 (N_32706,N_31625,N_31447);
xor U32707 (N_32707,N_31631,N_31200);
or U32708 (N_32708,N_31417,N_31155);
or U32709 (N_32709,N_31952,N_31778);
and U32710 (N_32710,N_31082,N_31111);
or U32711 (N_32711,N_31569,N_31297);
nand U32712 (N_32712,N_31855,N_31384);
nand U32713 (N_32713,N_31449,N_31053);
or U32714 (N_32714,N_31402,N_31278);
nor U32715 (N_32715,N_31533,N_31327);
or U32716 (N_32716,N_31342,N_31566);
nor U32717 (N_32717,N_31751,N_31687);
nand U32718 (N_32718,N_31608,N_31488);
nand U32719 (N_32719,N_31472,N_31969);
nand U32720 (N_32720,N_31641,N_31819);
nand U32721 (N_32721,N_31624,N_31098);
and U32722 (N_32722,N_31205,N_31425);
xor U32723 (N_32723,N_31275,N_31179);
or U32724 (N_32724,N_31389,N_31928);
xnor U32725 (N_32725,N_31578,N_31881);
nand U32726 (N_32726,N_31933,N_31534);
xor U32727 (N_32727,N_31420,N_31804);
xnor U32728 (N_32728,N_31609,N_31545);
nand U32729 (N_32729,N_31179,N_31142);
nand U32730 (N_32730,N_31538,N_31945);
nor U32731 (N_32731,N_31895,N_31708);
xnor U32732 (N_32732,N_31864,N_31780);
nand U32733 (N_32733,N_31637,N_31769);
and U32734 (N_32734,N_31216,N_31412);
nor U32735 (N_32735,N_31027,N_31857);
or U32736 (N_32736,N_31719,N_31972);
nor U32737 (N_32737,N_31249,N_31558);
nand U32738 (N_32738,N_31597,N_31531);
nand U32739 (N_32739,N_31495,N_31891);
xor U32740 (N_32740,N_31111,N_31743);
and U32741 (N_32741,N_31647,N_31785);
and U32742 (N_32742,N_31689,N_31050);
xor U32743 (N_32743,N_31666,N_31323);
nand U32744 (N_32744,N_31059,N_31001);
nor U32745 (N_32745,N_31771,N_31579);
or U32746 (N_32746,N_31411,N_31074);
or U32747 (N_32747,N_31345,N_31360);
or U32748 (N_32748,N_31243,N_31011);
nor U32749 (N_32749,N_31248,N_31105);
or U32750 (N_32750,N_31628,N_31689);
nand U32751 (N_32751,N_31298,N_31755);
nor U32752 (N_32752,N_31891,N_31635);
xor U32753 (N_32753,N_31400,N_31360);
xnor U32754 (N_32754,N_31264,N_31700);
or U32755 (N_32755,N_31110,N_31752);
xnor U32756 (N_32756,N_31100,N_31040);
nor U32757 (N_32757,N_31900,N_31054);
and U32758 (N_32758,N_31885,N_31324);
nand U32759 (N_32759,N_31327,N_31603);
and U32760 (N_32760,N_31073,N_31013);
xor U32761 (N_32761,N_31381,N_31585);
xor U32762 (N_32762,N_31065,N_31800);
xnor U32763 (N_32763,N_31755,N_31768);
xor U32764 (N_32764,N_31182,N_31844);
or U32765 (N_32765,N_31026,N_31642);
nand U32766 (N_32766,N_31630,N_31961);
nor U32767 (N_32767,N_31929,N_31897);
xor U32768 (N_32768,N_31491,N_31769);
nor U32769 (N_32769,N_31384,N_31893);
nor U32770 (N_32770,N_31949,N_31049);
nand U32771 (N_32771,N_31730,N_31562);
xor U32772 (N_32772,N_31233,N_31748);
nor U32773 (N_32773,N_31590,N_31468);
nand U32774 (N_32774,N_31008,N_31222);
or U32775 (N_32775,N_31930,N_31559);
and U32776 (N_32776,N_31832,N_31685);
nand U32777 (N_32777,N_31938,N_31531);
nand U32778 (N_32778,N_31678,N_31754);
and U32779 (N_32779,N_31201,N_31533);
and U32780 (N_32780,N_31917,N_31826);
and U32781 (N_32781,N_31250,N_31838);
nand U32782 (N_32782,N_31141,N_31131);
nor U32783 (N_32783,N_31620,N_31659);
or U32784 (N_32784,N_31724,N_31697);
or U32785 (N_32785,N_31660,N_31310);
xnor U32786 (N_32786,N_31070,N_31846);
xor U32787 (N_32787,N_31107,N_31093);
xnor U32788 (N_32788,N_31868,N_31114);
xor U32789 (N_32789,N_31193,N_31130);
xor U32790 (N_32790,N_31576,N_31007);
xor U32791 (N_32791,N_31540,N_31188);
nor U32792 (N_32792,N_31636,N_31734);
xnor U32793 (N_32793,N_31454,N_31868);
and U32794 (N_32794,N_31349,N_31764);
and U32795 (N_32795,N_31689,N_31040);
and U32796 (N_32796,N_31714,N_31843);
nor U32797 (N_32797,N_31037,N_31305);
nor U32798 (N_32798,N_31280,N_31938);
and U32799 (N_32799,N_31399,N_31618);
and U32800 (N_32800,N_31140,N_31740);
nor U32801 (N_32801,N_31657,N_31635);
xor U32802 (N_32802,N_31721,N_31297);
or U32803 (N_32803,N_31100,N_31208);
or U32804 (N_32804,N_31939,N_31415);
nand U32805 (N_32805,N_31386,N_31211);
xnor U32806 (N_32806,N_31002,N_31849);
nand U32807 (N_32807,N_31812,N_31896);
nor U32808 (N_32808,N_31999,N_31827);
or U32809 (N_32809,N_31964,N_31980);
nand U32810 (N_32810,N_31958,N_31526);
nand U32811 (N_32811,N_31148,N_31523);
xor U32812 (N_32812,N_31235,N_31920);
nor U32813 (N_32813,N_31926,N_31694);
and U32814 (N_32814,N_31712,N_31977);
and U32815 (N_32815,N_31997,N_31210);
nor U32816 (N_32816,N_31607,N_31851);
or U32817 (N_32817,N_31425,N_31579);
nor U32818 (N_32818,N_31778,N_31226);
or U32819 (N_32819,N_31313,N_31020);
nand U32820 (N_32820,N_31562,N_31092);
xor U32821 (N_32821,N_31263,N_31982);
xnor U32822 (N_32822,N_31850,N_31789);
or U32823 (N_32823,N_31178,N_31240);
nand U32824 (N_32824,N_31527,N_31718);
and U32825 (N_32825,N_31284,N_31058);
nand U32826 (N_32826,N_31092,N_31764);
or U32827 (N_32827,N_31833,N_31324);
and U32828 (N_32828,N_31043,N_31217);
nand U32829 (N_32829,N_31149,N_31048);
xor U32830 (N_32830,N_31778,N_31076);
nor U32831 (N_32831,N_31997,N_31381);
nor U32832 (N_32832,N_31001,N_31631);
and U32833 (N_32833,N_31573,N_31894);
nand U32834 (N_32834,N_31341,N_31059);
xor U32835 (N_32835,N_31446,N_31606);
nor U32836 (N_32836,N_31660,N_31022);
nand U32837 (N_32837,N_31506,N_31695);
nand U32838 (N_32838,N_31898,N_31080);
and U32839 (N_32839,N_31146,N_31698);
xnor U32840 (N_32840,N_31700,N_31455);
and U32841 (N_32841,N_31528,N_31340);
nand U32842 (N_32842,N_31451,N_31053);
or U32843 (N_32843,N_31520,N_31606);
xnor U32844 (N_32844,N_31619,N_31505);
or U32845 (N_32845,N_31854,N_31928);
nand U32846 (N_32846,N_31256,N_31919);
nand U32847 (N_32847,N_31454,N_31032);
xnor U32848 (N_32848,N_31203,N_31966);
xor U32849 (N_32849,N_31563,N_31873);
and U32850 (N_32850,N_31374,N_31031);
or U32851 (N_32851,N_31095,N_31705);
and U32852 (N_32852,N_31098,N_31970);
or U32853 (N_32853,N_31026,N_31698);
xor U32854 (N_32854,N_31634,N_31012);
nor U32855 (N_32855,N_31551,N_31423);
xnor U32856 (N_32856,N_31298,N_31193);
and U32857 (N_32857,N_31082,N_31381);
nand U32858 (N_32858,N_31151,N_31210);
nor U32859 (N_32859,N_31027,N_31561);
nor U32860 (N_32860,N_31834,N_31994);
or U32861 (N_32861,N_31309,N_31025);
or U32862 (N_32862,N_31490,N_31973);
nand U32863 (N_32863,N_31708,N_31475);
or U32864 (N_32864,N_31919,N_31814);
and U32865 (N_32865,N_31716,N_31496);
xnor U32866 (N_32866,N_31777,N_31027);
and U32867 (N_32867,N_31737,N_31274);
nand U32868 (N_32868,N_31327,N_31721);
or U32869 (N_32869,N_31643,N_31324);
or U32870 (N_32870,N_31812,N_31431);
nor U32871 (N_32871,N_31795,N_31132);
nor U32872 (N_32872,N_31078,N_31061);
and U32873 (N_32873,N_31359,N_31389);
and U32874 (N_32874,N_31164,N_31667);
nor U32875 (N_32875,N_31491,N_31999);
and U32876 (N_32876,N_31054,N_31184);
nand U32877 (N_32877,N_31185,N_31651);
and U32878 (N_32878,N_31044,N_31022);
nor U32879 (N_32879,N_31587,N_31333);
or U32880 (N_32880,N_31879,N_31809);
nand U32881 (N_32881,N_31392,N_31442);
or U32882 (N_32882,N_31156,N_31655);
or U32883 (N_32883,N_31714,N_31114);
and U32884 (N_32884,N_31486,N_31595);
xnor U32885 (N_32885,N_31360,N_31507);
nor U32886 (N_32886,N_31412,N_31297);
xnor U32887 (N_32887,N_31658,N_31899);
nand U32888 (N_32888,N_31475,N_31115);
xor U32889 (N_32889,N_31094,N_31645);
nand U32890 (N_32890,N_31940,N_31644);
xnor U32891 (N_32891,N_31588,N_31144);
or U32892 (N_32892,N_31248,N_31978);
or U32893 (N_32893,N_31541,N_31956);
nand U32894 (N_32894,N_31925,N_31127);
nand U32895 (N_32895,N_31795,N_31488);
nor U32896 (N_32896,N_31692,N_31142);
or U32897 (N_32897,N_31405,N_31213);
nand U32898 (N_32898,N_31103,N_31789);
nand U32899 (N_32899,N_31704,N_31966);
xor U32900 (N_32900,N_31680,N_31928);
nand U32901 (N_32901,N_31619,N_31264);
nor U32902 (N_32902,N_31235,N_31174);
nand U32903 (N_32903,N_31556,N_31680);
and U32904 (N_32904,N_31098,N_31215);
nor U32905 (N_32905,N_31522,N_31257);
or U32906 (N_32906,N_31376,N_31709);
nand U32907 (N_32907,N_31814,N_31654);
or U32908 (N_32908,N_31525,N_31561);
xnor U32909 (N_32909,N_31222,N_31255);
or U32910 (N_32910,N_31605,N_31763);
xor U32911 (N_32911,N_31107,N_31439);
nand U32912 (N_32912,N_31960,N_31464);
nand U32913 (N_32913,N_31296,N_31972);
and U32914 (N_32914,N_31130,N_31608);
and U32915 (N_32915,N_31950,N_31323);
xor U32916 (N_32916,N_31597,N_31000);
and U32917 (N_32917,N_31007,N_31622);
nor U32918 (N_32918,N_31879,N_31782);
nand U32919 (N_32919,N_31174,N_31029);
xor U32920 (N_32920,N_31856,N_31040);
nor U32921 (N_32921,N_31117,N_31867);
and U32922 (N_32922,N_31470,N_31301);
or U32923 (N_32923,N_31711,N_31959);
and U32924 (N_32924,N_31857,N_31025);
and U32925 (N_32925,N_31243,N_31192);
nor U32926 (N_32926,N_31790,N_31921);
nor U32927 (N_32927,N_31741,N_31510);
and U32928 (N_32928,N_31473,N_31996);
or U32929 (N_32929,N_31221,N_31280);
nor U32930 (N_32930,N_31486,N_31001);
xor U32931 (N_32931,N_31940,N_31357);
nor U32932 (N_32932,N_31377,N_31605);
nand U32933 (N_32933,N_31972,N_31183);
or U32934 (N_32934,N_31202,N_31861);
nor U32935 (N_32935,N_31311,N_31126);
nand U32936 (N_32936,N_31835,N_31860);
nand U32937 (N_32937,N_31247,N_31934);
or U32938 (N_32938,N_31748,N_31191);
nand U32939 (N_32939,N_31196,N_31248);
nor U32940 (N_32940,N_31877,N_31180);
and U32941 (N_32941,N_31874,N_31808);
nor U32942 (N_32942,N_31451,N_31640);
nor U32943 (N_32943,N_31348,N_31043);
xnor U32944 (N_32944,N_31760,N_31887);
xor U32945 (N_32945,N_31668,N_31955);
xor U32946 (N_32946,N_31863,N_31462);
nand U32947 (N_32947,N_31197,N_31483);
nand U32948 (N_32948,N_31962,N_31098);
nor U32949 (N_32949,N_31793,N_31720);
xor U32950 (N_32950,N_31037,N_31029);
xor U32951 (N_32951,N_31581,N_31109);
nand U32952 (N_32952,N_31024,N_31618);
xnor U32953 (N_32953,N_31753,N_31010);
or U32954 (N_32954,N_31712,N_31703);
xor U32955 (N_32955,N_31906,N_31175);
xor U32956 (N_32956,N_31232,N_31885);
or U32957 (N_32957,N_31175,N_31591);
or U32958 (N_32958,N_31165,N_31815);
and U32959 (N_32959,N_31631,N_31802);
xnor U32960 (N_32960,N_31266,N_31791);
nor U32961 (N_32961,N_31518,N_31288);
nor U32962 (N_32962,N_31443,N_31467);
nand U32963 (N_32963,N_31690,N_31078);
and U32964 (N_32964,N_31715,N_31145);
nand U32965 (N_32965,N_31847,N_31362);
nor U32966 (N_32966,N_31576,N_31764);
xor U32967 (N_32967,N_31346,N_31209);
and U32968 (N_32968,N_31878,N_31452);
and U32969 (N_32969,N_31431,N_31342);
nand U32970 (N_32970,N_31499,N_31084);
or U32971 (N_32971,N_31015,N_31180);
and U32972 (N_32972,N_31539,N_31454);
nor U32973 (N_32973,N_31064,N_31182);
and U32974 (N_32974,N_31892,N_31431);
nor U32975 (N_32975,N_31566,N_31163);
and U32976 (N_32976,N_31030,N_31587);
nand U32977 (N_32977,N_31414,N_31352);
nand U32978 (N_32978,N_31896,N_31536);
and U32979 (N_32979,N_31985,N_31507);
and U32980 (N_32980,N_31410,N_31734);
nor U32981 (N_32981,N_31732,N_31331);
nand U32982 (N_32982,N_31447,N_31371);
nand U32983 (N_32983,N_31398,N_31960);
xnor U32984 (N_32984,N_31032,N_31400);
xnor U32985 (N_32985,N_31865,N_31082);
or U32986 (N_32986,N_31145,N_31023);
or U32987 (N_32987,N_31236,N_31700);
nand U32988 (N_32988,N_31672,N_31657);
xnor U32989 (N_32989,N_31276,N_31183);
and U32990 (N_32990,N_31645,N_31459);
and U32991 (N_32991,N_31092,N_31717);
nand U32992 (N_32992,N_31197,N_31935);
and U32993 (N_32993,N_31324,N_31741);
nor U32994 (N_32994,N_31697,N_31672);
nand U32995 (N_32995,N_31069,N_31846);
xor U32996 (N_32996,N_31753,N_31149);
nand U32997 (N_32997,N_31963,N_31654);
or U32998 (N_32998,N_31195,N_31931);
nand U32999 (N_32999,N_31872,N_31862);
or U33000 (N_33000,N_32995,N_32975);
nor U33001 (N_33001,N_32184,N_32614);
xor U33002 (N_33002,N_32670,N_32831);
nand U33003 (N_33003,N_32113,N_32430);
or U33004 (N_33004,N_32931,N_32538);
nor U33005 (N_33005,N_32900,N_32007);
and U33006 (N_33006,N_32508,N_32862);
nor U33007 (N_33007,N_32445,N_32453);
nand U33008 (N_33008,N_32767,N_32652);
or U33009 (N_33009,N_32640,N_32258);
or U33010 (N_33010,N_32903,N_32738);
or U33011 (N_33011,N_32690,N_32618);
nand U33012 (N_33012,N_32298,N_32211);
nand U33013 (N_33013,N_32192,N_32491);
or U33014 (N_33014,N_32165,N_32342);
xor U33015 (N_33015,N_32979,N_32700);
nor U33016 (N_33016,N_32697,N_32511);
nor U33017 (N_33017,N_32300,N_32307);
and U33018 (N_33018,N_32568,N_32725);
nand U33019 (N_33019,N_32660,N_32658);
xor U33020 (N_33020,N_32191,N_32672);
nand U33021 (N_33021,N_32381,N_32205);
xnor U33022 (N_33022,N_32848,N_32504);
and U33023 (N_33023,N_32454,N_32262);
nor U33024 (N_33024,N_32280,N_32629);
or U33025 (N_33025,N_32040,N_32777);
nor U33026 (N_33026,N_32970,N_32460);
nor U33027 (N_33027,N_32632,N_32094);
xnor U33028 (N_33028,N_32240,N_32023);
nand U33029 (N_33029,N_32733,N_32420);
xnor U33030 (N_33030,N_32877,N_32325);
nand U33031 (N_33031,N_32013,N_32439);
nor U33032 (N_33032,N_32278,N_32625);
nor U33033 (N_33033,N_32729,N_32084);
and U33034 (N_33034,N_32691,N_32082);
nor U33035 (N_33035,N_32813,N_32047);
or U33036 (N_33036,N_32510,N_32586);
and U33037 (N_33037,N_32009,N_32748);
and U33038 (N_33038,N_32150,N_32461);
or U33039 (N_33039,N_32668,N_32999);
or U33040 (N_33040,N_32254,N_32261);
and U33041 (N_33041,N_32923,N_32216);
xnor U33042 (N_33042,N_32433,N_32214);
or U33043 (N_33043,N_32967,N_32768);
or U33044 (N_33044,N_32056,N_32869);
nand U33045 (N_33045,N_32621,N_32006);
and U33046 (N_33046,N_32126,N_32030);
nor U33047 (N_33047,N_32627,N_32789);
or U33048 (N_33048,N_32086,N_32277);
nor U33049 (N_33049,N_32354,N_32180);
xor U33050 (N_33050,N_32146,N_32512);
nand U33051 (N_33051,N_32236,N_32819);
nand U33052 (N_33052,N_32814,N_32521);
and U33053 (N_33053,N_32447,N_32498);
nor U33054 (N_33054,N_32939,N_32908);
xor U33055 (N_33055,N_32393,N_32032);
xor U33056 (N_33056,N_32707,N_32624);
xor U33057 (N_33057,N_32332,N_32988);
nand U33058 (N_33058,N_32615,N_32020);
nand U33059 (N_33059,N_32477,N_32158);
and U33060 (N_33060,N_32764,N_32513);
nand U33061 (N_33061,N_32699,N_32945);
xnor U33062 (N_33062,N_32693,N_32343);
nor U33063 (N_33063,N_32751,N_32390);
and U33064 (N_33064,N_32646,N_32626);
and U33065 (N_33065,N_32799,N_32259);
nor U33066 (N_33066,N_32688,N_32266);
xor U33067 (N_33067,N_32943,N_32299);
nor U33068 (N_33068,N_32893,N_32302);
or U33069 (N_33069,N_32228,N_32068);
nor U33070 (N_33070,N_32643,N_32283);
or U33071 (N_33071,N_32328,N_32352);
or U33072 (N_33072,N_32069,N_32155);
or U33073 (N_33073,N_32936,N_32090);
or U33074 (N_33074,N_32845,N_32924);
nand U33075 (N_33075,N_32832,N_32516);
nor U33076 (N_33076,N_32846,N_32217);
and U33077 (N_33077,N_32487,N_32589);
xnor U33078 (N_33078,N_32860,N_32138);
xnor U33079 (N_33079,N_32049,N_32909);
xnor U33080 (N_33080,N_32245,N_32617);
and U33081 (N_33081,N_32288,N_32530);
or U33082 (N_33082,N_32115,N_32152);
xor U33083 (N_33083,N_32054,N_32651);
nand U33084 (N_33084,N_32575,N_32244);
and U33085 (N_33085,N_32166,N_32061);
or U33086 (N_33086,N_32557,N_32016);
nor U33087 (N_33087,N_32494,N_32720);
nor U33088 (N_33088,N_32440,N_32297);
nor U33089 (N_33089,N_32935,N_32559);
nand U33090 (N_33090,N_32857,N_32647);
nand U33091 (N_33091,N_32329,N_32518);
or U33092 (N_33092,N_32687,N_32597);
nand U33093 (N_33093,N_32947,N_32224);
xnor U33094 (N_33094,N_32949,N_32401);
nor U33095 (N_33095,N_32196,N_32735);
nor U33096 (N_33096,N_32271,N_32787);
or U33097 (N_33097,N_32427,N_32823);
and U33098 (N_33098,N_32102,N_32983);
nand U33099 (N_33099,N_32728,N_32984);
nand U33100 (N_33100,N_32792,N_32774);
nand U33101 (N_33101,N_32019,N_32659);
and U33102 (N_33102,N_32482,N_32556);
nor U33103 (N_33103,N_32472,N_32035);
nand U33104 (N_33104,N_32669,N_32466);
xor U33105 (N_33105,N_32622,N_32143);
nand U33106 (N_33106,N_32847,N_32046);
nand U33107 (N_33107,N_32305,N_32679);
and U33108 (N_33108,N_32220,N_32083);
or U33109 (N_33109,N_32481,N_32136);
or U33110 (N_33110,N_32964,N_32114);
or U33111 (N_33111,N_32552,N_32858);
or U33112 (N_33112,N_32092,N_32279);
nor U33113 (N_33113,N_32957,N_32149);
and U33114 (N_33114,N_32921,N_32806);
and U33115 (N_33115,N_32140,N_32874);
nor U33116 (N_33116,N_32580,N_32844);
and U33117 (N_33117,N_32854,N_32934);
nand U33118 (N_33118,N_32418,N_32043);
nor U33119 (N_33119,N_32331,N_32375);
nand U33120 (N_33120,N_32930,N_32075);
and U33121 (N_33121,N_32800,N_32027);
xor U33122 (N_33122,N_32085,N_32241);
and U33123 (N_33123,N_32801,N_32443);
nor U33124 (N_33124,N_32260,N_32663);
and U33125 (N_33125,N_32937,N_32782);
nor U33126 (N_33126,N_32793,N_32605);
or U33127 (N_33127,N_32219,N_32435);
nor U33128 (N_33128,N_32692,N_32414);
or U33129 (N_33129,N_32028,N_32103);
xnor U33130 (N_33130,N_32355,N_32649);
nand U33131 (N_33131,N_32384,N_32594);
xnor U33132 (N_33132,N_32168,N_32110);
nand U33133 (N_33133,N_32486,N_32074);
or U33134 (N_33134,N_32592,N_32250);
and U33135 (N_33135,N_32497,N_32856);
nor U33136 (N_33136,N_32387,N_32717);
nor U33137 (N_33137,N_32958,N_32405);
nand U33138 (N_33138,N_32601,N_32509);
or U33139 (N_33139,N_32749,N_32351);
or U33140 (N_33140,N_32914,N_32173);
nor U33141 (N_33141,N_32213,N_32636);
and U33142 (N_33142,N_32225,N_32135);
nor U33143 (N_33143,N_32318,N_32628);
and U33144 (N_33144,N_32536,N_32826);
or U33145 (N_33145,N_32109,N_32662);
or U33146 (N_33146,N_32031,N_32133);
nand U33147 (N_33147,N_32992,N_32769);
nand U33148 (N_33148,N_32235,N_32422);
nand U33149 (N_33149,N_32489,N_32545);
nor U33150 (N_33150,N_32891,N_32177);
nand U33151 (N_33151,N_32711,N_32501);
or U33152 (N_33152,N_32033,N_32503);
and U33153 (N_33153,N_32396,N_32174);
and U33154 (N_33154,N_32522,N_32063);
or U33155 (N_33155,N_32452,N_32849);
nor U33156 (N_33156,N_32872,N_32505);
and U33157 (N_33157,N_32912,N_32765);
and U33158 (N_33158,N_32886,N_32423);
or U33159 (N_33159,N_32502,N_32195);
nor U33160 (N_33160,N_32336,N_32517);
nand U33161 (N_33161,N_32276,N_32760);
nand U33162 (N_33162,N_32602,N_32871);
nor U33163 (N_33163,N_32436,N_32327);
xnor U33164 (N_33164,N_32051,N_32383);
nor U33165 (N_33165,N_32002,N_32805);
nor U33166 (N_33166,N_32685,N_32001);
and U33167 (N_33167,N_32005,N_32493);
nor U33168 (N_33168,N_32755,N_32784);
and U33169 (N_33169,N_32229,N_32323);
nor U33170 (N_33170,N_32780,N_32012);
nor U33171 (N_33171,N_32052,N_32242);
nor U33172 (N_33172,N_32475,N_32314);
nand U33173 (N_33173,N_32956,N_32053);
nand U33174 (N_33174,N_32108,N_32585);
and U33175 (N_33175,N_32024,N_32121);
nor U33176 (N_33176,N_32710,N_32920);
or U33177 (N_33177,N_32918,N_32036);
xor U33178 (N_33178,N_32127,N_32570);
xnor U33179 (N_33179,N_32131,N_32123);
and U33180 (N_33180,N_32596,N_32320);
or U33181 (N_33181,N_32607,N_32471);
nor U33182 (N_33182,N_32850,N_32761);
nor U33183 (N_33183,N_32790,N_32441);
xnor U33184 (N_33184,N_32917,N_32786);
and U33185 (N_33185,N_32188,N_32535);
or U33186 (N_33186,N_32122,N_32011);
nor U33187 (N_33187,N_32997,N_32316);
and U33188 (N_33188,N_32894,N_32066);
nor U33189 (N_33189,N_32574,N_32932);
and U33190 (N_33190,N_32795,N_32137);
and U33191 (N_33191,N_32175,N_32204);
nor U33192 (N_33192,N_32953,N_32630);
nor U33193 (N_33193,N_32341,N_32546);
or U33194 (N_33194,N_32715,N_32081);
nand U33195 (N_33195,N_32008,N_32639);
or U33196 (N_33196,N_32419,N_32252);
nand U33197 (N_33197,N_32529,N_32201);
or U33198 (N_33198,N_32386,N_32408);
nand U33199 (N_33199,N_32994,N_32425);
xor U33200 (N_33200,N_32548,N_32695);
nor U33201 (N_33201,N_32657,N_32426);
or U33202 (N_33202,N_32785,N_32706);
nor U33203 (N_33203,N_32179,N_32286);
and U33204 (N_33204,N_32099,N_32678);
xnor U33205 (N_33205,N_32208,N_32634);
nor U33206 (N_33206,N_32349,N_32759);
and U33207 (N_33207,N_32287,N_32238);
or U33208 (N_33208,N_32340,N_32282);
xor U33209 (N_33209,N_32723,N_32274);
and U33210 (N_33210,N_32221,N_32797);
nand U33211 (N_33211,N_32904,N_32972);
and U33212 (N_33212,N_32551,N_32878);
nand U33213 (N_33213,N_32256,N_32484);
nor U33214 (N_33214,N_32257,N_32458);
nand U33215 (N_33215,N_32822,N_32273);
xor U33216 (N_33216,N_32233,N_32210);
xor U33217 (N_33217,N_32485,N_32993);
nand U33218 (N_33218,N_32112,N_32284);
or U33219 (N_33219,N_32772,N_32807);
or U33220 (N_33220,N_32434,N_32852);
or U33221 (N_33221,N_32916,N_32524);
nand U33222 (N_33222,N_32243,N_32062);
or U33223 (N_33223,N_32868,N_32808);
and U33224 (N_33224,N_32388,N_32358);
and U33225 (N_33225,N_32803,N_32281);
and U33226 (N_33226,N_32480,N_32673);
and U33227 (N_33227,N_32863,N_32335);
nand U33228 (N_33228,N_32413,N_32495);
and U33229 (N_33229,N_32896,N_32442);
and U33230 (N_33230,N_32468,N_32839);
xor U33231 (N_33231,N_32161,N_32778);
xor U33232 (N_33232,N_32398,N_32169);
xor U33233 (N_33233,N_32162,N_32264);
or U33234 (N_33234,N_32773,N_32843);
or U33235 (N_33235,N_32783,N_32523);
nor U33236 (N_33236,N_32952,N_32312);
xnor U33237 (N_33237,N_32534,N_32563);
or U33238 (N_33238,N_32378,N_32400);
nand U33239 (N_33239,N_32093,N_32724);
nor U33240 (N_33240,N_32719,N_32895);
or U33241 (N_33241,N_32206,N_32105);
and U33242 (N_33242,N_32057,N_32215);
and U33243 (N_33243,N_32731,N_32187);
nand U33244 (N_33244,N_32681,N_32752);
and U33245 (N_33245,N_32925,N_32290);
or U33246 (N_33246,N_32680,N_32567);
or U33247 (N_33247,N_32897,N_32721);
and U33248 (N_33248,N_32835,N_32569);
nand U33249 (N_33249,N_32412,N_32754);
and U33250 (N_33250,N_32541,N_32701);
or U33251 (N_33251,N_32553,N_32407);
or U33252 (N_33252,N_32488,N_32403);
nor U33253 (N_33253,N_32644,N_32247);
nand U33254 (N_33254,N_32665,N_32415);
nor U33255 (N_33255,N_32821,N_32326);
nor U33256 (N_33256,N_32620,N_32348);
and U33257 (N_33257,N_32160,N_32292);
or U33258 (N_33258,N_32989,N_32885);
and U33259 (N_33259,N_32543,N_32392);
nor U33260 (N_33260,N_32611,N_32128);
or U33261 (N_33261,N_32101,N_32587);
and U33262 (N_33262,N_32368,N_32479);
and U33263 (N_33263,N_32170,N_32591);
nand U33264 (N_33264,N_32653,N_32178);
nand U33265 (N_33265,N_32058,N_32365);
nand U33266 (N_33266,N_32042,N_32892);
or U33267 (N_33267,N_32406,N_32986);
nand U33268 (N_33268,N_32185,N_32671);
nand U33269 (N_33269,N_32294,N_32978);
nand U33270 (N_33270,N_32791,N_32740);
and U33271 (N_33271,N_32437,N_32927);
or U33272 (N_33272,N_32507,N_32391);
or U33273 (N_33273,N_32537,N_32815);
xnor U33274 (N_33274,N_32572,N_32990);
and U33275 (N_33275,N_32315,N_32026);
nor U33276 (N_33276,N_32705,N_32291);
and U33277 (N_33277,N_32802,N_32582);
xor U33278 (N_33278,N_32370,N_32593);
or U33279 (N_33279,N_32525,N_32842);
xor U33280 (N_33280,N_32041,N_32404);
xor U33281 (N_33281,N_32709,N_32189);
or U33282 (N_33282,N_32595,N_32684);
or U33283 (N_33283,N_32588,N_32890);
nand U33284 (N_33284,N_32411,N_32817);
nand U33285 (N_33285,N_32467,N_32533);
nor U33286 (N_33286,N_32638,N_32884);
nor U33287 (N_33287,N_32633,N_32267);
xnor U33288 (N_33288,N_32076,N_32203);
nand U33289 (N_33289,N_32377,N_32462);
nand U33290 (N_33290,N_32828,N_32876);
xor U33291 (N_33291,N_32116,N_32870);
or U33292 (N_33292,N_32132,N_32141);
and U33293 (N_33293,N_32337,N_32718);
nand U33294 (N_33294,N_32067,N_32139);
nor U33295 (N_33295,N_32003,N_32955);
nor U33296 (N_33296,N_32347,N_32741);
and U33297 (N_33297,N_32004,N_32528);
xor U33298 (N_33298,N_32478,N_32527);
or U33299 (N_33299,N_32492,N_32322);
and U33300 (N_33300,N_32324,N_32374);
or U33301 (N_33301,N_32641,N_32038);
or U33302 (N_33302,N_32227,N_32455);
nand U33303 (N_33303,N_32609,N_32014);
nor U33304 (N_33304,N_32416,N_32577);
xor U33305 (N_33305,N_32985,N_32645);
xnor U33306 (N_33306,N_32550,N_32199);
nand U33307 (N_33307,N_32350,N_32459);
nand U33308 (N_33308,N_32071,N_32410);
xor U33309 (N_33309,N_32451,N_32704);
xor U33310 (N_33310,N_32450,N_32500);
or U33311 (N_33311,N_32147,N_32861);
or U33312 (N_33312,N_32864,N_32654);
xnor U33313 (N_33313,N_32584,N_32382);
nor U33314 (N_33314,N_32303,N_32558);
or U33315 (N_33315,N_32186,N_32106);
xnor U33316 (N_33316,N_32376,N_32833);
xor U33317 (N_33317,N_32309,N_32853);
or U33318 (N_33318,N_32666,N_32674);
or U33319 (N_33319,N_32223,N_32334);
and U33320 (N_33320,N_32726,N_32739);
nand U33321 (N_33321,N_32851,N_32088);
or U33322 (N_33322,N_32825,N_32747);
nor U33323 (N_33323,N_32565,N_32465);
nand U33324 (N_33324,N_32766,N_32713);
or U33325 (N_33325,N_32855,N_32954);
xor U33326 (N_33326,N_32980,N_32018);
or U33327 (N_33327,N_32942,N_32623);
or U33328 (N_33328,N_32310,N_32712);
xor U33329 (N_33329,N_32603,N_32176);
and U33330 (N_33330,N_32838,N_32163);
xnor U33331 (N_33331,N_32330,N_32446);
nor U33332 (N_33332,N_32702,N_32910);
xor U33333 (N_33333,N_32125,N_32899);
nand U33334 (N_33334,N_32059,N_32490);
or U33335 (N_33335,N_32599,N_32432);
nand U33336 (N_33336,N_32564,N_32207);
xnor U33337 (N_33337,N_32218,N_32519);
xor U33338 (N_33338,N_32015,N_32022);
or U33339 (N_33339,N_32100,N_32532);
nor U33340 (N_33340,N_32246,N_32362);
nor U33341 (N_33341,N_32096,N_32514);
or U33342 (N_33342,N_32667,N_32742);
and U33343 (N_33343,N_32148,N_32963);
or U33344 (N_33344,N_32919,N_32034);
and U33345 (N_33345,N_32029,N_32431);
nand U33346 (N_33346,N_32880,N_32360);
xnor U33347 (N_33347,N_32976,N_32982);
xnor U33348 (N_33348,N_32873,N_32496);
xor U33349 (N_33349,N_32130,N_32159);
nor U33350 (N_33350,N_32198,N_32560);
nand U33351 (N_33351,N_32289,N_32397);
and U33352 (N_33352,N_32824,N_32399);
nand U33353 (N_33353,N_32077,N_32542);
and U33354 (N_33354,N_32590,N_32317);
and U33355 (N_33355,N_32065,N_32608);
or U33356 (N_33356,N_32356,N_32474);
nor U33357 (N_33357,N_32987,N_32212);
nor U33358 (N_33358,N_32762,N_32827);
nor U33359 (N_33359,N_32736,N_32193);
nor U33360 (N_33360,N_32463,N_32293);
nand U33361 (N_33361,N_32648,N_32369);
nor U33362 (N_33362,N_32157,N_32818);
or U33363 (N_33363,N_32239,N_32371);
xnor U33364 (N_33364,N_32222,N_32270);
and U33365 (N_33365,N_32859,N_32888);
or U33366 (N_33366,N_32714,N_32268);
nor U33367 (N_33367,N_32194,N_32091);
nand U33368 (N_33368,N_32010,N_32938);
nand U33369 (N_33369,N_32637,N_32750);
xnor U33370 (N_33370,N_32866,N_32961);
xnor U33371 (N_33371,N_32913,N_32424);
xnor U33372 (N_33372,N_32734,N_32037);
xor U33373 (N_33373,N_32579,N_32928);
and U33374 (N_33374,N_32120,N_32539);
or U33375 (N_33375,N_32867,N_32879);
or U33376 (N_33376,N_32794,N_32746);
nor U33377 (N_33377,N_32922,N_32064);
nand U33378 (N_33378,N_32576,N_32642);
or U33379 (N_33379,N_32156,N_32346);
and U33380 (N_33380,N_32313,N_32788);
xnor U33381 (N_33381,N_32991,N_32675);
or U33382 (N_33382,N_32696,N_32363);
or U33383 (N_33383,N_32732,N_32044);
nand U33384 (N_33384,N_32200,N_32929);
or U33385 (N_33385,N_32811,N_32448);
and U33386 (N_33386,N_32619,N_32809);
or U33387 (N_33387,N_32973,N_32578);
and U33388 (N_33388,N_32950,N_32145);
nand U33389 (N_33389,N_32359,N_32457);
and U33390 (N_33390,N_32758,N_32745);
nand U33391 (N_33391,N_32965,N_32962);
or U33392 (N_33392,N_32119,N_32840);
nor U33393 (N_33393,N_32107,N_32164);
and U33394 (N_33394,N_32689,N_32171);
nand U33395 (N_33395,N_32499,N_32249);
or U33396 (N_33396,N_32237,N_32781);
nand U33397 (N_33397,N_32875,N_32154);
nor U33398 (N_33398,N_32079,N_32757);
nor U33399 (N_33399,N_32295,N_32134);
or U33400 (N_33400,N_32664,N_32902);
and U33401 (N_33401,N_32798,N_32078);
nand U33402 (N_33402,N_32409,N_32181);
xor U33403 (N_33403,N_32946,N_32344);
or U33404 (N_33404,N_32060,N_32476);
nor U33405 (N_33405,N_32944,N_32703);
and U33406 (N_33406,N_32951,N_32661);
nor U33407 (N_33407,N_32470,N_32379);
xnor U33408 (N_33408,N_32039,N_32232);
or U33409 (N_33409,N_32153,N_32683);
or U33410 (N_33410,N_32686,N_32776);
or U33411 (N_33411,N_32357,N_32395);
nand U33412 (N_33412,N_32438,N_32421);
nand U33413 (N_33413,N_32562,N_32708);
and U33414 (N_33414,N_32183,N_32095);
nand U33415 (N_33415,N_32561,N_32142);
and U33416 (N_33416,N_32429,N_32339);
nor U33417 (N_33417,N_32255,N_32385);
xor U33418 (N_33418,N_32526,N_32977);
xor U33419 (N_33419,N_32650,N_32829);
or U33420 (N_33420,N_32655,N_32098);
and U33421 (N_33421,N_32000,N_32775);
xor U33422 (N_33422,N_32906,N_32959);
xor U33423 (N_33423,N_32926,N_32540);
xnor U33424 (N_33424,N_32272,N_32124);
and U33425 (N_33425,N_32981,N_32771);
xor U33426 (N_33426,N_32830,N_32402);
or U33427 (N_33427,N_32087,N_32190);
nand U33428 (N_33428,N_32070,N_32209);
nor U33429 (N_33429,N_32265,N_32616);
and U33430 (N_33430,N_32389,N_32367);
or U33431 (N_33431,N_32469,N_32968);
or U33432 (N_33432,N_32231,N_32333);
or U33433 (N_33433,N_32554,N_32167);
nand U33434 (N_33434,N_32915,N_32940);
xor U33435 (N_33435,N_32549,N_32072);
or U33436 (N_33436,N_32048,N_32373);
or U33437 (N_33437,N_32117,N_32045);
nor U33438 (N_33438,N_32882,N_32428);
nor U33439 (N_33439,N_32812,N_32531);
or U33440 (N_33440,N_32364,N_32129);
nor U33441 (N_33441,N_32635,N_32050);
and U33442 (N_33442,N_32456,N_32613);
nand U33443 (N_33443,N_32269,N_32361);
nand U33444 (N_33444,N_32417,N_32073);
or U33445 (N_33445,N_32394,N_32941);
nor U33446 (N_33446,N_32172,N_32151);
and U33447 (N_33447,N_32763,N_32969);
and U33448 (N_33448,N_32911,N_32308);
nand U33449 (N_33449,N_32581,N_32583);
xnor U33450 (N_33450,N_32722,N_32810);
or U33451 (N_33451,N_32089,N_32248);
or U33452 (N_33452,N_32600,N_32285);
and U33453 (N_33453,N_32933,N_32017);
nand U33454 (N_33454,N_32737,N_32694);
or U33455 (N_33455,N_32104,N_32727);
nor U33456 (N_33456,N_32837,N_32907);
nand U33457 (N_33457,N_32612,N_32473);
and U33458 (N_33458,N_32544,N_32555);
xor U33459 (N_33459,N_32226,N_32716);
xnor U33460 (N_33460,N_32515,N_32604);
nand U33461 (N_33461,N_32898,N_32566);
or U33462 (N_33462,N_32743,N_32960);
or U33463 (N_33463,N_32606,N_32676);
and U33464 (N_33464,N_32118,N_32197);
and U33465 (N_33465,N_32966,N_32234);
nand U33466 (N_33466,N_32834,N_32770);
nor U33467 (N_33467,N_32905,N_32338);
xnor U33468 (N_33468,N_32301,N_32571);
or U33469 (N_33469,N_32296,N_32055);
and U33470 (N_33470,N_32506,N_32321);
nor U33471 (N_33471,N_32796,N_32380);
xor U33472 (N_33472,N_32974,N_32865);
nor U33473 (N_33473,N_32573,N_32520);
xor U33474 (N_33474,N_32353,N_32304);
and U33475 (N_33475,N_32275,N_32111);
nor U33476 (N_33476,N_32230,N_32449);
nor U33477 (N_33477,N_32631,N_32779);
nor U33478 (N_33478,N_32547,N_32883);
nand U33479 (N_33479,N_32820,N_32251);
and U33480 (N_33480,N_32097,N_32698);
or U33481 (N_33481,N_32080,N_32464);
xnor U33482 (N_33482,N_32889,N_32366);
and U33483 (N_33483,N_32656,N_32306);
nor U33484 (N_33484,N_32887,N_32996);
nor U33485 (N_33485,N_32025,N_32756);
and U33486 (N_33486,N_32263,N_32744);
or U33487 (N_33487,N_32682,N_32444);
nor U33488 (N_33488,N_32730,N_32345);
xor U33489 (N_33489,N_32598,N_32753);
nand U33490 (N_33490,N_32948,N_32677);
and U33491 (N_33491,N_32971,N_32253);
xor U33492 (N_33492,N_32202,N_32841);
or U33493 (N_33493,N_32901,N_32021);
nor U33494 (N_33494,N_32319,N_32182);
nor U33495 (N_33495,N_32881,N_32804);
xnor U33496 (N_33496,N_32836,N_32372);
nand U33497 (N_33497,N_32816,N_32311);
or U33498 (N_33498,N_32998,N_32144);
xor U33499 (N_33499,N_32483,N_32610);
xnor U33500 (N_33500,N_32006,N_32081);
nor U33501 (N_33501,N_32504,N_32913);
nand U33502 (N_33502,N_32436,N_32408);
or U33503 (N_33503,N_32647,N_32061);
nand U33504 (N_33504,N_32679,N_32867);
nor U33505 (N_33505,N_32375,N_32016);
or U33506 (N_33506,N_32693,N_32750);
nor U33507 (N_33507,N_32719,N_32923);
nand U33508 (N_33508,N_32131,N_32419);
or U33509 (N_33509,N_32735,N_32160);
nor U33510 (N_33510,N_32458,N_32102);
or U33511 (N_33511,N_32081,N_32799);
and U33512 (N_33512,N_32994,N_32520);
or U33513 (N_33513,N_32329,N_32503);
nand U33514 (N_33514,N_32423,N_32234);
and U33515 (N_33515,N_32494,N_32292);
nand U33516 (N_33516,N_32262,N_32832);
xnor U33517 (N_33517,N_32459,N_32452);
nand U33518 (N_33518,N_32007,N_32922);
or U33519 (N_33519,N_32753,N_32461);
and U33520 (N_33520,N_32885,N_32800);
nor U33521 (N_33521,N_32961,N_32770);
and U33522 (N_33522,N_32565,N_32513);
and U33523 (N_33523,N_32099,N_32587);
nor U33524 (N_33524,N_32974,N_32554);
nand U33525 (N_33525,N_32127,N_32120);
nor U33526 (N_33526,N_32447,N_32358);
nor U33527 (N_33527,N_32575,N_32531);
nand U33528 (N_33528,N_32123,N_32471);
xnor U33529 (N_33529,N_32657,N_32905);
and U33530 (N_33530,N_32061,N_32962);
xnor U33531 (N_33531,N_32489,N_32715);
and U33532 (N_33532,N_32516,N_32860);
nand U33533 (N_33533,N_32613,N_32189);
or U33534 (N_33534,N_32382,N_32712);
nor U33535 (N_33535,N_32658,N_32115);
nor U33536 (N_33536,N_32951,N_32981);
or U33537 (N_33537,N_32503,N_32799);
or U33538 (N_33538,N_32369,N_32057);
xor U33539 (N_33539,N_32445,N_32877);
and U33540 (N_33540,N_32819,N_32565);
nor U33541 (N_33541,N_32456,N_32879);
and U33542 (N_33542,N_32987,N_32857);
and U33543 (N_33543,N_32555,N_32975);
xnor U33544 (N_33544,N_32190,N_32646);
nand U33545 (N_33545,N_32710,N_32374);
nor U33546 (N_33546,N_32953,N_32112);
nand U33547 (N_33547,N_32877,N_32585);
and U33548 (N_33548,N_32588,N_32059);
xnor U33549 (N_33549,N_32206,N_32932);
nand U33550 (N_33550,N_32665,N_32187);
nand U33551 (N_33551,N_32533,N_32118);
nand U33552 (N_33552,N_32295,N_32458);
nor U33553 (N_33553,N_32524,N_32159);
nor U33554 (N_33554,N_32233,N_32527);
and U33555 (N_33555,N_32405,N_32385);
nor U33556 (N_33556,N_32665,N_32066);
nand U33557 (N_33557,N_32735,N_32329);
nor U33558 (N_33558,N_32936,N_32347);
nand U33559 (N_33559,N_32349,N_32051);
or U33560 (N_33560,N_32727,N_32057);
nor U33561 (N_33561,N_32634,N_32394);
nand U33562 (N_33562,N_32087,N_32717);
xnor U33563 (N_33563,N_32363,N_32249);
and U33564 (N_33564,N_32446,N_32645);
nand U33565 (N_33565,N_32728,N_32387);
nand U33566 (N_33566,N_32449,N_32108);
nand U33567 (N_33567,N_32270,N_32477);
nand U33568 (N_33568,N_32860,N_32798);
nor U33569 (N_33569,N_32305,N_32015);
nor U33570 (N_33570,N_32884,N_32606);
nor U33571 (N_33571,N_32772,N_32630);
or U33572 (N_33572,N_32179,N_32259);
or U33573 (N_33573,N_32287,N_32391);
nand U33574 (N_33574,N_32236,N_32593);
or U33575 (N_33575,N_32582,N_32446);
nand U33576 (N_33576,N_32465,N_32044);
or U33577 (N_33577,N_32160,N_32618);
and U33578 (N_33578,N_32732,N_32389);
xor U33579 (N_33579,N_32270,N_32891);
xor U33580 (N_33580,N_32024,N_32674);
nor U33581 (N_33581,N_32444,N_32154);
and U33582 (N_33582,N_32040,N_32718);
xnor U33583 (N_33583,N_32542,N_32829);
nand U33584 (N_33584,N_32123,N_32893);
nor U33585 (N_33585,N_32717,N_32562);
nor U33586 (N_33586,N_32957,N_32602);
or U33587 (N_33587,N_32558,N_32114);
and U33588 (N_33588,N_32806,N_32657);
or U33589 (N_33589,N_32516,N_32843);
nand U33590 (N_33590,N_32088,N_32247);
or U33591 (N_33591,N_32179,N_32688);
xor U33592 (N_33592,N_32419,N_32320);
and U33593 (N_33593,N_32393,N_32017);
xnor U33594 (N_33594,N_32435,N_32643);
xor U33595 (N_33595,N_32596,N_32457);
and U33596 (N_33596,N_32511,N_32129);
nand U33597 (N_33597,N_32475,N_32608);
nand U33598 (N_33598,N_32970,N_32542);
and U33599 (N_33599,N_32360,N_32128);
nor U33600 (N_33600,N_32744,N_32934);
nand U33601 (N_33601,N_32851,N_32099);
xnor U33602 (N_33602,N_32961,N_32711);
and U33603 (N_33603,N_32751,N_32179);
nand U33604 (N_33604,N_32841,N_32668);
nor U33605 (N_33605,N_32819,N_32271);
and U33606 (N_33606,N_32656,N_32349);
nand U33607 (N_33607,N_32790,N_32606);
xor U33608 (N_33608,N_32424,N_32429);
and U33609 (N_33609,N_32687,N_32628);
nand U33610 (N_33610,N_32813,N_32237);
nand U33611 (N_33611,N_32823,N_32895);
nand U33612 (N_33612,N_32095,N_32270);
or U33613 (N_33613,N_32544,N_32411);
xnor U33614 (N_33614,N_32955,N_32706);
nor U33615 (N_33615,N_32625,N_32929);
nor U33616 (N_33616,N_32025,N_32166);
xor U33617 (N_33617,N_32997,N_32185);
nand U33618 (N_33618,N_32945,N_32154);
and U33619 (N_33619,N_32798,N_32574);
or U33620 (N_33620,N_32082,N_32539);
nor U33621 (N_33621,N_32183,N_32031);
and U33622 (N_33622,N_32600,N_32387);
xnor U33623 (N_33623,N_32839,N_32280);
or U33624 (N_33624,N_32929,N_32441);
nand U33625 (N_33625,N_32137,N_32168);
xor U33626 (N_33626,N_32924,N_32435);
and U33627 (N_33627,N_32545,N_32955);
nor U33628 (N_33628,N_32057,N_32935);
xnor U33629 (N_33629,N_32240,N_32996);
nand U33630 (N_33630,N_32160,N_32185);
nand U33631 (N_33631,N_32499,N_32431);
nor U33632 (N_33632,N_32227,N_32364);
xnor U33633 (N_33633,N_32531,N_32806);
xor U33634 (N_33634,N_32826,N_32170);
nand U33635 (N_33635,N_32075,N_32567);
or U33636 (N_33636,N_32352,N_32810);
xnor U33637 (N_33637,N_32824,N_32768);
and U33638 (N_33638,N_32948,N_32855);
nand U33639 (N_33639,N_32703,N_32472);
xor U33640 (N_33640,N_32813,N_32909);
nor U33641 (N_33641,N_32851,N_32473);
nor U33642 (N_33642,N_32119,N_32567);
xor U33643 (N_33643,N_32185,N_32232);
nor U33644 (N_33644,N_32332,N_32325);
nor U33645 (N_33645,N_32510,N_32386);
nor U33646 (N_33646,N_32665,N_32822);
nand U33647 (N_33647,N_32128,N_32746);
nor U33648 (N_33648,N_32063,N_32358);
nor U33649 (N_33649,N_32261,N_32645);
xor U33650 (N_33650,N_32062,N_32065);
nor U33651 (N_33651,N_32559,N_32039);
and U33652 (N_33652,N_32126,N_32657);
nand U33653 (N_33653,N_32558,N_32238);
nand U33654 (N_33654,N_32565,N_32939);
and U33655 (N_33655,N_32574,N_32787);
and U33656 (N_33656,N_32234,N_32467);
nor U33657 (N_33657,N_32759,N_32797);
and U33658 (N_33658,N_32914,N_32809);
xnor U33659 (N_33659,N_32973,N_32982);
xnor U33660 (N_33660,N_32594,N_32518);
or U33661 (N_33661,N_32766,N_32383);
xnor U33662 (N_33662,N_32063,N_32262);
or U33663 (N_33663,N_32835,N_32703);
nor U33664 (N_33664,N_32296,N_32539);
xnor U33665 (N_33665,N_32652,N_32682);
nand U33666 (N_33666,N_32254,N_32573);
nor U33667 (N_33667,N_32574,N_32356);
nor U33668 (N_33668,N_32177,N_32768);
xor U33669 (N_33669,N_32526,N_32281);
nand U33670 (N_33670,N_32996,N_32164);
and U33671 (N_33671,N_32087,N_32468);
xnor U33672 (N_33672,N_32123,N_32450);
xnor U33673 (N_33673,N_32265,N_32325);
nor U33674 (N_33674,N_32006,N_32124);
nor U33675 (N_33675,N_32610,N_32920);
xnor U33676 (N_33676,N_32502,N_32441);
or U33677 (N_33677,N_32704,N_32423);
xor U33678 (N_33678,N_32404,N_32088);
nor U33679 (N_33679,N_32352,N_32892);
or U33680 (N_33680,N_32251,N_32033);
or U33681 (N_33681,N_32065,N_32878);
nand U33682 (N_33682,N_32999,N_32862);
xor U33683 (N_33683,N_32386,N_32878);
nand U33684 (N_33684,N_32362,N_32379);
or U33685 (N_33685,N_32615,N_32833);
nor U33686 (N_33686,N_32212,N_32332);
xor U33687 (N_33687,N_32523,N_32888);
nand U33688 (N_33688,N_32528,N_32131);
xnor U33689 (N_33689,N_32887,N_32653);
or U33690 (N_33690,N_32114,N_32659);
xor U33691 (N_33691,N_32675,N_32531);
xnor U33692 (N_33692,N_32923,N_32003);
xnor U33693 (N_33693,N_32367,N_32280);
nand U33694 (N_33694,N_32193,N_32392);
and U33695 (N_33695,N_32146,N_32940);
xnor U33696 (N_33696,N_32426,N_32436);
xor U33697 (N_33697,N_32002,N_32259);
nand U33698 (N_33698,N_32519,N_32377);
and U33699 (N_33699,N_32013,N_32495);
and U33700 (N_33700,N_32319,N_32974);
xnor U33701 (N_33701,N_32203,N_32092);
and U33702 (N_33702,N_32134,N_32052);
nand U33703 (N_33703,N_32185,N_32405);
xor U33704 (N_33704,N_32490,N_32258);
nor U33705 (N_33705,N_32497,N_32351);
and U33706 (N_33706,N_32269,N_32328);
or U33707 (N_33707,N_32151,N_32110);
or U33708 (N_33708,N_32405,N_32462);
nor U33709 (N_33709,N_32203,N_32341);
nand U33710 (N_33710,N_32748,N_32670);
nor U33711 (N_33711,N_32673,N_32169);
nand U33712 (N_33712,N_32138,N_32847);
and U33713 (N_33713,N_32740,N_32203);
or U33714 (N_33714,N_32013,N_32339);
and U33715 (N_33715,N_32962,N_32058);
and U33716 (N_33716,N_32508,N_32385);
and U33717 (N_33717,N_32789,N_32531);
xnor U33718 (N_33718,N_32369,N_32473);
or U33719 (N_33719,N_32740,N_32544);
nor U33720 (N_33720,N_32778,N_32310);
and U33721 (N_33721,N_32828,N_32277);
nand U33722 (N_33722,N_32546,N_32621);
nand U33723 (N_33723,N_32418,N_32449);
xor U33724 (N_33724,N_32673,N_32600);
and U33725 (N_33725,N_32265,N_32237);
nand U33726 (N_33726,N_32011,N_32121);
and U33727 (N_33727,N_32719,N_32055);
xor U33728 (N_33728,N_32770,N_32108);
or U33729 (N_33729,N_32719,N_32014);
and U33730 (N_33730,N_32930,N_32031);
nand U33731 (N_33731,N_32007,N_32255);
nand U33732 (N_33732,N_32675,N_32936);
nor U33733 (N_33733,N_32045,N_32326);
xor U33734 (N_33734,N_32610,N_32155);
or U33735 (N_33735,N_32639,N_32477);
and U33736 (N_33736,N_32092,N_32533);
nor U33737 (N_33737,N_32383,N_32203);
or U33738 (N_33738,N_32638,N_32227);
and U33739 (N_33739,N_32543,N_32486);
nand U33740 (N_33740,N_32667,N_32917);
xnor U33741 (N_33741,N_32980,N_32520);
xnor U33742 (N_33742,N_32215,N_32033);
and U33743 (N_33743,N_32554,N_32886);
nor U33744 (N_33744,N_32475,N_32612);
xor U33745 (N_33745,N_32246,N_32964);
and U33746 (N_33746,N_32324,N_32002);
or U33747 (N_33747,N_32466,N_32490);
nor U33748 (N_33748,N_32611,N_32815);
or U33749 (N_33749,N_32395,N_32284);
and U33750 (N_33750,N_32743,N_32883);
or U33751 (N_33751,N_32785,N_32656);
xnor U33752 (N_33752,N_32028,N_32634);
xnor U33753 (N_33753,N_32442,N_32963);
and U33754 (N_33754,N_32051,N_32381);
and U33755 (N_33755,N_32186,N_32852);
nor U33756 (N_33756,N_32564,N_32013);
or U33757 (N_33757,N_32929,N_32191);
nand U33758 (N_33758,N_32876,N_32932);
and U33759 (N_33759,N_32180,N_32016);
and U33760 (N_33760,N_32425,N_32879);
or U33761 (N_33761,N_32626,N_32131);
nor U33762 (N_33762,N_32821,N_32880);
or U33763 (N_33763,N_32972,N_32857);
and U33764 (N_33764,N_32856,N_32692);
and U33765 (N_33765,N_32718,N_32275);
xor U33766 (N_33766,N_32791,N_32795);
nor U33767 (N_33767,N_32304,N_32749);
and U33768 (N_33768,N_32347,N_32639);
nor U33769 (N_33769,N_32954,N_32848);
or U33770 (N_33770,N_32403,N_32850);
nor U33771 (N_33771,N_32713,N_32231);
xnor U33772 (N_33772,N_32313,N_32702);
or U33773 (N_33773,N_32855,N_32375);
or U33774 (N_33774,N_32912,N_32209);
nor U33775 (N_33775,N_32189,N_32933);
nand U33776 (N_33776,N_32776,N_32403);
nor U33777 (N_33777,N_32432,N_32908);
and U33778 (N_33778,N_32739,N_32412);
and U33779 (N_33779,N_32716,N_32087);
or U33780 (N_33780,N_32696,N_32199);
nand U33781 (N_33781,N_32129,N_32445);
and U33782 (N_33782,N_32573,N_32804);
nor U33783 (N_33783,N_32941,N_32971);
nor U33784 (N_33784,N_32431,N_32472);
xor U33785 (N_33785,N_32115,N_32804);
or U33786 (N_33786,N_32260,N_32159);
or U33787 (N_33787,N_32819,N_32668);
nor U33788 (N_33788,N_32011,N_32720);
and U33789 (N_33789,N_32364,N_32887);
nor U33790 (N_33790,N_32970,N_32642);
xnor U33791 (N_33791,N_32599,N_32811);
or U33792 (N_33792,N_32114,N_32326);
or U33793 (N_33793,N_32405,N_32176);
or U33794 (N_33794,N_32274,N_32581);
nor U33795 (N_33795,N_32506,N_32388);
nand U33796 (N_33796,N_32575,N_32183);
nand U33797 (N_33797,N_32024,N_32997);
or U33798 (N_33798,N_32631,N_32770);
nand U33799 (N_33799,N_32584,N_32897);
xnor U33800 (N_33800,N_32929,N_32920);
nor U33801 (N_33801,N_32313,N_32089);
xnor U33802 (N_33802,N_32397,N_32184);
and U33803 (N_33803,N_32977,N_32150);
and U33804 (N_33804,N_32730,N_32266);
xor U33805 (N_33805,N_32674,N_32056);
nor U33806 (N_33806,N_32484,N_32132);
nand U33807 (N_33807,N_32239,N_32254);
xnor U33808 (N_33808,N_32856,N_32549);
nand U33809 (N_33809,N_32955,N_32304);
xor U33810 (N_33810,N_32033,N_32439);
and U33811 (N_33811,N_32731,N_32039);
xnor U33812 (N_33812,N_32914,N_32345);
and U33813 (N_33813,N_32474,N_32548);
and U33814 (N_33814,N_32664,N_32289);
and U33815 (N_33815,N_32806,N_32710);
or U33816 (N_33816,N_32909,N_32500);
and U33817 (N_33817,N_32014,N_32254);
or U33818 (N_33818,N_32347,N_32037);
or U33819 (N_33819,N_32286,N_32953);
xnor U33820 (N_33820,N_32647,N_32409);
and U33821 (N_33821,N_32666,N_32374);
xnor U33822 (N_33822,N_32635,N_32317);
and U33823 (N_33823,N_32363,N_32739);
xor U33824 (N_33824,N_32465,N_32938);
or U33825 (N_33825,N_32797,N_32693);
xnor U33826 (N_33826,N_32483,N_32110);
nand U33827 (N_33827,N_32114,N_32248);
and U33828 (N_33828,N_32624,N_32158);
nand U33829 (N_33829,N_32252,N_32365);
and U33830 (N_33830,N_32458,N_32052);
xnor U33831 (N_33831,N_32917,N_32308);
nand U33832 (N_33832,N_32232,N_32865);
nor U33833 (N_33833,N_32064,N_32832);
nor U33834 (N_33834,N_32438,N_32032);
nor U33835 (N_33835,N_32711,N_32234);
nand U33836 (N_33836,N_32401,N_32732);
xnor U33837 (N_33837,N_32282,N_32679);
nor U33838 (N_33838,N_32165,N_32259);
nand U33839 (N_33839,N_32605,N_32442);
nor U33840 (N_33840,N_32899,N_32152);
nor U33841 (N_33841,N_32097,N_32548);
or U33842 (N_33842,N_32680,N_32409);
or U33843 (N_33843,N_32191,N_32452);
nor U33844 (N_33844,N_32461,N_32551);
or U33845 (N_33845,N_32492,N_32663);
and U33846 (N_33846,N_32080,N_32220);
or U33847 (N_33847,N_32184,N_32876);
nand U33848 (N_33848,N_32592,N_32307);
xnor U33849 (N_33849,N_32181,N_32182);
xnor U33850 (N_33850,N_32750,N_32781);
and U33851 (N_33851,N_32400,N_32099);
nand U33852 (N_33852,N_32138,N_32427);
nor U33853 (N_33853,N_32221,N_32468);
nand U33854 (N_33854,N_32162,N_32697);
xor U33855 (N_33855,N_32779,N_32978);
and U33856 (N_33856,N_32706,N_32560);
nand U33857 (N_33857,N_32708,N_32842);
nor U33858 (N_33858,N_32949,N_32813);
nor U33859 (N_33859,N_32916,N_32501);
nor U33860 (N_33860,N_32224,N_32983);
nor U33861 (N_33861,N_32212,N_32762);
and U33862 (N_33862,N_32904,N_32016);
xnor U33863 (N_33863,N_32642,N_32163);
xor U33864 (N_33864,N_32650,N_32950);
xor U33865 (N_33865,N_32143,N_32957);
or U33866 (N_33866,N_32741,N_32594);
and U33867 (N_33867,N_32992,N_32393);
nor U33868 (N_33868,N_32805,N_32783);
nand U33869 (N_33869,N_32105,N_32329);
and U33870 (N_33870,N_32831,N_32929);
xnor U33871 (N_33871,N_32665,N_32900);
nand U33872 (N_33872,N_32441,N_32808);
nand U33873 (N_33873,N_32821,N_32139);
or U33874 (N_33874,N_32477,N_32522);
nor U33875 (N_33875,N_32296,N_32996);
xor U33876 (N_33876,N_32382,N_32416);
and U33877 (N_33877,N_32286,N_32514);
nand U33878 (N_33878,N_32544,N_32934);
and U33879 (N_33879,N_32388,N_32002);
nor U33880 (N_33880,N_32015,N_32550);
xnor U33881 (N_33881,N_32356,N_32051);
nor U33882 (N_33882,N_32042,N_32719);
nor U33883 (N_33883,N_32054,N_32866);
or U33884 (N_33884,N_32740,N_32463);
or U33885 (N_33885,N_32645,N_32312);
or U33886 (N_33886,N_32985,N_32821);
nor U33887 (N_33887,N_32712,N_32757);
and U33888 (N_33888,N_32542,N_32964);
nand U33889 (N_33889,N_32778,N_32515);
nand U33890 (N_33890,N_32391,N_32717);
nor U33891 (N_33891,N_32685,N_32676);
and U33892 (N_33892,N_32819,N_32453);
and U33893 (N_33893,N_32593,N_32244);
or U33894 (N_33894,N_32185,N_32744);
xor U33895 (N_33895,N_32783,N_32953);
and U33896 (N_33896,N_32386,N_32005);
xor U33897 (N_33897,N_32067,N_32181);
nand U33898 (N_33898,N_32006,N_32058);
and U33899 (N_33899,N_32070,N_32212);
or U33900 (N_33900,N_32830,N_32150);
nor U33901 (N_33901,N_32275,N_32121);
or U33902 (N_33902,N_32228,N_32719);
nand U33903 (N_33903,N_32161,N_32404);
xnor U33904 (N_33904,N_32696,N_32677);
nand U33905 (N_33905,N_32136,N_32424);
nand U33906 (N_33906,N_32269,N_32166);
and U33907 (N_33907,N_32389,N_32664);
or U33908 (N_33908,N_32527,N_32537);
nor U33909 (N_33909,N_32273,N_32769);
or U33910 (N_33910,N_32056,N_32143);
or U33911 (N_33911,N_32514,N_32274);
nor U33912 (N_33912,N_32381,N_32722);
and U33913 (N_33913,N_32823,N_32958);
and U33914 (N_33914,N_32479,N_32842);
and U33915 (N_33915,N_32919,N_32117);
and U33916 (N_33916,N_32177,N_32257);
and U33917 (N_33917,N_32179,N_32057);
nor U33918 (N_33918,N_32223,N_32931);
nor U33919 (N_33919,N_32749,N_32711);
nor U33920 (N_33920,N_32068,N_32585);
xor U33921 (N_33921,N_32503,N_32655);
xnor U33922 (N_33922,N_32014,N_32214);
and U33923 (N_33923,N_32803,N_32283);
xor U33924 (N_33924,N_32639,N_32476);
xor U33925 (N_33925,N_32625,N_32044);
nor U33926 (N_33926,N_32337,N_32084);
and U33927 (N_33927,N_32424,N_32787);
xor U33928 (N_33928,N_32501,N_32854);
and U33929 (N_33929,N_32067,N_32363);
or U33930 (N_33930,N_32674,N_32315);
and U33931 (N_33931,N_32239,N_32788);
and U33932 (N_33932,N_32956,N_32267);
xnor U33933 (N_33933,N_32673,N_32065);
xnor U33934 (N_33934,N_32938,N_32986);
nor U33935 (N_33935,N_32336,N_32289);
or U33936 (N_33936,N_32321,N_32416);
nand U33937 (N_33937,N_32164,N_32745);
nor U33938 (N_33938,N_32265,N_32025);
nor U33939 (N_33939,N_32936,N_32142);
nor U33940 (N_33940,N_32494,N_32957);
or U33941 (N_33941,N_32346,N_32139);
nand U33942 (N_33942,N_32508,N_32953);
and U33943 (N_33943,N_32086,N_32694);
nor U33944 (N_33944,N_32397,N_32662);
or U33945 (N_33945,N_32877,N_32060);
nand U33946 (N_33946,N_32262,N_32372);
nand U33947 (N_33947,N_32410,N_32348);
nand U33948 (N_33948,N_32116,N_32707);
and U33949 (N_33949,N_32146,N_32393);
nand U33950 (N_33950,N_32069,N_32232);
xor U33951 (N_33951,N_32428,N_32964);
or U33952 (N_33952,N_32151,N_32849);
and U33953 (N_33953,N_32409,N_32402);
nor U33954 (N_33954,N_32858,N_32652);
and U33955 (N_33955,N_32761,N_32394);
or U33956 (N_33956,N_32969,N_32520);
xnor U33957 (N_33957,N_32791,N_32153);
and U33958 (N_33958,N_32292,N_32484);
nand U33959 (N_33959,N_32881,N_32260);
and U33960 (N_33960,N_32529,N_32820);
xnor U33961 (N_33961,N_32907,N_32367);
or U33962 (N_33962,N_32973,N_32365);
nand U33963 (N_33963,N_32249,N_32295);
xnor U33964 (N_33964,N_32666,N_32958);
nor U33965 (N_33965,N_32628,N_32716);
xor U33966 (N_33966,N_32039,N_32963);
nand U33967 (N_33967,N_32424,N_32942);
xor U33968 (N_33968,N_32507,N_32234);
nor U33969 (N_33969,N_32357,N_32642);
nor U33970 (N_33970,N_32293,N_32417);
xor U33971 (N_33971,N_32318,N_32129);
or U33972 (N_33972,N_32286,N_32988);
or U33973 (N_33973,N_32312,N_32794);
or U33974 (N_33974,N_32274,N_32357);
and U33975 (N_33975,N_32256,N_32840);
and U33976 (N_33976,N_32680,N_32863);
or U33977 (N_33977,N_32675,N_32036);
xnor U33978 (N_33978,N_32864,N_32932);
nor U33979 (N_33979,N_32460,N_32872);
nand U33980 (N_33980,N_32472,N_32630);
nor U33981 (N_33981,N_32843,N_32989);
nor U33982 (N_33982,N_32599,N_32998);
nand U33983 (N_33983,N_32426,N_32487);
and U33984 (N_33984,N_32671,N_32376);
and U33985 (N_33985,N_32532,N_32561);
nand U33986 (N_33986,N_32520,N_32187);
nor U33987 (N_33987,N_32028,N_32055);
or U33988 (N_33988,N_32998,N_32042);
or U33989 (N_33989,N_32898,N_32208);
xor U33990 (N_33990,N_32757,N_32069);
and U33991 (N_33991,N_32211,N_32808);
xnor U33992 (N_33992,N_32107,N_32936);
or U33993 (N_33993,N_32928,N_32261);
nand U33994 (N_33994,N_32928,N_32063);
nor U33995 (N_33995,N_32372,N_32275);
and U33996 (N_33996,N_32403,N_32566);
nor U33997 (N_33997,N_32006,N_32013);
nand U33998 (N_33998,N_32346,N_32467);
nand U33999 (N_33999,N_32165,N_32628);
nor U34000 (N_34000,N_33370,N_33369);
xnor U34001 (N_34001,N_33852,N_33669);
nor U34002 (N_34002,N_33440,N_33076);
or U34003 (N_34003,N_33567,N_33391);
and U34004 (N_34004,N_33051,N_33394);
nand U34005 (N_34005,N_33281,N_33138);
nand U34006 (N_34006,N_33916,N_33870);
nand U34007 (N_34007,N_33271,N_33697);
nor U34008 (N_34008,N_33695,N_33764);
or U34009 (N_34009,N_33667,N_33320);
or U34010 (N_34010,N_33274,N_33861);
nand U34011 (N_34011,N_33933,N_33278);
or U34012 (N_34012,N_33867,N_33902);
or U34013 (N_34013,N_33720,N_33186);
nor U34014 (N_34014,N_33445,N_33666);
nand U34015 (N_34015,N_33649,N_33079);
nor U34016 (N_34016,N_33622,N_33664);
nor U34017 (N_34017,N_33090,N_33277);
or U34018 (N_34018,N_33755,N_33737);
xor U34019 (N_34019,N_33127,N_33419);
nand U34020 (N_34020,N_33890,N_33174);
xor U34021 (N_34021,N_33789,N_33312);
xor U34022 (N_34022,N_33485,N_33774);
or U34023 (N_34023,N_33516,N_33395);
or U34024 (N_34024,N_33824,N_33712);
and U34025 (N_34025,N_33604,N_33122);
or U34026 (N_34026,N_33941,N_33055);
xor U34027 (N_34027,N_33182,N_33155);
nor U34028 (N_34028,N_33676,N_33771);
nor U34029 (N_34029,N_33524,N_33926);
and U34030 (N_34030,N_33725,N_33619);
and U34031 (N_34031,N_33585,N_33678);
and U34032 (N_34032,N_33806,N_33629);
nor U34033 (N_34033,N_33157,N_33814);
and U34034 (N_34034,N_33692,N_33504);
nor U34035 (N_34035,N_33473,N_33661);
nand U34036 (N_34036,N_33810,N_33544);
nor U34037 (N_34037,N_33466,N_33531);
or U34038 (N_34038,N_33995,N_33048);
and U34039 (N_34039,N_33860,N_33168);
nand U34040 (N_34040,N_33191,N_33791);
nand U34041 (N_34041,N_33235,N_33548);
and U34042 (N_34042,N_33602,N_33406);
and U34043 (N_34043,N_33547,N_33074);
xor U34044 (N_34044,N_33868,N_33259);
xor U34045 (N_34045,N_33311,N_33131);
xnor U34046 (N_34046,N_33533,N_33361);
and U34047 (N_34047,N_33433,N_33372);
nor U34048 (N_34048,N_33269,N_33951);
nor U34049 (N_34049,N_33637,N_33097);
or U34050 (N_34050,N_33804,N_33309);
xor U34051 (N_34051,N_33875,N_33173);
or U34052 (N_34052,N_33184,N_33889);
nor U34053 (N_34053,N_33794,N_33895);
nand U34054 (N_34054,N_33593,N_33257);
or U34055 (N_34055,N_33096,N_33244);
and U34056 (N_34056,N_33333,N_33210);
nor U34057 (N_34057,N_33701,N_33285);
nor U34058 (N_34058,N_33813,N_33935);
xnor U34059 (N_34059,N_33782,N_33106);
or U34060 (N_34060,N_33015,N_33592);
xor U34061 (N_34061,N_33345,N_33300);
nor U34062 (N_34062,N_33389,N_33657);
xnor U34063 (N_34063,N_33520,N_33289);
xnor U34064 (N_34064,N_33971,N_33439);
or U34065 (N_34065,N_33021,N_33359);
xnor U34066 (N_34066,N_33606,N_33491);
and U34067 (N_34067,N_33882,N_33011);
nand U34068 (N_34068,N_33343,N_33167);
or U34069 (N_34069,N_33338,N_33821);
nor U34070 (N_34070,N_33843,N_33348);
and U34071 (N_34071,N_33261,N_33352);
or U34072 (N_34072,N_33085,N_33213);
and U34073 (N_34073,N_33750,N_33723);
nor U34074 (N_34074,N_33613,N_33552);
xor U34075 (N_34075,N_33883,N_33736);
nor U34076 (N_34076,N_33724,N_33077);
and U34077 (N_34077,N_33022,N_33237);
nand U34078 (N_34078,N_33660,N_33068);
nand U34079 (N_34079,N_33912,N_33741);
or U34080 (N_34080,N_33205,N_33297);
and U34081 (N_34081,N_33508,N_33961);
or U34082 (N_34082,N_33831,N_33233);
nor U34083 (N_34083,N_33337,N_33950);
and U34084 (N_34084,N_33087,N_33621);
nor U34085 (N_34085,N_33994,N_33521);
and U34086 (N_34086,N_33020,N_33584);
xor U34087 (N_34087,N_33132,N_33542);
and U34088 (N_34088,N_33137,N_33790);
or U34089 (N_34089,N_33012,N_33116);
and U34090 (N_34090,N_33967,N_33047);
or U34091 (N_34091,N_33071,N_33492);
nand U34092 (N_34092,N_33973,N_33702);
or U34093 (N_34093,N_33714,N_33735);
or U34094 (N_34094,N_33513,N_33416);
and U34095 (N_34095,N_33907,N_33420);
nand U34096 (N_34096,N_33234,N_33566);
nand U34097 (N_34097,N_33962,N_33927);
or U34098 (N_34098,N_33769,N_33523);
xor U34099 (N_34099,N_33110,N_33545);
xnor U34100 (N_34100,N_33553,N_33862);
nand U34101 (N_34101,N_33105,N_33380);
xnor U34102 (N_34102,N_33054,N_33284);
and U34103 (N_34103,N_33581,N_33934);
nor U34104 (N_34104,N_33064,N_33917);
nand U34105 (N_34105,N_33480,N_33829);
or U34106 (N_34106,N_33826,N_33160);
and U34107 (N_34107,N_33373,N_33823);
xor U34108 (N_34108,N_33019,N_33031);
xnor U34109 (N_34109,N_33412,N_33392);
or U34110 (N_34110,N_33733,N_33872);
nand U34111 (N_34111,N_33476,N_33665);
xnor U34112 (N_34112,N_33554,N_33303);
or U34113 (N_34113,N_33564,N_33005);
or U34114 (N_34114,N_33422,N_33827);
xnor U34115 (N_34115,N_33414,N_33802);
nor U34116 (N_34116,N_33819,N_33878);
xnor U34117 (N_34117,N_33832,N_33267);
and U34118 (N_34118,N_33909,N_33757);
xor U34119 (N_34119,N_33753,N_33717);
xor U34120 (N_34120,N_33130,N_33080);
nand U34121 (N_34121,N_33589,N_33828);
and U34122 (N_34122,N_33401,N_33408);
xnor U34123 (N_34123,N_33728,N_33456);
xnor U34124 (N_34124,N_33441,N_33428);
nor U34125 (N_34125,N_33921,N_33196);
or U34126 (N_34126,N_33302,N_33838);
and U34127 (N_34127,N_33276,N_33029);
or U34128 (N_34128,N_33488,N_33586);
xor U34129 (N_34129,N_33915,N_33314);
or U34130 (N_34130,N_33652,N_33510);
nor U34131 (N_34131,N_33039,N_33481);
or U34132 (N_34132,N_33243,N_33207);
nor U34133 (N_34133,N_33221,N_33245);
nand U34134 (N_34134,N_33760,N_33742);
nor U34135 (N_34135,N_33651,N_33086);
or U34136 (N_34136,N_33318,N_33025);
and U34137 (N_34137,N_33159,N_33163);
or U34138 (N_34138,N_33407,N_33474);
and U34139 (N_34139,N_33193,N_33987);
xor U34140 (N_34140,N_33900,N_33966);
nor U34141 (N_34141,N_33968,N_33228);
or U34142 (N_34142,N_33161,N_33084);
xnor U34143 (N_34143,N_33489,N_33135);
xor U34144 (N_34144,N_33842,N_33885);
xnor U34145 (N_34145,N_33255,N_33363);
nor U34146 (N_34146,N_33177,N_33913);
or U34147 (N_34147,N_33282,N_33938);
xnor U34148 (N_34148,N_33594,N_33470);
nor U34149 (N_34149,N_33793,N_33214);
and U34150 (N_34150,N_33376,N_33156);
or U34151 (N_34151,N_33706,N_33448);
or U34152 (N_34152,N_33464,N_33129);
nand U34153 (N_34153,N_33579,N_33436);
xor U34154 (N_34154,N_33431,N_33426);
xor U34155 (N_34155,N_33319,N_33784);
xor U34156 (N_34156,N_33185,N_33527);
and U34157 (N_34157,N_33266,N_33946);
nor U34158 (N_34158,N_33743,N_33822);
nand U34159 (N_34159,N_33236,N_33601);
nor U34160 (N_34160,N_33050,N_33618);
or U34161 (N_34161,N_33796,N_33299);
xnor U34162 (N_34162,N_33707,N_33858);
xnor U34163 (N_34163,N_33328,N_33744);
or U34164 (N_34164,N_33176,N_33415);
or U34165 (N_34165,N_33010,N_33937);
or U34166 (N_34166,N_33180,N_33770);
and U34167 (N_34167,N_33324,N_33151);
and U34168 (N_34168,N_33242,N_33203);
or U34169 (N_34169,N_33730,N_33374);
or U34170 (N_34170,N_33171,N_33482);
xnor U34171 (N_34171,N_33381,N_33710);
nor U34172 (N_34172,N_33249,N_33053);
xor U34173 (N_34173,N_33911,N_33857);
nand U34174 (N_34174,N_33538,N_33444);
nor U34175 (N_34175,N_33647,N_33874);
nor U34176 (N_34176,N_33014,N_33451);
nor U34177 (N_34177,N_33797,N_33959);
or U34178 (N_34178,N_33356,N_33632);
nand U34179 (N_34179,N_33475,N_33816);
xor U34180 (N_34180,N_33434,N_33779);
xor U34181 (N_34181,N_33449,N_33202);
and U34182 (N_34182,N_33638,N_33777);
and U34183 (N_34183,N_33030,N_33317);
nand U34184 (N_34184,N_33294,N_33033);
xor U34185 (N_34185,N_33776,N_33371);
and U34186 (N_34186,N_33919,N_33027);
and U34187 (N_34187,N_33901,N_33837);
nand U34188 (N_34188,N_33026,N_33859);
xnor U34189 (N_34189,N_33037,N_33896);
nand U34190 (N_34190,N_33227,N_33974);
nand U34191 (N_34191,N_33204,N_33438);
or U34192 (N_34192,N_33910,N_33220);
nand U34193 (N_34193,N_33305,N_33229);
or U34194 (N_34194,N_33061,N_33943);
or U34195 (N_34195,N_33700,N_33673);
or U34196 (N_34196,N_33698,N_33898);
nand U34197 (N_34197,N_33198,N_33625);
xor U34198 (N_34198,N_33687,N_33947);
or U34199 (N_34199,N_33323,N_33975);
xor U34200 (N_34200,N_33384,N_33756);
or U34201 (N_34201,N_33864,N_33032);
and U34202 (N_34202,N_33383,N_33158);
xnor U34203 (N_34203,N_33344,N_33888);
nor U34204 (N_34204,N_33082,N_33002);
nor U34205 (N_34205,N_33607,N_33939);
and U34206 (N_34206,N_33217,N_33672);
xor U34207 (N_34207,N_33248,N_33931);
and U34208 (N_34208,N_33653,N_33003);
or U34209 (N_34209,N_33863,N_33216);
xnor U34210 (N_34210,N_33886,N_33590);
xnor U34211 (N_34211,N_33711,N_33405);
or U34212 (N_34212,N_33494,N_33550);
nand U34213 (N_34213,N_33583,N_33949);
xnor U34214 (N_34214,N_33803,N_33427);
nand U34215 (N_34215,N_33410,N_33360);
or U34216 (N_34216,N_33224,N_33335);
nand U34217 (N_34217,N_33630,N_33091);
nand U34218 (N_34218,N_33468,N_33238);
nand U34219 (N_34219,N_33460,N_33016);
nor U34220 (N_34220,N_33979,N_33529);
xnor U34221 (N_34221,N_33930,N_33659);
or U34222 (N_34222,N_33102,N_33377);
nor U34223 (N_34223,N_33845,N_33316);
xnor U34224 (N_34224,N_33693,N_33873);
and U34225 (N_34225,N_33346,N_33801);
and U34226 (N_34226,N_33708,N_33140);
nor U34227 (N_34227,N_33500,N_33189);
and U34228 (N_34228,N_33611,N_33293);
nand U34229 (N_34229,N_33866,N_33833);
nand U34230 (N_34230,N_33848,N_33049);
and U34231 (N_34231,N_33250,N_33972);
nor U34232 (N_34232,N_33617,N_33313);
and U34233 (N_34233,N_33932,N_33557);
nand U34234 (N_34234,N_33634,N_33515);
nor U34235 (N_34235,N_33639,N_33070);
and U34236 (N_34236,N_33169,N_33499);
xor U34237 (N_34237,N_33201,N_33713);
xnor U34238 (N_34238,N_33081,N_33800);
xor U34239 (N_34239,N_33009,N_33128);
and U34240 (N_34240,N_33175,N_33417);
nor U34241 (N_34241,N_33246,N_33479);
or U34242 (N_34242,N_33597,N_33413);
or U34243 (N_34243,N_33549,N_33892);
nand U34244 (N_34244,N_33679,N_33881);
xor U34245 (N_34245,N_33040,N_33044);
nor U34246 (N_34246,N_33501,N_33219);
and U34247 (N_34247,N_33880,N_33614);
nand U34248 (N_34248,N_33256,N_33336);
xor U34249 (N_34249,N_33462,N_33561);
nand U34250 (N_34250,N_33268,N_33654);
xor U34251 (N_34251,N_33688,N_33871);
and U34252 (N_34252,N_33326,N_33108);
or U34253 (N_34253,N_33435,N_33512);
or U34254 (N_34254,N_33808,N_33763);
xor U34255 (N_34255,N_33088,N_33283);
or U34256 (N_34256,N_33365,N_33573);
and U34257 (N_34257,N_33350,N_33452);
xnor U34258 (N_34258,N_33605,N_33188);
nand U34259 (N_34259,N_33310,N_33985);
nor U34260 (N_34260,N_33378,N_33855);
or U34261 (N_34261,N_33980,N_33197);
nor U34262 (N_34262,N_33626,N_33258);
nand U34263 (N_34263,N_33825,N_33555);
or U34264 (N_34264,N_33904,N_33556);
xor U34265 (N_34265,N_33572,N_33840);
xnor U34266 (N_34266,N_33989,N_33656);
or U34267 (N_34267,N_33785,N_33696);
nor U34268 (N_34268,N_33853,N_33341);
and U34269 (N_34269,N_33423,N_33298);
and U34270 (N_34270,N_33208,N_33493);
or U34271 (N_34271,N_33390,N_33856);
or U34272 (N_34272,N_33477,N_33920);
and U34273 (N_34273,N_33820,N_33006);
or U34274 (N_34274,N_33388,N_33113);
xor U34275 (N_34275,N_33056,N_33307);
nor U34276 (N_34276,N_33152,N_33729);
xor U34277 (N_34277,N_33775,N_33600);
and U34278 (N_34278,N_33537,N_33092);
and U34279 (N_34279,N_33690,N_33612);
or U34280 (N_34280,N_33633,N_33628);
or U34281 (N_34281,N_33458,N_33036);
and U34282 (N_34282,N_33746,N_33535);
nor U34283 (N_34283,N_33008,N_33970);
nor U34284 (N_34284,N_33063,N_33170);
nor U34285 (N_34285,N_33580,N_33954);
nand U34286 (N_34286,N_33603,N_33674);
nor U34287 (N_34287,N_33306,N_33936);
or U34288 (N_34288,N_33778,N_33211);
and U34289 (N_34289,N_33263,N_33929);
nor U34290 (N_34290,N_33773,N_33694);
nand U34291 (N_34291,N_33432,N_33045);
nor U34292 (N_34292,N_33984,N_33945);
nor U34293 (N_34293,N_33334,N_33286);
or U34294 (N_34294,N_33809,N_33799);
or U34295 (N_34295,N_33540,N_33719);
nor U34296 (N_34296,N_33588,N_33503);
nor U34297 (N_34297,N_33918,N_33232);
nand U34298 (N_34298,N_33218,N_33172);
nand U34299 (N_34299,N_33264,N_33215);
xor U34300 (N_34300,N_33490,N_33836);
nand U34301 (N_34301,N_33528,N_33965);
or U34302 (N_34302,N_33849,N_33745);
or U34303 (N_34303,N_33686,N_33339);
and U34304 (N_34304,N_33368,N_33705);
and U34305 (N_34305,N_33754,N_33715);
xor U34306 (N_34306,N_33519,N_33366);
or U34307 (N_34307,N_33766,N_33691);
xnor U34308 (N_34308,N_33495,N_33418);
and U34309 (N_34309,N_33469,N_33834);
nor U34310 (N_34310,N_33768,N_33891);
or U34311 (N_34311,N_33587,N_33367);
or U34312 (N_34312,N_33141,N_33330);
and U34313 (N_34313,N_33496,N_33807);
or U34314 (N_34314,N_33498,N_33685);
or U34315 (N_34315,N_33484,N_33627);
and U34316 (N_34316,N_33304,N_33999);
nand U34317 (N_34317,N_33532,N_33017);
nor U34318 (N_34318,N_33465,N_33677);
nor U34319 (N_34319,N_33844,N_33123);
xor U34320 (N_34320,N_33409,N_33903);
or U34321 (N_34321,N_33992,N_33578);
and U34322 (N_34322,N_33905,N_33065);
nor U34323 (N_34323,N_33575,N_33375);
or U34324 (N_34324,N_33199,N_33740);
and U34325 (N_34325,N_33212,N_33718);
xor U34326 (N_34326,N_33075,N_33570);
or U34327 (N_34327,N_33908,N_33024);
nor U34328 (N_34328,N_33223,N_33925);
or U34329 (N_34329,N_33977,N_33393);
nor U34330 (N_34330,N_33650,N_33013);
and U34331 (N_34331,N_33506,N_33897);
xor U34332 (N_34332,N_33164,N_33559);
and U34333 (N_34333,N_33379,N_33640);
nor U34334 (N_34334,N_33430,N_33192);
xnor U34335 (N_34335,N_33231,N_33471);
nand U34336 (N_34336,N_33681,N_33960);
or U34337 (N_34337,N_33209,N_33877);
nand U34338 (N_34338,N_33689,N_33400);
or U34339 (N_34339,N_33067,N_33560);
nor U34340 (N_34340,N_33150,N_33442);
or U34341 (N_34341,N_33525,N_33599);
xor U34342 (N_34342,N_33502,N_33507);
xnor U34343 (N_34343,N_33663,N_33200);
nor U34344 (N_34344,N_33812,N_33062);
nor U34345 (N_34345,N_33631,N_33758);
and U34346 (N_34346,N_33709,N_33112);
or U34347 (N_34347,N_33028,N_33331);
xor U34348 (N_34348,N_33162,N_33069);
and U34349 (N_34349,N_33817,N_33922);
nor U34350 (N_34350,N_33254,N_33230);
xor U34351 (N_34351,N_33906,N_33385);
and U34352 (N_34352,N_33118,N_33099);
xor U34353 (N_34353,N_33120,N_33315);
or U34354 (N_34354,N_33991,N_33787);
or U34355 (N_34355,N_33115,N_33762);
nor U34356 (N_34356,N_33225,N_33035);
nand U34357 (N_34357,N_33830,N_33624);
nor U34358 (N_34358,N_33788,N_33792);
xnor U34359 (N_34359,N_33990,N_33247);
xor U34360 (N_34360,N_33955,N_33292);
or U34361 (N_34361,N_33124,N_33342);
and U34362 (N_34362,N_33461,N_33321);
xor U34363 (N_34363,N_33329,N_33576);
or U34364 (N_34364,N_33958,N_33924);
nand U34365 (N_34365,N_33668,N_33957);
nand U34366 (N_34366,N_33239,N_33783);
nor U34367 (N_34367,N_33983,N_33811);
or U34368 (N_34368,N_33386,N_33530);
and U34369 (N_34369,N_33781,N_33747);
nor U34370 (N_34370,N_33398,N_33403);
nor U34371 (N_34371,N_33704,N_33125);
or U34372 (N_34372,N_33057,N_33988);
nand U34373 (N_34373,N_33038,N_33662);
or U34374 (N_34374,N_33450,N_33457);
nand U34375 (N_34375,N_33732,N_33683);
nand U34376 (N_34376,N_33699,N_33646);
nand U34377 (N_34377,N_33001,N_33739);
xor U34378 (N_34378,N_33382,N_33396);
nand U34379 (N_34379,N_33463,N_33487);
xnor U34380 (N_34380,N_33424,N_33635);
nand U34381 (N_34381,N_33308,N_33133);
nand U34382 (N_34382,N_33265,N_33928);
and U34383 (N_34383,N_33357,N_33147);
and U34384 (N_34384,N_33643,N_33296);
xnor U34385 (N_34385,N_33952,N_33749);
nand U34386 (N_34386,N_33060,N_33887);
nor U34387 (N_34387,N_33478,N_33000);
or U34388 (N_34388,N_33805,N_33251);
and U34389 (N_34389,N_33145,N_33884);
and U34390 (N_34390,N_33981,N_33759);
or U34391 (N_34391,N_33953,N_33121);
and U34392 (N_34392,N_33518,N_33565);
or U34393 (N_34393,N_33194,N_33486);
and U34394 (N_34394,N_33675,N_33066);
nand U34395 (N_34395,N_33222,N_33165);
nand U34396 (N_34396,N_33976,N_33986);
nor U34397 (N_34397,N_33322,N_33114);
nand U34398 (N_34398,N_33948,N_33563);
and U34399 (N_34399,N_33574,N_33095);
and U34400 (N_34400,N_33273,N_33358);
or U34401 (N_34401,N_33332,N_33636);
nand U34402 (N_34402,N_33731,N_33093);
and U34403 (N_34403,N_33136,N_33997);
nand U34404 (N_34404,N_33734,N_33149);
and U34405 (N_34405,N_33998,N_33364);
nand U34406 (N_34406,N_33046,N_33680);
nand U34407 (N_34407,N_33648,N_33272);
and U34408 (N_34408,N_33964,N_33658);
or U34409 (N_34409,N_33052,N_33671);
or U34410 (N_34410,N_33854,N_33072);
xnor U34411 (N_34411,N_33582,N_33101);
nand U34412 (N_34412,N_33351,N_33327);
and U34413 (N_34413,N_33421,N_33569);
xnor U34414 (N_34414,N_33134,N_33655);
nor U34415 (N_34415,N_33241,N_33270);
xor U34416 (N_34416,N_33818,N_33253);
or U34417 (N_34417,N_33616,N_33059);
xor U34418 (N_34418,N_33682,N_33847);
nor U34419 (N_34419,N_33761,N_33726);
and U34420 (N_34420,N_33262,N_33411);
nand U34421 (N_34421,N_33509,N_33869);
or U34422 (N_34422,N_33083,N_33260);
nand U34423 (N_34423,N_33178,N_33534);
xor U34424 (N_34424,N_33539,N_33993);
nand U34425 (N_34425,N_33146,N_33923);
xnor U34426 (N_34426,N_33429,N_33103);
or U34427 (N_34427,N_33287,N_33595);
nor U34428 (N_34428,N_33543,N_33455);
and U34429 (N_34429,N_33835,N_33541);
and U34430 (N_34430,N_33404,N_33148);
or U34431 (N_34431,N_33645,N_33179);
or U34432 (N_34432,N_33577,N_33841);
nor U34433 (N_34433,N_33511,N_33183);
or U34434 (N_34434,N_33982,N_33004);
nand U34435 (N_34435,N_33117,N_33139);
nand U34436 (N_34436,N_33362,N_33944);
and U34437 (N_34437,N_33684,N_33111);
or U34438 (N_34438,N_33893,N_33459);
nand U34439 (N_34439,N_33153,N_33591);
nor U34440 (N_34440,N_33240,N_33325);
xnor U34441 (N_34441,N_33772,N_33166);
nor U34442 (N_34442,N_33722,N_33107);
or U34443 (N_34443,N_33143,N_33279);
xor U34444 (N_34444,N_33615,N_33126);
xnor U34445 (N_34445,N_33446,N_33399);
xor U34446 (N_34446,N_33397,N_33914);
and U34447 (N_34447,N_33522,N_33252);
and U34448 (N_34448,N_33568,N_33098);
nand U34449 (N_34449,N_33144,N_33623);
nor U34450 (N_34450,N_33620,N_33598);
nand U34451 (N_34451,N_33876,N_33558);
nand U34452 (N_34452,N_33454,N_33109);
and U34453 (N_34453,N_33018,N_33041);
nand U34454 (N_34454,N_33447,N_33963);
nand U34455 (N_34455,N_33355,N_33517);
xor U34456 (N_34456,N_33942,N_33738);
xor U34457 (N_34457,N_33187,N_33894);
nand U34458 (N_34458,N_33280,N_33716);
or U34459 (N_34459,N_33996,N_33291);
and U34460 (N_34460,N_33644,N_33786);
nand U34461 (N_34461,N_33058,N_33154);
nor U34462 (N_34462,N_33354,N_33748);
or U34463 (N_34463,N_33505,N_33546);
nor U34464 (N_34464,N_33195,N_33703);
nor U34465 (N_34465,N_33295,N_33751);
and U34466 (N_34466,N_33536,N_33078);
nand U34467 (N_34467,N_33551,N_33206);
nor U34468 (N_34468,N_33275,N_33226);
nor U34469 (N_34469,N_33453,N_33425);
nor U34470 (N_34470,N_33767,N_33879);
and U34471 (N_34471,N_33353,N_33798);
nand U34472 (N_34472,N_33288,N_33181);
nand U34473 (N_34473,N_33846,N_33839);
and U34474 (N_34474,N_33642,N_33100);
nor U34475 (N_34475,N_33340,N_33562);
nand U34476 (N_34476,N_33571,N_33043);
xnor U34477 (N_34477,N_33190,N_33301);
or U34478 (N_34478,N_33865,N_33034);
and U34479 (N_34479,N_33073,N_33023);
nand U34480 (N_34480,N_33641,N_33851);
xnor U34481 (N_34481,N_33752,N_33007);
nand U34482 (N_34482,N_33094,N_33940);
xor U34483 (N_34483,N_33596,N_33437);
and U34484 (N_34484,N_33526,N_33815);
nand U34485 (N_34485,N_33142,N_33670);
or U34486 (N_34486,N_33721,N_33349);
nand U34487 (N_34487,N_33514,N_33978);
nand U34488 (N_34488,N_33042,N_33850);
and U34489 (N_34489,N_33443,N_33472);
nand U34490 (N_34490,N_33387,N_33402);
or U34491 (N_34491,N_33467,N_33119);
and U34492 (N_34492,N_33608,N_33483);
or U34493 (N_34493,N_33727,N_33290);
and U34494 (N_34494,N_33497,N_33609);
and U34495 (N_34495,N_33104,N_33899);
xnor U34496 (N_34496,N_33780,N_33347);
xor U34497 (N_34497,N_33765,N_33956);
xnor U34498 (N_34498,N_33610,N_33089);
nand U34499 (N_34499,N_33795,N_33969);
or U34500 (N_34500,N_33877,N_33116);
and U34501 (N_34501,N_33114,N_33808);
nand U34502 (N_34502,N_33042,N_33795);
nor U34503 (N_34503,N_33517,N_33534);
nor U34504 (N_34504,N_33957,N_33252);
xor U34505 (N_34505,N_33632,N_33839);
nor U34506 (N_34506,N_33235,N_33965);
nand U34507 (N_34507,N_33321,N_33510);
nand U34508 (N_34508,N_33395,N_33033);
nand U34509 (N_34509,N_33642,N_33036);
and U34510 (N_34510,N_33291,N_33149);
nand U34511 (N_34511,N_33745,N_33690);
nand U34512 (N_34512,N_33328,N_33024);
or U34513 (N_34513,N_33907,N_33062);
nor U34514 (N_34514,N_33836,N_33321);
and U34515 (N_34515,N_33613,N_33872);
or U34516 (N_34516,N_33387,N_33560);
or U34517 (N_34517,N_33048,N_33939);
xor U34518 (N_34518,N_33245,N_33483);
nor U34519 (N_34519,N_33591,N_33781);
or U34520 (N_34520,N_33761,N_33107);
xor U34521 (N_34521,N_33931,N_33265);
xor U34522 (N_34522,N_33726,N_33825);
nand U34523 (N_34523,N_33802,N_33944);
nand U34524 (N_34524,N_33817,N_33693);
xnor U34525 (N_34525,N_33009,N_33224);
nand U34526 (N_34526,N_33552,N_33342);
nor U34527 (N_34527,N_33545,N_33360);
and U34528 (N_34528,N_33256,N_33210);
xor U34529 (N_34529,N_33358,N_33063);
and U34530 (N_34530,N_33072,N_33646);
xnor U34531 (N_34531,N_33658,N_33609);
nand U34532 (N_34532,N_33150,N_33912);
or U34533 (N_34533,N_33735,N_33278);
or U34534 (N_34534,N_33703,N_33779);
and U34535 (N_34535,N_33273,N_33667);
and U34536 (N_34536,N_33582,N_33332);
xnor U34537 (N_34537,N_33391,N_33168);
and U34538 (N_34538,N_33932,N_33412);
nand U34539 (N_34539,N_33014,N_33007);
nor U34540 (N_34540,N_33391,N_33776);
or U34541 (N_34541,N_33980,N_33511);
or U34542 (N_34542,N_33551,N_33789);
and U34543 (N_34543,N_33243,N_33839);
nand U34544 (N_34544,N_33862,N_33273);
nand U34545 (N_34545,N_33595,N_33816);
nand U34546 (N_34546,N_33325,N_33169);
and U34547 (N_34547,N_33647,N_33723);
or U34548 (N_34548,N_33639,N_33597);
or U34549 (N_34549,N_33506,N_33057);
xor U34550 (N_34550,N_33987,N_33228);
xor U34551 (N_34551,N_33547,N_33414);
nor U34552 (N_34552,N_33711,N_33801);
nand U34553 (N_34553,N_33328,N_33437);
and U34554 (N_34554,N_33682,N_33114);
xor U34555 (N_34555,N_33400,N_33897);
and U34556 (N_34556,N_33349,N_33287);
nor U34557 (N_34557,N_33534,N_33696);
xnor U34558 (N_34558,N_33990,N_33361);
and U34559 (N_34559,N_33437,N_33279);
xor U34560 (N_34560,N_33498,N_33464);
or U34561 (N_34561,N_33104,N_33266);
and U34562 (N_34562,N_33960,N_33134);
nand U34563 (N_34563,N_33868,N_33062);
xor U34564 (N_34564,N_33155,N_33407);
xnor U34565 (N_34565,N_33983,N_33142);
nand U34566 (N_34566,N_33475,N_33281);
or U34567 (N_34567,N_33053,N_33661);
xnor U34568 (N_34568,N_33432,N_33677);
and U34569 (N_34569,N_33249,N_33290);
and U34570 (N_34570,N_33613,N_33436);
or U34571 (N_34571,N_33655,N_33929);
nand U34572 (N_34572,N_33215,N_33558);
nor U34573 (N_34573,N_33342,N_33121);
xor U34574 (N_34574,N_33791,N_33677);
nand U34575 (N_34575,N_33501,N_33490);
or U34576 (N_34576,N_33267,N_33504);
nand U34577 (N_34577,N_33078,N_33531);
xor U34578 (N_34578,N_33379,N_33869);
nand U34579 (N_34579,N_33200,N_33268);
nand U34580 (N_34580,N_33515,N_33792);
or U34581 (N_34581,N_33474,N_33918);
and U34582 (N_34582,N_33175,N_33287);
or U34583 (N_34583,N_33505,N_33489);
nand U34584 (N_34584,N_33038,N_33472);
nor U34585 (N_34585,N_33935,N_33806);
and U34586 (N_34586,N_33291,N_33590);
and U34587 (N_34587,N_33885,N_33739);
xor U34588 (N_34588,N_33294,N_33345);
xor U34589 (N_34589,N_33726,N_33183);
xor U34590 (N_34590,N_33005,N_33391);
nand U34591 (N_34591,N_33172,N_33223);
or U34592 (N_34592,N_33679,N_33867);
or U34593 (N_34593,N_33505,N_33102);
or U34594 (N_34594,N_33028,N_33017);
or U34595 (N_34595,N_33235,N_33358);
and U34596 (N_34596,N_33742,N_33558);
and U34597 (N_34597,N_33486,N_33749);
or U34598 (N_34598,N_33444,N_33613);
and U34599 (N_34599,N_33196,N_33312);
and U34600 (N_34600,N_33007,N_33342);
and U34601 (N_34601,N_33674,N_33278);
xnor U34602 (N_34602,N_33373,N_33968);
or U34603 (N_34603,N_33619,N_33494);
xnor U34604 (N_34604,N_33813,N_33698);
or U34605 (N_34605,N_33938,N_33783);
xor U34606 (N_34606,N_33165,N_33853);
xor U34607 (N_34607,N_33987,N_33999);
nand U34608 (N_34608,N_33911,N_33757);
nor U34609 (N_34609,N_33988,N_33915);
nand U34610 (N_34610,N_33602,N_33030);
or U34611 (N_34611,N_33994,N_33010);
xnor U34612 (N_34612,N_33122,N_33861);
nor U34613 (N_34613,N_33673,N_33142);
nor U34614 (N_34614,N_33555,N_33533);
and U34615 (N_34615,N_33789,N_33526);
and U34616 (N_34616,N_33223,N_33214);
and U34617 (N_34617,N_33747,N_33184);
xor U34618 (N_34618,N_33364,N_33671);
or U34619 (N_34619,N_33013,N_33542);
and U34620 (N_34620,N_33771,N_33729);
nor U34621 (N_34621,N_33407,N_33022);
and U34622 (N_34622,N_33109,N_33951);
and U34623 (N_34623,N_33259,N_33907);
and U34624 (N_34624,N_33963,N_33022);
or U34625 (N_34625,N_33840,N_33020);
or U34626 (N_34626,N_33556,N_33827);
nand U34627 (N_34627,N_33637,N_33586);
and U34628 (N_34628,N_33997,N_33995);
or U34629 (N_34629,N_33609,N_33405);
nand U34630 (N_34630,N_33228,N_33180);
and U34631 (N_34631,N_33954,N_33870);
and U34632 (N_34632,N_33988,N_33479);
nor U34633 (N_34633,N_33420,N_33127);
xnor U34634 (N_34634,N_33529,N_33245);
nor U34635 (N_34635,N_33986,N_33398);
nand U34636 (N_34636,N_33381,N_33757);
xnor U34637 (N_34637,N_33615,N_33481);
nor U34638 (N_34638,N_33726,N_33675);
or U34639 (N_34639,N_33669,N_33781);
or U34640 (N_34640,N_33480,N_33784);
nand U34641 (N_34641,N_33854,N_33257);
nor U34642 (N_34642,N_33045,N_33442);
nand U34643 (N_34643,N_33597,N_33031);
xor U34644 (N_34644,N_33450,N_33966);
xor U34645 (N_34645,N_33928,N_33136);
nor U34646 (N_34646,N_33865,N_33269);
and U34647 (N_34647,N_33089,N_33795);
nor U34648 (N_34648,N_33545,N_33211);
nor U34649 (N_34649,N_33325,N_33563);
nand U34650 (N_34650,N_33886,N_33523);
and U34651 (N_34651,N_33680,N_33389);
nand U34652 (N_34652,N_33206,N_33026);
or U34653 (N_34653,N_33992,N_33961);
nand U34654 (N_34654,N_33930,N_33873);
and U34655 (N_34655,N_33045,N_33006);
or U34656 (N_34656,N_33454,N_33803);
and U34657 (N_34657,N_33516,N_33114);
and U34658 (N_34658,N_33121,N_33425);
nor U34659 (N_34659,N_33625,N_33024);
nand U34660 (N_34660,N_33746,N_33285);
or U34661 (N_34661,N_33847,N_33000);
nor U34662 (N_34662,N_33284,N_33422);
or U34663 (N_34663,N_33021,N_33649);
xnor U34664 (N_34664,N_33220,N_33697);
or U34665 (N_34665,N_33726,N_33818);
or U34666 (N_34666,N_33523,N_33081);
nand U34667 (N_34667,N_33502,N_33562);
nor U34668 (N_34668,N_33493,N_33148);
nor U34669 (N_34669,N_33713,N_33584);
or U34670 (N_34670,N_33800,N_33123);
nor U34671 (N_34671,N_33373,N_33795);
or U34672 (N_34672,N_33825,N_33138);
nor U34673 (N_34673,N_33522,N_33138);
nand U34674 (N_34674,N_33555,N_33448);
nor U34675 (N_34675,N_33408,N_33911);
xnor U34676 (N_34676,N_33365,N_33513);
and U34677 (N_34677,N_33272,N_33466);
xor U34678 (N_34678,N_33237,N_33857);
xnor U34679 (N_34679,N_33698,N_33864);
or U34680 (N_34680,N_33230,N_33949);
xnor U34681 (N_34681,N_33799,N_33970);
nor U34682 (N_34682,N_33214,N_33655);
nand U34683 (N_34683,N_33678,N_33407);
nand U34684 (N_34684,N_33103,N_33854);
xnor U34685 (N_34685,N_33301,N_33013);
and U34686 (N_34686,N_33920,N_33230);
or U34687 (N_34687,N_33049,N_33246);
or U34688 (N_34688,N_33820,N_33744);
nor U34689 (N_34689,N_33645,N_33732);
nor U34690 (N_34690,N_33152,N_33916);
xnor U34691 (N_34691,N_33848,N_33152);
nor U34692 (N_34692,N_33561,N_33326);
xnor U34693 (N_34693,N_33556,N_33454);
or U34694 (N_34694,N_33467,N_33630);
xnor U34695 (N_34695,N_33741,N_33949);
nor U34696 (N_34696,N_33469,N_33085);
nand U34697 (N_34697,N_33187,N_33317);
nor U34698 (N_34698,N_33551,N_33010);
xor U34699 (N_34699,N_33023,N_33277);
or U34700 (N_34700,N_33281,N_33649);
nand U34701 (N_34701,N_33721,N_33701);
or U34702 (N_34702,N_33706,N_33663);
nor U34703 (N_34703,N_33421,N_33680);
nand U34704 (N_34704,N_33092,N_33915);
nand U34705 (N_34705,N_33557,N_33765);
nand U34706 (N_34706,N_33691,N_33546);
or U34707 (N_34707,N_33992,N_33478);
nor U34708 (N_34708,N_33742,N_33888);
and U34709 (N_34709,N_33013,N_33757);
nor U34710 (N_34710,N_33278,N_33981);
xnor U34711 (N_34711,N_33831,N_33204);
and U34712 (N_34712,N_33654,N_33688);
nor U34713 (N_34713,N_33602,N_33971);
nand U34714 (N_34714,N_33151,N_33726);
nor U34715 (N_34715,N_33656,N_33919);
nor U34716 (N_34716,N_33489,N_33991);
nand U34717 (N_34717,N_33430,N_33406);
nor U34718 (N_34718,N_33909,N_33432);
or U34719 (N_34719,N_33519,N_33130);
and U34720 (N_34720,N_33607,N_33995);
nor U34721 (N_34721,N_33365,N_33423);
nand U34722 (N_34722,N_33245,N_33777);
nor U34723 (N_34723,N_33761,N_33574);
and U34724 (N_34724,N_33122,N_33660);
or U34725 (N_34725,N_33403,N_33681);
nand U34726 (N_34726,N_33212,N_33716);
or U34727 (N_34727,N_33178,N_33877);
nand U34728 (N_34728,N_33231,N_33466);
xnor U34729 (N_34729,N_33702,N_33499);
xor U34730 (N_34730,N_33570,N_33992);
nor U34731 (N_34731,N_33336,N_33680);
xnor U34732 (N_34732,N_33254,N_33973);
nor U34733 (N_34733,N_33982,N_33692);
and U34734 (N_34734,N_33109,N_33306);
xor U34735 (N_34735,N_33090,N_33147);
or U34736 (N_34736,N_33743,N_33877);
nor U34737 (N_34737,N_33064,N_33828);
xnor U34738 (N_34738,N_33358,N_33665);
nor U34739 (N_34739,N_33945,N_33774);
and U34740 (N_34740,N_33342,N_33879);
xor U34741 (N_34741,N_33659,N_33354);
nand U34742 (N_34742,N_33927,N_33756);
nand U34743 (N_34743,N_33127,N_33035);
or U34744 (N_34744,N_33249,N_33207);
or U34745 (N_34745,N_33066,N_33970);
and U34746 (N_34746,N_33289,N_33672);
and U34747 (N_34747,N_33337,N_33694);
nor U34748 (N_34748,N_33444,N_33031);
nor U34749 (N_34749,N_33580,N_33898);
and U34750 (N_34750,N_33200,N_33189);
xor U34751 (N_34751,N_33367,N_33978);
and U34752 (N_34752,N_33223,N_33806);
xnor U34753 (N_34753,N_33583,N_33041);
xnor U34754 (N_34754,N_33049,N_33851);
xnor U34755 (N_34755,N_33185,N_33081);
xor U34756 (N_34756,N_33261,N_33973);
nand U34757 (N_34757,N_33426,N_33665);
xnor U34758 (N_34758,N_33219,N_33982);
or U34759 (N_34759,N_33603,N_33345);
and U34760 (N_34760,N_33937,N_33228);
nor U34761 (N_34761,N_33827,N_33642);
xnor U34762 (N_34762,N_33607,N_33494);
and U34763 (N_34763,N_33217,N_33274);
xnor U34764 (N_34764,N_33226,N_33461);
nor U34765 (N_34765,N_33352,N_33127);
xnor U34766 (N_34766,N_33984,N_33110);
or U34767 (N_34767,N_33146,N_33369);
nand U34768 (N_34768,N_33178,N_33600);
xnor U34769 (N_34769,N_33399,N_33550);
nor U34770 (N_34770,N_33412,N_33380);
and U34771 (N_34771,N_33020,N_33205);
and U34772 (N_34772,N_33316,N_33745);
nand U34773 (N_34773,N_33150,N_33928);
xor U34774 (N_34774,N_33001,N_33514);
nand U34775 (N_34775,N_33187,N_33337);
and U34776 (N_34776,N_33725,N_33069);
and U34777 (N_34777,N_33285,N_33876);
nor U34778 (N_34778,N_33028,N_33830);
xor U34779 (N_34779,N_33053,N_33788);
or U34780 (N_34780,N_33310,N_33698);
and U34781 (N_34781,N_33385,N_33045);
nor U34782 (N_34782,N_33475,N_33164);
nor U34783 (N_34783,N_33477,N_33298);
and U34784 (N_34784,N_33728,N_33871);
nand U34785 (N_34785,N_33235,N_33799);
xor U34786 (N_34786,N_33927,N_33127);
nand U34787 (N_34787,N_33467,N_33402);
nor U34788 (N_34788,N_33989,N_33192);
and U34789 (N_34789,N_33798,N_33473);
or U34790 (N_34790,N_33551,N_33076);
nor U34791 (N_34791,N_33973,N_33496);
or U34792 (N_34792,N_33182,N_33003);
and U34793 (N_34793,N_33847,N_33219);
xnor U34794 (N_34794,N_33799,N_33105);
xnor U34795 (N_34795,N_33628,N_33414);
nand U34796 (N_34796,N_33145,N_33246);
and U34797 (N_34797,N_33879,N_33654);
and U34798 (N_34798,N_33967,N_33806);
and U34799 (N_34799,N_33285,N_33800);
or U34800 (N_34800,N_33675,N_33751);
and U34801 (N_34801,N_33635,N_33329);
nor U34802 (N_34802,N_33649,N_33763);
xnor U34803 (N_34803,N_33675,N_33216);
nand U34804 (N_34804,N_33638,N_33440);
or U34805 (N_34805,N_33088,N_33211);
nand U34806 (N_34806,N_33589,N_33569);
or U34807 (N_34807,N_33633,N_33860);
xnor U34808 (N_34808,N_33118,N_33615);
or U34809 (N_34809,N_33201,N_33528);
nand U34810 (N_34810,N_33304,N_33728);
and U34811 (N_34811,N_33053,N_33894);
or U34812 (N_34812,N_33852,N_33060);
or U34813 (N_34813,N_33036,N_33985);
nor U34814 (N_34814,N_33576,N_33948);
xor U34815 (N_34815,N_33134,N_33558);
and U34816 (N_34816,N_33447,N_33246);
nor U34817 (N_34817,N_33413,N_33819);
nor U34818 (N_34818,N_33270,N_33815);
nand U34819 (N_34819,N_33506,N_33836);
nor U34820 (N_34820,N_33762,N_33861);
or U34821 (N_34821,N_33404,N_33361);
or U34822 (N_34822,N_33150,N_33328);
and U34823 (N_34823,N_33675,N_33271);
and U34824 (N_34824,N_33189,N_33455);
and U34825 (N_34825,N_33887,N_33550);
nand U34826 (N_34826,N_33359,N_33985);
nor U34827 (N_34827,N_33080,N_33423);
nand U34828 (N_34828,N_33218,N_33460);
nand U34829 (N_34829,N_33843,N_33797);
or U34830 (N_34830,N_33570,N_33796);
nand U34831 (N_34831,N_33287,N_33817);
and U34832 (N_34832,N_33435,N_33916);
nor U34833 (N_34833,N_33855,N_33026);
xnor U34834 (N_34834,N_33400,N_33798);
nand U34835 (N_34835,N_33217,N_33467);
nand U34836 (N_34836,N_33276,N_33840);
or U34837 (N_34837,N_33569,N_33704);
nand U34838 (N_34838,N_33177,N_33455);
nor U34839 (N_34839,N_33713,N_33281);
and U34840 (N_34840,N_33593,N_33689);
xor U34841 (N_34841,N_33589,N_33676);
nor U34842 (N_34842,N_33307,N_33047);
nor U34843 (N_34843,N_33875,N_33200);
nand U34844 (N_34844,N_33356,N_33724);
or U34845 (N_34845,N_33497,N_33335);
nand U34846 (N_34846,N_33023,N_33025);
or U34847 (N_34847,N_33636,N_33480);
xor U34848 (N_34848,N_33693,N_33810);
or U34849 (N_34849,N_33130,N_33943);
xor U34850 (N_34850,N_33358,N_33218);
xor U34851 (N_34851,N_33288,N_33360);
nor U34852 (N_34852,N_33209,N_33253);
nand U34853 (N_34853,N_33472,N_33597);
xnor U34854 (N_34854,N_33431,N_33719);
nand U34855 (N_34855,N_33488,N_33285);
nand U34856 (N_34856,N_33906,N_33283);
nand U34857 (N_34857,N_33666,N_33148);
xor U34858 (N_34858,N_33630,N_33353);
nand U34859 (N_34859,N_33265,N_33448);
or U34860 (N_34860,N_33748,N_33515);
and U34861 (N_34861,N_33934,N_33549);
nand U34862 (N_34862,N_33875,N_33614);
nor U34863 (N_34863,N_33029,N_33266);
or U34864 (N_34864,N_33553,N_33386);
xnor U34865 (N_34865,N_33191,N_33043);
nor U34866 (N_34866,N_33839,N_33967);
nor U34867 (N_34867,N_33423,N_33945);
or U34868 (N_34868,N_33710,N_33964);
nand U34869 (N_34869,N_33039,N_33048);
nand U34870 (N_34870,N_33626,N_33817);
nor U34871 (N_34871,N_33312,N_33835);
and U34872 (N_34872,N_33191,N_33396);
nor U34873 (N_34873,N_33438,N_33667);
or U34874 (N_34874,N_33334,N_33683);
xnor U34875 (N_34875,N_33092,N_33694);
nand U34876 (N_34876,N_33166,N_33135);
and U34877 (N_34877,N_33435,N_33668);
and U34878 (N_34878,N_33210,N_33235);
or U34879 (N_34879,N_33282,N_33830);
nand U34880 (N_34880,N_33796,N_33426);
nand U34881 (N_34881,N_33379,N_33561);
or U34882 (N_34882,N_33887,N_33789);
nor U34883 (N_34883,N_33327,N_33206);
and U34884 (N_34884,N_33311,N_33245);
nand U34885 (N_34885,N_33042,N_33041);
or U34886 (N_34886,N_33893,N_33372);
nand U34887 (N_34887,N_33255,N_33633);
xor U34888 (N_34888,N_33584,N_33980);
nand U34889 (N_34889,N_33010,N_33440);
or U34890 (N_34890,N_33305,N_33718);
and U34891 (N_34891,N_33546,N_33519);
nor U34892 (N_34892,N_33198,N_33780);
xnor U34893 (N_34893,N_33480,N_33833);
nor U34894 (N_34894,N_33210,N_33900);
xor U34895 (N_34895,N_33775,N_33193);
nand U34896 (N_34896,N_33053,N_33142);
or U34897 (N_34897,N_33492,N_33894);
nand U34898 (N_34898,N_33230,N_33141);
xor U34899 (N_34899,N_33005,N_33331);
and U34900 (N_34900,N_33432,N_33022);
and U34901 (N_34901,N_33268,N_33414);
nor U34902 (N_34902,N_33947,N_33333);
nand U34903 (N_34903,N_33918,N_33803);
nor U34904 (N_34904,N_33807,N_33936);
nor U34905 (N_34905,N_33541,N_33550);
or U34906 (N_34906,N_33405,N_33347);
nand U34907 (N_34907,N_33461,N_33295);
xor U34908 (N_34908,N_33062,N_33920);
xnor U34909 (N_34909,N_33432,N_33796);
nor U34910 (N_34910,N_33812,N_33502);
nand U34911 (N_34911,N_33258,N_33242);
xnor U34912 (N_34912,N_33924,N_33199);
or U34913 (N_34913,N_33383,N_33082);
nand U34914 (N_34914,N_33872,N_33465);
or U34915 (N_34915,N_33760,N_33525);
or U34916 (N_34916,N_33112,N_33534);
nand U34917 (N_34917,N_33405,N_33101);
xor U34918 (N_34918,N_33208,N_33289);
nand U34919 (N_34919,N_33354,N_33236);
and U34920 (N_34920,N_33461,N_33783);
and U34921 (N_34921,N_33633,N_33376);
or U34922 (N_34922,N_33839,N_33899);
or U34923 (N_34923,N_33592,N_33916);
nand U34924 (N_34924,N_33626,N_33279);
nor U34925 (N_34925,N_33340,N_33952);
nor U34926 (N_34926,N_33752,N_33083);
nor U34927 (N_34927,N_33902,N_33996);
xor U34928 (N_34928,N_33058,N_33200);
xnor U34929 (N_34929,N_33729,N_33553);
xnor U34930 (N_34930,N_33150,N_33350);
and U34931 (N_34931,N_33699,N_33417);
and U34932 (N_34932,N_33838,N_33095);
or U34933 (N_34933,N_33289,N_33436);
xor U34934 (N_34934,N_33414,N_33240);
nor U34935 (N_34935,N_33586,N_33171);
nand U34936 (N_34936,N_33225,N_33713);
nand U34937 (N_34937,N_33923,N_33418);
xnor U34938 (N_34938,N_33470,N_33194);
and U34939 (N_34939,N_33742,N_33573);
nand U34940 (N_34940,N_33213,N_33443);
and U34941 (N_34941,N_33032,N_33074);
or U34942 (N_34942,N_33567,N_33446);
nor U34943 (N_34943,N_33030,N_33982);
nor U34944 (N_34944,N_33121,N_33895);
nand U34945 (N_34945,N_33863,N_33676);
nor U34946 (N_34946,N_33698,N_33732);
xor U34947 (N_34947,N_33671,N_33640);
and U34948 (N_34948,N_33112,N_33089);
and U34949 (N_34949,N_33421,N_33664);
nand U34950 (N_34950,N_33761,N_33152);
nand U34951 (N_34951,N_33281,N_33612);
or U34952 (N_34952,N_33323,N_33509);
or U34953 (N_34953,N_33597,N_33738);
xor U34954 (N_34954,N_33404,N_33462);
and U34955 (N_34955,N_33871,N_33130);
and U34956 (N_34956,N_33570,N_33029);
nand U34957 (N_34957,N_33565,N_33340);
xnor U34958 (N_34958,N_33921,N_33266);
or U34959 (N_34959,N_33629,N_33065);
or U34960 (N_34960,N_33532,N_33241);
or U34961 (N_34961,N_33018,N_33948);
nand U34962 (N_34962,N_33503,N_33126);
or U34963 (N_34963,N_33965,N_33783);
nor U34964 (N_34964,N_33005,N_33579);
nand U34965 (N_34965,N_33429,N_33698);
nand U34966 (N_34966,N_33540,N_33554);
and U34967 (N_34967,N_33417,N_33464);
or U34968 (N_34968,N_33910,N_33581);
and U34969 (N_34969,N_33576,N_33117);
nor U34970 (N_34970,N_33126,N_33322);
nand U34971 (N_34971,N_33506,N_33347);
or U34972 (N_34972,N_33139,N_33029);
xnor U34973 (N_34973,N_33026,N_33931);
nand U34974 (N_34974,N_33437,N_33142);
nor U34975 (N_34975,N_33478,N_33761);
or U34976 (N_34976,N_33910,N_33338);
and U34977 (N_34977,N_33935,N_33244);
nor U34978 (N_34978,N_33487,N_33127);
or U34979 (N_34979,N_33489,N_33517);
and U34980 (N_34980,N_33467,N_33070);
or U34981 (N_34981,N_33678,N_33857);
and U34982 (N_34982,N_33508,N_33642);
nor U34983 (N_34983,N_33121,N_33549);
and U34984 (N_34984,N_33257,N_33125);
and U34985 (N_34985,N_33745,N_33405);
nor U34986 (N_34986,N_33606,N_33784);
nand U34987 (N_34987,N_33511,N_33710);
and U34988 (N_34988,N_33819,N_33653);
xor U34989 (N_34989,N_33463,N_33835);
or U34990 (N_34990,N_33107,N_33078);
nor U34991 (N_34991,N_33347,N_33996);
xor U34992 (N_34992,N_33764,N_33689);
xnor U34993 (N_34993,N_33561,N_33907);
xor U34994 (N_34994,N_33949,N_33253);
and U34995 (N_34995,N_33921,N_33310);
xor U34996 (N_34996,N_33545,N_33227);
nand U34997 (N_34997,N_33383,N_33857);
nor U34998 (N_34998,N_33648,N_33047);
nor U34999 (N_34999,N_33668,N_33981);
or U35000 (N_35000,N_34921,N_34405);
nor U35001 (N_35001,N_34995,N_34880);
nand U35002 (N_35002,N_34330,N_34485);
xor U35003 (N_35003,N_34558,N_34067);
xnor U35004 (N_35004,N_34990,N_34229);
nand U35005 (N_35005,N_34607,N_34453);
or U35006 (N_35006,N_34134,N_34821);
nand U35007 (N_35007,N_34370,N_34554);
xor U35008 (N_35008,N_34731,N_34970);
and U35009 (N_35009,N_34872,N_34513);
nor U35010 (N_35010,N_34075,N_34559);
or U35011 (N_35011,N_34522,N_34155);
nor U35012 (N_35012,N_34501,N_34357);
or U35013 (N_35013,N_34673,N_34956);
or U35014 (N_35014,N_34749,N_34534);
nor U35015 (N_35015,N_34805,N_34244);
or U35016 (N_35016,N_34191,N_34841);
nand U35017 (N_35017,N_34910,N_34593);
and U35018 (N_35018,N_34350,N_34263);
nand U35019 (N_35019,N_34630,N_34683);
or U35020 (N_35020,N_34437,N_34313);
nor U35021 (N_35021,N_34410,N_34972);
or U35022 (N_35022,N_34891,N_34419);
and U35023 (N_35023,N_34792,N_34707);
xor U35024 (N_35024,N_34069,N_34623);
xor U35025 (N_35025,N_34871,N_34709);
nor U35026 (N_35026,N_34601,N_34220);
or U35027 (N_35027,N_34675,N_34704);
and U35028 (N_35028,N_34374,N_34271);
or U35029 (N_35029,N_34449,N_34609);
nor U35030 (N_35030,N_34729,N_34467);
or U35031 (N_35031,N_34482,N_34552);
xor U35032 (N_35032,N_34119,N_34298);
nand U35033 (N_35033,N_34603,N_34829);
or U35034 (N_35034,N_34176,N_34939);
xor U35035 (N_35035,N_34963,N_34632);
nand U35036 (N_35036,N_34373,N_34865);
xnor U35037 (N_35037,N_34351,N_34051);
or U35038 (N_35038,N_34053,N_34787);
and U35039 (N_35039,N_34786,N_34917);
or U35040 (N_35040,N_34376,N_34145);
nand U35041 (N_35041,N_34780,N_34907);
nor U35042 (N_35042,N_34836,N_34671);
nand U35043 (N_35043,N_34483,N_34008);
nor U35044 (N_35044,N_34743,N_34183);
nor U35045 (N_35045,N_34906,N_34817);
and U35046 (N_35046,N_34532,N_34884);
xnor U35047 (N_35047,N_34269,N_34988);
nand U35048 (N_35048,N_34202,N_34904);
nand U35049 (N_35049,N_34864,N_34457);
nor U35050 (N_35050,N_34063,N_34839);
or U35051 (N_35051,N_34934,N_34153);
nor U35052 (N_35052,N_34040,N_34944);
xor U35053 (N_35053,N_34626,N_34504);
nor U35054 (N_35054,N_34463,N_34827);
nand U35055 (N_35055,N_34898,N_34021);
and U35056 (N_35056,N_34336,N_34814);
nand U35057 (N_35057,N_34149,N_34451);
nor U35058 (N_35058,N_34052,N_34819);
and U35059 (N_35059,N_34016,N_34143);
nor U35060 (N_35060,N_34117,N_34126);
and U35061 (N_35061,N_34505,N_34318);
nand U35062 (N_35062,N_34658,N_34869);
xor U35063 (N_35063,N_34835,N_34033);
xor U35064 (N_35064,N_34035,N_34049);
nor U35065 (N_35065,N_34672,N_34068);
and U35066 (N_35066,N_34642,N_34338);
nor U35067 (N_35067,N_34386,N_34677);
xnor U35068 (N_35068,N_34618,N_34546);
xor U35069 (N_35069,N_34659,N_34822);
xor U35070 (N_35070,N_34364,N_34388);
or U35071 (N_35071,N_34916,N_34863);
nor U35072 (N_35072,N_34039,N_34484);
and U35073 (N_35073,N_34550,N_34566);
nor U35074 (N_35074,N_34693,N_34181);
and U35075 (N_35075,N_34684,N_34197);
or U35076 (N_35076,N_34846,N_34694);
nor U35077 (N_35077,N_34250,N_34077);
or U35078 (N_35078,N_34238,N_34310);
or U35079 (N_35079,N_34895,N_34273);
and U35080 (N_35080,N_34661,N_34211);
xnor U35081 (N_35081,N_34538,N_34432);
and U35082 (N_35082,N_34306,N_34133);
and U35083 (N_35083,N_34643,N_34424);
nor U35084 (N_35084,N_34740,N_34480);
nand U35085 (N_35085,N_34175,N_34032);
and U35086 (N_35086,N_34936,N_34109);
xor U35087 (N_35087,N_34790,N_34201);
and U35088 (N_35088,N_34699,N_34043);
xor U35089 (N_35089,N_34314,N_34442);
xor U35090 (N_35090,N_34520,N_34966);
or U35091 (N_35091,N_34355,N_34565);
or U35092 (N_35092,N_34443,N_34678);
or U35093 (N_35093,N_34938,N_34870);
xnor U35094 (N_35094,N_34209,N_34610);
nor U35095 (N_35095,N_34685,N_34163);
or U35096 (N_35096,N_34222,N_34637);
nor U35097 (N_35097,N_34901,N_34070);
or U35098 (N_35098,N_34369,N_34418);
nand U35099 (N_35099,N_34396,N_34038);
and U35100 (N_35100,N_34084,N_34257);
nand U35101 (N_35101,N_34947,N_34812);
nand U35102 (N_35102,N_34606,N_34025);
or U35103 (N_35103,N_34706,N_34539);
nor U35104 (N_35104,N_34614,N_34845);
or U35105 (N_35105,N_34085,N_34312);
nor U35106 (N_35106,N_34695,N_34274);
and U35107 (N_35107,N_34890,N_34826);
or U35108 (N_35108,N_34104,N_34221);
nor U35109 (N_35109,N_34042,N_34524);
nand U35110 (N_35110,N_34189,N_34590);
xor U35111 (N_35111,N_34304,N_34877);
or U35112 (N_35112,N_34582,N_34150);
nand U35113 (N_35113,N_34624,N_34363);
xnor U35114 (N_35114,N_34154,N_34999);
nand U35115 (N_35115,N_34592,N_34608);
nor U35116 (N_35116,N_34708,N_34783);
or U35117 (N_35117,N_34952,N_34237);
or U35118 (N_35118,N_34848,N_34978);
nor U35119 (N_35119,N_34561,N_34296);
nand U35120 (N_35120,N_34256,N_34406);
xor U35121 (N_35121,N_34896,N_34733);
or U35122 (N_35122,N_34616,N_34118);
xor U35123 (N_35123,N_34245,N_34454);
nand U35124 (N_35124,N_34665,N_34108);
nor U35125 (N_35125,N_34439,N_34862);
nor U35126 (N_35126,N_34859,N_34303);
and U35127 (N_35127,N_34487,N_34844);
or U35128 (N_35128,N_34146,N_34900);
xnor U35129 (N_35129,N_34161,N_34588);
xor U35130 (N_35130,N_34098,N_34837);
and U35131 (N_35131,N_34726,N_34991);
or U35132 (N_35132,N_34090,N_34998);
xor U35133 (N_35133,N_34850,N_34131);
nor U35134 (N_35134,N_34493,N_34761);
xnor U35135 (N_35135,N_34377,N_34171);
or U35136 (N_35136,N_34361,N_34022);
nand U35137 (N_35137,N_34002,N_34205);
nand U35138 (N_35138,N_34739,N_34088);
nor U35139 (N_35139,N_34302,N_34169);
or U35140 (N_35140,N_34969,N_34390);
or U35141 (N_35141,N_34751,N_34430);
nor U35142 (N_35142,N_34691,N_34241);
or U35143 (N_35143,N_34387,N_34286);
or U35144 (N_35144,N_34563,N_34889);
xnor U35145 (N_35145,N_34359,N_34931);
nand U35146 (N_35146,N_34120,N_34213);
nand U35147 (N_35147,N_34472,N_34311);
or U35148 (N_35148,N_34544,N_34059);
xnor U35149 (N_35149,N_34247,N_34315);
and U35150 (N_35150,N_34649,N_34885);
or U35151 (N_35151,N_34955,N_34433);
and U35152 (N_35152,N_34778,N_34329);
or U35153 (N_35153,N_34922,N_34662);
or U35154 (N_35154,N_34072,N_34349);
nor U35155 (N_35155,N_34692,N_34689);
or U35156 (N_35156,N_34818,N_34977);
or U35157 (N_35157,N_34718,N_34356);
and U35158 (N_35158,N_34249,N_34734);
xnor U35159 (N_35159,N_34946,N_34748);
and U35160 (N_35160,N_34100,N_34317);
and U35161 (N_35161,N_34802,N_34490);
xor U35162 (N_35162,N_34326,N_34801);
and U35163 (N_35163,N_34168,N_34669);
or U35164 (N_35164,N_34055,N_34010);
nor U35165 (N_35165,N_34989,N_34855);
nand U35166 (N_35166,N_34144,N_34741);
nand U35167 (N_35167,N_34687,N_34767);
or U35168 (N_35168,N_34288,N_34861);
and U35169 (N_35169,N_34064,N_34525);
xor U35170 (N_35170,N_34402,N_34605);
nand U35171 (N_35171,N_34560,N_34325);
nand U35172 (N_35172,N_34172,N_34395);
and U35173 (N_35173,N_34236,N_34346);
or U35174 (N_35174,N_34058,N_34887);
nand U35175 (N_35175,N_34368,N_34389);
nor U35176 (N_35176,N_34879,N_34591);
or U35177 (N_35177,N_34795,N_34971);
or U35178 (N_35178,N_34347,N_34755);
xnor U35179 (N_35179,N_34994,N_34173);
nand U35180 (N_35180,N_34653,N_34166);
nand U35181 (N_35181,N_34737,N_34182);
and U35182 (N_35182,N_34019,N_34625);
nor U35183 (N_35183,N_34383,N_34526);
xor U35184 (N_35184,N_34148,N_34644);
or U35185 (N_35185,N_34597,N_34730);
nand U35186 (N_35186,N_34132,N_34057);
and U35187 (N_35187,N_34567,N_34461);
or U35188 (N_35188,N_34757,N_34471);
xor U35189 (N_35189,N_34226,N_34178);
or U35190 (N_35190,N_34345,N_34655);
or U35191 (N_35191,N_34506,N_34151);
nor U35192 (N_35192,N_34335,N_34681);
nor U35193 (N_35193,N_34280,N_34445);
xor U35194 (N_35194,N_34727,N_34140);
and U35195 (N_35195,N_34823,N_34092);
nor U35196 (N_35196,N_34029,N_34961);
and U35197 (N_35197,N_34001,N_34628);
xor U35198 (N_35198,N_34409,N_34268);
and U35199 (N_35199,N_34803,N_34005);
and U35200 (N_35200,N_34078,N_34459);
nand U35201 (N_35201,N_34287,N_34414);
nand U35202 (N_35202,N_34279,N_34997);
nand U35203 (N_35203,N_34519,N_34631);
and U35204 (N_35204,N_34056,N_34198);
xnor U35205 (N_35205,N_34788,N_34228);
nand U35206 (N_35206,N_34412,N_34596);
or U35207 (N_35207,N_34000,N_34224);
nand U35208 (N_35208,N_34400,N_34696);
and U35209 (N_35209,N_34572,N_34720);
xnor U35210 (N_35210,N_34436,N_34050);
or U35211 (N_35211,N_34425,N_34621);
or U35212 (N_35212,N_34307,N_34768);
nand U35213 (N_35213,N_34779,N_34750);
or U35214 (N_35214,N_34996,N_34340);
nor U35215 (N_35215,N_34458,N_34545);
nand U35216 (N_35216,N_34796,N_34640);
or U35217 (N_35217,N_34259,N_34045);
or U35218 (N_35218,N_34600,N_34937);
nor U35219 (N_35219,N_34551,N_34509);
xor U35220 (N_35220,N_34018,N_34212);
or U35221 (N_35221,N_34984,N_34832);
or U35222 (N_35222,N_34371,N_34107);
xnor U35223 (N_35223,N_34281,N_34617);
nor U35224 (N_35224,N_34030,N_34867);
or U35225 (N_35225,N_34242,N_34785);
nand U35226 (N_35226,N_34702,N_34004);
or U35227 (N_35227,N_34820,N_34494);
or U35228 (N_35228,N_34073,N_34926);
nor U35229 (N_35229,N_34929,N_34752);
nand U35230 (N_35230,N_34114,N_34930);
or U35231 (N_35231,N_34523,N_34246);
nor U35232 (N_35232,N_34127,N_34394);
and U35233 (N_35233,N_34782,N_34128);
nor U35234 (N_35234,N_34948,N_34012);
nand U35235 (N_35235,N_34079,N_34612);
or U35236 (N_35236,N_34511,N_34456);
xor U35237 (N_35237,N_34137,N_34636);
or U35238 (N_35238,N_34499,N_34091);
nor U35239 (N_35239,N_34489,N_34428);
xnor U35240 (N_35240,N_34736,N_34646);
nand U35241 (N_35241,N_34233,N_34446);
nor U35242 (N_35242,N_34711,N_34024);
nand U35243 (N_35243,N_34275,N_34103);
or U35244 (N_35244,N_34267,N_34099);
or U35245 (N_35245,N_34670,N_34219);
xor U35246 (N_35246,N_34611,N_34903);
nor U35247 (N_35247,N_34775,N_34847);
nand U35248 (N_35248,N_34676,N_34352);
nand U35249 (N_35249,N_34116,N_34076);
nor U35250 (N_35250,N_34299,N_34066);
and U35251 (N_35251,N_34083,N_34744);
nand U35252 (N_35252,N_34682,N_34422);
xnor U35253 (N_35253,N_34578,N_34272);
nor U35254 (N_35254,N_34397,N_34933);
and U35255 (N_35255,N_34697,N_34897);
and U35256 (N_35256,N_34911,N_34048);
and U35257 (N_35257,N_34343,N_34794);
and U35258 (N_35258,N_34065,N_34964);
or U35259 (N_35259,N_34654,N_34633);
or U35260 (N_35260,N_34300,N_34874);
nor U35261 (N_35261,N_34027,N_34124);
nor U35262 (N_35262,N_34285,N_34838);
nor U35263 (N_35263,N_34095,N_34136);
and U35264 (N_35264,N_34913,N_34585);
xnor U35265 (N_35265,N_34765,N_34810);
xnor U35266 (N_35266,N_34575,N_34378);
xnor U35267 (N_35267,N_34725,N_34138);
and U35268 (N_35268,N_34615,N_34622);
or U35269 (N_35269,N_34723,N_34411);
and U35270 (N_35270,N_34759,N_34417);
xnor U35271 (N_35271,N_34094,N_34570);
and U35272 (N_35272,N_34160,N_34382);
nand U35273 (N_35273,N_34721,N_34714);
and U35274 (N_35274,N_34619,N_34258);
xor U35275 (N_35275,N_34892,N_34452);
or U35276 (N_35276,N_34421,N_34753);
xor U35277 (N_35277,N_34594,N_34193);
nor U35278 (N_35278,N_34252,N_34992);
xor U35279 (N_35279,N_34980,N_34983);
xnor U35280 (N_35280,N_34147,N_34123);
xnor U35281 (N_35281,N_34517,N_34294);
nor U35282 (N_35282,N_34974,N_34715);
nand U35283 (N_35283,N_34036,N_34014);
nand U35284 (N_35284,N_34284,N_34062);
nand U35285 (N_35285,N_34139,N_34320);
xor U35286 (N_35286,N_34840,N_34404);
and U35287 (N_35287,N_34899,N_34293);
xnor U35288 (N_35288,N_34037,N_34440);
nor U35289 (N_35289,N_34508,N_34557);
nand U35290 (N_35290,N_34398,N_34297);
nor U35291 (N_35291,N_34235,N_34918);
or U35292 (N_35292,N_34192,N_34112);
nand U35293 (N_35293,N_34074,N_34690);
or U35294 (N_35294,N_34825,N_34031);
nor U35295 (N_35295,N_34738,N_34549);
nor U35296 (N_35296,N_34354,N_34122);
and U35297 (N_35297,N_34384,N_34333);
nand U35298 (N_35298,N_34555,N_34113);
and U35299 (N_35299,N_34415,N_34876);
and U35300 (N_35300,N_34009,N_34516);
nor U35301 (N_35301,N_34510,N_34190);
or U35302 (N_35302,N_34660,N_34215);
nand U35303 (N_35303,N_34322,N_34015);
xor U35304 (N_35304,N_34060,N_34679);
and U35305 (N_35305,N_34089,N_34196);
nand U35306 (N_35306,N_34344,N_34957);
or U35307 (N_35307,N_34833,N_34204);
nor U35308 (N_35308,N_34959,N_34776);
or U35309 (N_35309,N_34573,N_34656);
nand U35310 (N_35310,N_34366,N_34973);
and U35311 (N_35311,N_34081,N_34629);
nor U35312 (N_35312,N_34564,N_34981);
nand U35313 (N_35313,N_34717,N_34745);
and U35314 (N_35314,N_34502,N_34919);
and U35315 (N_35315,N_34486,N_34875);
nand U35316 (N_35316,N_34466,N_34843);
and U35317 (N_35317,N_34162,N_34993);
nor U35318 (N_35318,N_34834,N_34853);
nand U35319 (N_35319,N_34071,N_34831);
xor U35320 (N_35320,N_34760,N_34866);
and U35321 (N_35321,N_34521,N_34928);
and U35322 (N_35322,N_34087,N_34470);
and U35323 (N_35323,N_34231,N_34571);
nand U35324 (N_35324,N_34447,N_34905);
nor U35325 (N_35325,N_34023,N_34185);
or U35326 (N_35326,N_34492,N_34399);
or U35327 (N_35327,N_34982,N_34547);
or U35328 (N_35328,N_34710,N_34791);
nand U35329 (N_35329,N_34082,N_34054);
nand U35330 (N_35330,N_34518,N_34479);
and U35331 (N_35331,N_34945,N_34854);
nor U35332 (N_35332,N_34769,N_34497);
nor U35333 (N_35333,N_34713,N_34806);
nand U35334 (N_35334,N_34968,N_34141);
xnor U35335 (N_35335,N_34650,N_34225);
xnor U35336 (N_35336,N_34540,N_34353);
or U35337 (N_35337,N_34041,N_34503);
nand U35338 (N_35338,N_34979,N_34758);
nand U35339 (N_35339,N_34438,N_34584);
xnor U35340 (N_35340,N_34495,N_34548);
nor U35341 (N_35341,N_34341,N_34883);
xnor U35342 (N_35342,N_34276,N_34308);
and U35343 (N_35343,N_34260,N_34535);
and U35344 (N_35344,N_34652,N_34908);
or U35345 (N_35345,N_34924,N_34180);
nand U35346 (N_35346,N_34253,N_34179);
and U35347 (N_35347,N_34770,N_34809);
and U35348 (N_35348,N_34536,N_34125);
xor U35349 (N_35349,N_34638,N_34849);
xor U35350 (N_35350,N_34476,N_34747);
xor U35351 (N_35351,N_34232,N_34047);
nor U35352 (N_35352,N_34342,N_34932);
or U35353 (N_35353,N_34531,N_34771);
xnor U35354 (N_35354,N_34960,N_34651);
and U35355 (N_35355,N_34407,N_34746);
xor U35356 (N_35356,N_34429,N_34214);
or U35357 (N_35357,N_34102,N_34950);
xnor U35358 (N_35358,N_34381,N_34589);
nand U35359 (N_35359,N_34339,N_34949);
nor U35360 (N_35360,N_34556,N_34164);
and U35361 (N_35361,N_34774,N_34888);
and U35362 (N_35362,N_34987,N_34732);
xnor U35363 (N_35363,N_34360,N_34923);
xnor U35364 (N_35364,N_34915,N_34334);
or U35365 (N_35365,N_34188,N_34159);
nand U35366 (N_35366,N_34784,N_34115);
or U35367 (N_35367,N_34323,N_34886);
or U35368 (N_35368,N_34647,N_34627);
and U35369 (N_35369,N_34097,N_34441);
and U35370 (N_35370,N_34290,N_34431);
nor U35371 (N_35371,N_34044,N_34562);
nand U35372 (N_35372,N_34240,N_34719);
and U35373 (N_35373,N_34265,N_34580);
and U35374 (N_35374,N_34537,N_34261);
xor U35375 (N_35375,N_34423,N_34724);
nand U35376 (N_35376,N_34909,N_34203);
xnor U35377 (N_35377,N_34688,N_34797);
and U35378 (N_35378,N_34365,N_34645);
and U35379 (N_35379,N_34291,N_34427);
or U35380 (N_35380,N_34583,N_34498);
and U35381 (N_35381,N_34210,N_34170);
and U35382 (N_35382,N_34587,N_34216);
nand U35383 (N_35383,N_34003,N_34804);
nand U35384 (N_35384,N_34375,N_34868);
and U35385 (N_35385,N_34800,N_34327);
nand U35386 (N_35386,N_34264,N_34105);
nor U35387 (N_35387,N_34664,N_34129);
xnor U35388 (N_35388,N_34251,N_34852);
or U35389 (N_35389,N_34324,N_34912);
nor U35390 (N_35390,N_34700,N_34954);
or U35391 (N_35391,N_34301,N_34234);
nand U35392 (N_35392,N_34332,N_34475);
and U35393 (N_35393,N_34528,N_34766);
nand U35394 (N_35394,N_34953,N_34860);
nor U35395 (N_35395,N_34507,N_34393);
and U35396 (N_35396,N_34135,N_34667);
nand U35397 (N_35397,N_34789,N_34028);
xor U35398 (N_35398,N_34481,N_34914);
nor U35399 (N_35399,N_34392,N_34529);
xnor U35400 (N_35400,N_34533,N_34469);
nor U35401 (N_35401,N_34080,N_34680);
nand U35402 (N_35402,N_34735,N_34195);
xor U35403 (N_35403,N_34277,N_34061);
nor U35404 (N_35404,N_34106,N_34086);
xnor U35405 (N_35405,N_34174,N_34362);
nand U35406 (N_35406,N_34292,N_34530);
xnor U35407 (N_35407,N_34478,N_34894);
xnor U35408 (N_35408,N_34828,N_34416);
xnor U35409 (N_35409,N_34046,N_34882);
nand U35410 (N_35410,N_34270,N_34965);
xor U35411 (N_35411,N_34305,N_34595);
nand U35412 (N_35412,N_34703,N_34975);
nand U35413 (N_35413,N_34319,N_34756);
and U35414 (N_35414,N_34130,N_34798);
nor U35415 (N_35415,N_34579,N_34674);
nand U35416 (N_35416,N_34426,N_34208);
or U35417 (N_35417,N_34764,N_34401);
and U35418 (N_35418,N_34206,N_34553);
or U35419 (N_35419,N_34613,N_34142);
nor U35420 (N_35420,N_34266,N_34167);
nor U35421 (N_35421,N_34006,N_34278);
and U35422 (N_35422,N_34096,N_34468);
nand U35423 (N_35423,N_34824,N_34477);
and U35424 (N_35424,N_34460,N_34728);
nand U35425 (N_35425,N_34013,N_34420);
nor U35426 (N_35426,N_34121,N_34586);
nand U35427 (N_35427,N_34316,N_34199);
nor U35428 (N_35428,N_34435,N_34663);
and U35429 (N_35429,N_34391,N_34465);
or U35430 (N_35430,N_34379,N_34496);
nor U35431 (N_35431,N_34902,N_34712);
or U35432 (N_35432,N_34927,N_34218);
xor U35433 (N_35433,N_34985,N_34295);
or U35434 (N_35434,N_34413,N_34254);
and U35435 (N_35435,N_34742,N_34576);
xor U35436 (N_35436,N_34668,N_34514);
nor U35437 (N_35437,N_34156,N_34815);
or U35438 (N_35438,N_34289,N_34110);
xnor U35439 (N_35439,N_34858,N_34158);
and U35440 (N_35440,N_34941,N_34604);
nor U35441 (N_35441,N_34958,N_34230);
and U35442 (N_35442,N_34793,N_34473);
xor U35443 (N_35443,N_34657,N_34830);
and U35444 (N_35444,N_34722,N_34194);
and U35445 (N_35445,N_34177,N_34569);
nor U35446 (N_35446,N_34026,N_34328);
nor U35447 (N_35447,N_34434,N_34856);
or U35448 (N_35448,N_34842,N_34186);
nor U35449 (N_35449,N_34873,N_34007);
xor U35450 (N_35450,N_34925,N_34701);
nand U35451 (N_35451,N_34634,N_34034);
or U35452 (N_35452,N_34641,N_34282);
nor U35453 (N_35453,N_34309,N_34541);
xor U35454 (N_35454,N_34635,N_34337);
and U35455 (N_35455,N_34450,N_34200);
nand U35456 (N_35456,N_34799,N_34878);
nor U35457 (N_35457,N_34358,N_34620);
nor U35458 (N_35458,N_34942,N_34372);
and U35459 (N_35459,N_34542,N_34403);
xor U35460 (N_35460,N_34772,N_34262);
or U35461 (N_35461,N_34811,N_34602);
or U35462 (N_35462,N_34808,N_34935);
xnor U35463 (N_35463,N_34283,N_34348);
nor U35464 (N_35464,N_34816,N_34331);
and U35465 (N_35465,N_34639,N_34217);
or U35466 (N_35466,N_34599,N_34951);
nand U35467 (N_35467,N_34754,N_34101);
or U35468 (N_35468,N_34491,N_34207);
nand U35469 (N_35469,N_34515,N_34581);
and U35470 (N_35470,N_34111,N_34763);
and U35471 (N_35471,N_34574,N_34686);
nor U35472 (N_35472,N_34321,N_34385);
xor U35473 (N_35473,N_34474,N_34017);
xnor U35474 (N_35474,N_34187,N_34512);
or U35475 (N_35475,N_34962,N_34444);
xnor U35476 (N_35476,N_34857,N_34976);
xor U35477 (N_35477,N_34152,N_34940);
or U35478 (N_35478,N_34255,N_34227);
or U35479 (N_35479,N_34380,N_34464);
nor U35480 (N_35480,N_34967,N_34157);
or U35481 (N_35481,N_34705,N_34543);
and U35482 (N_35482,N_34568,N_34462);
or U35483 (N_35483,N_34093,N_34527);
nand U35484 (N_35484,N_34851,N_34020);
nor U35485 (N_35485,N_34920,N_34243);
and U35486 (N_35486,N_34408,N_34777);
and U35487 (N_35487,N_34666,N_34500);
nor U35488 (N_35488,N_34223,N_34698);
xor U35489 (N_35489,N_34239,N_34184);
xnor U35490 (N_35490,N_34488,N_34893);
xnor U35491 (N_35491,N_34943,N_34248);
and U35492 (N_35492,N_34807,N_34455);
and U35493 (N_35493,N_34762,N_34367);
nand U35494 (N_35494,N_34881,N_34448);
nand U35495 (N_35495,N_34165,N_34781);
and U35496 (N_35496,N_34598,N_34648);
xnor U35497 (N_35497,N_34773,N_34986);
or U35498 (N_35498,N_34716,N_34813);
and U35499 (N_35499,N_34577,N_34011);
nand U35500 (N_35500,N_34011,N_34000);
and U35501 (N_35501,N_34711,N_34795);
nand U35502 (N_35502,N_34771,N_34951);
and U35503 (N_35503,N_34361,N_34235);
xor U35504 (N_35504,N_34113,N_34607);
and U35505 (N_35505,N_34509,N_34908);
nand U35506 (N_35506,N_34143,N_34658);
or U35507 (N_35507,N_34000,N_34609);
or U35508 (N_35508,N_34119,N_34294);
nor U35509 (N_35509,N_34182,N_34670);
or U35510 (N_35510,N_34657,N_34648);
or U35511 (N_35511,N_34055,N_34948);
or U35512 (N_35512,N_34692,N_34289);
and U35513 (N_35513,N_34444,N_34350);
and U35514 (N_35514,N_34299,N_34883);
nand U35515 (N_35515,N_34169,N_34495);
nand U35516 (N_35516,N_34379,N_34372);
and U35517 (N_35517,N_34219,N_34904);
or U35518 (N_35518,N_34836,N_34277);
xor U35519 (N_35519,N_34767,N_34404);
or U35520 (N_35520,N_34361,N_34482);
or U35521 (N_35521,N_34829,N_34914);
nand U35522 (N_35522,N_34667,N_34724);
or U35523 (N_35523,N_34076,N_34428);
xor U35524 (N_35524,N_34960,N_34887);
and U35525 (N_35525,N_34111,N_34261);
nand U35526 (N_35526,N_34383,N_34399);
and U35527 (N_35527,N_34940,N_34617);
xnor U35528 (N_35528,N_34745,N_34386);
or U35529 (N_35529,N_34912,N_34146);
and U35530 (N_35530,N_34179,N_34709);
and U35531 (N_35531,N_34927,N_34144);
or U35532 (N_35532,N_34849,N_34892);
nand U35533 (N_35533,N_34824,N_34132);
nor U35534 (N_35534,N_34465,N_34894);
or U35535 (N_35535,N_34110,N_34525);
nand U35536 (N_35536,N_34801,N_34775);
xor U35537 (N_35537,N_34679,N_34213);
or U35538 (N_35538,N_34199,N_34852);
nand U35539 (N_35539,N_34059,N_34616);
and U35540 (N_35540,N_34778,N_34594);
and U35541 (N_35541,N_34906,N_34719);
nand U35542 (N_35542,N_34278,N_34835);
nor U35543 (N_35543,N_34221,N_34720);
xor U35544 (N_35544,N_34408,N_34710);
nor U35545 (N_35545,N_34573,N_34011);
xnor U35546 (N_35546,N_34395,N_34053);
nor U35547 (N_35547,N_34659,N_34044);
or U35548 (N_35548,N_34071,N_34492);
and U35549 (N_35549,N_34289,N_34284);
or U35550 (N_35550,N_34479,N_34033);
and U35551 (N_35551,N_34148,N_34960);
xnor U35552 (N_35552,N_34116,N_34703);
nor U35553 (N_35553,N_34276,N_34312);
nor U35554 (N_35554,N_34990,N_34276);
xor U35555 (N_35555,N_34757,N_34021);
nand U35556 (N_35556,N_34823,N_34369);
or U35557 (N_35557,N_34218,N_34308);
xnor U35558 (N_35558,N_34950,N_34454);
xnor U35559 (N_35559,N_34881,N_34019);
xor U35560 (N_35560,N_34839,N_34149);
and U35561 (N_35561,N_34173,N_34049);
xor U35562 (N_35562,N_34493,N_34487);
xnor U35563 (N_35563,N_34650,N_34477);
nand U35564 (N_35564,N_34961,N_34687);
xnor U35565 (N_35565,N_34926,N_34257);
nand U35566 (N_35566,N_34891,N_34311);
or U35567 (N_35567,N_34661,N_34985);
xor U35568 (N_35568,N_34499,N_34362);
nand U35569 (N_35569,N_34667,N_34283);
nor U35570 (N_35570,N_34285,N_34877);
and U35571 (N_35571,N_34544,N_34423);
or U35572 (N_35572,N_34233,N_34881);
xnor U35573 (N_35573,N_34297,N_34069);
xor U35574 (N_35574,N_34777,N_34839);
xor U35575 (N_35575,N_34013,N_34997);
nand U35576 (N_35576,N_34585,N_34398);
and U35577 (N_35577,N_34959,N_34884);
nand U35578 (N_35578,N_34764,N_34046);
nor U35579 (N_35579,N_34166,N_34503);
or U35580 (N_35580,N_34746,N_34956);
and U35581 (N_35581,N_34524,N_34064);
xnor U35582 (N_35582,N_34992,N_34189);
and U35583 (N_35583,N_34023,N_34479);
or U35584 (N_35584,N_34707,N_34521);
and U35585 (N_35585,N_34866,N_34614);
or U35586 (N_35586,N_34446,N_34067);
nand U35587 (N_35587,N_34034,N_34651);
nand U35588 (N_35588,N_34116,N_34503);
nor U35589 (N_35589,N_34321,N_34665);
xnor U35590 (N_35590,N_34576,N_34628);
nand U35591 (N_35591,N_34270,N_34211);
xor U35592 (N_35592,N_34474,N_34762);
nand U35593 (N_35593,N_34794,N_34045);
xor U35594 (N_35594,N_34724,N_34149);
and U35595 (N_35595,N_34399,N_34528);
or U35596 (N_35596,N_34748,N_34386);
nand U35597 (N_35597,N_34451,N_34713);
nor U35598 (N_35598,N_34784,N_34043);
nand U35599 (N_35599,N_34042,N_34780);
nand U35600 (N_35600,N_34161,N_34006);
xnor U35601 (N_35601,N_34794,N_34002);
nand U35602 (N_35602,N_34877,N_34555);
or U35603 (N_35603,N_34651,N_34326);
xnor U35604 (N_35604,N_34093,N_34761);
xnor U35605 (N_35605,N_34843,N_34012);
xor U35606 (N_35606,N_34507,N_34597);
xor U35607 (N_35607,N_34066,N_34756);
and U35608 (N_35608,N_34606,N_34852);
or U35609 (N_35609,N_34228,N_34186);
xor U35610 (N_35610,N_34362,N_34896);
xnor U35611 (N_35611,N_34621,N_34994);
nand U35612 (N_35612,N_34876,N_34345);
nor U35613 (N_35613,N_34490,N_34247);
or U35614 (N_35614,N_34539,N_34627);
or U35615 (N_35615,N_34816,N_34404);
nor U35616 (N_35616,N_34918,N_34939);
nand U35617 (N_35617,N_34104,N_34082);
or U35618 (N_35618,N_34853,N_34262);
and U35619 (N_35619,N_34177,N_34500);
nand U35620 (N_35620,N_34007,N_34366);
and U35621 (N_35621,N_34426,N_34682);
or U35622 (N_35622,N_34808,N_34413);
nand U35623 (N_35623,N_34555,N_34207);
xor U35624 (N_35624,N_34141,N_34455);
nor U35625 (N_35625,N_34987,N_34027);
and U35626 (N_35626,N_34983,N_34550);
and U35627 (N_35627,N_34684,N_34185);
nor U35628 (N_35628,N_34793,N_34426);
and U35629 (N_35629,N_34768,N_34537);
or U35630 (N_35630,N_34223,N_34218);
or U35631 (N_35631,N_34202,N_34664);
xnor U35632 (N_35632,N_34035,N_34044);
and U35633 (N_35633,N_34943,N_34741);
or U35634 (N_35634,N_34734,N_34341);
nand U35635 (N_35635,N_34460,N_34994);
nor U35636 (N_35636,N_34871,N_34275);
nor U35637 (N_35637,N_34907,N_34831);
nand U35638 (N_35638,N_34245,N_34310);
nand U35639 (N_35639,N_34887,N_34996);
nor U35640 (N_35640,N_34318,N_34379);
and U35641 (N_35641,N_34332,N_34254);
or U35642 (N_35642,N_34573,N_34138);
or U35643 (N_35643,N_34534,N_34898);
nor U35644 (N_35644,N_34710,N_34809);
and U35645 (N_35645,N_34253,N_34915);
nor U35646 (N_35646,N_34965,N_34984);
xnor U35647 (N_35647,N_34582,N_34176);
nor U35648 (N_35648,N_34857,N_34537);
nand U35649 (N_35649,N_34982,N_34526);
nand U35650 (N_35650,N_34168,N_34235);
nor U35651 (N_35651,N_34381,N_34739);
nand U35652 (N_35652,N_34064,N_34864);
and U35653 (N_35653,N_34469,N_34266);
or U35654 (N_35654,N_34011,N_34841);
and U35655 (N_35655,N_34903,N_34933);
nor U35656 (N_35656,N_34039,N_34422);
nand U35657 (N_35657,N_34688,N_34199);
or U35658 (N_35658,N_34421,N_34902);
and U35659 (N_35659,N_34213,N_34336);
xor U35660 (N_35660,N_34382,N_34935);
nand U35661 (N_35661,N_34052,N_34047);
nand U35662 (N_35662,N_34364,N_34684);
and U35663 (N_35663,N_34420,N_34583);
nor U35664 (N_35664,N_34265,N_34963);
and U35665 (N_35665,N_34938,N_34233);
and U35666 (N_35666,N_34968,N_34338);
and U35667 (N_35667,N_34465,N_34811);
xnor U35668 (N_35668,N_34697,N_34477);
xor U35669 (N_35669,N_34553,N_34674);
and U35670 (N_35670,N_34599,N_34152);
and U35671 (N_35671,N_34505,N_34155);
nor U35672 (N_35672,N_34009,N_34552);
xor U35673 (N_35673,N_34929,N_34134);
nand U35674 (N_35674,N_34261,N_34234);
nand U35675 (N_35675,N_34622,N_34638);
nand U35676 (N_35676,N_34845,N_34045);
and U35677 (N_35677,N_34028,N_34794);
nor U35678 (N_35678,N_34875,N_34842);
nand U35679 (N_35679,N_34291,N_34827);
nand U35680 (N_35680,N_34085,N_34869);
xnor U35681 (N_35681,N_34122,N_34370);
and U35682 (N_35682,N_34050,N_34233);
nor U35683 (N_35683,N_34202,N_34248);
or U35684 (N_35684,N_34248,N_34868);
nand U35685 (N_35685,N_34474,N_34348);
xor U35686 (N_35686,N_34295,N_34787);
nand U35687 (N_35687,N_34446,N_34095);
nor U35688 (N_35688,N_34999,N_34458);
nand U35689 (N_35689,N_34901,N_34483);
xnor U35690 (N_35690,N_34996,N_34796);
and U35691 (N_35691,N_34859,N_34438);
xor U35692 (N_35692,N_34879,N_34201);
nor U35693 (N_35693,N_34487,N_34107);
xnor U35694 (N_35694,N_34959,N_34231);
xnor U35695 (N_35695,N_34417,N_34050);
and U35696 (N_35696,N_34851,N_34447);
nand U35697 (N_35697,N_34605,N_34058);
nor U35698 (N_35698,N_34655,N_34711);
nand U35699 (N_35699,N_34431,N_34464);
xor U35700 (N_35700,N_34655,N_34904);
and U35701 (N_35701,N_34588,N_34753);
and U35702 (N_35702,N_34501,N_34240);
xnor U35703 (N_35703,N_34669,N_34166);
or U35704 (N_35704,N_34112,N_34062);
nor U35705 (N_35705,N_34074,N_34202);
nor U35706 (N_35706,N_34403,N_34237);
xor U35707 (N_35707,N_34900,N_34744);
and U35708 (N_35708,N_34620,N_34424);
or U35709 (N_35709,N_34510,N_34973);
or U35710 (N_35710,N_34697,N_34854);
and U35711 (N_35711,N_34897,N_34797);
or U35712 (N_35712,N_34674,N_34431);
and U35713 (N_35713,N_34697,N_34667);
xor U35714 (N_35714,N_34090,N_34965);
nand U35715 (N_35715,N_34206,N_34933);
and U35716 (N_35716,N_34168,N_34475);
or U35717 (N_35717,N_34275,N_34984);
xnor U35718 (N_35718,N_34554,N_34572);
nand U35719 (N_35719,N_34763,N_34002);
and U35720 (N_35720,N_34319,N_34170);
and U35721 (N_35721,N_34899,N_34177);
and U35722 (N_35722,N_34712,N_34000);
or U35723 (N_35723,N_34368,N_34700);
and U35724 (N_35724,N_34498,N_34647);
xor U35725 (N_35725,N_34525,N_34384);
nor U35726 (N_35726,N_34186,N_34901);
and U35727 (N_35727,N_34373,N_34097);
or U35728 (N_35728,N_34614,N_34137);
or U35729 (N_35729,N_34327,N_34622);
or U35730 (N_35730,N_34039,N_34660);
nand U35731 (N_35731,N_34492,N_34356);
and U35732 (N_35732,N_34062,N_34317);
nand U35733 (N_35733,N_34330,N_34949);
nand U35734 (N_35734,N_34485,N_34309);
and U35735 (N_35735,N_34858,N_34620);
nand U35736 (N_35736,N_34980,N_34816);
and U35737 (N_35737,N_34272,N_34796);
nor U35738 (N_35738,N_34401,N_34377);
nand U35739 (N_35739,N_34483,N_34135);
or U35740 (N_35740,N_34903,N_34014);
or U35741 (N_35741,N_34531,N_34845);
or U35742 (N_35742,N_34559,N_34816);
or U35743 (N_35743,N_34705,N_34779);
or U35744 (N_35744,N_34104,N_34165);
xor U35745 (N_35745,N_34257,N_34336);
nor U35746 (N_35746,N_34046,N_34512);
or U35747 (N_35747,N_34727,N_34803);
and U35748 (N_35748,N_34107,N_34297);
nor U35749 (N_35749,N_34078,N_34574);
or U35750 (N_35750,N_34026,N_34251);
and U35751 (N_35751,N_34159,N_34420);
nand U35752 (N_35752,N_34638,N_34468);
nor U35753 (N_35753,N_34308,N_34972);
nor U35754 (N_35754,N_34584,N_34848);
nor U35755 (N_35755,N_34315,N_34451);
and U35756 (N_35756,N_34315,N_34554);
or U35757 (N_35757,N_34860,N_34032);
nand U35758 (N_35758,N_34483,N_34568);
xnor U35759 (N_35759,N_34388,N_34550);
nor U35760 (N_35760,N_34947,N_34559);
nand U35761 (N_35761,N_34066,N_34143);
xnor U35762 (N_35762,N_34684,N_34878);
and U35763 (N_35763,N_34011,N_34243);
nor U35764 (N_35764,N_34979,N_34636);
nor U35765 (N_35765,N_34364,N_34090);
or U35766 (N_35766,N_34322,N_34688);
xnor U35767 (N_35767,N_34677,N_34409);
nand U35768 (N_35768,N_34210,N_34146);
or U35769 (N_35769,N_34659,N_34569);
nand U35770 (N_35770,N_34431,N_34377);
or U35771 (N_35771,N_34343,N_34220);
nor U35772 (N_35772,N_34923,N_34306);
xor U35773 (N_35773,N_34251,N_34772);
or U35774 (N_35774,N_34427,N_34539);
and U35775 (N_35775,N_34066,N_34282);
xor U35776 (N_35776,N_34358,N_34424);
or U35777 (N_35777,N_34522,N_34639);
or U35778 (N_35778,N_34238,N_34811);
and U35779 (N_35779,N_34969,N_34498);
or U35780 (N_35780,N_34696,N_34543);
or U35781 (N_35781,N_34105,N_34240);
nor U35782 (N_35782,N_34570,N_34952);
or U35783 (N_35783,N_34842,N_34654);
nor U35784 (N_35784,N_34620,N_34041);
nor U35785 (N_35785,N_34345,N_34374);
nand U35786 (N_35786,N_34198,N_34206);
xnor U35787 (N_35787,N_34279,N_34489);
or U35788 (N_35788,N_34307,N_34989);
nor U35789 (N_35789,N_34332,N_34012);
nor U35790 (N_35790,N_34217,N_34625);
nor U35791 (N_35791,N_34866,N_34523);
or U35792 (N_35792,N_34154,N_34553);
or U35793 (N_35793,N_34082,N_34577);
or U35794 (N_35794,N_34638,N_34528);
and U35795 (N_35795,N_34695,N_34410);
xor U35796 (N_35796,N_34938,N_34030);
or U35797 (N_35797,N_34389,N_34189);
nand U35798 (N_35798,N_34732,N_34064);
xor U35799 (N_35799,N_34316,N_34975);
and U35800 (N_35800,N_34041,N_34978);
or U35801 (N_35801,N_34190,N_34585);
nor U35802 (N_35802,N_34094,N_34400);
or U35803 (N_35803,N_34833,N_34121);
nand U35804 (N_35804,N_34145,N_34372);
nand U35805 (N_35805,N_34446,N_34778);
nand U35806 (N_35806,N_34283,N_34104);
or U35807 (N_35807,N_34371,N_34313);
nand U35808 (N_35808,N_34989,N_34513);
and U35809 (N_35809,N_34592,N_34841);
or U35810 (N_35810,N_34723,N_34819);
nand U35811 (N_35811,N_34444,N_34887);
xnor U35812 (N_35812,N_34638,N_34788);
nand U35813 (N_35813,N_34010,N_34151);
xor U35814 (N_35814,N_34741,N_34009);
nor U35815 (N_35815,N_34722,N_34421);
nor U35816 (N_35816,N_34516,N_34423);
nand U35817 (N_35817,N_34275,N_34155);
nor U35818 (N_35818,N_34072,N_34558);
nand U35819 (N_35819,N_34982,N_34306);
and U35820 (N_35820,N_34960,N_34033);
xor U35821 (N_35821,N_34222,N_34710);
xnor U35822 (N_35822,N_34880,N_34500);
and U35823 (N_35823,N_34758,N_34956);
or U35824 (N_35824,N_34990,N_34447);
nand U35825 (N_35825,N_34892,N_34507);
and U35826 (N_35826,N_34585,N_34807);
nor U35827 (N_35827,N_34014,N_34470);
nand U35828 (N_35828,N_34623,N_34935);
nand U35829 (N_35829,N_34325,N_34688);
xnor U35830 (N_35830,N_34957,N_34529);
or U35831 (N_35831,N_34771,N_34092);
nor U35832 (N_35832,N_34168,N_34156);
nand U35833 (N_35833,N_34392,N_34561);
and U35834 (N_35834,N_34416,N_34841);
xnor U35835 (N_35835,N_34302,N_34653);
nor U35836 (N_35836,N_34343,N_34213);
nand U35837 (N_35837,N_34694,N_34934);
xor U35838 (N_35838,N_34709,N_34512);
xor U35839 (N_35839,N_34404,N_34268);
nand U35840 (N_35840,N_34301,N_34862);
nor U35841 (N_35841,N_34125,N_34122);
and U35842 (N_35842,N_34531,N_34930);
xnor U35843 (N_35843,N_34001,N_34160);
xor U35844 (N_35844,N_34208,N_34028);
xor U35845 (N_35845,N_34419,N_34225);
xnor U35846 (N_35846,N_34954,N_34067);
nand U35847 (N_35847,N_34418,N_34822);
or U35848 (N_35848,N_34232,N_34803);
xnor U35849 (N_35849,N_34073,N_34940);
nand U35850 (N_35850,N_34812,N_34899);
nor U35851 (N_35851,N_34779,N_34211);
xnor U35852 (N_35852,N_34978,N_34632);
and U35853 (N_35853,N_34656,N_34856);
and U35854 (N_35854,N_34636,N_34403);
nor U35855 (N_35855,N_34941,N_34675);
and U35856 (N_35856,N_34881,N_34828);
xnor U35857 (N_35857,N_34163,N_34975);
or U35858 (N_35858,N_34718,N_34620);
and U35859 (N_35859,N_34594,N_34954);
xor U35860 (N_35860,N_34094,N_34050);
nand U35861 (N_35861,N_34613,N_34794);
nor U35862 (N_35862,N_34031,N_34458);
and U35863 (N_35863,N_34373,N_34061);
nand U35864 (N_35864,N_34862,N_34034);
xnor U35865 (N_35865,N_34175,N_34413);
nand U35866 (N_35866,N_34214,N_34159);
nor U35867 (N_35867,N_34591,N_34018);
and U35868 (N_35868,N_34835,N_34653);
or U35869 (N_35869,N_34917,N_34234);
xor U35870 (N_35870,N_34055,N_34932);
nand U35871 (N_35871,N_34160,N_34690);
and U35872 (N_35872,N_34161,N_34816);
and U35873 (N_35873,N_34484,N_34951);
nand U35874 (N_35874,N_34070,N_34622);
nand U35875 (N_35875,N_34986,N_34044);
and U35876 (N_35876,N_34193,N_34085);
and U35877 (N_35877,N_34300,N_34409);
nor U35878 (N_35878,N_34299,N_34008);
xor U35879 (N_35879,N_34748,N_34383);
xor U35880 (N_35880,N_34299,N_34939);
xnor U35881 (N_35881,N_34670,N_34940);
nor U35882 (N_35882,N_34162,N_34142);
and U35883 (N_35883,N_34324,N_34246);
xor U35884 (N_35884,N_34528,N_34442);
nand U35885 (N_35885,N_34982,N_34009);
or U35886 (N_35886,N_34091,N_34154);
nor U35887 (N_35887,N_34343,N_34255);
or U35888 (N_35888,N_34185,N_34493);
and U35889 (N_35889,N_34578,N_34912);
nor U35890 (N_35890,N_34849,N_34609);
nand U35891 (N_35891,N_34620,N_34220);
xor U35892 (N_35892,N_34452,N_34730);
or U35893 (N_35893,N_34031,N_34102);
xor U35894 (N_35894,N_34546,N_34219);
nor U35895 (N_35895,N_34300,N_34754);
and U35896 (N_35896,N_34196,N_34740);
nor U35897 (N_35897,N_34048,N_34906);
nand U35898 (N_35898,N_34319,N_34556);
xnor U35899 (N_35899,N_34101,N_34425);
nor U35900 (N_35900,N_34249,N_34607);
nand U35901 (N_35901,N_34787,N_34964);
nand U35902 (N_35902,N_34272,N_34725);
or U35903 (N_35903,N_34774,N_34443);
and U35904 (N_35904,N_34208,N_34438);
or U35905 (N_35905,N_34496,N_34739);
nor U35906 (N_35906,N_34038,N_34436);
and U35907 (N_35907,N_34797,N_34961);
and U35908 (N_35908,N_34093,N_34427);
and U35909 (N_35909,N_34331,N_34080);
nand U35910 (N_35910,N_34145,N_34964);
nand U35911 (N_35911,N_34351,N_34906);
nor U35912 (N_35912,N_34152,N_34099);
nand U35913 (N_35913,N_34888,N_34295);
and U35914 (N_35914,N_34880,N_34065);
xor U35915 (N_35915,N_34606,N_34727);
or U35916 (N_35916,N_34016,N_34918);
or U35917 (N_35917,N_34699,N_34027);
nand U35918 (N_35918,N_34459,N_34407);
and U35919 (N_35919,N_34597,N_34397);
and U35920 (N_35920,N_34310,N_34398);
and U35921 (N_35921,N_34065,N_34815);
and U35922 (N_35922,N_34874,N_34157);
nand U35923 (N_35923,N_34275,N_34681);
xor U35924 (N_35924,N_34726,N_34008);
nand U35925 (N_35925,N_34446,N_34014);
nand U35926 (N_35926,N_34647,N_34138);
and U35927 (N_35927,N_34793,N_34217);
nand U35928 (N_35928,N_34233,N_34930);
nand U35929 (N_35929,N_34836,N_34878);
nor U35930 (N_35930,N_34203,N_34530);
xnor U35931 (N_35931,N_34478,N_34719);
nor U35932 (N_35932,N_34205,N_34569);
xnor U35933 (N_35933,N_34326,N_34170);
nor U35934 (N_35934,N_34155,N_34818);
nand U35935 (N_35935,N_34505,N_34102);
or U35936 (N_35936,N_34485,N_34529);
and U35937 (N_35937,N_34360,N_34633);
xnor U35938 (N_35938,N_34595,N_34972);
nand U35939 (N_35939,N_34695,N_34042);
xor U35940 (N_35940,N_34832,N_34479);
nand U35941 (N_35941,N_34804,N_34085);
and U35942 (N_35942,N_34329,N_34737);
or U35943 (N_35943,N_34931,N_34695);
nor U35944 (N_35944,N_34761,N_34221);
nand U35945 (N_35945,N_34702,N_34764);
nor U35946 (N_35946,N_34881,N_34501);
xor U35947 (N_35947,N_34575,N_34443);
and U35948 (N_35948,N_34497,N_34220);
nand U35949 (N_35949,N_34510,N_34935);
nand U35950 (N_35950,N_34004,N_34075);
nand U35951 (N_35951,N_34611,N_34194);
nand U35952 (N_35952,N_34470,N_34773);
nor U35953 (N_35953,N_34849,N_34832);
or U35954 (N_35954,N_34663,N_34913);
and U35955 (N_35955,N_34695,N_34515);
xor U35956 (N_35956,N_34916,N_34560);
and U35957 (N_35957,N_34200,N_34140);
nand U35958 (N_35958,N_34244,N_34861);
xnor U35959 (N_35959,N_34984,N_34312);
or U35960 (N_35960,N_34472,N_34463);
nand U35961 (N_35961,N_34553,N_34215);
or U35962 (N_35962,N_34940,N_34270);
or U35963 (N_35963,N_34711,N_34147);
nor U35964 (N_35964,N_34744,N_34277);
and U35965 (N_35965,N_34234,N_34757);
nand U35966 (N_35966,N_34755,N_34423);
nor U35967 (N_35967,N_34697,N_34880);
xor U35968 (N_35968,N_34089,N_34242);
xnor U35969 (N_35969,N_34935,N_34733);
nand U35970 (N_35970,N_34538,N_34923);
nand U35971 (N_35971,N_34614,N_34287);
and U35972 (N_35972,N_34100,N_34603);
nand U35973 (N_35973,N_34620,N_34178);
nand U35974 (N_35974,N_34511,N_34758);
or U35975 (N_35975,N_34737,N_34219);
nand U35976 (N_35976,N_34580,N_34888);
and U35977 (N_35977,N_34021,N_34157);
and U35978 (N_35978,N_34409,N_34744);
or U35979 (N_35979,N_34856,N_34677);
xor U35980 (N_35980,N_34198,N_34683);
nand U35981 (N_35981,N_34781,N_34075);
and U35982 (N_35982,N_34536,N_34318);
and U35983 (N_35983,N_34042,N_34265);
nand U35984 (N_35984,N_34526,N_34890);
or U35985 (N_35985,N_34154,N_34600);
xor U35986 (N_35986,N_34684,N_34398);
nor U35987 (N_35987,N_34505,N_34671);
nand U35988 (N_35988,N_34928,N_34382);
nor U35989 (N_35989,N_34470,N_34338);
xor U35990 (N_35990,N_34758,N_34645);
and U35991 (N_35991,N_34030,N_34620);
nand U35992 (N_35992,N_34648,N_34411);
xor U35993 (N_35993,N_34126,N_34574);
or U35994 (N_35994,N_34850,N_34430);
xor U35995 (N_35995,N_34881,N_34270);
xnor U35996 (N_35996,N_34734,N_34013);
xor U35997 (N_35997,N_34694,N_34920);
and U35998 (N_35998,N_34273,N_34721);
or U35999 (N_35999,N_34593,N_34213);
nand U36000 (N_36000,N_35696,N_35355);
nand U36001 (N_36001,N_35318,N_35503);
nor U36002 (N_36002,N_35501,N_35829);
and U36003 (N_36003,N_35329,N_35723);
nor U36004 (N_36004,N_35281,N_35908);
and U36005 (N_36005,N_35132,N_35474);
and U36006 (N_36006,N_35458,N_35207);
nor U36007 (N_36007,N_35983,N_35114);
nand U36008 (N_36008,N_35016,N_35764);
nor U36009 (N_36009,N_35015,N_35813);
and U36010 (N_36010,N_35367,N_35586);
nand U36011 (N_36011,N_35164,N_35344);
xor U36012 (N_36012,N_35333,N_35285);
nand U36013 (N_36013,N_35427,N_35748);
or U36014 (N_36014,N_35537,N_35794);
nor U36015 (N_36015,N_35403,N_35663);
or U36016 (N_36016,N_35293,N_35969);
nor U36017 (N_36017,N_35664,N_35235);
or U36018 (N_36018,N_35528,N_35411);
xnor U36019 (N_36019,N_35430,N_35718);
nor U36020 (N_36020,N_35328,N_35496);
nand U36021 (N_36021,N_35311,N_35962);
xnor U36022 (N_36022,N_35163,N_35985);
and U36023 (N_36023,N_35593,N_35107);
and U36024 (N_36024,N_35340,N_35565);
and U36025 (N_36025,N_35850,N_35279);
or U36026 (N_36026,N_35881,N_35704);
nand U36027 (N_36027,N_35889,N_35765);
xor U36028 (N_36028,N_35870,N_35459);
or U36029 (N_36029,N_35486,N_35776);
nor U36030 (N_36030,N_35788,N_35898);
or U36031 (N_36031,N_35313,N_35090);
xnor U36032 (N_36032,N_35131,N_35084);
nand U36033 (N_36033,N_35577,N_35861);
and U36034 (N_36034,N_35797,N_35187);
nand U36035 (N_36035,N_35575,N_35173);
and U36036 (N_36036,N_35552,N_35215);
xnor U36037 (N_36037,N_35771,N_35386);
xor U36038 (N_36038,N_35493,N_35737);
and U36039 (N_36039,N_35315,N_35607);
xor U36040 (N_36040,N_35997,N_35860);
nor U36041 (N_36041,N_35683,N_35820);
and U36042 (N_36042,N_35888,N_35843);
or U36043 (N_36043,N_35609,N_35021);
and U36044 (N_36044,N_35373,N_35990);
nand U36045 (N_36045,N_35183,N_35716);
and U36046 (N_36046,N_35991,N_35128);
xnor U36047 (N_36047,N_35753,N_35446);
xor U36048 (N_36048,N_35227,N_35561);
nand U36049 (N_36049,N_35289,N_35648);
and U36050 (N_36050,N_35694,N_35316);
and U36051 (N_36051,N_35017,N_35801);
nand U36052 (N_36052,N_35996,N_35229);
nor U36053 (N_36053,N_35886,N_35249);
nand U36054 (N_36054,N_35910,N_35245);
or U36055 (N_36055,N_35721,N_35049);
and U36056 (N_36056,N_35484,N_35087);
or U36057 (N_36057,N_35169,N_35959);
nor U36058 (N_36058,N_35652,N_35709);
and U36059 (N_36059,N_35202,N_35225);
or U36060 (N_36060,N_35504,N_35407);
nand U36061 (N_36061,N_35780,N_35011);
nor U36062 (N_36062,N_35795,N_35179);
and U36063 (N_36063,N_35511,N_35489);
or U36064 (N_36064,N_35634,N_35302);
and U36065 (N_36065,N_35751,N_35897);
and U36066 (N_36066,N_35196,N_35295);
nand U36067 (N_36067,N_35693,N_35519);
nor U36068 (N_36068,N_35884,N_35433);
xnor U36069 (N_36069,N_35826,N_35914);
xor U36070 (N_36070,N_35548,N_35998);
nand U36071 (N_36071,N_35608,N_35953);
and U36072 (N_36072,N_35863,N_35812);
and U36073 (N_36073,N_35426,N_35480);
and U36074 (N_36074,N_35122,N_35724);
nand U36075 (N_36075,N_35450,N_35174);
and U36076 (N_36076,N_35182,N_35442);
nor U36077 (N_36077,N_35256,N_35934);
and U36078 (N_36078,N_35680,N_35729);
and U36079 (N_36079,N_35060,N_35097);
nor U36080 (N_36080,N_35554,N_35611);
nor U36081 (N_36081,N_35534,N_35530);
or U36082 (N_36082,N_35138,N_35014);
nor U36083 (N_36083,N_35009,N_35117);
xnor U36084 (N_36084,N_35346,N_35973);
nor U36085 (N_36085,N_35500,N_35210);
nand U36086 (N_36086,N_35181,N_35744);
and U36087 (N_36087,N_35698,N_35774);
nor U36088 (N_36088,N_35789,N_35306);
xor U36089 (N_36089,N_35516,N_35292);
nand U36090 (N_36090,N_35628,N_35214);
nand U36091 (N_36091,N_35241,N_35613);
nor U36092 (N_36092,N_35713,N_35896);
nor U36093 (N_36093,N_35779,N_35986);
or U36094 (N_36094,N_35601,N_35802);
and U36095 (N_36095,N_35301,N_35799);
and U36096 (N_36096,N_35380,N_35655);
and U36097 (N_36097,N_35363,N_35247);
or U36098 (N_36098,N_35465,N_35250);
nor U36099 (N_36099,N_35871,N_35102);
and U36100 (N_36100,N_35069,N_35599);
or U36101 (N_36101,N_35029,N_35665);
nand U36102 (N_36102,N_35522,N_35982);
or U36103 (N_36103,N_35948,N_35711);
nand U36104 (N_36104,N_35167,N_35445);
xnor U36105 (N_36105,N_35630,N_35785);
or U36106 (N_36106,N_35391,N_35644);
xor U36107 (N_36107,N_35510,N_35993);
nor U36108 (N_36108,N_35273,N_35255);
or U36109 (N_36109,N_35464,N_35587);
or U36110 (N_36110,N_35862,N_35398);
xor U36111 (N_36111,N_35457,N_35712);
xor U36112 (N_36112,N_35777,N_35217);
and U36113 (N_36113,N_35961,N_35835);
nand U36114 (N_36114,N_35922,N_35947);
xor U36115 (N_36115,N_35974,N_35451);
nor U36116 (N_36116,N_35823,N_35880);
nor U36117 (N_36117,N_35824,N_35950);
xnor U36118 (N_36118,N_35640,N_35846);
or U36119 (N_36119,N_35538,N_35852);
nand U36120 (N_36120,N_35116,N_35001);
or U36121 (N_36121,N_35702,N_35524);
and U36122 (N_36122,N_35645,N_35578);
nand U36123 (N_36123,N_35019,N_35024);
and U36124 (N_36124,N_35347,N_35335);
xor U36125 (N_36125,N_35471,N_35497);
and U36126 (N_36126,N_35343,N_35514);
or U36127 (N_36127,N_35394,N_35473);
and U36128 (N_36128,N_35485,N_35405);
nor U36129 (N_36129,N_35410,N_35671);
nand U36130 (N_36130,N_35752,N_35858);
nand U36131 (N_36131,N_35298,N_35264);
nand U36132 (N_36132,N_35282,N_35643);
and U36133 (N_36133,N_35818,N_35689);
nor U36134 (N_36134,N_35192,N_35606);
nand U36135 (N_36135,N_35821,N_35906);
and U36136 (N_36136,N_35261,N_35568);
and U36137 (N_36137,N_35072,N_35113);
nor U36138 (N_36138,N_35422,N_35787);
nand U36139 (N_36139,N_35589,N_35415);
or U36140 (N_36140,N_35409,N_35104);
xor U36141 (N_36141,N_35866,N_35618);
xnor U36142 (N_36142,N_35622,N_35044);
xnor U36143 (N_36143,N_35936,N_35436);
xnor U36144 (N_36144,N_35275,N_35656);
and U36145 (N_36145,N_35957,N_35749);
nand U36146 (N_36146,N_35266,N_35231);
nor U36147 (N_36147,N_35833,N_35495);
and U36148 (N_36148,N_35847,N_35195);
nor U36149 (N_36149,N_35203,N_35526);
or U36150 (N_36150,N_35269,N_35762);
nand U36151 (N_36151,N_35073,N_35757);
nand U36152 (N_36152,N_35909,N_35345);
nor U36153 (N_36153,N_35375,N_35383);
nand U36154 (N_36154,N_35389,N_35460);
nand U36155 (N_36155,N_35262,N_35219);
xor U36156 (N_36156,N_35374,N_35356);
or U36157 (N_36157,N_35124,N_35056);
or U36158 (N_36158,N_35837,N_35531);
and U36159 (N_36159,N_35189,N_35088);
or U36160 (N_36160,N_35070,N_35722);
xor U36161 (N_36161,N_35440,N_35542);
nand U36162 (N_36162,N_35617,N_35031);
nor U36163 (N_36163,N_35304,N_35756);
nand U36164 (N_36164,N_35941,N_35105);
nand U36165 (N_36165,N_35632,N_35929);
or U36166 (N_36166,N_35276,N_35498);
nand U36167 (N_36167,N_35958,N_35491);
and U36168 (N_36168,N_35964,N_35421);
or U36169 (N_36169,N_35616,N_35137);
or U36170 (N_36170,N_35218,N_35074);
xnor U36171 (N_36171,N_35152,N_35400);
or U36172 (N_36172,N_35067,N_35574);
xor U36173 (N_36173,N_35651,N_35690);
nor U36174 (N_36174,N_35717,N_35604);
or U36175 (N_36175,N_35584,N_35239);
nor U36176 (N_36176,N_35760,N_35792);
and U36177 (N_36177,N_35778,N_35654);
and U36178 (N_36178,N_35591,N_35359);
or U36179 (N_36179,N_35900,N_35629);
xnor U36180 (N_36180,N_35224,N_35399);
or U36181 (N_36181,N_35803,N_35106);
nor U36182 (N_36182,N_35018,N_35994);
nor U36183 (N_36183,N_35253,N_35170);
nand U36184 (N_36184,N_35223,N_35815);
and U36185 (N_36185,N_35481,N_35585);
or U36186 (N_36186,N_35463,N_35793);
xor U36187 (N_36187,N_35461,N_35423);
or U36188 (N_36188,N_35034,N_35559);
nor U36189 (N_36189,N_35502,N_35057);
or U36190 (N_36190,N_35631,N_35902);
nand U36191 (N_36191,N_35872,N_35290);
xor U36192 (N_36192,N_35819,N_35598);
nand U36193 (N_36193,N_35715,N_35194);
or U36194 (N_36194,N_35669,N_35746);
nor U36195 (N_36195,N_35428,N_35636);
nor U36196 (N_36196,N_35323,N_35236);
xor U36197 (N_36197,N_35545,N_35319);
xnor U36198 (N_36198,N_35177,N_35977);
and U36199 (N_36199,N_35257,N_35842);
and U36200 (N_36200,N_35523,N_35267);
or U36201 (N_36201,N_35555,N_35877);
and U36202 (N_36202,N_35462,N_35414);
nand U36203 (N_36203,N_35377,N_35707);
or U36204 (N_36204,N_35602,N_35342);
nor U36205 (N_36205,N_35350,N_35047);
and U36206 (N_36206,N_35658,N_35995);
or U36207 (N_36207,N_35317,N_35036);
nand U36208 (N_36208,N_35068,N_35556);
nand U36209 (N_36209,N_35867,N_35638);
or U36210 (N_36210,N_35730,N_35701);
xor U36211 (N_36211,N_35784,N_35954);
xor U36212 (N_36212,N_35408,N_35988);
xnor U36213 (N_36213,N_35123,N_35197);
or U36214 (N_36214,N_35558,N_35238);
nor U36215 (N_36215,N_35190,N_35360);
or U36216 (N_36216,N_35331,N_35392);
nand U36217 (N_36217,N_35120,N_35817);
or U36218 (N_36218,N_35930,N_35684);
xnor U36219 (N_36219,N_35620,N_35938);
or U36220 (N_36220,N_35868,N_35506);
nand U36221 (N_36221,N_35726,N_35755);
or U36222 (N_36222,N_35551,N_35564);
xor U36223 (N_36223,N_35062,N_35332);
and U36224 (N_36224,N_35145,N_35844);
and U36225 (N_36225,N_35469,N_35401);
nor U36226 (N_36226,N_35198,N_35066);
xor U36227 (N_36227,N_35322,N_35963);
or U36228 (N_36228,N_35920,N_35614);
nor U36229 (N_36229,N_35854,N_35259);
or U36230 (N_36230,N_35143,N_35810);
xnor U36231 (N_36231,N_35149,N_35184);
xnor U36232 (N_36232,N_35252,N_35926);
or U36233 (N_36233,N_35907,N_35085);
or U36234 (N_36234,N_35121,N_35937);
nand U36235 (N_36235,N_35970,N_35200);
nor U36236 (N_36236,N_35494,N_35595);
nor U36237 (N_36237,N_35045,N_35082);
and U36238 (N_36238,N_35178,N_35507);
nand U36239 (N_36239,N_35895,N_35439);
xnor U36240 (N_36240,N_35093,N_35492);
and U36241 (N_36241,N_35175,N_35912);
and U36242 (N_36242,N_35839,N_35384);
or U36243 (N_36243,N_35321,N_35659);
and U36244 (N_36244,N_35488,N_35096);
nor U36245 (N_36245,N_35625,N_35244);
and U36246 (N_36246,N_35134,N_35213);
nand U36247 (N_36247,N_35869,N_35008);
and U36248 (N_36248,N_35058,N_35467);
xor U36249 (N_36249,N_35532,N_35918);
or U36250 (N_36250,N_35547,N_35432);
or U36251 (N_36251,N_35129,N_35791);
or U36252 (N_36252,N_35845,N_35940);
xor U36253 (N_36253,N_35822,N_35666);
or U36254 (N_36254,N_35188,N_35418);
xor U36255 (N_36255,N_35441,N_35650);
or U36256 (N_36256,N_35657,N_35125);
or U36257 (N_36257,N_35233,N_35515);
and U36258 (N_36258,N_35118,N_35841);
or U36259 (N_36259,N_35443,N_35254);
nor U36260 (N_36260,N_35621,N_35543);
xor U36261 (N_36261,N_35291,N_35126);
nor U36262 (N_36262,N_35274,N_35027);
and U36263 (N_36263,N_35849,N_35059);
and U36264 (N_36264,N_35892,N_35588);
and U36265 (N_36265,N_35052,N_35747);
or U36266 (N_36266,N_35228,N_35061);
and U36267 (N_36267,N_35280,N_35827);
and U36268 (N_36268,N_35299,N_35560);
nor U36269 (N_36269,N_35536,N_35449);
xnor U36270 (N_36270,N_35296,N_35221);
or U36271 (N_36271,N_35590,N_35674);
nor U36272 (N_36272,N_35733,N_35284);
xor U36273 (N_36273,N_35686,N_35240);
nor U36274 (N_36274,N_35055,N_35743);
and U36275 (N_36275,N_35859,N_35978);
nor U36276 (N_36276,N_35155,N_35679);
xnor U36277 (N_36277,N_35147,N_35452);
nor U36278 (N_36278,N_35942,N_35438);
nor U36279 (N_36279,N_35050,N_35487);
nand U36280 (N_36280,N_35670,N_35688);
nor U36281 (N_36281,N_35212,N_35153);
or U36282 (N_36282,N_35731,N_35369);
or U36283 (N_36283,N_35447,N_35740);
or U36284 (N_36284,N_35376,N_35268);
nor U36285 (N_36285,N_35078,N_35208);
and U36286 (N_36286,N_35148,N_35136);
nor U36287 (N_36287,N_35358,N_35265);
xor U36288 (N_36288,N_35853,N_35040);
nor U36289 (N_36289,N_35133,N_35703);
nor U36290 (N_36290,N_35115,N_35165);
and U36291 (N_36291,N_35992,N_35579);
and U36292 (N_36292,N_35150,N_35278);
nor U36293 (N_36293,N_35417,N_35303);
nand U36294 (N_36294,N_35945,N_35808);
or U36295 (N_36295,N_35162,N_35570);
or U36296 (N_36296,N_35790,N_35873);
xor U36297 (N_36297,N_35234,N_35848);
or U36298 (N_36298,N_35573,N_35626);
or U36299 (N_36299,N_35310,N_35309);
xor U36300 (N_36300,N_35566,N_35135);
xnor U36301 (N_36301,N_35226,N_35395);
and U36302 (N_36302,N_35834,N_35569);
or U36303 (N_36303,N_35028,N_35048);
xor U36304 (N_36304,N_35033,N_35939);
nor U36305 (N_36305,N_35357,N_35529);
xnor U36306 (N_36306,N_35007,N_35004);
nor U36307 (N_36307,N_35110,N_35572);
nand U36308 (N_36308,N_35080,N_35071);
nand U36309 (N_36309,N_35075,N_35286);
nor U36310 (N_36310,N_35378,N_35952);
nor U36311 (N_36311,N_35742,N_35020);
or U36312 (N_36312,N_35037,N_35161);
xor U36313 (N_36313,N_35781,N_35989);
xnor U36314 (N_36314,N_35600,N_35928);
and U36315 (N_36315,N_35307,N_35141);
nor U36316 (N_36316,N_35220,N_35766);
or U36317 (N_36317,N_35385,N_35581);
or U36318 (N_36318,N_35258,N_35130);
xnor U36319 (N_36319,N_35975,N_35038);
xnor U36320 (N_36320,N_35270,N_35923);
nand U36321 (N_36321,N_35468,N_35856);
nor U36322 (N_36322,N_35878,N_35882);
or U36323 (N_36323,N_35919,N_35230);
nand U36324 (N_36324,N_35372,N_35435);
and U36325 (N_36325,N_35246,N_35100);
and U36326 (N_36326,N_35580,N_35466);
nand U36327 (N_36327,N_35687,N_35624);
or U36328 (N_36328,N_35754,N_35348);
nand U36329 (N_36329,N_35379,N_35429);
nand U36330 (N_36330,N_35444,N_35805);
nor U36331 (N_36331,N_35035,N_35685);
nand U36332 (N_36332,N_35763,N_35193);
nand U36333 (N_36333,N_35855,N_35662);
and U36334 (N_36334,N_35661,N_35112);
and U36335 (N_36335,N_35916,N_35211);
and U36336 (N_36336,N_35697,N_35352);
xor U36337 (N_36337,N_35158,N_35098);
nor U36338 (N_36338,N_35927,N_35157);
and U36339 (N_36339,N_35944,N_35732);
nand U36340 (N_36340,N_35984,N_35140);
xnor U36341 (N_36341,N_35678,N_35010);
xnor U36342 (N_36342,N_35054,N_35750);
or U36343 (N_36343,N_35980,N_35330);
xor U36344 (N_36344,N_35741,N_35089);
or U36345 (N_36345,N_35368,N_35816);
nand U36346 (N_36346,N_35022,N_35739);
xnor U36347 (N_36347,N_35456,N_35677);
nand U36348 (N_36348,N_35773,N_35758);
nor U36349 (N_36349,N_35828,N_35204);
and U36350 (N_36350,N_35396,N_35705);
xor U36351 (N_36351,N_35243,N_35943);
or U36352 (N_36352,N_35111,N_35904);
and U36353 (N_36353,N_35119,N_35840);
and U36354 (N_36354,N_35594,N_35478);
xor U36355 (N_36355,N_35382,N_35637);
xor U36356 (N_36356,N_35633,N_35647);
xor U36357 (N_36357,N_35349,N_35404);
and U36358 (N_36358,N_35046,N_35475);
and U36359 (N_36359,N_35546,N_35911);
nand U36360 (N_36360,N_35351,N_35798);
xor U36361 (N_36361,N_35025,N_35370);
or U36362 (N_36362,N_35476,N_35783);
nor U36363 (N_36363,N_35354,N_35005);
nor U36364 (N_36364,N_35935,N_35030);
nor U36365 (N_36365,N_35921,N_35099);
or U36366 (N_36366,N_35431,N_35412);
and U36367 (N_36367,N_35003,N_35761);
xnor U36368 (N_36368,N_35232,N_35272);
nand U36369 (N_36369,N_35216,N_35171);
or U36370 (N_36370,N_35660,N_35972);
or U36371 (N_36371,N_35672,N_35520);
and U36372 (N_36372,N_35681,N_35767);
nand U36373 (N_36373,N_35371,N_35108);
or U36374 (N_36374,N_35308,N_35894);
and U36375 (N_36375,N_35700,N_35393);
or U36376 (N_36376,N_35668,N_35879);
or U36377 (N_36377,N_35336,N_35472);
or U36378 (N_36378,N_35676,N_35032);
nor U36379 (N_36379,N_35453,N_35364);
nor U36380 (N_36380,N_35339,N_35425);
xnor U36381 (N_36381,N_35933,N_35361);
or U36382 (N_36382,N_35571,N_35806);
or U36383 (N_36383,N_35260,N_35237);
nor U36384 (N_36384,N_35146,N_35518);
or U36385 (N_36385,N_35151,N_35682);
nor U36386 (N_36386,N_35277,N_35782);
nand U36387 (N_36387,N_35720,N_35925);
or U36388 (N_36388,N_35312,N_35814);
and U36389 (N_36389,N_35470,N_35127);
and U36390 (N_36390,N_35406,N_35201);
nand U36391 (N_36391,N_35159,N_35831);
nand U36392 (N_36392,N_35390,N_35583);
nor U36393 (N_36393,N_35081,N_35337);
and U36394 (N_36394,N_35166,N_35951);
and U36395 (N_36395,N_35796,N_35772);
xor U36396 (N_36396,N_35455,N_35041);
and U36397 (N_36397,N_35101,N_35109);
nand U36398 (N_36398,N_35582,N_35710);
or U36399 (N_36399,N_35728,N_35800);
xor U36400 (N_36400,N_35508,N_35283);
nor U36401 (N_36401,N_35699,N_35890);
xnor U36402 (N_36402,N_35499,N_35051);
or U36403 (N_36403,N_35490,N_35857);
and U36404 (N_36404,N_35366,N_35077);
or U36405 (N_36405,N_35320,N_35987);
xnor U36406 (N_36406,N_35932,N_35966);
or U36407 (N_36407,N_35000,N_35026);
or U36408 (N_36408,N_35769,N_35971);
or U36409 (N_36409,N_35263,N_35525);
and U36410 (N_36410,N_35735,N_35002);
nand U36411 (N_36411,N_35915,N_35300);
nand U36412 (N_36412,N_35513,N_35725);
nand U36413 (N_36413,N_35338,N_35965);
xor U36414 (N_36414,N_35901,N_35649);
nor U36415 (N_36415,N_35541,N_35825);
nor U36416 (N_36416,N_35738,N_35905);
and U36417 (N_36417,N_35615,N_35079);
and U36418 (N_36418,N_35365,N_35064);
and U36419 (N_36419,N_35039,N_35251);
nand U36420 (N_36420,N_35832,N_35448);
xnor U36421 (N_36421,N_35642,N_35838);
nor U36422 (N_36422,N_35186,N_35612);
nand U36423 (N_36423,N_35675,N_35521);
or U36424 (N_36424,N_35592,N_35402);
and U36425 (N_36425,N_35734,N_35271);
or U36426 (N_36426,N_35042,N_35563);
nor U36427 (N_36427,N_35596,N_35065);
xnor U36428 (N_36428,N_35185,N_35597);
and U36429 (N_36429,N_35619,N_35567);
or U36430 (N_36430,N_35786,N_35479);
nor U36431 (N_36431,N_35692,N_35836);
and U36432 (N_36432,N_35539,N_35885);
xor U36433 (N_36433,N_35326,N_35544);
nor U36434 (N_36434,N_35086,N_35206);
nand U36435 (N_36435,N_35397,N_35416);
nor U36436 (N_36436,N_35549,N_35981);
or U36437 (N_36437,N_35509,N_35811);
nand U36438 (N_36438,N_35770,N_35413);
xnor U36439 (N_36439,N_35759,N_35768);
nor U36440 (N_36440,N_35635,N_35388);
or U36441 (N_36441,N_35875,N_35013);
nor U36442 (N_36442,N_35899,N_35830);
and U36443 (N_36443,N_35362,N_35420);
nor U36444 (N_36444,N_35695,N_35540);
nor U36445 (N_36445,N_35887,N_35477);
xor U36446 (N_36446,N_35864,N_35437);
nand U36447 (N_36447,N_35653,N_35727);
nand U36448 (N_36448,N_35483,N_35550);
nand U36449 (N_36449,N_35248,N_35381);
xor U36450 (N_36450,N_35706,N_35083);
or U36451 (N_36451,N_35979,N_35903);
nand U36452 (N_36452,N_35527,N_35095);
nand U36453 (N_36453,N_35891,N_35673);
xnor U36454 (N_36454,N_35324,N_35931);
and U36455 (N_36455,N_35314,N_35053);
and U36456 (N_36456,N_35142,N_35168);
nand U36457 (N_36457,N_35512,N_35623);
nand U36458 (N_36458,N_35865,N_35063);
nand U36459 (N_36459,N_35809,N_35139);
xor U36460 (N_36460,N_35976,N_35288);
nor U36461 (N_36461,N_35199,N_35023);
or U36462 (N_36462,N_35736,N_35876);
and U36463 (N_36463,N_35144,N_35641);
and U36464 (N_36464,N_35043,N_35160);
or U36465 (N_36465,N_35387,N_35960);
nand U36466 (N_36466,N_35419,N_35610);
and U36467 (N_36467,N_35434,N_35924);
nor U36468 (N_36468,N_35667,N_35719);
or U36469 (N_36469,N_35745,N_35505);
nor U36470 (N_36470,N_35454,N_35557);
and U36471 (N_36471,N_35176,N_35334);
nand U36472 (N_36472,N_35603,N_35297);
xor U36473 (N_36473,N_35012,N_35424);
and U36474 (N_36474,N_35807,N_35341);
or U36475 (N_36475,N_35287,N_35242);
xnor U36476 (N_36476,N_35103,N_35094);
xor U36477 (N_36477,N_35956,N_35156);
and U36478 (N_36478,N_35691,N_35006);
or U36479 (N_36479,N_35172,N_35327);
nor U36480 (N_36480,N_35605,N_35946);
xor U36481 (N_36481,N_35576,N_35209);
or U36482 (N_36482,N_35076,N_35955);
nand U36483 (N_36483,N_35714,N_35325);
xor U36484 (N_36484,N_35968,N_35646);
nor U36485 (N_36485,N_35205,N_35917);
and U36486 (N_36486,N_35874,N_35883);
nor U36487 (N_36487,N_35533,N_35949);
xnor U36488 (N_36488,N_35775,N_35708);
or U36489 (N_36489,N_35562,N_35535);
and U36490 (N_36490,N_35180,N_35999);
xnor U36491 (N_36491,N_35517,N_35092);
or U36492 (N_36492,N_35851,N_35305);
nand U36493 (N_36493,N_35294,N_35191);
nand U36494 (N_36494,N_35639,N_35804);
nand U36495 (N_36495,N_35553,N_35893);
xor U36496 (N_36496,N_35627,N_35913);
nand U36497 (N_36497,N_35154,N_35353);
and U36498 (N_36498,N_35482,N_35091);
and U36499 (N_36499,N_35222,N_35967);
xnor U36500 (N_36500,N_35131,N_35342);
and U36501 (N_36501,N_35445,N_35965);
and U36502 (N_36502,N_35286,N_35858);
nor U36503 (N_36503,N_35718,N_35048);
and U36504 (N_36504,N_35352,N_35624);
nand U36505 (N_36505,N_35367,N_35670);
or U36506 (N_36506,N_35973,N_35945);
and U36507 (N_36507,N_35276,N_35426);
or U36508 (N_36508,N_35722,N_35236);
nor U36509 (N_36509,N_35558,N_35027);
nand U36510 (N_36510,N_35564,N_35725);
or U36511 (N_36511,N_35350,N_35836);
nor U36512 (N_36512,N_35699,N_35050);
and U36513 (N_36513,N_35690,N_35283);
or U36514 (N_36514,N_35854,N_35635);
or U36515 (N_36515,N_35336,N_35438);
xnor U36516 (N_36516,N_35099,N_35611);
nor U36517 (N_36517,N_35633,N_35386);
or U36518 (N_36518,N_35900,N_35225);
nand U36519 (N_36519,N_35859,N_35659);
xor U36520 (N_36520,N_35280,N_35931);
nand U36521 (N_36521,N_35528,N_35495);
and U36522 (N_36522,N_35263,N_35782);
nand U36523 (N_36523,N_35032,N_35511);
nor U36524 (N_36524,N_35533,N_35997);
or U36525 (N_36525,N_35555,N_35022);
nor U36526 (N_36526,N_35332,N_35366);
nand U36527 (N_36527,N_35460,N_35213);
nand U36528 (N_36528,N_35451,N_35624);
nand U36529 (N_36529,N_35061,N_35905);
nor U36530 (N_36530,N_35300,N_35885);
nor U36531 (N_36531,N_35673,N_35360);
nor U36532 (N_36532,N_35243,N_35818);
nand U36533 (N_36533,N_35394,N_35229);
and U36534 (N_36534,N_35504,N_35736);
and U36535 (N_36535,N_35756,N_35133);
xnor U36536 (N_36536,N_35721,N_35911);
xor U36537 (N_36537,N_35391,N_35577);
nand U36538 (N_36538,N_35277,N_35096);
and U36539 (N_36539,N_35096,N_35968);
or U36540 (N_36540,N_35187,N_35486);
xor U36541 (N_36541,N_35949,N_35342);
xor U36542 (N_36542,N_35706,N_35983);
or U36543 (N_36543,N_35973,N_35465);
nand U36544 (N_36544,N_35593,N_35077);
nand U36545 (N_36545,N_35665,N_35577);
nand U36546 (N_36546,N_35931,N_35651);
or U36547 (N_36547,N_35723,N_35982);
nor U36548 (N_36548,N_35101,N_35370);
nor U36549 (N_36549,N_35310,N_35690);
nand U36550 (N_36550,N_35175,N_35661);
xnor U36551 (N_36551,N_35508,N_35607);
nand U36552 (N_36552,N_35819,N_35926);
or U36553 (N_36553,N_35436,N_35443);
and U36554 (N_36554,N_35496,N_35227);
xor U36555 (N_36555,N_35268,N_35662);
nand U36556 (N_36556,N_35754,N_35003);
nor U36557 (N_36557,N_35198,N_35641);
nand U36558 (N_36558,N_35383,N_35334);
nand U36559 (N_36559,N_35335,N_35199);
and U36560 (N_36560,N_35874,N_35811);
nor U36561 (N_36561,N_35935,N_35123);
or U36562 (N_36562,N_35686,N_35745);
and U36563 (N_36563,N_35899,N_35528);
xnor U36564 (N_36564,N_35086,N_35796);
xnor U36565 (N_36565,N_35913,N_35620);
nand U36566 (N_36566,N_35908,N_35042);
or U36567 (N_36567,N_35436,N_35578);
or U36568 (N_36568,N_35790,N_35889);
or U36569 (N_36569,N_35213,N_35120);
xor U36570 (N_36570,N_35249,N_35172);
xor U36571 (N_36571,N_35883,N_35109);
nor U36572 (N_36572,N_35171,N_35300);
or U36573 (N_36573,N_35313,N_35305);
nor U36574 (N_36574,N_35240,N_35345);
nand U36575 (N_36575,N_35125,N_35405);
xor U36576 (N_36576,N_35076,N_35375);
or U36577 (N_36577,N_35212,N_35778);
or U36578 (N_36578,N_35515,N_35170);
nand U36579 (N_36579,N_35203,N_35581);
or U36580 (N_36580,N_35399,N_35330);
nor U36581 (N_36581,N_35731,N_35376);
or U36582 (N_36582,N_35870,N_35413);
nor U36583 (N_36583,N_35614,N_35840);
nand U36584 (N_36584,N_35762,N_35329);
and U36585 (N_36585,N_35881,N_35020);
or U36586 (N_36586,N_35182,N_35441);
xnor U36587 (N_36587,N_35318,N_35159);
nor U36588 (N_36588,N_35074,N_35822);
nand U36589 (N_36589,N_35297,N_35574);
xnor U36590 (N_36590,N_35297,N_35715);
and U36591 (N_36591,N_35461,N_35877);
xnor U36592 (N_36592,N_35972,N_35733);
nor U36593 (N_36593,N_35235,N_35945);
nor U36594 (N_36594,N_35360,N_35776);
nor U36595 (N_36595,N_35242,N_35290);
or U36596 (N_36596,N_35580,N_35790);
xor U36597 (N_36597,N_35569,N_35457);
and U36598 (N_36598,N_35566,N_35753);
or U36599 (N_36599,N_35054,N_35067);
nor U36600 (N_36600,N_35874,N_35689);
nor U36601 (N_36601,N_35494,N_35819);
nor U36602 (N_36602,N_35474,N_35175);
nand U36603 (N_36603,N_35082,N_35466);
nor U36604 (N_36604,N_35276,N_35762);
nor U36605 (N_36605,N_35471,N_35102);
nand U36606 (N_36606,N_35285,N_35008);
or U36607 (N_36607,N_35622,N_35654);
xor U36608 (N_36608,N_35408,N_35964);
nand U36609 (N_36609,N_35460,N_35277);
nor U36610 (N_36610,N_35314,N_35007);
xnor U36611 (N_36611,N_35077,N_35263);
nor U36612 (N_36612,N_35988,N_35975);
and U36613 (N_36613,N_35037,N_35171);
or U36614 (N_36614,N_35328,N_35221);
and U36615 (N_36615,N_35113,N_35150);
nand U36616 (N_36616,N_35155,N_35114);
nor U36617 (N_36617,N_35967,N_35970);
xnor U36618 (N_36618,N_35578,N_35082);
nand U36619 (N_36619,N_35547,N_35151);
nor U36620 (N_36620,N_35794,N_35532);
nor U36621 (N_36621,N_35940,N_35772);
and U36622 (N_36622,N_35502,N_35892);
nand U36623 (N_36623,N_35265,N_35512);
or U36624 (N_36624,N_35447,N_35755);
or U36625 (N_36625,N_35498,N_35706);
nand U36626 (N_36626,N_35466,N_35170);
and U36627 (N_36627,N_35157,N_35485);
or U36628 (N_36628,N_35201,N_35975);
and U36629 (N_36629,N_35608,N_35090);
and U36630 (N_36630,N_35214,N_35799);
nand U36631 (N_36631,N_35703,N_35191);
nor U36632 (N_36632,N_35202,N_35211);
nor U36633 (N_36633,N_35043,N_35382);
nor U36634 (N_36634,N_35959,N_35470);
and U36635 (N_36635,N_35095,N_35202);
nor U36636 (N_36636,N_35706,N_35097);
or U36637 (N_36637,N_35213,N_35671);
nor U36638 (N_36638,N_35941,N_35510);
and U36639 (N_36639,N_35202,N_35061);
nand U36640 (N_36640,N_35825,N_35289);
xnor U36641 (N_36641,N_35054,N_35303);
nor U36642 (N_36642,N_35558,N_35244);
xnor U36643 (N_36643,N_35851,N_35270);
nor U36644 (N_36644,N_35658,N_35418);
nand U36645 (N_36645,N_35012,N_35676);
and U36646 (N_36646,N_35009,N_35241);
or U36647 (N_36647,N_35326,N_35754);
nand U36648 (N_36648,N_35391,N_35461);
nor U36649 (N_36649,N_35862,N_35285);
nand U36650 (N_36650,N_35903,N_35136);
xnor U36651 (N_36651,N_35768,N_35305);
nor U36652 (N_36652,N_35479,N_35095);
or U36653 (N_36653,N_35063,N_35124);
nor U36654 (N_36654,N_35706,N_35868);
xnor U36655 (N_36655,N_35419,N_35930);
xor U36656 (N_36656,N_35362,N_35031);
nand U36657 (N_36657,N_35195,N_35504);
or U36658 (N_36658,N_35156,N_35810);
xor U36659 (N_36659,N_35051,N_35819);
and U36660 (N_36660,N_35827,N_35636);
xnor U36661 (N_36661,N_35354,N_35311);
xnor U36662 (N_36662,N_35628,N_35033);
nand U36663 (N_36663,N_35371,N_35149);
or U36664 (N_36664,N_35600,N_35696);
nand U36665 (N_36665,N_35114,N_35818);
nand U36666 (N_36666,N_35760,N_35778);
nor U36667 (N_36667,N_35853,N_35254);
nand U36668 (N_36668,N_35141,N_35186);
nand U36669 (N_36669,N_35095,N_35425);
nor U36670 (N_36670,N_35405,N_35186);
nand U36671 (N_36671,N_35897,N_35652);
nand U36672 (N_36672,N_35096,N_35049);
or U36673 (N_36673,N_35686,N_35724);
xnor U36674 (N_36674,N_35179,N_35463);
nand U36675 (N_36675,N_35282,N_35904);
and U36676 (N_36676,N_35889,N_35491);
or U36677 (N_36677,N_35190,N_35370);
xor U36678 (N_36678,N_35534,N_35344);
nand U36679 (N_36679,N_35752,N_35005);
nor U36680 (N_36680,N_35371,N_35977);
or U36681 (N_36681,N_35898,N_35576);
nand U36682 (N_36682,N_35384,N_35489);
or U36683 (N_36683,N_35090,N_35773);
and U36684 (N_36684,N_35247,N_35184);
and U36685 (N_36685,N_35278,N_35332);
or U36686 (N_36686,N_35573,N_35967);
and U36687 (N_36687,N_35207,N_35967);
and U36688 (N_36688,N_35407,N_35189);
nand U36689 (N_36689,N_35640,N_35589);
or U36690 (N_36690,N_35056,N_35359);
nor U36691 (N_36691,N_35208,N_35838);
xnor U36692 (N_36692,N_35203,N_35141);
nand U36693 (N_36693,N_35245,N_35924);
or U36694 (N_36694,N_35994,N_35841);
nand U36695 (N_36695,N_35188,N_35235);
or U36696 (N_36696,N_35425,N_35490);
xor U36697 (N_36697,N_35182,N_35481);
xnor U36698 (N_36698,N_35773,N_35114);
nand U36699 (N_36699,N_35092,N_35319);
or U36700 (N_36700,N_35201,N_35475);
and U36701 (N_36701,N_35014,N_35136);
and U36702 (N_36702,N_35679,N_35011);
xnor U36703 (N_36703,N_35148,N_35838);
nor U36704 (N_36704,N_35250,N_35957);
xor U36705 (N_36705,N_35402,N_35315);
nor U36706 (N_36706,N_35842,N_35819);
xnor U36707 (N_36707,N_35934,N_35543);
nor U36708 (N_36708,N_35491,N_35797);
or U36709 (N_36709,N_35784,N_35859);
nor U36710 (N_36710,N_35854,N_35602);
nor U36711 (N_36711,N_35993,N_35860);
and U36712 (N_36712,N_35131,N_35876);
nor U36713 (N_36713,N_35873,N_35552);
nor U36714 (N_36714,N_35323,N_35371);
and U36715 (N_36715,N_35874,N_35302);
or U36716 (N_36716,N_35410,N_35951);
xor U36717 (N_36717,N_35150,N_35651);
nor U36718 (N_36718,N_35774,N_35143);
xor U36719 (N_36719,N_35731,N_35462);
xnor U36720 (N_36720,N_35756,N_35416);
or U36721 (N_36721,N_35806,N_35787);
and U36722 (N_36722,N_35297,N_35852);
nand U36723 (N_36723,N_35485,N_35946);
and U36724 (N_36724,N_35045,N_35682);
nor U36725 (N_36725,N_35566,N_35207);
and U36726 (N_36726,N_35317,N_35716);
nand U36727 (N_36727,N_35168,N_35505);
nand U36728 (N_36728,N_35584,N_35882);
xnor U36729 (N_36729,N_35040,N_35390);
nor U36730 (N_36730,N_35953,N_35454);
xor U36731 (N_36731,N_35253,N_35020);
nand U36732 (N_36732,N_35627,N_35850);
xnor U36733 (N_36733,N_35750,N_35845);
nand U36734 (N_36734,N_35476,N_35008);
nand U36735 (N_36735,N_35798,N_35304);
and U36736 (N_36736,N_35715,N_35532);
or U36737 (N_36737,N_35081,N_35054);
nor U36738 (N_36738,N_35205,N_35974);
or U36739 (N_36739,N_35054,N_35903);
nor U36740 (N_36740,N_35515,N_35444);
and U36741 (N_36741,N_35053,N_35784);
xnor U36742 (N_36742,N_35432,N_35973);
or U36743 (N_36743,N_35924,N_35143);
xor U36744 (N_36744,N_35987,N_35462);
nor U36745 (N_36745,N_35191,N_35138);
xnor U36746 (N_36746,N_35282,N_35774);
xnor U36747 (N_36747,N_35374,N_35734);
or U36748 (N_36748,N_35926,N_35726);
and U36749 (N_36749,N_35934,N_35383);
nand U36750 (N_36750,N_35501,N_35049);
and U36751 (N_36751,N_35622,N_35644);
nand U36752 (N_36752,N_35297,N_35020);
xnor U36753 (N_36753,N_35534,N_35047);
or U36754 (N_36754,N_35408,N_35462);
and U36755 (N_36755,N_35873,N_35693);
or U36756 (N_36756,N_35863,N_35440);
and U36757 (N_36757,N_35909,N_35419);
nand U36758 (N_36758,N_35327,N_35993);
nor U36759 (N_36759,N_35282,N_35630);
nor U36760 (N_36760,N_35433,N_35529);
nor U36761 (N_36761,N_35465,N_35858);
nand U36762 (N_36762,N_35001,N_35561);
and U36763 (N_36763,N_35338,N_35466);
nor U36764 (N_36764,N_35404,N_35898);
or U36765 (N_36765,N_35418,N_35078);
xnor U36766 (N_36766,N_35857,N_35899);
xor U36767 (N_36767,N_35269,N_35170);
or U36768 (N_36768,N_35117,N_35556);
nor U36769 (N_36769,N_35126,N_35612);
and U36770 (N_36770,N_35465,N_35319);
xnor U36771 (N_36771,N_35345,N_35262);
or U36772 (N_36772,N_35766,N_35408);
and U36773 (N_36773,N_35126,N_35851);
nand U36774 (N_36774,N_35635,N_35658);
nor U36775 (N_36775,N_35172,N_35448);
and U36776 (N_36776,N_35608,N_35954);
nand U36777 (N_36777,N_35566,N_35557);
nor U36778 (N_36778,N_35141,N_35052);
nor U36779 (N_36779,N_35397,N_35777);
and U36780 (N_36780,N_35938,N_35139);
nor U36781 (N_36781,N_35960,N_35923);
or U36782 (N_36782,N_35620,N_35305);
and U36783 (N_36783,N_35954,N_35551);
xnor U36784 (N_36784,N_35345,N_35601);
or U36785 (N_36785,N_35549,N_35669);
and U36786 (N_36786,N_35191,N_35392);
xor U36787 (N_36787,N_35644,N_35819);
or U36788 (N_36788,N_35511,N_35568);
and U36789 (N_36789,N_35830,N_35144);
nor U36790 (N_36790,N_35010,N_35004);
or U36791 (N_36791,N_35185,N_35751);
nor U36792 (N_36792,N_35840,N_35692);
nand U36793 (N_36793,N_35577,N_35969);
xor U36794 (N_36794,N_35006,N_35756);
and U36795 (N_36795,N_35025,N_35260);
xnor U36796 (N_36796,N_35696,N_35416);
or U36797 (N_36797,N_35671,N_35714);
nand U36798 (N_36798,N_35441,N_35422);
nor U36799 (N_36799,N_35783,N_35239);
xor U36800 (N_36800,N_35450,N_35065);
nand U36801 (N_36801,N_35169,N_35117);
or U36802 (N_36802,N_35822,N_35368);
nand U36803 (N_36803,N_35945,N_35366);
xor U36804 (N_36804,N_35371,N_35633);
and U36805 (N_36805,N_35426,N_35685);
nand U36806 (N_36806,N_35137,N_35959);
nor U36807 (N_36807,N_35291,N_35769);
xor U36808 (N_36808,N_35783,N_35215);
nand U36809 (N_36809,N_35838,N_35146);
nor U36810 (N_36810,N_35399,N_35810);
nor U36811 (N_36811,N_35176,N_35805);
nand U36812 (N_36812,N_35249,N_35298);
and U36813 (N_36813,N_35881,N_35258);
xor U36814 (N_36814,N_35990,N_35725);
xor U36815 (N_36815,N_35856,N_35242);
or U36816 (N_36816,N_35607,N_35732);
and U36817 (N_36817,N_35841,N_35418);
nand U36818 (N_36818,N_35059,N_35012);
xor U36819 (N_36819,N_35726,N_35635);
xor U36820 (N_36820,N_35645,N_35004);
nor U36821 (N_36821,N_35291,N_35979);
nor U36822 (N_36822,N_35289,N_35829);
or U36823 (N_36823,N_35020,N_35555);
and U36824 (N_36824,N_35818,N_35361);
nand U36825 (N_36825,N_35985,N_35494);
xor U36826 (N_36826,N_35135,N_35596);
or U36827 (N_36827,N_35346,N_35820);
or U36828 (N_36828,N_35338,N_35233);
nor U36829 (N_36829,N_35756,N_35004);
nor U36830 (N_36830,N_35867,N_35377);
and U36831 (N_36831,N_35761,N_35744);
nor U36832 (N_36832,N_35323,N_35376);
and U36833 (N_36833,N_35752,N_35837);
and U36834 (N_36834,N_35180,N_35207);
nor U36835 (N_36835,N_35612,N_35032);
xor U36836 (N_36836,N_35817,N_35949);
nor U36837 (N_36837,N_35496,N_35282);
nor U36838 (N_36838,N_35814,N_35513);
nand U36839 (N_36839,N_35369,N_35806);
nor U36840 (N_36840,N_35907,N_35630);
nand U36841 (N_36841,N_35204,N_35782);
or U36842 (N_36842,N_35257,N_35097);
and U36843 (N_36843,N_35303,N_35591);
xor U36844 (N_36844,N_35296,N_35039);
nor U36845 (N_36845,N_35955,N_35180);
nand U36846 (N_36846,N_35418,N_35032);
and U36847 (N_36847,N_35572,N_35407);
and U36848 (N_36848,N_35348,N_35418);
or U36849 (N_36849,N_35912,N_35502);
and U36850 (N_36850,N_35488,N_35952);
xor U36851 (N_36851,N_35076,N_35336);
xor U36852 (N_36852,N_35878,N_35306);
and U36853 (N_36853,N_35307,N_35193);
or U36854 (N_36854,N_35248,N_35557);
and U36855 (N_36855,N_35619,N_35295);
nor U36856 (N_36856,N_35634,N_35367);
or U36857 (N_36857,N_35779,N_35858);
xnor U36858 (N_36858,N_35690,N_35421);
or U36859 (N_36859,N_35934,N_35846);
nand U36860 (N_36860,N_35345,N_35930);
nand U36861 (N_36861,N_35042,N_35122);
nand U36862 (N_36862,N_35913,N_35808);
nand U36863 (N_36863,N_35594,N_35694);
nor U36864 (N_36864,N_35779,N_35235);
nor U36865 (N_36865,N_35736,N_35149);
nand U36866 (N_36866,N_35255,N_35679);
nor U36867 (N_36867,N_35176,N_35731);
and U36868 (N_36868,N_35903,N_35012);
nor U36869 (N_36869,N_35573,N_35318);
xor U36870 (N_36870,N_35679,N_35135);
nor U36871 (N_36871,N_35077,N_35929);
xor U36872 (N_36872,N_35236,N_35801);
and U36873 (N_36873,N_35648,N_35566);
or U36874 (N_36874,N_35666,N_35915);
nand U36875 (N_36875,N_35318,N_35708);
xnor U36876 (N_36876,N_35720,N_35480);
xnor U36877 (N_36877,N_35904,N_35754);
nor U36878 (N_36878,N_35793,N_35226);
xor U36879 (N_36879,N_35814,N_35065);
nor U36880 (N_36880,N_35435,N_35969);
xor U36881 (N_36881,N_35875,N_35270);
or U36882 (N_36882,N_35737,N_35285);
nand U36883 (N_36883,N_35555,N_35286);
nand U36884 (N_36884,N_35788,N_35197);
nand U36885 (N_36885,N_35191,N_35372);
nor U36886 (N_36886,N_35954,N_35614);
or U36887 (N_36887,N_35762,N_35976);
and U36888 (N_36888,N_35975,N_35497);
and U36889 (N_36889,N_35797,N_35138);
nor U36890 (N_36890,N_35465,N_35690);
xor U36891 (N_36891,N_35122,N_35513);
or U36892 (N_36892,N_35416,N_35952);
nor U36893 (N_36893,N_35294,N_35432);
xor U36894 (N_36894,N_35939,N_35104);
nor U36895 (N_36895,N_35000,N_35167);
nor U36896 (N_36896,N_35002,N_35443);
xor U36897 (N_36897,N_35019,N_35414);
xnor U36898 (N_36898,N_35858,N_35109);
nor U36899 (N_36899,N_35415,N_35259);
or U36900 (N_36900,N_35515,N_35036);
or U36901 (N_36901,N_35651,N_35212);
or U36902 (N_36902,N_35984,N_35267);
nand U36903 (N_36903,N_35504,N_35182);
and U36904 (N_36904,N_35231,N_35250);
xnor U36905 (N_36905,N_35848,N_35413);
nor U36906 (N_36906,N_35736,N_35318);
nor U36907 (N_36907,N_35616,N_35787);
xnor U36908 (N_36908,N_35533,N_35539);
or U36909 (N_36909,N_35351,N_35508);
nor U36910 (N_36910,N_35208,N_35786);
xor U36911 (N_36911,N_35609,N_35764);
nand U36912 (N_36912,N_35232,N_35514);
and U36913 (N_36913,N_35842,N_35630);
or U36914 (N_36914,N_35534,N_35513);
or U36915 (N_36915,N_35187,N_35876);
nor U36916 (N_36916,N_35887,N_35043);
or U36917 (N_36917,N_35398,N_35167);
and U36918 (N_36918,N_35776,N_35841);
or U36919 (N_36919,N_35668,N_35568);
nor U36920 (N_36920,N_35179,N_35187);
or U36921 (N_36921,N_35759,N_35584);
and U36922 (N_36922,N_35631,N_35963);
nand U36923 (N_36923,N_35800,N_35133);
xor U36924 (N_36924,N_35170,N_35984);
nand U36925 (N_36925,N_35510,N_35311);
or U36926 (N_36926,N_35308,N_35713);
nand U36927 (N_36927,N_35969,N_35332);
and U36928 (N_36928,N_35366,N_35587);
and U36929 (N_36929,N_35176,N_35503);
nand U36930 (N_36930,N_35301,N_35064);
nor U36931 (N_36931,N_35718,N_35915);
xnor U36932 (N_36932,N_35848,N_35658);
nand U36933 (N_36933,N_35243,N_35357);
xnor U36934 (N_36934,N_35590,N_35821);
or U36935 (N_36935,N_35457,N_35385);
nand U36936 (N_36936,N_35432,N_35628);
and U36937 (N_36937,N_35278,N_35042);
xnor U36938 (N_36938,N_35676,N_35076);
or U36939 (N_36939,N_35576,N_35532);
nor U36940 (N_36940,N_35739,N_35108);
and U36941 (N_36941,N_35820,N_35192);
nand U36942 (N_36942,N_35973,N_35131);
nor U36943 (N_36943,N_35664,N_35765);
and U36944 (N_36944,N_35125,N_35833);
nand U36945 (N_36945,N_35760,N_35361);
xor U36946 (N_36946,N_35007,N_35196);
nand U36947 (N_36947,N_35624,N_35155);
xor U36948 (N_36948,N_35194,N_35367);
and U36949 (N_36949,N_35580,N_35873);
nor U36950 (N_36950,N_35621,N_35706);
and U36951 (N_36951,N_35690,N_35491);
nand U36952 (N_36952,N_35303,N_35926);
or U36953 (N_36953,N_35646,N_35881);
and U36954 (N_36954,N_35862,N_35102);
nor U36955 (N_36955,N_35132,N_35015);
and U36956 (N_36956,N_35399,N_35072);
or U36957 (N_36957,N_35070,N_35764);
and U36958 (N_36958,N_35259,N_35665);
and U36959 (N_36959,N_35379,N_35967);
or U36960 (N_36960,N_35982,N_35146);
or U36961 (N_36961,N_35295,N_35285);
nand U36962 (N_36962,N_35533,N_35760);
nor U36963 (N_36963,N_35534,N_35602);
nor U36964 (N_36964,N_35266,N_35696);
or U36965 (N_36965,N_35433,N_35198);
xor U36966 (N_36966,N_35283,N_35613);
nand U36967 (N_36967,N_35240,N_35528);
or U36968 (N_36968,N_35245,N_35596);
xnor U36969 (N_36969,N_35585,N_35337);
xnor U36970 (N_36970,N_35454,N_35201);
or U36971 (N_36971,N_35632,N_35307);
and U36972 (N_36972,N_35026,N_35512);
nand U36973 (N_36973,N_35654,N_35308);
nor U36974 (N_36974,N_35593,N_35065);
nand U36975 (N_36975,N_35972,N_35351);
and U36976 (N_36976,N_35773,N_35565);
or U36977 (N_36977,N_35870,N_35254);
or U36978 (N_36978,N_35660,N_35059);
and U36979 (N_36979,N_35672,N_35353);
xnor U36980 (N_36980,N_35316,N_35185);
and U36981 (N_36981,N_35831,N_35936);
xor U36982 (N_36982,N_35736,N_35935);
nor U36983 (N_36983,N_35841,N_35629);
or U36984 (N_36984,N_35766,N_35670);
nor U36985 (N_36985,N_35952,N_35036);
and U36986 (N_36986,N_35421,N_35633);
and U36987 (N_36987,N_35413,N_35038);
nand U36988 (N_36988,N_35967,N_35646);
nor U36989 (N_36989,N_35738,N_35180);
nor U36990 (N_36990,N_35730,N_35918);
and U36991 (N_36991,N_35481,N_35567);
xnor U36992 (N_36992,N_35806,N_35611);
nand U36993 (N_36993,N_35805,N_35527);
nor U36994 (N_36994,N_35736,N_35475);
or U36995 (N_36995,N_35390,N_35399);
and U36996 (N_36996,N_35515,N_35985);
nor U36997 (N_36997,N_35216,N_35336);
xnor U36998 (N_36998,N_35881,N_35380);
nor U36999 (N_36999,N_35953,N_35324);
and U37000 (N_37000,N_36867,N_36295);
nor U37001 (N_37001,N_36610,N_36501);
nor U37002 (N_37002,N_36690,N_36017);
or U37003 (N_37003,N_36891,N_36816);
and U37004 (N_37004,N_36351,N_36492);
nor U37005 (N_37005,N_36794,N_36776);
or U37006 (N_37006,N_36222,N_36323);
nand U37007 (N_37007,N_36919,N_36881);
and U37008 (N_37008,N_36616,N_36317);
or U37009 (N_37009,N_36280,N_36830);
nand U37010 (N_37010,N_36143,N_36694);
xor U37011 (N_37011,N_36325,N_36730);
nor U37012 (N_37012,N_36927,N_36573);
nor U37013 (N_37013,N_36402,N_36117);
or U37014 (N_37014,N_36487,N_36465);
nand U37015 (N_37015,N_36734,N_36807);
nor U37016 (N_37016,N_36532,N_36828);
nand U37017 (N_37017,N_36874,N_36952);
xnor U37018 (N_37018,N_36498,N_36368);
nor U37019 (N_37019,N_36126,N_36844);
or U37020 (N_37020,N_36750,N_36618);
nor U37021 (N_37021,N_36561,N_36588);
and U37022 (N_37022,N_36652,N_36053);
or U37023 (N_37023,N_36739,N_36803);
nor U37024 (N_37024,N_36673,N_36175);
nor U37025 (N_37025,N_36084,N_36507);
nand U37026 (N_37026,N_36451,N_36626);
nor U37027 (N_37027,N_36068,N_36591);
or U37028 (N_37028,N_36050,N_36130);
nor U37029 (N_37029,N_36493,N_36788);
nor U37030 (N_37030,N_36944,N_36847);
xnor U37031 (N_37031,N_36306,N_36703);
and U37032 (N_37032,N_36848,N_36202);
xnor U37033 (N_37033,N_36283,N_36406);
and U37034 (N_37034,N_36933,N_36934);
and U37035 (N_37035,N_36634,N_36504);
nand U37036 (N_37036,N_36370,N_36288);
and U37037 (N_37037,N_36369,N_36834);
and U37038 (N_37038,N_36420,N_36469);
nor U37039 (N_37039,N_36007,N_36954);
and U37040 (N_37040,N_36430,N_36333);
or U37041 (N_37041,N_36679,N_36005);
or U37042 (N_37042,N_36411,N_36015);
xor U37043 (N_37043,N_36965,N_36581);
or U37044 (N_37044,N_36708,N_36879);
and U37045 (N_37045,N_36461,N_36963);
and U37046 (N_37046,N_36232,N_36884);
xnor U37047 (N_37047,N_36820,N_36653);
nor U37048 (N_37048,N_36531,N_36990);
nand U37049 (N_37049,N_36211,N_36003);
or U37050 (N_37050,N_36758,N_36320);
nor U37051 (N_37051,N_36046,N_36726);
xor U37052 (N_37052,N_36772,N_36304);
nand U37053 (N_37053,N_36100,N_36332);
or U37054 (N_37054,N_36725,N_36782);
or U37055 (N_37055,N_36253,N_36098);
or U37056 (N_37056,N_36960,N_36548);
or U37057 (N_37057,N_36227,N_36199);
xnor U37058 (N_37058,N_36571,N_36900);
xor U37059 (N_37059,N_36145,N_36951);
xor U37060 (N_37060,N_36310,N_36683);
nor U37061 (N_37061,N_36208,N_36804);
and U37062 (N_37062,N_36414,N_36206);
xnor U37063 (N_37063,N_36519,N_36181);
nor U37064 (N_37064,N_36836,N_36045);
or U37065 (N_37065,N_36685,N_36445);
nor U37066 (N_37066,N_36632,N_36104);
and U37067 (N_37067,N_36404,N_36686);
or U37068 (N_37068,N_36291,N_36779);
or U37069 (N_37069,N_36715,N_36854);
or U37070 (N_37070,N_36355,N_36247);
xnor U37071 (N_37071,N_36521,N_36264);
or U37072 (N_37072,N_36929,N_36850);
and U37073 (N_37073,N_36274,N_36584);
or U37074 (N_37074,N_36378,N_36946);
nand U37075 (N_37075,N_36322,N_36853);
or U37076 (N_37076,N_36263,N_36416);
and U37077 (N_37077,N_36078,N_36517);
nand U37078 (N_37078,N_36550,N_36284);
or U37079 (N_37079,N_36641,N_36137);
and U37080 (N_37080,N_36440,N_36043);
and U37081 (N_37081,N_36585,N_36379);
nor U37082 (N_37082,N_36949,N_36637);
nor U37083 (N_37083,N_36018,N_36747);
nor U37084 (N_37084,N_36169,N_36497);
nor U37085 (N_37085,N_36470,N_36059);
or U37086 (N_37086,N_36133,N_36185);
nand U37087 (N_37087,N_36760,N_36530);
and U37088 (N_37088,N_36062,N_36873);
nand U37089 (N_37089,N_36866,N_36156);
xnor U37090 (N_37090,N_36432,N_36869);
and U37091 (N_37091,N_36887,N_36744);
and U37092 (N_37092,N_36533,N_36746);
and U37093 (N_37093,N_36525,N_36364);
and U37094 (N_37094,N_36090,N_36553);
nand U37095 (N_37095,N_36153,N_36657);
nand U37096 (N_37096,N_36871,N_36889);
nor U37097 (N_37097,N_36361,N_36148);
and U37098 (N_37098,N_36347,N_36923);
nand U37099 (N_37099,N_36814,N_36974);
nor U37100 (N_37100,N_36054,N_36796);
xnor U37101 (N_37101,N_36818,N_36051);
and U37102 (N_37102,N_36823,N_36383);
nand U37103 (N_37103,N_36099,N_36462);
xnor U37104 (N_37104,N_36542,N_36987);
nor U37105 (N_37105,N_36700,N_36733);
nand U37106 (N_37106,N_36680,N_36075);
and U37107 (N_37107,N_36736,N_36773);
or U37108 (N_37108,N_36142,N_36729);
nor U37109 (N_37109,N_36862,N_36040);
or U37110 (N_37110,N_36109,N_36431);
or U37111 (N_37111,N_36508,N_36048);
xnor U37112 (N_37112,N_36982,N_36287);
and U37113 (N_37113,N_36556,N_36908);
or U37114 (N_37114,N_36707,N_36036);
xnor U37115 (N_37115,N_36286,N_36030);
and U37116 (N_37116,N_36119,N_36318);
nor U37117 (N_37117,N_36975,N_36904);
or U37118 (N_37118,N_36595,N_36230);
nand U37119 (N_37119,N_36528,N_36204);
and U37120 (N_37120,N_36842,N_36621);
xor U37121 (N_37121,N_36094,N_36745);
or U37122 (N_37122,N_36910,N_36723);
nand U37123 (N_37123,N_36245,N_36833);
or U37124 (N_37124,N_36524,N_36205);
and U37125 (N_37125,N_36356,N_36164);
xnor U37126 (N_37126,N_36695,N_36315);
and U37127 (N_37127,N_36489,N_36234);
nand U37128 (N_37128,N_36254,N_36579);
nand U37129 (N_37129,N_36592,N_36444);
nand U37130 (N_37130,N_36622,N_36631);
nand U37131 (N_37131,N_36165,N_36551);
xor U37132 (N_37132,N_36022,N_36615);
and U37133 (N_37133,N_36924,N_36605);
or U37134 (N_37134,N_36238,N_36226);
nor U37135 (N_37135,N_36486,N_36698);
xor U37136 (N_37136,N_36568,N_36589);
nor U37137 (N_37137,N_36380,N_36895);
nand U37138 (N_37138,N_36638,N_36539);
xnor U37139 (N_37139,N_36429,N_36674);
xor U37140 (N_37140,N_36074,N_36372);
or U37141 (N_37141,N_36768,N_36962);
nor U37142 (N_37142,N_36838,N_36738);
xnor U37143 (N_37143,N_36327,N_36063);
or U37144 (N_37144,N_36855,N_36037);
nand U37145 (N_37145,N_36023,N_36650);
nand U37146 (N_37146,N_36986,N_36580);
and U37147 (N_37147,N_36405,N_36308);
nand U37148 (N_37148,N_36473,N_36611);
or U37149 (N_37149,N_36600,N_36565);
nor U37150 (N_37150,N_36968,N_36442);
nor U37151 (N_37151,N_36251,N_36755);
nand U37152 (N_37152,N_36647,N_36623);
and U37153 (N_37153,N_36790,N_36374);
or U37154 (N_37154,N_36464,N_36389);
and U37155 (N_37155,N_36417,N_36192);
xnor U37156 (N_37156,N_36856,N_36116);
and U37157 (N_37157,N_36453,N_36135);
nor U37158 (N_37158,N_36067,N_36147);
and U37159 (N_37159,N_36302,N_36756);
nand U37160 (N_37160,N_36583,N_36179);
xor U37161 (N_37161,N_36049,N_36978);
nor U37162 (N_37162,N_36221,N_36363);
and U37163 (N_37163,N_36696,N_36194);
nand U37164 (N_37164,N_36992,N_36178);
or U37165 (N_37165,N_36780,N_36681);
nand U37166 (N_37166,N_36993,N_36273);
xnor U37167 (N_37167,N_36909,N_36103);
nor U37168 (N_37168,N_36841,N_36307);
xor U37169 (N_37169,N_36984,N_36971);
xnor U37170 (N_37170,N_36961,N_36385);
xor U37171 (N_37171,N_36146,N_36367);
or U37172 (N_37172,N_36223,N_36570);
nand U37173 (N_37173,N_36678,N_36025);
nor U37174 (N_37174,N_36705,N_36651);
or U37175 (N_37175,N_36233,N_36603);
and U37176 (N_37176,N_36159,N_36382);
nor U37177 (N_37177,N_36316,N_36460);
xnor U37178 (N_37178,N_36922,N_36477);
nand U37179 (N_37179,N_36475,N_36012);
or U37180 (N_37180,N_36256,N_36265);
nor U37181 (N_37181,N_36170,N_36242);
or U37182 (N_37182,N_36764,N_36885);
or U37183 (N_37183,N_36035,N_36714);
xor U37184 (N_37184,N_36294,N_36858);
and U37185 (N_37185,N_36576,N_36391);
nand U37186 (N_37186,N_36193,N_36536);
or U37187 (N_37187,N_36502,N_36371);
nand U37188 (N_37188,N_36267,N_36888);
nor U37189 (N_37189,N_36709,N_36912);
and U37190 (N_37190,N_36898,N_36518);
and U37191 (N_37191,N_36339,N_36452);
nand U37192 (N_37192,N_36947,N_36200);
nor U37193 (N_37193,N_36625,N_36795);
or U37194 (N_37194,N_36218,N_36161);
xor U37195 (N_37195,N_36289,N_36645);
nor U37196 (N_37196,N_36976,N_36552);
nor U37197 (N_37197,N_36311,N_36813);
nand U37198 (N_37198,N_36967,N_36829);
and U37199 (N_37199,N_36476,N_36825);
and U37200 (N_37200,N_36753,N_36138);
nand U37201 (N_37201,N_36352,N_36914);
nand U37202 (N_37202,N_36213,N_36127);
nand U37203 (N_37203,N_36152,N_36071);
xnor U37204 (N_37204,N_36546,N_36029);
nor U37205 (N_37205,N_36314,N_36044);
and U37206 (N_37206,N_36666,N_36831);
xor U37207 (N_37207,N_36643,N_36168);
and U37208 (N_37208,N_36207,N_36506);
and U37209 (N_37209,N_36697,N_36281);
and U37210 (N_37210,N_36996,N_36824);
and U37211 (N_37211,N_36184,N_36392);
or U37212 (N_37212,N_36977,N_36056);
and U37213 (N_37213,N_36627,N_36878);
or U37214 (N_37214,N_36344,N_36742);
and U37215 (N_37215,N_36991,N_36896);
nand U37216 (N_37216,N_36144,N_36203);
or U37217 (N_37217,N_36341,N_36549);
xor U37218 (N_37218,N_36220,N_36636);
and U37219 (N_37219,N_36935,N_36166);
xor U37220 (N_37220,N_36481,N_36886);
and U37221 (N_37221,N_36587,N_36437);
xor U37222 (N_37222,N_36474,N_36959);
xor U37223 (N_37223,N_36375,N_36102);
and U37224 (N_37224,N_36120,N_36767);
nand U37225 (N_37225,N_36901,N_36198);
nand U37226 (N_37226,N_36268,N_36937);
or U37227 (N_37227,N_36926,N_36249);
nor U37228 (N_37228,N_36279,N_36132);
or U37229 (N_37229,N_36248,N_36224);
xor U37230 (N_37230,N_36969,N_36956);
nor U37231 (N_37231,N_36513,N_36649);
nand U37232 (N_37232,N_36598,N_36483);
xnor U37233 (N_37233,N_36210,N_36523);
or U37234 (N_37234,N_36309,N_36938);
and U37235 (N_37235,N_36269,N_36069);
and U37236 (N_37236,N_36763,N_36365);
nor U37237 (N_37237,N_36010,N_36731);
and U37238 (N_37238,N_36073,N_36512);
xnor U37239 (N_37239,N_36577,N_36943);
nor U37240 (N_37240,N_36122,N_36157);
xor U37241 (N_37241,N_36957,N_36418);
and U37242 (N_37242,N_36630,N_36260);
or U37243 (N_37243,N_36865,N_36660);
nand U37244 (N_37244,N_36907,N_36435);
or U37245 (N_37245,N_36955,N_36290);
and U37246 (N_37246,N_36353,N_36270);
and U37247 (N_37247,N_36136,N_36154);
and U37248 (N_37248,N_36762,N_36628);
xnor U37249 (N_37249,N_36262,N_36711);
or U37250 (N_37250,N_36097,N_36413);
nand U37251 (N_37251,N_36401,N_36663);
nor U37252 (N_37252,N_36540,N_36409);
xnor U37253 (N_37253,N_36348,N_36761);
xnor U37254 (N_37254,N_36032,N_36123);
nor U37255 (N_37255,N_36384,N_36293);
nor U37256 (N_37256,N_36349,N_36272);
or U37257 (N_37257,N_36151,N_36303);
nor U37258 (N_37258,N_36601,N_36484);
or U37259 (N_37259,N_36713,N_36387);
nor U37260 (N_37260,N_36520,N_36002);
and U37261 (N_37261,N_36196,N_36607);
and U37262 (N_37262,N_36602,N_36438);
nor U37263 (N_37263,N_36390,N_36070);
and U37264 (N_37264,N_36875,N_36215);
nor U37265 (N_37265,N_36691,N_36061);
nor U37266 (N_37266,N_36769,N_36160);
nor U37267 (N_37267,N_36225,N_36633);
nand U37268 (N_37268,N_36244,N_36766);
and U37269 (N_37269,N_36613,N_36083);
nor U37270 (N_37270,N_36671,N_36500);
xor U37271 (N_37271,N_36155,N_36080);
xor U37272 (N_37272,N_36522,N_36899);
and U37273 (N_37273,N_36011,N_36282);
nand U37274 (N_37274,N_36942,N_36183);
nor U37275 (N_37275,N_36350,N_36743);
xor U37276 (N_37276,N_36190,N_36134);
xor U37277 (N_37277,N_36271,N_36024);
and U37278 (N_37278,N_36876,N_36792);
nor U37279 (N_37279,N_36342,N_36863);
xor U37280 (N_37280,N_36688,N_36091);
xnor U37281 (N_37281,N_36751,N_36994);
xnor U37282 (N_37282,N_36981,N_36689);
xor U37283 (N_37283,N_36042,N_36459);
or U37284 (N_37284,N_36027,N_36261);
and U37285 (N_37285,N_36988,N_36354);
nand U37286 (N_37286,N_36543,N_36737);
nor U37287 (N_37287,N_36216,N_36490);
nor U37288 (N_37288,N_36276,N_36920);
nor U37289 (N_37289,N_36236,N_36574);
xor U37290 (N_37290,N_36827,N_36789);
xnor U37291 (N_37291,N_36423,N_36381);
nor U37292 (N_37292,N_36659,N_36106);
and U37293 (N_37293,N_36259,N_36357);
or U37294 (N_37294,N_36554,N_36403);
nor U37295 (N_37295,N_36958,N_36336);
xnor U37296 (N_37296,N_36692,N_36687);
nand U37297 (N_37297,N_36456,N_36212);
nor U37298 (N_37298,N_36101,N_36439);
nor U37299 (N_37299,N_36640,N_36243);
and U37300 (N_37300,N_36534,N_36324);
or U37301 (N_37301,N_36408,N_36433);
and U37302 (N_37302,N_36826,N_36578);
and U37303 (N_37303,N_36089,N_36400);
and U37304 (N_37304,N_36412,N_36038);
xnor U37305 (N_37305,N_36979,N_36458);
and U37306 (N_37306,N_36020,N_36706);
nor U37307 (N_37307,N_36906,N_36079);
xnor U37308 (N_37308,N_36864,N_36559);
nand U37309 (N_37309,N_36593,N_36511);
nand U37310 (N_37310,N_36077,N_36187);
and U37311 (N_37311,N_36677,N_36158);
or U37312 (N_37312,N_36599,N_36092);
xnor U37313 (N_37313,N_36407,N_36312);
xor U37314 (N_37314,N_36802,N_36699);
xnor U37315 (N_37315,N_36340,N_36941);
nand U37316 (N_37316,N_36052,N_36441);
nand U37317 (N_37317,N_36890,N_36376);
xor U37318 (N_37318,N_36514,N_36060);
nand U37319 (N_37319,N_36195,N_36781);
nor U37320 (N_37320,N_36008,N_36572);
nand U37321 (N_37321,N_36893,N_36031);
or U37322 (N_37322,N_36180,N_36110);
xnor U37323 (N_37323,N_36569,N_36149);
nor U37324 (N_37324,N_36805,N_36921);
nor U37325 (N_37325,N_36778,N_36877);
nand U37326 (N_37326,N_36845,N_36811);
nand U37327 (N_37327,N_36292,N_36016);
xnor U37328 (N_37328,N_36426,N_36837);
and U37329 (N_37329,N_36614,N_36727);
nor U37330 (N_37330,N_36278,N_36125);
xor U37331 (N_37331,N_36812,N_36188);
and U37332 (N_37332,N_36467,N_36173);
or U37333 (N_37333,N_36594,N_36197);
nor U37334 (N_37334,N_36801,N_36620);
and U37335 (N_37335,N_36819,N_36480);
and U37336 (N_37336,N_36162,N_36629);
nand U37337 (N_37337,N_36396,N_36646);
nor U37338 (N_37338,N_36735,N_36642);
xor U37339 (N_37339,N_36905,N_36472);
nand U37340 (N_37340,N_36596,N_36201);
nor U37341 (N_37341,N_36186,N_36485);
or U37342 (N_37342,N_36740,N_36980);
or U37343 (N_37343,N_36868,N_36777);
nand U37344 (N_37344,N_36305,N_36930);
or U37345 (N_37345,N_36562,N_36081);
and U37346 (N_37346,N_36606,N_36343);
or U37347 (N_37347,N_36752,N_36377);
xor U37348 (N_37348,N_36466,N_36505);
nand U37349 (N_37349,N_36566,N_36997);
or U37350 (N_37350,N_36085,N_36107);
xnor U37351 (N_37351,N_36373,N_36872);
or U37352 (N_37352,N_36478,N_36034);
xnor U37353 (N_37353,N_36258,N_36076);
or U37354 (N_37354,N_36555,N_36970);
nor U37355 (N_37355,N_36228,N_36301);
nor U37356 (N_37356,N_36721,N_36704);
nand U37357 (N_37357,N_36009,N_36529);
nor U37358 (N_37358,N_36808,N_36182);
nand U37359 (N_37359,N_36928,N_36214);
nand U37360 (N_37360,N_36945,N_36682);
nor U37361 (N_37361,N_36932,N_36006);
nand U37362 (N_37362,N_36880,N_36319);
or U37363 (N_37363,N_36985,N_36167);
xnor U37364 (N_37364,N_36547,N_36774);
nor U37365 (N_37365,N_36112,N_36086);
nand U37366 (N_37366,N_36421,N_36757);
or U37367 (N_37367,N_36998,N_36624);
nand U37368 (N_37368,N_36619,N_36019);
or U37369 (N_37369,N_36821,N_36612);
and U37370 (N_37370,N_36277,N_36939);
xor U37371 (N_37371,N_36668,N_36329);
xnor U37372 (N_37372,N_36915,N_36235);
and U37373 (N_37373,N_36330,N_36499);
xnor U37374 (N_37374,N_36770,N_36299);
or U37375 (N_37375,N_36468,N_36693);
nor U37376 (N_37376,N_36793,N_36172);
nor U37377 (N_37377,N_36503,N_36419);
or U37378 (N_37378,N_36791,N_36118);
xor U37379 (N_37379,N_36732,N_36131);
nor U37380 (N_37380,N_36455,N_36916);
nand U37381 (N_37381,N_36346,N_36973);
nor U37382 (N_37382,N_36093,N_36515);
nor U37383 (N_37383,N_36749,N_36115);
and U37384 (N_37384,N_36257,N_36237);
nand U37385 (N_37385,N_36719,N_36799);
nand U37386 (N_37386,N_36775,N_36014);
nor U37387 (N_37387,N_36718,N_36806);
and U37388 (N_37388,N_36434,N_36150);
nor U37389 (N_37389,N_36328,N_36496);
nor U37390 (N_37390,N_36999,N_36479);
nor U37391 (N_37391,N_36676,N_36717);
nand U37392 (N_37392,N_36388,N_36544);
or U37393 (N_37393,N_36013,N_36360);
and U37394 (N_37394,N_36454,N_36482);
and U37395 (N_37395,N_36443,N_36139);
or U37396 (N_37396,N_36728,N_36004);
nor U37397 (N_37397,N_36298,N_36491);
and U37398 (N_37398,N_36557,N_36564);
nor U37399 (N_37399,N_36000,N_36722);
nor U37400 (N_37400,N_36065,N_36297);
nor U37401 (N_37401,N_36672,N_36447);
nand U37402 (N_37402,N_36966,N_36664);
nand U37403 (N_37403,N_36712,N_36894);
nor U37404 (N_37404,N_36953,N_36658);
nand U37405 (N_37405,N_36702,N_36840);
or U37406 (N_37406,N_36174,N_36424);
and U37407 (N_37407,N_36334,N_36028);
nand U37408 (N_37408,N_36883,N_36798);
nor U37409 (N_37409,N_36141,N_36095);
xor U37410 (N_37410,N_36335,N_36494);
nor U37411 (N_37411,N_36121,N_36140);
or U37412 (N_37412,N_36989,N_36541);
and U37413 (N_37413,N_36033,N_36832);
or U37414 (N_37414,N_36321,N_36058);
xnor U37415 (N_37415,N_36701,N_36537);
xor U37416 (N_37416,N_36285,N_36720);
nor U37417 (N_37417,N_36082,N_36096);
and U37418 (N_37418,N_36582,N_36608);
and U37419 (N_37419,N_36662,N_36001);
nand U37420 (N_37420,N_36545,N_36255);
and U37421 (N_37421,N_36239,N_36724);
xor U37422 (N_37422,N_36538,N_36860);
and U37423 (N_37423,N_36567,N_36846);
or U37424 (N_37424,N_36655,N_36488);
nor U37425 (N_37425,N_36366,N_36563);
nand U37426 (N_37426,N_36331,N_36219);
nand U37427 (N_37427,N_36057,N_36240);
nor U37428 (N_37428,N_36422,N_36415);
nand U37429 (N_37429,N_36326,N_36066);
xnor U37430 (N_37430,N_36670,N_36784);
or U37431 (N_37431,N_36338,N_36797);
xor U37432 (N_37432,N_36635,N_36857);
nand U37433 (N_37433,N_36604,N_36936);
nand U37434 (N_37434,N_36560,N_36463);
or U37435 (N_37435,N_36394,N_36748);
xnor U37436 (N_37436,N_36039,N_36983);
or U37437 (N_37437,N_36189,N_36124);
and U37438 (N_37438,N_36822,N_36710);
and U37439 (N_37439,N_36972,N_36471);
nand U37440 (N_37440,N_36667,N_36800);
nor U37441 (N_37441,N_36558,N_36783);
xnor U37442 (N_37442,N_36948,N_36362);
nor U37443 (N_37443,N_36849,N_36765);
nor U37444 (N_37444,N_36644,N_36105);
nand U37445 (N_37445,N_36231,N_36399);
xor U37446 (N_37446,N_36395,N_36410);
xnor U37447 (N_37447,N_36759,N_36026);
and U37448 (N_37448,N_36918,N_36064);
nand U37449 (N_37449,N_36892,N_36516);
xor U37450 (N_37450,N_36654,N_36171);
nor U37451 (N_37451,N_36510,N_36250);
nand U37452 (N_37452,N_36527,N_36684);
xnor U37453 (N_37453,N_36386,N_36176);
and U37454 (N_37454,N_36785,N_36457);
nor U37455 (N_37455,N_36843,N_36754);
xnor U37456 (N_37456,N_36526,N_36448);
nand U37457 (N_37457,N_36809,N_36656);
nand U37458 (N_37458,N_36397,N_36446);
or U37459 (N_37459,N_36041,N_36449);
and U37460 (N_37460,N_36931,N_36337);
nor U37461 (N_37461,N_36902,N_36897);
nor U37462 (N_37462,N_36427,N_36741);
and U37463 (N_37463,N_36586,N_36590);
and U37464 (N_37464,N_36669,N_36597);
or U37465 (N_37465,N_36639,N_36246);
and U37466 (N_37466,N_36917,N_36810);
or U37467 (N_37467,N_36163,N_36209);
or U37468 (N_37468,N_36911,N_36252);
and U37469 (N_37469,N_36129,N_36913);
nor U37470 (N_37470,N_36114,N_36786);
and U37471 (N_37471,N_36108,N_36425);
or U37472 (N_37472,N_36940,N_36995);
nor U37473 (N_37473,N_36229,N_36436);
or U37474 (N_37474,N_36882,N_36903);
and U37475 (N_37475,N_36870,N_36617);
xnor U37476 (N_37476,N_36217,N_36113);
xnor U37477 (N_37477,N_36111,N_36359);
xnor U37478 (N_37478,N_36839,N_36535);
or U37479 (N_37479,N_36495,N_36313);
or U37480 (N_37480,N_36665,N_36047);
and U37481 (N_37481,N_36398,N_36393);
or U37482 (N_37482,N_36925,N_36771);
or U37483 (N_37483,N_36266,N_36950);
or U37484 (N_37484,N_36191,N_36648);
or U37485 (N_37485,N_36241,N_36815);
nand U37486 (N_37486,N_36358,N_36275);
nor U37487 (N_37487,N_36817,N_36787);
or U37488 (N_37488,N_36609,N_36296);
nand U37489 (N_37489,N_36450,N_36088);
nor U37490 (N_37490,N_36661,N_36087);
nor U37491 (N_37491,N_36851,N_36177);
nand U37492 (N_37492,N_36345,N_36835);
nor U37493 (N_37493,N_36861,N_36675);
xnor U37494 (N_37494,N_36021,N_36072);
and U37495 (N_37495,N_36575,N_36964);
and U37496 (N_37496,N_36509,N_36128);
and U37497 (N_37497,N_36300,N_36852);
xor U37498 (N_37498,N_36055,N_36716);
xor U37499 (N_37499,N_36428,N_36859);
and U37500 (N_37500,N_36997,N_36219);
nor U37501 (N_37501,N_36650,N_36890);
or U37502 (N_37502,N_36104,N_36944);
or U37503 (N_37503,N_36711,N_36339);
or U37504 (N_37504,N_36782,N_36372);
or U37505 (N_37505,N_36581,N_36022);
and U37506 (N_37506,N_36124,N_36318);
xnor U37507 (N_37507,N_36147,N_36907);
nand U37508 (N_37508,N_36557,N_36081);
or U37509 (N_37509,N_36706,N_36092);
nand U37510 (N_37510,N_36934,N_36308);
xnor U37511 (N_37511,N_36034,N_36730);
xor U37512 (N_37512,N_36054,N_36777);
and U37513 (N_37513,N_36186,N_36571);
or U37514 (N_37514,N_36769,N_36946);
and U37515 (N_37515,N_36361,N_36916);
nor U37516 (N_37516,N_36302,N_36121);
nand U37517 (N_37517,N_36872,N_36135);
and U37518 (N_37518,N_36593,N_36103);
xor U37519 (N_37519,N_36538,N_36025);
nand U37520 (N_37520,N_36486,N_36813);
nand U37521 (N_37521,N_36026,N_36436);
and U37522 (N_37522,N_36943,N_36874);
xnor U37523 (N_37523,N_36642,N_36438);
or U37524 (N_37524,N_36668,N_36281);
nand U37525 (N_37525,N_36250,N_36515);
nor U37526 (N_37526,N_36316,N_36193);
nor U37527 (N_37527,N_36267,N_36873);
or U37528 (N_37528,N_36901,N_36114);
xnor U37529 (N_37529,N_36405,N_36547);
or U37530 (N_37530,N_36432,N_36731);
nand U37531 (N_37531,N_36036,N_36135);
nand U37532 (N_37532,N_36625,N_36767);
xor U37533 (N_37533,N_36123,N_36953);
xor U37534 (N_37534,N_36620,N_36366);
nand U37535 (N_37535,N_36082,N_36812);
nor U37536 (N_37536,N_36150,N_36006);
xor U37537 (N_37537,N_36924,N_36123);
nor U37538 (N_37538,N_36594,N_36952);
xor U37539 (N_37539,N_36095,N_36805);
xnor U37540 (N_37540,N_36210,N_36549);
and U37541 (N_37541,N_36470,N_36543);
nand U37542 (N_37542,N_36307,N_36673);
and U37543 (N_37543,N_36437,N_36315);
xnor U37544 (N_37544,N_36983,N_36468);
and U37545 (N_37545,N_36202,N_36404);
xnor U37546 (N_37546,N_36010,N_36688);
or U37547 (N_37547,N_36945,N_36348);
xnor U37548 (N_37548,N_36027,N_36343);
nor U37549 (N_37549,N_36078,N_36672);
nand U37550 (N_37550,N_36762,N_36558);
nor U37551 (N_37551,N_36868,N_36807);
xnor U37552 (N_37552,N_36862,N_36992);
and U37553 (N_37553,N_36933,N_36117);
or U37554 (N_37554,N_36968,N_36099);
or U37555 (N_37555,N_36059,N_36736);
and U37556 (N_37556,N_36184,N_36179);
xnor U37557 (N_37557,N_36126,N_36039);
nand U37558 (N_37558,N_36065,N_36926);
or U37559 (N_37559,N_36950,N_36007);
nor U37560 (N_37560,N_36417,N_36064);
or U37561 (N_37561,N_36067,N_36616);
and U37562 (N_37562,N_36564,N_36441);
xor U37563 (N_37563,N_36780,N_36395);
xnor U37564 (N_37564,N_36885,N_36315);
and U37565 (N_37565,N_36401,N_36278);
and U37566 (N_37566,N_36807,N_36253);
xnor U37567 (N_37567,N_36406,N_36991);
and U37568 (N_37568,N_36971,N_36377);
or U37569 (N_37569,N_36241,N_36873);
and U37570 (N_37570,N_36337,N_36049);
xnor U37571 (N_37571,N_36171,N_36161);
nand U37572 (N_37572,N_36980,N_36004);
nand U37573 (N_37573,N_36261,N_36944);
nor U37574 (N_37574,N_36311,N_36355);
or U37575 (N_37575,N_36487,N_36970);
nand U37576 (N_37576,N_36495,N_36839);
xnor U37577 (N_37577,N_36808,N_36585);
xnor U37578 (N_37578,N_36571,N_36501);
or U37579 (N_37579,N_36873,N_36331);
and U37580 (N_37580,N_36805,N_36893);
or U37581 (N_37581,N_36263,N_36850);
nor U37582 (N_37582,N_36200,N_36426);
and U37583 (N_37583,N_36284,N_36406);
or U37584 (N_37584,N_36226,N_36956);
nand U37585 (N_37585,N_36640,N_36212);
and U37586 (N_37586,N_36247,N_36205);
and U37587 (N_37587,N_36318,N_36726);
and U37588 (N_37588,N_36151,N_36449);
xor U37589 (N_37589,N_36528,N_36036);
or U37590 (N_37590,N_36358,N_36391);
and U37591 (N_37591,N_36635,N_36971);
xor U37592 (N_37592,N_36587,N_36891);
and U37593 (N_37593,N_36276,N_36407);
and U37594 (N_37594,N_36440,N_36544);
and U37595 (N_37595,N_36142,N_36635);
nor U37596 (N_37596,N_36601,N_36127);
xnor U37597 (N_37597,N_36204,N_36682);
or U37598 (N_37598,N_36865,N_36171);
and U37599 (N_37599,N_36707,N_36898);
nand U37600 (N_37600,N_36318,N_36860);
and U37601 (N_37601,N_36319,N_36060);
nand U37602 (N_37602,N_36839,N_36477);
xnor U37603 (N_37603,N_36837,N_36215);
nor U37604 (N_37604,N_36062,N_36936);
and U37605 (N_37605,N_36607,N_36704);
or U37606 (N_37606,N_36027,N_36989);
nand U37607 (N_37607,N_36105,N_36729);
or U37608 (N_37608,N_36997,N_36168);
and U37609 (N_37609,N_36688,N_36760);
nor U37610 (N_37610,N_36917,N_36470);
xnor U37611 (N_37611,N_36385,N_36663);
or U37612 (N_37612,N_36920,N_36993);
or U37613 (N_37613,N_36276,N_36755);
xnor U37614 (N_37614,N_36766,N_36215);
and U37615 (N_37615,N_36385,N_36939);
nand U37616 (N_37616,N_36458,N_36189);
or U37617 (N_37617,N_36782,N_36991);
nor U37618 (N_37618,N_36900,N_36679);
nand U37619 (N_37619,N_36358,N_36225);
or U37620 (N_37620,N_36238,N_36319);
or U37621 (N_37621,N_36918,N_36065);
nand U37622 (N_37622,N_36544,N_36831);
and U37623 (N_37623,N_36676,N_36197);
or U37624 (N_37624,N_36556,N_36366);
or U37625 (N_37625,N_36554,N_36164);
and U37626 (N_37626,N_36367,N_36931);
or U37627 (N_37627,N_36158,N_36954);
xnor U37628 (N_37628,N_36566,N_36541);
or U37629 (N_37629,N_36893,N_36003);
or U37630 (N_37630,N_36619,N_36207);
nand U37631 (N_37631,N_36031,N_36158);
xor U37632 (N_37632,N_36049,N_36547);
or U37633 (N_37633,N_36609,N_36953);
and U37634 (N_37634,N_36488,N_36542);
nand U37635 (N_37635,N_36875,N_36620);
nor U37636 (N_37636,N_36273,N_36312);
and U37637 (N_37637,N_36757,N_36859);
xnor U37638 (N_37638,N_36438,N_36650);
nand U37639 (N_37639,N_36933,N_36119);
xnor U37640 (N_37640,N_36265,N_36761);
nor U37641 (N_37641,N_36199,N_36355);
nor U37642 (N_37642,N_36744,N_36889);
or U37643 (N_37643,N_36898,N_36367);
xnor U37644 (N_37644,N_36979,N_36484);
xor U37645 (N_37645,N_36931,N_36866);
or U37646 (N_37646,N_36104,N_36920);
nand U37647 (N_37647,N_36637,N_36195);
and U37648 (N_37648,N_36085,N_36813);
nand U37649 (N_37649,N_36668,N_36855);
and U37650 (N_37650,N_36646,N_36229);
and U37651 (N_37651,N_36810,N_36354);
or U37652 (N_37652,N_36542,N_36082);
and U37653 (N_37653,N_36068,N_36763);
or U37654 (N_37654,N_36856,N_36145);
or U37655 (N_37655,N_36896,N_36030);
and U37656 (N_37656,N_36463,N_36826);
nand U37657 (N_37657,N_36618,N_36282);
or U37658 (N_37658,N_36913,N_36529);
nor U37659 (N_37659,N_36793,N_36768);
or U37660 (N_37660,N_36010,N_36701);
and U37661 (N_37661,N_36393,N_36649);
nand U37662 (N_37662,N_36900,N_36139);
or U37663 (N_37663,N_36028,N_36246);
and U37664 (N_37664,N_36175,N_36257);
nor U37665 (N_37665,N_36450,N_36313);
nand U37666 (N_37666,N_36744,N_36595);
nor U37667 (N_37667,N_36089,N_36159);
or U37668 (N_37668,N_36804,N_36382);
or U37669 (N_37669,N_36756,N_36789);
or U37670 (N_37670,N_36614,N_36183);
or U37671 (N_37671,N_36006,N_36400);
nor U37672 (N_37672,N_36552,N_36768);
nor U37673 (N_37673,N_36962,N_36732);
or U37674 (N_37674,N_36318,N_36765);
xnor U37675 (N_37675,N_36962,N_36920);
and U37676 (N_37676,N_36001,N_36859);
and U37677 (N_37677,N_36740,N_36025);
xor U37678 (N_37678,N_36411,N_36827);
or U37679 (N_37679,N_36921,N_36058);
and U37680 (N_37680,N_36820,N_36889);
nand U37681 (N_37681,N_36753,N_36342);
nand U37682 (N_37682,N_36918,N_36715);
or U37683 (N_37683,N_36932,N_36038);
or U37684 (N_37684,N_36255,N_36013);
nor U37685 (N_37685,N_36625,N_36573);
or U37686 (N_37686,N_36870,N_36604);
or U37687 (N_37687,N_36164,N_36950);
nor U37688 (N_37688,N_36060,N_36401);
nor U37689 (N_37689,N_36070,N_36209);
and U37690 (N_37690,N_36868,N_36356);
xor U37691 (N_37691,N_36634,N_36015);
xnor U37692 (N_37692,N_36967,N_36229);
nand U37693 (N_37693,N_36531,N_36091);
nand U37694 (N_37694,N_36939,N_36240);
nand U37695 (N_37695,N_36387,N_36385);
or U37696 (N_37696,N_36060,N_36763);
or U37697 (N_37697,N_36275,N_36002);
xnor U37698 (N_37698,N_36431,N_36123);
and U37699 (N_37699,N_36660,N_36555);
xnor U37700 (N_37700,N_36273,N_36724);
nor U37701 (N_37701,N_36462,N_36134);
or U37702 (N_37702,N_36960,N_36660);
xor U37703 (N_37703,N_36481,N_36283);
nand U37704 (N_37704,N_36051,N_36284);
nor U37705 (N_37705,N_36589,N_36416);
nand U37706 (N_37706,N_36679,N_36665);
xnor U37707 (N_37707,N_36040,N_36675);
xnor U37708 (N_37708,N_36131,N_36489);
or U37709 (N_37709,N_36336,N_36441);
xor U37710 (N_37710,N_36492,N_36348);
nand U37711 (N_37711,N_36469,N_36579);
nand U37712 (N_37712,N_36818,N_36463);
nor U37713 (N_37713,N_36822,N_36068);
nor U37714 (N_37714,N_36970,N_36079);
nand U37715 (N_37715,N_36629,N_36126);
xor U37716 (N_37716,N_36802,N_36729);
or U37717 (N_37717,N_36711,N_36964);
xor U37718 (N_37718,N_36588,N_36548);
or U37719 (N_37719,N_36557,N_36799);
nand U37720 (N_37720,N_36397,N_36778);
and U37721 (N_37721,N_36536,N_36569);
nand U37722 (N_37722,N_36611,N_36105);
nor U37723 (N_37723,N_36457,N_36362);
nand U37724 (N_37724,N_36385,N_36274);
and U37725 (N_37725,N_36625,N_36245);
xnor U37726 (N_37726,N_36771,N_36853);
xnor U37727 (N_37727,N_36191,N_36881);
xnor U37728 (N_37728,N_36221,N_36883);
nor U37729 (N_37729,N_36707,N_36749);
nor U37730 (N_37730,N_36448,N_36224);
or U37731 (N_37731,N_36316,N_36822);
and U37732 (N_37732,N_36018,N_36456);
or U37733 (N_37733,N_36115,N_36626);
nand U37734 (N_37734,N_36919,N_36752);
nor U37735 (N_37735,N_36513,N_36125);
nor U37736 (N_37736,N_36322,N_36811);
and U37737 (N_37737,N_36487,N_36509);
nand U37738 (N_37738,N_36461,N_36458);
or U37739 (N_37739,N_36736,N_36531);
nand U37740 (N_37740,N_36643,N_36297);
nand U37741 (N_37741,N_36784,N_36583);
nand U37742 (N_37742,N_36152,N_36177);
and U37743 (N_37743,N_36667,N_36768);
or U37744 (N_37744,N_36964,N_36362);
and U37745 (N_37745,N_36215,N_36442);
xor U37746 (N_37746,N_36058,N_36266);
and U37747 (N_37747,N_36219,N_36494);
xnor U37748 (N_37748,N_36843,N_36333);
nor U37749 (N_37749,N_36603,N_36550);
or U37750 (N_37750,N_36842,N_36925);
xor U37751 (N_37751,N_36006,N_36296);
nor U37752 (N_37752,N_36685,N_36251);
and U37753 (N_37753,N_36208,N_36818);
and U37754 (N_37754,N_36336,N_36797);
and U37755 (N_37755,N_36373,N_36011);
xnor U37756 (N_37756,N_36150,N_36226);
xor U37757 (N_37757,N_36273,N_36450);
nor U37758 (N_37758,N_36109,N_36200);
nor U37759 (N_37759,N_36126,N_36204);
and U37760 (N_37760,N_36627,N_36680);
and U37761 (N_37761,N_36336,N_36315);
nor U37762 (N_37762,N_36641,N_36760);
nand U37763 (N_37763,N_36341,N_36036);
nor U37764 (N_37764,N_36373,N_36255);
and U37765 (N_37765,N_36440,N_36656);
nand U37766 (N_37766,N_36519,N_36723);
nor U37767 (N_37767,N_36596,N_36123);
nand U37768 (N_37768,N_36696,N_36523);
nor U37769 (N_37769,N_36614,N_36818);
xor U37770 (N_37770,N_36339,N_36085);
or U37771 (N_37771,N_36733,N_36582);
or U37772 (N_37772,N_36227,N_36146);
xor U37773 (N_37773,N_36766,N_36451);
or U37774 (N_37774,N_36343,N_36095);
or U37775 (N_37775,N_36490,N_36701);
or U37776 (N_37776,N_36795,N_36067);
xnor U37777 (N_37777,N_36674,N_36951);
nor U37778 (N_37778,N_36486,N_36557);
or U37779 (N_37779,N_36445,N_36315);
or U37780 (N_37780,N_36305,N_36454);
and U37781 (N_37781,N_36069,N_36379);
or U37782 (N_37782,N_36570,N_36181);
nand U37783 (N_37783,N_36964,N_36838);
nand U37784 (N_37784,N_36181,N_36806);
nor U37785 (N_37785,N_36591,N_36664);
xnor U37786 (N_37786,N_36421,N_36877);
nor U37787 (N_37787,N_36714,N_36943);
and U37788 (N_37788,N_36862,N_36504);
xnor U37789 (N_37789,N_36333,N_36650);
nor U37790 (N_37790,N_36109,N_36313);
xnor U37791 (N_37791,N_36860,N_36965);
nand U37792 (N_37792,N_36960,N_36000);
nor U37793 (N_37793,N_36421,N_36370);
and U37794 (N_37794,N_36936,N_36505);
xnor U37795 (N_37795,N_36029,N_36982);
nor U37796 (N_37796,N_36793,N_36537);
xor U37797 (N_37797,N_36414,N_36522);
or U37798 (N_37798,N_36320,N_36502);
xor U37799 (N_37799,N_36103,N_36013);
nand U37800 (N_37800,N_36518,N_36047);
or U37801 (N_37801,N_36636,N_36654);
nor U37802 (N_37802,N_36459,N_36037);
nand U37803 (N_37803,N_36242,N_36705);
nor U37804 (N_37804,N_36009,N_36441);
or U37805 (N_37805,N_36255,N_36154);
or U37806 (N_37806,N_36651,N_36075);
xnor U37807 (N_37807,N_36196,N_36581);
nor U37808 (N_37808,N_36288,N_36123);
nor U37809 (N_37809,N_36615,N_36961);
nor U37810 (N_37810,N_36303,N_36264);
xnor U37811 (N_37811,N_36177,N_36864);
nor U37812 (N_37812,N_36030,N_36420);
and U37813 (N_37813,N_36894,N_36438);
or U37814 (N_37814,N_36448,N_36796);
nor U37815 (N_37815,N_36515,N_36607);
nor U37816 (N_37816,N_36612,N_36386);
xor U37817 (N_37817,N_36856,N_36306);
nor U37818 (N_37818,N_36886,N_36173);
or U37819 (N_37819,N_36037,N_36959);
nor U37820 (N_37820,N_36683,N_36660);
or U37821 (N_37821,N_36123,N_36675);
and U37822 (N_37822,N_36124,N_36390);
nand U37823 (N_37823,N_36709,N_36358);
and U37824 (N_37824,N_36725,N_36059);
nand U37825 (N_37825,N_36356,N_36977);
or U37826 (N_37826,N_36601,N_36062);
nand U37827 (N_37827,N_36765,N_36749);
nand U37828 (N_37828,N_36013,N_36414);
nand U37829 (N_37829,N_36936,N_36707);
or U37830 (N_37830,N_36022,N_36332);
nand U37831 (N_37831,N_36012,N_36300);
nor U37832 (N_37832,N_36346,N_36178);
xor U37833 (N_37833,N_36378,N_36867);
or U37834 (N_37834,N_36366,N_36323);
and U37835 (N_37835,N_36329,N_36826);
nor U37836 (N_37836,N_36681,N_36244);
nand U37837 (N_37837,N_36747,N_36820);
xnor U37838 (N_37838,N_36253,N_36630);
or U37839 (N_37839,N_36451,N_36419);
nor U37840 (N_37840,N_36792,N_36429);
or U37841 (N_37841,N_36057,N_36964);
nand U37842 (N_37842,N_36840,N_36904);
nor U37843 (N_37843,N_36347,N_36280);
or U37844 (N_37844,N_36787,N_36152);
nand U37845 (N_37845,N_36490,N_36655);
or U37846 (N_37846,N_36046,N_36405);
nor U37847 (N_37847,N_36438,N_36312);
nor U37848 (N_37848,N_36760,N_36568);
xnor U37849 (N_37849,N_36142,N_36488);
and U37850 (N_37850,N_36742,N_36260);
xor U37851 (N_37851,N_36439,N_36250);
nand U37852 (N_37852,N_36393,N_36924);
xor U37853 (N_37853,N_36204,N_36640);
or U37854 (N_37854,N_36163,N_36190);
xor U37855 (N_37855,N_36465,N_36761);
or U37856 (N_37856,N_36793,N_36986);
and U37857 (N_37857,N_36726,N_36214);
and U37858 (N_37858,N_36652,N_36410);
or U37859 (N_37859,N_36409,N_36248);
or U37860 (N_37860,N_36042,N_36492);
and U37861 (N_37861,N_36287,N_36600);
or U37862 (N_37862,N_36060,N_36919);
or U37863 (N_37863,N_36355,N_36071);
xnor U37864 (N_37864,N_36568,N_36630);
nor U37865 (N_37865,N_36867,N_36968);
or U37866 (N_37866,N_36055,N_36951);
xnor U37867 (N_37867,N_36050,N_36565);
and U37868 (N_37868,N_36914,N_36704);
nor U37869 (N_37869,N_36105,N_36542);
xnor U37870 (N_37870,N_36545,N_36306);
xor U37871 (N_37871,N_36722,N_36678);
and U37872 (N_37872,N_36625,N_36609);
nand U37873 (N_37873,N_36404,N_36358);
nand U37874 (N_37874,N_36665,N_36197);
xnor U37875 (N_37875,N_36240,N_36966);
or U37876 (N_37876,N_36576,N_36780);
xor U37877 (N_37877,N_36188,N_36205);
nand U37878 (N_37878,N_36868,N_36622);
and U37879 (N_37879,N_36578,N_36844);
xor U37880 (N_37880,N_36603,N_36485);
nor U37881 (N_37881,N_36848,N_36768);
nand U37882 (N_37882,N_36357,N_36949);
nand U37883 (N_37883,N_36059,N_36602);
and U37884 (N_37884,N_36550,N_36363);
nand U37885 (N_37885,N_36347,N_36573);
xnor U37886 (N_37886,N_36902,N_36708);
and U37887 (N_37887,N_36193,N_36716);
xor U37888 (N_37888,N_36546,N_36858);
or U37889 (N_37889,N_36334,N_36557);
xnor U37890 (N_37890,N_36853,N_36078);
nor U37891 (N_37891,N_36033,N_36284);
nand U37892 (N_37892,N_36556,N_36860);
nand U37893 (N_37893,N_36591,N_36201);
xor U37894 (N_37894,N_36701,N_36522);
and U37895 (N_37895,N_36533,N_36058);
nor U37896 (N_37896,N_36333,N_36627);
and U37897 (N_37897,N_36839,N_36440);
nand U37898 (N_37898,N_36259,N_36962);
and U37899 (N_37899,N_36891,N_36032);
or U37900 (N_37900,N_36815,N_36963);
nand U37901 (N_37901,N_36885,N_36124);
and U37902 (N_37902,N_36587,N_36468);
nand U37903 (N_37903,N_36324,N_36907);
or U37904 (N_37904,N_36596,N_36239);
or U37905 (N_37905,N_36344,N_36847);
or U37906 (N_37906,N_36989,N_36076);
nor U37907 (N_37907,N_36289,N_36988);
nand U37908 (N_37908,N_36229,N_36215);
nor U37909 (N_37909,N_36772,N_36098);
xnor U37910 (N_37910,N_36142,N_36293);
xor U37911 (N_37911,N_36105,N_36374);
and U37912 (N_37912,N_36484,N_36527);
or U37913 (N_37913,N_36231,N_36479);
and U37914 (N_37914,N_36489,N_36727);
xor U37915 (N_37915,N_36344,N_36400);
or U37916 (N_37916,N_36270,N_36124);
xnor U37917 (N_37917,N_36909,N_36071);
or U37918 (N_37918,N_36492,N_36186);
nor U37919 (N_37919,N_36614,N_36764);
nor U37920 (N_37920,N_36107,N_36613);
and U37921 (N_37921,N_36782,N_36362);
nand U37922 (N_37922,N_36135,N_36443);
or U37923 (N_37923,N_36111,N_36622);
and U37924 (N_37924,N_36756,N_36233);
nand U37925 (N_37925,N_36637,N_36470);
nor U37926 (N_37926,N_36020,N_36312);
nor U37927 (N_37927,N_36870,N_36430);
nor U37928 (N_37928,N_36890,N_36876);
nor U37929 (N_37929,N_36819,N_36292);
or U37930 (N_37930,N_36887,N_36159);
nor U37931 (N_37931,N_36374,N_36843);
xor U37932 (N_37932,N_36172,N_36936);
and U37933 (N_37933,N_36575,N_36563);
nor U37934 (N_37934,N_36059,N_36511);
nand U37935 (N_37935,N_36171,N_36902);
and U37936 (N_37936,N_36019,N_36965);
nand U37937 (N_37937,N_36151,N_36506);
nand U37938 (N_37938,N_36436,N_36902);
nor U37939 (N_37939,N_36485,N_36149);
and U37940 (N_37940,N_36059,N_36390);
xor U37941 (N_37941,N_36587,N_36386);
or U37942 (N_37942,N_36864,N_36101);
xnor U37943 (N_37943,N_36301,N_36551);
xnor U37944 (N_37944,N_36275,N_36421);
or U37945 (N_37945,N_36858,N_36280);
nor U37946 (N_37946,N_36615,N_36306);
or U37947 (N_37947,N_36974,N_36720);
xnor U37948 (N_37948,N_36760,N_36299);
nor U37949 (N_37949,N_36898,N_36420);
and U37950 (N_37950,N_36979,N_36513);
xnor U37951 (N_37951,N_36406,N_36618);
nand U37952 (N_37952,N_36822,N_36662);
or U37953 (N_37953,N_36570,N_36310);
nor U37954 (N_37954,N_36462,N_36590);
or U37955 (N_37955,N_36801,N_36130);
nand U37956 (N_37956,N_36569,N_36162);
or U37957 (N_37957,N_36877,N_36551);
or U37958 (N_37958,N_36151,N_36071);
and U37959 (N_37959,N_36407,N_36675);
xnor U37960 (N_37960,N_36195,N_36152);
xor U37961 (N_37961,N_36170,N_36809);
xor U37962 (N_37962,N_36513,N_36790);
nor U37963 (N_37963,N_36939,N_36567);
nor U37964 (N_37964,N_36324,N_36385);
nor U37965 (N_37965,N_36014,N_36919);
or U37966 (N_37966,N_36445,N_36092);
nor U37967 (N_37967,N_36247,N_36937);
nand U37968 (N_37968,N_36895,N_36955);
and U37969 (N_37969,N_36052,N_36059);
and U37970 (N_37970,N_36274,N_36888);
nor U37971 (N_37971,N_36264,N_36008);
or U37972 (N_37972,N_36411,N_36960);
and U37973 (N_37973,N_36289,N_36966);
nor U37974 (N_37974,N_36646,N_36603);
nand U37975 (N_37975,N_36761,N_36426);
xor U37976 (N_37976,N_36832,N_36332);
or U37977 (N_37977,N_36634,N_36613);
nand U37978 (N_37978,N_36087,N_36064);
nor U37979 (N_37979,N_36199,N_36449);
nor U37980 (N_37980,N_36201,N_36837);
or U37981 (N_37981,N_36180,N_36923);
nor U37982 (N_37982,N_36376,N_36193);
or U37983 (N_37983,N_36342,N_36029);
or U37984 (N_37984,N_36315,N_36378);
nor U37985 (N_37985,N_36737,N_36243);
and U37986 (N_37986,N_36213,N_36712);
xor U37987 (N_37987,N_36157,N_36521);
nand U37988 (N_37988,N_36222,N_36769);
nor U37989 (N_37989,N_36766,N_36020);
and U37990 (N_37990,N_36675,N_36296);
nand U37991 (N_37991,N_36905,N_36713);
and U37992 (N_37992,N_36134,N_36668);
and U37993 (N_37993,N_36325,N_36584);
xor U37994 (N_37994,N_36181,N_36659);
nand U37995 (N_37995,N_36173,N_36607);
nand U37996 (N_37996,N_36094,N_36158);
and U37997 (N_37997,N_36195,N_36578);
or U37998 (N_37998,N_36816,N_36259);
xnor U37999 (N_37999,N_36327,N_36649);
xnor U38000 (N_38000,N_37538,N_37055);
or U38001 (N_38001,N_37799,N_37548);
and U38002 (N_38002,N_37401,N_37661);
xor U38003 (N_38003,N_37985,N_37839);
xnor U38004 (N_38004,N_37859,N_37279);
and U38005 (N_38005,N_37696,N_37339);
or U38006 (N_38006,N_37184,N_37711);
xnor U38007 (N_38007,N_37207,N_37603);
or U38008 (N_38008,N_37892,N_37775);
or U38009 (N_38009,N_37131,N_37011);
or U38010 (N_38010,N_37641,N_37836);
nand U38011 (N_38011,N_37426,N_37257);
nor U38012 (N_38012,N_37460,N_37769);
nor U38013 (N_38013,N_37183,N_37567);
or U38014 (N_38014,N_37116,N_37719);
nor U38015 (N_38015,N_37613,N_37221);
nor U38016 (N_38016,N_37351,N_37561);
nand U38017 (N_38017,N_37518,N_37447);
nor U38018 (N_38018,N_37380,N_37188);
and U38019 (N_38019,N_37552,N_37192);
nand U38020 (N_38020,N_37699,N_37141);
nand U38021 (N_38021,N_37424,N_37559);
xor U38022 (N_38022,N_37582,N_37675);
nand U38023 (N_38023,N_37085,N_37557);
or U38024 (N_38024,N_37509,N_37466);
nor U38025 (N_38025,N_37077,N_37313);
or U38026 (N_38026,N_37956,N_37366);
nand U38027 (N_38027,N_37653,N_37076);
nand U38028 (N_38028,N_37996,N_37064);
or U38029 (N_38029,N_37473,N_37340);
and U38030 (N_38030,N_37525,N_37484);
xor U38031 (N_38031,N_37623,N_37949);
xor U38032 (N_38032,N_37234,N_37970);
or U38033 (N_38033,N_37274,N_37140);
xnor U38034 (N_38034,N_37530,N_37852);
and U38035 (N_38035,N_37453,N_37843);
nand U38036 (N_38036,N_37199,N_37702);
nand U38037 (N_38037,N_37521,N_37701);
xor U38038 (N_38038,N_37007,N_37413);
or U38039 (N_38039,N_37408,N_37478);
or U38040 (N_38040,N_37019,N_37901);
xnor U38041 (N_38041,N_37244,N_37186);
and U38042 (N_38042,N_37658,N_37531);
or U38043 (N_38043,N_37025,N_37747);
xnor U38044 (N_38044,N_37382,N_37179);
xnor U38045 (N_38045,N_37500,N_37662);
nand U38046 (N_38046,N_37685,N_37938);
nor U38047 (N_38047,N_37941,N_37931);
xnor U38048 (N_38048,N_37158,N_37648);
nand U38049 (N_38049,N_37590,N_37533);
xor U38050 (N_38050,N_37565,N_37487);
nor U38051 (N_38051,N_37580,N_37194);
and U38052 (N_38052,N_37456,N_37438);
xnor U38053 (N_38053,N_37224,N_37047);
and U38054 (N_38054,N_37588,N_37520);
or U38055 (N_38055,N_37905,N_37877);
nand U38056 (N_38056,N_37316,N_37104);
nor U38057 (N_38057,N_37650,N_37618);
nand U38058 (N_38058,N_37228,N_37512);
or U38059 (N_38059,N_37440,N_37082);
and U38060 (N_38060,N_37793,N_37361);
xnor U38061 (N_38061,N_37247,N_37123);
nor U38062 (N_38062,N_37665,N_37300);
and U38063 (N_38063,N_37527,N_37948);
or U38064 (N_38064,N_37091,N_37803);
xnor U38065 (N_38065,N_37833,N_37563);
nand U38066 (N_38066,N_37503,N_37804);
nor U38067 (N_38067,N_37286,N_37871);
xor U38068 (N_38068,N_37133,N_37819);
nor U38069 (N_38069,N_37881,N_37318);
nand U38070 (N_38070,N_37823,N_37489);
xnor U38071 (N_38071,N_37687,N_37258);
xor U38072 (N_38072,N_37939,N_37672);
nor U38073 (N_38073,N_37443,N_37093);
nand U38074 (N_38074,N_37848,N_37309);
and U38075 (N_38075,N_37607,N_37004);
nand U38076 (N_38076,N_37295,N_37343);
nand U38077 (N_38077,N_37846,N_37034);
xnor U38078 (N_38078,N_37777,N_37075);
xnor U38079 (N_38079,N_37005,N_37491);
and U38080 (N_38080,N_37227,N_37389);
or U38081 (N_38081,N_37157,N_37037);
and U38082 (N_38082,N_37673,N_37828);
xor U38083 (N_38083,N_37425,N_37288);
and U38084 (N_38084,N_37337,N_37811);
nor U38085 (N_38085,N_37358,N_37649);
nand U38086 (N_38086,N_37807,N_37414);
nand U38087 (N_38087,N_37462,N_37853);
nand U38088 (N_38088,N_37904,N_37180);
nand U38089 (N_38089,N_37142,N_37721);
and U38090 (N_38090,N_37051,N_37950);
nand U38091 (N_38091,N_37237,N_37962);
and U38092 (N_38092,N_37558,N_37910);
nor U38093 (N_38093,N_37212,N_37148);
nor U38094 (N_38094,N_37292,N_37139);
nand U38095 (N_38095,N_37677,N_37523);
nor U38096 (N_38096,N_37454,N_37597);
nand U38097 (N_38097,N_37394,N_37378);
and U38098 (N_38098,N_37448,N_37411);
or U38099 (N_38099,N_37726,N_37089);
nand U38100 (N_38100,N_37418,N_37544);
nor U38101 (N_38101,N_37385,N_37165);
nand U38102 (N_38102,N_37050,N_37020);
xor U38103 (N_38103,N_37119,N_37009);
and U38104 (N_38104,N_37336,N_37112);
nand U38105 (N_38105,N_37253,N_37357);
nor U38106 (N_38106,N_37018,N_37345);
nor U38107 (N_38107,N_37554,N_37164);
xnor U38108 (N_38108,N_37707,N_37344);
and U38109 (N_38109,N_37121,N_37074);
nand U38110 (N_38110,N_37543,N_37774);
nor U38111 (N_38111,N_37392,N_37102);
or U38112 (N_38112,N_37922,N_37980);
nor U38113 (N_38113,N_37639,N_37039);
nand U38114 (N_38114,N_37746,N_37880);
and U38115 (N_38115,N_37486,N_37753);
or U38116 (N_38116,N_37961,N_37697);
or U38117 (N_38117,N_37878,N_37727);
nand U38118 (N_38118,N_37783,N_37206);
or U38119 (N_38119,N_37973,N_37428);
or U38120 (N_38120,N_37920,N_37876);
or U38121 (N_38121,N_37480,N_37749);
xor U38122 (N_38122,N_37252,N_37373);
nand U38123 (N_38123,N_37259,N_37153);
or U38124 (N_38124,N_37238,N_37107);
nor U38125 (N_38125,N_37912,N_37269);
or U38126 (N_38126,N_37126,N_37755);
nand U38127 (N_38127,N_37383,N_37045);
or U38128 (N_38128,N_37936,N_37763);
xnor U38129 (N_38129,N_37888,N_37611);
xnor U38130 (N_38130,N_37223,N_37120);
nor U38131 (N_38131,N_37869,N_37000);
or U38132 (N_38132,N_37481,N_37850);
or U38133 (N_38133,N_37229,N_37315);
and U38134 (N_38134,N_37797,N_37322);
nand U38135 (N_38135,N_37609,N_37870);
and U38136 (N_38136,N_37855,N_37713);
xnor U38137 (N_38137,N_37765,N_37187);
nand U38138 (N_38138,N_37268,N_37568);
nand U38139 (N_38139,N_37222,N_37532);
or U38140 (N_38140,N_37935,N_37502);
and U38141 (N_38141,N_37759,N_37863);
or U38142 (N_38142,N_37628,N_37715);
or U38143 (N_38143,N_37474,N_37993);
nand U38144 (N_38144,N_37205,N_37255);
xnor U38145 (N_38145,N_37813,N_37978);
xnor U38146 (N_38146,N_37325,N_37267);
and U38147 (N_38147,N_37780,N_37737);
nand U38148 (N_38148,N_37926,N_37808);
nand U38149 (N_38149,N_37692,N_37147);
xor U38150 (N_38150,N_37306,N_37958);
or U38151 (N_38151,N_37354,N_37844);
nor U38152 (N_38152,N_37412,N_37356);
nor U38153 (N_38153,N_37537,N_37113);
xnor U38154 (N_38154,N_37465,N_37856);
xnor U38155 (N_38155,N_37493,N_37396);
nand U38156 (N_38156,N_37998,N_37136);
nand U38157 (N_38157,N_37895,N_37505);
nor U38158 (N_38158,N_37917,N_37647);
nor U38159 (N_38159,N_37211,N_37435);
and U38160 (N_38160,N_37553,N_37096);
nor U38161 (N_38161,N_37353,N_37163);
or U38162 (N_38162,N_37111,N_37053);
and U38163 (N_38163,N_37442,N_37738);
nor U38164 (N_38164,N_37766,N_37627);
nand U38165 (N_38165,N_37457,N_37049);
nor U38166 (N_38166,N_37417,N_37029);
nor U38167 (N_38167,N_37214,N_37256);
nor U38168 (N_38168,N_37193,N_37964);
nor U38169 (N_38169,N_37884,N_37115);
xnor U38170 (N_38170,N_37872,N_37646);
or U38171 (N_38171,N_37798,N_37556);
or U38172 (N_38172,N_37346,N_37273);
or U38173 (N_38173,N_37535,N_37511);
nor U38174 (N_38174,N_37965,N_37861);
nand U38175 (N_38175,N_37695,N_37177);
nor U38176 (N_38176,N_37534,N_37812);
nand U38177 (N_38177,N_37591,N_37002);
xor U38178 (N_38178,N_37945,N_37232);
nand U38179 (N_38179,N_37874,N_37235);
nor U38180 (N_38180,N_37916,N_37144);
nand U38181 (N_38181,N_37156,N_37249);
and U38182 (N_38182,N_37513,N_37372);
and U38183 (N_38183,N_37562,N_37573);
nand U38184 (N_38184,N_37399,N_37427);
nand U38185 (N_38185,N_37515,N_37990);
xor U38186 (N_38186,N_37040,N_37752);
or U38187 (N_38187,N_37445,N_37303);
nand U38188 (N_38188,N_37831,N_37065);
nor U38189 (N_38189,N_37925,N_37734);
or U38190 (N_38190,N_37150,N_37429);
xor U38191 (N_38191,N_37643,N_37976);
nand U38192 (N_38192,N_37175,N_37494);
nand U38193 (N_38193,N_37678,N_37555);
xor U38194 (N_38194,N_37003,N_37791);
xnor U38195 (N_38195,N_37407,N_37772);
xnor U38196 (N_38196,N_37826,N_37578);
nor U38197 (N_38197,N_37934,N_37094);
and U38198 (N_38198,N_37127,N_37472);
nand U38199 (N_38199,N_37806,N_37265);
nor U38200 (N_38200,N_37446,N_37246);
xnor U38201 (N_38201,N_37391,N_37704);
nor U38202 (N_38202,N_37195,N_37744);
xor U38203 (N_38203,N_37860,N_37248);
or U38204 (N_38204,N_37196,N_37287);
nand U38205 (N_38205,N_37624,N_37317);
nand U38206 (N_38206,N_37682,N_37422);
xnor U38207 (N_38207,N_37071,N_37689);
nand U38208 (N_38208,N_37108,N_37785);
nand U38209 (N_38209,N_37197,N_37341);
nand U38210 (N_38210,N_37760,N_37078);
nand U38211 (N_38211,N_37619,N_37656);
nand U38212 (N_38212,N_37169,N_37906);
nor U38213 (N_38213,N_37593,N_37595);
xnor U38214 (N_38214,N_37444,N_37911);
nand U38215 (N_38215,N_37270,N_37644);
xor U38216 (N_38216,N_37514,N_37581);
or U38217 (N_38217,N_37092,N_37600);
xnor U38218 (N_38218,N_37751,N_37101);
nand U38219 (N_38219,N_37430,N_37740);
xnor U38220 (N_38220,N_37266,N_37893);
xnor U38221 (N_38221,N_37483,N_37988);
nand U38222 (N_38222,N_37868,N_37606);
or U38223 (N_38223,N_37103,N_37277);
and U38224 (N_38224,N_37659,N_37902);
nand U38225 (N_38225,N_37681,N_37733);
nand U38226 (N_38226,N_37016,N_37773);
or U38227 (N_38227,N_37290,N_37146);
nor U38228 (N_38228,N_37858,N_37564);
and U38229 (N_38229,N_37889,N_37132);
nand U38230 (N_38230,N_37084,N_37294);
or U38231 (N_38231,N_37940,N_37170);
nand U38232 (N_38232,N_37099,N_37308);
nor U38233 (N_38233,N_37347,N_37981);
and U38234 (N_38234,N_37621,N_37008);
nand U38235 (N_38235,N_37021,N_37652);
nand U38236 (N_38236,N_37517,N_37161);
and U38237 (N_38237,N_37134,N_37991);
and U38238 (N_38238,N_37128,N_37043);
and U38239 (N_38239,N_37023,N_37063);
nand U38240 (N_38240,N_37790,N_37959);
xnor U38241 (N_38241,N_37060,N_37510);
and U38242 (N_38242,N_37311,N_37296);
or U38243 (N_38243,N_37485,N_37952);
and U38244 (N_38244,N_37731,N_37540);
xor U38245 (N_38245,N_37592,N_37708);
xnor U38246 (N_38246,N_37706,N_37690);
nor U38247 (N_38247,N_37897,N_37006);
and U38248 (N_38248,N_37820,N_37894);
nor U38249 (N_38249,N_37464,N_37622);
nand U38250 (N_38250,N_37620,N_37499);
xor U38251 (N_38251,N_37371,N_37587);
nand U38252 (N_38252,N_37670,N_37913);
and U38253 (N_38253,N_37864,N_37814);
nand U38254 (N_38254,N_37730,N_37566);
or U38255 (N_38255,N_37374,N_37079);
nand U38256 (N_38256,N_37743,N_37421);
nand U38257 (N_38257,N_37468,N_37506);
nor U38258 (N_38258,N_37027,N_37929);
xor U38259 (N_38259,N_37986,N_37569);
xnor U38260 (N_38260,N_37403,N_37957);
and U38261 (N_38261,N_37320,N_37887);
and U38262 (N_38262,N_37219,N_37381);
nand U38263 (N_38263,N_37189,N_37038);
or U38264 (N_38264,N_37914,N_37987);
or U38265 (N_38265,N_37151,N_37182);
nand U38266 (N_38266,N_37469,N_37918);
nand U38267 (N_38267,N_37634,N_37997);
or U38268 (N_38268,N_37254,N_37405);
or U38269 (N_38269,N_37933,N_37654);
nor U38270 (N_38270,N_37028,N_37989);
nor U38271 (N_38271,N_37501,N_37233);
xor U38272 (N_38272,N_37285,N_37459);
or U38273 (N_38273,N_37278,N_37896);
or U38274 (N_38274,N_37334,N_37736);
or U38275 (N_38275,N_37398,N_37610);
nand U38276 (N_38276,N_37676,N_37393);
xnor U38277 (N_38277,N_37498,N_37795);
xor U38278 (N_38278,N_37898,N_37827);
nand U38279 (N_38279,N_37226,N_37824);
or U38280 (N_38280,N_37630,N_37200);
xor U38281 (N_38281,N_37969,N_37434);
xnor U38282 (N_38282,N_37671,N_37764);
nor U38283 (N_38283,N_37907,N_37845);
nor U38284 (N_38284,N_37415,N_37416);
xor U38285 (N_38285,N_37741,N_37208);
nand U38286 (N_38286,N_37041,N_37106);
nor U38287 (N_38287,N_37838,N_37655);
xnor U38288 (N_38288,N_37974,N_37576);
nand U38289 (N_38289,N_37349,N_37342);
nor U38290 (N_38290,N_37335,N_37130);
xor U38291 (N_38291,N_37667,N_37081);
and U38292 (N_38292,N_37362,N_37810);
nor U38293 (N_38293,N_37923,N_37014);
nor U38294 (N_38294,N_37504,N_37241);
and U38295 (N_38295,N_37299,N_37999);
xor U38296 (N_38296,N_37327,N_37080);
or U38297 (N_38297,N_37044,N_37100);
and U38298 (N_38298,N_37026,N_37022);
or U38299 (N_38299,N_37301,N_37449);
nand U38300 (N_38300,N_37482,N_37031);
nand U38301 (N_38301,N_37717,N_37612);
or U38302 (N_38302,N_37842,N_37384);
and U38303 (N_38303,N_37251,N_37062);
xnor U38304 (N_38304,N_37754,N_37761);
xnor U38305 (N_38305,N_37802,N_37585);
nor U38306 (N_38306,N_37930,N_37352);
nand U38307 (N_38307,N_37275,N_37614);
or U38308 (N_38308,N_37599,N_37225);
xnor U38309 (N_38309,N_37982,N_37046);
or U38310 (N_38310,N_37291,N_37605);
nor U38311 (N_38311,N_37718,N_37596);
or U38312 (N_38312,N_37475,N_37983);
nand U38313 (N_38313,N_37488,N_37323);
and U38314 (N_38314,N_37979,N_37883);
or U38315 (N_38315,N_37160,N_37589);
and U38316 (N_38316,N_37069,N_37572);
and U38317 (N_38317,N_37947,N_37851);
nand U38318 (N_38318,N_37546,N_37015);
nand U38319 (N_38319,N_37307,N_37172);
and U38320 (N_38320,N_37549,N_37326);
nor U38321 (N_38321,N_37789,N_37700);
or U38322 (N_38322,N_37668,N_37202);
nor U38323 (N_38323,N_37159,N_37243);
and U38324 (N_38324,N_37276,N_37209);
or U38325 (N_38325,N_37875,N_37397);
nor U38326 (N_38326,N_37272,N_37735);
nand U38327 (N_38327,N_37282,N_37732);
and U38328 (N_38328,N_37879,N_37890);
and U38329 (N_38329,N_37162,N_37057);
xor U38330 (N_38330,N_37679,N_37355);
nor U38331 (N_38331,N_37545,N_37536);
or U38332 (N_38332,N_37691,N_37458);
or U38333 (N_38333,N_37857,N_37310);
nor U38334 (N_38334,N_37402,N_37470);
nor U38335 (N_38335,N_37097,N_37400);
xor U38336 (N_38336,N_37350,N_37263);
nor U38337 (N_38337,N_37837,N_37835);
xnor U38338 (N_38338,N_37036,N_37056);
nor U38339 (N_38339,N_37068,N_37758);
and U38340 (N_38340,N_37284,N_37645);
nand U38341 (N_38341,N_37995,N_37762);
nor U38342 (N_38342,N_37867,N_37637);
and U38343 (N_38343,N_37756,N_37001);
nand U38344 (N_38344,N_37967,N_37786);
nand U38345 (N_38345,N_37866,N_37017);
nand U38346 (N_38346,N_37467,N_37862);
and U38347 (N_38347,N_37145,N_37370);
or U38348 (N_38348,N_37210,N_37579);
xor U38349 (N_38349,N_37377,N_37240);
nand U38350 (N_38350,N_37185,N_37348);
and U38351 (N_38351,N_37739,N_37954);
and U38352 (N_38352,N_37794,N_37865);
nor U38353 (N_38353,N_37124,N_37575);
nand U38354 (N_38354,N_37943,N_37250);
xnor U38355 (N_38355,N_37771,N_37830);
or U38356 (N_38356,N_37975,N_37432);
nor U38357 (N_38357,N_37683,N_37406);
xnor U38358 (N_38358,N_37010,N_37757);
or U38359 (N_38359,N_37386,N_37154);
nand U38360 (N_38360,N_37698,N_37924);
or U38361 (N_38361,N_37490,N_37138);
or U38362 (N_38362,N_37090,N_37834);
and U38363 (N_38363,N_37776,N_37477);
xor U38364 (N_38364,N_37946,N_37321);
xor U38365 (N_38365,N_37629,N_37242);
nor U38366 (N_38366,N_37067,N_37927);
nand U38367 (N_38367,N_37849,N_37059);
and U38368 (N_38368,N_37712,N_37479);
xor U38369 (N_38369,N_37423,N_37451);
nand U38370 (N_38370,N_37114,N_37095);
xor U38371 (N_38371,N_37178,N_37239);
xor U38372 (N_38372,N_37714,N_37439);
nand U38373 (N_38373,N_37441,N_37953);
nand U38374 (N_38374,N_37635,N_37168);
xor U38375 (N_38375,N_37135,N_37539);
nor U38376 (N_38376,N_37173,N_37261);
nand U38377 (N_38377,N_37686,N_37725);
xor U38378 (N_38378,N_37217,N_37507);
and U38379 (N_38379,N_37052,N_37304);
and U38380 (N_38380,N_37364,N_37604);
nand U38381 (N_38381,N_37742,N_37395);
and U38382 (N_38382,N_37433,N_37626);
xnor U38383 (N_38383,N_37297,N_37784);
nand U38384 (N_38384,N_37452,N_37289);
xnor U38385 (N_38385,N_37110,N_37387);
xor U38386 (N_38386,N_37745,N_37632);
nor U38387 (N_38387,N_37528,N_37633);
xor U38388 (N_38388,N_37616,N_37577);
nor U38389 (N_38389,N_37657,N_37463);
and U38390 (N_38390,N_37617,N_37365);
or U38391 (N_38391,N_37174,N_37710);
nor U38392 (N_38392,N_37782,N_37903);
and U38393 (N_38393,N_37171,N_37886);
and U38394 (N_38394,N_37942,N_37450);
xor U38395 (N_38395,N_37722,N_37822);
xor U38396 (N_38396,N_37293,N_37329);
nand U38397 (N_38397,N_37109,N_37368);
xor U38398 (N_38398,N_37680,N_37314);
nor U38399 (N_38399,N_37013,N_37571);
xnor U38400 (N_38400,N_37963,N_37181);
nand U38401 (N_38401,N_37496,N_37709);
or U38402 (N_38402,N_37035,N_37821);
nand U38403 (N_38403,N_37972,N_37608);
nor U38404 (N_38404,N_37420,N_37792);
nand U38405 (N_38405,N_37817,N_37215);
xor U38406 (N_38406,N_37167,N_37779);
and U38407 (N_38407,N_37332,N_37281);
or U38408 (N_38408,N_37770,N_37213);
nor U38409 (N_38409,N_37176,N_37885);
nor U38410 (N_38410,N_37663,N_37873);
or U38411 (N_38411,N_37636,N_37330);
or U38412 (N_38412,N_37117,N_37932);
nand U38413 (N_38413,N_37305,N_37058);
xnor U38414 (N_38414,N_37149,N_37264);
or U38415 (N_38415,N_37919,N_37431);
nand U38416 (N_38416,N_37818,N_37550);
or U38417 (N_38417,N_37570,N_37542);
and U38418 (N_38418,N_37705,N_37367);
nor U38419 (N_38419,N_37640,N_37541);
nand U38420 (N_38420,N_37809,N_37966);
nor U38421 (N_38421,N_37497,N_37781);
nor U38422 (N_38422,N_37921,N_37841);
xor U38423 (N_38423,N_37066,N_37230);
nor U38424 (N_38424,N_37220,N_37012);
nand U38425 (N_38425,N_37360,N_37992);
and U38426 (N_38426,N_37476,N_37083);
nor U38427 (N_38427,N_37048,N_37033);
nor U38428 (N_38428,N_37198,N_37376);
or U38429 (N_38429,N_37522,N_37087);
nand U38430 (N_38430,N_37271,N_37319);
nor U38431 (N_38431,N_37908,N_37098);
and U38432 (N_38432,N_37832,N_37201);
xnor U38433 (N_38433,N_37615,N_37436);
nand U38434 (N_38434,N_37660,N_37602);
and U38435 (N_38435,N_37125,N_37369);
or U38436 (N_38436,N_37994,N_37388);
nor U38437 (N_38437,N_37152,N_37086);
nand U38438 (N_38438,N_37105,N_37236);
nand U38439 (N_38439,N_37669,N_37166);
xnor U38440 (N_38440,N_37410,N_37216);
and U38441 (N_38441,N_37333,N_37815);
nor U38442 (N_38442,N_37495,N_37338);
nor U38443 (N_38443,N_37245,N_37122);
nand U38444 (N_38444,N_37716,N_37519);
or U38445 (N_38445,N_37840,N_37703);
xnor U38446 (N_38446,N_37203,N_37379);
nand U38447 (N_38447,N_37955,N_37638);
or U38448 (N_38448,N_37787,N_37801);
nand U38449 (N_38449,N_37891,N_37129);
or U38450 (N_38450,N_37684,N_37526);
nor U38451 (N_38451,N_37260,N_37800);
and U38452 (N_38452,N_37231,N_37032);
xor U38453 (N_38453,N_37547,N_37190);
nand U38454 (N_38454,N_37461,N_37944);
or U38455 (N_38455,N_37601,N_37724);
or U38456 (N_38456,N_37899,N_37328);
nand U38457 (N_38457,N_37359,N_37584);
and U38458 (N_38458,N_37298,N_37977);
and U38459 (N_38459,N_37796,N_37586);
xnor U38460 (N_38460,N_37788,N_37778);
or U38461 (N_38461,N_37723,N_37302);
xnor U38462 (N_38462,N_37805,N_37375);
nor U38463 (N_38463,N_37631,N_37331);
or U38464 (N_38464,N_37960,N_37583);
nor U38465 (N_38465,N_37390,N_37455);
nand U38466 (N_38466,N_37218,N_37666);
nand U38467 (N_38467,N_37024,N_37508);
xor U38468 (N_38468,N_37598,N_37882);
nor U38469 (N_38469,N_37054,N_37909);
and U38470 (N_38470,N_37551,N_37204);
or U38471 (N_38471,N_37030,N_37191);
nor U38472 (N_38472,N_37971,N_37750);
xnor U38473 (N_38473,N_37073,N_37143);
nand U38474 (N_38474,N_37529,N_37061);
xor U38475 (N_38475,N_37951,N_37312);
and U38476 (N_38476,N_37404,N_37928);
or U38477 (N_38477,N_37748,N_37283);
and U38478 (N_38478,N_37693,N_37829);
xnor U38479 (N_38479,N_37674,N_37419);
or U38480 (N_38480,N_37574,N_37594);
and U38481 (N_38481,N_37437,N_37625);
xnor U38482 (N_38482,N_37728,N_37492);
or U38483 (N_38483,N_37984,N_37847);
and U38484 (N_38484,N_37694,N_37768);
and U38485 (N_38485,N_37324,N_37280);
or U38486 (N_38486,N_37720,N_37651);
and U38487 (N_38487,N_37642,N_37825);
nor U38488 (N_38488,N_37088,N_37042);
nor U38489 (N_38489,N_37900,N_37471);
nor U38490 (N_38490,N_37664,N_37137);
or U38491 (N_38491,N_37915,N_37118);
or U38492 (N_38492,N_37262,N_37937);
nor U38493 (N_38493,N_37524,N_37155);
nand U38494 (N_38494,N_37767,N_37729);
and U38495 (N_38495,N_37968,N_37409);
or U38496 (N_38496,N_37560,N_37688);
and U38497 (N_38497,N_37363,N_37072);
or U38498 (N_38498,N_37516,N_37816);
xnor U38499 (N_38499,N_37070,N_37854);
nor U38500 (N_38500,N_37149,N_37772);
or U38501 (N_38501,N_37061,N_37660);
nand U38502 (N_38502,N_37007,N_37639);
or U38503 (N_38503,N_37516,N_37670);
and U38504 (N_38504,N_37444,N_37878);
nor U38505 (N_38505,N_37000,N_37259);
or U38506 (N_38506,N_37256,N_37725);
nand U38507 (N_38507,N_37369,N_37350);
nor U38508 (N_38508,N_37767,N_37868);
nor U38509 (N_38509,N_37738,N_37325);
xnor U38510 (N_38510,N_37951,N_37310);
and U38511 (N_38511,N_37703,N_37157);
nand U38512 (N_38512,N_37358,N_37333);
xor U38513 (N_38513,N_37082,N_37911);
or U38514 (N_38514,N_37463,N_37234);
nor U38515 (N_38515,N_37404,N_37408);
nor U38516 (N_38516,N_37450,N_37371);
nand U38517 (N_38517,N_37517,N_37573);
nor U38518 (N_38518,N_37990,N_37842);
xnor U38519 (N_38519,N_37927,N_37625);
or U38520 (N_38520,N_37110,N_37371);
nand U38521 (N_38521,N_37904,N_37626);
nor U38522 (N_38522,N_37606,N_37436);
nor U38523 (N_38523,N_37665,N_37226);
nor U38524 (N_38524,N_37029,N_37218);
nand U38525 (N_38525,N_37103,N_37642);
and U38526 (N_38526,N_37404,N_37701);
nand U38527 (N_38527,N_37678,N_37567);
xor U38528 (N_38528,N_37949,N_37278);
xor U38529 (N_38529,N_37766,N_37658);
xnor U38530 (N_38530,N_37546,N_37068);
nand U38531 (N_38531,N_37772,N_37217);
nand U38532 (N_38532,N_37867,N_37325);
or U38533 (N_38533,N_37443,N_37626);
nor U38534 (N_38534,N_37878,N_37511);
or U38535 (N_38535,N_37478,N_37151);
and U38536 (N_38536,N_37990,N_37355);
and U38537 (N_38537,N_37805,N_37961);
xnor U38538 (N_38538,N_37855,N_37204);
nor U38539 (N_38539,N_37373,N_37184);
nor U38540 (N_38540,N_37305,N_37224);
nor U38541 (N_38541,N_37702,N_37038);
and U38542 (N_38542,N_37904,N_37576);
and U38543 (N_38543,N_37936,N_37982);
nor U38544 (N_38544,N_37361,N_37227);
nor U38545 (N_38545,N_37074,N_37997);
nand U38546 (N_38546,N_37693,N_37362);
or U38547 (N_38547,N_37073,N_37252);
and U38548 (N_38548,N_37701,N_37602);
xnor U38549 (N_38549,N_37637,N_37590);
or U38550 (N_38550,N_37352,N_37092);
xnor U38551 (N_38551,N_37407,N_37692);
xor U38552 (N_38552,N_37926,N_37631);
or U38553 (N_38553,N_37981,N_37829);
and U38554 (N_38554,N_37063,N_37579);
nor U38555 (N_38555,N_37210,N_37085);
nor U38556 (N_38556,N_37603,N_37325);
nand U38557 (N_38557,N_37837,N_37463);
nor U38558 (N_38558,N_37559,N_37723);
nand U38559 (N_38559,N_37166,N_37443);
nand U38560 (N_38560,N_37192,N_37611);
nor U38561 (N_38561,N_37391,N_37869);
nand U38562 (N_38562,N_37098,N_37884);
nand U38563 (N_38563,N_37150,N_37149);
nand U38564 (N_38564,N_37287,N_37400);
nand U38565 (N_38565,N_37078,N_37336);
nor U38566 (N_38566,N_37895,N_37852);
or U38567 (N_38567,N_37305,N_37966);
xor U38568 (N_38568,N_37201,N_37495);
or U38569 (N_38569,N_37679,N_37896);
or U38570 (N_38570,N_37200,N_37893);
and U38571 (N_38571,N_37283,N_37556);
or U38572 (N_38572,N_37809,N_37329);
nand U38573 (N_38573,N_37138,N_37332);
nand U38574 (N_38574,N_37113,N_37044);
and U38575 (N_38575,N_37379,N_37600);
xnor U38576 (N_38576,N_37005,N_37998);
nor U38577 (N_38577,N_37492,N_37498);
or U38578 (N_38578,N_37189,N_37601);
nor U38579 (N_38579,N_37827,N_37784);
nand U38580 (N_38580,N_37318,N_37551);
nor U38581 (N_38581,N_37121,N_37798);
nor U38582 (N_38582,N_37583,N_37231);
xor U38583 (N_38583,N_37546,N_37325);
and U38584 (N_38584,N_37361,N_37547);
nor U38585 (N_38585,N_37807,N_37501);
xor U38586 (N_38586,N_37353,N_37617);
nand U38587 (N_38587,N_37386,N_37732);
nor U38588 (N_38588,N_37755,N_37227);
or U38589 (N_38589,N_37488,N_37552);
xnor U38590 (N_38590,N_37208,N_37568);
and U38591 (N_38591,N_37504,N_37525);
or U38592 (N_38592,N_37287,N_37039);
and U38593 (N_38593,N_37158,N_37989);
nor U38594 (N_38594,N_37863,N_37689);
and U38595 (N_38595,N_37644,N_37584);
nor U38596 (N_38596,N_37408,N_37539);
or U38597 (N_38597,N_37619,N_37074);
and U38598 (N_38598,N_37760,N_37648);
or U38599 (N_38599,N_37396,N_37661);
nand U38600 (N_38600,N_37010,N_37454);
and U38601 (N_38601,N_37732,N_37322);
and U38602 (N_38602,N_37023,N_37209);
nor U38603 (N_38603,N_37767,N_37159);
nand U38604 (N_38604,N_37873,N_37722);
xnor U38605 (N_38605,N_37016,N_37716);
xor U38606 (N_38606,N_37304,N_37838);
nor U38607 (N_38607,N_37983,N_37067);
and U38608 (N_38608,N_37445,N_37278);
and U38609 (N_38609,N_37026,N_37698);
or U38610 (N_38610,N_37675,N_37743);
or U38611 (N_38611,N_37034,N_37762);
xnor U38612 (N_38612,N_37012,N_37972);
nand U38613 (N_38613,N_37326,N_37436);
or U38614 (N_38614,N_37852,N_37334);
and U38615 (N_38615,N_37094,N_37828);
and U38616 (N_38616,N_37270,N_37432);
xnor U38617 (N_38617,N_37573,N_37114);
nor U38618 (N_38618,N_37561,N_37837);
xor U38619 (N_38619,N_37464,N_37050);
xnor U38620 (N_38620,N_37925,N_37720);
or U38621 (N_38621,N_37940,N_37075);
xnor U38622 (N_38622,N_37308,N_37979);
or U38623 (N_38623,N_37931,N_37671);
and U38624 (N_38624,N_37933,N_37204);
xor U38625 (N_38625,N_37914,N_37766);
nand U38626 (N_38626,N_37565,N_37324);
nor U38627 (N_38627,N_37873,N_37746);
xor U38628 (N_38628,N_37321,N_37222);
or U38629 (N_38629,N_37909,N_37292);
nand U38630 (N_38630,N_37931,N_37147);
nand U38631 (N_38631,N_37022,N_37704);
nor U38632 (N_38632,N_37700,N_37549);
xnor U38633 (N_38633,N_37568,N_37665);
xnor U38634 (N_38634,N_37354,N_37805);
xnor U38635 (N_38635,N_37158,N_37349);
nand U38636 (N_38636,N_37543,N_37595);
nand U38637 (N_38637,N_37372,N_37651);
or U38638 (N_38638,N_37666,N_37672);
and U38639 (N_38639,N_37623,N_37879);
nor U38640 (N_38640,N_37681,N_37775);
xnor U38641 (N_38641,N_37162,N_37549);
nand U38642 (N_38642,N_37031,N_37746);
nor U38643 (N_38643,N_37863,N_37542);
xnor U38644 (N_38644,N_37261,N_37560);
or U38645 (N_38645,N_37017,N_37297);
and U38646 (N_38646,N_37159,N_37003);
or U38647 (N_38647,N_37559,N_37113);
nor U38648 (N_38648,N_37427,N_37177);
nor U38649 (N_38649,N_37445,N_37932);
and U38650 (N_38650,N_37628,N_37374);
xnor U38651 (N_38651,N_37127,N_37616);
xnor U38652 (N_38652,N_37196,N_37463);
or U38653 (N_38653,N_37721,N_37089);
and U38654 (N_38654,N_37605,N_37870);
nor U38655 (N_38655,N_37162,N_37816);
xor U38656 (N_38656,N_37956,N_37757);
nor U38657 (N_38657,N_37524,N_37647);
nand U38658 (N_38658,N_37951,N_37091);
or U38659 (N_38659,N_37652,N_37514);
or U38660 (N_38660,N_37221,N_37301);
nand U38661 (N_38661,N_37300,N_37643);
and U38662 (N_38662,N_37251,N_37153);
nand U38663 (N_38663,N_37261,N_37506);
nand U38664 (N_38664,N_37662,N_37948);
and U38665 (N_38665,N_37826,N_37499);
nand U38666 (N_38666,N_37720,N_37787);
nor U38667 (N_38667,N_37370,N_37161);
or U38668 (N_38668,N_37271,N_37849);
nor U38669 (N_38669,N_37374,N_37173);
xnor U38670 (N_38670,N_37608,N_37838);
nor U38671 (N_38671,N_37288,N_37599);
nand U38672 (N_38672,N_37561,N_37388);
xor U38673 (N_38673,N_37875,N_37613);
nor U38674 (N_38674,N_37669,N_37624);
nand U38675 (N_38675,N_37092,N_37895);
xor U38676 (N_38676,N_37132,N_37198);
nor U38677 (N_38677,N_37337,N_37203);
xnor U38678 (N_38678,N_37436,N_37174);
nor U38679 (N_38679,N_37192,N_37242);
nand U38680 (N_38680,N_37532,N_37430);
nand U38681 (N_38681,N_37009,N_37861);
nor U38682 (N_38682,N_37096,N_37176);
and U38683 (N_38683,N_37718,N_37906);
or U38684 (N_38684,N_37342,N_37310);
xor U38685 (N_38685,N_37755,N_37652);
and U38686 (N_38686,N_37914,N_37840);
xor U38687 (N_38687,N_37444,N_37518);
nand U38688 (N_38688,N_37951,N_37098);
and U38689 (N_38689,N_37421,N_37276);
nor U38690 (N_38690,N_37321,N_37548);
xnor U38691 (N_38691,N_37573,N_37506);
nor U38692 (N_38692,N_37653,N_37987);
or U38693 (N_38693,N_37791,N_37036);
or U38694 (N_38694,N_37507,N_37003);
and U38695 (N_38695,N_37259,N_37845);
and U38696 (N_38696,N_37259,N_37740);
xnor U38697 (N_38697,N_37805,N_37757);
nor U38698 (N_38698,N_37738,N_37682);
xnor U38699 (N_38699,N_37959,N_37423);
nand U38700 (N_38700,N_37869,N_37402);
and U38701 (N_38701,N_37023,N_37141);
nor U38702 (N_38702,N_37848,N_37835);
or U38703 (N_38703,N_37637,N_37426);
and U38704 (N_38704,N_37489,N_37607);
and U38705 (N_38705,N_37844,N_37777);
nor U38706 (N_38706,N_37923,N_37884);
xnor U38707 (N_38707,N_37980,N_37585);
and U38708 (N_38708,N_37384,N_37429);
or U38709 (N_38709,N_37546,N_37798);
nor U38710 (N_38710,N_37998,N_37479);
xnor U38711 (N_38711,N_37943,N_37327);
nor U38712 (N_38712,N_37573,N_37385);
nor U38713 (N_38713,N_37512,N_37601);
or U38714 (N_38714,N_37583,N_37552);
or U38715 (N_38715,N_37859,N_37061);
and U38716 (N_38716,N_37532,N_37163);
nor U38717 (N_38717,N_37317,N_37575);
or U38718 (N_38718,N_37713,N_37200);
and U38719 (N_38719,N_37752,N_37312);
or U38720 (N_38720,N_37861,N_37550);
xor U38721 (N_38721,N_37585,N_37468);
xor U38722 (N_38722,N_37099,N_37337);
and U38723 (N_38723,N_37885,N_37878);
xor U38724 (N_38724,N_37816,N_37034);
nor U38725 (N_38725,N_37120,N_37638);
or U38726 (N_38726,N_37094,N_37573);
nor U38727 (N_38727,N_37691,N_37217);
or U38728 (N_38728,N_37568,N_37939);
xor U38729 (N_38729,N_37842,N_37042);
nand U38730 (N_38730,N_37308,N_37775);
or U38731 (N_38731,N_37036,N_37272);
and U38732 (N_38732,N_37592,N_37861);
xnor U38733 (N_38733,N_37373,N_37615);
nor U38734 (N_38734,N_37943,N_37587);
and U38735 (N_38735,N_37919,N_37496);
or U38736 (N_38736,N_37529,N_37911);
and U38737 (N_38737,N_37629,N_37654);
xnor U38738 (N_38738,N_37128,N_37549);
xnor U38739 (N_38739,N_37936,N_37729);
or U38740 (N_38740,N_37317,N_37146);
xor U38741 (N_38741,N_37414,N_37523);
nor U38742 (N_38742,N_37776,N_37979);
nand U38743 (N_38743,N_37961,N_37233);
and U38744 (N_38744,N_37745,N_37979);
xnor U38745 (N_38745,N_37241,N_37691);
nor U38746 (N_38746,N_37088,N_37771);
nand U38747 (N_38747,N_37554,N_37283);
nand U38748 (N_38748,N_37014,N_37657);
xor U38749 (N_38749,N_37645,N_37195);
nand U38750 (N_38750,N_37700,N_37820);
nand U38751 (N_38751,N_37661,N_37940);
or U38752 (N_38752,N_37496,N_37091);
or U38753 (N_38753,N_37171,N_37824);
nor U38754 (N_38754,N_37413,N_37048);
xor U38755 (N_38755,N_37428,N_37684);
nand U38756 (N_38756,N_37997,N_37667);
nor U38757 (N_38757,N_37489,N_37267);
nor U38758 (N_38758,N_37421,N_37803);
and U38759 (N_38759,N_37191,N_37269);
or U38760 (N_38760,N_37927,N_37021);
nor U38761 (N_38761,N_37007,N_37495);
nand U38762 (N_38762,N_37353,N_37911);
nor U38763 (N_38763,N_37297,N_37116);
or U38764 (N_38764,N_37385,N_37614);
or U38765 (N_38765,N_37217,N_37427);
xnor U38766 (N_38766,N_37204,N_37526);
or U38767 (N_38767,N_37036,N_37569);
or U38768 (N_38768,N_37494,N_37858);
or U38769 (N_38769,N_37265,N_37720);
nand U38770 (N_38770,N_37124,N_37759);
xnor U38771 (N_38771,N_37992,N_37379);
or U38772 (N_38772,N_37589,N_37109);
nand U38773 (N_38773,N_37090,N_37161);
or U38774 (N_38774,N_37914,N_37759);
nor U38775 (N_38775,N_37564,N_37222);
nor U38776 (N_38776,N_37974,N_37529);
nor U38777 (N_38777,N_37679,N_37787);
xnor U38778 (N_38778,N_37299,N_37007);
nand U38779 (N_38779,N_37496,N_37233);
or U38780 (N_38780,N_37136,N_37984);
xor U38781 (N_38781,N_37289,N_37333);
xnor U38782 (N_38782,N_37299,N_37649);
or U38783 (N_38783,N_37645,N_37502);
and U38784 (N_38784,N_37208,N_37091);
or U38785 (N_38785,N_37760,N_37797);
xor U38786 (N_38786,N_37169,N_37248);
xnor U38787 (N_38787,N_37907,N_37903);
nand U38788 (N_38788,N_37941,N_37223);
or U38789 (N_38789,N_37884,N_37655);
nand U38790 (N_38790,N_37848,N_37932);
xnor U38791 (N_38791,N_37217,N_37892);
nand U38792 (N_38792,N_37330,N_37058);
nor U38793 (N_38793,N_37996,N_37629);
nand U38794 (N_38794,N_37345,N_37327);
nand U38795 (N_38795,N_37391,N_37807);
or U38796 (N_38796,N_37952,N_37687);
xor U38797 (N_38797,N_37049,N_37202);
nor U38798 (N_38798,N_37385,N_37477);
nand U38799 (N_38799,N_37463,N_37082);
xor U38800 (N_38800,N_37324,N_37291);
nand U38801 (N_38801,N_37918,N_37649);
and U38802 (N_38802,N_37196,N_37985);
nand U38803 (N_38803,N_37398,N_37199);
xnor U38804 (N_38804,N_37815,N_37229);
nand U38805 (N_38805,N_37449,N_37504);
xor U38806 (N_38806,N_37051,N_37912);
and U38807 (N_38807,N_37078,N_37202);
xnor U38808 (N_38808,N_37782,N_37133);
nand U38809 (N_38809,N_37621,N_37323);
nor U38810 (N_38810,N_37644,N_37540);
nand U38811 (N_38811,N_37533,N_37679);
nand U38812 (N_38812,N_37010,N_37053);
xnor U38813 (N_38813,N_37949,N_37997);
nor U38814 (N_38814,N_37573,N_37720);
nor U38815 (N_38815,N_37010,N_37402);
nor U38816 (N_38816,N_37207,N_37720);
xnor U38817 (N_38817,N_37316,N_37010);
nor U38818 (N_38818,N_37818,N_37085);
xor U38819 (N_38819,N_37169,N_37323);
or U38820 (N_38820,N_37548,N_37537);
nor U38821 (N_38821,N_37652,N_37314);
nand U38822 (N_38822,N_37241,N_37559);
nor U38823 (N_38823,N_37704,N_37178);
nand U38824 (N_38824,N_37003,N_37294);
xnor U38825 (N_38825,N_37441,N_37070);
xnor U38826 (N_38826,N_37569,N_37847);
nor U38827 (N_38827,N_37018,N_37961);
or U38828 (N_38828,N_37990,N_37294);
or U38829 (N_38829,N_37770,N_37949);
or U38830 (N_38830,N_37383,N_37137);
nor U38831 (N_38831,N_37119,N_37383);
xor U38832 (N_38832,N_37543,N_37958);
or U38833 (N_38833,N_37934,N_37544);
nor U38834 (N_38834,N_37845,N_37531);
nor U38835 (N_38835,N_37446,N_37073);
nor U38836 (N_38836,N_37725,N_37639);
nand U38837 (N_38837,N_37041,N_37429);
nand U38838 (N_38838,N_37211,N_37729);
nor U38839 (N_38839,N_37252,N_37270);
xor U38840 (N_38840,N_37188,N_37319);
nor U38841 (N_38841,N_37132,N_37348);
xor U38842 (N_38842,N_37256,N_37781);
and U38843 (N_38843,N_37732,N_37141);
xnor U38844 (N_38844,N_37195,N_37921);
or U38845 (N_38845,N_37381,N_37501);
and U38846 (N_38846,N_37450,N_37511);
nand U38847 (N_38847,N_37042,N_37271);
and U38848 (N_38848,N_37061,N_37408);
or U38849 (N_38849,N_37350,N_37743);
xnor U38850 (N_38850,N_37571,N_37965);
or U38851 (N_38851,N_37074,N_37641);
or U38852 (N_38852,N_37199,N_37549);
and U38853 (N_38853,N_37359,N_37285);
xor U38854 (N_38854,N_37006,N_37482);
xor U38855 (N_38855,N_37098,N_37207);
and U38856 (N_38856,N_37967,N_37769);
and U38857 (N_38857,N_37617,N_37701);
nor U38858 (N_38858,N_37761,N_37034);
and U38859 (N_38859,N_37987,N_37113);
xnor U38860 (N_38860,N_37774,N_37458);
and U38861 (N_38861,N_37294,N_37000);
or U38862 (N_38862,N_37224,N_37055);
nor U38863 (N_38863,N_37617,N_37624);
and U38864 (N_38864,N_37718,N_37525);
xnor U38865 (N_38865,N_37630,N_37381);
or U38866 (N_38866,N_37585,N_37010);
nor U38867 (N_38867,N_37351,N_37249);
nor U38868 (N_38868,N_37958,N_37055);
or U38869 (N_38869,N_37210,N_37862);
nand U38870 (N_38870,N_37624,N_37385);
nand U38871 (N_38871,N_37835,N_37318);
xnor U38872 (N_38872,N_37711,N_37574);
nor U38873 (N_38873,N_37849,N_37643);
nand U38874 (N_38874,N_37356,N_37940);
and U38875 (N_38875,N_37255,N_37917);
nand U38876 (N_38876,N_37450,N_37427);
or U38877 (N_38877,N_37687,N_37792);
xnor U38878 (N_38878,N_37804,N_37422);
xnor U38879 (N_38879,N_37769,N_37928);
or U38880 (N_38880,N_37041,N_37698);
nand U38881 (N_38881,N_37989,N_37692);
nor U38882 (N_38882,N_37881,N_37632);
xor U38883 (N_38883,N_37690,N_37661);
and U38884 (N_38884,N_37071,N_37540);
nor U38885 (N_38885,N_37778,N_37851);
nor U38886 (N_38886,N_37118,N_37384);
and U38887 (N_38887,N_37141,N_37230);
or U38888 (N_38888,N_37453,N_37002);
xnor U38889 (N_38889,N_37434,N_37526);
nor U38890 (N_38890,N_37630,N_37431);
xnor U38891 (N_38891,N_37879,N_37091);
nor U38892 (N_38892,N_37112,N_37120);
xnor U38893 (N_38893,N_37021,N_37381);
nand U38894 (N_38894,N_37206,N_37252);
and U38895 (N_38895,N_37434,N_37860);
and U38896 (N_38896,N_37982,N_37592);
xor U38897 (N_38897,N_37678,N_37108);
nor U38898 (N_38898,N_37580,N_37088);
and U38899 (N_38899,N_37563,N_37328);
nand U38900 (N_38900,N_37836,N_37962);
xnor U38901 (N_38901,N_37122,N_37139);
xnor U38902 (N_38902,N_37592,N_37733);
nand U38903 (N_38903,N_37549,N_37450);
and U38904 (N_38904,N_37909,N_37012);
and U38905 (N_38905,N_37633,N_37282);
xor U38906 (N_38906,N_37629,N_37740);
nand U38907 (N_38907,N_37827,N_37335);
xnor U38908 (N_38908,N_37193,N_37881);
nor U38909 (N_38909,N_37518,N_37658);
nand U38910 (N_38910,N_37718,N_37394);
nor U38911 (N_38911,N_37794,N_37166);
or U38912 (N_38912,N_37248,N_37920);
nand U38913 (N_38913,N_37674,N_37024);
or U38914 (N_38914,N_37607,N_37520);
xor U38915 (N_38915,N_37082,N_37606);
xor U38916 (N_38916,N_37597,N_37652);
and U38917 (N_38917,N_37253,N_37562);
xor U38918 (N_38918,N_37437,N_37171);
xor U38919 (N_38919,N_37065,N_37752);
nand U38920 (N_38920,N_37060,N_37961);
nand U38921 (N_38921,N_37105,N_37829);
xor U38922 (N_38922,N_37150,N_37074);
or U38923 (N_38923,N_37001,N_37803);
nand U38924 (N_38924,N_37479,N_37495);
and U38925 (N_38925,N_37423,N_37212);
and U38926 (N_38926,N_37946,N_37165);
nand U38927 (N_38927,N_37466,N_37288);
nor U38928 (N_38928,N_37912,N_37786);
and U38929 (N_38929,N_37233,N_37916);
nand U38930 (N_38930,N_37057,N_37463);
or U38931 (N_38931,N_37092,N_37178);
nand U38932 (N_38932,N_37607,N_37820);
xor U38933 (N_38933,N_37552,N_37278);
xnor U38934 (N_38934,N_37836,N_37143);
and U38935 (N_38935,N_37669,N_37742);
xnor U38936 (N_38936,N_37110,N_37240);
nor U38937 (N_38937,N_37228,N_37939);
nand U38938 (N_38938,N_37562,N_37410);
and U38939 (N_38939,N_37790,N_37625);
nor U38940 (N_38940,N_37714,N_37301);
or U38941 (N_38941,N_37518,N_37915);
nand U38942 (N_38942,N_37192,N_37323);
or U38943 (N_38943,N_37456,N_37378);
and U38944 (N_38944,N_37346,N_37954);
or U38945 (N_38945,N_37692,N_37338);
nor U38946 (N_38946,N_37370,N_37026);
nand U38947 (N_38947,N_37110,N_37190);
or U38948 (N_38948,N_37765,N_37984);
or U38949 (N_38949,N_37602,N_37798);
nor U38950 (N_38950,N_37461,N_37496);
or U38951 (N_38951,N_37929,N_37183);
nand U38952 (N_38952,N_37923,N_37302);
and U38953 (N_38953,N_37217,N_37101);
and U38954 (N_38954,N_37619,N_37348);
xnor U38955 (N_38955,N_37241,N_37259);
nor U38956 (N_38956,N_37938,N_37846);
nand U38957 (N_38957,N_37512,N_37155);
xnor U38958 (N_38958,N_37903,N_37104);
and U38959 (N_38959,N_37817,N_37925);
nand U38960 (N_38960,N_37610,N_37177);
xnor U38961 (N_38961,N_37954,N_37413);
nor U38962 (N_38962,N_37868,N_37489);
and U38963 (N_38963,N_37053,N_37264);
and U38964 (N_38964,N_37950,N_37227);
nand U38965 (N_38965,N_37614,N_37373);
nand U38966 (N_38966,N_37982,N_37367);
and U38967 (N_38967,N_37085,N_37611);
nor U38968 (N_38968,N_37332,N_37405);
nand U38969 (N_38969,N_37691,N_37594);
or U38970 (N_38970,N_37954,N_37016);
nor U38971 (N_38971,N_37093,N_37068);
and U38972 (N_38972,N_37111,N_37215);
nand U38973 (N_38973,N_37299,N_37866);
nand U38974 (N_38974,N_37885,N_37803);
nor U38975 (N_38975,N_37575,N_37383);
or U38976 (N_38976,N_37155,N_37133);
or U38977 (N_38977,N_37621,N_37700);
and U38978 (N_38978,N_37325,N_37365);
nor U38979 (N_38979,N_37866,N_37091);
and U38980 (N_38980,N_37973,N_37402);
or U38981 (N_38981,N_37314,N_37084);
and U38982 (N_38982,N_37876,N_37555);
xor U38983 (N_38983,N_37207,N_37734);
and U38984 (N_38984,N_37958,N_37830);
nand U38985 (N_38985,N_37400,N_37860);
nor U38986 (N_38986,N_37757,N_37289);
nand U38987 (N_38987,N_37434,N_37404);
nand U38988 (N_38988,N_37328,N_37228);
or U38989 (N_38989,N_37295,N_37857);
and U38990 (N_38990,N_37663,N_37555);
xnor U38991 (N_38991,N_37570,N_37643);
and U38992 (N_38992,N_37522,N_37508);
or U38993 (N_38993,N_37743,N_37626);
nand U38994 (N_38994,N_37233,N_37357);
nand U38995 (N_38995,N_37121,N_37909);
nor U38996 (N_38996,N_37193,N_37445);
nand U38997 (N_38997,N_37019,N_37167);
xnor U38998 (N_38998,N_37222,N_37170);
nand U38999 (N_38999,N_37860,N_37640);
nor U39000 (N_39000,N_38311,N_38372);
or U39001 (N_39001,N_38367,N_38738);
nand U39002 (N_39002,N_38499,N_38930);
and U39003 (N_39003,N_38170,N_38585);
or U39004 (N_39004,N_38080,N_38235);
nor U39005 (N_39005,N_38378,N_38414);
or U39006 (N_39006,N_38716,N_38489);
or U39007 (N_39007,N_38121,N_38990);
and U39008 (N_39008,N_38377,N_38838);
or U39009 (N_39009,N_38784,N_38652);
and U39010 (N_39010,N_38016,N_38409);
and U39011 (N_39011,N_38219,N_38146);
and U39012 (N_39012,N_38233,N_38978);
or U39013 (N_39013,N_38393,N_38073);
or U39014 (N_39014,N_38906,N_38256);
and U39015 (N_39015,N_38917,N_38529);
or U39016 (N_39016,N_38515,N_38159);
nor U39017 (N_39017,N_38565,N_38018);
xor U39018 (N_39018,N_38316,N_38480);
nand U39019 (N_39019,N_38063,N_38005);
xnor U39020 (N_39020,N_38527,N_38718);
and U39021 (N_39021,N_38120,N_38833);
nor U39022 (N_39022,N_38555,N_38521);
xor U39023 (N_39023,N_38925,N_38487);
xnor U39024 (N_39024,N_38750,N_38607);
nor U39025 (N_39025,N_38991,N_38425);
nor U39026 (N_39026,N_38344,N_38180);
or U39027 (N_39027,N_38185,N_38891);
nand U39028 (N_39028,N_38024,N_38104);
xor U39029 (N_39029,N_38950,N_38254);
xnor U39030 (N_39030,N_38835,N_38376);
xor U39031 (N_39031,N_38786,N_38528);
or U39032 (N_39032,N_38986,N_38910);
nand U39033 (N_39033,N_38899,N_38079);
nor U39034 (N_39034,N_38535,N_38503);
xnor U39035 (N_39035,N_38187,N_38280);
and U39036 (N_39036,N_38215,N_38475);
nor U39037 (N_39037,N_38935,N_38782);
and U39038 (N_39038,N_38894,N_38176);
and U39039 (N_39039,N_38457,N_38613);
and U39040 (N_39040,N_38646,N_38711);
and U39041 (N_39041,N_38143,N_38203);
or U39042 (N_39042,N_38883,N_38597);
and U39043 (N_39043,N_38395,N_38186);
xor U39044 (N_39044,N_38987,N_38774);
nand U39045 (N_39045,N_38325,N_38928);
and U39046 (N_39046,N_38798,N_38920);
nor U39047 (N_39047,N_38516,N_38023);
and U39048 (N_39048,N_38275,N_38569);
nand U39049 (N_39049,N_38916,N_38909);
nor U39050 (N_39050,N_38098,N_38568);
or U39051 (N_39051,N_38757,N_38197);
and U39052 (N_39052,N_38412,N_38262);
xor U39053 (N_39053,N_38322,N_38857);
nor U39054 (N_39054,N_38831,N_38299);
nand U39055 (N_39055,N_38217,N_38710);
or U39056 (N_39056,N_38057,N_38856);
and U39057 (N_39057,N_38611,N_38670);
and U39058 (N_39058,N_38240,N_38164);
or U39059 (N_39059,N_38058,N_38125);
xor U39060 (N_39060,N_38596,N_38654);
nand U39061 (N_39061,N_38735,N_38175);
nor U39062 (N_39062,N_38394,N_38476);
or U39063 (N_39063,N_38216,N_38497);
and U39064 (N_39064,N_38531,N_38207);
nand U39065 (N_39065,N_38327,N_38470);
xor U39066 (N_39066,N_38971,N_38149);
xor U39067 (N_39067,N_38934,N_38863);
nand U39068 (N_39068,N_38099,N_38313);
nor U39069 (N_39069,N_38865,N_38882);
nor U39070 (N_39070,N_38763,N_38255);
nor U39071 (N_39071,N_38000,N_38446);
or U39072 (N_39072,N_38343,N_38397);
nand U39073 (N_39073,N_38131,N_38672);
xnor U39074 (N_39074,N_38329,N_38214);
nand U39075 (N_39075,N_38498,N_38723);
and U39076 (N_39076,N_38403,N_38806);
and U39077 (N_39077,N_38491,N_38382);
xor U39078 (N_39078,N_38231,N_38713);
nand U39079 (N_39079,N_38967,N_38730);
nand U39080 (N_39080,N_38158,N_38250);
or U39081 (N_39081,N_38020,N_38705);
and U39082 (N_39082,N_38418,N_38651);
nand U39083 (N_39083,N_38224,N_38247);
or U39084 (N_39084,N_38668,N_38827);
xnor U39085 (N_39085,N_38828,N_38427);
xor U39086 (N_39086,N_38054,N_38939);
and U39087 (N_39087,N_38157,N_38717);
nor U39088 (N_39088,N_38604,N_38629);
and U39089 (N_39089,N_38993,N_38793);
nand U39090 (N_39090,N_38444,N_38645);
xor U39091 (N_39091,N_38051,N_38896);
nor U39092 (N_39092,N_38663,N_38421);
nand U39093 (N_39093,N_38765,N_38434);
or U39094 (N_39094,N_38577,N_38252);
nor U39095 (N_39095,N_38291,N_38388);
nand U39096 (N_39096,N_38892,N_38748);
xor U39097 (N_39097,N_38573,N_38901);
or U39098 (N_39098,N_38257,N_38505);
xnor U39099 (N_39099,N_38832,N_38044);
nand U39100 (N_39100,N_38741,N_38830);
and U39101 (N_39101,N_38969,N_38155);
xnor U39102 (N_39102,N_38558,N_38113);
nor U39103 (N_39103,N_38360,N_38603);
nand U39104 (N_39104,N_38649,N_38996);
nor U39105 (N_39105,N_38511,N_38606);
nand U39106 (N_39106,N_38460,N_38465);
xnor U39107 (N_39107,N_38681,N_38324);
xor U39108 (N_39108,N_38734,N_38998);
nand U39109 (N_39109,N_38053,N_38799);
xnor U39110 (N_39110,N_38072,N_38789);
or U39111 (N_39111,N_38762,N_38512);
xnor U39112 (N_39112,N_38825,N_38405);
nand U39113 (N_39113,N_38453,N_38593);
xor U39114 (N_39114,N_38130,N_38241);
or U39115 (N_39115,N_38972,N_38030);
and U39116 (N_39116,N_38223,N_38204);
nand U39117 (N_39117,N_38251,N_38253);
nand U39118 (N_39118,N_38638,N_38068);
nand U39119 (N_39119,N_38980,N_38676);
nand U39120 (N_39120,N_38188,N_38191);
xor U39121 (N_39121,N_38644,N_38945);
xor U39122 (N_39122,N_38635,N_38881);
or U39123 (N_39123,N_38974,N_38583);
nand U39124 (N_39124,N_38225,N_38055);
nor U39125 (N_39125,N_38123,N_38334);
and U39126 (N_39126,N_38486,N_38745);
xor U39127 (N_39127,N_38727,N_38504);
nand U39128 (N_39128,N_38743,N_38625);
or U39129 (N_39129,N_38539,N_38703);
or U39130 (N_39130,N_38758,N_38348);
nor U39131 (N_39131,N_38318,N_38586);
or U39132 (N_39132,N_38809,N_38085);
nor U39133 (N_39133,N_38093,N_38747);
or U39134 (N_39134,N_38228,N_38979);
or U39135 (N_39135,N_38541,N_38420);
xor U39136 (N_39136,N_38634,N_38728);
or U39137 (N_39137,N_38379,N_38074);
or U39138 (N_39138,N_38419,N_38006);
xor U39139 (N_39139,N_38648,N_38818);
nor U39140 (N_39140,N_38477,N_38566);
and U39141 (N_39141,N_38304,N_38069);
and U39142 (N_39142,N_38374,N_38326);
nor U39143 (N_39143,N_38685,N_38265);
nand U39144 (N_39144,N_38689,N_38742);
or U39145 (N_39145,N_38801,N_38153);
or U39146 (N_39146,N_38036,N_38732);
or U39147 (N_39147,N_38872,N_38154);
or U39148 (N_39148,N_38813,N_38640);
or U39149 (N_39149,N_38542,N_38824);
and U39150 (N_39150,N_38242,N_38234);
and U39151 (N_39151,N_38462,N_38870);
nand U39152 (N_39152,N_38563,N_38594);
nor U39153 (N_39153,N_38683,N_38712);
nand U39154 (N_39154,N_38954,N_38790);
nor U39155 (N_39155,N_38864,N_38009);
and U39156 (N_39156,N_38315,N_38688);
nor U39157 (N_39157,N_38959,N_38112);
or U39158 (N_39158,N_38867,N_38684);
and U39159 (N_39159,N_38513,N_38178);
and U39160 (N_39160,N_38386,N_38336);
and U39161 (N_39161,N_38821,N_38694);
xor U39162 (N_39162,N_38796,N_38706);
nor U39163 (N_39163,N_38693,N_38229);
nor U39164 (N_39164,N_38519,N_38246);
nand U39165 (N_39165,N_38862,N_38854);
or U39166 (N_39166,N_38353,N_38171);
xnor U39167 (N_39167,N_38321,N_38720);
xor U39168 (N_39168,N_38888,N_38089);
nor U39169 (N_39169,N_38087,N_38855);
nor U39170 (N_39170,N_38754,N_38064);
nor U39171 (N_39171,N_38352,N_38822);
xor U39172 (N_39172,N_38687,N_38298);
nor U39173 (N_39173,N_38135,N_38236);
or U39174 (N_39174,N_38346,N_38340);
or U39175 (N_39175,N_38387,N_38680);
and U39176 (N_39176,N_38037,N_38780);
and U39177 (N_39177,N_38156,N_38042);
and U39178 (N_39178,N_38576,N_38468);
nand U39179 (N_39179,N_38788,N_38454);
and U39180 (N_39180,N_38495,N_38942);
xnor U39181 (N_39181,N_38391,N_38205);
nor U39182 (N_39182,N_38385,N_38759);
or U39183 (N_39183,N_38050,N_38110);
nand U39184 (N_39184,N_38721,N_38808);
nand U39185 (N_39185,N_38261,N_38551);
or U39186 (N_39186,N_38861,N_38218);
or U39187 (N_39187,N_38898,N_38239);
and U39188 (N_39188,N_38283,N_38267);
or U39189 (N_39189,N_38627,N_38438);
and U39190 (N_39190,N_38200,N_38666);
nor U39191 (N_39191,N_38905,N_38097);
xnor U39192 (N_39192,N_38816,N_38167);
nand U39193 (N_39193,N_38548,N_38132);
and U39194 (N_39194,N_38616,N_38027);
nand U39195 (N_39195,N_38608,N_38570);
or U39196 (N_39196,N_38595,N_38332);
and U39197 (N_39197,N_38396,N_38567);
and U39198 (N_39198,N_38671,N_38260);
xor U39199 (N_39199,N_38289,N_38624);
xor U39200 (N_39200,N_38605,N_38556);
or U39201 (N_39201,N_38658,N_38949);
and U39202 (N_39202,N_38049,N_38739);
nand U39203 (N_39203,N_38227,N_38589);
and U39204 (N_39204,N_38439,N_38659);
and U39205 (N_39205,N_38467,N_38614);
xnor U39206 (N_39206,N_38284,N_38105);
or U39207 (N_39207,N_38632,N_38033);
or U39208 (N_39208,N_38363,N_38957);
xor U39209 (N_39209,N_38066,N_38895);
xor U39210 (N_39210,N_38435,N_38769);
and U39211 (N_39211,N_38046,N_38929);
and U39212 (N_39212,N_38746,N_38984);
nor U39213 (N_39213,N_38364,N_38075);
nand U39214 (N_39214,N_38017,N_38545);
and U39215 (N_39215,N_38002,N_38911);
xor U39216 (N_39216,N_38931,N_38041);
nor U39217 (N_39217,N_38494,N_38884);
or U39218 (N_39218,N_38483,N_38966);
nor U39219 (N_39219,N_38664,N_38650);
xnor U39220 (N_39220,N_38781,N_38936);
and U39221 (N_39221,N_38887,N_38144);
nand U39222 (N_39222,N_38775,N_38787);
or U39223 (N_39223,N_38406,N_38707);
and U39224 (N_39224,N_38923,N_38243);
or U39225 (N_39225,N_38198,N_38731);
nor U39226 (N_39226,N_38965,N_38564);
or U39227 (N_39227,N_38709,N_38274);
xnor U39228 (N_39228,N_38698,N_38482);
xor U39229 (N_39229,N_38067,N_38416);
nand U39230 (N_39230,N_38471,N_38797);
nor U39231 (N_39231,N_38128,N_38874);
xor U39232 (N_39232,N_38873,N_38783);
xnor U39233 (N_39233,N_38653,N_38791);
or U39234 (N_39234,N_38669,N_38392);
and U39235 (N_39235,N_38096,N_38270);
nor U39236 (N_39236,N_38590,N_38455);
xor U39237 (N_39237,N_38310,N_38839);
nand U39238 (N_39238,N_38165,N_38485);
or U39239 (N_39239,N_38195,N_38866);
nor U39240 (N_39240,N_38601,N_38244);
and U39241 (N_39241,N_38772,N_38286);
nor U39242 (N_39242,N_38273,N_38598);
nand U39243 (N_39243,N_38922,N_38502);
xnor U39244 (N_39244,N_38660,N_38963);
or U39245 (N_39245,N_38778,N_38411);
nand U39246 (N_39246,N_38724,N_38043);
and U39247 (N_39247,N_38103,N_38501);
nand U39248 (N_39248,N_38140,N_38269);
nand U39249 (N_39249,N_38852,N_38578);
xnor U39250 (N_39250,N_38259,N_38375);
or U39251 (N_39251,N_38450,N_38587);
xor U39252 (N_39252,N_38268,N_38860);
xor U39253 (N_39253,N_38636,N_38021);
xnor U39254 (N_39254,N_38029,N_38859);
and U39255 (N_39255,N_38958,N_38297);
nor U39256 (N_39256,N_38083,N_38961);
xor U39257 (N_39257,N_38662,N_38767);
nor U39258 (N_39258,N_38115,N_38447);
nor U39259 (N_39259,N_38700,N_38600);
nor U39260 (N_39260,N_38307,N_38122);
nand U39261 (N_39261,N_38858,N_38701);
xor U39262 (N_39262,N_38168,N_38179);
or U39263 (N_39263,N_38533,N_38160);
or U39264 (N_39264,N_38880,N_38517);
or U39265 (N_39265,N_38572,N_38071);
xnor U39266 (N_39266,N_38761,N_38014);
nor U39267 (N_39267,N_38915,N_38362);
xor U39268 (N_39268,N_38960,N_38359);
and U39269 (N_39269,N_38696,N_38019);
nand U39270 (N_39270,N_38056,N_38383);
xnor U39271 (N_39271,N_38999,N_38803);
nor U39272 (N_39272,N_38815,N_38506);
nand U39273 (N_39273,N_38704,N_38038);
or U39274 (N_39274,N_38534,N_38845);
nor U39275 (N_39275,N_38619,N_38559);
and U39276 (N_39276,N_38174,N_38912);
nor U39277 (N_39277,N_38190,N_38955);
or U39278 (N_39278,N_38937,N_38312);
and U39279 (N_39279,N_38523,N_38507);
and U39280 (N_39280,N_38118,N_38647);
and U39281 (N_39281,N_38509,N_38389);
xor U39282 (N_39282,N_38903,N_38526);
nor U39283 (N_39283,N_38342,N_38290);
nand U39284 (N_39284,N_38621,N_38970);
nor U39285 (N_39285,N_38161,N_38040);
and U39286 (N_39286,N_38561,N_38337);
and U39287 (N_39287,N_38878,N_38983);
or U39288 (N_39288,N_38520,N_38760);
nand U39289 (N_39289,N_38582,N_38035);
nor U39290 (N_39290,N_38111,N_38012);
nor U39291 (N_39291,N_38641,N_38975);
and U39292 (N_39292,N_38610,N_38390);
nor U39293 (N_39293,N_38142,N_38126);
xor U39294 (N_39294,N_38695,N_38264);
nor U39295 (N_39295,N_38319,N_38442);
xor U39296 (N_39296,N_38794,N_38620);
and U39297 (N_39297,N_38886,N_38380);
and U39298 (N_39298,N_38940,N_38722);
and U39299 (N_39299,N_38443,N_38992);
or U39300 (N_39300,N_38877,N_38220);
nand U39301 (N_39301,N_38173,N_38810);
nor U39302 (N_39302,N_38084,N_38368);
xor U39303 (N_39303,N_38407,N_38719);
and U39304 (N_39304,N_38048,N_38714);
or U39305 (N_39305,N_38306,N_38885);
or U39306 (N_39306,N_38740,N_38773);
and U39307 (N_39307,N_38404,N_38811);
xor U39308 (N_39308,N_38847,N_38221);
or U39309 (N_39309,N_38301,N_38656);
xor U39310 (N_39310,N_38138,N_38061);
and U39311 (N_39311,N_38938,N_38599);
or U39312 (N_39312,N_38837,N_38147);
nor U39313 (N_39313,N_38484,N_38114);
nand U39314 (N_39314,N_38356,N_38472);
nand U39315 (N_39315,N_38779,N_38544);
nand U39316 (N_39316,N_38150,N_38571);
or U39317 (N_39317,N_38557,N_38039);
and U39318 (N_39318,N_38317,N_38490);
nand U39319 (N_39319,N_38091,N_38820);
nor U39320 (N_39320,N_38626,N_38488);
and U39321 (N_39321,N_38550,N_38088);
and U39322 (N_39322,N_38532,N_38423);
nand U39323 (N_39323,N_38162,N_38276);
and U39324 (N_39324,N_38101,N_38819);
nand U39325 (N_39325,N_38366,N_38371);
xnor U39326 (N_39326,N_38851,N_38524);
and U39327 (N_39327,N_38107,N_38744);
or U39328 (N_39328,N_38102,N_38817);
nor U39329 (N_39329,N_38547,N_38538);
nand U39330 (N_39330,N_38622,N_38546);
nor U39331 (N_39331,N_38358,N_38904);
xor U39332 (N_39332,N_38010,N_38031);
or U39333 (N_39333,N_38025,N_38725);
xnor U39334 (N_39334,N_38258,N_38575);
nor U39335 (N_39335,N_38117,N_38052);
and U39336 (N_39336,N_38194,N_38537);
nor U39337 (N_39337,N_38508,N_38034);
nand U39338 (N_39338,N_38733,N_38560);
and U39339 (N_39339,N_38848,N_38410);
and U39340 (N_39340,N_38172,N_38287);
nand U39341 (N_39341,N_38729,N_38417);
xnor U39342 (N_39342,N_38077,N_38481);
nor U39343 (N_39343,N_38095,N_38708);
nand U39344 (N_39344,N_38897,N_38631);
and U39345 (N_39345,N_38726,N_38871);
nor U39346 (N_39346,N_38305,N_38384);
and U39347 (N_39347,N_38690,N_38602);
nor U39348 (N_39348,N_38691,N_38308);
nand U39349 (N_39349,N_38081,N_38633);
nand U39350 (N_39350,N_38953,N_38768);
and U39351 (N_39351,N_38908,N_38090);
or U39352 (N_39352,N_38209,N_38751);
or U39353 (N_39353,N_38500,N_38330);
nand U39354 (N_39354,N_38770,N_38333);
nand U39355 (N_39355,N_38295,N_38426);
or U39356 (N_39356,N_38134,N_38617);
nor U39357 (N_39357,N_38677,N_38540);
or U39358 (N_39358,N_38169,N_38285);
nor U39359 (N_39359,N_38673,N_38192);
nand U39360 (N_39360,N_38588,N_38338);
nand U39361 (N_39361,N_38182,N_38562);
nor U39362 (N_39362,N_38355,N_38226);
nor U39363 (N_39363,N_38238,N_38350);
nor U39364 (N_39364,N_38919,N_38615);
xor U39365 (N_39365,N_38109,N_38682);
and U39366 (N_39366,N_38674,N_38947);
or U39367 (N_39367,N_38357,N_38932);
nor U39368 (N_39368,N_38373,N_38753);
xor U39369 (N_39369,N_38145,N_38479);
or U39370 (N_39370,N_38011,N_38116);
and U39371 (N_39371,N_38849,N_38232);
or U39372 (N_39372,N_38004,N_38846);
and U39373 (N_39373,N_38292,N_38492);
or U39374 (N_39374,N_38944,N_38853);
nand U39375 (N_39375,N_38844,N_38510);
or U39376 (N_39376,N_38459,N_38400);
nor U39377 (N_39377,N_38248,N_38592);
or U39378 (N_39378,N_38771,N_38893);
and U39379 (N_39379,N_38060,N_38948);
nand U39380 (N_39380,N_38591,N_38973);
or U39381 (N_39381,N_38678,N_38493);
and U39382 (N_39382,N_38402,N_38166);
nor U39383 (N_39383,N_38094,N_38989);
and U39384 (N_39384,N_38136,N_38059);
xnor U39385 (N_39385,N_38177,N_38320);
or U39386 (N_39386,N_38804,N_38463);
or U39387 (N_39387,N_38213,N_38433);
xor U39388 (N_39388,N_38702,N_38826);
or U39389 (N_39389,N_38752,N_38875);
nand U39390 (N_39390,N_38536,N_38092);
or U39391 (N_39391,N_38108,N_38464);
or U39392 (N_39392,N_38137,N_38335);
nor U39393 (N_39393,N_38345,N_38288);
nor U39394 (N_39394,N_38941,N_38070);
xnor U39395 (N_39395,N_38294,N_38764);
nor U39396 (N_39396,N_38869,N_38628);
nand U39397 (N_39397,N_38840,N_38293);
nand U39398 (N_39398,N_38062,N_38119);
nand U39399 (N_39399,N_38580,N_38977);
nor U39400 (N_39400,N_38451,N_38314);
and U39401 (N_39401,N_38913,N_38212);
xor U39402 (N_39402,N_38436,N_38282);
xnor U39403 (N_39403,N_38876,N_38065);
nand U39404 (N_39404,N_38263,N_38834);
nand U39405 (N_39405,N_38210,N_38655);
xnor U39406 (N_39406,N_38163,N_38800);
or U39407 (N_39407,N_38657,N_38047);
nor U39408 (N_39408,N_38206,N_38981);
nand U39409 (N_39409,N_38401,N_38202);
xor U39410 (N_39410,N_38995,N_38127);
and U39411 (N_39411,N_38441,N_38007);
and U39412 (N_39412,N_38581,N_38032);
nand U39413 (N_39413,N_38148,N_38579);
nand U39414 (N_39414,N_38328,N_38956);
nand U39415 (N_39415,N_38365,N_38199);
or U39416 (N_39416,N_38045,N_38082);
xor U39417 (N_39417,N_38461,N_38124);
or U39418 (N_39418,N_38349,N_38921);
and U39419 (N_39419,N_38623,N_38230);
or U39420 (N_39420,N_38184,N_38807);
nand U39421 (N_39421,N_38474,N_38952);
or U39422 (N_39422,N_38988,N_38982);
nor U39423 (N_39423,N_38927,N_38208);
nor U39424 (N_39424,N_38424,N_38151);
and U39425 (N_39425,N_38452,N_38440);
xor U39426 (N_39426,N_38183,N_38422);
nand U39427 (N_39427,N_38968,N_38133);
nand U39428 (N_39428,N_38639,N_38271);
and U39429 (N_39429,N_38331,N_38802);
and U39430 (N_39430,N_38078,N_38369);
or U39431 (N_39431,N_38445,N_38842);
nor U39432 (N_39432,N_38964,N_38994);
xnor U39433 (N_39433,N_38785,N_38466);
and U39434 (N_39434,N_38829,N_38850);
nand U39435 (N_39435,N_38086,N_38022);
nor U39436 (N_39436,N_38630,N_38398);
xnor U39437 (N_39437,N_38889,N_38951);
or U39438 (N_39438,N_38667,N_38997);
or U39439 (N_39439,N_38249,N_38609);
or U39440 (N_39440,N_38554,N_38697);
or U39441 (N_39441,N_38478,N_38429);
or U39442 (N_39442,N_38812,N_38522);
nand U39443 (N_39443,N_38943,N_38665);
nor U39444 (N_39444,N_38675,N_38303);
nor U39445 (N_39445,N_38841,N_38279);
nor U39446 (N_39446,N_38843,N_38196);
nor U39447 (N_39447,N_38496,N_38437);
xor U39448 (N_39448,N_38428,N_38448);
nor U39449 (N_39449,N_38792,N_38013);
nand U39450 (N_39450,N_38518,N_38795);
and U39451 (N_39451,N_38514,N_38637);
and U39452 (N_39452,N_38347,N_38805);
nand U39453 (N_39453,N_38309,N_38914);
xnor U39454 (N_39454,N_38766,N_38736);
and U39455 (N_39455,N_38237,N_38553);
and U39456 (N_39456,N_38879,N_38777);
nor U39457 (N_39457,N_38415,N_38413);
or U39458 (N_39458,N_38549,N_38692);
nand U39459 (N_39459,N_38266,N_38900);
and U39460 (N_39460,N_38642,N_38026);
xnor U39461 (N_39461,N_38469,N_38201);
nand U39462 (N_39462,N_38661,N_38868);
and U39463 (N_39463,N_38543,N_38432);
and U39464 (N_39464,N_38525,N_38749);
and U39465 (N_39465,N_38907,N_38530);
or U39466 (N_39466,N_38612,N_38141);
and U39467 (N_39467,N_38100,N_38339);
nand U39468 (N_39468,N_38902,N_38924);
xor U39469 (N_39469,N_38755,N_38003);
and U39470 (N_39470,N_38245,N_38281);
nor U39471 (N_39471,N_38976,N_38361);
or U39472 (N_39472,N_38679,N_38354);
nand U39473 (N_39473,N_38222,N_38737);
or U39474 (N_39474,N_38574,N_38946);
nand U39475 (N_39475,N_38008,N_38552);
nor U39476 (N_39476,N_38918,N_38686);
xnor U39477 (N_39477,N_38028,N_38277);
nor U39478 (N_39478,N_38458,N_38193);
or U39479 (N_39479,N_38189,N_38473);
xor U39480 (N_39480,N_38456,N_38323);
xor U39481 (N_39481,N_38985,N_38106);
xor U39482 (N_39482,N_38836,N_38408);
and U39483 (N_39483,N_38076,N_38302);
nand U39484 (N_39484,N_38211,N_38381);
nor U39485 (N_39485,N_38129,N_38181);
or U39486 (N_39486,N_38823,N_38015);
xnor U39487 (N_39487,N_38618,N_38584);
nor U39488 (N_39488,N_38351,N_38139);
and U39489 (N_39489,N_38449,N_38001);
nand U39490 (N_39490,N_38715,N_38756);
nand U39491 (N_39491,N_38430,N_38272);
and U39492 (N_39492,N_38370,N_38431);
xor U39493 (N_39493,N_38152,N_38890);
or U39494 (N_39494,N_38776,N_38643);
nand U39495 (N_39495,N_38399,N_38296);
nand U39496 (N_39496,N_38962,N_38699);
nand U39497 (N_39497,N_38341,N_38278);
and U39498 (N_39498,N_38926,N_38300);
or U39499 (N_39499,N_38933,N_38814);
nor U39500 (N_39500,N_38263,N_38671);
xnor U39501 (N_39501,N_38587,N_38525);
xnor U39502 (N_39502,N_38670,N_38403);
nand U39503 (N_39503,N_38101,N_38817);
nor U39504 (N_39504,N_38019,N_38826);
and U39505 (N_39505,N_38458,N_38777);
and U39506 (N_39506,N_38441,N_38332);
xnor U39507 (N_39507,N_38735,N_38463);
and U39508 (N_39508,N_38942,N_38707);
xnor U39509 (N_39509,N_38727,N_38349);
nor U39510 (N_39510,N_38227,N_38771);
or U39511 (N_39511,N_38768,N_38368);
nand U39512 (N_39512,N_38644,N_38809);
or U39513 (N_39513,N_38059,N_38252);
nand U39514 (N_39514,N_38638,N_38796);
or U39515 (N_39515,N_38332,N_38780);
xnor U39516 (N_39516,N_38132,N_38184);
or U39517 (N_39517,N_38329,N_38960);
nor U39518 (N_39518,N_38282,N_38593);
nor U39519 (N_39519,N_38337,N_38986);
or U39520 (N_39520,N_38859,N_38491);
nor U39521 (N_39521,N_38024,N_38261);
nand U39522 (N_39522,N_38809,N_38819);
and U39523 (N_39523,N_38342,N_38823);
or U39524 (N_39524,N_38623,N_38797);
nor U39525 (N_39525,N_38157,N_38209);
nand U39526 (N_39526,N_38021,N_38715);
xnor U39527 (N_39527,N_38251,N_38228);
and U39528 (N_39528,N_38415,N_38760);
nor U39529 (N_39529,N_38356,N_38374);
nor U39530 (N_39530,N_38350,N_38751);
xor U39531 (N_39531,N_38074,N_38187);
xor U39532 (N_39532,N_38710,N_38716);
nand U39533 (N_39533,N_38561,N_38984);
and U39534 (N_39534,N_38536,N_38125);
xor U39535 (N_39535,N_38233,N_38127);
xor U39536 (N_39536,N_38696,N_38381);
or U39537 (N_39537,N_38780,N_38744);
nand U39538 (N_39538,N_38913,N_38242);
or U39539 (N_39539,N_38195,N_38780);
nand U39540 (N_39540,N_38837,N_38926);
nand U39541 (N_39541,N_38575,N_38639);
and U39542 (N_39542,N_38844,N_38916);
and U39543 (N_39543,N_38651,N_38224);
or U39544 (N_39544,N_38324,N_38266);
and U39545 (N_39545,N_38227,N_38907);
and U39546 (N_39546,N_38492,N_38953);
and U39547 (N_39547,N_38547,N_38246);
nor U39548 (N_39548,N_38549,N_38388);
nand U39549 (N_39549,N_38456,N_38011);
or U39550 (N_39550,N_38646,N_38793);
and U39551 (N_39551,N_38310,N_38318);
and U39552 (N_39552,N_38075,N_38944);
or U39553 (N_39553,N_38861,N_38853);
nor U39554 (N_39554,N_38640,N_38471);
or U39555 (N_39555,N_38417,N_38755);
nor U39556 (N_39556,N_38450,N_38066);
and U39557 (N_39557,N_38729,N_38595);
nand U39558 (N_39558,N_38277,N_38529);
xnor U39559 (N_39559,N_38076,N_38383);
and U39560 (N_39560,N_38571,N_38294);
nand U39561 (N_39561,N_38823,N_38769);
nor U39562 (N_39562,N_38328,N_38197);
nand U39563 (N_39563,N_38659,N_38353);
or U39564 (N_39564,N_38629,N_38650);
or U39565 (N_39565,N_38307,N_38245);
nand U39566 (N_39566,N_38456,N_38918);
and U39567 (N_39567,N_38757,N_38201);
and U39568 (N_39568,N_38698,N_38502);
nor U39569 (N_39569,N_38115,N_38426);
or U39570 (N_39570,N_38780,N_38897);
nand U39571 (N_39571,N_38832,N_38639);
nor U39572 (N_39572,N_38196,N_38665);
and U39573 (N_39573,N_38127,N_38040);
and U39574 (N_39574,N_38738,N_38695);
xnor U39575 (N_39575,N_38814,N_38896);
xor U39576 (N_39576,N_38305,N_38799);
or U39577 (N_39577,N_38571,N_38739);
nor U39578 (N_39578,N_38973,N_38665);
nor U39579 (N_39579,N_38037,N_38308);
nand U39580 (N_39580,N_38784,N_38462);
xnor U39581 (N_39581,N_38579,N_38904);
nand U39582 (N_39582,N_38951,N_38885);
xnor U39583 (N_39583,N_38327,N_38453);
and U39584 (N_39584,N_38394,N_38756);
xnor U39585 (N_39585,N_38935,N_38981);
xnor U39586 (N_39586,N_38424,N_38857);
and U39587 (N_39587,N_38670,N_38837);
nand U39588 (N_39588,N_38024,N_38566);
nor U39589 (N_39589,N_38395,N_38964);
and U39590 (N_39590,N_38145,N_38041);
or U39591 (N_39591,N_38403,N_38496);
xnor U39592 (N_39592,N_38091,N_38359);
nor U39593 (N_39593,N_38207,N_38386);
nand U39594 (N_39594,N_38747,N_38710);
nand U39595 (N_39595,N_38376,N_38150);
and U39596 (N_39596,N_38964,N_38168);
nor U39597 (N_39597,N_38326,N_38151);
or U39598 (N_39598,N_38759,N_38180);
or U39599 (N_39599,N_38173,N_38702);
nand U39600 (N_39600,N_38312,N_38321);
xor U39601 (N_39601,N_38550,N_38199);
xor U39602 (N_39602,N_38352,N_38741);
xor U39603 (N_39603,N_38276,N_38311);
xor U39604 (N_39604,N_38337,N_38108);
xor U39605 (N_39605,N_38548,N_38391);
xor U39606 (N_39606,N_38855,N_38140);
or U39607 (N_39607,N_38379,N_38703);
or U39608 (N_39608,N_38745,N_38430);
xor U39609 (N_39609,N_38536,N_38754);
or U39610 (N_39610,N_38532,N_38255);
and U39611 (N_39611,N_38182,N_38788);
nand U39612 (N_39612,N_38984,N_38350);
nor U39613 (N_39613,N_38338,N_38372);
nor U39614 (N_39614,N_38300,N_38254);
xnor U39615 (N_39615,N_38659,N_38942);
nand U39616 (N_39616,N_38404,N_38261);
nor U39617 (N_39617,N_38615,N_38472);
and U39618 (N_39618,N_38937,N_38263);
or U39619 (N_39619,N_38966,N_38884);
and U39620 (N_39620,N_38371,N_38094);
and U39621 (N_39621,N_38223,N_38087);
and U39622 (N_39622,N_38094,N_38213);
nor U39623 (N_39623,N_38733,N_38393);
xnor U39624 (N_39624,N_38806,N_38547);
and U39625 (N_39625,N_38692,N_38481);
xor U39626 (N_39626,N_38967,N_38797);
or U39627 (N_39627,N_38983,N_38872);
or U39628 (N_39628,N_38369,N_38124);
nand U39629 (N_39629,N_38850,N_38338);
and U39630 (N_39630,N_38446,N_38767);
nor U39631 (N_39631,N_38951,N_38595);
nor U39632 (N_39632,N_38372,N_38476);
and U39633 (N_39633,N_38876,N_38091);
nand U39634 (N_39634,N_38787,N_38941);
nor U39635 (N_39635,N_38884,N_38071);
xor U39636 (N_39636,N_38148,N_38209);
nor U39637 (N_39637,N_38092,N_38309);
nand U39638 (N_39638,N_38805,N_38190);
and U39639 (N_39639,N_38117,N_38213);
or U39640 (N_39640,N_38805,N_38754);
xnor U39641 (N_39641,N_38782,N_38968);
xnor U39642 (N_39642,N_38253,N_38372);
and U39643 (N_39643,N_38034,N_38574);
xor U39644 (N_39644,N_38103,N_38520);
nor U39645 (N_39645,N_38578,N_38819);
nand U39646 (N_39646,N_38422,N_38521);
or U39647 (N_39647,N_38537,N_38513);
nor U39648 (N_39648,N_38674,N_38711);
nor U39649 (N_39649,N_38105,N_38603);
and U39650 (N_39650,N_38533,N_38694);
xor U39651 (N_39651,N_38417,N_38692);
nor U39652 (N_39652,N_38310,N_38557);
and U39653 (N_39653,N_38458,N_38985);
or U39654 (N_39654,N_38448,N_38810);
and U39655 (N_39655,N_38829,N_38345);
xnor U39656 (N_39656,N_38237,N_38563);
nand U39657 (N_39657,N_38807,N_38695);
and U39658 (N_39658,N_38439,N_38368);
nor U39659 (N_39659,N_38288,N_38594);
and U39660 (N_39660,N_38266,N_38389);
nand U39661 (N_39661,N_38285,N_38048);
nand U39662 (N_39662,N_38797,N_38813);
or U39663 (N_39663,N_38187,N_38370);
or U39664 (N_39664,N_38965,N_38921);
nor U39665 (N_39665,N_38993,N_38705);
xor U39666 (N_39666,N_38776,N_38989);
or U39667 (N_39667,N_38290,N_38982);
and U39668 (N_39668,N_38504,N_38921);
and U39669 (N_39669,N_38498,N_38309);
and U39670 (N_39670,N_38020,N_38028);
nand U39671 (N_39671,N_38922,N_38219);
nor U39672 (N_39672,N_38019,N_38627);
nand U39673 (N_39673,N_38714,N_38983);
nand U39674 (N_39674,N_38002,N_38427);
nor U39675 (N_39675,N_38161,N_38772);
nor U39676 (N_39676,N_38615,N_38775);
xnor U39677 (N_39677,N_38519,N_38549);
and U39678 (N_39678,N_38126,N_38255);
nor U39679 (N_39679,N_38106,N_38474);
xor U39680 (N_39680,N_38210,N_38311);
or U39681 (N_39681,N_38701,N_38868);
and U39682 (N_39682,N_38050,N_38225);
nand U39683 (N_39683,N_38573,N_38669);
and U39684 (N_39684,N_38880,N_38640);
or U39685 (N_39685,N_38453,N_38962);
and U39686 (N_39686,N_38261,N_38784);
nor U39687 (N_39687,N_38772,N_38282);
and U39688 (N_39688,N_38620,N_38856);
and U39689 (N_39689,N_38534,N_38375);
nand U39690 (N_39690,N_38387,N_38928);
or U39691 (N_39691,N_38205,N_38979);
xnor U39692 (N_39692,N_38170,N_38108);
or U39693 (N_39693,N_38245,N_38035);
and U39694 (N_39694,N_38916,N_38047);
nor U39695 (N_39695,N_38665,N_38506);
nor U39696 (N_39696,N_38680,N_38591);
nand U39697 (N_39697,N_38822,N_38195);
and U39698 (N_39698,N_38487,N_38196);
nor U39699 (N_39699,N_38017,N_38925);
xnor U39700 (N_39700,N_38111,N_38616);
and U39701 (N_39701,N_38965,N_38526);
xor U39702 (N_39702,N_38776,N_38613);
nor U39703 (N_39703,N_38962,N_38927);
nor U39704 (N_39704,N_38420,N_38292);
nor U39705 (N_39705,N_38007,N_38244);
or U39706 (N_39706,N_38172,N_38041);
nand U39707 (N_39707,N_38457,N_38301);
nor U39708 (N_39708,N_38853,N_38264);
xnor U39709 (N_39709,N_38169,N_38492);
or U39710 (N_39710,N_38263,N_38293);
or U39711 (N_39711,N_38577,N_38432);
xor U39712 (N_39712,N_38352,N_38592);
nor U39713 (N_39713,N_38746,N_38541);
nor U39714 (N_39714,N_38801,N_38696);
xnor U39715 (N_39715,N_38659,N_38409);
xnor U39716 (N_39716,N_38496,N_38906);
or U39717 (N_39717,N_38202,N_38250);
nand U39718 (N_39718,N_38378,N_38786);
or U39719 (N_39719,N_38250,N_38261);
xnor U39720 (N_39720,N_38336,N_38353);
nor U39721 (N_39721,N_38207,N_38663);
nand U39722 (N_39722,N_38164,N_38565);
nor U39723 (N_39723,N_38834,N_38100);
nor U39724 (N_39724,N_38469,N_38744);
or U39725 (N_39725,N_38781,N_38426);
nor U39726 (N_39726,N_38900,N_38442);
nand U39727 (N_39727,N_38501,N_38191);
and U39728 (N_39728,N_38781,N_38451);
nand U39729 (N_39729,N_38530,N_38272);
and U39730 (N_39730,N_38576,N_38622);
or U39731 (N_39731,N_38323,N_38336);
or U39732 (N_39732,N_38822,N_38909);
nor U39733 (N_39733,N_38201,N_38519);
xnor U39734 (N_39734,N_38545,N_38337);
xnor U39735 (N_39735,N_38407,N_38335);
or U39736 (N_39736,N_38079,N_38262);
xnor U39737 (N_39737,N_38787,N_38717);
xor U39738 (N_39738,N_38337,N_38196);
nand U39739 (N_39739,N_38063,N_38981);
or U39740 (N_39740,N_38767,N_38018);
nor U39741 (N_39741,N_38917,N_38019);
nand U39742 (N_39742,N_38016,N_38620);
or U39743 (N_39743,N_38532,N_38103);
xor U39744 (N_39744,N_38607,N_38380);
nand U39745 (N_39745,N_38168,N_38638);
and U39746 (N_39746,N_38246,N_38073);
and U39747 (N_39747,N_38737,N_38429);
or U39748 (N_39748,N_38113,N_38271);
or U39749 (N_39749,N_38936,N_38718);
nor U39750 (N_39750,N_38391,N_38298);
and U39751 (N_39751,N_38293,N_38453);
xnor U39752 (N_39752,N_38204,N_38980);
xnor U39753 (N_39753,N_38316,N_38861);
nor U39754 (N_39754,N_38855,N_38770);
and U39755 (N_39755,N_38996,N_38222);
and U39756 (N_39756,N_38284,N_38021);
nand U39757 (N_39757,N_38419,N_38926);
xnor U39758 (N_39758,N_38486,N_38380);
or U39759 (N_39759,N_38828,N_38246);
nand U39760 (N_39760,N_38970,N_38656);
and U39761 (N_39761,N_38874,N_38518);
xor U39762 (N_39762,N_38752,N_38854);
or U39763 (N_39763,N_38774,N_38451);
or U39764 (N_39764,N_38532,N_38490);
or U39765 (N_39765,N_38907,N_38868);
nor U39766 (N_39766,N_38657,N_38220);
xor U39767 (N_39767,N_38111,N_38512);
nor U39768 (N_39768,N_38239,N_38048);
or U39769 (N_39769,N_38198,N_38381);
or U39770 (N_39770,N_38393,N_38382);
or U39771 (N_39771,N_38185,N_38871);
nand U39772 (N_39772,N_38949,N_38703);
or U39773 (N_39773,N_38281,N_38950);
nand U39774 (N_39774,N_38759,N_38091);
xor U39775 (N_39775,N_38280,N_38344);
xor U39776 (N_39776,N_38293,N_38580);
nor U39777 (N_39777,N_38097,N_38495);
xnor U39778 (N_39778,N_38956,N_38020);
nand U39779 (N_39779,N_38570,N_38603);
nand U39780 (N_39780,N_38626,N_38830);
or U39781 (N_39781,N_38108,N_38687);
xor U39782 (N_39782,N_38436,N_38441);
or U39783 (N_39783,N_38983,N_38448);
xor U39784 (N_39784,N_38099,N_38880);
nor U39785 (N_39785,N_38855,N_38669);
nand U39786 (N_39786,N_38396,N_38587);
xor U39787 (N_39787,N_38695,N_38863);
and U39788 (N_39788,N_38813,N_38347);
nor U39789 (N_39789,N_38446,N_38308);
and U39790 (N_39790,N_38282,N_38638);
or U39791 (N_39791,N_38535,N_38807);
nand U39792 (N_39792,N_38153,N_38197);
or U39793 (N_39793,N_38494,N_38333);
nor U39794 (N_39794,N_38410,N_38808);
or U39795 (N_39795,N_38354,N_38745);
xnor U39796 (N_39796,N_38864,N_38851);
or U39797 (N_39797,N_38466,N_38203);
or U39798 (N_39798,N_38745,N_38240);
xnor U39799 (N_39799,N_38627,N_38870);
and U39800 (N_39800,N_38478,N_38441);
nor U39801 (N_39801,N_38058,N_38518);
nand U39802 (N_39802,N_38999,N_38533);
and U39803 (N_39803,N_38175,N_38913);
xnor U39804 (N_39804,N_38056,N_38642);
nand U39805 (N_39805,N_38432,N_38367);
xnor U39806 (N_39806,N_38155,N_38764);
or U39807 (N_39807,N_38512,N_38877);
nand U39808 (N_39808,N_38312,N_38727);
nor U39809 (N_39809,N_38824,N_38933);
xor U39810 (N_39810,N_38148,N_38986);
or U39811 (N_39811,N_38409,N_38312);
xnor U39812 (N_39812,N_38691,N_38591);
and U39813 (N_39813,N_38114,N_38336);
xnor U39814 (N_39814,N_38293,N_38438);
xnor U39815 (N_39815,N_38355,N_38372);
and U39816 (N_39816,N_38249,N_38363);
xor U39817 (N_39817,N_38728,N_38220);
or U39818 (N_39818,N_38974,N_38845);
or U39819 (N_39819,N_38652,N_38191);
and U39820 (N_39820,N_38923,N_38673);
and U39821 (N_39821,N_38943,N_38541);
nor U39822 (N_39822,N_38097,N_38926);
and U39823 (N_39823,N_38050,N_38415);
or U39824 (N_39824,N_38292,N_38867);
nor U39825 (N_39825,N_38715,N_38952);
xnor U39826 (N_39826,N_38596,N_38696);
nor U39827 (N_39827,N_38706,N_38549);
xor U39828 (N_39828,N_38784,N_38779);
or U39829 (N_39829,N_38510,N_38240);
nand U39830 (N_39830,N_38967,N_38986);
or U39831 (N_39831,N_38553,N_38179);
nor U39832 (N_39832,N_38040,N_38065);
nand U39833 (N_39833,N_38447,N_38429);
nand U39834 (N_39834,N_38879,N_38546);
nand U39835 (N_39835,N_38239,N_38126);
nor U39836 (N_39836,N_38399,N_38805);
xnor U39837 (N_39837,N_38981,N_38751);
and U39838 (N_39838,N_38571,N_38062);
or U39839 (N_39839,N_38681,N_38791);
xor U39840 (N_39840,N_38188,N_38580);
or U39841 (N_39841,N_38659,N_38651);
and U39842 (N_39842,N_38428,N_38324);
xor U39843 (N_39843,N_38545,N_38668);
nand U39844 (N_39844,N_38027,N_38817);
and U39845 (N_39845,N_38220,N_38498);
and U39846 (N_39846,N_38838,N_38902);
xor U39847 (N_39847,N_38038,N_38271);
and U39848 (N_39848,N_38806,N_38117);
or U39849 (N_39849,N_38895,N_38214);
and U39850 (N_39850,N_38980,N_38822);
xnor U39851 (N_39851,N_38246,N_38724);
xor U39852 (N_39852,N_38231,N_38766);
xor U39853 (N_39853,N_38477,N_38373);
or U39854 (N_39854,N_38810,N_38406);
nor U39855 (N_39855,N_38471,N_38666);
or U39856 (N_39856,N_38926,N_38663);
or U39857 (N_39857,N_38140,N_38076);
xor U39858 (N_39858,N_38678,N_38343);
xnor U39859 (N_39859,N_38195,N_38956);
or U39860 (N_39860,N_38630,N_38980);
or U39861 (N_39861,N_38902,N_38998);
or U39862 (N_39862,N_38072,N_38412);
or U39863 (N_39863,N_38303,N_38369);
xor U39864 (N_39864,N_38382,N_38169);
and U39865 (N_39865,N_38633,N_38603);
or U39866 (N_39866,N_38429,N_38138);
nand U39867 (N_39867,N_38033,N_38684);
and U39868 (N_39868,N_38438,N_38708);
nand U39869 (N_39869,N_38783,N_38940);
or U39870 (N_39870,N_38559,N_38909);
nor U39871 (N_39871,N_38626,N_38739);
xor U39872 (N_39872,N_38432,N_38967);
xnor U39873 (N_39873,N_38713,N_38595);
nand U39874 (N_39874,N_38529,N_38208);
or U39875 (N_39875,N_38503,N_38340);
nand U39876 (N_39876,N_38522,N_38204);
and U39877 (N_39877,N_38308,N_38953);
or U39878 (N_39878,N_38653,N_38268);
and U39879 (N_39879,N_38264,N_38985);
nor U39880 (N_39880,N_38908,N_38584);
xor U39881 (N_39881,N_38240,N_38962);
nor U39882 (N_39882,N_38340,N_38069);
and U39883 (N_39883,N_38962,N_38086);
or U39884 (N_39884,N_38168,N_38461);
nor U39885 (N_39885,N_38605,N_38332);
and U39886 (N_39886,N_38367,N_38400);
xnor U39887 (N_39887,N_38639,N_38835);
nor U39888 (N_39888,N_38038,N_38222);
nand U39889 (N_39889,N_38306,N_38571);
and U39890 (N_39890,N_38974,N_38255);
or U39891 (N_39891,N_38121,N_38706);
nor U39892 (N_39892,N_38349,N_38586);
and U39893 (N_39893,N_38503,N_38770);
nand U39894 (N_39894,N_38062,N_38510);
nor U39895 (N_39895,N_38060,N_38918);
and U39896 (N_39896,N_38857,N_38431);
nor U39897 (N_39897,N_38022,N_38554);
or U39898 (N_39898,N_38772,N_38666);
xnor U39899 (N_39899,N_38592,N_38518);
or U39900 (N_39900,N_38167,N_38625);
nand U39901 (N_39901,N_38738,N_38648);
nand U39902 (N_39902,N_38612,N_38999);
nand U39903 (N_39903,N_38700,N_38207);
nor U39904 (N_39904,N_38640,N_38491);
nand U39905 (N_39905,N_38401,N_38565);
nand U39906 (N_39906,N_38820,N_38211);
or U39907 (N_39907,N_38558,N_38690);
nand U39908 (N_39908,N_38781,N_38259);
or U39909 (N_39909,N_38949,N_38750);
xor U39910 (N_39910,N_38248,N_38452);
xor U39911 (N_39911,N_38862,N_38833);
and U39912 (N_39912,N_38580,N_38366);
and U39913 (N_39913,N_38081,N_38564);
xnor U39914 (N_39914,N_38644,N_38355);
or U39915 (N_39915,N_38677,N_38671);
and U39916 (N_39916,N_38507,N_38868);
xnor U39917 (N_39917,N_38966,N_38095);
nand U39918 (N_39918,N_38731,N_38523);
or U39919 (N_39919,N_38815,N_38978);
and U39920 (N_39920,N_38167,N_38421);
xor U39921 (N_39921,N_38480,N_38042);
xnor U39922 (N_39922,N_38555,N_38975);
or U39923 (N_39923,N_38432,N_38359);
xor U39924 (N_39924,N_38547,N_38302);
or U39925 (N_39925,N_38014,N_38817);
nand U39926 (N_39926,N_38099,N_38142);
xnor U39927 (N_39927,N_38131,N_38342);
nor U39928 (N_39928,N_38816,N_38555);
nor U39929 (N_39929,N_38931,N_38532);
xor U39930 (N_39930,N_38637,N_38967);
nor U39931 (N_39931,N_38942,N_38679);
xor U39932 (N_39932,N_38051,N_38799);
xor U39933 (N_39933,N_38515,N_38450);
nand U39934 (N_39934,N_38875,N_38888);
xnor U39935 (N_39935,N_38444,N_38079);
nand U39936 (N_39936,N_38016,N_38998);
nand U39937 (N_39937,N_38982,N_38207);
and U39938 (N_39938,N_38056,N_38265);
and U39939 (N_39939,N_38029,N_38607);
and U39940 (N_39940,N_38367,N_38407);
or U39941 (N_39941,N_38651,N_38571);
xor U39942 (N_39942,N_38478,N_38909);
xor U39943 (N_39943,N_38278,N_38989);
nand U39944 (N_39944,N_38044,N_38815);
and U39945 (N_39945,N_38545,N_38498);
nand U39946 (N_39946,N_38605,N_38049);
xor U39947 (N_39947,N_38339,N_38956);
xnor U39948 (N_39948,N_38301,N_38017);
or U39949 (N_39949,N_38730,N_38338);
or U39950 (N_39950,N_38147,N_38997);
or U39951 (N_39951,N_38413,N_38924);
nor U39952 (N_39952,N_38058,N_38375);
nor U39953 (N_39953,N_38784,N_38486);
nor U39954 (N_39954,N_38967,N_38735);
nand U39955 (N_39955,N_38553,N_38400);
xnor U39956 (N_39956,N_38533,N_38592);
and U39957 (N_39957,N_38773,N_38035);
and U39958 (N_39958,N_38870,N_38720);
nand U39959 (N_39959,N_38712,N_38921);
xor U39960 (N_39960,N_38967,N_38563);
nor U39961 (N_39961,N_38805,N_38075);
xor U39962 (N_39962,N_38135,N_38052);
xor U39963 (N_39963,N_38335,N_38195);
and U39964 (N_39964,N_38268,N_38905);
or U39965 (N_39965,N_38470,N_38286);
and U39966 (N_39966,N_38532,N_38847);
nand U39967 (N_39967,N_38167,N_38728);
nor U39968 (N_39968,N_38106,N_38294);
or U39969 (N_39969,N_38101,N_38493);
or U39970 (N_39970,N_38134,N_38268);
nand U39971 (N_39971,N_38018,N_38607);
xor U39972 (N_39972,N_38547,N_38403);
and U39973 (N_39973,N_38194,N_38660);
and U39974 (N_39974,N_38822,N_38121);
nor U39975 (N_39975,N_38307,N_38686);
xor U39976 (N_39976,N_38837,N_38288);
nand U39977 (N_39977,N_38060,N_38935);
and U39978 (N_39978,N_38555,N_38381);
or U39979 (N_39979,N_38484,N_38709);
xor U39980 (N_39980,N_38269,N_38209);
or U39981 (N_39981,N_38894,N_38051);
nor U39982 (N_39982,N_38969,N_38714);
nor U39983 (N_39983,N_38348,N_38251);
and U39984 (N_39984,N_38095,N_38094);
and U39985 (N_39985,N_38062,N_38698);
nand U39986 (N_39986,N_38425,N_38788);
nand U39987 (N_39987,N_38069,N_38581);
xor U39988 (N_39988,N_38486,N_38517);
nand U39989 (N_39989,N_38470,N_38166);
xor U39990 (N_39990,N_38208,N_38908);
or U39991 (N_39991,N_38086,N_38959);
and U39992 (N_39992,N_38168,N_38264);
nor U39993 (N_39993,N_38391,N_38024);
xor U39994 (N_39994,N_38488,N_38314);
xnor U39995 (N_39995,N_38825,N_38413);
nor U39996 (N_39996,N_38535,N_38643);
nand U39997 (N_39997,N_38850,N_38017);
xnor U39998 (N_39998,N_38918,N_38541);
nor U39999 (N_39999,N_38485,N_38204);
and U40000 (N_40000,N_39542,N_39940);
and U40001 (N_40001,N_39789,N_39502);
or U40002 (N_40002,N_39939,N_39090);
xor U40003 (N_40003,N_39345,N_39161);
nor U40004 (N_40004,N_39109,N_39145);
nand U40005 (N_40005,N_39653,N_39120);
and U40006 (N_40006,N_39630,N_39261);
or U40007 (N_40007,N_39840,N_39674);
nor U40008 (N_40008,N_39773,N_39903);
nor U40009 (N_40009,N_39995,N_39246);
nand U40010 (N_40010,N_39131,N_39938);
and U40011 (N_40011,N_39990,N_39069);
xnor U40012 (N_40012,N_39479,N_39035);
or U40013 (N_40013,N_39066,N_39176);
or U40014 (N_40014,N_39981,N_39805);
nor U40015 (N_40015,N_39321,N_39920);
xor U40016 (N_40016,N_39156,N_39974);
xnor U40017 (N_40017,N_39948,N_39216);
nor U40018 (N_40018,N_39725,N_39856);
nand U40019 (N_40019,N_39271,N_39633);
or U40020 (N_40020,N_39683,N_39512);
or U40021 (N_40021,N_39579,N_39217);
xor U40022 (N_40022,N_39941,N_39178);
or U40023 (N_40023,N_39332,N_39115);
and U40024 (N_40024,N_39590,N_39010);
nand U40025 (N_40025,N_39838,N_39614);
or U40026 (N_40026,N_39053,N_39736);
xnor U40027 (N_40027,N_39196,N_39097);
or U40028 (N_40028,N_39154,N_39572);
xnor U40029 (N_40029,N_39235,N_39787);
nand U40030 (N_40030,N_39365,N_39682);
nand U40031 (N_40031,N_39786,N_39025);
and U40032 (N_40032,N_39622,N_39909);
nand U40033 (N_40033,N_39484,N_39922);
or U40034 (N_40034,N_39804,N_39781);
nand U40035 (N_40035,N_39983,N_39259);
xor U40036 (N_40036,N_39467,N_39262);
nor U40037 (N_40037,N_39244,N_39518);
or U40038 (N_40038,N_39666,N_39000);
nor U40039 (N_40039,N_39458,N_39863);
nor U40040 (N_40040,N_39075,N_39972);
xnor U40041 (N_40041,N_39900,N_39629);
nor U40042 (N_40042,N_39135,N_39390);
nand U40043 (N_40043,N_39207,N_39347);
or U40044 (N_40044,N_39383,N_39762);
and U40045 (N_40045,N_39334,N_39959);
and U40046 (N_40046,N_39788,N_39628);
and U40047 (N_40047,N_39558,N_39224);
nor U40048 (N_40048,N_39050,N_39247);
nor U40049 (N_40049,N_39078,N_39330);
and U40050 (N_40050,N_39077,N_39453);
nand U40051 (N_40051,N_39891,N_39521);
nand U40052 (N_40052,N_39464,N_39545);
or U40053 (N_40053,N_39290,N_39327);
nand U40054 (N_40054,N_39204,N_39764);
nand U40055 (N_40055,N_39181,N_39855);
or U40056 (N_40056,N_39094,N_39228);
and U40057 (N_40057,N_39304,N_39954);
or U40058 (N_40058,N_39753,N_39122);
xor U40059 (N_40059,N_39231,N_39236);
and U40060 (N_40060,N_39032,N_39285);
nor U40061 (N_40061,N_39210,N_39192);
nand U40062 (N_40062,N_39401,N_39612);
or U40063 (N_40063,N_39520,N_39733);
nand U40064 (N_40064,N_39564,N_39143);
and U40065 (N_40065,N_39585,N_39607);
nor U40066 (N_40066,N_39643,N_39623);
nor U40067 (N_40067,N_39041,N_39289);
nor U40068 (N_40068,N_39870,N_39960);
xnor U40069 (N_40069,N_39012,N_39867);
xor U40070 (N_40070,N_39408,N_39309);
or U40071 (N_40071,N_39134,N_39428);
or U40072 (N_40072,N_39841,N_39646);
xnor U40073 (N_40073,N_39311,N_39644);
or U40074 (N_40074,N_39926,N_39727);
or U40075 (N_40075,N_39839,N_39076);
nor U40076 (N_40076,N_39242,N_39996);
nor U40077 (N_40077,N_39864,N_39305);
or U40078 (N_40078,N_39673,N_39744);
nor U40079 (N_40079,N_39694,N_39267);
nor U40080 (N_40080,N_39952,N_39544);
nand U40081 (N_40081,N_39515,N_39601);
xor U40082 (N_40082,N_39089,N_39671);
nand U40083 (N_40083,N_39913,N_39800);
and U40084 (N_40084,N_39584,N_39536);
or U40085 (N_40085,N_39606,N_39317);
nor U40086 (N_40086,N_39269,N_39381);
or U40087 (N_40087,N_39424,N_39185);
xor U40088 (N_40088,N_39164,N_39924);
and U40089 (N_40089,N_39306,N_39979);
nand U40090 (N_40090,N_39885,N_39649);
nor U40091 (N_40091,N_39255,N_39582);
or U40092 (N_40092,N_39491,N_39883);
xor U40093 (N_40093,N_39591,N_39895);
nor U40094 (N_40094,N_39240,N_39237);
or U40095 (N_40095,N_39563,N_39626);
and U40096 (N_40096,N_39794,N_39522);
xor U40097 (N_40097,N_39982,N_39052);
nand U40098 (N_40098,N_39608,N_39004);
nor U40099 (N_40099,N_39248,N_39229);
nand U40100 (N_40100,N_39619,N_39046);
or U40101 (N_40101,N_39746,N_39758);
or U40102 (N_40102,N_39524,N_39132);
and U40103 (N_40103,N_39958,N_39659);
nor U40104 (N_40104,N_39929,N_39118);
and U40105 (N_40105,N_39138,N_39947);
xnor U40106 (N_40106,N_39447,N_39557);
nor U40107 (N_40107,N_39897,N_39396);
or U40108 (N_40108,N_39051,N_39356);
or U40109 (N_40109,N_39818,N_39587);
nand U40110 (N_40110,N_39807,N_39421);
nor U40111 (N_40111,N_39548,N_39976);
or U40112 (N_40112,N_39469,N_39160);
and U40113 (N_40113,N_39495,N_39583);
nor U40114 (N_40114,N_39253,N_39632);
and U40115 (N_40115,N_39711,N_39042);
or U40116 (N_40116,N_39657,N_39946);
xnor U40117 (N_40117,N_39905,N_39441);
nor U40118 (N_40118,N_39654,N_39700);
nor U40119 (N_40119,N_39760,N_39373);
nand U40120 (N_40120,N_39136,N_39106);
nor U40121 (N_40121,N_39193,N_39568);
and U40122 (N_40122,N_39021,N_39956);
xnor U40123 (N_40123,N_39037,N_39497);
xor U40124 (N_40124,N_39426,N_39079);
nor U40125 (N_40125,N_39882,N_39346);
nand U40126 (N_40126,N_39281,N_39716);
nor U40127 (N_40127,N_39177,N_39553);
or U40128 (N_40128,N_39690,N_39452);
nand U40129 (N_40129,N_39937,N_39412);
or U40130 (N_40130,N_39470,N_39574);
nand U40131 (N_40131,N_39901,N_39577);
nor U40132 (N_40132,N_39935,N_39696);
nand U40133 (N_40133,N_39481,N_39064);
nor U40134 (N_40134,N_39222,N_39312);
and U40135 (N_40135,N_39057,N_39977);
nand U40136 (N_40136,N_39575,N_39689);
nand U40137 (N_40137,N_39308,N_39962);
nand U40138 (N_40138,N_39351,N_39872);
nand U40139 (N_40139,N_39845,N_39265);
xor U40140 (N_40140,N_39105,N_39985);
or U40141 (N_40141,N_39344,N_39743);
nand U40142 (N_40142,N_39934,N_39123);
and U40143 (N_40143,N_39769,N_39993);
or U40144 (N_40144,N_39742,N_39245);
xnor U40145 (N_40145,N_39496,N_39567);
xor U40146 (N_40146,N_39755,N_39017);
nand U40147 (N_40147,N_39793,N_39436);
or U40148 (N_40148,N_39813,N_39268);
xnor U40149 (N_40149,N_39018,N_39302);
nor U40150 (N_40150,N_39911,N_39752);
nor U40151 (N_40151,N_39029,N_39249);
or U40152 (N_40152,N_39537,N_39892);
nand U40153 (N_40153,N_39338,N_39896);
nor U40154 (N_40154,N_39824,N_39505);
or U40155 (N_40155,N_39218,N_39174);
xnor U40156 (N_40156,N_39811,N_39296);
xor U40157 (N_40157,N_39792,N_39234);
or U40158 (N_40158,N_39765,N_39648);
or U40159 (N_40159,N_39595,N_39006);
nand U40160 (N_40160,N_39779,N_39343);
xor U40161 (N_40161,N_39511,N_39149);
or U40162 (N_40162,N_39377,N_39331);
nor U40163 (N_40163,N_39420,N_39501);
or U40164 (N_40164,N_39631,N_39555);
and U40165 (N_40165,N_39028,N_39251);
and U40166 (N_40166,N_39641,N_39117);
xor U40167 (N_40167,N_39226,N_39637);
xor U40168 (N_40168,N_39039,N_39573);
nand U40169 (N_40169,N_39363,N_39741);
nand U40170 (N_40170,N_39635,N_39551);
and U40171 (N_40171,N_39780,N_39560);
and U40172 (N_40172,N_39385,N_39359);
and U40173 (N_40173,N_39086,N_39093);
nor U40174 (N_40174,N_39307,N_39071);
nor U40175 (N_40175,N_39547,N_39655);
nand U40176 (N_40176,N_39706,N_39499);
and U40177 (N_40177,N_39483,N_39494);
or U40178 (N_40178,N_39975,N_39904);
and U40179 (N_40179,N_39315,N_39023);
or U40180 (N_40180,N_39927,N_39814);
nor U40181 (N_40181,N_39707,N_39702);
xor U40182 (N_40182,N_39239,N_39188);
nor U40183 (N_40183,N_39214,N_39677);
and U40184 (N_40184,N_39451,N_39433);
or U40185 (N_40185,N_39802,N_39594);
or U40186 (N_40186,N_39930,N_39152);
nor U40187 (N_40187,N_39531,N_39823);
xor U40188 (N_40188,N_39367,N_39517);
or U40189 (N_40189,N_39917,N_39737);
nand U40190 (N_40190,N_39316,N_39387);
or U40191 (N_40191,N_39906,N_39774);
xnor U40192 (N_40192,N_39445,N_39507);
nor U40193 (N_40193,N_39527,N_39820);
xnor U40194 (N_40194,N_39953,N_39658);
nor U40195 (N_40195,N_39931,N_39036);
and U40196 (N_40196,N_39205,N_39394);
xnor U40197 (N_40197,N_39328,N_39799);
nor U40198 (N_40198,N_39124,N_39910);
nand U40199 (N_40199,N_39020,N_39144);
or U40200 (N_40200,N_39171,N_39999);
xnor U40201 (N_40201,N_39907,N_39357);
xor U40202 (N_40202,N_39663,N_39335);
nor U40203 (N_40203,N_39809,N_39528);
and U40204 (N_40204,N_39615,N_39301);
nor U40205 (N_40205,N_39513,N_39102);
nor U40206 (N_40206,N_39266,N_39260);
nand U40207 (N_40207,N_39191,N_39008);
or U40208 (N_40208,N_39718,N_39691);
or U40209 (N_40209,N_39202,N_39611);
or U40210 (N_40210,N_39790,N_39912);
or U40211 (N_40211,N_39148,N_39063);
nor U40212 (N_40212,N_39073,N_39704);
or U40213 (N_40213,N_39617,N_39681);
and U40214 (N_40214,N_39352,N_39854);
nand U40215 (N_40215,N_39389,N_39701);
or U40216 (N_40216,N_39678,N_39825);
xnor U40217 (N_40217,N_39766,N_39988);
xor U40218 (N_40218,N_39430,N_39116);
or U40219 (N_40219,N_39961,N_39443);
xnor U40220 (N_40220,N_39158,N_39431);
and U40221 (N_40221,N_39273,N_39139);
or U40222 (N_40222,N_39729,N_39096);
or U40223 (N_40223,N_39044,N_39288);
and U40224 (N_40224,N_39916,N_39853);
and U40225 (N_40225,N_39561,N_39002);
nand U40226 (N_40226,N_39687,N_39293);
nand U40227 (N_40227,N_39830,N_39552);
or U40228 (N_40228,N_39605,N_39759);
and U40229 (N_40229,N_39984,N_39461);
nand U40230 (N_40230,N_39219,N_39169);
and U40231 (N_40231,N_39437,N_39326);
and U40232 (N_40232,N_39535,N_39364);
nand U40233 (N_40233,N_39569,N_39879);
xnor U40234 (N_40234,N_39101,N_39033);
or U40235 (N_40235,N_39889,N_39350);
or U40236 (N_40236,N_39730,N_39429);
nor U40237 (N_40237,N_39446,N_39503);
or U40238 (N_40238,N_39195,N_39936);
and U40239 (N_40239,N_39890,N_39989);
xor U40240 (N_40240,N_39358,N_39460);
or U40241 (N_40241,N_39566,N_39713);
nand U40242 (N_40242,N_39416,N_39850);
and U40243 (N_40243,N_39091,N_39874);
and U40244 (N_40244,N_39014,N_39703);
and U40245 (N_40245,N_39324,N_39360);
or U40246 (N_40246,N_39740,N_39233);
xnor U40247 (N_40247,N_39369,N_39486);
nand U40248 (N_40248,N_39925,N_39844);
or U40249 (N_40249,N_39529,N_39852);
nand U40250 (N_40250,N_39448,N_39969);
nor U40251 (N_40251,N_39717,N_39592);
nand U40252 (N_40252,N_39015,N_39045);
xnor U40253 (N_40253,N_39603,N_39846);
xor U40254 (N_40254,N_39209,N_39963);
nor U40255 (N_40255,N_39337,N_39627);
nand U40256 (N_40256,N_39955,N_39862);
and U40257 (N_40257,N_39581,N_39624);
nand U40258 (N_40258,N_39510,N_39980);
xnor U40259 (N_40259,N_39059,N_39944);
nor U40260 (N_40260,N_39128,N_39411);
or U40261 (N_40261,N_39061,N_39998);
nor U40262 (N_40262,N_39942,N_39320);
or U40263 (N_40263,N_39898,N_39082);
nand U40264 (N_40264,N_39415,N_39048);
nor U40265 (N_40265,N_39213,N_39586);
xor U40266 (N_40266,N_39291,N_39914);
nand U40267 (N_40267,N_39419,N_39843);
xnor U40268 (N_40268,N_39571,N_39992);
and U40269 (N_40269,N_39908,N_39422);
xor U40270 (N_40270,N_39887,N_39991);
xor U40271 (N_40271,N_39761,N_39822);
nand U40272 (N_40272,N_39263,N_39153);
and U40273 (N_40273,N_39857,N_39967);
or U40274 (N_40274,N_39187,N_39466);
xor U40275 (N_40275,N_39899,N_39200);
xor U40276 (N_40276,N_39593,N_39554);
xor U40277 (N_40277,N_39785,N_39815);
nand U40278 (N_40278,N_39757,N_39651);
xor U40279 (N_40279,N_39580,N_39860);
nor U40280 (N_40280,N_39837,N_39489);
nor U40281 (N_40281,N_39866,N_39147);
and U40282 (N_40282,N_39477,N_39523);
or U40283 (N_40283,N_39928,N_39965);
or U40284 (N_40284,N_39264,N_39256);
nor U40285 (N_40285,N_39923,N_39111);
nand U40286 (N_40286,N_39221,N_39405);
nor U40287 (N_40287,N_39054,N_39182);
nor U40288 (N_40288,N_39126,N_39533);
xnor U40289 (N_40289,N_39276,N_39386);
xor U40290 (N_40290,N_39541,N_39709);
or U40291 (N_40291,N_39684,N_39362);
and U40292 (N_40292,N_39693,N_39819);
xor U40293 (N_40293,N_39201,N_39747);
and U40294 (N_40294,N_39970,N_39831);
or U40295 (N_40295,N_39720,N_39013);
nor U40296 (N_40296,N_39414,N_39650);
and U40297 (N_40297,N_39616,N_39672);
or U40298 (N_40298,N_39994,N_39519);
or U40299 (N_40299,N_39026,N_39129);
xor U40300 (N_40300,N_39159,N_39639);
nor U40301 (N_40301,N_39068,N_39966);
xnor U40302 (N_40302,N_39668,N_39859);
xor U40303 (N_40303,N_39664,N_39190);
nand U40304 (N_40304,N_39058,N_39024);
nor U40305 (N_40305,N_39243,N_39763);
nor U40306 (N_40306,N_39220,N_39738);
nand U40307 (N_40307,N_39098,N_39865);
xor U40308 (N_40308,N_39333,N_39697);
nor U40309 (N_40309,N_39642,N_39427);
and U40310 (N_40310,N_39679,N_39768);
nand U40311 (N_40311,N_39721,N_39810);
or U40312 (N_40312,N_39797,N_39669);
nand U40313 (N_40313,N_39816,N_39485);
or U40314 (N_40314,N_39771,N_39978);
or U40315 (N_40315,N_39060,N_39151);
or U40316 (N_40316,N_39016,N_39848);
nand U40317 (N_40317,N_39439,N_39971);
nor U40318 (N_40318,N_39832,N_39157);
nand U40319 (N_40319,N_39348,N_39784);
nand U40320 (N_40320,N_39119,N_39685);
xor U40321 (N_40321,N_39272,N_39215);
nand U40322 (N_40322,N_39254,N_39107);
nand U40323 (N_40323,N_39748,N_39660);
or U40324 (N_40324,N_39777,N_39661);
xor U40325 (N_40325,N_39722,N_39380);
nor U40326 (N_40326,N_39104,N_39735);
nor U40327 (N_40327,N_39776,N_39125);
nand U40328 (N_40328,N_39180,N_39007);
nor U40329 (N_40329,N_39062,N_39835);
nor U40330 (N_40330,N_39951,N_39932);
xnor U40331 (N_40331,N_39406,N_39425);
or U40332 (N_40332,N_39067,N_39791);
nand U40333 (N_40333,N_39886,N_39827);
or U40334 (N_40334,N_39403,N_39183);
and U40335 (N_40335,N_39508,N_39141);
or U40336 (N_40336,N_39699,N_39588);
nand U40337 (N_40337,N_39550,N_39092);
xnor U40338 (N_40338,N_39388,N_39698);
nand U40339 (N_40339,N_39888,N_39705);
nand U40340 (N_40340,N_39110,N_39604);
xor U40341 (N_40341,N_39770,N_39894);
nor U40342 (N_40342,N_39223,N_39487);
or U40343 (N_40343,N_39184,N_39277);
or U40344 (N_40344,N_39796,N_39714);
nor U40345 (N_40345,N_39457,N_39875);
xnor U40346 (N_40346,N_39353,N_39287);
nand U40347 (N_40347,N_39950,N_39084);
nand U40348 (N_40348,N_39478,N_39103);
nand U40349 (N_40349,N_39884,N_39099);
and U40350 (N_40350,N_39756,N_39434);
nand U40351 (N_40351,N_39456,N_39121);
xor U40352 (N_40352,N_39806,N_39278);
and U40353 (N_40353,N_39162,N_39949);
xor U40354 (N_40354,N_39303,N_39801);
xnor U40355 (N_40355,N_39795,N_39313);
and U40356 (N_40356,N_39918,N_39565);
nand U40357 (N_40357,N_39179,N_39284);
or U40358 (N_40358,N_39986,N_39283);
and U40359 (N_40359,N_39475,N_39973);
xnor U40360 (N_40360,N_39462,N_39197);
or U40361 (N_40361,N_39600,N_39166);
xnor U40362 (N_40362,N_39130,N_39645);
xnor U40363 (N_40363,N_39395,N_39500);
xnor U40364 (N_40364,N_39397,N_39150);
and U40365 (N_40365,N_39598,N_39413);
xnor U40366 (N_40366,N_39323,N_39556);
and U40367 (N_40367,N_39675,N_39376);
nor U40368 (N_40368,N_39821,N_39945);
xor U40369 (N_40369,N_39728,N_39878);
and U40370 (N_40370,N_39172,N_39108);
nor U40371 (N_40371,N_39782,N_39921);
or U40372 (N_40372,N_39286,N_39435);
nor U40373 (N_40373,N_39933,N_39578);
xnor U40374 (N_40374,N_39391,N_39371);
or U40375 (N_40375,N_39418,N_39964);
and U40376 (N_40376,N_39379,N_39208);
or U40377 (N_40377,N_39250,N_39167);
or U40378 (N_40378,N_39539,N_39238);
nand U40379 (N_40379,N_39186,N_39056);
and U40380 (N_40380,N_39189,N_39576);
nand U40381 (N_40381,N_39997,N_39410);
or U40382 (N_40382,N_39175,N_39695);
or U40383 (N_40383,N_39772,N_39636);
nor U40384 (N_40384,N_39667,N_39080);
nand U40385 (N_40385,N_39361,N_39597);
and U40386 (N_40386,N_39198,N_39530);
or U40387 (N_40387,N_39423,N_39957);
or U40388 (N_40388,N_39734,N_39402);
nor U40389 (N_40389,N_39043,N_39710);
xnor U40390 (N_40390,N_39532,N_39803);
nand U40391 (N_40391,N_39444,N_39754);
or U40392 (N_40392,N_39609,N_39009);
or U40393 (N_40393,N_39919,N_39506);
xor U40394 (N_40394,N_39270,N_39298);
nand U40395 (N_40395,N_39034,N_39847);
nand U40396 (N_40396,N_39339,N_39168);
and U40397 (N_40397,N_39088,N_39318);
nand U40398 (N_40398,N_39194,N_39493);
nor U40399 (N_40399,N_39055,N_39440);
nor U40400 (N_40400,N_39602,N_39432);
xnor U40401 (N_40401,N_39112,N_39399);
nor U40402 (N_40402,N_39341,N_39274);
or U40403 (N_40403,N_39022,N_39340);
nor U40404 (N_40404,N_39516,N_39449);
nand U40405 (N_40405,N_39232,N_39065);
xnor U40406 (N_40406,N_39375,N_39712);
and U40407 (N_40407,N_39355,N_39817);
and U40408 (N_40408,N_39001,N_39005);
nand U40409 (N_40409,N_39750,N_39670);
or U40410 (N_40410,N_39828,N_39325);
or U40411 (N_40411,N_39534,N_39072);
or U40412 (N_40412,N_39472,N_39459);
xor U40413 (N_40413,N_39027,N_39031);
nand U40414 (N_40414,N_39384,N_39620);
nand U40415 (N_40415,N_39310,N_39538);
or U40416 (N_40416,N_39858,N_39943);
xnor U40417 (N_40417,N_39319,N_39812);
and U40418 (N_40418,N_39030,N_39767);
nor U40419 (N_40419,N_39137,N_39011);
nor U40420 (N_40420,N_39474,N_39442);
xor U40421 (N_40421,N_39127,N_39662);
nand U40422 (N_40422,N_39074,N_39625);
or U40423 (N_40423,N_39211,N_39829);
xnor U40424 (N_40424,N_39775,N_39834);
nor U40425 (N_40425,N_39083,N_39783);
or U40426 (N_40426,N_39146,N_39656);
nor U40427 (N_40427,N_39640,N_39163);
xnor U40428 (N_40428,N_39095,N_39562);
nor U40429 (N_40429,N_39230,N_39724);
nor U40430 (N_40430,N_39299,N_39842);
and U40431 (N_40431,N_39851,N_39665);
and U40432 (N_40432,N_39808,N_39087);
nor U40433 (N_40433,N_39492,N_39599);
nor U40434 (N_40434,N_39374,N_39473);
or U40435 (N_40435,N_39294,N_39400);
or U40436 (N_40436,N_39778,N_39114);
xor U40437 (N_40437,N_39915,N_39173);
nor U40438 (N_40438,N_39468,N_39300);
xor U40439 (N_40439,N_39257,N_39241);
nand U40440 (N_40440,N_39404,N_39732);
or U40441 (N_40441,N_39525,N_39454);
nor U40442 (N_40442,N_39354,N_39490);
and U40443 (N_40443,N_39019,N_39081);
nand U40444 (N_40444,N_39652,N_39417);
nor U40445 (N_40445,N_39745,N_39372);
nor U40446 (N_40446,N_39849,N_39155);
nand U40447 (N_40447,N_39049,N_39570);
and U40448 (N_40448,N_39621,N_39723);
nor U40449 (N_40449,N_39407,N_39543);
nor U40450 (N_40450,N_39589,N_39258);
nand U40451 (N_40451,N_39968,N_39280);
nor U40452 (N_40452,N_39170,N_39199);
or U40453 (N_40453,N_39610,N_39739);
nand U40454 (N_40454,N_39225,N_39861);
or U40455 (N_40455,N_39140,N_39370);
xor U40456 (N_40456,N_39833,N_39336);
nor U40457 (N_40457,N_39368,N_39366);
nor U40458 (N_40458,N_39726,N_39038);
xnor U40459 (N_40459,N_39686,N_39540);
xor U40460 (N_40460,N_39393,N_39692);
xor U40461 (N_40461,N_39549,N_39227);
nor U40462 (N_40462,N_39322,N_39040);
xnor U40463 (N_40463,N_39482,N_39869);
nand U40464 (N_40464,N_39480,N_39613);
nand U40465 (N_40465,N_39476,N_39455);
xnor U40466 (N_40466,N_39871,N_39113);
xor U40467 (N_40467,N_39297,N_39392);
nand U40468 (N_40468,N_39881,N_39731);
nor U40469 (N_40469,N_39295,N_39133);
nor U40470 (N_40470,N_39471,N_39559);
xnor U40471 (N_40471,N_39378,N_39826);
nand U40472 (N_40472,N_39987,N_39047);
nand U40473 (N_40473,N_39546,N_39680);
nor U40474 (N_40474,N_39596,N_39398);
or U40475 (N_40475,N_39876,N_39836);
and U40476 (N_40476,N_39514,N_39409);
or U40477 (N_40477,N_39634,N_39085);
xor U40478 (N_40478,N_39488,N_39450);
nand U40479 (N_40479,N_39498,N_39275);
xnor U40480 (N_40480,N_39206,N_39212);
nand U40481 (N_40481,N_39873,N_39638);
and U40482 (N_40482,N_39751,N_39314);
or U40483 (N_40483,N_39715,N_39003);
nor U40484 (N_40484,N_39880,N_39438);
nand U40485 (N_40485,N_39165,N_39100);
nand U40486 (N_40486,N_39279,N_39382);
nand U40487 (N_40487,N_39509,N_39282);
and U40488 (N_40488,N_39142,N_39465);
nor U40489 (N_40489,N_39893,N_39749);
nand U40490 (N_40490,N_39526,N_39708);
nor U40491 (N_40491,N_39463,N_39676);
and U40492 (N_40492,N_39349,N_39618);
xnor U40493 (N_40493,N_39719,N_39877);
nand U40494 (N_40494,N_39688,N_39070);
or U40495 (N_40495,N_39868,N_39647);
nor U40496 (N_40496,N_39252,N_39329);
or U40497 (N_40497,N_39902,N_39203);
and U40498 (N_40498,N_39798,N_39504);
nor U40499 (N_40499,N_39292,N_39342);
xnor U40500 (N_40500,N_39910,N_39896);
nor U40501 (N_40501,N_39349,N_39249);
xor U40502 (N_40502,N_39129,N_39289);
nor U40503 (N_40503,N_39505,N_39393);
and U40504 (N_40504,N_39511,N_39476);
or U40505 (N_40505,N_39325,N_39517);
or U40506 (N_40506,N_39297,N_39295);
nand U40507 (N_40507,N_39908,N_39560);
xnor U40508 (N_40508,N_39527,N_39884);
xnor U40509 (N_40509,N_39461,N_39301);
and U40510 (N_40510,N_39350,N_39557);
nand U40511 (N_40511,N_39357,N_39318);
nand U40512 (N_40512,N_39530,N_39965);
xnor U40513 (N_40513,N_39673,N_39163);
and U40514 (N_40514,N_39149,N_39460);
or U40515 (N_40515,N_39456,N_39619);
or U40516 (N_40516,N_39570,N_39044);
and U40517 (N_40517,N_39524,N_39417);
and U40518 (N_40518,N_39934,N_39286);
or U40519 (N_40519,N_39465,N_39482);
or U40520 (N_40520,N_39020,N_39329);
nand U40521 (N_40521,N_39854,N_39692);
and U40522 (N_40522,N_39749,N_39676);
nor U40523 (N_40523,N_39821,N_39103);
nand U40524 (N_40524,N_39292,N_39548);
nand U40525 (N_40525,N_39305,N_39612);
nand U40526 (N_40526,N_39768,N_39261);
nand U40527 (N_40527,N_39491,N_39466);
xnor U40528 (N_40528,N_39274,N_39069);
or U40529 (N_40529,N_39856,N_39445);
nor U40530 (N_40530,N_39541,N_39765);
nor U40531 (N_40531,N_39905,N_39906);
nand U40532 (N_40532,N_39656,N_39446);
and U40533 (N_40533,N_39903,N_39749);
nor U40534 (N_40534,N_39826,N_39402);
nor U40535 (N_40535,N_39822,N_39635);
or U40536 (N_40536,N_39516,N_39192);
or U40537 (N_40537,N_39186,N_39078);
xor U40538 (N_40538,N_39969,N_39418);
or U40539 (N_40539,N_39031,N_39733);
xor U40540 (N_40540,N_39363,N_39121);
and U40541 (N_40541,N_39840,N_39666);
and U40542 (N_40542,N_39067,N_39122);
nor U40543 (N_40543,N_39912,N_39418);
xnor U40544 (N_40544,N_39258,N_39683);
nand U40545 (N_40545,N_39031,N_39001);
xnor U40546 (N_40546,N_39659,N_39546);
xor U40547 (N_40547,N_39720,N_39279);
and U40548 (N_40548,N_39169,N_39713);
or U40549 (N_40549,N_39900,N_39395);
or U40550 (N_40550,N_39360,N_39182);
or U40551 (N_40551,N_39197,N_39060);
nand U40552 (N_40552,N_39780,N_39719);
or U40553 (N_40553,N_39394,N_39217);
or U40554 (N_40554,N_39655,N_39121);
nand U40555 (N_40555,N_39636,N_39073);
or U40556 (N_40556,N_39830,N_39740);
and U40557 (N_40557,N_39347,N_39904);
or U40558 (N_40558,N_39809,N_39811);
nand U40559 (N_40559,N_39423,N_39078);
and U40560 (N_40560,N_39962,N_39555);
or U40561 (N_40561,N_39489,N_39442);
nor U40562 (N_40562,N_39660,N_39688);
or U40563 (N_40563,N_39289,N_39799);
nor U40564 (N_40564,N_39013,N_39152);
and U40565 (N_40565,N_39063,N_39636);
xor U40566 (N_40566,N_39287,N_39420);
and U40567 (N_40567,N_39562,N_39536);
or U40568 (N_40568,N_39048,N_39189);
and U40569 (N_40569,N_39656,N_39668);
xnor U40570 (N_40570,N_39847,N_39594);
nor U40571 (N_40571,N_39876,N_39211);
or U40572 (N_40572,N_39708,N_39471);
xnor U40573 (N_40573,N_39413,N_39555);
nand U40574 (N_40574,N_39178,N_39790);
and U40575 (N_40575,N_39356,N_39702);
nand U40576 (N_40576,N_39462,N_39140);
xor U40577 (N_40577,N_39552,N_39174);
or U40578 (N_40578,N_39092,N_39212);
nand U40579 (N_40579,N_39291,N_39707);
nor U40580 (N_40580,N_39302,N_39443);
nor U40581 (N_40581,N_39199,N_39629);
nand U40582 (N_40582,N_39564,N_39226);
or U40583 (N_40583,N_39714,N_39061);
xor U40584 (N_40584,N_39143,N_39544);
nand U40585 (N_40585,N_39063,N_39588);
or U40586 (N_40586,N_39948,N_39592);
xor U40587 (N_40587,N_39374,N_39418);
nor U40588 (N_40588,N_39229,N_39811);
or U40589 (N_40589,N_39895,N_39353);
nand U40590 (N_40590,N_39497,N_39717);
and U40591 (N_40591,N_39213,N_39188);
xnor U40592 (N_40592,N_39863,N_39032);
nand U40593 (N_40593,N_39223,N_39383);
nand U40594 (N_40594,N_39045,N_39334);
or U40595 (N_40595,N_39482,N_39085);
and U40596 (N_40596,N_39174,N_39279);
nand U40597 (N_40597,N_39920,N_39144);
nor U40598 (N_40598,N_39366,N_39627);
or U40599 (N_40599,N_39815,N_39261);
and U40600 (N_40600,N_39768,N_39075);
nand U40601 (N_40601,N_39860,N_39438);
nand U40602 (N_40602,N_39873,N_39448);
or U40603 (N_40603,N_39001,N_39505);
xnor U40604 (N_40604,N_39794,N_39248);
xnor U40605 (N_40605,N_39078,N_39448);
nand U40606 (N_40606,N_39288,N_39119);
nand U40607 (N_40607,N_39718,N_39523);
xor U40608 (N_40608,N_39057,N_39297);
or U40609 (N_40609,N_39882,N_39288);
or U40610 (N_40610,N_39976,N_39869);
and U40611 (N_40611,N_39933,N_39085);
xnor U40612 (N_40612,N_39288,N_39245);
or U40613 (N_40613,N_39208,N_39436);
xor U40614 (N_40614,N_39809,N_39233);
xor U40615 (N_40615,N_39444,N_39250);
xor U40616 (N_40616,N_39446,N_39498);
and U40617 (N_40617,N_39084,N_39291);
xor U40618 (N_40618,N_39045,N_39954);
xnor U40619 (N_40619,N_39402,N_39877);
nor U40620 (N_40620,N_39590,N_39991);
nor U40621 (N_40621,N_39130,N_39997);
or U40622 (N_40622,N_39875,N_39825);
nand U40623 (N_40623,N_39957,N_39863);
or U40624 (N_40624,N_39489,N_39586);
nor U40625 (N_40625,N_39413,N_39404);
nor U40626 (N_40626,N_39029,N_39037);
nand U40627 (N_40627,N_39717,N_39393);
nand U40628 (N_40628,N_39015,N_39215);
or U40629 (N_40629,N_39828,N_39592);
and U40630 (N_40630,N_39601,N_39322);
xnor U40631 (N_40631,N_39891,N_39153);
nand U40632 (N_40632,N_39334,N_39973);
or U40633 (N_40633,N_39486,N_39050);
nand U40634 (N_40634,N_39300,N_39641);
nand U40635 (N_40635,N_39661,N_39197);
nand U40636 (N_40636,N_39670,N_39845);
nand U40637 (N_40637,N_39772,N_39199);
and U40638 (N_40638,N_39269,N_39748);
nand U40639 (N_40639,N_39239,N_39850);
or U40640 (N_40640,N_39851,N_39666);
xnor U40641 (N_40641,N_39111,N_39871);
nor U40642 (N_40642,N_39343,N_39680);
and U40643 (N_40643,N_39051,N_39506);
nor U40644 (N_40644,N_39753,N_39622);
nor U40645 (N_40645,N_39757,N_39642);
nand U40646 (N_40646,N_39115,N_39358);
and U40647 (N_40647,N_39335,N_39938);
nand U40648 (N_40648,N_39000,N_39079);
nor U40649 (N_40649,N_39578,N_39086);
or U40650 (N_40650,N_39634,N_39277);
xor U40651 (N_40651,N_39156,N_39883);
xor U40652 (N_40652,N_39557,N_39800);
xnor U40653 (N_40653,N_39639,N_39874);
and U40654 (N_40654,N_39836,N_39300);
nor U40655 (N_40655,N_39650,N_39623);
nand U40656 (N_40656,N_39831,N_39287);
and U40657 (N_40657,N_39599,N_39531);
xnor U40658 (N_40658,N_39894,N_39742);
nand U40659 (N_40659,N_39291,N_39019);
or U40660 (N_40660,N_39861,N_39830);
or U40661 (N_40661,N_39831,N_39073);
nor U40662 (N_40662,N_39689,N_39499);
nor U40663 (N_40663,N_39988,N_39969);
nand U40664 (N_40664,N_39997,N_39617);
and U40665 (N_40665,N_39813,N_39551);
or U40666 (N_40666,N_39762,N_39015);
xor U40667 (N_40667,N_39754,N_39855);
and U40668 (N_40668,N_39788,N_39204);
and U40669 (N_40669,N_39228,N_39794);
or U40670 (N_40670,N_39906,N_39918);
nor U40671 (N_40671,N_39999,N_39820);
xnor U40672 (N_40672,N_39056,N_39297);
nor U40673 (N_40673,N_39112,N_39703);
nor U40674 (N_40674,N_39892,N_39318);
and U40675 (N_40675,N_39127,N_39031);
and U40676 (N_40676,N_39439,N_39358);
nor U40677 (N_40677,N_39864,N_39166);
or U40678 (N_40678,N_39951,N_39916);
or U40679 (N_40679,N_39029,N_39853);
or U40680 (N_40680,N_39298,N_39474);
and U40681 (N_40681,N_39661,N_39973);
nor U40682 (N_40682,N_39223,N_39832);
nor U40683 (N_40683,N_39435,N_39227);
or U40684 (N_40684,N_39994,N_39546);
nor U40685 (N_40685,N_39937,N_39875);
nand U40686 (N_40686,N_39988,N_39568);
and U40687 (N_40687,N_39608,N_39026);
and U40688 (N_40688,N_39959,N_39693);
and U40689 (N_40689,N_39181,N_39476);
xor U40690 (N_40690,N_39409,N_39431);
xor U40691 (N_40691,N_39813,N_39300);
xnor U40692 (N_40692,N_39351,N_39502);
nor U40693 (N_40693,N_39768,N_39315);
or U40694 (N_40694,N_39511,N_39254);
nand U40695 (N_40695,N_39318,N_39715);
and U40696 (N_40696,N_39520,N_39959);
nor U40697 (N_40697,N_39007,N_39394);
or U40698 (N_40698,N_39201,N_39884);
nand U40699 (N_40699,N_39728,N_39827);
and U40700 (N_40700,N_39548,N_39484);
or U40701 (N_40701,N_39594,N_39515);
nor U40702 (N_40702,N_39123,N_39333);
nand U40703 (N_40703,N_39898,N_39890);
nor U40704 (N_40704,N_39036,N_39942);
xnor U40705 (N_40705,N_39501,N_39634);
xor U40706 (N_40706,N_39291,N_39405);
nand U40707 (N_40707,N_39425,N_39796);
nand U40708 (N_40708,N_39212,N_39476);
or U40709 (N_40709,N_39096,N_39233);
or U40710 (N_40710,N_39532,N_39527);
nand U40711 (N_40711,N_39837,N_39612);
nor U40712 (N_40712,N_39517,N_39894);
nand U40713 (N_40713,N_39895,N_39966);
and U40714 (N_40714,N_39287,N_39876);
or U40715 (N_40715,N_39228,N_39579);
or U40716 (N_40716,N_39123,N_39731);
or U40717 (N_40717,N_39211,N_39744);
or U40718 (N_40718,N_39158,N_39913);
or U40719 (N_40719,N_39151,N_39303);
or U40720 (N_40720,N_39269,N_39425);
nand U40721 (N_40721,N_39535,N_39840);
xnor U40722 (N_40722,N_39991,N_39079);
and U40723 (N_40723,N_39514,N_39847);
nor U40724 (N_40724,N_39680,N_39399);
nor U40725 (N_40725,N_39762,N_39730);
nor U40726 (N_40726,N_39641,N_39739);
nor U40727 (N_40727,N_39135,N_39773);
or U40728 (N_40728,N_39391,N_39752);
xor U40729 (N_40729,N_39935,N_39872);
xnor U40730 (N_40730,N_39596,N_39671);
or U40731 (N_40731,N_39218,N_39368);
nand U40732 (N_40732,N_39230,N_39226);
and U40733 (N_40733,N_39980,N_39604);
xnor U40734 (N_40734,N_39839,N_39114);
nand U40735 (N_40735,N_39131,N_39902);
nor U40736 (N_40736,N_39678,N_39316);
and U40737 (N_40737,N_39325,N_39366);
xnor U40738 (N_40738,N_39116,N_39613);
nand U40739 (N_40739,N_39431,N_39147);
nor U40740 (N_40740,N_39133,N_39902);
or U40741 (N_40741,N_39747,N_39104);
or U40742 (N_40742,N_39192,N_39543);
nand U40743 (N_40743,N_39318,N_39026);
xnor U40744 (N_40744,N_39978,N_39695);
nor U40745 (N_40745,N_39275,N_39970);
and U40746 (N_40746,N_39571,N_39079);
nand U40747 (N_40747,N_39309,N_39346);
xnor U40748 (N_40748,N_39301,N_39730);
xnor U40749 (N_40749,N_39477,N_39126);
and U40750 (N_40750,N_39901,N_39693);
and U40751 (N_40751,N_39925,N_39284);
nand U40752 (N_40752,N_39232,N_39928);
and U40753 (N_40753,N_39228,N_39332);
nand U40754 (N_40754,N_39909,N_39574);
nand U40755 (N_40755,N_39126,N_39947);
or U40756 (N_40756,N_39189,N_39914);
nor U40757 (N_40757,N_39606,N_39833);
or U40758 (N_40758,N_39315,N_39488);
and U40759 (N_40759,N_39740,N_39503);
or U40760 (N_40760,N_39653,N_39673);
nand U40761 (N_40761,N_39066,N_39117);
nor U40762 (N_40762,N_39017,N_39498);
and U40763 (N_40763,N_39361,N_39227);
xor U40764 (N_40764,N_39576,N_39748);
or U40765 (N_40765,N_39101,N_39032);
or U40766 (N_40766,N_39083,N_39409);
nand U40767 (N_40767,N_39922,N_39167);
nor U40768 (N_40768,N_39126,N_39643);
and U40769 (N_40769,N_39731,N_39744);
nand U40770 (N_40770,N_39377,N_39794);
nand U40771 (N_40771,N_39588,N_39204);
and U40772 (N_40772,N_39220,N_39058);
xor U40773 (N_40773,N_39885,N_39872);
and U40774 (N_40774,N_39772,N_39648);
xor U40775 (N_40775,N_39911,N_39928);
or U40776 (N_40776,N_39953,N_39321);
xor U40777 (N_40777,N_39384,N_39181);
nand U40778 (N_40778,N_39763,N_39718);
nor U40779 (N_40779,N_39062,N_39706);
nand U40780 (N_40780,N_39421,N_39680);
and U40781 (N_40781,N_39678,N_39752);
and U40782 (N_40782,N_39528,N_39618);
nand U40783 (N_40783,N_39599,N_39444);
or U40784 (N_40784,N_39415,N_39431);
and U40785 (N_40785,N_39356,N_39219);
nand U40786 (N_40786,N_39696,N_39946);
xor U40787 (N_40787,N_39636,N_39209);
and U40788 (N_40788,N_39139,N_39591);
nor U40789 (N_40789,N_39884,N_39958);
and U40790 (N_40790,N_39787,N_39683);
nand U40791 (N_40791,N_39974,N_39219);
and U40792 (N_40792,N_39200,N_39987);
and U40793 (N_40793,N_39646,N_39462);
and U40794 (N_40794,N_39275,N_39652);
nand U40795 (N_40795,N_39749,N_39516);
xnor U40796 (N_40796,N_39527,N_39044);
and U40797 (N_40797,N_39272,N_39744);
xor U40798 (N_40798,N_39280,N_39342);
nand U40799 (N_40799,N_39659,N_39462);
and U40800 (N_40800,N_39220,N_39890);
nor U40801 (N_40801,N_39112,N_39294);
nand U40802 (N_40802,N_39309,N_39642);
xnor U40803 (N_40803,N_39534,N_39673);
xnor U40804 (N_40804,N_39678,N_39020);
xor U40805 (N_40805,N_39872,N_39077);
nand U40806 (N_40806,N_39650,N_39367);
nor U40807 (N_40807,N_39293,N_39508);
nor U40808 (N_40808,N_39934,N_39939);
nand U40809 (N_40809,N_39789,N_39526);
and U40810 (N_40810,N_39187,N_39228);
or U40811 (N_40811,N_39191,N_39598);
nor U40812 (N_40812,N_39617,N_39414);
nor U40813 (N_40813,N_39293,N_39195);
xnor U40814 (N_40814,N_39193,N_39478);
and U40815 (N_40815,N_39754,N_39879);
nand U40816 (N_40816,N_39598,N_39652);
or U40817 (N_40817,N_39616,N_39487);
nand U40818 (N_40818,N_39130,N_39349);
nor U40819 (N_40819,N_39755,N_39384);
or U40820 (N_40820,N_39893,N_39947);
or U40821 (N_40821,N_39755,N_39176);
nor U40822 (N_40822,N_39983,N_39374);
nor U40823 (N_40823,N_39919,N_39893);
and U40824 (N_40824,N_39045,N_39322);
nand U40825 (N_40825,N_39492,N_39724);
nand U40826 (N_40826,N_39645,N_39529);
and U40827 (N_40827,N_39634,N_39362);
nor U40828 (N_40828,N_39098,N_39320);
nor U40829 (N_40829,N_39146,N_39751);
nand U40830 (N_40830,N_39495,N_39015);
nor U40831 (N_40831,N_39370,N_39275);
xnor U40832 (N_40832,N_39756,N_39204);
and U40833 (N_40833,N_39406,N_39423);
xnor U40834 (N_40834,N_39687,N_39336);
and U40835 (N_40835,N_39096,N_39577);
nand U40836 (N_40836,N_39182,N_39716);
nand U40837 (N_40837,N_39633,N_39514);
nor U40838 (N_40838,N_39853,N_39543);
nand U40839 (N_40839,N_39747,N_39999);
nand U40840 (N_40840,N_39435,N_39225);
and U40841 (N_40841,N_39167,N_39372);
or U40842 (N_40842,N_39464,N_39906);
xor U40843 (N_40843,N_39858,N_39143);
nand U40844 (N_40844,N_39991,N_39432);
xor U40845 (N_40845,N_39070,N_39801);
or U40846 (N_40846,N_39755,N_39770);
and U40847 (N_40847,N_39824,N_39569);
or U40848 (N_40848,N_39051,N_39109);
nor U40849 (N_40849,N_39827,N_39691);
and U40850 (N_40850,N_39089,N_39756);
nor U40851 (N_40851,N_39307,N_39652);
nor U40852 (N_40852,N_39031,N_39290);
nor U40853 (N_40853,N_39892,N_39888);
or U40854 (N_40854,N_39501,N_39059);
nand U40855 (N_40855,N_39226,N_39416);
nor U40856 (N_40856,N_39953,N_39387);
nor U40857 (N_40857,N_39335,N_39549);
xor U40858 (N_40858,N_39721,N_39806);
xor U40859 (N_40859,N_39279,N_39376);
xnor U40860 (N_40860,N_39758,N_39375);
nand U40861 (N_40861,N_39910,N_39120);
nor U40862 (N_40862,N_39612,N_39304);
xnor U40863 (N_40863,N_39298,N_39946);
nand U40864 (N_40864,N_39639,N_39229);
nor U40865 (N_40865,N_39424,N_39128);
nand U40866 (N_40866,N_39161,N_39615);
nand U40867 (N_40867,N_39016,N_39373);
and U40868 (N_40868,N_39931,N_39881);
nor U40869 (N_40869,N_39113,N_39119);
xor U40870 (N_40870,N_39516,N_39568);
or U40871 (N_40871,N_39755,N_39304);
or U40872 (N_40872,N_39801,N_39769);
or U40873 (N_40873,N_39506,N_39426);
nor U40874 (N_40874,N_39093,N_39939);
nand U40875 (N_40875,N_39910,N_39349);
and U40876 (N_40876,N_39217,N_39462);
xor U40877 (N_40877,N_39077,N_39798);
or U40878 (N_40878,N_39876,N_39850);
or U40879 (N_40879,N_39554,N_39136);
nand U40880 (N_40880,N_39148,N_39396);
or U40881 (N_40881,N_39818,N_39333);
or U40882 (N_40882,N_39844,N_39901);
or U40883 (N_40883,N_39486,N_39896);
and U40884 (N_40884,N_39993,N_39001);
or U40885 (N_40885,N_39286,N_39859);
nand U40886 (N_40886,N_39863,N_39656);
or U40887 (N_40887,N_39445,N_39522);
xnor U40888 (N_40888,N_39613,N_39002);
nand U40889 (N_40889,N_39097,N_39559);
nand U40890 (N_40890,N_39324,N_39162);
nand U40891 (N_40891,N_39840,N_39620);
and U40892 (N_40892,N_39654,N_39838);
nand U40893 (N_40893,N_39979,N_39389);
or U40894 (N_40894,N_39285,N_39511);
and U40895 (N_40895,N_39615,N_39177);
xor U40896 (N_40896,N_39606,N_39797);
xor U40897 (N_40897,N_39148,N_39397);
and U40898 (N_40898,N_39438,N_39504);
or U40899 (N_40899,N_39911,N_39573);
or U40900 (N_40900,N_39738,N_39443);
xor U40901 (N_40901,N_39759,N_39193);
and U40902 (N_40902,N_39019,N_39549);
xnor U40903 (N_40903,N_39502,N_39515);
nand U40904 (N_40904,N_39222,N_39293);
or U40905 (N_40905,N_39213,N_39495);
nand U40906 (N_40906,N_39056,N_39443);
or U40907 (N_40907,N_39221,N_39392);
nand U40908 (N_40908,N_39700,N_39804);
xnor U40909 (N_40909,N_39960,N_39017);
nor U40910 (N_40910,N_39484,N_39491);
nor U40911 (N_40911,N_39033,N_39596);
nand U40912 (N_40912,N_39984,N_39464);
xnor U40913 (N_40913,N_39080,N_39908);
or U40914 (N_40914,N_39493,N_39933);
and U40915 (N_40915,N_39364,N_39406);
and U40916 (N_40916,N_39593,N_39486);
xnor U40917 (N_40917,N_39601,N_39195);
xor U40918 (N_40918,N_39671,N_39781);
nor U40919 (N_40919,N_39424,N_39959);
or U40920 (N_40920,N_39495,N_39262);
and U40921 (N_40921,N_39025,N_39345);
nand U40922 (N_40922,N_39095,N_39810);
and U40923 (N_40923,N_39006,N_39787);
and U40924 (N_40924,N_39220,N_39243);
nand U40925 (N_40925,N_39625,N_39619);
or U40926 (N_40926,N_39141,N_39485);
or U40927 (N_40927,N_39066,N_39518);
and U40928 (N_40928,N_39912,N_39745);
nand U40929 (N_40929,N_39554,N_39024);
or U40930 (N_40930,N_39730,N_39909);
and U40931 (N_40931,N_39834,N_39121);
nand U40932 (N_40932,N_39163,N_39621);
nand U40933 (N_40933,N_39842,N_39953);
nand U40934 (N_40934,N_39853,N_39279);
nor U40935 (N_40935,N_39474,N_39273);
and U40936 (N_40936,N_39727,N_39693);
and U40937 (N_40937,N_39025,N_39137);
xnor U40938 (N_40938,N_39499,N_39245);
and U40939 (N_40939,N_39701,N_39343);
and U40940 (N_40940,N_39875,N_39242);
and U40941 (N_40941,N_39554,N_39713);
nor U40942 (N_40942,N_39697,N_39277);
or U40943 (N_40943,N_39911,N_39382);
nor U40944 (N_40944,N_39304,N_39515);
or U40945 (N_40945,N_39859,N_39569);
nand U40946 (N_40946,N_39011,N_39270);
xnor U40947 (N_40947,N_39327,N_39208);
or U40948 (N_40948,N_39071,N_39406);
or U40949 (N_40949,N_39963,N_39531);
nor U40950 (N_40950,N_39654,N_39159);
and U40951 (N_40951,N_39086,N_39163);
nand U40952 (N_40952,N_39530,N_39173);
xor U40953 (N_40953,N_39155,N_39311);
and U40954 (N_40954,N_39521,N_39859);
nand U40955 (N_40955,N_39624,N_39843);
nand U40956 (N_40956,N_39525,N_39841);
xnor U40957 (N_40957,N_39471,N_39120);
nand U40958 (N_40958,N_39487,N_39139);
nand U40959 (N_40959,N_39880,N_39230);
nor U40960 (N_40960,N_39848,N_39840);
or U40961 (N_40961,N_39855,N_39829);
and U40962 (N_40962,N_39211,N_39395);
and U40963 (N_40963,N_39419,N_39041);
xor U40964 (N_40964,N_39993,N_39751);
or U40965 (N_40965,N_39757,N_39252);
or U40966 (N_40966,N_39422,N_39309);
nand U40967 (N_40967,N_39586,N_39508);
nor U40968 (N_40968,N_39291,N_39395);
or U40969 (N_40969,N_39510,N_39033);
xor U40970 (N_40970,N_39666,N_39906);
nand U40971 (N_40971,N_39972,N_39101);
xor U40972 (N_40972,N_39669,N_39621);
nand U40973 (N_40973,N_39844,N_39361);
and U40974 (N_40974,N_39562,N_39649);
nand U40975 (N_40975,N_39222,N_39158);
xor U40976 (N_40976,N_39247,N_39219);
nor U40977 (N_40977,N_39707,N_39348);
and U40978 (N_40978,N_39767,N_39278);
or U40979 (N_40979,N_39480,N_39311);
xor U40980 (N_40980,N_39808,N_39918);
xor U40981 (N_40981,N_39398,N_39629);
xor U40982 (N_40982,N_39832,N_39370);
and U40983 (N_40983,N_39760,N_39611);
and U40984 (N_40984,N_39657,N_39526);
and U40985 (N_40985,N_39129,N_39602);
or U40986 (N_40986,N_39785,N_39124);
xor U40987 (N_40987,N_39808,N_39020);
nand U40988 (N_40988,N_39804,N_39047);
and U40989 (N_40989,N_39557,N_39068);
or U40990 (N_40990,N_39503,N_39897);
nor U40991 (N_40991,N_39669,N_39905);
and U40992 (N_40992,N_39810,N_39403);
or U40993 (N_40993,N_39399,N_39088);
nand U40994 (N_40994,N_39815,N_39533);
or U40995 (N_40995,N_39545,N_39444);
nand U40996 (N_40996,N_39448,N_39860);
xor U40997 (N_40997,N_39639,N_39362);
xnor U40998 (N_40998,N_39622,N_39060);
and U40999 (N_40999,N_39746,N_39834);
nand U41000 (N_41000,N_40898,N_40648);
nand U41001 (N_41001,N_40727,N_40938);
and U41002 (N_41002,N_40665,N_40435);
xor U41003 (N_41003,N_40960,N_40602);
or U41004 (N_41004,N_40145,N_40097);
or U41005 (N_41005,N_40300,N_40293);
nor U41006 (N_41006,N_40258,N_40715);
xnor U41007 (N_41007,N_40362,N_40691);
nand U41008 (N_41008,N_40378,N_40206);
nor U41009 (N_41009,N_40353,N_40538);
xor U41010 (N_41010,N_40979,N_40773);
nand U41011 (N_41011,N_40395,N_40970);
and U41012 (N_41012,N_40430,N_40038);
and U41013 (N_41013,N_40163,N_40758);
nor U41014 (N_41014,N_40320,N_40613);
and U41015 (N_41015,N_40630,N_40984);
nand U41016 (N_41016,N_40085,N_40713);
nand U41017 (N_41017,N_40906,N_40029);
nand U41018 (N_41018,N_40487,N_40221);
and U41019 (N_41019,N_40263,N_40025);
or U41020 (N_41020,N_40990,N_40522);
nor U41021 (N_41021,N_40809,N_40335);
nand U41022 (N_41022,N_40241,N_40526);
or U41023 (N_41023,N_40500,N_40352);
nor U41024 (N_41024,N_40683,N_40657);
and U41025 (N_41025,N_40739,N_40053);
nor U41026 (N_41026,N_40190,N_40316);
nor U41027 (N_41027,N_40942,N_40868);
nand U41028 (N_41028,N_40696,N_40034);
xor U41029 (N_41029,N_40975,N_40342);
or U41030 (N_41030,N_40746,N_40688);
or U41031 (N_41031,N_40872,N_40826);
and U41032 (N_41032,N_40076,N_40548);
xnor U41033 (N_41033,N_40349,N_40518);
or U41034 (N_41034,N_40059,N_40434);
nor U41035 (N_41035,N_40892,N_40109);
or U41036 (N_41036,N_40457,N_40172);
nand U41037 (N_41037,N_40618,N_40155);
and U41038 (N_41038,N_40649,N_40233);
nand U41039 (N_41039,N_40794,N_40503);
nand U41040 (N_41040,N_40302,N_40895);
and U41041 (N_41041,N_40592,N_40346);
and U41042 (N_41042,N_40420,N_40994);
xnor U41043 (N_41043,N_40472,N_40819);
nand U41044 (N_41044,N_40020,N_40069);
nor U41045 (N_41045,N_40308,N_40561);
or U41046 (N_41046,N_40900,N_40041);
xor U41047 (N_41047,N_40622,N_40735);
nor U41048 (N_41048,N_40778,N_40184);
or U41049 (N_41049,N_40763,N_40644);
xor U41050 (N_41050,N_40875,N_40912);
nand U41051 (N_41051,N_40516,N_40927);
xnor U41052 (N_41052,N_40901,N_40540);
and U41053 (N_41053,N_40929,N_40252);
nor U41054 (N_41054,N_40078,N_40523);
and U41055 (N_41055,N_40579,N_40358);
and U41056 (N_41056,N_40936,N_40808);
nand U41057 (N_41057,N_40517,N_40571);
nand U41058 (N_41058,N_40425,N_40963);
and U41059 (N_41059,N_40139,N_40314);
nor U41060 (N_41060,N_40507,N_40603);
and U41061 (N_41061,N_40806,N_40123);
nor U41062 (N_41062,N_40108,N_40598);
xor U41063 (N_41063,N_40610,N_40187);
or U41064 (N_41064,N_40676,N_40541);
xnor U41065 (N_41065,N_40110,N_40026);
nand U41066 (N_41066,N_40708,N_40064);
nand U41067 (N_41067,N_40762,N_40724);
nor U41068 (N_41068,N_40336,N_40721);
or U41069 (N_41069,N_40646,N_40181);
nand U41070 (N_41070,N_40334,N_40061);
nor U41071 (N_41071,N_40832,N_40031);
nand U41072 (N_41072,N_40364,N_40889);
and U41073 (N_41073,N_40261,N_40931);
nor U41074 (N_41074,N_40429,N_40392);
and U41075 (N_41075,N_40847,N_40703);
nor U41076 (N_41076,N_40286,N_40619);
xor U41077 (N_41077,N_40193,N_40318);
nor U41078 (N_41078,N_40483,N_40752);
and U41079 (N_41079,N_40486,N_40611);
xor U41080 (N_41080,N_40654,N_40480);
nor U41081 (N_41081,N_40478,N_40641);
and U41082 (N_41082,N_40958,N_40355);
or U41083 (N_41083,N_40527,N_40961);
nand U41084 (N_41084,N_40831,N_40192);
nor U41085 (N_41085,N_40780,N_40073);
nand U41086 (N_41086,N_40771,N_40423);
or U41087 (N_41087,N_40582,N_40617);
nor U41088 (N_41088,N_40162,N_40276);
and U41089 (N_41089,N_40573,N_40751);
and U41090 (N_41090,N_40666,N_40514);
xor U41091 (N_41091,N_40462,N_40825);
xor U41092 (N_41092,N_40852,N_40873);
and U41093 (N_41093,N_40081,N_40294);
nand U41094 (N_41094,N_40917,N_40481);
nand U41095 (N_41095,N_40333,N_40273);
or U41096 (N_41096,N_40543,N_40655);
and U41097 (N_41097,N_40063,N_40600);
xor U41098 (N_41098,N_40608,N_40547);
xor U41099 (N_41099,N_40301,N_40940);
and U41100 (N_41100,N_40419,N_40207);
xor U41101 (N_41101,N_40813,N_40783);
or U41102 (N_41102,N_40640,N_40304);
nand U41103 (N_41103,N_40374,N_40397);
nand U41104 (N_41104,N_40874,N_40521);
nor U41105 (N_41105,N_40891,N_40581);
and U41106 (N_41106,N_40839,N_40008);
nand U41107 (N_41107,N_40861,N_40638);
nand U41108 (N_41108,N_40989,N_40270);
nor U41109 (N_41109,N_40987,N_40766);
nor U41110 (N_41110,N_40645,N_40475);
and U41111 (N_41111,N_40634,N_40685);
xor U41112 (N_41112,N_40636,N_40256);
or U41113 (N_41113,N_40673,N_40052);
or U41114 (N_41114,N_40091,N_40531);
xnor U41115 (N_41115,N_40047,N_40787);
nand U41116 (N_41116,N_40653,N_40099);
nand U41117 (N_41117,N_40790,N_40601);
nor U41118 (N_41118,N_40152,N_40709);
and U41119 (N_41119,N_40268,N_40552);
nand U41120 (N_41120,N_40629,N_40862);
nand U41121 (N_41121,N_40197,N_40344);
and U41122 (N_41122,N_40239,N_40479);
nand U41123 (N_41123,N_40111,N_40465);
or U41124 (N_41124,N_40476,N_40447);
or U41125 (N_41125,N_40921,N_40381);
nor U41126 (N_41126,N_40048,N_40911);
nand U41127 (N_41127,N_40754,N_40855);
and U41128 (N_41128,N_40528,N_40730);
nand U41129 (N_41129,N_40216,N_40106);
nor U41130 (N_41130,N_40098,N_40606);
and U41131 (N_41131,N_40916,N_40818);
xnor U41132 (N_41132,N_40815,N_40237);
and U41133 (N_41133,N_40325,N_40198);
or U41134 (N_41134,N_40731,N_40222);
nand U41135 (N_41135,N_40712,N_40575);
nor U41136 (N_41136,N_40774,N_40442);
and U41137 (N_41137,N_40386,N_40050);
and U41138 (N_41138,N_40698,N_40201);
nand U41139 (N_41139,N_40443,N_40105);
xnor U41140 (N_41140,N_40343,N_40559);
and U41141 (N_41141,N_40717,N_40729);
or U41142 (N_41142,N_40436,N_40983);
nor U41143 (N_41143,N_40804,N_40032);
and U41144 (N_41144,N_40781,N_40793);
and U41145 (N_41145,N_40279,N_40812);
nor U41146 (N_41146,N_40470,N_40148);
and U41147 (N_41147,N_40136,N_40426);
or U41148 (N_41148,N_40980,N_40962);
nor U41149 (N_41149,N_40287,N_40096);
nor U41150 (N_41150,N_40623,N_40460);
xor U41151 (N_41151,N_40449,N_40332);
or U41152 (N_41152,N_40800,N_40492);
nor U41153 (N_41153,N_40121,N_40577);
xor U41154 (N_41154,N_40628,N_40632);
or U41155 (N_41155,N_40599,N_40382);
nor U41156 (N_41156,N_40350,N_40095);
nand U41157 (N_41157,N_40992,N_40694);
and U41158 (N_41158,N_40493,N_40094);
nor U41159 (N_41159,N_40950,N_40066);
or U41160 (N_41160,N_40775,N_40525);
nor U41161 (N_41161,N_40421,N_40678);
and U41162 (N_41162,N_40118,N_40489);
nor U41163 (N_41163,N_40651,N_40253);
nor U41164 (N_41164,N_40883,N_40033);
or U41165 (N_41165,N_40896,N_40652);
or U41166 (N_41166,N_40292,N_40376);
nor U41167 (N_41167,N_40843,N_40802);
nand U41168 (N_41168,N_40338,N_40505);
or U41169 (N_41169,N_40904,N_40718);
or U41170 (N_41170,N_40330,N_40490);
nor U41171 (N_41171,N_40488,N_40639);
and U41172 (N_41172,N_40250,N_40871);
or U41173 (N_41173,N_40377,N_40366);
or U41174 (N_41174,N_40669,N_40520);
nor U41175 (N_41175,N_40633,N_40035);
or U41176 (N_41176,N_40170,N_40563);
nor U41177 (N_41177,N_40814,N_40532);
nor U41178 (N_41178,N_40161,N_40022);
xor U41179 (N_41179,N_40234,N_40977);
nor U41180 (N_41180,N_40680,N_40733);
or U41181 (N_41181,N_40251,N_40930);
nor U41182 (N_41182,N_40908,N_40863);
and U41183 (N_41183,N_40589,N_40844);
nand U41184 (N_41184,N_40278,N_40011);
nand U41185 (N_41185,N_40012,N_40555);
or U41186 (N_41186,N_40671,N_40760);
and U41187 (N_41187,N_40837,N_40084);
nor U41188 (N_41188,N_40845,N_40051);
or U41189 (N_41189,N_40219,N_40755);
nor U41190 (N_41190,N_40941,N_40913);
nor U41191 (N_41191,N_40448,N_40792);
and U41192 (N_41192,N_40211,N_40565);
nor U41193 (N_41193,N_40959,N_40295);
xnor U41194 (N_41194,N_40890,N_40827);
or U41195 (N_41195,N_40070,N_40180);
nor U41196 (N_41196,N_40003,N_40922);
and U41197 (N_41197,N_40248,N_40176);
or U41198 (N_41198,N_40939,N_40955);
and U41199 (N_41199,N_40328,N_40568);
xor U41200 (N_41200,N_40112,N_40807);
and U41201 (N_41201,N_40113,N_40867);
and U41202 (N_41202,N_40074,N_40393);
and U41203 (N_41203,N_40667,N_40734);
nand U41204 (N_41204,N_40410,N_40985);
nor U41205 (N_41205,N_40409,N_40329);
xnor U41206 (N_41206,N_40438,N_40836);
and U41207 (N_41207,N_40972,N_40714);
xor U41208 (N_41208,N_40923,N_40976);
nand U41209 (N_41209,N_40864,N_40662);
nand U41210 (N_41210,N_40511,N_40828);
xnor U41211 (N_41211,N_40779,N_40595);
nor U41212 (N_41212,N_40010,N_40798);
or U41213 (N_41213,N_40590,N_40146);
or U41214 (N_41214,N_40782,N_40236);
and U41215 (N_41215,N_40786,N_40834);
nor U41216 (N_41216,N_40416,N_40030);
nor U41217 (N_41217,N_40143,N_40466);
nor U41218 (N_41218,N_40040,N_40124);
nand U41219 (N_41219,N_40439,N_40083);
and U41220 (N_41220,N_40171,N_40303);
and U41221 (N_41221,N_40705,N_40291);
xor U41222 (N_41222,N_40089,N_40337);
nand U41223 (N_41223,N_40816,N_40150);
nor U41224 (N_41224,N_40805,N_40103);
and U41225 (N_41225,N_40627,N_40907);
and U41226 (N_41226,N_40137,N_40860);
or U41227 (N_41227,N_40365,N_40056);
or U41228 (N_41228,N_40188,N_40620);
nand U41229 (N_41229,N_40557,N_40427);
nor U41230 (N_41230,N_40943,N_40138);
xor U41231 (N_41231,N_40995,N_40933);
and U41232 (N_41232,N_40659,N_40529);
xnor U41233 (N_41233,N_40037,N_40341);
or U41234 (N_41234,N_40903,N_40130);
and U41235 (N_41235,N_40888,N_40288);
nor U41236 (N_41236,N_40272,N_40497);
and U41237 (N_41237,N_40367,N_40700);
and U41238 (N_41238,N_40177,N_40550);
and U41239 (N_41239,N_40530,N_40125);
nand U41240 (N_41240,N_40887,N_40668);
nand U41241 (N_41241,N_40701,N_40626);
or U41242 (N_41242,N_40591,N_40249);
nand U41243 (N_41243,N_40881,N_40928);
nand U41244 (N_41244,N_40723,N_40495);
xnor U41245 (N_41245,N_40937,N_40686);
or U41246 (N_41246,N_40379,N_40046);
or U41247 (N_41247,N_40042,N_40978);
nand U41248 (N_41248,N_40405,N_40494);
nand U41249 (N_41249,N_40126,N_40504);
xnor U41250 (N_41250,N_40820,N_40092);
nand U41251 (N_41251,N_40660,N_40450);
nor U41252 (N_41252,N_40182,N_40326);
or U41253 (N_41253,N_40391,N_40658);
nor U41254 (N_41254,N_40886,N_40833);
xnor U41255 (N_41255,N_40689,N_40157);
nor U41256 (N_41256,N_40100,N_40323);
and U41257 (N_41257,N_40297,N_40502);
nor U41258 (N_41258,N_40310,N_40934);
or U41259 (N_41259,N_40885,N_40266);
nor U41260 (N_41260,N_40451,N_40537);
or U41261 (N_41261,N_40741,N_40803);
and U41262 (N_41262,N_40461,N_40199);
nand U41263 (N_41263,N_40684,N_40210);
and U41264 (N_41264,N_40607,N_40021);
or U41265 (N_41265,N_40414,N_40850);
and U41266 (N_41266,N_40422,N_40919);
nand U41267 (N_41267,N_40749,N_40104);
nand U41268 (N_41268,N_40956,N_40799);
nand U41269 (N_41269,N_40005,N_40851);
and U41270 (N_41270,N_40158,N_40404);
and U41271 (N_41271,N_40156,N_40769);
xnor U41272 (N_41272,N_40072,N_40508);
and U41273 (N_41273,N_40880,N_40213);
and U41274 (N_41274,N_40356,N_40870);
nand U41275 (N_41275,N_40675,N_40394);
nand U41276 (N_41276,N_40133,N_40093);
nand U41277 (N_41277,N_40569,N_40604);
nor U41278 (N_41278,N_40687,N_40372);
nand U41279 (N_41279,N_40214,N_40817);
xnor U41280 (N_41280,N_40361,N_40299);
nand U41281 (N_41281,N_40765,N_40593);
and U41282 (N_41282,N_40255,N_40631);
nor U41283 (N_41283,N_40560,N_40240);
nand U41284 (N_41284,N_40464,N_40597);
nor U41285 (N_41285,N_40045,N_40585);
nor U41286 (N_41286,N_40609,N_40722);
nand U41287 (N_41287,N_40202,N_40468);
and U41288 (N_41288,N_40205,N_40235);
xor U41289 (N_41289,N_40002,N_40244);
nand U41290 (N_41290,N_40168,N_40884);
and U41291 (N_41291,N_40067,N_40265);
and U41292 (N_41292,N_40354,N_40305);
xor U41293 (N_41293,N_40153,N_40122);
and U41294 (N_41294,N_40981,N_40043);
xor U41295 (N_41295,N_40742,N_40544);
xor U41296 (N_41296,N_40179,N_40313);
xnor U41297 (N_41297,N_40456,N_40716);
xor U41298 (N_41298,N_40183,N_40120);
nor U41299 (N_41299,N_40062,N_40797);
and U41300 (N_41300,N_40140,N_40801);
and U41301 (N_41301,N_40951,N_40228);
nand U41302 (N_41302,N_40196,N_40661);
xor U41303 (N_41303,N_40194,N_40612);
nand U41304 (N_41304,N_40107,N_40952);
and U41305 (N_41305,N_40396,N_40079);
or U41306 (N_41306,N_40406,N_40699);
or U41307 (N_41307,N_40259,N_40877);
or U41308 (N_41308,N_40398,N_40368);
or U41309 (N_41309,N_40102,N_40643);
and U41310 (N_41310,N_40509,N_40835);
nand U41311 (N_41311,N_40088,N_40208);
nor U41312 (N_41312,N_40348,N_40428);
or U41313 (N_41313,N_40160,N_40949);
and U41314 (N_41314,N_40647,N_40650);
nand U41315 (N_41315,N_40412,N_40954);
and U41316 (N_41316,N_40535,N_40151);
and U41317 (N_41317,N_40369,N_40849);
and U41318 (N_41318,N_40223,N_40229);
nand U41319 (N_41319,N_40562,N_40411);
nor U41320 (N_41320,N_40238,N_40656);
and U41321 (N_41321,N_40173,N_40384);
or U41322 (N_41322,N_40080,N_40914);
and U41323 (N_41323,N_40446,N_40246);
and U41324 (N_41324,N_40371,N_40473);
or U41325 (N_41325,N_40791,N_40496);
and U41326 (N_41326,N_40424,N_40498);
xnor U41327 (N_41327,N_40576,N_40621);
xor U41328 (N_41328,N_40925,N_40924);
xnor U41329 (N_41329,N_40129,N_40857);
and U41330 (N_41330,N_40269,N_40232);
nor U41331 (N_41331,N_40719,N_40454);
and U41332 (N_41332,N_40400,N_40387);
nand U41333 (N_41333,N_40433,N_40345);
and U41334 (N_41334,N_40225,N_40471);
and U41335 (N_41335,N_40477,N_40389);
xor U41336 (N_41336,N_40524,N_40677);
xnor U41337 (N_41337,N_40039,N_40191);
nor U41338 (N_41338,N_40309,N_40044);
or U41339 (N_41339,N_40262,N_40853);
and U41340 (N_41340,N_40932,N_40566);
nor U41341 (N_41341,N_40909,N_40131);
xnor U41342 (N_41342,N_40280,N_40534);
nor U41343 (N_41343,N_40578,N_40247);
and U41344 (N_41344,N_40926,N_40664);
nand U41345 (N_41345,N_40770,N_40014);
and U41346 (N_41346,N_40441,N_40065);
xnor U41347 (N_41347,N_40811,N_40215);
nand U41348 (N_41348,N_40728,N_40823);
nand U41349 (N_41349,N_40738,N_40681);
or U41350 (N_41350,N_40347,N_40966);
nor U41351 (N_41351,N_40403,N_40615);
xor U41352 (N_41352,N_40127,N_40154);
nor U41353 (N_41353,N_40455,N_40948);
nand U41354 (N_41354,N_40218,N_40245);
or U41355 (N_41355,N_40277,N_40558);
or U41356 (N_41356,N_40854,N_40554);
and U41357 (N_41357,N_40087,N_40401);
or U41358 (N_41358,N_40788,N_40458);
or U41359 (N_41359,N_40946,N_40075);
and U41360 (N_41360,N_40117,N_40306);
xnor U41361 (N_41361,N_40467,N_40474);
nor U41362 (N_41362,N_40842,N_40999);
nor U41363 (N_41363,N_40663,N_40296);
or U41364 (N_41364,N_40973,N_40281);
or U41365 (N_41365,N_40408,N_40822);
xnor U41366 (N_41366,N_40785,N_40830);
and U41367 (N_41367,N_40546,N_40415);
nand U41368 (N_41368,N_40690,N_40726);
and U41369 (N_41369,N_40167,N_40918);
nand U41370 (N_41370,N_40082,N_40230);
nand U41371 (N_41371,N_40128,N_40789);
xor U41372 (N_41372,N_40290,N_40119);
nand U41373 (N_41373,N_40795,N_40242);
nor U41374 (N_41374,N_40897,N_40549);
nor U41375 (N_41375,N_40567,N_40957);
or U41376 (N_41376,N_40370,N_40536);
nand U41377 (N_41377,N_40209,N_40407);
or U41378 (N_41378,N_40399,N_40178);
and U41379 (N_41379,N_40444,N_40510);
nor U41380 (N_41380,N_40596,N_40697);
or U41381 (N_41381,N_40587,N_40380);
and U41382 (N_41382,N_40777,N_40635);
and U41383 (N_41383,N_40231,N_40899);
xnor U41384 (N_41384,N_40289,N_40588);
or U41385 (N_41385,N_40796,N_40418);
xor U41386 (N_41386,N_40616,N_40055);
nand U41387 (N_41387,N_40169,N_40768);
or U41388 (N_41388,N_40840,N_40203);
or U41389 (N_41389,N_40311,N_40116);
xor U41390 (N_41390,N_40743,N_40077);
xor U41391 (N_41391,N_40315,N_40463);
xnor U41392 (N_41392,N_40969,N_40115);
nand U41393 (N_41393,N_40340,N_40737);
or U41394 (N_41394,N_40865,N_40114);
nand U41395 (N_41395,N_40267,N_40375);
and U41396 (N_41396,N_40431,N_40132);
nor U41397 (N_41397,N_40693,N_40711);
and U41398 (N_41398,N_40545,N_40185);
xor U41399 (N_41399,N_40945,N_40485);
xnor U41400 (N_41400,N_40134,N_40846);
nand U41401 (N_41401,N_40905,N_40829);
nor U41402 (N_41402,N_40226,N_40482);
and U41403 (N_41403,N_40810,N_40953);
nand U41404 (N_41404,N_40284,N_40821);
xnor U41405 (N_41405,N_40858,N_40260);
nand U41406 (N_41406,N_40965,N_40570);
and U41407 (N_41407,N_40533,N_40838);
xnor U41408 (N_41408,N_40707,N_40227);
or U41409 (N_41409,N_40982,N_40710);
or U41410 (N_41410,N_40893,N_40748);
nor U41411 (N_41411,N_40702,N_40841);
or U41412 (N_41412,N_40204,N_40432);
nor U41413 (N_41413,N_40357,N_40772);
nand U41414 (N_41414,N_40704,N_40679);
nor U41415 (N_41415,N_40776,N_40915);
nor U41416 (N_41416,N_40007,N_40017);
and U41417 (N_41417,N_40165,N_40740);
xnor U41418 (N_41418,N_40993,N_40019);
and U41419 (N_41419,N_40383,N_40583);
nand U41420 (N_41420,N_40220,N_40445);
nand U41421 (N_41421,N_40317,N_40339);
xor U41422 (N_41422,N_40642,N_40186);
xnor U41423 (N_41423,N_40388,N_40417);
nand U41424 (N_41424,N_40506,N_40068);
nand U41425 (N_41425,N_40254,N_40024);
nand U41426 (N_41426,N_40257,N_40876);
nor U41427 (N_41427,N_40501,N_40513);
and U41428 (N_41428,N_40453,N_40920);
or U41429 (N_41429,N_40016,N_40373);
xor U41430 (N_41430,N_40149,N_40910);
nor U41431 (N_41431,N_40968,N_40164);
and U41432 (N_41432,N_40060,N_40000);
nand U41433 (N_41433,N_40013,N_40224);
and U41434 (N_41434,N_40351,N_40159);
or U41435 (N_41435,N_40624,N_40009);
or U41436 (N_41436,N_40878,N_40243);
nor U41437 (N_41437,N_40459,N_40848);
or U41438 (N_41438,N_40135,N_40499);
xor U41439 (N_41439,N_40580,N_40036);
nand U41440 (N_41440,N_40745,N_40469);
or U41441 (N_41441,N_40586,N_40264);
and U41442 (N_41442,N_40312,N_40553);
xnor U41443 (N_41443,N_40556,N_40166);
and U41444 (N_41444,N_40331,N_40764);
nand U41445 (N_41445,N_40856,N_40452);
and U41446 (N_41446,N_40058,N_40935);
nor U41447 (N_41447,N_40001,N_40998);
or U41448 (N_41448,N_40988,N_40512);
nand U41449 (N_41449,N_40997,N_40141);
nor U41450 (N_41450,N_40319,N_40195);
xnor U41451 (N_41451,N_40967,N_40271);
nand U41452 (N_41452,N_40437,N_40637);
or U41453 (N_41453,N_40732,N_40584);
nor U41454 (N_41454,N_40006,N_40614);
nor U41455 (N_41455,N_40744,N_40484);
nor U41456 (N_41456,N_40018,N_40757);
nand U41457 (N_41457,N_40519,N_40200);
xnor U41458 (N_41458,N_40071,N_40625);
nor U41459 (N_41459,N_40147,N_40307);
or U41460 (N_41460,N_40275,N_40101);
and U41461 (N_41461,N_40359,N_40682);
and U41462 (N_41462,N_40725,N_40015);
or U41463 (N_41463,N_40144,N_40974);
nor U41464 (N_41464,N_40217,N_40282);
and U41465 (N_41465,N_40574,N_40327);
or U41466 (N_41466,N_40515,N_40023);
and U41467 (N_41467,N_40736,N_40706);
nand U41468 (N_41468,N_40539,N_40759);
xor U41469 (N_41469,N_40004,N_40944);
or U41470 (N_41470,N_40054,N_40321);
and U41471 (N_41471,N_40142,N_40440);
or U41472 (N_41472,N_40283,N_40090);
nor U41473 (N_41473,N_40996,N_40363);
and U41474 (N_41474,N_40413,N_40285);
or U41475 (N_41475,N_40385,N_40298);
and U41476 (N_41476,N_40866,N_40964);
xor U41477 (N_41477,N_40027,N_40894);
and U41478 (N_41478,N_40189,N_40986);
xnor U41479 (N_41479,N_40784,N_40761);
xor U41480 (N_41480,N_40542,N_40753);
xor U41481 (N_41481,N_40674,N_40947);
nand U41482 (N_41482,N_40057,N_40750);
xor U41483 (N_41483,N_40869,N_40971);
xor U41484 (N_41484,N_40274,N_40692);
and U41485 (N_41485,N_40672,N_40491);
xnor U41486 (N_41486,N_40991,N_40572);
xnor U41487 (N_41487,N_40551,N_40756);
nand U41488 (N_41488,N_40594,N_40882);
nor U41489 (N_41489,N_40390,N_40360);
nand U41490 (N_41490,N_40902,N_40174);
nor U41491 (N_41491,N_40564,N_40028);
xor U41492 (N_41492,N_40695,N_40049);
nor U41493 (N_41493,N_40322,N_40324);
xnor U41494 (N_41494,N_40086,N_40767);
nand U41495 (N_41495,N_40212,N_40720);
and U41496 (N_41496,N_40824,N_40175);
or U41497 (N_41497,N_40670,N_40747);
xor U41498 (N_41498,N_40605,N_40879);
or U41499 (N_41499,N_40402,N_40859);
nand U41500 (N_41500,N_40263,N_40324);
nand U41501 (N_41501,N_40084,N_40121);
or U41502 (N_41502,N_40346,N_40933);
nand U41503 (N_41503,N_40795,N_40515);
nor U41504 (N_41504,N_40936,N_40572);
nor U41505 (N_41505,N_40180,N_40676);
xnor U41506 (N_41506,N_40230,N_40981);
nor U41507 (N_41507,N_40672,N_40179);
or U41508 (N_41508,N_40475,N_40744);
or U41509 (N_41509,N_40164,N_40066);
or U41510 (N_41510,N_40473,N_40873);
and U41511 (N_41511,N_40068,N_40099);
or U41512 (N_41512,N_40558,N_40823);
xor U41513 (N_41513,N_40745,N_40951);
xor U41514 (N_41514,N_40587,N_40320);
nor U41515 (N_41515,N_40773,N_40583);
or U41516 (N_41516,N_40802,N_40872);
nor U41517 (N_41517,N_40301,N_40165);
or U41518 (N_41518,N_40444,N_40653);
xor U41519 (N_41519,N_40028,N_40613);
nor U41520 (N_41520,N_40941,N_40435);
nor U41521 (N_41521,N_40774,N_40062);
nor U41522 (N_41522,N_40812,N_40377);
nor U41523 (N_41523,N_40830,N_40332);
nand U41524 (N_41524,N_40668,N_40240);
nand U41525 (N_41525,N_40579,N_40248);
and U41526 (N_41526,N_40238,N_40130);
and U41527 (N_41527,N_40821,N_40002);
xor U41528 (N_41528,N_40353,N_40573);
nand U41529 (N_41529,N_40109,N_40593);
nor U41530 (N_41530,N_40646,N_40999);
and U41531 (N_41531,N_40992,N_40943);
nand U41532 (N_41532,N_40074,N_40649);
xnor U41533 (N_41533,N_40842,N_40743);
or U41534 (N_41534,N_40543,N_40427);
xor U41535 (N_41535,N_40890,N_40779);
xnor U41536 (N_41536,N_40994,N_40675);
or U41537 (N_41537,N_40087,N_40772);
or U41538 (N_41538,N_40874,N_40492);
or U41539 (N_41539,N_40176,N_40035);
xor U41540 (N_41540,N_40563,N_40095);
nor U41541 (N_41541,N_40708,N_40453);
nor U41542 (N_41542,N_40921,N_40232);
nor U41543 (N_41543,N_40927,N_40735);
xnor U41544 (N_41544,N_40025,N_40131);
xnor U41545 (N_41545,N_40753,N_40393);
nand U41546 (N_41546,N_40791,N_40452);
or U41547 (N_41547,N_40514,N_40698);
xor U41548 (N_41548,N_40792,N_40953);
xor U41549 (N_41549,N_40569,N_40726);
and U41550 (N_41550,N_40992,N_40377);
xor U41551 (N_41551,N_40724,N_40212);
nand U41552 (N_41552,N_40364,N_40938);
or U41553 (N_41553,N_40887,N_40994);
and U41554 (N_41554,N_40722,N_40281);
and U41555 (N_41555,N_40126,N_40114);
nand U41556 (N_41556,N_40793,N_40601);
or U41557 (N_41557,N_40401,N_40573);
nand U41558 (N_41558,N_40317,N_40334);
xor U41559 (N_41559,N_40660,N_40482);
nor U41560 (N_41560,N_40198,N_40428);
and U41561 (N_41561,N_40547,N_40271);
nor U41562 (N_41562,N_40341,N_40665);
nand U41563 (N_41563,N_40032,N_40317);
nand U41564 (N_41564,N_40202,N_40791);
or U41565 (N_41565,N_40797,N_40686);
nor U41566 (N_41566,N_40064,N_40744);
or U41567 (N_41567,N_40555,N_40281);
xnor U41568 (N_41568,N_40159,N_40562);
xnor U41569 (N_41569,N_40180,N_40904);
nor U41570 (N_41570,N_40801,N_40914);
xnor U41571 (N_41571,N_40019,N_40656);
xnor U41572 (N_41572,N_40016,N_40660);
xnor U41573 (N_41573,N_40700,N_40960);
nand U41574 (N_41574,N_40687,N_40953);
and U41575 (N_41575,N_40572,N_40077);
nor U41576 (N_41576,N_40605,N_40854);
nor U41577 (N_41577,N_40295,N_40473);
and U41578 (N_41578,N_40334,N_40300);
or U41579 (N_41579,N_40375,N_40088);
nand U41580 (N_41580,N_40894,N_40475);
or U41581 (N_41581,N_40808,N_40549);
xor U41582 (N_41582,N_40920,N_40770);
nor U41583 (N_41583,N_40962,N_40341);
or U41584 (N_41584,N_40250,N_40202);
or U41585 (N_41585,N_40573,N_40015);
xor U41586 (N_41586,N_40564,N_40598);
or U41587 (N_41587,N_40607,N_40837);
and U41588 (N_41588,N_40263,N_40863);
nor U41589 (N_41589,N_40324,N_40032);
and U41590 (N_41590,N_40917,N_40953);
nor U41591 (N_41591,N_40524,N_40003);
nand U41592 (N_41592,N_40822,N_40142);
and U41593 (N_41593,N_40549,N_40112);
and U41594 (N_41594,N_40574,N_40753);
and U41595 (N_41595,N_40447,N_40401);
xnor U41596 (N_41596,N_40262,N_40101);
nand U41597 (N_41597,N_40522,N_40038);
or U41598 (N_41598,N_40738,N_40763);
and U41599 (N_41599,N_40663,N_40425);
and U41600 (N_41600,N_40491,N_40917);
and U41601 (N_41601,N_40071,N_40080);
nand U41602 (N_41602,N_40134,N_40380);
xor U41603 (N_41603,N_40655,N_40455);
or U41604 (N_41604,N_40294,N_40474);
nor U41605 (N_41605,N_40348,N_40000);
nor U41606 (N_41606,N_40538,N_40247);
xnor U41607 (N_41607,N_40761,N_40303);
xnor U41608 (N_41608,N_40603,N_40369);
or U41609 (N_41609,N_40370,N_40236);
and U41610 (N_41610,N_40876,N_40757);
or U41611 (N_41611,N_40877,N_40134);
and U41612 (N_41612,N_40807,N_40340);
nor U41613 (N_41613,N_40507,N_40532);
xnor U41614 (N_41614,N_40300,N_40305);
nand U41615 (N_41615,N_40880,N_40740);
or U41616 (N_41616,N_40973,N_40582);
and U41617 (N_41617,N_40246,N_40809);
or U41618 (N_41618,N_40635,N_40337);
and U41619 (N_41619,N_40646,N_40667);
nor U41620 (N_41620,N_40682,N_40191);
nor U41621 (N_41621,N_40009,N_40693);
xor U41622 (N_41622,N_40218,N_40307);
nand U41623 (N_41623,N_40710,N_40579);
or U41624 (N_41624,N_40215,N_40064);
and U41625 (N_41625,N_40626,N_40731);
and U41626 (N_41626,N_40221,N_40532);
or U41627 (N_41627,N_40860,N_40055);
and U41628 (N_41628,N_40746,N_40309);
nand U41629 (N_41629,N_40564,N_40463);
nor U41630 (N_41630,N_40242,N_40228);
nand U41631 (N_41631,N_40567,N_40638);
nand U41632 (N_41632,N_40808,N_40752);
or U41633 (N_41633,N_40350,N_40523);
and U41634 (N_41634,N_40955,N_40600);
nor U41635 (N_41635,N_40156,N_40415);
and U41636 (N_41636,N_40609,N_40841);
and U41637 (N_41637,N_40918,N_40577);
xnor U41638 (N_41638,N_40122,N_40096);
nand U41639 (N_41639,N_40217,N_40606);
nand U41640 (N_41640,N_40727,N_40514);
nor U41641 (N_41641,N_40297,N_40589);
and U41642 (N_41642,N_40927,N_40066);
nand U41643 (N_41643,N_40461,N_40023);
xnor U41644 (N_41644,N_40581,N_40658);
nor U41645 (N_41645,N_40847,N_40356);
and U41646 (N_41646,N_40436,N_40683);
nand U41647 (N_41647,N_40246,N_40099);
xor U41648 (N_41648,N_40111,N_40398);
nand U41649 (N_41649,N_40747,N_40034);
and U41650 (N_41650,N_40501,N_40813);
xor U41651 (N_41651,N_40338,N_40168);
nor U41652 (N_41652,N_40174,N_40017);
nand U41653 (N_41653,N_40991,N_40759);
or U41654 (N_41654,N_40538,N_40813);
xor U41655 (N_41655,N_40066,N_40864);
or U41656 (N_41656,N_40027,N_40808);
xnor U41657 (N_41657,N_40388,N_40657);
and U41658 (N_41658,N_40026,N_40130);
nor U41659 (N_41659,N_40503,N_40857);
nor U41660 (N_41660,N_40500,N_40997);
xor U41661 (N_41661,N_40431,N_40845);
nand U41662 (N_41662,N_40559,N_40607);
xor U41663 (N_41663,N_40706,N_40635);
or U41664 (N_41664,N_40055,N_40812);
nor U41665 (N_41665,N_40965,N_40095);
and U41666 (N_41666,N_40172,N_40087);
nand U41667 (N_41667,N_40288,N_40634);
and U41668 (N_41668,N_40630,N_40189);
or U41669 (N_41669,N_40329,N_40889);
xor U41670 (N_41670,N_40270,N_40235);
or U41671 (N_41671,N_40409,N_40289);
nand U41672 (N_41672,N_40906,N_40762);
and U41673 (N_41673,N_40050,N_40302);
nand U41674 (N_41674,N_40060,N_40588);
xnor U41675 (N_41675,N_40390,N_40357);
nand U41676 (N_41676,N_40813,N_40842);
xor U41677 (N_41677,N_40460,N_40448);
nor U41678 (N_41678,N_40392,N_40369);
and U41679 (N_41679,N_40970,N_40061);
xor U41680 (N_41680,N_40927,N_40252);
or U41681 (N_41681,N_40150,N_40881);
or U41682 (N_41682,N_40630,N_40721);
or U41683 (N_41683,N_40894,N_40119);
and U41684 (N_41684,N_40360,N_40861);
and U41685 (N_41685,N_40646,N_40767);
or U41686 (N_41686,N_40383,N_40766);
and U41687 (N_41687,N_40579,N_40722);
xor U41688 (N_41688,N_40634,N_40862);
xor U41689 (N_41689,N_40544,N_40046);
or U41690 (N_41690,N_40063,N_40385);
nor U41691 (N_41691,N_40303,N_40498);
nand U41692 (N_41692,N_40938,N_40432);
and U41693 (N_41693,N_40737,N_40697);
nand U41694 (N_41694,N_40660,N_40021);
nor U41695 (N_41695,N_40888,N_40136);
xor U41696 (N_41696,N_40201,N_40877);
nor U41697 (N_41697,N_40556,N_40090);
and U41698 (N_41698,N_40198,N_40033);
nor U41699 (N_41699,N_40972,N_40419);
nand U41700 (N_41700,N_40391,N_40972);
nand U41701 (N_41701,N_40612,N_40641);
xor U41702 (N_41702,N_40793,N_40904);
nand U41703 (N_41703,N_40364,N_40581);
xor U41704 (N_41704,N_40527,N_40497);
nand U41705 (N_41705,N_40387,N_40281);
nor U41706 (N_41706,N_40533,N_40710);
and U41707 (N_41707,N_40883,N_40580);
nor U41708 (N_41708,N_40882,N_40496);
nand U41709 (N_41709,N_40401,N_40426);
and U41710 (N_41710,N_40620,N_40184);
nor U41711 (N_41711,N_40955,N_40495);
nor U41712 (N_41712,N_40758,N_40276);
nor U41713 (N_41713,N_40227,N_40090);
xnor U41714 (N_41714,N_40739,N_40164);
and U41715 (N_41715,N_40439,N_40255);
and U41716 (N_41716,N_40465,N_40942);
or U41717 (N_41717,N_40363,N_40229);
xor U41718 (N_41718,N_40696,N_40960);
xor U41719 (N_41719,N_40992,N_40330);
nor U41720 (N_41720,N_40411,N_40370);
nor U41721 (N_41721,N_40677,N_40186);
nor U41722 (N_41722,N_40523,N_40730);
nand U41723 (N_41723,N_40525,N_40176);
or U41724 (N_41724,N_40304,N_40798);
or U41725 (N_41725,N_40935,N_40688);
nand U41726 (N_41726,N_40037,N_40215);
nand U41727 (N_41727,N_40696,N_40857);
and U41728 (N_41728,N_40989,N_40646);
and U41729 (N_41729,N_40446,N_40156);
or U41730 (N_41730,N_40736,N_40109);
or U41731 (N_41731,N_40149,N_40688);
or U41732 (N_41732,N_40356,N_40329);
nor U41733 (N_41733,N_40368,N_40612);
or U41734 (N_41734,N_40088,N_40319);
and U41735 (N_41735,N_40663,N_40420);
xnor U41736 (N_41736,N_40028,N_40542);
or U41737 (N_41737,N_40632,N_40540);
or U41738 (N_41738,N_40122,N_40532);
nand U41739 (N_41739,N_40309,N_40040);
xnor U41740 (N_41740,N_40559,N_40427);
xor U41741 (N_41741,N_40369,N_40794);
or U41742 (N_41742,N_40599,N_40668);
nand U41743 (N_41743,N_40269,N_40998);
xnor U41744 (N_41744,N_40734,N_40983);
nor U41745 (N_41745,N_40020,N_40140);
xor U41746 (N_41746,N_40116,N_40020);
and U41747 (N_41747,N_40798,N_40847);
nand U41748 (N_41748,N_40054,N_40197);
xnor U41749 (N_41749,N_40256,N_40240);
and U41750 (N_41750,N_40095,N_40834);
nand U41751 (N_41751,N_40703,N_40256);
or U41752 (N_41752,N_40021,N_40447);
nand U41753 (N_41753,N_40329,N_40778);
or U41754 (N_41754,N_40952,N_40942);
and U41755 (N_41755,N_40777,N_40904);
and U41756 (N_41756,N_40050,N_40647);
nand U41757 (N_41757,N_40108,N_40943);
nand U41758 (N_41758,N_40920,N_40339);
or U41759 (N_41759,N_40041,N_40127);
nor U41760 (N_41760,N_40581,N_40462);
or U41761 (N_41761,N_40936,N_40191);
nor U41762 (N_41762,N_40641,N_40681);
or U41763 (N_41763,N_40483,N_40753);
or U41764 (N_41764,N_40709,N_40570);
xnor U41765 (N_41765,N_40367,N_40540);
nor U41766 (N_41766,N_40606,N_40584);
nand U41767 (N_41767,N_40422,N_40415);
nand U41768 (N_41768,N_40151,N_40917);
or U41769 (N_41769,N_40300,N_40136);
nand U41770 (N_41770,N_40419,N_40061);
or U41771 (N_41771,N_40259,N_40796);
and U41772 (N_41772,N_40258,N_40366);
xor U41773 (N_41773,N_40605,N_40585);
or U41774 (N_41774,N_40399,N_40817);
and U41775 (N_41775,N_40967,N_40750);
nor U41776 (N_41776,N_40763,N_40514);
nand U41777 (N_41777,N_40914,N_40881);
and U41778 (N_41778,N_40487,N_40047);
and U41779 (N_41779,N_40070,N_40189);
nor U41780 (N_41780,N_40627,N_40812);
and U41781 (N_41781,N_40954,N_40827);
xor U41782 (N_41782,N_40056,N_40258);
xnor U41783 (N_41783,N_40701,N_40093);
nand U41784 (N_41784,N_40487,N_40993);
or U41785 (N_41785,N_40025,N_40770);
or U41786 (N_41786,N_40867,N_40192);
nor U41787 (N_41787,N_40927,N_40995);
nor U41788 (N_41788,N_40990,N_40205);
and U41789 (N_41789,N_40887,N_40843);
nor U41790 (N_41790,N_40261,N_40680);
xnor U41791 (N_41791,N_40557,N_40971);
and U41792 (N_41792,N_40128,N_40841);
nand U41793 (N_41793,N_40298,N_40900);
nand U41794 (N_41794,N_40431,N_40912);
nand U41795 (N_41795,N_40904,N_40586);
nand U41796 (N_41796,N_40350,N_40942);
nor U41797 (N_41797,N_40765,N_40162);
or U41798 (N_41798,N_40573,N_40953);
or U41799 (N_41799,N_40691,N_40191);
nand U41800 (N_41800,N_40366,N_40785);
and U41801 (N_41801,N_40363,N_40590);
nor U41802 (N_41802,N_40878,N_40846);
nor U41803 (N_41803,N_40620,N_40055);
nand U41804 (N_41804,N_40426,N_40608);
and U41805 (N_41805,N_40175,N_40648);
or U41806 (N_41806,N_40316,N_40385);
xor U41807 (N_41807,N_40229,N_40847);
nand U41808 (N_41808,N_40108,N_40780);
xnor U41809 (N_41809,N_40246,N_40918);
nor U41810 (N_41810,N_40660,N_40759);
xnor U41811 (N_41811,N_40220,N_40178);
and U41812 (N_41812,N_40963,N_40370);
and U41813 (N_41813,N_40325,N_40088);
and U41814 (N_41814,N_40085,N_40497);
nand U41815 (N_41815,N_40093,N_40669);
nor U41816 (N_41816,N_40727,N_40197);
nand U41817 (N_41817,N_40059,N_40628);
nor U41818 (N_41818,N_40787,N_40825);
nor U41819 (N_41819,N_40512,N_40585);
and U41820 (N_41820,N_40521,N_40672);
xnor U41821 (N_41821,N_40589,N_40313);
nor U41822 (N_41822,N_40006,N_40801);
or U41823 (N_41823,N_40755,N_40502);
nor U41824 (N_41824,N_40001,N_40135);
or U41825 (N_41825,N_40296,N_40497);
nand U41826 (N_41826,N_40776,N_40334);
xor U41827 (N_41827,N_40639,N_40513);
nor U41828 (N_41828,N_40275,N_40899);
xnor U41829 (N_41829,N_40254,N_40620);
nand U41830 (N_41830,N_40823,N_40618);
nand U41831 (N_41831,N_40339,N_40787);
nor U41832 (N_41832,N_40117,N_40042);
xor U41833 (N_41833,N_40376,N_40169);
nor U41834 (N_41834,N_40127,N_40855);
and U41835 (N_41835,N_40083,N_40226);
nand U41836 (N_41836,N_40513,N_40440);
or U41837 (N_41837,N_40169,N_40648);
or U41838 (N_41838,N_40242,N_40080);
or U41839 (N_41839,N_40714,N_40007);
xnor U41840 (N_41840,N_40386,N_40279);
xnor U41841 (N_41841,N_40984,N_40569);
and U41842 (N_41842,N_40035,N_40989);
or U41843 (N_41843,N_40163,N_40387);
and U41844 (N_41844,N_40619,N_40778);
nand U41845 (N_41845,N_40314,N_40865);
nor U41846 (N_41846,N_40855,N_40010);
or U41847 (N_41847,N_40846,N_40671);
nor U41848 (N_41848,N_40323,N_40021);
nand U41849 (N_41849,N_40116,N_40562);
and U41850 (N_41850,N_40740,N_40785);
and U41851 (N_41851,N_40212,N_40391);
nand U41852 (N_41852,N_40767,N_40732);
xor U41853 (N_41853,N_40259,N_40109);
or U41854 (N_41854,N_40423,N_40051);
xnor U41855 (N_41855,N_40242,N_40914);
xor U41856 (N_41856,N_40557,N_40107);
and U41857 (N_41857,N_40129,N_40640);
nand U41858 (N_41858,N_40776,N_40221);
nand U41859 (N_41859,N_40260,N_40685);
xor U41860 (N_41860,N_40730,N_40980);
or U41861 (N_41861,N_40701,N_40196);
and U41862 (N_41862,N_40555,N_40942);
xor U41863 (N_41863,N_40503,N_40094);
nor U41864 (N_41864,N_40016,N_40786);
and U41865 (N_41865,N_40567,N_40318);
nand U41866 (N_41866,N_40683,N_40191);
nand U41867 (N_41867,N_40897,N_40378);
nor U41868 (N_41868,N_40336,N_40692);
xor U41869 (N_41869,N_40248,N_40386);
nor U41870 (N_41870,N_40575,N_40861);
and U41871 (N_41871,N_40265,N_40720);
and U41872 (N_41872,N_40901,N_40645);
nand U41873 (N_41873,N_40799,N_40828);
xnor U41874 (N_41874,N_40353,N_40523);
nor U41875 (N_41875,N_40609,N_40566);
nand U41876 (N_41876,N_40160,N_40907);
nand U41877 (N_41877,N_40744,N_40984);
xnor U41878 (N_41878,N_40080,N_40796);
nand U41879 (N_41879,N_40444,N_40929);
and U41880 (N_41880,N_40218,N_40851);
and U41881 (N_41881,N_40902,N_40613);
or U41882 (N_41882,N_40125,N_40771);
or U41883 (N_41883,N_40021,N_40543);
and U41884 (N_41884,N_40896,N_40975);
and U41885 (N_41885,N_40894,N_40273);
xnor U41886 (N_41886,N_40642,N_40528);
nand U41887 (N_41887,N_40495,N_40683);
and U41888 (N_41888,N_40043,N_40730);
nand U41889 (N_41889,N_40502,N_40013);
nand U41890 (N_41890,N_40332,N_40839);
nor U41891 (N_41891,N_40070,N_40895);
nand U41892 (N_41892,N_40187,N_40955);
and U41893 (N_41893,N_40039,N_40639);
or U41894 (N_41894,N_40557,N_40420);
and U41895 (N_41895,N_40447,N_40450);
and U41896 (N_41896,N_40554,N_40787);
nand U41897 (N_41897,N_40077,N_40641);
nor U41898 (N_41898,N_40558,N_40865);
and U41899 (N_41899,N_40258,N_40036);
and U41900 (N_41900,N_40750,N_40217);
xor U41901 (N_41901,N_40002,N_40316);
or U41902 (N_41902,N_40091,N_40803);
xnor U41903 (N_41903,N_40517,N_40101);
nor U41904 (N_41904,N_40778,N_40084);
xor U41905 (N_41905,N_40254,N_40603);
xnor U41906 (N_41906,N_40991,N_40664);
or U41907 (N_41907,N_40893,N_40435);
and U41908 (N_41908,N_40199,N_40872);
nor U41909 (N_41909,N_40843,N_40653);
xnor U41910 (N_41910,N_40613,N_40016);
or U41911 (N_41911,N_40050,N_40831);
and U41912 (N_41912,N_40772,N_40710);
or U41913 (N_41913,N_40503,N_40030);
nand U41914 (N_41914,N_40844,N_40018);
or U41915 (N_41915,N_40799,N_40886);
xnor U41916 (N_41916,N_40068,N_40753);
or U41917 (N_41917,N_40186,N_40093);
xnor U41918 (N_41918,N_40850,N_40078);
xnor U41919 (N_41919,N_40736,N_40128);
nand U41920 (N_41920,N_40197,N_40781);
and U41921 (N_41921,N_40391,N_40066);
and U41922 (N_41922,N_40138,N_40561);
or U41923 (N_41923,N_40378,N_40382);
nand U41924 (N_41924,N_40077,N_40623);
xor U41925 (N_41925,N_40241,N_40350);
xnor U41926 (N_41926,N_40370,N_40660);
xnor U41927 (N_41927,N_40129,N_40400);
and U41928 (N_41928,N_40591,N_40620);
xnor U41929 (N_41929,N_40866,N_40506);
nor U41930 (N_41930,N_40485,N_40300);
or U41931 (N_41931,N_40994,N_40717);
and U41932 (N_41932,N_40633,N_40063);
nand U41933 (N_41933,N_40575,N_40893);
and U41934 (N_41934,N_40684,N_40000);
nand U41935 (N_41935,N_40111,N_40861);
nand U41936 (N_41936,N_40132,N_40935);
and U41937 (N_41937,N_40760,N_40011);
or U41938 (N_41938,N_40909,N_40946);
xor U41939 (N_41939,N_40705,N_40543);
or U41940 (N_41940,N_40539,N_40983);
or U41941 (N_41941,N_40947,N_40301);
nand U41942 (N_41942,N_40334,N_40808);
nand U41943 (N_41943,N_40929,N_40113);
and U41944 (N_41944,N_40476,N_40954);
xor U41945 (N_41945,N_40635,N_40238);
or U41946 (N_41946,N_40330,N_40600);
or U41947 (N_41947,N_40189,N_40510);
xor U41948 (N_41948,N_40298,N_40255);
nor U41949 (N_41949,N_40317,N_40201);
nand U41950 (N_41950,N_40142,N_40489);
nor U41951 (N_41951,N_40136,N_40992);
xnor U41952 (N_41952,N_40149,N_40881);
nand U41953 (N_41953,N_40448,N_40990);
and U41954 (N_41954,N_40625,N_40227);
xnor U41955 (N_41955,N_40666,N_40383);
xor U41956 (N_41956,N_40453,N_40577);
xnor U41957 (N_41957,N_40174,N_40018);
nor U41958 (N_41958,N_40351,N_40199);
nor U41959 (N_41959,N_40520,N_40907);
nor U41960 (N_41960,N_40409,N_40472);
or U41961 (N_41961,N_40213,N_40247);
xnor U41962 (N_41962,N_40010,N_40748);
nand U41963 (N_41963,N_40976,N_40868);
and U41964 (N_41964,N_40840,N_40120);
or U41965 (N_41965,N_40790,N_40702);
or U41966 (N_41966,N_40303,N_40787);
xor U41967 (N_41967,N_40642,N_40177);
or U41968 (N_41968,N_40794,N_40767);
or U41969 (N_41969,N_40678,N_40251);
or U41970 (N_41970,N_40454,N_40876);
or U41971 (N_41971,N_40478,N_40679);
and U41972 (N_41972,N_40946,N_40939);
and U41973 (N_41973,N_40947,N_40653);
nor U41974 (N_41974,N_40333,N_40940);
nand U41975 (N_41975,N_40141,N_40455);
xnor U41976 (N_41976,N_40013,N_40527);
and U41977 (N_41977,N_40213,N_40374);
xnor U41978 (N_41978,N_40125,N_40685);
or U41979 (N_41979,N_40566,N_40153);
nor U41980 (N_41980,N_40064,N_40216);
nor U41981 (N_41981,N_40923,N_40418);
nand U41982 (N_41982,N_40437,N_40064);
nor U41983 (N_41983,N_40343,N_40678);
nor U41984 (N_41984,N_40718,N_40908);
xor U41985 (N_41985,N_40585,N_40195);
or U41986 (N_41986,N_40575,N_40970);
xor U41987 (N_41987,N_40770,N_40487);
or U41988 (N_41988,N_40425,N_40758);
nor U41989 (N_41989,N_40242,N_40359);
or U41990 (N_41990,N_40120,N_40305);
or U41991 (N_41991,N_40053,N_40063);
and U41992 (N_41992,N_40962,N_40553);
or U41993 (N_41993,N_40400,N_40604);
and U41994 (N_41994,N_40163,N_40130);
or U41995 (N_41995,N_40747,N_40020);
nand U41996 (N_41996,N_40612,N_40811);
nand U41997 (N_41997,N_40938,N_40482);
or U41998 (N_41998,N_40565,N_40667);
nand U41999 (N_41999,N_40602,N_40255);
xor U42000 (N_42000,N_41233,N_41913);
xnor U42001 (N_42001,N_41114,N_41561);
nor U42002 (N_42002,N_41470,N_41627);
and U42003 (N_42003,N_41001,N_41088);
nand U42004 (N_42004,N_41006,N_41829);
nor U42005 (N_42005,N_41574,N_41304);
or U42006 (N_42006,N_41038,N_41839);
and U42007 (N_42007,N_41336,N_41931);
xor U42008 (N_42008,N_41965,N_41184);
and U42009 (N_42009,N_41365,N_41337);
and U42010 (N_42010,N_41824,N_41711);
nor U42011 (N_42011,N_41348,N_41558);
and U42012 (N_42012,N_41515,N_41925);
nor U42013 (N_42013,N_41548,N_41709);
and U42014 (N_42014,N_41897,N_41194);
nor U42015 (N_42015,N_41275,N_41953);
nand U42016 (N_42016,N_41540,N_41320);
xor U42017 (N_42017,N_41232,N_41325);
xnor U42018 (N_42018,N_41361,N_41922);
nor U42019 (N_42019,N_41085,N_41732);
xor U42020 (N_42020,N_41706,N_41154);
xor U42021 (N_42021,N_41899,N_41794);
nand U42022 (N_42022,N_41370,N_41591);
xor U42023 (N_42023,N_41151,N_41921);
and U42024 (N_42024,N_41625,N_41052);
nor U42025 (N_42025,N_41780,N_41496);
nand U42026 (N_42026,N_41411,N_41293);
and U42027 (N_42027,N_41251,N_41074);
nand U42028 (N_42028,N_41754,N_41613);
nor U42029 (N_42029,N_41306,N_41248);
nor U42030 (N_42030,N_41908,N_41107);
nor U42031 (N_42031,N_41472,N_41047);
nor U42032 (N_42032,N_41919,N_41125);
or U42033 (N_42033,N_41405,N_41281);
or U42034 (N_42034,N_41299,N_41997);
nor U42035 (N_42035,N_41105,N_41934);
and U42036 (N_42036,N_41420,N_41791);
nand U42037 (N_42037,N_41900,N_41367);
and U42038 (N_42038,N_41970,N_41830);
and U42039 (N_42039,N_41172,N_41401);
xor U42040 (N_42040,N_41433,N_41021);
nor U42041 (N_42041,N_41977,N_41297);
nor U42042 (N_42042,N_41759,N_41529);
and U42043 (N_42043,N_41744,N_41728);
and U42044 (N_42044,N_41139,N_41643);
or U42045 (N_42045,N_41078,N_41395);
or U42046 (N_42046,N_41158,N_41661);
nand U42047 (N_42047,N_41784,N_41523);
and U42048 (N_42048,N_41875,N_41214);
or U42049 (N_42049,N_41017,N_41926);
nor U42050 (N_42050,N_41327,N_41901);
and U42051 (N_42051,N_41705,N_41222);
nor U42052 (N_42052,N_41659,N_41115);
and U42053 (N_42053,N_41487,N_41537);
nor U42054 (N_42054,N_41013,N_41493);
or U42055 (N_42055,N_41841,N_41007);
nand U42056 (N_42056,N_41328,N_41140);
and U42057 (N_42057,N_41174,N_41520);
and U42058 (N_42058,N_41510,N_41255);
nand U42059 (N_42059,N_41695,N_41192);
and U42060 (N_42060,N_41800,N_41112);
xnor U42061 (N_42061,N_41102,N_41747);
or U42062 (N_42062,N_41024,N_41851);
and U42063 (N_42063,N_41513,N_41447);
nand U42064 (N_42064,N_41768,N_41729);
and U42065 (N_42065,N_41873,N_41188);
nor U42066 (N_42066,N_41681,N_41850);
and U42067 (N_42067,N_41062,N_41952);
and U42068 (N_42068,N_41628,N_41687);
xor U42069 (N_42069,N_41059,N_41334);
or U42070 (N_42070,N_41782,N_41189);
xnor U42071 (N_42071,N_41355,N_41212);
or U42072 (N_42072,N_41670,N_41050);
and U42073 (N_42073,N_41415,N_41616);
or U42074 (N_42074,N_41950,N_41371);
and U42075 (N_42075,N_41620,N_41864);
xor U42076 (N_42076,N_41083,N_41402);
nor U42077 (N_42077,N_41142,N_41905);
nand U42078 (N_42078,N_41823,N_41976);
and U42079 (N_42079,N_41476,N_41404);
xnor U42080 (N_42080,N_41565,N_41081);
xor U42081 (N_42081,N_41508,N_41097);
and U42082 (N_42082,N_41571,N_41482);
or U42083 (N_42083,N_41204,N_41494);
or U42084 (N_42084,N_41036,N_41291);
nand U42085 (N_42085,N_41180,N_41126);
xor U42086 (N_42086,N_41497,N_41086);
or U42087 (N_42087,N_41621,N_41844);
nand U42088 (N_42088,N_41141,N_41727);
nor U42089 (N_42089,N_41303,N_41505);
xor U42090 (N_42090,N_41846,N_41169);
or U42091 (N_42091,N_41506,N_41671);
and U42092 (N_42092,N_41243,N_41985);
nand U42093 (N_42093,N_41301,N_41279);
nor U42094 (N_42094,N_41998,N_41409);
xnor U42095 (N_42095,N_41993,N_41321);
xnor U42096 (N_42096,N_41544,N_41040);
xnor U42097 (N_42097,N_41018,N_41449);
or U42098 (N_42098,N_41489,N_41596);
nor U42099 (N_42099,N_41814,N_41752);
and U42100 (N_42100,N_41957,N_41623);
nor U42101 (N_42101,N_41208,N_41015);
xor U42102 (N_42102,N_41210,N_41207);
nand U42103 (N_42103,N_41758,N_41278);
xor U42104 (N_42104,N_41426,N_41444);
and U42105 (N_42105,N_41676,N_41556);
nor U42106 (N_42106,N_41032,N_41329);
xor U42107 (N_42107,N_41090,N_41111);
nand U42108 (N_42108,N_41884,N_41324);
and U42109 (N_42109,N_41165,N_41516);
nor U42110 (N_42110,N_41481,N_41969);
xor U42111 (N_42111,N_41295,N_41309);
nor U42112 (N_42112,N_41029,N_41091);
and U42113 (N_42113,N_41491,N_41842);
or U42114 (N_42114,N_41332,N_41138);
nor U42115 (N_42115,N_41719,N_41722);
and U42116 (N_42116,N_41099,N_41200);
nor U42117 (N_42117,N_41594,N_41354);
nor U42118 (N_42118,N_41294,N_41073);
or U42119 (N_42119,N_41615,N_41464);
xor U42120 (N_42120,N_41642,N_41445);
nand U42121 (N_42121,N_41166,N_41912);
nor U42122 (N_42122,N_41937,N_41767);
and U42123 (N_42123,N_41252,N_41714);
or U42124 (N_42124,N_41492,N_41638);
xor U42125 (N_42125,N_41810,N_41080);
nand U42126 (N_42126,N_41503,N_41265);
xnor U42127 (N_42127,N_41490,N_41406);
and U42128 (N_42128,N_41225,N_41807);
or U42129 (N_42129,N_41739,N_41101);
nand U42130 (N_42130,N_41688,N_41231);
nand U42131 (N_42131,N_41622,N_41173);
or U42132 (N_42132,N_41096,N_41757);
or U42133 (N_42133,N_41109,N_41702);
and U42134 (N_42134,N_41575,N_41219);
nor U42135 (N_42135,N_41742,N_41879);
or U42136 (N_42136,N_41820,N_41907);
and U42137 (N_42137,N_41347,N_41462);
nor U42138 (N_42138,N_41534,N_41763);
xor U42139 (N_42139,N_41284,N_41037);
nand U42140 (N_42140,N_41813,N_41734);
xor U42141 (N_42141,N_41022,N_41667);
or U42142 (N_42142,N_41778,N_41197);
and U42143 (N_42143,N_41185,N_41634);
xor U42144 (N_42144,N_41205,N_41906);
nor U42145 (N_42145,N_41010,N_41753);
nor U42146 (N_42146,N_41887,N_41104);
xnor U42147 (N_42147,N_41836,N_41587);
nor U42148 (N_42148,N_41193,N_41771);
and U42149 (N_42149,N_41443,N_41726);
nand U42150 (N_42150,N_41809,N_41240);
or U42151 (N_42151,N_41380,N_41379);
and U42152 (N_42152,N_41150,N_41927);
and U42153 (N_42153,N_41382,N_41220);
nor U42154 (N_42154,N_41647,N_41894);
nand U42155 (N_42155,N_41811,N_41176);
and U42156 (N_42156,N_41880,N_41501);
nand U42157 (N_42157,N_41393,N_41968);
xor U42158 (N_42158,N_41499,N_41788);
and U42159 (N_42159,N_41226,N_41941);
and U42160 (N_42160,N_41322,N_41290);
nand U42161 (N_42161,N_41580,N_41025);
or U42162 (N_42162,N_41590,N_41979);
xnor U42163 (N_42163,N_41770,N_41860);
xnor U42164 (N_42164,N_41692,N_41133);
nor U42165 (N_42165,N_41902,N_41439);
nand U42166 (N_42166,N_41127,N_41773);
xnor U42167 (N_42167,N_41572,N_41678);
nand U42168 (N_42168,N_41690,N_41391);
and U42169 (N_42169,N_41145,N_41498);
xor U42170 (N_42170,N_41626,N_41871);
nor U42171 (N_42171,N_41701,N_41458);
nand U42172 (N_42172,N_41817,N_41377);
nand U42173 (N_42173,N_41507,N_41808);
or U42174 (N_42174,N_41256,N_41271);
nor U42175 (N_42175,N_41478,N_41488);
xnor U42176 (N_42176,N_41543,N_41630);
nor U42177 (N_42177,N_41500,N_41044);
nand U42178 (N_42178,N_41341,N_41241);
nor U42179 (N_42179,N_41253,N_41796);
xnor U42180 (N_42180,N_41518,N_41170);
nand U42181 (N_42181,N_41117,N_41054);
xor U42182 (N_42182,N_41190,N_41751);
nand U42183 (N_42183,N_41463,N_41581);
nand U42184 (N_42184,N_41582,N_41885);
or U42185 (N_42185,N_41373,N_41664);
nand U42186 (N_42186,N_41629,N_41954);
xor U42187 (N_42187,N_41455,N_41124);
xnor U42188 (N_42188,N_41797,N_41110);
nor U42189 (N_42189,N_41378,N_41855);
nor U42190 (N_42190,N_41635,N_41364);
nor U42191 (N_42191,N_41994,N_41394);
xnor U42192 (N_42192,N_41883,N_41662);
or U42193 (N_42193,N_41223,N_41895);
and U42194 (N_42194,N_41749,N_41002);
or U42195 (N_42195,N_41057,N_41483);
and U42196 (N_42196,N_41031,N_41552);
xor U42197 (N_42197,N_41183,N_41238);
nand U42198 (N_42198,N_41358,N_41438);
and U42199 (N_42199,N_41260,N_41048);
and U42200 (N_42200,N_41199,N_41425);
nor U42201 (N_42201,N_41624,N_41106);
nand U42202 (N_42202,N_41089,N_41264);
nor U42203 (N_42203,N_41446,N_41051);
and U42204 (N_42204,N_41870,N_41452);
nand U42205 (N_42205,N_41178,N_41202);
nor U42206 (N_42206,N_41655,N_41863);
xnor U42207 (N_42207,N_41563,N_41063);
or U42208 (N_42208,N_41689,N_41266);
nand U42209 (N_42209,N_41802,N_41362);
nand U42210 (N_42210,N_41612,N_41512);
nor U42211 (N_42211,N_41995,N_41318);
or U42212 (N_42212,N_41056,N_41718);
and U42213 (N_42213,N_41019,N_41277);
and U42214 (N_42214,N_41603,N_41053);
xor U42215 (N_42215,N_41929,N_41453);
xnor U42216 (N_42216,N_41514,N_41245);
nor U42217 (N_42217,N_41974,N_41387);
nand U42218 (N_42218,N_41177,N_41323);
or U42219 (N_42219,N_41351,N_41805);
nand U42220 (N_42220,N_41485,N_41632);
nand U42221 (N_42221,N_41822,N_41866);
nor U42222 (N_42222,N_41878,N_41413);
nand U42223 (N_42223,N_41748,N_41967);
or U42224 (N_42224,N_41691,N_41546);
nor U42225 (N_42225,N_41082,N_41641);
nand U42226 (N_42226,N_41132,N_41148);
xnor U42227 (N_42227,N_41710,N_41774);
nor U42228 (N_42228,N_41588,N_41239);
or U42229 (N_42229,N_41388,N_41084);
or U42230 (N_42230,N_41665,N_41923);
nand U42231 (N_42231,N_41298,N_41285);
or U42232 (N_42232,N_41799,N_41416);
nand U42233 (N_42233,N_41567,N_41254);
nor U42234 (N_42234,N_41123,N_41595);
nor U42235 (N_42235,N_41731,N_41903);
nand U42236 (N_42236,N_41960,N_41168);
or U42237 (N_42237,N_41509,N_41660);
nor U42238 (N_42238,N_41242,N_41831);
nor U42239 (N_42239,N_41760,N_41636);
or U42240 (N_42240,N_41466,N_41435);
nor U42241 (N_42241,N_41221,N_41717);
xor U42242 (N_42242,N_41686,N_41064);
nor U42243 (N_42243,N_41834,N_41975);
nand U42244 (N_42244,N_41874,N_41450);
xnor U42245 (N_42245,N_41033,N_41209);
or U42246 (N_42246,N_41619,N_41585);
nand U42247 (N_42247,N_41973,N_41989);
nand U42248 (N_42248,N_41704,N_41777);
nor U42249 (N_42249,N_41972,N_41889);
nor U42250 (N_42250,N_41026,N_41034);
nor U42251 (N_42251,N_41495,N_41217);
xnor U42252 (N_42252,N_41943,N_41418);
nand U42253 (N_42253,N_41288,N_41287);
xor U42254 (N_42254,N_41521,N_41745);
nor U42255 (N_42255,N_41683,N_41386);
xnor U42256 (N_42256,N_41949,N_41804);
or U42257 (N_42257,N_41366,N_41042);
xnor U42258 (N_42258,N_41790,N_41892);
nand U42259 (N_42259,N_41849,N_41633);
nand U42260 (N_42260,N_41750,N_41740);
and U42261 (N_42261,N_41360,N_41584);
or U42262 (N_42262,N_41668,N_41611);
and U42263 (N_42263,N_41396,N_41795);
and U42264 (N_42264,N_41988,N_41631);
or U42265 (N_42265,N_41357,N_41312);
xor U42266 (N_42266,N_41310,N_41964);
nand U42267 (N_42267,N_41087,N_41832);
xor U42268 (N_42268,N_41069,N_41996);
and U42269 (N_42269,N_41261,N_41282);
or U42270 (N_42270,N_41039,N_41076);
nor U42271 (N_42271,N_41385,N_41144);
nand U42272 (N_42272,N_41314,N_41249);
nand U42273 (N_42273,N_41606,N_41666);
nand U42274 (N_42274,N_41349,N_41502);
xnor U42275 (N_42275,N_41825,N_41372);
nor U42276 (N_42276,N_41339,N_41600);
nand U42277 (N_42277,N_41955,N_41566);
or U42278 (N_42278,N_41736,N_41030);
nand U42279 (N_42279,N_41715,N_41067);
and U42280 (N_42280,N_41335,N_41916);
xor U42281 (N_42281,N_41545,N_41761);
and U42282 (N_42282,N_41143,N_41129);
nor U42283 (N_42283,N_41776,N_41557);
and U42284 (N_42284,N_41685,N_41441);
or U42285 (N_42285,N_41161,N_41077);
nor U42286 (N_42286,N_41066,N_41363);
and U42287 (N_42287,N_41837,N_41191);
or U42288 (N_42288,N_41990,N_41187);
nand U42289 (N_42289,N_41610,N_41517);
and U42290 (N_42290,N_41697,N_41227);
nand U42291 (N_42291,N_41307,N_41898);
nand U42292 (N_42292,N_41999,N_41422);
nor U42293 (N_42293,N_41987,N_41663);
nand U42294 (N_42294,N_41856,N_41340);
xnor U42295 (N_42295,N_41308,N_41963);
and U42296 (N_42296,N_41986,N_41300);
or U42297 (N_42297,N_41043,N_41068);
nand U42298 (N_42298,N_41716,N_41136);
or U42299 (N_42299,N_41060,N_41932);
xnor U42300 (N_42300,N_41682,N_41146);
or U42301 (N_42301,N_41707,N_41005);
nor U42302 (N_42302,N_41576,N_41381);
or U42303 (N_42303,N_41270,N_41951);
nand U42304 (N_42304,N_41764,N_41779);
nand U42305 (N_42305,N_41984,N_41302);
xor U42306 (N_42306,N_41946,N_41467);
or U42307 (N_42307,N_41474,N_41838);
xnor U42308 (N_42308,N_41679,N_41504);
nand U42309 (N_42309,N_41675,N_41792);
xnor U42310 (N_42310,N_41672,N_41945);
xor U42311 (N_42311,N_41128,N_41234);
xnor U42312 (N_42312,N_41599,N_41201);
or U42313 (N_42313,N_41374,N_41762);
nor U42314 (N_42314,N_41465,N_41915);
nor U42315 (N_42315,N_41211,N_41156);
or U42316 (N_42316,N_41434,N_41135);
nor U42317 (N_42317,N_41421,N_41738);
or U42318 (N_42318,N_41100,N_41654);
nor U42319 (N_42319,N_41843,N_41353);
xnor U42320 (N_42320,N_41547,N_41167);
xnor U42321 (N_42321,N_41930,N_41533);
nand U42322 (N_42322,N_41645,N_41833);
and U42323 (N_42323,N_41528,N_41646);
xnor U42324 (N_42324,N_41392,N_41819);
or U42325 (N_42325,N_41818,N_41657);
nor U42326 (N_42326,N_41121,N_41028);
and U42327 (N_42327,N_41317,N_41120);
nand U42328 (N_42328,N_41586,N_41027);
nand U42329 (N_42329,N_41648,N_41947);
xnor U42330 (N_42330,N_41075,N_41562);
or U42331 (N_42331,N_41847,N_41787);
nor U42332 (N_42332,N_41730,N_41541);
and U42333 (N_42333,N_41250,N_41700);
xnor U42334 (N_42334,N_41246,N_41338);
xor U42335 (N_42335,N_41094,N_41958);
nand U42336 (N_42336,N_41538,N_41186);
nor U42337 (N_42337,N_41607,N_41213);
nor U42338 (N_42338,N_41786,N_41971);
nand U42339 (N_42339,N_41555,N_41652);
and U42340 (N_42340,N_41536,N_41583);
and U42341 (N_42341,N_41263,N_41535);
or U42342 (N_42342,N_41229,N_41480);
xnor U42343 (N_42343,N_41737,N_41342);
nor U42344 (N_42344,N_41609,N_41755);
nand U42345 (N_42345,N_41525,N_41982);
xor U42346 (N_42346,N_41359,N_41431);
xor U42347 (N_42347,N_41769,N_41673);
nor U42348 (N_42348,N_41092,N_41400);
and U42349 (N_42349,N_41840,N_41602);
nand U42350 (N_42350,N_41980,N_41313);
nor U42351 (N_42351,N_41430,N_41333);
and U42352 (N_42352,N_41526,N_41775);
and U42353 (N_42353,N_41933,N_41134);
and U42354 (N_42354,N_41639,N_41798);
nand U42355 (N_42355,N_41460,N_41551);
nand U42356 (N_42356,N_41071,N_41981);
and U42357 (N_42357,N_41414,N_41826);
or U42358 (N_42358,N_41868,N_41821);
xor U42359 (N_42359,N_41131,N_41041);
and U42360 (N_42360,N_41095,N_41137);
nor U42361 (N_42361,N_41049,N_41407);
nor U42362 (N_42362,N_41854,N_41806);
nor U42363 (N_42363,N_41848,N_41924);
xor U42364 (N_42364,N_41549,N_41108);
xor U42365 (N_42365,N_41274,N_41983);
or U42366 (N_42366,N_41532,N_41914);
and U42367 (N_42367,N_41319,N_41326);
nand U42368 (N_42368,N_41772,N_41157);
xnor U42369 (N_42369,N_41936,N_41230);
or U42370 (N_42370,N_41098,N_41789);
nand U42371 (N_42371,N_41247,N_41605);
nor U42372 (N_42372,N_41195,N_41542);
and U42373 (N_42373,N_41257,N_41862);
nand U42374 (N_42374,N_41218,N_41920);
or U42375 (N_42375,N_41289,N_41035);
or U42376 (N_42376,N_41079,N_41948);
nand U42377 (N_42377,N_41153,N_41781);
xnor U42378 (N_42378,N_41577,N_41559);
nand U42379 (N_42379,N_41020,N_41011);
xnor U42380 (N_42380,N_41162,N_41429);
xor U42381 (N_42381,N_41045,N_41680);
or U42382 (N_42382,N_41944,N_41723);
nand U42383 (N_42383,N_41305,N_41940);
xnor U42384 (N_42384,N_41592,N_41262);
nor U42385 (N_42385,N_41070,N_41093);
nor U42386 (N_42386,N_41935,N_41276);
nor U42387 (N_42387,N_41065,N_41910);
xor U42388 (N_42388,N_41442,N_41658);
xor U42389 (N_42389,N_41149,N_41331);
nand U42390 (N_42390,N_41244,N_41383);
and U42391 (N_42391,N_41296,N_41113);
or U42392 (N_42392,N_41292,N_41427);
nor U42393 (N_42393,N_41375,N_41468);
or U42394 (N_42394,N_41828,N_41432);
and U42395 (N_42395,N_41942,N_41486);
and U42396 (N_42396,N_41656,N_41216);
nor U42397 (N_42397,N_41403,N_41876);
xnor U42398 (N_42398,N_41014,N_41962);
and U42399 (N_42399,N_41012,N_41783);
or U42400 (N_42400,N_41477,N_41785);
and U42401 (N_42401,N_41259,N_41286);
xnor U42402 (N_42402,N_41280,N_41741);
or U42403 (N_42403,N_41424,N_41911);
xor U42404 (N_42404,N_41206,N_41966);
xor U42405 (N_42405,N_41845,N_41961);
or U42406 (N_42406,N_41356,N_41684);
nor U42407 (N_42407,N_41175,N_41398);
xnor U42408 (N_42408,N_41344,N_41454);
nand U42409 (N_42409,N_41568,N_41519);
nand U42410 (N_42410,N_41917,N_41569);
nand U42411 (N_42411,N_41369,N_41699);
and U42412 (N_42412,N_41058,N_41694);
xnor U42413 (N_42413,N_41119,N_41617);
xnor U42414 (N_42414,N_41816,N_41882);
nor U42415 (N_42415,N_41578,N_41475);
or U42416 (N_42416,N_41550,N_41203);
or U42417 (N_42417,N_41459,N_41956);
nand U42418 (N_42418,N_41909,N_41440);
and U42419 (N_42419,N_41147,N_41593);
and U42420 (N_42420,N_41160,N_41696);
or U42421 (N_42421,N_41721,N_41608);
nor U42422 (N_42422,N_41573,N_41428);
nor U42423 (N_42423,N_41765,N_41315);
nand U42424 (N_42424,N_41992,N_41597);
nand U42425 (N_42425,N_41614,N_41674);
or U42426 (N_42426,N_41938,N_41928);
nor U42427 (N_42427,N_41163,N_41016);
nand U42428 (N_42428,N_41473,N_41417);
nand U42429 (N_42429,N_41756,N_41368);
or U42430 (N_42430,N_41530,N_41072);
xor U42431 (N_42431,N_41461,N_41893);
nor U42432 (N_42432,N_41236,N_41869);
and U42433 (N_42433,N_41003,N_41196);
and U42434 (N_42434,N_41235,N_41531);
or U42435 (N_42435,N_41399,N_41725);
nor U42436 (N_42436,N_41618,N_41735);
or U42437 (N_42437,N_41554,N_41258);
or U42438 (N_42438,N_41766,N_41733);
nor U42439 (N_42439,N_41410,N_41269);
xor U42440 (N_42440,N_41881,N_41346);
or U42441 (N_42441,N_41835,N_41812);
and U42442 (N_42442,N_41511,N_41524);
or U42443 (N_42443,N_41479,N_41330);
xnor U42444 (N_42444,N_41598,N_41877);
xor U42445 (N_42445,N_41743,N_41273);
and U42446 (N_42446,N_41861,N_41886);
nor U42447 (N_42447,N_41283,N_41852);
and U42448 (N_42448,N_41939,N_41698);
and U42449 (N_42449,N_41376,N_41703);
and U42450 (N_42450,N_41669,N_41122);
nor U42451 (N_42451,N_41159,N_41055);
or U42452 (N_42452,N_41004,N_41272);
nor U42453 (N_42453,N_41640,N_41224);
nor U42454 (N_42454,N_41539,N_41389);
or U42455 (N_42455,N_41397,N_41553);
and U42456 (N_42456,N_41130,N_41215);
or U42457 (N_42457,N_41182,N_41437);
and U42458 (N_42458,N_41228,N_41522);
and U42459 (N_42459,N_41471,N_41152);
nand U42460 (N_42460,N_41644,N_41316);
or U42461 (N_42461,N_41859,N_41008);
nor U42462 (N_42462,N_41527,N_41350);
nor U42463 (N_42463,N_41103,N_41896);
or U42464 (N_42464,N_41746,N_41023);
and U42465 (N_42465,N_41171,N_41918);
and U42466 (N_42466,N_41046,N_41352);
xnor U42467 (N_42467,N_41815,N_41451);
xor U42468 (N_42468,N_41803,N_41858);
nor U42469 (N_42469,N_41891,N_41865);
nor U42470 (N_42470,N_41198,N_41457);
xnor U42471 (N_42471,N_41857,N_41423);
nor U42472 (N_42472,N_41564,N_41181);
and U42473 (N_42473,N_41116,N_41724);
nor U42474 (N_42474,N_41384,N_41000);
nor U42475 (N_42475,N_41118,N_41604);
nor U42476 (N_42476,N_41456,N_41579);
and U42477 (N_42477,N_41408,N_41888);
or U42478 (N_42478,N_41978,N_41484);
nor U42479 (N_42479,N_41720,N_41708);
and U42480 (N_42480,N_41650,N_41448);
and U42481 (N_42481,N_41991,N_41793);
xnor U42482 (N_42482,N_41653,N_41637);
xor U42483 (N_42483,N_41827,N_41179);
nand U42484 (N_42484,N_41959,N_41853);
nor U42485 (N_42485,N_41419,N_41436);
and U42486 (N_42486,N_41601,N_41009);
and U42487 (N_42487,N_41649,N_41890);
xnor U42488 (N_42488,N_41801,N_41343);
or U42489 (N_42489,N_41693,N_41651);
nand U42490 (N_42490,N_41390,N_41867);
xor U42491 (N_42491,N_41345,N_41268);
and U42492 (N_42492,N_41237,N_41061);
nor U42493 (N_42493,N_41311,N_41904);
nor U42494 (N_42494,N_41469,N_41267);
nand U42495 (N_42495,N_41560,N_41589);
or U42496 (N_42496,N_41164,N_41155);
xnor U42497 (N_42497,N_41412,N_41570);
or U42498 (N_42498,N_41712,N_41872);
and U42499 (N_42499,N_41713,N_41677);
and U42500 (N_42500,N_41834,N_41066);
and U42501 (N_42501,N_41189,N_41182);
nand U42502 (N_42502,N_41951,N_41566);
nand U42503 (N_42503,N_41250,N_41483);
xor U42504 (N_42504,N_41513,N_41664);
or U42505 (N_42505,N_41098,N_41091);
xnor U42506 (N_42506,N_41569,N_41857);
or U42507 (N_42507,N_41243,N_41305);
xor U42508 (N_42508,N_41126,N_41072);
nand U42509 (N_42509,N_41741,N_41927);
xor U42510 (N_42510,N_41703,N_41454);
or U42511 (N_42511,N_41080,N_41635);
xnor U42512 (N_42512,N_41303,N_41349);
or U42513 (N_42513,N_41997,N_41015);
and U42514 (N_42514,N_41397,N_41943);
xnor U42515 (N_42515,N_41601,N_41905);
xor U42516 (N_42516,N_41266,N_41950);
or U42517 (N_42517,N_41515,N_41675);
nand U42518 (N_42518,N_41945,N_41716);
and U42519 (N_42519,N_41139,N_41991);
xor U42520 (N_42520,N_41520,N_41243);
or U42521 (N_42521,N_41530,N_41893);
nor U42522 (N_42522,N_41441,N_41466);
nor U42523 (N_42523,N_41499,N_41091);
nand U42524 (N_42524,N_41112,N_41743);
nand U42525 (N_42525,N_41784,N_41380);
or U42526 (N_42526,N_41080,N_41242);
nor U42527 (N_42527,N_41152,N_41617);
or U42528 (N_42528,N_41487,N_41530);
nand U42529 (N_42529,N_41940,N_41329);
or U42530 (N_42530,N_41945,N_41620);
or U42531 (N_42531,N_41530,N_41736);
or U42532 (N_42532,N_41529,N_41730);
and U42533 (N_42533,N_41818,N_41790);
xor U42534 (N_42534,N_41516,N_41367);
nand U42535 (N_42535,N_41076,N_41961);
and U42536 (N_42536,N_41434,N_41515);
or U42537 (N_42537,N_41867,N_41238);
or U42538 (N_42538,N_41495,N_41162);
nand U42539 (N_42539,N_41474,N_41371);
xor U42540 (N_42540,N_41470,N_41751);
nand U42541 (N_42541,N_41710,N_41033);
or U42542 (N_42542,N_41656,N_41979);
nor U42543 (N_42543,N_41539,N_41342);
or U42544 (N_42544,N_41937,N_41608);
nand U42545 (N_42545,N_41080,N_41201);
and U42546 (N_42546,N_41086,N_41513);
and U42547 (N_42547,N_41787,N_41661);
xor U42548 (N_42548,N_41303,N_41131);
and U42549 (N_42549,N_41381,N_41186);
or U42550 (N_42550,N_41085,N_41484);
xnor U42551 (N_42551,N_41444,N_41458);
nor U42552 (N_42552,N_41099,N_41137);
and U42553 (N_42553,N_41501,N_41552);
nand U42554 (N_42554,N_41914,N_41750);
nand U42555 (N_42555,N_41020,N_41396);
xnor U42556 (N_42556,N_41989,N_41869);
or U42557 (N_42557,N_41534,N_41999);
and U42558 (N_42558,N_41299,N_41816);
xnor U42559 (N_42559,N_41471,N_41123);
and U42560 (N_42560,N_41057,N_41138);
nor U42561 (N_42561,N_41333,N_41259);
nand U42562 (N_42562,N_41496,N_41271);
nand U42563 (N_42563,N_41615,N_41768);
and U42564 (N_42564,N_41697,N_41476);
nor U42565 (N_42565,N_41053,N_41876);
nand U42566 (N_42566,N_41514,N_41090);
nand U42567 (N_42567,N_41667,N_41973);
nor U42568 (N_42568,N_41342,N_41398);
xor U42569 (N_42569,N_41235,N_41511);
or U42570 (N_42570,N_41039,N_41467);
nand U42571 (N_42571,N_41963,N_41585);
and U42572 (N_42572,N_41350,N_41335);
nor U42573 (N_42573,N_41297,N_41984);
and U42574 (N_42574,N_41827,N_41310);
or U42575 (N_42575,N_41504,N_41225);
and U42576 (N_42576,N_41285,N_41478);
nor U42577 (N_42577,N_41925,N_41230);
nand U42578 (N_42578,N_41332,N_41142);
or U42579 (N_42579,N_41226,N_41560);
nand U42580 (N_42580,N_41696,N_41586);
nor U42581 (N_42581,N_41708,N_41963);
nor U42582 (N_42582,N_41197,N_41294);
and U42583 (N_42583,N_41831,N_41282);
and U42584 (N_42584,N_41952,N_41614);
nor U42585 (N_42585,N_41978,N_41238);
xnor U42586 (N_42586,N_41520,N_41007);
xnor U42587 (N_42587,N_41388,N_41509);
nor U42588 (N_42588,N_41593,N_41817);
and U42589 (N_42589,N_41428,N_41343);
nand U42590 (N_42590,N_41128,N_41571);
or U42591 (N_42591,N_41351,N_41084);
and U42592 (N_42592,N_41518,N_41857);
and U42593 (N_42593,N_41036,N_41502);
or U42594 (N_42594,N_41170,N_41095);
xor U42595 (N_42595,N_41542,N_41073);
and U42596 (N_42596,N_41059,N_41089);
nand U42597 (N_42597,N_41758,N_41755);
and U42598 (N_42598,N_41060,N_41031);
or U42599 (N_42599,N_41256,N_41224);
or U42600 (N_42600,N_41222,N_41136);
xnor U42601 (N_42601,N_41328,N_41437);
and U42602 (N_42602,N_41920,N_41489);
and U42603 (N_42603,N_41237,N_41977);
and U42604 (N_42604,N_41174,N_41004);
nor U42605 (N_42605,N_41621,N_41198);
nor U42606 (N_42606,N_41208,N_41790);
nand U42607 (N_42607,N_41245,N_41832);
xnor U42608 (N_42608,N_41032,N_41730);
nand U42609 (N_42609,N_41019,N_41591);
xnor U42610 (N_42610,N_41040,N_41485);
nand U42611 (N_42611,N_41836,N_41430);
nor U42612 (N_42612,N_41757,N_41945);
nor U42613 (N_42613,N_41386,N_41884);
or U42614 (N_42614,N_41006,N_41096);
or U42615 (N_42615,N_41082,N_41677);
and U42616 (N_42616,N_41133,N_41072);
or U42617 (N_42617,N_41177,N_41022);
nand U42618 (N_42618,N_41944,N_41293);
or U42619 (N_42619,N_41954,N_41121);
xnor U42620 (N_42620,N_41988,N_41715);
xnor U42621 (N_42621,N_41224,N_41965);
or U42622 (N_42622,N_41504,N_41460);
xnor U42623 (N_42623,N_41494,N_41144);
xnor U42624 (N_42624,N_41675,N_41064);
or U42625 (N_42625,N_41996,N_41733);
nor U42626 (N_42626,N_41178,N_41281);
or U42627 (N_42627,N_41624,N_41457);
and U42628 (N_42628,N_41193,N_41167);
nand U42629 (N_42629,N_41967,N_41379);
nor U42630 (N_42630,N_41299,N_41496);
xnor U42631 (N_42631,N_41919,N_41781);
nand U42632 (N_42632,N_41669,N_41170);
or U42633 (N_42633,N_41779,N_41404);
nor U42634 (N_42634,N_41755,N_41975);
nor U42635 (N_42635,N_41850,N_41958);
or U42636 (N_42636,N_41075,N_41887);
xnor U42637 (N_42637,N_41838,N_41922);
and U42638 (N_42638,N_41259,N_41636);
or U42639 (N_42639,N_41119,N_41797);
xnor U42640 (N_42640,N_41709,N_41875);
and U42641 (N_42641,N_41492,N_41483);
nand U42642 (N_42642,N_41504,N_41657);
xor U42643 (N_42643,N_41273,N_41194);
and U42644 (N_42644,N_41437,N_41649);
or U42645 (N_42645,N_41141,N_41406);
or U42646 (N_42646,N_41591,N_41244);
xor U42647 (N_42647,N_41814,N_41029);
or U42648 (N_42648,N_41135,N_41550);
nand U42649 (N_42649,N_41526,N_41571);
and U42650 (N_42650,N_41438,N_41480);
xnor U42651 (N_42651,N_41792,N_41472);
nor U42652 (N_42652,N_41608,N_41216);
xnor U42653 (N_42653,N_41229,N_41447);
nor U42654 (N_42654,N_41786,N_41029);
nor U42655 (N_42655,N_41026,N_41022);
xor U42656 (N_42656,N_41309,N_41906);
nand U42657 (N_42657,N_41635,N_41312);
nand U42658 (N_42658,N_41222,N_41974);
nor U42659 (N_42659,N_41576,N_41916);
nand U42660 (N_42660,N_41807,N_41015);
or U42661 (N_42661,N_41672,N_41394);
or U42662 (N_42662,N_41810,N_41001);
xor U42663 (N_42663,N_41140,N_41933);
nand U42664 (N_42664,N_41942,N_41972);
nor U42665 (N_42665,N_41727,N_41333);
xnor U42666 (N_42666,N_41685,N_41011);
nand U42667 (N_42667,N_41867,N_41421);
nand U42668 (N_42668,N_41311,N_41280);
xor U42669 (N_42669,N_41854,N_41389);
and U42670 (N_42670,N_41531,N_41001);
nor U42671 (N_42671,N_41765,N_41970);
or U42672 (N_42672,N_41406,N_41033);
and U42673 (N_42673,N_41706,N_41013);
and U42674 (N_42674,N_41866,N_41435);
and U42675 (N_42675,N_41755,N_41317);
xnor U42676 (N_42676,N_41954,N_41762);
nand U42677 (N_42677,N_41266,N_41987);
nor U42678 (N_42678,N_41539,N_41680);
and U42679 (N_42679,N_41581,N_41218);
nor U42680 (N_42680,N_41274,N_41555);
and U42681 (N_42681,N_41081,N_41553);
xnor U42682 (N_42682,N_41342,N_41049);
nor U42683 (N_42683,N_41495,N_41360);
xor U42684 (N_42684,N_41671,N_41865);
or U42685 (N_42685,N_41531,N_41156);
and U42686 (N_42686,N_41218,N_41150);
or U42687 (N_42687,N_41666,N_41370);
and U42688 (N_42688,N_41375,N_41401);
nand U42689 (N_42689,N_41482,N_41084);
xnor U42690 (N_42690,N_41644,N_41155);
or U42691 (N_42691,N_41117,N_41388);
and U42692 (N_42692,N_41619,N_41789);
xnor U42693 (N_42693,N_41457,N_41492);
nor U42694 (N_42694,N_41697,N_41012);
nand U42695 (N_42695,N_41864,N_41725);
nand U42696 (N_42696,N_41680,N_41177);
or U42697 (N_42697,N_41648,N_41694);
or U42698 (N_42698,N_41118,N_41783);
xor U42699 (N_42699,N_41320,N_41868);
or U42700 (N_42700,N_41487,N_41733);
or U42701 (N_42701,N_41135,N_41310);
nor U42702 (N_42702,N_41251,N_41243);
xnor U42703 (N_42703,N_41428,N_41394);
nand U42704 (N_42704,N_41919,N_41787);
nor U42705 (N_42705,N_41367,N_41589);
xnor U42706 (N_42706,N_41633,N_41266);
xor U42707 (N_42707,N_41971,N_41359);
or U42708 (N_42708,N_41768,N_41427);
or U42709 (N_42709,N_41659,N_41827);
or U42710 (N_42710,N_41219,N_41311);
nor U42711 (N_42711,N_41048,N_41605);
xnor U42712 (N_42712,N_41882,N_41340);
nand U42713 (N_42713,N_41608,N_41289);
or U42714 (N_42714,N_41748,N_41202);
or U42715 (N_42715,N_41033,N_41512);
xnor U42716 (N_42716,N_41537,N_41639);
nor U42717 (N_42717,N_41007,N_41035);
or U42718 (N_42718,N_41444,N_41582);
or U42719 (N_42719,N_41456,N_41000);
or U42720 (N_42720,N_41340,N_41993);
and U42721 (N_42721,N_41513,N_41310);
nand U42722 (N_42722,N_41322,N_41724);
xnor U42723 (N_42723,N_41672,N_41907);
nor U42724 (N_42724,N_41614,N_41898);
nand U42725 (N_42725,N_41695,N_41575);
xnor U42726 (N_42726,N_41699,N_41411);
and U42727 (N_42727,N_41037,N_41587);
nand U42728 (N_42728,N_41830,N_41465);
nand U42729 (N_42729,N_41869,N_41661);
nor U42730 (N_42730,N_41641,N_41199);
and U42731 (N_42731,N_41423,N_41925);
xor U42732 (N_42732,N_41611,N_41837);
xnor U42733 (N_42733,N_41195,N_41312);
or U42734 (N_42734,N_41675,N_41570);
nor U42735 (N_42735,N_41154,N_41365);
nand U42736 (N_42736,N_41279,N_41501);
or U42737 (N_42737,N_41470,N_41172);
nor U42738 (N_42738,N_41383,N_41176);
and U42739 (N_42739,N_41942,N_41702);
and U42740 (N_42740,N_41904,N_41441);
xor U42741 (N_42741,N_41803,N_41180);
and U42742 (N_42742,N_41347,N_41353);
xor U42743 (N_42743,N_41313,N_41116);
or U42744 (N_42744,N_41340,N_41326);
nor U42745 (N_42745,N_41148,N_41119);
nand U42746 (N_42746,N_41576,N_41502);
nand U42747 (N_42747,N_41100,N_41973);
xor U42748 (N_42748,N_41318,N_41063);
nand U42749 (N_42749,N_41863,N_41883);
nand U42750 (N_42750,N_41954,N_41056);
and U42751 (N_42751,N_41579,N_41947);
nand U42752 (N_42752,N_41837,N_41250);
nand U42753 (N_42753,N_41254,N_41166);
or U42754 (N_42754,N_41469,N_41819);
or U42755 (N_42755,N_41523,N_41538);
or U42756 (N_42756,N_41827,N_41271);
and U42757 (N_42757,N_41751,N_41228);
xnor U42758 (N_42758,N_41386,N_41188);
or U42759 (N_42759,N_41239,N_41163);
nand U42760 (N_42760,N_41997,N_41096);
nand U42761 (N_42761,N_41133,N_41963);
or U42762 (N_42762,N_41189,N_41299);
or U42763 (N_42763,N_41254,N_41232);
xor U42764 (N_42764,N_41748,N_41024);
or U42765 (N_42765,N_41709,N_41462);
xnor U42766 (N_42766,N_41524,N_41545);
and U42767 (N_42767,N_41526,N_41539);
xnor U42768 (N_42768,N_41370,N_41121);
or U42769 (N_42769,N_41330,N_41280);
xnor U42770 (N_42770,N_41943,N_41343);
nand U42771 (N_42771,N_41578,N_41723);
xor U42772 (N_42772,N_41368,N_41634);
nand U42773 (N_42773,N_41637,N_41687);
nand U42774 (N_42774,N_41987,N_41989);
and U42775 (N_42775,N_41895,N_41891);
or U42776 (N_42776,N_41026,N_41032);
nand U42777 (N_42777,N_41589,N_41363);
or U42778 (N_42778,N_41180,N_41451);
or U42779 (N_42779,N_41179,N_41918);
nand U42780 (N_42780,N_41352,N_41557);
and U42781 (N_42781,N_41707,N_41061);
and U42782 (N_42782,N_41917,N_41852);
nand U42783 (N_42783,N_41231,N_41426);
xor U42784 (N_42784,N_41285,N_41714);
xnor U42785 (N_42785,N_41068,N_41268);
nor U42786 (N_42786,N_41493,N_41188);
nor U42787 (N_42787,N_41083,N_41305);
nor U42788 (N_42788,N_41294,N_41014);
and U42789 (N_42789,N_41320,N_41144);
nand U42790 (N_42790,N_41610,N_41992);
and U42791 (N_42791,N_41228,N_41153);
nor U42792 (N_42792,N_41469,N_41489);
or U42793 (N_42793,N_41571,N_41455);
or U42794 (N_42794,N_41924,N_41176);
and U42795 (N_42795,N_41976,N_41480);
xnor U42796 (N_42796,N_41178,N_41001);
nand U42797 (N_42797,N_41903,N_41289);
xnor U42798 (N_42798,N_41029,N_41535);
nor U42799 (N_42799,N_41470,N_41968);
nor U42800 (N_42800,N_41777,N_41802);
nor U42801 (N_42801,N_41593,N_41581);
nor U42802 (N_42802,N_41360,N_41773);
xor U42803 (N_42803,N_41763,N_41433);
and U42804 (N_42804,N_41807,N_41153);
and U42805 (N_42805,N_41626,N_41885);
and U42806 (N_42806,N_41737,N_41153);
nand U42807 (N_42807,N_41283,N_41187);
and U42808 (N_42808,N_41022,N_41839);
nand U42809 (N_42809,N_41713,N_41380);
or U42810 (N_42810,N_41663,N_41224);
nand U42811 (N_42811,N_41563,N_41037);
nand U42812 (N_42812,N_41875,N_41128);
nor U42813 (N_42813,N_41655,N_41803);
nor U42814 (N_42814,N_41714,N_41732);
xnor U42815 (N_42815,N_41291,N_41874);
xor U42816 (N_42816,N_41879,N_41730);
and U42817 (N_42817,N_41169,N_41689);
xnor U42818 (N_42818,N_41166,N_41082);
nor U42819 (N_42819,N_41099,N_41612);
nor U42820 (N_42820,N_41191,N_41561);
nand U42821 (N_42821,N_41129,N_41849);
and U42822 (N_42822,N_41519,N_41309);
xnor U42823 (N_42823,N_41147,N_41764);
and U42824 (N_42824,N_41062,N_41179);
and U42825 (N_42825,N_41017,N_41344);
nor U42826 (N_42826,N_41199,N_41820);
or U42827 (N_42827,N_41864,N_41055);
nor U42828 (N_42828,N_41523,N_41594);
nand U42829 (N_42829,N_41884,N_41937);
nor U42830 (N_42830,N_41423,N_41160);
nor U42831 (N_42831,N_41680,N_41311);
xor U42832 (N_42832,N_41525,N_41696);
nand U42833 (N_42833,N_41207,N_41808);
nand U42834 (N_42834,N_41916,N_41154);
nand U42835 (N_42835,N_41226,N_41649);
or U42836 (N_42836,N_41537,N_41319);
nand U42837 (N_42837,N_41983,N_41158);
xor U42838 (N_42838,N_41766,N_41746);
or U42839 (N_42839,N_41486,N_41868);
or U42840 (N_42840,N_41645,N_41632);
nand U42841 (N_42841,N_41086,N_41200);
and U42842 (N_42842,N_41562,N_41901);
nand U42843 (N_42843,N_41701,N_41510);
nand U42844 (N_42844,N_41176,N_41352);
nor U42845 (N_42845,N_41136,N_41916);
or U42846 (N_42846,N_41635,N_41704);
or U42847 (N_42847,N_41513,N_41809);
or U42848 (N_42848,N_41707,N_41197);
nor U42849 (N_42849,N_41011,N_41532);
and U42850 (N_42850,N_41803,N_41834);
nand U42851 (N_42851,N_41996,N_41377);
xnor U42852 (N_42852,N_41786,N_41708);
nor U42853 (N_42853,N_41925,N_41394);
nor U42854 (N_42854,N_41608,N_41572);
and U42855 (N_42855,N_41842,N_41208);
and U42856 (N_42856,N_41002,N_41222);
nor U42857 (N_42857,N_41416,N_41389);
and U42858 (N_42858,N_41714,N_41828);
or U42859 (N_42859,N_41541,N_41634);
or U42860 (N_42860,N_41056,N_41434);
nand U42861 (N_42861,N_41888,N_41710);
or U42862 (N_42862,N_41348,N_41617);
nor U42863 (N_42863,N_41235,N_41351);
and U42864 (N_42864,N_41823,N_41025);
nand U42865 (N_42865,N_41104,N_41051);
nand U42866 (N_42866,N_41540,N_41601);
xnor U42867 (N_42867,N_41947,N_41793);
xor U42868 (N_42868,N_41889,N_41619);
or U42869 (N_42869,N_41978,N_41151);
nor U42870 (N_42870,N_41415,N_41853);
or U42871 (N_42871,N_41510,N_41506);
xor U42872 (N_42872,N_41670,N_41584);
nand U42873 (N_42873,N_41437,N_41664);
or U42874 (N_42874,N_41459,N_41208);
xor U42875 (N_42875,N_41982,N_41824);
nand U42876 (N_42876,N_41789,N_41724);
xnor U42877 (N_42877,N_41077,N_41924);
xnor U42878 (N_42878,N_41708,N_41802);
or U42879 (N_42879,N_41464,N_41238);
and U42880 (N_42880,N_41480,N_41376);
or U42881 (N_42881,N_41626,N_41315);
nor U42882 (N_42882,N_41222,N_41042);
or U42883 (N_42883,N_41206,N_41608);
xnor U42884 (N_42884,N_41452,N_41676);
nand U42885 (N_42885,N_41284,N_41699);
or U42886 (N_42886,N_41295,N_41254);
nor U42887 (N_42887,N_41540,N_41227);
and U42888 (N_42888,N_41603,N_41425);
or U42889 (N_42889,N_41054,N_41244);
or U42890 (N_42890,N_41457,N_41377);
or U42891 (N_42891,N_41097,N_41441);
xor U42892 (N_42892,N_41023,N_41474);
or U42893 (N_42893,N_41427,N_41253);
xnor U42894 (N_42894,N_41725,N_41977);
xnor U42895 (N_42895,N_41239,N_41400);
xor U42896 (N_42896,N_41059,N_41142);
nand U42897 (N_42897,N_41267,N_41218);
or U42898 (N_42898,N_41221,N_41328);
nor U42899 (N_42899,N_41344,N_41453);
nor U42900 (N_42900,N_41742,N_41417);
or U42901 (N_42901,N_41695,N_41674);
nand U42902 (N_42902,N_41544,N_41508);
nor U42903 (N_42903,N_41332,N_41037);
and U42904 (N_42904,N_41231,N_41257);
nor U42905 (N_42905,N_41386,N_41646);
and U42906 (N_42906,N_41954,N_41897);
and U42907 (N_42907,N_41453,N_41100);
nand U42908 (N_42908,N_41031,N_41249);
and U42909 (N_42909,N_41161,N_41263);
or U42910 (N_42910,N_41162,N_41941);
xnor U42911 (N_42911,N_41568,N_41763);
nor U42912 (N_42912,N_41142,N_41464);
and U42913 (N_42913,N_41621,N_41692);
or U42914 (N_42914,N_41570,N_41797);
nand U42915 (N_42915,N_41235,N_41372);
nor U42916 (N_42916,N_41729,N_41401);
nand U42917 (N_42917,N_41032,N_41666);
and U42918 (N_42918,N_41469,N_41754);
nand U42919 (N_42919,N_41042,N_41170);
or U42920 (N_42920,N_41876,N_41084);
nor U42921 (N_42921,N_41855,N_41876);
nor U42922 (N_42922,N_41237,N_41436);
and U42923 (N_42923,N_41240,N_41257);
or U42924 (N_42924,N_41543,N_41225);
nand U42925 (N_42925,N_41550,N_41312);
and U42926 (N_42926,N_41969,N_41896);
and U42927 (N_42927,N_41054,N_41447);
and U42928 (N_42928,N_41338,N_41758);
xnor U42929 (N_42929,N_41159,N_41221);
or U42930 (N_42930,N_41297,N_41407);
or U42931 (N_42931,N_41400,N_41040);
nor U42932 (N_42932,N_41729,N_41145);
and U42933 (N_42933,N_41545,N_41598);
nand U42934 (N_42934,N_41853,N_41424);
nor U42935 (N_42935,N_41560,N_41617);
and U42936 (N_42936,N_41328,N_41726);
or U42937 (N_42937,N_41263,N_41567);
and U42938 (N_42938,N_41985,N_41117);
or U42939 (N_42939,N_41185,N_41301);
xnor U42940 (N_42940,N_41297,N_41508);
and U42941 (N_42941,N_41020,N_41308);
xnor U42942 (N_42942,N_41086,N_41483);
and U42943 (N_42943,N_41540,N_41798);
and U42944 (N_42944,N_41881,N_41517);
nand U42945 (N_42945,N_41586,N_41658);
nand U42946 (N_42946,N_41150,N_41566);
xnor U42947 (N_42947,N_41332,N_41981);
nor U42948 (N_42948,N_41353,N_41228);
nand U42949 (N_42949,N_41448,N_41496);
xnor U42950 (N_42950,N_41856,N_41138);
nor U42951 (N_42951,N_41063,N_41431);
nor U42952 (N_42952,N_41736,N_41402);
xnor U42953 (N_42953,N_41281,N_41587);
nand U42954 (N_42954,N_41795,N_41916);
nand U42955 (N_42955,N_41100,N_41780);
xor U42956 (N_42956,N_41023,N_41569);
or U42957 (N_42957,N_41963,N_41473);
xor U42958 (N_42958,N_41393,N_41913);
and U42959 (N_42959,N_41762,N_41385);
and U42960 (N_42960,N_41157,N_41675);
or U42961 (N_42961,N_41321,N_41491);
and U42962 (N_42962,N_41237,N_41894);
nor U42963 (N_42963,N_41034,N_41122);
or U42964 (N_42964,N_41731,N_41015);
xnor U42965 (N_42965,N_41870,N_41808);
xnor U42966 (N_42966,N_41247,N_41138);
nor U42967 (N_42967,N_41998,N_41669);
xnor U42968 (N_42968,N_41921,N_41696);
or U42969 (N_42969,N_41149,N_41568);
or U42970 (N_42970,N_41682,N_41371);
or U42971 (N_42971,N_41635,N_41902);
or U42972 (N_42972,N_41169,N_41589);
or U42973 (N_42973,N_41241,N_41369);
xor U42974 (N_42974,N_41673,N_41442);
or U42975 (N_42975,N_41587,N_41523);
nor U42976 (N_42976,N_41576,N_41738);
xnor U42977 (N_42977,N_41401,N_41188);
or U42978 (N_42978,N_41009,N_41166);
nand U42979 (N_42979,N_41052,N_41268);
xnor U42980 (N_42980,N_41619,N_41667);
or U42981 (N_42981,N_41657,N_41572);
nand U42982 (N_42982,N_41498,N_41448);
or U42983 (N_42983,N_41543,N_41756);
nor U42984 (N_42984,N_41250,N_41018);
xnor U42985 (N_42985,N_41633,N_41041);
and U42986 (N_42986,N_41966,N_41743);
and U42987 (N_42987,N_41637,N_41904);
nand U42988 (N_42988,N_41203,N_41128);
nand U42989 (N_42989,N_41018,N_41144);
or U42990 (N_42990,N_41888,N_41663);
xnor U42991 (N_42991,N_41476,N_41893);
or U42992 (N_42992,N_41730,N_41192);
and U42993 (N_42993,N_41551,N_41433);
or U42994 (N_42994,N_41998,N_41996);
or U42995 (N_42995,N_41047,N_41642);
or U42996 (N_42996,N_41782,N_41528);
xnor U42997 (N_42997,N_41949,N_41635);
and U42998 (N_42998,N_41507,N_41617);
nor U42999 (N_42999,N_41953,N_41260);
nor U43000 (N_43000,N_42264,N_42063);
and U43001 (N_43001,N_42571,N_42251);
and U43002 (N_43002,N_42947,N_42411);
and U43003 (N_43003,N_42835,N_42305);
nor U43004 (N_43004,N_42952,N_42638);
nor U43005 (N_43005,N_42909,N_42170);
nand U43006 (N_43006,N_42678,N_42279);
nand U43007 (N_43007,N_42395,N_42373);
or U43008 (N_43008,N_42477,N_42957);
and U43009 (N_43009,N_42766,N_42345);
or U43010 (N_43010,N_42534,N_42507);
xnor U43011 (N_43011,N_42794,N_42203);
nor U43012 (N_43012,N_42996,N_42245);
and U43013 (N_43013,N_42887,N_42662);
xor U43014 (N_43014,N_42030,N_42595);
and U43015 (N_43015,N_42764,N_42856);
nor U43016 (N_43016,N_42554,N_42062);
nor U43017 (N_43017,N_42441,N_42017);
nor U43018 (N_43018,N_42447,N_42162);
or U43019 (N_43019,N_42043,N_42734);
or U43020 (N_43020,N_42956,N_42562);
nand U43021 (N_43021,N_42448,N_42701);
nor U43022 (N_43022,N_42895,N_42605);
nand U43023 (N_43023,N_42616,N_42660);
or U43024 (N_43024,N_42904,N_42212);
nor U43025 (N_43025,N_42682,N_42827);
nor U43026 (N_43026,N_42593,N_42387);
nor U43027 (N_43027,N_42284,N_42500);
and U43028 (N_43028,N_42729,N_42445);
or U43029 (N_43029,N_42304,N_42107);
xnor U43030 (N_43030,N_42462,N_42153);
nor U43031 (N_43031,N_42992,N_42749);
and U43032 (N_43032,N_42903,N_42070);
nor U43033 (N_43033,N_42577,N_42006);
nand U43034 (N_43034,N_42053,N_42287);
or U43035 (N_43035,N_42988,N_42491);
nand U43036 (N_43036,N_42423,N_42647);
nand U43037 (N_43037,N_42602,N_42514);
and U43038 (N_43038,N_42269,N_42843);
xor U43039 (N_43039,N_42228,N_42220);
or U43040 (N_43040,N_42041,N_42513);
nor U43041 (N_43041,N_42670,N_42855);
and U43042 (N_43042,N_42607,N_42922);
nor U43043 (N_43043,N_42389,N_42669);
xnor U43044 (N_43044,N_42675,N_42710);
xnor U43045 (N_43045,N_42780,N_42049);
nor U43046 (N_43046,N_42892,N_42092);
nor U43047 (N_43047,N_42340,N_42591);
nand U43048 (N_43048,N_42801,N_42680);
and U43049 (N_43049,N_42972,N_42370);
or U43050 (N_43050,N_42074,N_42271);
or U43051 (N_43051,N_42350,N_42531);
and U43052 (N_43052,N_42820,N_42257);
or U43053 (N_43053,N_42005,N_42886);
nand U43054 (N_43054,N_42981,N_42024);
nand U43055 (N_43055,N_42877,N_42526);
xor U43056 (N_43056,N_42243,N_42953);
nand U43057 (N_43057,N_42560,N_42103);
nor U43058 (N_43058,N_42578,N_42424);
nor U43059 (N_43059,N_42604,N_42708);
nor U43060 (N_43060,N_42376,N_42367);
xnor U43061 (N_43061,N_42803,N_42382);
and U43062 (N_43062,N_42893,N_42664);
nor U43063 (N_43063,N_42108,N_42214);
and U43064 (N_43064,N_42480,N_42036);
nand U43065 (N_43065,N_42700,N_42039);
nor U43066 (N_43066,N_42880,N_42227);
nor U43067 (N_43067,N_42949,N_42038);
nand U43068 (N_43068,N_42505,N_42207);
nor U43069 (N_43069,N_42929,N_42589);
or U43070 (N_43070,N_42289,N_42584);
nor U43071 (N_43071,N_42319,N_42672);
xnor U43072 (N_43072,N_42961,N_42774);
nand U43073 (N_43073,N_42919,N_42649);
nand U43074 (N_43074,N_42733,N_42113);
or U43075 (N_43075,N_42739,N_42658);
nor U43076 (N_43076,N_42335,N_42252);
and U43077 (N_43077,N_42709,N_42457);
xnor U43078 (N_43078,N_42550,N_42191);
and U43079 (N_43079,N_42202,N_42366);
nor U43080 (N_43080,N_42555,N_42283);
nor U43081 (N_43081,N_42330,N_42422);
xor U43082 (N_43082,N_42337,N_42781);
or U43083 (N_43083,N_42438,N_42426);
nor U43084 (N_43084,N_42194,N_42711);
xor U43085 (N_43085,N_42322,N_42148);
nor U43086 (N_43086,N_42506,N_42280);
xnor U43087 (N_43087,N_42659,N_42222);
nor U43088 (N_43088,N_42008,N_42580);
nand U43089 (N_43089,N_42343,N_42421);
or U43090 (N_43090,N_42095,N_42752);
nand U43091 (N_43091,N_42718,N_42540);
or U43092 (N_43092,N_42090,N_42631);
nand U43093 (N_43093,N_42233,N_42535);
and U43094 (N_43094,N_42529,N_42465);
or U43095 (N_43095,N_42692,N_42303);
and U43096 (N_43096,N_42863,N_42037);
or U43097 (N_43097,N_42104,N_42695);
and U43098 (N_43098,N_42282,N_42728);
and U43099 (N_43099,N_42862,N_42163);
xnor U43100 (N_43100,N_42768,N_42634);
or U43101 (N_43101,N_42374,N_42481);
nand U43102 (N_43102,N_42861,N_42434);
xnor U43103 (N_43103,N_42045,N_42564);
and U43104 (N_43104,N_42250,N_42157);
xnor U43105 (N_43105,N_42727,N_42516);
or U43106 (N_43106,N_42991,N_42115);
nand U43107 (N_43107,N_42548,N_42750);
or U43108 (N_43108,N_42181,N_42811);
or U43109 (N_43109,N_42642,N_42574);
or U43110 (N_43110,N_42489,N_42666);
and U43111 (N_43111,N_42042,N_42152);
or U43112 (N_43112,N_42690,N_42779);
or U43113 (N_43113,N_42351,N_42195);
or U43114 (N_43114,N_42380,N_42312);
nand U43115 (N_43115,N_42263,N_42234);
xnor U43116 (N_43116,N_42760,N_42939);
and U43117 (N_43117,N_42098,N_42132);
and U43118 (N_43118,N_42703,N_42427);
nor U43119 (N_43119,N_42393,N_42072);
and U43120 (N_43120,N_42783,N_42479);
or U43121 (N_43121,N_42379,N_42874);
or U43122 (N_43122,N_42353,N_42256);
nor U43123 (N_43123,N_42915,N_42511);
or U43124 (N_43124,N_42001,N_42192);
nor U43125 (N_43125,N_42297,N_42354);
nor U43126 (N_43126,N_42216,N_42057);
or U43127 (N_43127,N_42133,N_42249);
nand U43128 (N_43128,N_42276,N_42990);
nand U43129 (N_43129,N_42224,N_42334);
nand U43130 (N_43130,N_42964,N_42097);
nor U43131 (N_43131,N_42625,N_42247);
nor U43132 (N_43132,N_42628,N_42795);
and U43133 (N_43133,N_42583,N_42646);
nor U43134 (N_43134,N_42822,N_42325);
and U43135 (N_43135,N_42211,N_42888);
nor U43136 (N_43136,N_42557,N_42410);
and U43137 (N_43137,N_42673,N_42572);
xnor U43138 (N_43138,N_42923,N_42854);
or U43139 (N_43139,N_42167,N_42873);
and U43140 (N_43140,N_42352,N_42079);
nand U43141 (N_43141,N_42911,N_42654);
and U43142 (N_43142,N_42592,N_42525);
xnor U43143 (N_43143,N_42657,N_42521);
and U43144 (N_43144,N_42492,N_42896);
xnor U43145 (N_43145,N_42890,N_42339);
nor U43146 (N_43146,N_42544,N_42897);
or U43147 (N_43147,N_42603,N_42145);
and U43148 (N_43148,N_42661,N_42016);
and U43149 (N_43149,N_42310,N_42165);
nor U43150 (N_43150,N_42720,N_42111);
and U43151 (N_43151,N_42546,N_42429);
xnor U43152 (N_43152,N_42503,N_42292);
nand U43153 (N_43153,N_42433,N_42905);
nor U43154 (N_43154,N_42139,N_42770);
nand U43155 (N_43155,N_42123,N_42937);
xnor U43156 (N_43156,N_42180,N_42117);
nand U43157 (N_43157,N_42796,N_42128);
nor U43158 (N_43158,N_42782,N_42866);
nor U43159 (N_43159,N_42771,N_42620);
xor U43160 (N_43160,N_42081,N_42294);
xor U43161 (N_43161,N_42997,N_42933);
and U43162 (N_43162,N_42528,N_42600);
or U43163 (N_43163,N_42959,N_42968);
xor U43164 (N_43164,N_42640,N_42627);
and U43165 (N_43165,N_42437,N_42813);
nor U43166 (N_43166,N_42327,N_42809);
or U43167 (N_43167,N_42118,N_42364);
or U43168 (N_43168,N_42826,N_42740);
or U43169 (N_43169,N_42934,N_42706);
xor U43170 (N_43170,N_42832,N_42808);
nand U43171 (N_43171,N_42461,N_42684);
or U43172 (N_43172,N_42597,N_42716);
nand U43173 (N_43173,N_42552,N_42587);
and U43174 (N_43174,N_42838,N_42205);
or U43175 (N_43175,N_42527,N_42231);
xnor U43176 (N_43176,N_42920,N_42935);
nor U43177 (N_43177,N_42401,N_42449);
or U43178 (N_43178,N_42260,N_42786);
xnor U43179 (N_43179,N_42792,N_42386);
nor U43180 (N_43180,N_42772,N_42825);
xor U43181 (N_43181,N_42917,N_42171);
or U43182 (N_43182,N_42463,N_42721);
or U43183 (N_43183,N_42295,N_42164);
or U43184 (N_43184,N_42056,N_42565);
nand U43185 (N_43185,N_42416,N_42044);
nor U43186 (N_43186,N_42394,N_42083);
and U43187 (N_43187,N_42026,N_42773);
nor U43188 (N_43188,N_42435,N_42836);
and U43189 (N_43189,N_42758,N_42302);
nor U43190 (N_43190,N_42160,N_42120);
nor U43191 (N_43191,N_42267,N_42306);
nor U43192 (N_43192,N_42313,N_42331);
xnor U43193 (N_43193,N_42954,N_42648);
and U43194 (N_43194,N_42136,N_42004);
and U43195 (N_43195,N_42454,N_42431);
xor U43196 (N_43196,N_42129,N_42573);
nor U43197 (N_43197,N_42459,N_42722);
and U43198 (N_43198,N_42549,N_42018);
or U43199 (N_43199,N_42847,N_42530);
nor U43200 (N_43200,N_42860,N_42409);
or U43201 (N_43201,N_42747,N_42124);
nor U43202 (N_43202,N_42293,N_42737);
nor U43203 (N_43203,N_42029,N_42439);
and U43204 (N_43204,N_42741,N_42858);
nor U43205 (N_43205,N_42109,N_42859);
or U43206 (N_43206,N_42208,N_42520);
and U43207 (N_43207,N_42408,N_42360);
nand U43208 (N_43208,N_42348,N_42980);
nor U43209 (N_43209,N_42450,N_42496);
xor U43210 (N_43210,N_42946,N_42599);
or U43211 (N_43211,N_42522,N_42715);
and U43212 (N_43212,N_42291,N_42106);
nand U43213 (N_43213,N_42196,N_42846);
or U43214 (N_43214,N_42100,N_42730);
or U43215 (N_43215,N_42080,N_42748);
xnor U43216 (N_43216,N_42144,N_42876);
nand U43217 (N_43217,N_42869,N_42432);
or U43218 (N_43218,N_42865,N_42742);
or U43219 (N_43219,N_42059,N_42501);
or U43220 (N_43220,N_42932,N_42105);
and U43221 (N_43221,N_42928,N_42912);
and U43222 (N_43222,N_42753,N_42763);
nand U43223 (N_43223,N_42576,N_42681);
nand U43224 (N_43224,N_42143,N_42891);
or U43225 (N_43225,N_42732,N_42655);
nand U43226 (N_43226,N_42842,N_42713);
nand U43227 (N_43227,N_42281,N_42135);
xor U43228 (N_43228,N_42785,N_42745);
and U43229 (N_43229,N_42615,N_42235);
xor U43230 (N_43230,N_42201,N_42907);
or U43231 (N_43231,N_42736,N_42719);
xnor U43232 (N_43232,N_42543,N_42537);
or U43233 (N_43233,N_42965,N_42702);
nor U43234 (N_43234,N_42040,N_42467);
nor U43235 (N_43235,N_42868,N_42962);
nor U43236 (N_43236,N_42391,N_42498);
xnor U43237 (N_43237,N_42582,N_42581);
nand U43238 (N_43238,N_42769,N_42242);
nand U43239 (N_43239,N_42977,N_42096);
or U43240 (N_43240,N_42641,N_42762);
nand U43241 (N_43241,N_42342,N_42472);
nand U43242 (N_43242,N_42091,N_42705);
nand U43243 (N_43243,N_42948,N_42995);
xnor U43244 (N_43244,N_42927,N_42551);
or U43245 (N_43245,N_42140,N_42332);
nor U43246 (N_43246,N_42372,N_42147);
nand U43247 (N_43247,N_42047,N_42188);
and U43248 (N_43248,N_42073,N_42324);
nand U43249 (N_43249,N_42493,N_42969);
and U43250 (N_43250,N_42320,N_42189);
or U43251 (N_43251,N_42598,N_42942);
nor U43252 (N_43252,N_42967,N_42979);
nand U43253 (N_43253,N_42093,N_42071);
nor U43254 (N_43254,N_42341,N_42226);
and U43255 (N_43255,N_42823,N_42683);
and U43256 (N_43256,N_42048,N_42914);
or U43257 (N_43257,N_42025,N_42517);
and U43258 (N_43258,N_42428,N_42679);
and U43259 (N_43259,N_42412,N_42130);
xor U43260 (N_43260,N_42687,N_42608);
nand U43261 (N_43261,N_42442,N_42588);
nand U43262 (N_43262,N_42663,N_42436);
or U43263 (N_43263,N_42755,N_42989);
or U43264 (N_43264,N_42817,N_42495);
nor U43265 (N_43265,N_42176,N_42368);
or U43266 (N_43266,N_42757,N_42206);
nand U43267 (N_43267,N_42022,N_42034);
or U43268 (N_43268,N_42767,N_42458);
or U43269 (N_43269,N_42744,N_42971);
or U43270 (N_43270,N_42329,N_42547);
or U43271 (N_43271,N_42487,N_42430);
or U43272 (N_43272,N_42694,N_42805);
nand U43273 (N_43273,N_42788,N_42221);
xnor U43274 (N_43274,N_42328,N_42689);
xnor U43275 (N_43275,N_42944,N_42926);
xnor U43276 (N_43276,N_42656,N_42898);
or U43277 (N_43277,N_42204,N_42812);
xnor U43278 (N_43278,N_42563,N_42532);
or U43279 (N_43279,N_42943,N_42168);
or U43280 (N_43280,N_42405,N_42975);
and U43281 (N_43281,N_42921,N_42845);
nor U43282 (N_43282,N_42468,N_42725);
xor U43283 (N_43283,N_42347,N_42759);
or U43284 (N_43284,N_42945,N_42173);
or U43285 (N_43285,N_42850,N_42830);
xor U43286 (N_43286,N_42955,N_42032);
and U43287 (N_43287,N_42624,N_42596);
and U43288 (N_43288,N_42629,N_42940);
and U43289 (N_43289,N_42963,N_42966);
nor U43290 (N_43290,N_42797,N_42668);
nand U43291 (N_43291,N_42166,N_42285);
nand U43292 (N_43292,N_42693,N_42613);
nand U43293 (N_43293,N_42645,N_42978);
or U43294 (N_43294,N_42985,N_42723);
nand U43295 (N_43295,N_42027,N_42262);
nor U43296 (N_43296,N_42466,N_42611);
xor U43297 (N_43297,N_42632,N_42076);
and U43298 (N_43298,N_42916,N_42483);
nand U43299 (N_43299,N_42253,N_42161);
or U43300 (N_43300,N_42307,N_42355);
and U43301 (N_43301,N_42010,N_42622);
nor U43302 (N_43302,N_42158,N_42002);
or U43303 (N_43303,N_42069,N_42390);
and U43304 (N_43304,N_42185,N_42635);
nor U43305 (N_43305,N_42538,N_42277);
and U43306 (N_43306,N_42998,N_42003);
or U43307 (N_43307,N_42743,N_42114);
nand U43308 (N_43308,N_42712,N_42137);
or U43309 (N_43309,N_42248,N_42925);
nor U43310 (N_43310,N_42035,N_42519);
xnor U43311 (N_43311,N_42504,N_42317);
xor U43312 (N_43312,N_42052,N_42831);
nand U43313 (N_43313,N_42169,N_42473);
nor U43314 (N_43314,N_42960,N_42704);
nor U43315 (N_43315,N_42088,N_42485);
xor U43316 (N_43316,N_42486,N_42901);
or U43317 (N_43317,N_42884,N_42023);
and U43318 (N_43318,N_42761,N_42218);
nand U43319 (N_43319,N_42399,N_42275);
xnor U43320 (N_43320,N_42417,N_42906);
xor U43321 (N_43321,N_42314,N_42122);
and U43322 (N_43322,N_42346,N_42545);
and U43323 (N_43323,N_42470,N_42751);
xor U43324 (N_43324,N_42879,N_42406);
and U43325 (N_43325,N_42610,N_42397);
and U43326 (N_43326,N_42902,N_42717);
nand U43327 (N_43327,N_42777,N_42614);
nor U43328 (N_43328,N_42084,N_42286);
or U43329 (N_43329,N_42033,N_42146);
or U43330 (N_43330,N_42881,N_42566);
xor U43331 (N_43331,N_42864,N_42296);
or U43332 (N_43332,N_42125,N_42951);
or U43333 (N_43333,N_42061,N_42174);
nand U43334 (N_43334,N_42046,N_42970);
or U43335 (N_43335,N_42223,N_42619);
nand U43336 (N_43336,N_42800,N_42236);
or U43337 (N_43337,N_42244,N_42403);
nand U43338 (N_43338,N_42494,N_42810);
nand U43339 (N_43339,N_42217,N_42142);
and U43340 (N_43340,N_42198,N_42400);
nand U43341 (N_43341,N_42665,N_42899);
nand U43342 (N_43342,N_42254,N_42112);
or U43343 (N_43343,N_42013,N_42308);
or U43344 (N_43344,N_42210,N_42674);
and U43345 (N_43345,N_42054,N_42315);
nand U43346 (N_43346,N_42606,N_42011);
xor U43347 (N_43347,N_42938,N_42568);
nand U43348 (N_43348,N_42579,N_42490);
xor U43349 (N_43349,N_42818,N_42478);
xor U43350 (N_43350,N_42502,N_42585);
xnor U43351 (N_43351,N_42378,N_42488);
or U43352 (N_43352,N_42425,N_42676);
and U43353 (N_43353,N_42453,N_42793);
xor U43354 (N_43354,N_42650,N_42735);
nor U43355 (N_43355,N_42311,N_42515);
nand U43356 (N_43356,N_42338,N_42802);
nand U43357 (N_43357,N_42418,N_42178);
and U43358 (N_43358,N_42184,N_42626);
and U43359 (N_43359,N_42396,N_42055);
and U43360 (N_43360,N_42357,N_42870);
nor U43361 (N_43361,N_42982,N_42193);
nor U43362 (N_43362,N_42241,N_42984);
nor U43363 (N_43363,N_42110,N_42082);
xnor U43364 (N_43364,N_42677,N_42569);
xor U43365 (N_43365,N_42950,N_42509);
or U43366 (N_43366,N_42099,N_42816);
and U43367 (N_43367,N_42958,N_42298);
nor U43368 (N_43368,N_42644,N_42882);
xor U43369 (N_43369,N_42089,N_42190);
or U43370 (N_43370,N_42398,N_42651);
and U43371 (N_43371,N_42512,N_42183);
and U43372 (N_43372,N_42561,N_42878);
and U43373 (N_43373,N_42476,N_42318);
nand U43374 (N_43374,N_42361,N_42362);
nand U43375 (N_43375,N_42617,N_42326);
nand U43376 (N_43376,N_42623,N_42219);
xor U43377 (N_43377,N_42799,N_42475);
or U43378 (N_43378,N_42238,N_42775);
or U43379 (N_43379,N_42924,N_42973);
or U43380 (N_43380,N_42413,N_42172);
and U43381 (N_43381,N_42000,N_42778);
or U43382 (N_43382,N_42134,N_42225);
and U43383 (N_43383,N_42536,N_42232);
nor U43384 (N_43384,N_42230,N_42215);
or U43385 (N_43385,N_42094,N_42829);
xor U43386 (N_43386,N_42187,N_42246);
or U43387 (N_43387,N_42154,N_42051);
xor U43388 (N_43388,N_42381,N_42848);
and U43389 (N_43389,N_42983,N_42553);
or U43390 (N_43390,N_42685,N_42075);
xnor U43391 (N_43391,N_42559,N_42363);
and U43392 (N_43392,N_42787,N_42078);
nor U43393 (N_43393,N_42844,N_42871);
nor U43394 (N_43394,N_42691,N_42857);
and U43395 (N_43395,N_42067,N_42612);
nand U43396 (N_43396,N_42474,N_42452);
or U43397 (N_43397,N_42636,N_42765);
xnor U43398 (N_43398,N_42301,N_42852);
or U43399 (N_43399,N_42804,N_42918);
and U43400 (N_43400,N_42499,N_42014);
and U43401 (N_43401,N_42375,N_42789);
or U43402 (N_43402,N_42278,N_42179);
nor U43403 (N_43403,N_42349,N_42814);
nor U43404 (N_43404,N_42265,N_42385);
and U43405 (N_43405,N_42883,N_42068);
xnor U43406 (N_43406,N_42268,N_42671);
nor U43407 (N_43407,N_42101,N_42261);
nor U43408 (N_43408,N_42446,N_42309);
or U43409 (N_43409,N_42266,N_42460);
and U43410 (N_43410,N_42159,N_42255);
or U43411 (N_43411,N_42853,N_42542);
xnor U43412 (N_43412,N_42012,N_42618);
or U43413 (N_43413,N_42533,N_42686);
or U43414 (N_43414,N_42116,N_42875);
xnor U43415 (N_43415,N_42819,N_42471);
nand U43416 (N_43416,N_42126,N_42087);
nand U43417 (N_43417,N_42455,N_42889);
nor U43418 (N_43418,N_42273,N_42894);
xor U43419 (N_43419,N_42833,N_42197);
nor U43420 (N_43420,N_42066,N_42443);
nor U43421 (N_43421,N_42239,N_42175);
nor U43422 (N_43422,N_42867,N_42383);
and U43423 (N_43423,N_42637,N_42299);
or U43424 (N_43424,N_42667,N_42974);
xor U43425 (N_43425,N_42186,N_42064);
nand U43426 (N_43426,N_42415,N_42523);
nand U43427 (N_43427,N_42288,N_42177);
and U43428 (N_43428,N_42791,N_42077);
and U43429 (N_43429,N_42839,N_42999);
nand U43430 (N_43430,N_42590,N_42594);
or U43431 (N_43431,N_42524,N_42086);
nand U43432 (N_43432,N_42127,N_42824);
and U43433 (N_43433,N_42402,N_42102);
and U43434 (N_43434,N_42652,N_42085);
xor U43435 (N_43435,N_42119,N_42698);
or U43436 (N_43436,N_42015,N_42815);
nor U43437 (N_43437,N_42258,N_42541);
xor U43438 (N_43438,N_42058,N_42776);
nand U43439 (N_43439,N_42031,N_42518);
or U43440 (N_43440,N_42688,N_42456);
and U43441 (N_43441,N_42993,N_42806);
nor U43442 (N_43442,N_42567,N_42404);
and U43443 (N_43443,N_42724,N_42316);
nor U43444 (N_43444,N_42707,N_42451);
nor U43445 (N_43445,N_42731,N_42601);
or U43446 (N_43446,N_42392,N_42575);
and U43447 (N_43447,N_42908,N_42021);
and U43448 (N_43448,N_42300,N_42910);
or U43449 (N_43449,N_42290,N_42828);
xnor U43450 (N_43450,N_42259,N_42420);
nand U43451 (N_43451,N_42323,N_42790);
or U43452 (N_43452,N_42643,N_42754);
nor U43453 (N_43453,N_42994,N_42182);
xnor U43454 (N_43454,N_42333,N_42019);
and U43455 (N_43455,N_42849,N_42229);
xnor U43456 (N_43456,N_42028,N_42936);
nor U43457 (N_43457,N_42209,N_42274);
or U43458 (N_43458,N_42414,N_42821);
nand U43459 (N_43459,N_42482,N_42986);
or U43460 (N_43460,N_42138,N_42726);
nand U43461 (N_43461,N_42941,N_42344);
xor U43462 (N_43462,N_42639,N_42699);
and U43463 (N_43463,N_42356,N_42050);
nand U43464 (N_43464,N_42156,N_42798);
or U43465 (N_43465,N_42151,N_42930);
and U43466 (N_43466,N_42237,N_42913);
nor U43467 (N_43467,N_42586,N_42556);
or U43468 (N_43468,N_42840,N_42837);
nand U43469 (N_43469,N_42009,N_42653);
or U43470 (N_43470,N_42060,N_42807);
xor U43471 (N_43471,N_42444,N_42377);
or U43472 (N_43472,N_42885,N_42469);
xnor U43473 (N_43473,N_42141,N_42834);
and U43474 (N_43474,N_42369,N_42419);
nor U43475 (N_43475,N_42131,N_42440);
and U43476 (N_43476,N_42558,N_42407);
nor U43477 (N_43477,N_42358,N_42359);
nor U43478 (N_43478,N_42539,N_42150);
nand U43479 (N_43479,N_42388,N_42872);
or U43480 (N_43480,N_42570,N_42336);
nand U43481 (N_43481,N_42065,N_42149);
or U43482 (N_43482,N_42696,N_42213);
xor U43483 (N_43483,N_42738,N_42199);
nand U43484 (N_43484,N_42508,N_42510);
or U43485 (N_43485,N_42900,N_42746);
nand U43486 (N_43486,N_42272,N_42714);
or U43487 (N_43487,N_42007,N_42784);
xor U43488 (N_43488,N_42321,N_42976);
nor U43489 (N_43489,N_42371,N_42931);
xor U43490 (N_43490,N_42240,N_42121);
nor U43491 (N_43491,N_42851,N_42841);
xnor U43492 (N_43492,N_42484,N_42633);
nand U43493 (N_43493,N_42609,N_42497);
and U43494 (N_43494,N_42200,N_42987);
xnor U43495 (N_43495,N_42384,N_42365);
and U43496 (N_43496,N_42020,N_42270);
or U43497 (N_43497,N_42630,N_42155);
nand U43498 (N_43498,N_42756,N_42464);
nand U43499 (N_43499,N_42697,N_42621);
and U43500 (N_43500,N_42395,N_42425);
and U43501 (N_43501,N_42558,N_42517);
nand U43502 (N_43502,N_42029,N_42440);
nand U43503 (N_43503,N_42620,N_42033);
nand U43504 (N_43504,N_42505,N_42639);
or U43505 (N_43505,N_42972,N_42948);
nand U43506 (N_43506,N_42761,N_42635);
nand U43507 (N_43507,N_42601,N_42775);
nand U43508 (N_43508,N_42665,N_42117);
or U43509 (N_43509,N_42996,N_42375);
nor U43510 (N_43510,N_42490,N_42312);
and U43511 (N_43511,N_42762,N_42107);
xnor U43512 (N_43512,N_42644,N_42237);
and U43513 (N_43513,N_42954,N_42349);
xor U43514 (N_43514,N_42578,N_42438);
and U43515 (N_43515,N_42986,N_42381);
xnor U43516 (N_43516,N_42101,N_42714);
nor U43517 (N_43517,N_42753,N_42818);
and U43518 (N_43518,N_42703,N_42153);
nor U43519 (N_43519,N_42302,N_42592);
xor U43520 (N_43520,N_42142,N_42498);
nand U43521 (N_43521,N_42008,N_42307);
nor U43522 (N_43522,N_42297,N_42689);
nand U43523 (N_43523,N_42458,N_42357);
and U43524 (N_43524,N_42076,N_42277);
and U43525 (N_43525,N_42247,N_42033);
and U43526 (N_43526,N_42086,N_42327);
nand U43527 (N_43527,N_42252,N_42768);
nor U43528 (N_43528,N_42132,N_42801);
xor U43529 (N_43529,N_42088,N_42636);
or U43530 (N_43530,N_42084,N_42318);
xor U43531 (N_43531,N_42942,N_42989);
or U43532 (N_43532,N_42565,N_42641);
or U43533 (N_43533,N_42670,N_42144);
nor U43534 (N_43534,N_42137,N_42422);
and U43535 (N_43535,N_42132,N_42027);
nor U43536 (N_43536,N_42896,N_42999);
and U43537 (N_43537,N_42782,N_42026);
nand U43538 (N_43538,N_42880,N_42800);
xor U43539 (N_43539,N_42889,N_42356);
xnor U43540 (N_43540,N_42340,N_42174);
nand U43541 (N_43541,N_42404,N_42135);
xor U43542 (N_43542,N_42868,N_42994);
and U43543 (N_43543,N_42873,N_42845);
nand U43544 (N_43544,N_42833,N_42224);
and U43545 (N_43545,N_42670,N_42477);
or U43546 (N_43546,N_42354,N_42096);
nand U43547 (N_43547,N_42988,N_42553);
or U43548 (N_43548,N_42411,N_42349);
nor U43549 (N_43549,N_42560,N_42136);
and U43550 (N_43550,N_42641,N_42872);
nand U43551 (N_43551,N_42364,N_42036);
xor U43552 (N_43552,N_42373,N_42667);
or U43553 (N_43553,N_42868,N_42328);
nor U43554 (N_43554,N_42634,N_42415);
or U43555 (N_43555,N_42355,N_42328);
nor U43556 (N_43556,N_42745,N_42630);
xor U43557 (N_43557,N_42222,N_42750);
xnor U43558 (N_43558,N_42200,N_42398);
nand U43559 (N_43559,N_42578,N_42125);
or U43560 (N_43560,N_42304,N_42617);
and U43561 (N_43561,N_42705,N_42890);
nand U43562 (N_43562,N_42638,N_42291);
nand U43563 (N_43563,N_42475,N_42895);
nand U43564 (N_43564,N_42609,N_42089);
nor U43565 (N_43565,N_42604,N_42443);
xnor U43566 (N_43566,N_42111,N_42996);
nand U43567 (N_43567,N_42269,N_42994);
xor U43568 (N_43568,N_42066,N_42846);
xor U43569 (N_43569,N_42321,N_42659);
xor U43570 (N_43570,N_42827,N_42315);
or U43571 (N_43571,N_42726,N_42948);
or U43572 (N_43572,N_42891,N_42544);
nand U43573 (N_43573,N_42010,N_42318);
nand U43574 (N_43574,N_42471,N_42735);
nor U43575 (N_43575,N_42825,N_42808);
or U43576 (N_43576,N_42198,N_42320);
nand U43577 (N_43577,N_42866,N_42084);
or U43578 (N_43578,N_42104,N_42531);
xnor U43579 (N_43579,N_42516,N_42721);
and U43580 (N_43580,N_42212,N_42245);
and U43581 (N_43581,N_42366,N_42784);
and U43582 (N_43582,N_42324,N_42517);
or U43583 (N_43583,N_42481,N_42340);
or U43584 (N_43584,N_42240,N_42632);
nor U43585 (N_43585,N_42895,N_42694);
or U43586 (N_43586,N_42449,N_42015);
nor U43587 (N_43587,N_42530,N_42462);
xor U43588 (N_43588,N_42413,N_42612);
nand U43589 (N_43589,N_42213,N_42132);
nand U43590 (N_43590,N_42750,N_42846);
and U43591 (N_43591,N_42142,N_42600);
and U43592 (N_43592,N_42762,N_42598);
nor U43593 (N_43593,N_42171,N_42215);
and U43594 (N_43594,N_42743,N_42054);
and U43595 (N_43595,N_42903,N_42448);
xor U43596 (N_43596,N_42825,N_42369);
xor U43597 (N_43597,N_42167,N_42953);
and U43598 (N_43598,N_42249,N_42711);
xnor U43599 (N_43599,N_42852,N_42890);
xor U43600 (N_43600,N_42886,N_42129);
or U43601 (N_43601,N_42368,N_42578);
and U43602 (N_43602,N_42847,N_42038);
nor U43603 (N_43603,N_42179,N_42205);
and U43604 (N_43604,N_42222,N_42849);
nor U43605 (N_43605,N_42412,N_42291);
and U43606 (N_43606,N_42631,N_42293);
or U43607 (N_43607,N_42635,N_42352);
nor U43608 (N_43608,N_42526,N_42584);
and U43609 (N_43609,N_42864,N_42631);
xnor U43610 (N_43610,N_42862,N_42858);
nor U43611 (N_43611,N_42598,N_42979);
or U43612 (N_43612,N_42514,N_42596);
xnor U43613 (N_43613,N_42537,N_42045);
or U43614 (N_43614,N_42198,N_42156);
or U43615 (N_43615,N_42958,N_42677);
xor U43616 (N_43616,N_42523,N_42076);
nand U43617 (N_43617,N_42435,N_42047);
nor U43618 (N_43618,N_42736,N_42901);
nand U43619 (N_43619,N_42504,N_42399);
or U43620 (N_43620,N_42584,N_42478);
nor U43621 (N_43621,N_42237,N_42931);
nor U43622 (N_43622,N_42533,N_42913);
nor U43623 (N_43623,N_42519,N_42427);
and U43624 (N_43624,N_42010,N_42228);
or U43625 (N_43625,N_42109,N_42999);
nand U43626 (N_43626,N_42428,N_42425);
nor U43627 (N_43627,N_42997,N_42132);
nand U43628 (N_43628,N_42309,N_42418);
nor U43629 (N_43629,N_42902,N_42491);
nand U43630 (N_43630,N_42069,N_42472);
and U43631 (N_43631,N_42148,N_42707);
or U43632 (N_43632,N_42998,N_42744);
nand U43633 (N_43633,N_42644,N_42519);
nor U43634 (N_43634,N_42332,N_42498);
or U43635 (N_43635,N_42780,N_42138);
or U43636 (N_43636,N_42468,N_42633);
xnor U43637 (N_43637,N_42320,N_42720);
and U43638 (N_43638,N_42531,N_42565);
and U43639 (N_43639,N_42674,N_42719);
or U43640 (N_43640,N_42035,N_42962);
nor U43641 (N_43641,N_42565,N_42126);
or U43642 (N_43642,N_42550,N_42955);
nor U43643 (N_43643,N_42393,N_42235);
nand U43644 (N_43644,N_42883,N_42237);
xnor U43645 (N_43645,N_42174,N_42787);
nand U43646 (N_43646,N_42851,N_42875);
nor U43647 (N_43647,N_42257,N_42833);
and U43648 (N_43648,N_42425,N_42650);
nand U43649 (N_43649,N_42373,N_42181);
nor U43650 (N_43650,N_42494,N_42536);
or U43651 (N_43651,N_42013,N_42733);
xnor U43652 (N_43652,N_42258,N_42441);
and U43653 (N_43653,N_42063,N_42921);
nand U43654 (N_43654,N_42539,N_42394);
or U43655 (N_43655,N_42969,N_42241);
nor U43656 (N_43656,N_42626,N_42598);
and U43657 (N_43657,N_42757,N_42317);
nand U43658 (N_43658,N_42529,N_42374);
and U43659 (N_43659,N_42743,N_42517);
and U43660 (N_43660,N_42501,N_42582);
and U43661 (N_43661,N_42365,N_42284);
and U43662 (N_43662,N_42920,N_42067);
nor U43663 (N_43663,N_42631,N_42132);
nor U43664 (N_43664,N_42232,N_42021);
and U43665 (N_43665,N_42720,N_42226);
or U43666 (N_43666,N_42194,N_42521);
or U43667 (N_43667,N_42980,N_42655);
xor U43668 (N_43668,N_42354,N_42101);
nor U43669 (N_43669,N_42835,N_42184);
and U43670 (N_43670,N_42077,N_42789);
and U43671 (N_43671,N_42857,N_42092);
xnor U43672 (N_43672,N_42197,N_42944);
nor U43673 (N_43673,N_42129,N_42637);
nor U43674 (N_43674,N_42647,N_42495);
and U43675 (N_43675,N_42160,N_42888);
nor U43676 (N_43676,N_42995,N_42865);
nand U43677 (N_43677,N_42261,N_42586);
nor U43678 (N_43678,N_42928,N_42450);
nor U43679 (N_43679,N_42291,N_42741);
xor U43680 (N_43680,N_42521,N_42216);
xnor U43681 (N_43681,N_42719,N_42439);
nand U43682 (N_43682,N_42860,N_42635);
nor U43683 (N_43683,N_42998,N_42071);
and U43684 (N_43684,N_42766,N_42478);
nor U43685 (N_43685,N_42316,N_42052);
or U43686 (N_43686,N_42248,N_42753);
or U43687 (N_43687,N_42091,N_42999);
xnor U43688 (N_43688,N_42248,N_42499);
nor U43689 (N_43689,N_42631,N_42159);
nor U43690 (N_43690,N_42427,N_42587);
xor U43691 (N_43691,N_42762,N_42716);
nor U43692 (N_43692,N_42693,N_42931);
nor U43693 (N_43693,N_42329,N_42322);
and U43694 (N_43694,N_42730,N_42718);
and U43695 (N_43695,N_42216,N_42766);
and U43696 (N_43696,N_42781,N_42936);
nand U43697 (N_43697,N_42676,N_42387);
or U43698 (N_43698,N_42201,N_42840);
or U43699 (N_43699,N_42770,N_42418);
or U43700 (N_43700,N_42214,N_42137);
nor U43701 (N_43701,N_42706,N_42161);
nor U43702 (N_43702,N_42107,N_42612);
xnor U43703 (N_43703,N_42008,N_42271);
nor U43704 (N_43704,N_42376,N_42621);
nand U43705 (N_43705,N_42244,N_42622);
xnor U43706 (N_43706,N_42360,N_42233);
and U43707 (N_43707,N_42097,N_42697);
xor U43708 (N_43708,N_42520,N_42790);
nor U43709 (N_43709,N_42301,N_42866);
nand U43710 (N_43710,N_42216,N_42326);
or U43711 (N_43711,N_42127,N_42884);
and U43712 (N_43712,N_42771,N_42250);
and U43713 (N_43713,N_42747,N_42151);
nand U43714 (N_43714,N_42269,N_42673);
nor U43715 (N_43715,N_42421,N_42933);
and U43716 (N_43716,N_42250,N_42320);
or U43717 (N_43717,N_42440,N_42322);
xnor U43718 (N_43718,N_42077,N_42827);
and U43719 (N_43719,N_42747,N_42780);
xor U43720 (N_43720,N_42935,N_42241);
or U43721 (N_43721,N_42467,N_42733);
nor U43722 (N_43722,N_42912,N_42639);
and U43723 (N_43723,N_42115,N_42864);
or U43724 (N_43724,N_42838,N_42197);
or U43725 (N_43725,N_42806,N_42866);
xnor U43726 (N_43726,N_42445,N_42094);
nor U43727 (N_43727,N_42084,N_42949);
and U43728 (N_43728,N_42678,N_42470);
and U43729 (N_43729,N_42931,N_42712);
xor U43730 (N_43730,N_42109,N_42758);
nor U43731 (N_43731,N_42578,N_42552);
nor U43732 (N_43732,N_42167,N_42521);
and U43733 (N_43733,N_42325,N_42311);
and U43734 (N_43734,N_42621,N_42331);
nor U43735 (N_43735,N_42588,N_42581);
or U43736 (N_43736,N_42995,N_42889);
or U43737 (N_43737,N_42965,N_42604);
xnor U43738 (N_43738,N_42241,N_42523);
nor U43739 (N_43739,N_42227,N_42107);
or U43740 (N_43740,N_42362,N_42244);
nor U43741 (N_43741,N_42576,N_42520);
or U43742 (N_43742,N_42109,N_42625);
nor U43743 (N_43743,N_42139,N_42505);
nor U43744 (N_43744,N_42345,N_42750);
nor U43745 (N_43745,N_42483,N_42433);
nand U43746 (N_43746,N_42376,N_42260);
nand U43747 (N_43747,N_42116,N_42103);
nor U43748 (N_43748,N_42196,N_42358);
or U43749 (N_43749,N_42619,N_42617);
nand U43750 (N_43750,N_42379,N_42165);
or U43751 (N_43751,N_42777,N_42682);
or U43752 (N_43752,N_42623,N_42499);
xnor U43753 (N_43753,N_42274,N_42943);
and U43754 (N_43754,N_42178,N_42552);
and U43755 (N_43755,N_42469,N_42723);
or U43756 (N_43756,N_42650,N_42368);
xor U43757 (N_43757,N_42130,N_42094);
xnor U43758 (N_43758,N_42207,N_42211);
or U43759 (N_43759,N_42426,N_42327);
nand U43760 (N_43760,N_42683,N_42851);
nand U43761 (N_43761,N_42330,N_42497);
or U43762 (N_43762,N_42204,N_42556);
xnor U43763 (N_43763,N_42542,N_42982);
or U43764 (N_43764,N_42538,N_42579);
or U43765 (N_43765,N_42808,N_42950);
or U43766 (N_43766,N_42779,N_42466);
nor U43767 (N_43767,N_42656,N_42429);
or U43768 (N_43768,N_42669,N_42364);
nor U43769 (N_43769,N_42330,N_42232);
or U43770 (N_43770,N_42328,N_42114);
nand U43771 (N_43771,N_42888,N_42238);
nor U43772 (N_43772,N_42459,N_42670);
or U43773 (N_43773,N_42427,N_42061);
nand U43774 (N_43774,N_42965,N_42697);
nand U43775 (N_43775,N_42224,N_42805);
or U43776 (N_43776,N_42079,N_42215);
and U43777 (N_43777,N_42714,N_42153);
and U43778 (N_43778,N_42231,N_42546);
and U43779 (N_43779,N_42705,N_42160);
or U43780 (N_43780,N_42117,N_42056);
and U43781 (N_43781,N_42823,N_42831);
xor U43782 (N_43782,N_42651,N_42149);
or U43783 (N_43783,N_42678,N_42205);
or U43784 (N_43784,N_42984,N_42261);
nand U43785 (N_43785,N_42255,N_42757);
nand U43786 (N_43786,N_42582,N_42744);
nand U43787 (N_43787,N_42523,N_42993);
nand U43788 (N_43788,N_42024,N_42552);
and U43789 (N_43789,N_42009,N_42057);
or U43790 (N_43790,N_42750,N_42586);
nor U43791 (N_43791,N_42649,N_42143);
nand U43792 (N_43792,N_42940,N_42666);
nor U43793 (N_43793,N_42903,N_42981);
nand U43794 (N_43794,N_42520,N_42267);
nor U43795 (N_43795,N_42626,N_42202);
or U43796 (N_43796,N_42333,N_42891);
and U43797 (N_43797,N_42596,N_42008);
or U43798 (N_43798,N_42778,N_42429);
and U43799 (N_43799,N_42596,N_42905);
or U43800 (N_43800,N_42629,N_42216);
or U43801 (N_43801,N_42706,N_42092);
or U43802 (N_43802,N_42050,N_42468);
nor U43803 (N_43803,N_42096,N_42109);
and U43804 (N_43804,N_42890,N_42421);
and U43805 (N_43805,N_42048,N_42338);
xor U43806 (N_43806,N_42624,N_42035);
and U43807 (N_43807,N_42085,N_42764);
nand U43808 (N_43808,N_42965,N_42474);
nor U43809 (N_43809,N_42293,N_42268);
or U43810 (N_43810,N_42323,N_42653);
xnor U43811 (N_43811,N_42441,N_42676);
and U43812 (N_43812,N_42042,N_42315);
or U43813 (N_43813,N_42884,N_42650);
xor U43814 (N_43814,N_42521,N_42483);
xnor U43815 (N_43815,N_42140,N_42230);
nor U43816 (N_43816,N_42070,N_42499);
and U43817 (N_43817,N_42641,N_42260);
xor U43818 (N_43818,N_42373,N_42215);
nand U43819 (N_43819,N_42530,N_42546);
nor U43820 (N_43820,N_42428,N_42015);
nand U43821 (N_43821,N_42749,N_42773);
nand U43822 (N_43822,N_42378,N_42326);
or U43823 (N_43823,N_42221,N_42133);
nor U43824 (N_43824,N_42772,N_42349);
xnor U43825 (N_43825,N_42611,N_42098);
nor U43826 (N_43826,N_42661,N_42373);
and U43827 (N_43827,N_42525,N_42563);
and U43828 (N_43828,N_42512,N_42995);
nor U43829 (N_43829,N_42082,N_42996);
nand U43830 (N_43830,N_42617,N_42116);
and U43831 (N_43831,N_42875,N_42725);
nand U43832 (N_43832,N_42426,N_42995);
and U43833 (N_43833,N_42275,N_42453);
nor U43834 (N_43834,N_42771,N_42995);
or U43835 (N_43835,N_42447,N_42913);
and U43836 (N_43836,N_42117,N_42184);
nor U43837 (N_43837,N_42475,N_42703);
nand U43838 (N_43838,N_42501,N_42067);
or U43839 (N_43839,N_42306,N_42867);
and U43840 (N_43840,N_42279,N_42324);
and U43841 (N_43841,N_42237,N_42219);
and U43842 (N_43842,N_42952,N_42417);
or U43843 (N_43843,N_42492,N_42308);
xnor U43844 (N_43844,N_42811,N_42969);
xnor U43845 (N_43845,N_42093,N_42568);
nor U43846 (N_43846,N_42604,N_42364);
nand U43847 (N_43847,N_42737,N_42490);
xor U43848 (N_43848,N_42320,N_42451);
xor U43849 (N_43849,N_42769,N_42098);
nand U43850 (N_43850,N_42167,N_42243);
and U43851 (N_43851,N_42066,N_42239);
and U43852 (N_43852,N_42840,N_42430);
or U43853 (N_43853,N_42816,N_42950);
or U43854 (N_43854,N_42107,N_42186);
nor U43855 (N_43855,N_42105,N_42349);
xor U43856 (N_43856,N_42572,N_42005);
or U43857 (N_43857,N_42182,N_42550);
nand U43858 (N_43858,N_42461,N_42717);
nand U43859 (N_43859,N_42306,N_42779);
nor U43860 (N_43860,N_42986,N_42899);
or U43861 (N_43861,N_42047,N_42725);
or U43862 (N_43862,N_42321,N_42650);
xor U43863 (N_43863,N_42502,N_42733);
xnor U43864 (N_43864,N_42864,N_42072);
or U43865 (N_43865,N_42566,N_42232);
nand U43866 (N_43866,N_42347,N_42683);
nor U43867 (N_43867,N_42514,N_42343);
nor U43868 (N_43868,N_42528,N_42503);
nor U43869 (N_43869,N_42550,N_42508);
or U43870 (N_43870,N_42284,N_42476);
or U43871 (N_43871,N_42556,N_42060);
or U43872 (N_43872,N_42770,N_42025);
xor U43873 (N_43873,N_42107,N_42649);
xor U43874 (N_43874,N_42879,N_42955);
nor U43875 (N_43875,N_42982,N_42620);
or U43876 (N_43876,N_42324,N_42139);
and U43877 (N_43877,N_42609,N_42776);
or U43878 (N_43878,N_42449,N_42217);
or U43879 (N_43879,N_42763,N_42563);
nor U43880 (N_43880,N_42159,N_42734);
xnor U43881 (N_43881,N_42946,N_42215);
nand U43882 (N_43882,N_42414,N_42707);
nand U43883 (N_43883,N_42766,N_42122);
nand U43884 (N_43884,N_42894,N_42953);
nand U43885 (N_43885,N_42517,N_42672);
nor U43886 (N_43886,N_42210,N_42936);
xnor U43887 (N_43887,N_42500,N_42891);
xor U43888 (N_43888,N_42442,N_42044);
nand U43889 (N_43889,N_42608,N_42275);
or U43890 (N_43890,N_42340,N_42170);
nand U43891 (N_43891,N_42404,N_42821);
xor U43892 (N_43892,N_42917,N_42049);
and U43893 (N_43893,N_42284,N_42184);
nand U43894 (N_43894,N_42445,N_42989);
and U43895 (N_43895,N_42340,N_42772);
or U43896 (N_43896,N_42062,N_42559);
nand U43897 (N_43897,N_42058,N_42370);
xnor U43898 (N_43898,N_42905,N_42010);
and U43899 (N_43899,N_42643,N_42475);
nand U43900 (N_43900,N_42721,N_42990);
nor U43901 (N_43901,N_42808,N_42958);
xor U43902 (N_43902,N_42270,N_42904);
nand U43903 (N_43903,N_42807,N_42927);
or U43904 (N_43904,N_42174,N_42268);
nand U43905 (N_43905,N_42931,N_42202);
xnor U43906 (N_43906,N_42265,N_42551);
or U43907 (N_43907,N_42454,N_42864);
nand U43908 (N_43908,N_42118,N_42557);
or U43909 (N_43909,N_42667,N_42676);
nor U43910 (N_43910,N_42772,N_42846);
xnor U43911 (N_43911,N_42970,N_42179);
or U43912 (N_43912,N_42161,N_42877);
nor U43913 (N_43913,N_42117,N_42344);
and U43914 (N_43914,N_42804,N_42356);
nand U43915 (N_43915,N_42836,N_42594);
or U43916 (N_43916,N_42835,N_42091);
and U43917 (N_43917,N_42770,N_42081);
nand U43918 (N_43918,N_42640,N_42292);
and U43919 (N_43919,N_42558,N_42707);
nor U43920 (N_43920,N_42589,N_42484);
or U43921 (N_43921,N_42383,N_42955);
nor U43922 (N_43922,N_42737,N_42966);
xor U43923 (N_43923,N_42998,N_42159);
xnor U43924 (N_43924,N_42004,N_42420);
nor U43925 (N_43925,N_42904,N_42041);
and U43926 (N_43926,N_42204,N_42607);
or U43927 (N_43927,N_42565,N_42917);
and U43928 (N_43928,N_42985,N_42954);
or U43929 (N_43929,N_42796,N_42773);
or U43930 (N_43930,N_42892,N_42511);
xor U43931 (N_43931,N_42046,N_42529);
nor U43932 (N_43932,N_42479,N_42009);
xnor U43933 (N_43933,N_42099,N_42697);
xor U43934 (N_43934,N_42211,N_42567);
nor U43935 (N_43935,N_42806,N_42104);
xnor U43936 (N_43936,N_42605,N_42566);
xnor U43937 (N_43937,N_42512,N_42481);
nor U43938 (N_43938,N_42638,N_42919);
nor U43939 (N_43939,N_42765,N_42367);
or U43940 (N_43940,N_42171,N_42182);
nand U43941 (N_43941,N_42994,N_42679);
nor U43942 (N_43942,N_42158,N_42339);
and U43943 (N_43943,N_42432,N_42593);
and U43944 (N_43944,N_42914,N_42891);
nor U43945 (N_43945,N_42279,N_42207);
nor U43946 (N_43946,N_42594,N_42972);
nand U43947 (N_43947,N_42610,N_42429);
xnor U43948 (N_43948,N_42809,N_42136);
xor U43949 (N_43949,N_42712,N_42606);
or U43950 (N_43950,N_42372,N_42523);
nor U43951 (N_43951,N_42535,N_42234);
nor U43952 (N_43952,N_42063,N_42054);
nor U43953 (N_43953,N_42604,N_42351);
nand U43954 (N_43954,N_42728,N_42675);
nand U43955 (N_43955,N_42707,N_42789);
or U43956 (N_43956,N_42176,N_42385);
and U43957 (N_43957,N_42771,N_42937);
nor U43958 (N_43958,N_42832,N_42715);
xor U43959 (N_43959,N_42429,N_42255);
xnor U43960 (N_43960,N_42277,N_42225);
nand U43961 (N_43961,N_42697,N_42344);
and U43962 (N_43962,N_42932,N_42425);
nand U43963 (N_43963,N_42388,N_42140);
or U43964 (N_43964,N_42603,N_42242);
nor U43965 (N_43965,N_42307,N_42874);
xnor U43966 (N_43966,N_42533,N_42312);
nand U43967 (N_43967,N_42555,N_42426);
nand U43968 (N_43968,N_42319,N_42121);
or U43969 (N_43969,N_42438,N_42115);
or U43970 (N_43970,N_42344,N_42217);
or U43971 (N_43971,N_42695,N_42318);
or U43972 (N_43972,N_42974,N_42102);
or U43973 (N_43973,N_42142,N_42090);
nor U43974 (N_43974,N_42914,N_42829);
or U43975 (N_43975,N_42056,N_42087);
or U43976 (N_43976,N_42408,N_42431);
or U43977 (N_43977,N_42095,N_42268);
xnor U43978 (N_43978,N_42884,N_42548);
or U43979 (N_43979,N_42136,N_42411);
and U43980 (N_43980,N_42168,N_42672);
and U43981 (N_43981,N_42973,N_42673);
or U43982 (N_43982,N_42569,N_42039);
nor U43983 (N_43983,N_42812,N_42617);
and U43984 (N_43984,N_42698,N_42678);
or U43985 (N_43985,N_42037,N_42365);
or U43986 (N_43986,N_42584,N_42097);
nor U43987 (N_43987,N_42165,N_42864);
nand U43988 (N_43988,N_42560,N_42201);
or U43989 (N_43989,N_42808,N_42763);
nor U43990 (N_43990,N_42961,N_42138);
and U43991 (N_43991,N_42986,N_42062);
or U43992 (N_43992,N_42469,N_42543);
xnor U43993 (N_43993,N_42079,N_42807);
and U43994 (N_43994,N_42871,N_42020);
and U43995 (N_43995,N_42998,N_42386);
nor U43996 (N_43996,N_42155,N_42108);
and U43997 (N_43997,N_42428,N_42301);
xor U43998 (N_43998,N_42190,N_42420);
or U43999 (N_43999,N_42795,N_42290);
and U44000 (N_44000,N_43784,N_43175);
or U44001 (N_44001,N_43874,N_43883);
nand U44002 (N_44002,N_43765,N_43952);
xnor U44003 (N_44003,N_43377,N_43168);
nor U44004 (N_44004,N_43145,N_43225);
nor U44005 (N_44005,N_43212,N_43663);
xnor U44006 (N_44006,N_43977,N_43871);
nand U44007 (N_44007,N_43019,N_43155);
and U44008 (N_44008,N_43656,N_43343);
nand U44009 (N_44009,N_43443,N_43901);
xnor U44010 (N_44010,N_43555,N_43709);
xnor U44011 (N_44011,N_43713,N_43915);
and U44012 (N_44012,N_43889,N_43353);
and U44013 (N_44013,N_43109,N_43851);
and U44014 (N_44014,N_43916,N_43919);
xnor U44015 (N_44015,N_43446,N_43480);
and U44016 (N_44016,N_43575,N_43869);
and U44017 (N_44017,N_43960,N_43131);
and U44018 (N_44018,N_43689,N_43124);
nor U44019 (N_44019,N_43270,N_43737);
nor U44020 (N_44020,N_43537,N_43974);
or U44021 (N_44021,N_43422,N_43299);
or U44022 (N_44022,N_43303,N_43870);
nand U44023 (N_44023,N_43267,N_43676);
nor U44024 (N_44024,N_43039,N_43272);
xor U44025 (N_44025,N_43886,N_43126);
xnor U44026 (N_44026,N_43804,N_43077);
and U44027 (N_44027,N_43875,N_43240);
or U44028 (N_44028,N_43018,N_43056);
or U44029 (N_44029,N_43242,N_43605);
nor U44030 (N_44030,N_43021,N_43690);
nand U44031 (N_44031,N_43582,N_43652);
xnor U44032 (N_44032,N_43583,N_43858);
xnor U44033 (N_44033,N_43328,N_43466);
xor U44034 (N_44034,N_43815,N_43708);
and U44035 (N_44035,N_43771,N_43301);
and U44036 (N_44036,N_43230,N_43619);
and U44037 (N_44037,N_43630,N_43520);
xnor U44038 (N_44038,N_43667,N_43703);
nand U44039 (N_44039,N_43584,N_43662);
xor U44040 (N_44040,N_43360,N_43534);
and U44041 (N_44041,N_43167,N_43203);
or U44042 (N_44042,N_43472,N_43772);
nand U44043 (N_44043,N_43705,N_43518);
nor U44044 (N_44044,N_43551,N_43087);
and U44045 (N_44045,N_43751,N_43361);
or U44046 (N_44046,N_43146,N_43941);
and U44047 (N_44047,N_43214,N_43532);
nand U44048 (N_44048,N_43906,N_43052);
or U44049 (N_44049,N_43005,N_43330);
and U44050 (N_44050,N_43528,N_43151);
nand U44051 (N_44051,N_43339,N_43793);
or U44052 (N_44052,N_43856,N_43269);
nor U44053 (N_44053,N_43276,N_43921);
nand U44054 (N_44054,N_43476,N_43779);
or U44055 (N_44055,N_43591,N_43295);
and U44056 (N_44056,N_43562,N_43973);
xor U44057 (N_44057,N_43491,N_43133);
nor U44058 (N_44058,N_43334,N_43780);
nand U44059 (N_44059,N_43154,N_43937);
nor U44060 (N_44060,N_43899,N_43435);
nor U44061 (N_44061,N_43069,N_43986);
xor U44062 (N_44062,N_43064,N_43351);
and U44063 (N_44063,N_43822,N_43816);
xnor U44064 (N_44064,N_43580,N_43226);
xnor U44065 (N_44065,N_43454,N_43402);
xor U44066 (N_44066,N_43910,N_43695);
or U44067 (N_44067,N_43818,N_43726);
nor U44068 (N_44068,N_43523,N_43278);
nor U44069 (N_44069,N_43691,N_43075);
nand U44070 (N_44070,N_43437,N_43012);
nor U44071 (N_44071,N_43011,N_43380);
nor U44072 (N_44072,N_43794,N_43680);
nand U44073 (N_44073,N_43204,N_43354);
xnor U44074 (N_44074,N_43633,N_43451);
nand U44075 (N_44075,N_43231,N_43594);
and U44076 (N_44076,N_43588,N_43376);
and U44077 (N_44077,N_43678,N_43529);
xor U44078 (N_44078,N_43622,N_43478);
nor U44079 (N_44079,N_43470,N_43929);
nand U44080 (N_44080,N_43090,N_43103);
nand U44081 (N_44081,N_43248,N_43623);
and U44082 (N_44082,N_43408,N_43542);
and U44083 (N_44083,N_43441,N_43258);
nor U44084 (N_44084,N_43785,N_43911);
or U44085 (N_44085,N_43234,N_43833);
nor U44086 (N_44086,N_43597,N_43552);
and U44087 (N_44087,N_43569,N_43010);
nand U44088 (N_44088,N_43586,N_43671);
and U44089 (N_44089,N_43461,N_43022);
xor U44090 (N_44090,N_43504,N_43876);
nor U44091 (N_44091,N_43958,N_43367);
or U44092 (N_44092,N_43798,N_43349);
nor U44093 (N_44093,N_43199,N_43745);
or U44094 (N_44094,N_43388,N_43163);
xnor U44095 (N_44095,N_43836,N_43089);
and U44096 (N_44096,N_43266,N_43420);
or U44097 (N_44097,N_43953,N_43967);
nand U44098 (N_44098,N_43501,N_43307);
xor U44099 (N_44099,N_43099,N_43912);
xor U44100 (N_44100,N_43280,N_43762);
xnor U44101 (N_44101,N_43608,N_43355);
or U44102 (N_44102,N_43326,N_43810);
nand U44103 (N_44103,N_43140,N_43189);
and U44104 (N_44104,N_43999,N_43174);
xor U44105 (N_44105,N_43202,N_43603);
or U44106 (N_44106,N_43766,N_43421);
nand U44107 (N_44107,N_43365,N_43992);
nor U44108 (N_44108,N_43842,N_43527);
nand U44109 (N_44109,N_43313,N_43809);
xor U44110 (N_44110,N_43302,N_43926);
xnor U44111 (N_44111,N_43814,N_43268);
nor U44112 (N_44112,N_43627,N_43497);
nor U44113 (N_44113,N_43065,N_43935);
xnor U44114 (N_44114,N_43393,N_43561);
xnor U44115 (N_44115,N_43185,N_43639);
and U44116 (N_44116,N_43878,N_43255);
nor U44117 (N_44117,N_43898,N_43978);
and U44118 (N_44118,N_43522,N_43544);
or U44119 (N_44119,N_43796,N_43572);
or U44120 (N_44120,N_43318,N_43288);
nor U44121 (N_44121,N_43642,N_43070);
nor U44122 (N_44122,N_43853,N_43673);
or U44123 (N_44123,N_43382,N_43001);
and U44124 (N_44124,N_43492,N_43533);
xor U44125 (N_44125,N_43100,N_43754);
or U44126 (N_44126,N_43803,N_43505);
or U44127 (N_44127,N_43949,N_43985);
and U44128 (N_44128,N_43548,N_43828);
or U44129 (N_44129,N_43494,N_43710);
xnor U44130 (N_44130,N_43568,N_43612);
nor U44131 (N_44131,N_43291,N_43027);
or U44132 (N_44132,N_43183,N_43062);
nand U44133 (N_44133,N_43757,N_43991);
nand U44134 (N_44134,N_43681,N_43625);
nor U44135 (N_44135,N_43315,N_43909);
nor U44136 (N_44136,N_43609,N_43936);
or U44137 (N_44137,N_43257,N_43932);
nor U44138 (N_44138,N_43008,N_43723);
or U44139 (N_44139,N_43375,N_43473);
nor U44140 (N_44140,N_43106,N_43650);
and U44141 (N_44141,N_43186,N_43546);
nor U44142 (N_44142,N_43325,N_43054);
or U44143 (N_44143,N_43989,N_43442);
xor U44144 (N_44144,N_43023,N_43033);
xnor U44145 (N_44145,N_43788,N_43968);
xor U44146 (N_44146,N_43517,N_43811);
nor U44147 (N_44147,N_43802,N_43373);
or U44148 (N_44148,N_43409,N_43670);
and U44149 (N_44149,N_43756,N_43127);
or U44150 (N_44150,N_43073,N_43223);
nand U44151 (N_44151,N_43825,N_43787);
nand U44152 (N_44152,N_43347,N_43035);
nand U44153 (N_44153,N_43434,N_43948);
or U44154 (N_44154,N_43120,N_43419);
and U44155 (N_44155,N_43162,N_43563);
nor U44156 (N_44156,N_43698,N_43342);
nand U44157 (N_44157,N_43245,N_43463);
nand U44158 (N_44158,N_43465,N_43975);
nand U44159 (N_44159,N_43007,N_43640);
and U44160 (N_44160,N_43942,N_43835);
nand U44161 (N_44161,N_43507,N_43746);
nor U44162 (N_44162,N_43452,N_43674);
nor U44163 (N_44163,N_43567,N_43239);
nor U44164 (N_44164,N_43966,N_43381);
xnor U44165 (N_44165,N_43574,N_43558);
nor U44166 (N_44166,N_43317,N_43116);
nand U44167 (N_44167,N_43982,N_43888);
nor U44168 (N_44168,N_43571,N_43436);
nand U44169 (N_44169,N_43564,N_43078);
nor U44170 (N_44170,N_43237,N_43006);
nand U44171 (N_44171,N_43806,N_43407);
nor U44172 (N_44172,N_43016,N_43866);
nand U44173 (N_44173,N_43045,N_43512);
nand U44174 (N_44174,N_43515,N_43444);
nor U44175 (N_44175,N_43995,N_43128);
or U44176 (N_44176,N_43294,N_43720);
nor U44177 (N_44177,N_43727,N_43538);
nor U44178 (N_44178,N_43323,N_43955);
nor U44179 (N_44179,N_43651,N_43867);
or U44180 (N_44180,N_43410,N_43243);
or U44181 (N_44181,N_43536,N_43819);
nand U44182 (N_44182,N_43617,N_43577);
xor U44183 (N_44183,N_43578,N_43646);
nand U44184 (N_44184,N_43755,N_43110);
or U44185 (N_44185,N_43715,N_43770);
xor U44186 (N_44186,N_43438,N_43246);
or U44187 (N_44187,N_43404,N_43406);
or U44188 (N_44188,N_43644,N_43287);
nand U44189 (N_44189,N_43098,N_43777);
xnor U44190 (N_44190,N_43359,N_43554);
nor U44191 (N_44191,N_43807,N_43907);
or U44192 (N_44192,N_43138,N_43044);
and U44193 (N_44193,N_43002,N_43618);
xnor U44194 (N_44194,N_43930,N_43774);
nor U44195 (N_44195,N_43686,N_43259);
xor U44196 (N_44196,N_43232,N_43954);
or U44197 (N_44197,N_43289,N_43742);
and U44198 (N_44198,N_43813,N_43635);
nor U44199 (N_44199,N_43606,N_43193);
nor U44200 (N_44200,N_43150,N_43111);
nor U44201 (N_44201,N_43769,N_43573);
nor U44202 (N_44202,N_43412,N_43540);
nand U44203 (N_44203,N_43397,N_43498);
and U44204 (N_44204,N_43081,N_43217);
or U44205 (N_44205,N_43366,N_43880);
xnor U44206 (N_44206,N_43384,N_43735);
nand U44207 (N_44207,N_43961,N_43104);
nor U44208 (N_44208,N_43697,N_43047);
or U44209 (N_44209,N_43363,N_43352);
xor U44210 (N_44210,N_43068,N_43215);
or U44211 (N_44211,N_43261,N_43998);
nor U44212 (N_44212,N_43645,N_43132);
and U44213 (N_44213,N_43487,N_43071);
and U44214 (N_44214,N_43170,N_43320);
nand U44215 (N_44215,N_43972,N_43097);
xnor U44216 (N_44216,N_43621,N_43218);
nand U44217 (N_44217,N_43331,N_43864);
and U44218 (N_44218,N_43728,N_43643);
nand U44219 (N_44219,N_43519,N_43539);
xnor U44220 (N_44220,N_43130,N_43036);
nand U44221 (N_44221,N_43172,N_43666);
and U44222 (N_44222,N_43076,N_43620);
and U44223 (N_44223,N_43198,N_43611);
nor U44224 (N_44224,N_43395,N_43252);
nor U44225 (N_44225,N_43971,N_43928);
or U44226 (N_44226,N_43768,N_43565);
or U44227 (N_44227,N_43030,N_43700);
nor U44228 (N_44228,N_43485,N_43776);
nor U44229 (N_44229,N_43238,N_43702);
nor U44230 (N_44230,N_43416,N_43368);
xnor U44231 (N_44231,N_43500,N_43468);
nor U44232 (N_44232,N_43009,N_43590);
or U44233 (N_44233,N_43153,N_43043);
nand U44234 (N_44234,N_43877,N_43450);
nand U44235 (N_44235,N_43696,N_43309);
and U44236 (N_44236,N_43729,N_43525);
nor U44237 (N_44237,N_43830,N_43904);
or U44238 (N_44238,N_43418,N_43271);
nor U44239 (N_44239,N_43843,N_43587);
xor U44240 (N_44240,N_43891,N_43903);
or U44241 (N_44241,N_43469,N_43987);
or U44242 (N_44242,N_43939,N_43984);
or U44243 (N_44243,N_43134,N_43428);
xnor U44244 (N_44244,N_43905,N_43080);
nand U44245 (N_44245,N_43514,N_43764);
xor U44246 (N_44246,N_43283,N_43029);
xnor U44247 (N_44247,N_43661,N_43460);
nand U44248 (N_44248,N_43881,N_43837);
or U44249 (N_44249,N_43508,N_43171);
xnor U44250 (N_44250,N_43657,N_43279);
nand U44251 (N_44251,N_43306,N_43964);
and U44252 (N_44252,N_43464,N_43371);
or U44253 (N_44253,N_43254,N_43415);
nand U44254 (N_44254,N_43628,N_43601);
or U44255 (N_44255,N_43716,N_43216);
nand U44256 (N_44256,N_43838,N_43829);
or U44257 (N_44257,N_43297,N_43839);
nor U44258 (N_44258,N_43337,N_43499);
and U44259 (N_44259,N_43025,N_43761);
xor U44260 (N_44260,N_43176,N_43191);
and U44261 (N_44261,N_43117,N_43453);
nor U44262 (N_44262,N_43447,N_43626);
and U44263 (N_44263,N_43970,N_43826);
xor U44264 (N_44264,N_43892,N_43273);
nand U44265 (N_44265,N_43137,N_43227);
xnor U44266 (N_44266,N_43413,N_43850);
xnor U44267 (N_44267,N_43918,N_43253);
xnor U44268 (N_44268,N_43310,N_43139);
xnor U44269 (N_44269,N_43722,N_43086);
and U44270 (N_44270,N_43900,N_43741);
xnor U44271 (N_44271,N_43855,N_43861);
nand U44272 (N_44272,N_43182,N_43882);
xnor U44273 (N_44273,N_43341,N_43229);
nor U44274 (N_44274,N_43456,N_43530);
nand U44275 (N_44275,N_43792,N_43061);
nor U44276 (N_44276,N_43604,N_43108);
and U44277 (N_44277,N_43057,N_43541);
nand U44278 (N_44278,N_43902,N_43988);
xnor U44279 (N_44279,N_43083,N_43896);
nor U44280 (N_44280,N_43526,N_43687);
xnor U44281 (N_44281,N_43660,N_43192);
nand U44282 (N_44282,N_43405,N_43429);
and U44283 (N_44283,N_43831,N_43015);
nand U44284 (N_44284,N_43922,N_43783);
nand U44285 (N_44285,N_43679,N_43758);
xor U44286 (N_44286,N_43024,N_43040);
or U44287 (N_44287,N_43647,N_43118);
nand U44288 (N_44288,N_43908,N_43285);
and U44289 (N_44289,N_43060,N_43250);
nand U44290 (N_44290,N_43496,N_43951);
nor U44291 (N_44291,N_43684,N_43734);
nand U44292 (N_44292,N_43105,N_43322);
nor U44293 (N_44293,N_43220,N_43072);
nand U44294 (N_44294,N_43164,N_43767);
and U44295 (N_44295,N_43445,N_43917);
or U44296 (N_44296,N_43790,N_43812);
or U44297 (N_44297,N_43993,N_43031);
nand U44298 (N_44298,N_43550,N_43378);
nor U44299 (N_44299,N_43744,N_43669);
or U44300 (N_44300,N_43332,N_43599);
or U44301 (N_44301,N_43712,N_43311);
nand U44302 (N_44302,N_43516,N_43335);
xnor U44303 (N_44303,N_43041,N_43503);
xor U44304 (N_44304,N_43860,N_43188);
nand U44305 (N_44305,N_43894,N_43913);
and U44306 (N_44306,N_43324,N_43281);
xnor U44307 (N_44307,N_43113,N_43732);
and U44308 (N_44308,N_43067,N_43423);
nor U44309 (N_44309,N_43286,N_43114);
and U44310 (N_44310,N_43034,N_43969);
xnor U44311 (N_44311,N_43648,N_43383);
xnor U44312 (N_44312,N_43208,N_43275);
and U44313 (N_44313,N_43593,N_43400);
nand U44314 (N_44314,N_43166,N_43221);
nor U44315 (N_44315,N_43672,N_43931);
nor U44316 (N_44316,N_43179,N_43760);
nor U44317 (N_44317,N_43211,N_43959);
xor U44318 (N_44318,N_43885,N_43282);
xor U44319 (N_44319,N_43848,N_43718);
xor U44320 (N_44320,N_43293,N_43654);
and U44321 (N_44321,N_43598,N_43050);
and U44322 (N_44322,N_43032,N_43940);
and U44323 (N_44323,N_43859,N_43136);
nand U44324 (N_44324,N_43391,N_43739);
nor U44325 (N_44325,N_43602,N_43135);
or U44326 (N_44326,N_43187,N_43846);
or U44327 (N_44327,N_43013,N_43095);
xor U44328 (N_44328,N_43028,N_43659);
and U44329 (N_44329,N_43592,N_43414);
or U44330 (N_44330,N_43510,N_43990);
or U44331 (N_44331,N_43631,N_43224);
or U44332 (N_44332,N_43431,N_43731);
or U44333 (N_44333,N_43209,N_43570);
nand U44334 (N_44334,N_43738,N_43596);
nor U44335 (N_44335,N_43983,N_43115);
nand U44336 (N_44336,N_43079,N_43426);
and U44337 (N_44337,N_43566,N_43290);
nand U44338 (N_44338,N_43805,N_43157);
nor U44339 (N_44339,N_43477,N_43724);
and U44340 (N_44340,N_43161,N_43641);
nor U44341 (N_44341,N_43759,N_43688);
nand U44342 (N_44342,N_43439,N_43945);
and U44343 (N_44343,N_43148,N_43506);
nor U44344 (N_44344,N_43425,N_43943);
xnor U44345 (N_44345,N_43747,N_43462);
nand U44346 (N_44346,N_43997,N_43123);
or U44347 (N_44347,N_43256,N_43743);
or U44348 (N_44348,N_43247,N_43251);
nor U44349 (N_44349,N_43177,N_43677);
and U44350 (N_44350,N_43344,N_43160);
nand U44351 (N_44351,N_43956,N_43692);
or U44352 (N_44352,N_43298,N_43263);
or U44353 (N_44353,N_43038,N_43675);
and U44354 (N_44354,N_43719,N_43017);
xnor U44355 (N_44355,N_43336,N_43051);
xor U44356 (N_44356,N_43312,N_43556);
xnor U44357 (N_44357,N_43553,N_43386);
nor U44358 (N_44358,N_43321,N_43965);
xor U44359 (N_44359,N_43236,N_43066);
xnor U44360 (N_44360,N_43055,N_43664);
xnor U44361 (N_44361,N_43004,N_43222);
nor U44362 (N_44362,N_43093,N_43775);
xnor U44363 (N_44363,N_43857,N_43957);
or U44364 (N_44364,N_43795,N_43610);
nand U44365 (N_44365,N_43781,N_43156);
nor U44366 (N_44366,N_43338,N_43490);
nand U44367 (N_44367,N_43084,N_43370);
and U44368 (N_44368,N_43165,N_43852);
or U44369 (N_44369,N_43158,N_43356);
or U44370 (N_44370,N_43292,N_43707);
nor U44371 (N_44371,N_43181,N_43459);
and U44372 (N_44372,N_43101,N_43392);
and U44373 (N_44373,N_43950,N_43683);
nor U44374 (N_44374,N_43348,N_43228);
or U44375 (N_44375,N_43305,N_43364);
nor U44376 (N_44376,N_43827,N_43091);
nor U44377 (N_44377,N_43053,N_43037);
nor U44378 (N_44378,N_43914,N_43748);
nand U44379 (N_44379,N_43560,N_43197);
nor U44380 (N_44380,N_43200,N_43927);
nor U44381 (N_44381,N_43482,N_43387);
and U44382 (N_44382,N_43721,N_43399);
nand U44383 (N_44383,N_43063,N_43862);
or U44384 (N_44384,N_43773,N_43403);
xnor U44385 (N_44385,N_43058,N_43107);
or U44386 (N_44386,N_43433,N_43241);
or U44387 (N_44387,N_43868,N_43873);
and U44388 (N_44388,N_43449,N_43682);
or U44389 (N_44389,N_43390,N_43196);
xor U44390 (N_44390,N_43430,N_43455);
nand U44391 (N_44391,N_43865,N_43180);
xnor U44392 (N_44392,N_43920,N_43634);
or U44393 (N_44393,N_43979,N_43521);
or U44394 (N_44394,N_43733,N_43394);
or U44395 (N_44395,N_43304,N_43730);
or U44396 (N_44396,N_43753,N_43963);
xor U44397 (N_44397,N_43195,N_43653);
nand U44398 (N_44398,N_43474,N_43600);
nand U44399 (N_44399,N_43147,N_43996);
or U44400 (N_44400,N_43854,N_43471);
and U44401 (N_44401,N_43260,N_43595);
or U44402 (N_44402,N_43346,N_43210);
xor U44403 (N_44403,N_43495,N_43725);
and U44404 (N_44404,N_43589,N_43944);
nor U44405 (N_44405,N_43934,N_43946);
nand U44406 (N_44406,N_43475,N_43924);
nand U44407 (N_44407,N_43750,N_43668);
and U44408 (N_44408,N_43749,N_43636);
or U44409 (N_44409,N_43884,N_43457);
and U44410 (N_44410,N_43863,N_43481);
nor U44411 (N_44411,N_43049,N_43493);
nor U44412 (N_44412,N_43129,N_43340);
or U44413 (N_44413,N_43938,N_43308);
and U44414 (N_44414,N_43821,N_43092);
nor U44415 (N_44415,N_43849,N_43840);
nand U44416 (N_44416,N_43014,N_43094);
nand U44417 (N_44417,N_43887,N_43637);
and U44418 (N_44418,N_43121,N_43923);
or U44419 (N_44419,N_43141,N_43427);
nand U44420 (N_44420,N_43976,N_43194);
and U44421 (N_44421,N_43143,N_43706);
nor U44422 (N_44422,N_43778,N_43531);
or U44423 (N_44423,N_43265,N_43694);
xor U44424 (N_44424,N_43358,N_43169);
nand U44425 (N_44425,N_43799,N_43219);
xor U44426 (N_44426,N_43003,N_43801);
xnor U44427 (N_44427,N_43581,N_43897);
nand U44428 (N_44428,N_43059,N_43088);
and U44429 (N_44429,N_43832,N_43484);
nor U44430 (N_44430,N_43144,N_43119);
xnor U44431 (N_44431,N_43752,N_43205);
nor U44432 (N_44432,N_43557,N_43206);
nand U44433 (N_44433,N_43947,N_43693);
or U44434 (N_44434,N_43740,N_43613);
or U44435 (N_44435,N_43699,N_43329);
nand U44436 (N_44436,N_43685,N_43649);
xnor U44437 (N_44437,N_43233,N_43797);
nor U44438 (N_44438,N_43327,N_43547);
nand U44439 (N_44439,N_43314,N_43980);
nand U44440 (N_44440,N_43277,N_43479);
and U44441 (N_44441,N_43300,N_43411);
nand U44442 (N_44442,N_43879,N_43834);
nor U44443 (N_44443,N_43658,N_43458);
xnor U44444 (N_44444,N_43559,N_43389);
nor U44445 (N_44445,N_43489,N_43190);
or U44446 (N_44446,N_43149,N_43244);
nand U44447 (N_44447,N_43082,N_43000);
and U44448 (N_44448,N_43576,N_43513);
nor U44449 (N_44449,N_43890,N_43509);
nand U44450 (N_44450,N_43424,N_43096);
xnor U44451 (N_44451,N_43369,N_43274);
nor U44452 (N_44452,N_43417,N_43872);
and U44453 (N_44453,N_43159,N_43026);
or U44454 (N_44454,N_43374,N_43152);
xnor U44455 (N_44455,N_43893,N_43398);
nand U44456 (N_44456,N_43800,N_43345);
xor U44457 (N_44457,N_43085,N_43362);
nor U44458 (N_44458,N_43467,N_43440);
xor U44459 (N_44459,N_43173,N_43213);
xnor U44460 (N_44460,N_43020,N_43820);
xnor U44461 (N_44461,N_43046,N_43847);
or U44462 (N_44462,N_43629,N_43549);
nor U44463 (N_44463,N_43655,N_43235);
nor U44464 (N_44464,N_43841,N_43178);
nand U44465 (N_44465,N_43379,N_43184);
nand U44466 (N_44466,N_43048,N_43432);
or U44467 (N_44467,N_43665,N_43579);
or U44468 (N_44468,N_43502,N_43616);
nor U44469 (N_44469,N_43264,N_43717);
nand U44470 (N_44470,N_43791,N_43333);
nand U44471 (N_44471,N_43786,N_43789);
and U44472 (N_44472,N_43201,N_43102);
nor U44473 (N_44473,N_43925,N_43249);
xnor U44474 (N_44474,N_43823,N_43845);
or U44475 (N_44475,N_43714,N_43962);
or U44476 (N_44476,N_43994,N_43316);
or U44477 (N_44477,N_43207,N_43483);
nand U44478 (N_44478,N_43511,N_43585);
nand U44479 (N_44479,N_43486,N_43817);
nor U44480 (N_44480,N_43933,N_43782);
nand U44481 (N_44481,N_43372,N_43632);
or U44482 (N_44482,N_43763,N_43704);
and U44483 (N_44483,N_43122,N_43543);
xor U44484 (N_44484,N_43448,N_43524);
or U44485 (N_44485,N_43711,N_43701);
nor U44486 (N_44486,N_43385,N_43488);
and U44487 (N_44487,N_43042,N_43607);
or U44488 (N_44488,N_43824,N_43125);
or U44489 (N_44489,N_43401,N_43350);
nor U44490 (N_44490,N_43614,N_43112);
and U44491 (N_44491,N_43736,N_43396);
nor U44492 (N_44492,N_43981,N_43615);
nand U44493 (N_44493,N_43357,N_43319);
or U44494 (N_44494,N_43545,N_43074);
or U44495 (N_44495,N_43535,N_43808);
nor U44496 (N_44496,N_43624,N_43284);
or U44497 (N_44497,N_43895,N_43296);
and U44498 (N_44498,N_43844,N_43638);
nor U44499 (N_44499,N_43262,N_43142);
xor U44500 (N_44500,N_43637,N_43451);
or U44501 (N_44501,N_43359,N_43092);
xor U44502 (N_44502,N_43069,N_43595);
nor U44503 (N_44503,N_43087,N_43440);
and U44504 (N_44504,N_43930,N_43254);
xnor U44505 (N_44505,N_43277,N_43088);
or U44506 (N_44506,N_43170,N_43129);
nor U44507 (N_44507,N_43806,N_43940);
nand U44508 (N_44508,N_43981,N_43326);
or U44509 (N_44509,N_43138,N_43344);
nor U44510 (N_44510,N_43919,N_43804);
or U44511 (N_44511,N_43247,N_43035);
nor U44512 (N_44512,N_43535,N_43673);
nor U44513 (N_44513,N_43528,N_43329);
nand U44514 (N_44514,N_43240,N_43562);
and U44515 (N_44515,N_43895,N_43960);
nand U44516 (N_44516,N_43571,N_43599);
or U44517 (N_44517,N_43289,N_43508);
xnor U44518 (N_44518,N_43208,N_43013);
or U44519 (N_44519,N_43201,N_43293);
nand U44520 (N_44520,N_43294,N_43757);
xnor U44521 (N_44521,N_43131,N_43512);
xor U44522 (N_44522,N_43477,N_43917);
or U44523 (N_44523,N_43246,N_43187);
nand U44524 (N_44524,N_43238,N_43884);
and U44525 (N_44525,N_43463,N_43302);
xnor U44526 (N_44526,N_43557,N_43052);
xor U44527 (N_44527,N_43278,N_43792);
and U44528 (N_44528,N_43551,N_43090);
nand U44529 (N_44529,N_43901,N_43829);
or U44530 (N_44530,N_43855,N_43857);
or U44531 (N_44531,N_43679,N_43461);
nor U44532 (N_44532,N_43641,N_43494);
nand U44533 (N_44533,N_43025,N_43449);
nand U44534 (N_44534,N_43430,N_43370);
nand U44535 (N_44535,N_43081,N_43396);
nand U44536 (N_44536,N_43371,N_43064);
nand U44537 (N_44537,N_43617,N_43286);
nand U44538 (N_44538,N_43658,N_43991);
xnor U44539 (N_44539,N_43319,N_43293);
nor U44540 (N_44540,N_43966,N_43324);
xnor U44541 (N_44541,N_43855,N_43209);
nand U44542 (N_44542,N_43042,N_43418);
or U44543 (N_44543,N_43103,N_43869);
xor U44544 (N_44544,N_43919,N_43681);
nor U44545 (N_44545,N_43179,N_43349);
xor U44546 (N_44546,N_43462,N_43215);
xor U44547 (N_44547,N_43496,N_43624);
and U44548 (N_44548,N_43820,N_43689);
nand U44549 (N_44549,N_43813,N_43248);
xnor U44550 (N_44550,N_43958,N_43212);
nor U44551 (N_44551,N_43317,N_43460);
and U44552 (N_44552,N_43824,N_43949);
nand U44553 (N_44553,N_43214,N_43201);
or U44554 (N_44554,N_43412,N_43760);
xnor U44555 (N_44555,N_43761,N_43045);
and U44556 (N_44556,N_43858,N_43573);
nor U44557 (N_44557,N_43738,N_43607);
xor U44558 (N_44558,N_43265,N_43180);
nor U44559 (N_44559,N_43300,N_43677);
nand U44560 (N_44560,N_43510,N_43925);
and U44561 (N_44561,N_43910,N_43639);
nand U44562 (N_44562,N_43771,N_43239);
or U44563 (N_44563,N_43507,N_43016);
nor U44564 (N_44564,N_43534,N_43025);
or U44565 (N_44565,N_43673,N_43507);
and U44566 (N_44566,N_43897,N_43605);
or U44567 (N_44567,N_43226,N_43748);
xnor U44568 (N_44568,N_43307,N_43162);
nor U44569 (N_44569,N_43502,N_43565);
xor U44570 (N_44570,N_43515,N_43961);
and U44571 (N_44571,N_43919,N_43990);
or U44572 (N_44572,N_43781,N_43723);
xnor U44573 (N_44573,N_43229,N_43213);
and U44574 (N_44574,N_43061,N_43249);
nor U44575 (N_44575,N_43197,N_43564);
and U44576 (N_44576,N_43643,N_43391);
xor U44577 (N_44577,N_43348,N_43051);
nor U44578 (N_44578,N_43202,N_43055);
nand U44579 (N_44579,N_43382,N_43303);
or U44580 (N_44580,N_43929,N_43844);
xor U44581 (N_44581,N_43489,N_43957);
and U44582 (N_44582,N_43942,N_43547);
and U44583 (N_44583,N_43852,N_43244);
nand U44584 (N_44584,N_43805,N_43670);
nand U44585 (N_44585,N_43787,N_43899);
and U44586 (N_44586,N_43639,N_43036);
or U44587 (N_44587,N_43156,N_43522);
nand U44588 (N_44588,N_43314,N_43498);
or U44589 (N_44589,N_43554,N_43942);
nor U44590 (N_44590,N_43734,N_43819);
and U44591 (N_44591,N_43848,N_43000);
or U44592 (N_44592,N_43849,N_43678);
and U44593 (N_44593,N_43334,N_43410);
xor U44594 (N_44594,N_43108,N_43710);
nor U44595 (N_44595,N_43563,N_43694);
and U44596 (N_44596,N_43124,N_43395);
nand U44597 (N_44597,N_43932,N_43163);
nor U44598 (N_44598,N_43538,N_43467);
nor U44599 (N_44599,N_43367,N_43287);
and U44600 (N_44600,N_43099,N_43153);
nand U44601 (N_44601,N_43741,N_43740);
and U44602 (N_44602,N_43355,N_43714);
xnor U44603 (N_44603,N_43359,N_43475);
nor U44604 (N_44604,N_43481,N_43373);
nand U44605 (N_44605,N_43624,N_43592);
xnor U44606 (N_44606,N_43880,N_43065);
or U44607 (N_44607,N_43934,N_43942);
xnor U44608 (N_44608,N_43730,N_43768);
nand U44609 (N_44609,N_43676,N_43165);
nand U44610 (N_44610,N_43540,N_43696);
xnor U44611 (N_44611,N_43711,N_43074);
nor U44612 (N_44612,N_43359,N_43264);
nor U44613 (N_44613,N_43017,N_43891);
and U44614 (N_44614,N_43385,N_43775);
and U44615 (N_44615,N_43930,N_43676);
xnor U44616 (N_44616,N_43825,N_43051);
or U44617 (N_44617,N_43548,N_43418);
and U44618 (N_44618,N_43678,N_43623);
or U44619 (N_44619,N_43292,N_43865);
xnor U44620 (N_44620,N_43163,N_43844);
or U44621 (N_44621,N_43114,N_43350);
nand U44622 (N_44622,N_43630,N_43588);
and U44623 (N_44623,N_43820,N_43522);
nand U44624 (N_44624,N_43076,N_43458);
and U44625 (N_44625,N_43512,N_43187);
nor U44626 (N_44626,N_43907,N_43683);
nand U44627 (N_44627,N_43254,N_43886);
nor U44628 (N_44628,N_43016,N_43442);
nor U44629 (N_44629,N_43694,N_43890);
nor U44630 (N_44630,N_43976,N_43266);
xnor U44631 (N_44631,N_43846,N_43964);
nand U44632 (N_44632,N_43455,N_43591);
or U44633 (N_44633,N_43405,N_43068);
nor U44634 (N_44634,N_43679,N_43837);
xnor U44635 (N_44635,N_43276,N_43308);
xor U44636 (N_44636,N_43341,N_43045);
nor U44637 (N_44637,N_43230,N_43537);
nand U44638 (N_44638,N_43441,N_43700);
nor U44639 (N_44639,N_43273,N_43318);
nor U44640 (N_44640,N_43614,N_43219);
nor U44641 (N_44641,N_43844,N_43536);
nand U44642 (N_44642,N_43267,N_43350);
and U44643 (N_44643,N_43204,N_43772);
nor U44644 (N_44644,N_43571,N_43573);
and U44645 (N_44645,N_43522,N_43884);
xnor U44646 (N_44646,N_43722,N_43131);
nand U44647 (N_44647,N_43536,N_43865);
nor U44648 (N_44648,N_43173,N_43147);
nand U44649 (N_44649,N_43022,N_43867);
or U44650 (N_44650,N_43926,N_43463);
nor U44651 (N_44651,N_43051,N_43663);
nand U44652 (N_44652,N_43058,N_43804);
nand U44653 (N_44653,N_43948,N_43975);
and U44654 (N_44654,N_43614,N_43296);
nand U44655 (N_44655,N_43016,N_43566);
and U44656 (N_44656,N_43329,N_43681);
or U44657 (N_44657,N_43737,N_43081);
nand U44658 (N_44658,N_43167,N_43786);
nor U44659 (N_44659,N_43422,N_43194);
and U44660 (N_44660,N_43034,N_43298);
nand U44661 (N_44661,N_43064,N_43354);
nand U44662 (N_44662,N_43673,N_43633);
nand U44663 (N_44663,N_43727,N_43515);
xnor U44664 (N_44664,N_43691,N_43167);
or U44665 (N_44665,N_43164,N_43728);
and U44666 (N_44666,N_43985,N_43001);
and U44667 (N_44667,N_43062,N_43761);
or U44668 (N_44668,N_43447,N_43324);
nand U44669 (N_44669,N_43687,N_43173);
and U44670 (N_44670,N_43053,N_43308);
nor U44671 (N_44671,N_43632,N_43931);
or U44672 (N_44672,N_43112,N_43908);
nor U44673 (N_44673,N_43791,N_43571);
xor U44674 (N_44674,N_43143,N_43624);
and U44675 (N_44675,N_43302,N_43574);
nor U44676 (N_44676,N_43765,N_43433);
xor U44677 (N_44677,N_43933,N_43629);
and U44678 (N_44678,N_43440,N_43565);
xor U44679 (N_44679,N_43760,N_43690);
xor U44680 (N_44680,N_43450,N_43393);
or U44681 (N_44681,N_43709,N_43319);
xnor U44682 (N_44682,N_43292,N_43133);
and U44683 (N_44683,N_43304,N_43635);
or U44684 (N_44684,N_43526,N_43189);
nor U44685 (N_44685,N_43919,N_43385);
nand U44686 (N_44686,N_43194,N_43699);
xor U44687 (N_44687,N_43863,N_43273);
nand U44688 (N_44688,N_43960,N_43715);
or U44689 (N_44689,N_43633,N_43197);
xnor U44690 (N_44690,N_43181,N_43331);
nand U44691 (N_44691,N_43128,N_43060);
nor U44692 (N_44692,N_43150,N_43748);
or U44693 (N_44693,N_43298,N_43328);
and U44694 (N_44694,N_43873,N_43923);
and U44695 (N_44695,N_43015,N_43193);
or U44696 (N_44696,N_43052,N_43922);
nor U44697 (N_44697,N_43681,N_43966);
nor U44698 (N_44698,N_43734,N_43727);
and U44699 (N_44699,N_43661,N_43393);
xnor U44700 (N_44700,N_43030,N_43650);
or U44701 (N_44701,N_43372,N_43762);
and U44702 (N_44702,N_43278,N_43928);
nor U44703 (N_44703,N_43213,N_43584);
and U44704 (N_44704,N_43796,N_43788);
xnor U44705 (N_44705,N_43745,N_43054);
nand U44706 (N_44706,N_43696,N_43962);
xor U44707 (N_44707,N_43995,N_43105);
nor U44708 (N_44708,N_43116,N_43825);
nor U44709 (N_44709,N_43542,N_43495);
nand U44710 (N_44710,N_43073,N_43817);
nor U44711 (N_44711,N_43752,N_43917);
or U44712 (N_44712,N_43703,N_43466);
nor U44713 (N_44713,N_43199,N_43050);
nand U44714 (N_44714,N_43198,N_43101);
nand U44715 (N_44715,N_43716,N_43194);
nor U44716 (N_44716,N_43347,N_43223);
nand U44717 (N_44717,N_43861,N_43678);
xor U44718 (N_44718,N_43213,N_43849);
nor U44719 (N_44719,N_43788,N_43933);
nor U44720 (N_44720,N_43869,N_43180);
or U44721 (N_44721,N_43265,N_43629);
nand U44722 (N_44722,N_43404,N_43433);
nand U44723 (N_44723,N_43842,N_43279);
nand U44724 (N_44724,N_43946,N_43466);
nor U44725 (N_44725,N_43713,N_43671);
xor U44726 (N_44726,N_43166,N_43896);
or U44727 (N_44727,N_43249,N_43334);
or U44728 (N_44728,N_43727,N_43614);
and U44729 (N_44729,N_43762,N_43979);
nor U44730 (N_44730,N_43964,N_43677);
nand U44731 (N_44731,N_43775,N_43112);
nor U44732 (N_44732,N_43732,N_43326);
or U44733 (N_44733,N_43371,N_43265);
nor U44734 (N_44734,N_43175,N_43600);
and U44735 (N_44735,N_43859,N_43333);
or U44736 (N_44736,N_43022,N_43665);
nand U44737 (N_44737,N_43562,N_43733);
xnor U44738 (N_44738,N_43330,N_43840);
xnor U44739 (N_44739,N_43051,N_43581);
or U44740 (N_44740,N_43186,N_43531);
nor U44741 (N_44741,N_43971,N_43183);
nor U44742 (N_44742,N_43196,N_43509);
nand U44743 (N_44743,N_43309,N_43848);
xnor U44744 (N_44744,N_43306,N_43317);
xor U44745 (N_44745,N_43377,N_43802);
and U44746 (N_44746,N_43280,N_43949);
nand U44747 (N_44747,N_43877,N_43527);
or U44748 (N_44748,N_43101,N_43102);
and U44749 (N_44749,N_43468,N_43007);
nand U44750 (N_44750,N_43702,N_43348);
nand U44751 (N_44751,N_43683,N_43522);
or U44752 (N_44752,N_43550,N_43129);
and U44753 (N_44753,N_43474,N_43793);
nand U44754 (N_44754,N_43449,N_43387);
xnor U44755 (N_44755,N_43696,N_43672);
and U44756 (N_44756,N_43502,N_43973);
nor U44757 (N_44757,N_43158,N_43962);
nor U44758 (N_44758,N_43902,N_43799);
nor U44759 (N_44759,N_43187,N_43548);
xnor U44760 (N_44760,N_43063,N_43020);
xnor U44761 (N_44761,N_43304,N_43362);
xor U44762 (N_44762,N_43515,N_43209);
xnor U44763 (N_44763,N_43325,N_43234);
nand U44764 (N_44764,N_43098,N_43101);
nand U44765 (N_44765,N_43192,N_43236);
and U44766 (N_44766,N_43577,N_43712);
nand U44767 (N_44767,N_43497,N_43749);
or U44768 (N_44768,N_43148,N_43869);
nor U44769 (N_44769,N_43592,N_43929);
and U44770 (N_44770,N_43101,N_43386);
nor U44771 (N_44771,N_43452,N_43898);
nand U44772 (N_44772,N_43999,N_43448);
or U44773 (N_44773,N_43078,N_43993);
nor U44774 (N_44774,N_43175,N_43232);
and U44775 (N_44775,N_43615,N_43104);
nor U44776 (N_44776,N_43478,N_43777);
nor U44777 (N_44777,N_43291,N_43502);
nand U44778 (N_44778,N_43910,N_43431);
or U44779 (N_44779,N_43003,N_43894);
and U44780 (N_44780,N_43602,N_43585);
nand U44781 (N_44781,N_43904,N_43832);
nand U44782 (N_44782,N_43236,N_43777);
and U44783 (N_44783,N_43357,N_43724);
xnor U44784 (N_44784,N_43426,N_43815);
nand U44785 (N_44785,N_43983,N_43662);
and U44786 (N_44786,N_43302,N_43879);
and U44787 (N_44787,N_43827,N_43887);
nor U44788 (N_44788,N_43788,N_43983);
or U44789 (N_44789,N_43459,N_43138);
and U44790 (N_44790,N_43528,N_43250);
nand U44791 (N_44791,N_43547,N_43053);
xor U44792 (N_44792,N_43271,N_43311);
and U44793 (N_44793,N_43769,N_43497);
or U44794 (N_44794,N_43474,N_43212);
or U44795 (N_44795,N_43273,N_43083);
xnor U44796 (N_44796,N_43559,N_43737);
nor U44797 (N_44797,N_43511,N_43277);
xnor U44798 (N_44798,N_43765,N_43887);
or U44799 (N_44799,N_43608,N_43354);
xor U44800 (N_44800,N_43801,N_43882);
and U44801 (N_44801,N_43877,N_43859);
nand U44802 (N_44802,N_43324,N_43777);
nor U44803 (N_44803,N_43414,N_43602);
xnor U44804 (N_44804,N_43132,N_43242);
xor U44805 (N_44805,N_43953,N_43673);
or U44806 (N_44806,N_43078,N_43829);
or U44807 (N_44807,N_43157,N_43419);
nand U44808 (N_44808,N_43680,N_43977);
nand U44809 (N_44809,N_43887,N_43657);
xor U44810 (N_44810,N_43003,N_43007);
or U44811 (N_44811,N_43176,N_43609);
nand U44812 (N_44812,N_43456,N_43649);
nand U44813 (N_44813,N_43682,N_43595);
xnor U44814 (N_44814,N_43227,N_43090);
or U44815 (N_44815,N_43537,N_43307);
or U44816 (N_44816,N_43504,N_43709);
nand U44817 (N_44817,N_43272,N_43380);
and U44818 (N_44818,N_43923,N_43038);
and U44819 (N_44819,N_43379,N_43886);
and U44820 (N_44820,N_43008,N_43761);
nor U44821 (N_44821,N_43840,N_43613);
nor U44822 (N_44822,N_43755,N_43773);
xor U44823 (N_44823,N_43774,N_43419);
nand U44824 (N_44824,N_43165,N_43542);
or U44825 (N_44825,N_43104,N_43766);
and U44826 (N_44826,N_43001,N_43958);
nand U44827 (N_44827,N_43517,N_43459);
nor U44828 (N_44828,N_43281,N_43385);
nand U44829 (N_44829,N_43729,N_43635);
nand U44830 (N_44830,N_43242,N_43627);
or U44831 (N_44831,N_43179,N_43806);
nand U44832 (N_44832,N_43448,N_43823);
nor U44833 (N_44833,N_43273,N_43878);
nand U44834 (N_44834,N_43624,N_43477);
nand U44835 (N_44835,N_43890,N_43193);
or U44836 (N_44836,N_43203,N_43959);
nand U44837 (N_44837,N_43285,N_43599);
xor U44838 (N_44838,N_43103,N_43373);
nand U44839 (N_44839,N_43956,N_43386);
or U44840 (N_44840,N_43598,N_43585);
and U44841 (N_44841,N_43704,N_43513);
nor U44842 (N_44842,N_43980,N_43603);
nor U44843 (N_44843,N_43841,N_43951);
and U44844 (N_44844,N_43662,N_43367);
nor U44845 (N_44845,N_43244,N_43493);
or U44846 (N_44846,N_43476,N_43917);
and U44847 (N_44847,N_43297,N_43057);
xor U44848 (N_44848,N_43325,N_43369);
nand U44849 (N_44849,N_43117,N_43160);
and U44850 (N_44850,N_43602,N_43679);
xor U44851 (N_44851,N_43471,N_43470);
or U44852 (N_44852,N_43403,N_43717);
and U44853 (N_44853,N_43556,N_43843);
or U44854 (N_44854,N_43897,N_43241);
xor U44855 (N_44855,N_43925,N_43356);
or U44856 (N_44856,N_43967,N_43571);
and U44857 (N_44857,N_43996,N_43405);
nor U44858 (N_44858,N_43912,N_43501);
or U44859 (N_44859,N_43985,N_43839);
nor U44860 (N_44860,N_43207,N_43585);
or U44861 (N_44861,N_43577,N_43046);
or U44862 (N_44862,N_43529,N_43575);
xor U44863 (N_44863,N_43515,N_43114);
and U44864 (N_44864,N_43061,N_43456);
nand U44865 (N_44865,N_43775,N_43863);
and U44866 (N_44866,N_43918,N_43954);
and U44867 (N_44867,N_43539,N_43656);
and U44868 (N_44868,N_43696,N_43933);
or U44869 (N_44869,N_43473,N_43449);
nor U44870 (N_44870,N_43061,N_43844);
nand U44871 (N_44871,N_43767,N_43992);
and U44872 (N_44872,N_43987,N_43435);
and U44873 (N_44873,N_43464,N_43297);
xor U44874 (N_44874,N_43788,N_43046);
xor U44875 (N_44875,N_43881,N_43562);
nand U44876 (N_44876,N_43478,N_43812);
or U44877 (N_44877,N_43172,N_43054);
and U44878 (N_44878,N_43626,N_43694);
nand U44879 (N_44879,N_43136,N_43640);
and U44880 (N_44880,N_43935,N_43407);
nand U44881 (N_44881,N_43929,N_43015);
xnor U44882 (N_44882,N_43916,N_43430);
or U44883 (N_44883,N_43486,N_43612);
or U44884 (N_44884,N_43112,N_43261);
and U44885 (N_44885,N_43485,N_43858);
and U44886 (N_44886,N_43015,N_43411);
xor U44887 (N_44887,N_43516,N_43083);
xnor U44888 (N_44888,N_43564,N_43620);
or U44889 (N_44889,N_43425,N_43992);
nand U44890 (N_44890,N_43875,N_43902);
or U44891 (N_44891,N_43592,N_43768);
and U44892 (N_44892,N_43746,N_43927);
nand U44893 (N_44893,N_43971,N_43006);
and U44894 (N_44894,N_43501,N_43222);
nand U44895 (N_44895,N_43870,N_43205);
or U44896 (N_44896,N_43308,N_43421);
and U44897 (N_44897,N_43339,N_43307);
xor U44898 (N_44898,N_43974,N_43686);
or U44899 (N_44899,N_43724,N_43699);
nand U44900 (N_44900,N_43146,N_43733);
nor U44901 (N_44901,N_43920,N_43621);
nand U44902 (N_44902,N_43197,N_43320);
or U44903 (N_44903,N_43852,N_43153);
or U44904 (N_44904,N_43434,N_43840);
nand U44905 (N_44905,N_43936,N_43155);
and U44906 (N_44906,N_43669,N_43899);
and U44907 (N_44907,N_43363,N_43010);
nor U44908 (N_44908,N_43263,N_43210);
nand U44909 (N_44909,N_43716,N_43890);
nor U44910 (N_44910,N_43581,N_43005);
nor U44911 (N_44911,N_43096,N_43858);
xor U44912 (N_44912,N_43572,N_43125);
nand U44913 (N_44913,N_43312,N_43477);
nor U44914 (N_44914,N_43677,N_43740);
nor U44915 (N_44915,N_43846,N_43836);
nor U44916 (N_44916,N_43577,N_43258);
xnor U44917 (N_44917,N_43879,N_43414);
and U44918 (N_44918,N_43982,N_43288);
xnor U44919 (N_44919,N_43781,N_43768);
nand U44920 (N_44920,N_43110,N_43468);
nor U44921 (N_44921,N_43591,N_43174);
or U44922 (N_44922,N_43503,N_43084);
and U44923 (N_44923,N_43031,N_43110);
nor U44924 (N_44924,N_43074,N_43323);
and U44925 (N_44925,N_43428,N_43532);
and U44926 (N_44926,N_43565,N_43528);
nor U44927 (N_44927,N_43073,N_43079);
or U44928 (N_44928,N_43795,N_43107);
xor U44929 (N_44929,N_43019,N_43632);
nand U44930 (N_44930,N_43506,N_43018);
or U44931 (N_44931,N_43572,N_43552);
nor U44932 (N_44932,N_43711,N_43106);
nor U44933 (N_44933,N_43185,N_43611);
nand U44934 (N_44934,N_43241,N_43343);
or U44935 (N_44935,N_43936,N_43474);
nor U44936 (N_44936,N_43196,N_43426);
and U44937 (N_44937,N_43532,N_43234);
nand U44938 (N_44938,N_43704,N_43449);
and U44939 (N_44939,N_43577,N_43579);
xor U44940 (N_44940,N_43863,N_43682);
and U44941 (N_44941,N_43412,N_43448);
nand U44942 (N_44942,N_43536,N_43347);
xor U44943 (N_44943,N_43386,N_43051);
and U44944 (N_44944,N_43660,N_43035);
and U44945 (N_44945,N_43011,N_43340);
xnor U44946 (N_44946,N_43255,N_43404);
xnor U44947 (N_44947,N_43875,N_43660);
nand U44948 (N_44948,N_43748,N_43510);
nor U44949 (N_44949,N_43722,N_43652);
nor U44950 (N_44950,N_43372,N_43054);
xnor U44951 (N_44951,N_43592,N_43154);
xnor U44952 (N_44952,N_43318,N_43796);
or U44953 (N_44953,N_43571,N_43060);
xor U44954 (N_44954,N_43258,N_43436);
xnor U44955 (N_44955,N_43871,N_43406);
nand U44956 (N_44956,N_43335,N_43660);
or U44957 (N_44957,N_43912,N_43457);
xor U44958 (N_44958,N_43598,N_43560);
nor U44959 (N_44959,N_43196,N_43413);
and U44960 (N_44960,N_43618,N_43455);
and U44961 (N_44961,N_43322,N_43242);
nor U44962 (N_44962,N_43500,N_43493);
nor U44963 (N_44963,N_43878,N_43508);
xor U44964 (N_44964,N_43850,N_43270);
xnor U44965 (N_44965,N_43821,N_43245);
xnor U44966 (N_44966,N_43091,N_43732);
or U44967 (N_44967,N_43185,N_43294);
xor U44968 (N_44968,N_43961,N_43369);
or U44969 (N_44969,N_43259,N_43627);
xor U44970 (N_44970,N_43259,N_43205);
xnor U44971 (N_44971,N_43825,N_43105);
or U44972 (N_44972,N_43880,N_43489);
nor U44973 (N_44973,N_43373,N_43139);
xnor U44974 (N_44974,N_43060,N_43553);
nor U44975 (N_44975,N_43488,N_43647);
or U44976 (N_44976,N_43325,N_43456);
nand U44977 (N_44977,N_43162,N_43598);
xor U44978 (N_44978,N_43157,N_43243);
nand U44979 (N_44979,N_43987,N_43166);
nor U44980 (N_44980,N_43558,N_43613);
and U44981 (N_44981,N_43898,N_43168);
and U44982 (N_44982,N_43332,N_43134);
nand U44983 (N_44983,N_43134,N_43604);
xnor U44984 (N_44984,N_43573,N_43112);
or U44985 (N_44985,N_43710,N_43884);
xor U44986 (N_44986,N_43992,N_43230);
nand U44987 (N_44987,N_43837,N_43587);
nor U44988 (N_44988,N_43052,N_43128);
and U44989 (N_44989,N_43278,N_43575);
or U44990 (N_44990,N_43105,N_43339);
nor U44991 (N_44991,N_43139,N_43132);
nor U44992 (N_44992,N_43207,N_43464);
or U44993 (N_44993,N_43321,N_43153);
xor U44994 (N_44994,N_43998,N_43860);
nand U44995 (N_44995,N_43935,N_43201);
nor U44996 (N_44996,N_43555,N_43877);
or U44997 (N_44997,N_43947,N_43251);
nand U44998 (N_44998,N_43051,N_43234);
nand U44999 (N_44999,N_43157,N_43937);
and U45000 (N_45000,N_44157,N_44768);
xor U45001 (N_45001,N_44687,N_44518);
xor U45002 (N_45002,N_44373,N_44326);
nor U45003 (N_45003,N_44495,N_44023);
nand U45004 (N_45004,N_44880,N_44771);
xnor U45005 (N_45005,N_44058,N_44201);
xnor U45006 (N_45006,N_44836,N_44904);
nand U45007 (N_45007,N_44247,N_44934);
and U45008 (N_45008,N_44966,N_44388);
and U45009 (N_45009,N_44869,N_44362);
or U45010 (N_45010,N_44781,N_44586);
and U45011 (N_45011,N_44713,N_44856);
xnor U45012 (N_45012,N_44772,N_44973);
or U45013 (N_45013,N_44867,N_44814);
and U45014 (N_45014,N_44854,N_44722);
xor U45015 (N_45015,N_44677,N_44892);
xor U45016 (N_45016,N_44274,N_44923);
nand U45017 (N_45017,N_44801,N_44327);
nor U45018 (N_45018,N_44844,N_44858);
and U45019 (N_45019,N_44673,N_44523);
or U45020 (N_45020,N_44669,N_44271);
xnor U45021 (N_45021,N_44333,N_44580);
and U45022 (N_45022,N_44114,N_44736);
xor U45023 (N_45023,N_44576,N_44916);
xnor U45024 (N_45024,N_44967,N_44453);
and U45025 (N_45025,N_44188,N_44016);
and U45026 (N_45026,N_44012,N_44314);
xor U45027 (N_45027,N_44600,N_44778);
xnor U45028 (N_45028,N_44352,N_44659);
and U45029 (N_45029,N_44229,N_44076);
nor U45030 (N_45030,N_44479,N_44286);
or U45031 (N_45031,N_44273,N_44711);
nand U45032 (N_45032,N_44275,N_44172);
nor U45033 (N_45033,N_44281,N_44402);
nand U45034 (N_45034,N_44039,N_44666);
xor U45035 (N_45035,N_44958,N_44884);
or U45036 (N_45036,N_44979,N_44940);
and U45037 (N_45037,N_44443,N_44227);
or U45038 (N_45038,N_44387,N_44099);
xor U45039 (N_45039,N_44299,N_44897);
nand U45040 (N_45040,N_44661,N_44716);
and U45041 (N_45041,N_44725,N_44888);
nor U45042 (N_45042,N_44260,N_44040);
or U45043 (N_45043,N_44909,N_44168);
and U45044 (N_45044,N_44835,N_44493);
and U45045 (N_45045,N_44862,N_44700);
or U45046 (N_45046,N_44442,N_44970);
nor U45047 (N_45047,N_44246,N_44968);
nor U45048 (N_45048,N_44222,N_44054);
nand U45049 (N_45049,N_44633,N_44512);
nor U45050 (N_45050,N_44432,N_44338);
nand U45051 (N_45051,N_44151,N_44808);
nand U45052 (N_45052,N_44800,N_44935);
xor U45053 (N_45053,N_44385,N_44397);
or U45054 (N_45054,N_44845,N_44186);
or U45055 (N_45055,N_44256,N_44272);
nand U45056 (N_45056,N_44573,N_44115);
nor U45057 (N_45057,N_44461,N_44637);
nand U45058 (N_45058,N_44320,N_44582);
or U45059 (N_45059,N_44851,N_44235);
or U45060 (N_45060,N_44802,N_44462);
nor U45061 (N_45061,N_44564,N_44568);
nand U45062 (N_45062,N_44008,N_44507);
nand U45063 (N_45063,N_44139,N_44847);
nor U45064 (N_45064,N_44752,N_44226);
or U45065 (N_45065,N_44457,N_44075);
and U45066 (N_45066,N_44822,N_44548);
nand U45067 (N_45067,N_44542,N_44720);
xor U45068 (N_45068,N_44212,N_44043);
and U45069 (N_45069,N_44945,N_44610);
and U45070 (N_45070,N_44855,N_44864);
or U45071 (N_45071,N_44307,N_44251);
and U45072 (N_45072,N_44565,N_44630);
or U45073 (N_45073,N_44863,N_44489);
nor U45074 (N_45074,N_44336,N_44430);
and U45075 (N_45075,N_44913,N_44823);
or U45076 (N_45076,N_44607,N_44120);
and U45077 (N_45077,N_44149,N_44960);
or U45078 (N_45078,N_44731,N_44224);
nor U45079 (N_45079,N_44985,N_44833);
nor U45080 (N_45080,N_44887,N_44150);
nor U45081 (N_45081,N_44324,N_44563);
nand U45082 (N_45082,N_44178,N_44981);
nor U45083 (N_45083,N_44963,N_44956);
nand U45084 (N_45084,N_44366,N_44560);
xnor U45085 (N_45085,N_44136,N_44350);
xor U45086 (N_45086,N_44127,N_44500);
xor U45087 (N_45087,N_44323,N_44287);
nor U45088 (N_45088,N_44313,N_44729);
nand U45089 (N_45089,N_44991,N_44773);
nor U45090 (N_45090,N_44303,N_44562);
xor U45091 (N_45091,N_44784,N_44519);
and U45092 (N_45092,N_44685,N_44705);
xnor U45093 (N_45093,N_44346,N_44029);
or U45094 (N_45094,N_44399,N_44253);
and U45095 (N_45095,N_44827,N_44045);
and U45096 (N_45096,N_44574,N_44471);
nor U45097 (N_45097,N_44347,N_44325);
nor U45098 (N_45098,N_44764,N_44905);
nand U45099 (N_45099,N_44976,N_44578);
nor U45100 (N_45100,N_44206,N_44690);
nor U45101 (N_45101,N_44555,N_44750);
nor U45102 (N_45102,N_44048,N_44143);
nand U45103 (N_45103,N_44357,N_44196);
or U45104 (N_45104,N_44077,N_44038);
or U45105 (N_45105,N_44917,N_44230);
nor U45106 (N_45106,N_44538,N_44369);
nand U45107 (N_45107,N_44549,N_44672);
or U45108 (N_45108,N_44872,N_44481);
xor U45109 (N_45109,N_44689,N_44603);
xnor U45110 (N_45110,N_44939,N_44796);
nand U45111 (N_45111,N_44421,N_44349);
xor U45112 (N_45112,N_44749,N_44765);
nor U45113 (N_45113,N_44436,N_44826);
nand U45114 (N_45114,N_44066,N_44769);
nor U45115 (N_45115,N_44737,N_44658);
nor U45116 (N_45116,N_44219,N_44181);
nand U45117 (N_45117,N_44546,N_44199);
and U45118 (N_45118,N_44113,N_44531);
nand U45119 (N_45119,N_44670,N_44448);
nor U45120 (N_45120,N_44930,N_44257);
xnor U45121 (N_45121,N_44541,N_44259);
nor U45122 (N_45122,N_44180,N_44176);
xor U45123 (N_45123,N_44123,N_44813);
and U45124 (N_45124,N_44965,N_44594);
xnor U45125 (N_45125,N_44002,N_44110);
nor U45126 (N_45126,N_44084,N_44783);
nand U45127 (N_45127,N_44730,N_44843);
nor U45128 (N_45128,N_44001,N_44019);
xnor U45129 (N_45129,N_44861,N_44638);
or U45130 (N_45130,N_44683,N_44393);
or U45131 (N_45131,N_44487,N_44400);
xnor U45132 (N_45132,N_44141,N_44550);
or U45133 (N_45133,N_44645,N_44424);
nand U45134 (N_45134,N_44680,N_44473);
or U45135 (N_45135,N_44153,N_44335);
or U45136 (N_45136,N_44679,N_44007);
nor U45137 (N_45137,N_44995,N_44992);
or U45138 (N_45138,N_44289,N_44572);
or U45139 (N_45139,N_44824,N_44951);
nand U45140 (N_45140,N_44947,N_44915);
xor U45141 (N_45141,N_44604,N_44418);
nand U45142 (N_45142,N_44821,N_44083);
xnor U45143 (N_45143,N_44641,N_44878);
and U45144 (N_45144,N_44390,N_44063);
and U45145 (N_45145,N_44948,N_44233);
xnor U45146 (N_45146,N_44697,N_44733);
or U45147 (N_45147,N_44760,N_44865);
xor U45148 (N_45148,N_44454,N_44944);
and U45149 (N_45149,N_44398,N_44041);
nor U45150 (N_45150,N_44318,N_44381);
nand U45151 (N_45151,N_44086,N_44559);
nand U45152 (N_45152,N_44619,N_44900);
nor U45153 (N_45153,N_44615,N_44354);
xor U45154 (N_45154,N_44691,N_44072);
nor U45155 (N_45155,N_44104,N_44167);
and U45156 (N_45156,N_44392,N_44282);
or U45157 (N_45157,N_44036,N_44606);
xor U45158 (N_45158,N_44870,N_44291);
or U45159 (N_45159,N_44655,N_44345);
nor U45160 (N_45160,N_44717,N_44830);
and U45161 (N_45161,N_44994,N_44522);
and U45162 (N_45162,N_44348,N_44617);
nand U45163 (N_45163,N_44311,N_44746);
and U45164 (N_45164,N_44194,N_44839);
xnor U45165 (N_45165,N_44065,N_44850);
xnor U45166 (N_45166,N_44420,N_44148);
and U45167 (N_45167,N_44152,N_44653);
nand U45168 (N_45168,N_44358,N_44243);
xor U45169 (N_45169,N_44015,N_44906);
nand U45170 (N_45170,N_44020,N_44384);
or U45171 (N_45171,N_44674,N_44359);
nand U45172 (N_45172,N_44988,N_44547);
and U45173 (N_45173,N_44187,N_44698);
or U45174 (N_45174,N_44306,N_44414);
and U45175 (N_45175,N_44647,N_44627);
xor U45176 (N_45176,N_44632,N_44488);
or U45177 (N_45177,N_44232,N_44807);
nand U45178 (N_45178,N_44070,N_44258);
xnor U45179 (N_45179,N_44654,N_44942);
and U45180 (N_45180,N_44774,N_44625);
nand U45181 (N_45181,N_44753,N_44678);
or U45182 (N_45182,N_44344,N_44031);
xnor U45183 (N_45183,N_44809,N_44191);
and U45184 (N_45184,N_44694,N_44221);
nand U45185 (N_45185,N_44050,N_44261);
xor U45186 (N_45186,N_44094,N_44445);
nand U45187 (N_45187,N_44005,N_44405);
xnor U45188 (N_45188,N_44118,N_44047);
nor U45189 (N_45189,N_44567,N_44440);
nor U45190 (N_45190,N_44696,N_44961);
xor U45191 (N_45191,N_44203,N_44021);
nand U45192 (N_45192,N_44812,N_44871);
or U45193 (N_45193,N_44447,N_44977);
and U45194 (N_45194,N_44928,N_44794);
nor U45195 (N_45195,N_44622,N_44513);
or U45196 (N_45196,N_44000,N_44278);
nor U45197 (N_45197,N_44776,N_44927);
nor U45198 (N_45198,N_44537,N_44220);
nand U45199 (N_45199,N_44561,N_44707);
or U45200 (N_45200,N_44726,N_44244);
xnor U45201 (N_45201,N_44789,N_44569);
and U45202 (N_45202,N_44290,N_44030);
xor U45203 (N_45203,N_44171,N_44211);
or U45204 (N_45204,N_44463,N_44093);
nor U45205 (N_45205,N_44551,N_44528);
xor U45206 (N_45206,N_44416,N_44996);
and U45207 (N_45207,N_44106,N_44508);
nor U45208 (N_45208,N_44929,N_44126);
and U45209 (N_45209,N_44492,N_44986);
and U45210 (N_45210,N_44074,N_44444);
nand U45211 (N_45211,N_44060,N_44319);
and U45212 (N_45212,N_44483,N_44946);
nand U45213 (N_45213,N_44890,N_44660);
nor U45214 (N_45214,N_44498,N_44704);
nor U45215 (N_45215,N_44342,N_44975);
or U45216 (N_45216,N_44302,N_44849);
nor U45217 (N_45217,N_44435,N_44974);
and U45218 (N_45218,N_44596,N_44484);
or U45219 (N_45219,N_44536,N_44252);
nor U45220 (N_45220,N_44124,N_44010);
nor U45221 (N_45221,N_44777,N_44734);
and U45222 (N_45222,N_44391,N_44267);
or U45223 (N_45223,N_44166,N_44408);
xor U45224 (N_45224,N_44057,N_44198);
xor U45225 (N_45225,N_44160,N_44702);
xnor U45226 (N_45226,N_44371,N_44853);
and U45227 (N_45227,N_44268,N_44980);
nand U45228 (N_45228,N_44245,N_44477);
and U45229 (N_45229,N_44082,N_44499);
and U45230 (N_45230,N_44936,N_44953);
or U45231 (N_45231,N_44533,N_44634);
and U45232 (N_45232,N_44640,N_44589);
nor U45233 (N_45233,N_44044,N_44575);
or U45234 (N_45234,N_44330,N_44091);
and U45235 (N_45235,N_44101,N_44540);
xnor U45236 (N_45236,N_44506,N_44207);
or U45237 (N_45237,N_44882,N_44503);
or U45238 (N_45238,N_44130,N_44714);
or U45239 (N_45239,N_44739,N_44061);
nand U45240 (N_45240,N_44684,N_44204);
nand U45241 (N_45241,N_44819,N_44626);
xor U45242 (N_45242,N_44406,N_44873);
or U45243 (N_45243,N_44553,N_44254);
and U45244 (N_45244,N_44059,N_44231);
nand U45245 (N_45245,N_44401,N_44249);
nand U45246 (N_45246,N_44363,N_44434);
or U45247 (N_45247,N_44437,N_44394);
nand U45248 (N_45248,N_44073,N_44741);
or U45249 (N_45249,N_44544,N_44411);
xnor U45250 (N_45250,N_44109,N_44079);
and U45251 (N_45251,N_44816,N_44591);
nand U45252 (N_45252,N_44228,N_44703);
or U45253 (N_45253,N_44621,N_44895);
or U45254 (N_45254,N_44999,N_44761);
xor U45255 (N_45255,N_44164,N_44998);
xor U45256 (N_45256,N_44962,N_44080);
or U45257 (N_45257,N_44068,N_44131);
nand U45258 (N_45258,N_44676,N_44334);
nor U45259 (N_45259,N_44642,N_44004);
xnor U45260 (N_45260,N_44601,N_44724);
and U45261 (N_45261,N_44154,N_44983);
nor U45262 (N_45262,N_44427,N_44592);
or U45263 (N_45263,N_44014,N_44779);
xnor U45264 (N_45264,N_44037,N_44718);
nor U45265 (N_45265,N_44085,N_44423);
nor U45266 (N_45266,N_44757,N_44545);
or U45267 (N_45267,N_44343,N_44460);
and U45268 (N_45268,N_44317,N_44543);
xor U45269 (N_45269,N_44791,N_44027);
or U45270 (N_45270,N_44024,N_44117);
xor U45271 (N_45271,N_44926,N_44693);
and U45272 (N_45272,N_44404,N_44766);
nand U45273 (N_45273,N_44524,N_44635);
or U45274 (N_45274,N_44908,N_44429);
nand U45275 (N_45275,N_44184,N_44351);
xor U45276 (N_45276,N_44129,N_44831);
nor U45277 (N_45277,N_44521,N_44145);
nand U45278 (N_45278,N_44571,N_44469);
and U45279 (N_45279,N_44223,N_44611);
nor U45280 (N_45280,N_44566,N_44389);
nor U45281 (N_45281,N_44209,N_44175);
or U45282 (N_45282,N_44284,N_44441);
and U45283 (N_45283,N_44896,N_44234);
and U45284 (N_45284,N_44785,N_44163);
or U45285 (N_45285,N_44138,N_44316);
and U45286 (N_45286,N_44375,N_44032);
and U45287 (N_45287,N_44439,N_44280);
nand U45288 (N_45288,N_44511,N_44098);
and U45289 (N_45289,N_44173,N_44517);
or U45290 (N_45290,N_44121,N_44377);
nand U45291 (N_45291,N_44860,N_44312);
and U45292 (N_45292,N_44266,N_44395);
nand U45293 (N_45293,N_44025,N_44431);
nand U45294 (N_45294,N_44409,N_44248);
nand U45295 (N_45295,N_44745,N_44593);
or U45296 (N_45296,N_44598,N_44475);
or U45297 (N_45297,N_44088,N_44662);
xnor U45298 (N_45298,N_44095,N_44918);
nand U45299 (N_45299,N_44142,N_44526);
xor U45300 (N_45300,N_44069,N_44894);
nor U45301 (N_45301,N_44588,N_44305);
and U45302 (N_45302,N_44195,N_44505);
nand U45303 (N_45303,N_44419,N_44668);
nor U45304 (N_45304,N_44467,N_44602);
xnor U45305 (N_45305,N_44744,N_44225);
xnor U45306 (N_45306,N_44552,N_44197);
or U45307 (N_45307,N_44509,N_44331);
nor U45308 (N_45308,N_44337,N_44957);
nand U45309 (N_45309,N_44775,N_44581);
or U45310 (N_45310,N_44842,N_44321);
and U45311 (N_45311,N_44156,N_44486);
nand U45312 (N_45312,N_44558,N_44190);
and U45313 (N_45313,N_44193,N_44332);
or U45314 (N_45314,N_44682,N_44504);
nand U45315 (N_45315,N_44925,N_44997);
or U45316 (N_45316,N_44017,N_44675);
xor U45317 (N_45317,N_44049,N_44815);
nor U45318 (N_45318,N_44786,N_44608);
or U45319 (N_45319,N_44643,N_44297);
xnor U45320 (N_45320,N_44046,N_44264);
nand U45321 (N_45321,N_44051,N_44215);
nand U45322 (N_45322,N_44449,N_44652);
nor U45323 (N_45323,N_44612,N_44650);
or U45324 (N_45324,N_44170,N_44210);
and U45325 (N_45325,N_44200,N_44780);
or U45326 (N_45326,N_44035,N_44656);
nand U45327 (N_45327,N_44422,N_44263);
nor U45328 (N_45328,N_44055,N_44214);
nand U45329 (N_45329,N_44361,N_44742);
or U45330 (N_45330,N_44797,N_44071);
xor U45331 (N_45331,N_44686,N_44743);
xor U45332 (N_45332,N_44554,N_44053);
and U45333 (N_45333,N_44159,N_44667);
nand U45334 (N_45334,N_44100,N_44382);
and U45335 (N_45335,N_44751,N_44959);
or U45336 (N_45336,N_44494,N_44183);
and U45337 (N_45337,N_44879,N_44782);
nor U45338 (N_45338,N_44125,N_44360);
and U45339 (N_45339,N_44587,N_44497);
nor U45340 (N_45340,N_44056,N_44112);
and U45341 (N_45341,N_44296,N_44396);
xor U45342 (N_45342,N_44456,N_44003);
xor U45343 (N_45343,N_44132,N_44695);
nor U45344 (N_45344,N_44426,N_44671);
nor U45345 (N_45345,N_44458,N_44579);
xor U45346 (N_45346,N_44480,N_44496);
nand U45347 (N_45347,N_44692,N_44365);
nand U45348 (N_45348,N_44620,N_44735);
nor U45349 (N_45349,N_44265,N_44340);
or U45350 (N_45350,N_44790,N_44535);
nand U45351 (N_45351,N_44699,N_44092);
xnor U45352 (N_45352,N_44920,N_44557);
and U45353 (N_45353,N_44754,N_44111);
and U45354 (N_45354,N_44978,N_44459);
nand U45355 (N_45355,N_44452,N_44681);
or U45356 (N_45356,N_44885,N_44174);
xnor U45357 (N_45357,N_44912,N_44628);
nand U45358 (N_45358,N_44308,N_44339);
xor U45359 (N_45359,N_44874,N_44514);
or U45360 (N_45360,N_44875,N_44989);
nand U45361 (N_45361,N_44646,N_44820);
or U45362 (N_45362,N_44848,N_44599);
or U45363 (N_45363,N_44446,N_44740);
nand U45364 (N_45364,N_44269,N_44428);
xnor U45365 (N_45365,N_44468,N_44107);
or U45366 (N_45366,N_44096,N_44018);
and U45367 (N_45367,N_44116,N_44993);
nor U45368 (N_45368,N_44134,N_44179);
and U45369 (N_45369,N_44241,N_44491);
and U45370 (N_45370,N_44728,N_44476);
or U45371 (N_45371,N_44664,N_44834);
xnor U45372 (N_45372,N_44597,N_44165);
nor U45373 (N_45373,N_44756,N_44710);
or U45374 (N_45374,N_44810,N_44034);
and U45375 (N_45375,N_44866,N_44262);
nor U45376 (N_45376,N_44964,N_44378);
and U45377 (N_45377,N_44955,N_44146);
or U45378 (N_45378,N_44943,N_44250);
nand U45379 (N_45379,N_44386,N_44285);
nand U45380 (N_45380,N_44712,N_44868);
or U45381 (N_45381,N_44931,N_44793);
or U45382 (N_45382,N_44087,N_44022);
or U45383 (N_45383,N_44723,N_44613);
xnor U45384 (N_45384,N_44438,N_44623);
nand U45385 (N_45385,N_44510,N_44817);
nor U45386 (N_45386,N_44938,N_44103);
nand U45387 (N_45387,N_44949,N_44276);
nor U45388 (N_45388,N_44825,N_44937);
or U45389 (N_45389,N_44876,N_44239);
and U45390 (N_45390,N_44984,N_44639);
nor U45391 (N_45391,N_44954,N_44356);
xor U45392 (N_45392,N_44144,N_44013);
nor U45393 (N_45393,N_44708,N_44950);
and U45394 (N_45394,N_44859,N_44889);
or U45395 (N_45395,N_44277,N_44255);
and U45396 (N_45396,N_44852,N_44648);
nor U45397 (N_45397,N_44614,N_44759);
or U45398 (N_45398,N_44837,N_44539);
nor U45399 (N_45399,N_44155,N_44413);
and U45400 (N_45400,N_44952,N_44886);
or U45401 (N_45401,N_44767,N_44624);
nand U45402 (N_45402,N_44715,N_44832);
nor U45403 (N_45403,N_44840,N_44605);
nand U45404 (N_45404,N_44105,N_44727);
or U45405 (N_45405,N_44236,N_44062);
and U45406 (N_45406,N_44738,N_44370);
xnor U45407 (N_45407,N_44770,N_44403);
and U45408 (N_45408,N_44914,N_44798);
nand U45409 (N_45409,N_44301,N_44485);
and U45410 (N_45410,N_44502,N_44294);
xor U45411 (N_45411,N_44971,N_44169);
or U45412 (N_45412,N_44629,N_44595);
or U45413 (N_45413,N_44147,N_44706);
xnor U45414 (N_45414,N_44933,N_44490);
nor U45415 (N_45415,N_44932,N_44911);
xor U45416 (N_45416,N_44202,N_44238);
xnor U45417 (N_45417,N_44465,N_44133);
and U45418 (N_45418,N_44616,N_44379);
xnor U45419 (N_45419,N_44412,N_44310);
or U45420 (N_45420,N_44924,N_44577);
or U45421 (N_45421,N_44732,N_44763);
and U45422 (N_45422,N_44585,N_44140);
and U45423 (N_45423,N_44828,N_44516);
xnor U45424 (N_45424,N_44636,N_44011);
nand U45425 (N_45425,N_44415,N_44122);
or U45426 (N_45426,N_44341,N_44161);
or U45427 (N_45427,N_44829,N_44811);
nand U45428 (N_45428,N_44529,N_44372);
nor U45429 (N_45429,N_44182,N_44067);
xor U45430 (N_45430,N_44584,N_44353);
nand U45431 (N_45431,N_44474,N_44097);
nor U45432 (N_45432,N_44185,N_44376);
nand U45433 (N_45433,N_44982,N_44901);
nand U45434 (N_45434,N_44322,N_44618);
nand U45435 (N_45435,N_44217,N_44237);
and U45436 (N_45436,N_44218,N_44451);
and U45437 (N_45437,N_44158,N_44857);
and U45438 (N_45438,N_44102,N_44270);
nor U45439 (N_45439,N_44530,N_44657);
and U45440 (N_45440,N_44192,N_44064);
xor U45441 (N_45441,N_44283,N_44838);
and U45442 (N_45442,N_44364,N_44033);
or U45443 (N_45443,N_44921,N_44177);
xor U45444 (N_45444,N_44162,N_44407);
and U45445 (N_45445,N_44877,N_44922);
and U45446 (N_45446,N_44425,N_44309);
or U45447 (N_45447,N_44028,N_44189);
or U45448 (N_45448,N_44799,N_44026);
and U45449 (N_45449,N_44374,N_44081);
xor U45450 (N_45450,N_44293,N_44907);
xor U45451 (N_45451,N_44367,N_44208);
or U45452 (N_45452,N_44520,N_44899);
nand U45453 (N_45453,N_44804,N_44570);
xor U45454 (N_45454,N_44478,N_44470);
or U45455 (N_45455,N_44410,N_44298);
and U45456 (N_45456,N_44532,N_44719);
or U45457 (N_45457,N_44910,N_44903);
nor U45458 (N_45458,N_44501,N_44279);
nor U45459 (N_45459,N_44137,N_44755);
or U45460 (N_45460,N_44433,N_44205);
xor U45461 (N_45461,N_44288,N_44792);
xor U45462 (N_45462,N_44846,N_44242);
nor U45463 (N_45463,N_44583,N_44515);
xor U45464 (N_45464,N_44748,N_44969);
and U45465 (N_45465,N_44119,N_44525);
nand U45466 (N_45466,N_44328,N_44383);
and U45467 (N_45467,N_44078,N_44009);
xor U45468 (N_45468,N_44380,N_44891);
xnor U45469 (N_45469,N_44990,N_44881);
nand U45470 (N_45470,N_44688,N_44987);
and U45471 (N_45471,N_44304,N_44466);
and U45472 (N_45472,N_44701,N_44329);
and U45473 (N_45473,N_44758,N_44644);
xnor U45474 (N_45474,N_44534,N_44788);
and U45475 (N_45475,N_44795,N_44649);
nand U45476 (N_45476,N_44919,N_44818);
or U45477 (N_45477,N_44883,N_44368);
nand U45478 (N_45478,N_44972,N_44893);
nand U45479 (N_45479,N_44090,N_44709);
and U45480 (N_45480,N_44482,N_44590);
and U45481 (N_45481,N_44803,N_44042);
xor U45482 (N_45482,N_44609,N_44006);
nand U45483 (N_45483,N_44527,N_44631);
nor U45484 (N_45484,N_44806,N_44898);
nand U45485 (N_45485,N_44417,N_44315);
or U45486 (N_45486,N_44787,N_44663);
nand U45487 (N_45487,N_44089,N_44455);
or U45488 (N_45488,N_44135,N_44902);
and U45489 (N_45489,N_44240,N_44665);
or U45490 (N_45490,N_44841,N_44747);
nand U45491 (N_45491,N_44213,N_44052);
and U45492 (N_45492,N_44450,N_44721);
and U45493 (N_45493,N_44805,N_44128);
or U45494 (N_45494,N_44292,N_44651);
xnor U45495 (N_45495,N_44108,N_44762);
or U45496 (N_45496,N_44941,N_44472);
or U45497 (N_45497,N_44216,N_44556);
xnor U45498 (N_45498,N_44300,N_44355);
nor U45499 (N_45499,N_44295,N_44464);
nand U45500 (N_45500,N_44874,N_44376);
or U45501 (N_45501,N_44459,N_44063);
or U45502 (N_45502,N_44680,N_44561);
or U45503 (N_45503,N_44287,N_44780);
and U45504 (N_45504,N_44412,N_44797);
and U45505 (N_45505,N_44698,N_44538);
xnor U45506 (N_45506,N_44726,N_44874);
xor U45507 (N_45507,N_44585,N_44926);
xnor U45508 (N_45508,N_44941,N_44175);
nor U45509 (N_45509,N_44906,N_44666);
xor U45510 (N_45510,N_44894,N_44484);
nand U45511 (N_45511,N_44678,N_44870);
or U45512 (N_45512,N_44135,N_44530);
and U45513 (N_45513,N_44643,N_44931);
or U45514 (N_45514,N_44037,N_44465);
nand U45515 (N_45515,N_44312,N_44391);
xnor U45516 (N_45516,N_44196,N_44360);
or U45517 (N_45517,N_44516,N_44280);
nand U45518 (N_45518,N_44475,N_44366);
xnor U45519 (N_45519,N_44969,N_44340);
xor U45520 (N_45520,N_44009,N_44960);
nor U45521 (N_45521,N_44608,N_44841);
nor U45522 (N_45522,N_44445,N_44679);
nand U45523 (N_45523,N_44011,N_44288);
and U45524 (N_45524,N_44434,N_44131);
and U45525 (N_45525,N_44488,N_44566);
nand U45526 (N_45526,N_44105,N_44220);
nor U45527 (N_45527,N_44003,N_44226);
xnor U45528 (N_45528,N_44604,N_44966);
nand U45529 (N_45529,N_44059,N_44485);
xnor U45530 (N_45530,N_44199,N_44216);
xor U45531 (N_45531,N_44459,N_44327);
and U45532 (N_45532,N_44730,N_44410);
or U45533 (N_45533,N_44220,N_44607);
and U45534 (N_45534,N_44129,N_44304);
or U45535 (N_45535,N_44848,N_44157);
or U45536 (N_45536,N_44237,N_44677);
nand U45537 (N_45537,N_44724,N_44595);
nand U45538 (N_45538,N_44249,N_44244);
nand U45539 (N_45539,N_44723,N_44322);
or U45540 (N_45540,N_44762,N_44170);
nor U45541 (N_45541,N_44999,N_44062);
or U45542 (N_45542,N_44228,N_44863);
xnor U45543 (N_45543,N_44795,N_44574);
or U45544 (N_45544,N_44154,N_44807);
nor U45545 (N_45545,N_44061,N_44858);
and U45546 (N_45546,N_44288,N_44571);
or U45547 (N_45547,N_44979,N_44384);
xnor U45548 (N_45548,N_44066,N_44724);
nand U45549 (N_45549,N_44445,N_44593);
or U45550 (N_45550,N_44788,N_44691);
or U45551 (N_45551,N_44793,N_44337);
xor U45552 (N_45552,N_44689,N_44197);
and U45553 (N_45553,N_44978,N_44531);
nand U45554 (N_45554,N_44813,N_44930);
or U45555 (N_45555,N_44424,N_44127);
nand U45556 (N_45556,N_44554,N_44119);
nor U45557 (N_45557,N_44683,N_44082);
and U45558 (N_45558,N_44509,N_44450);
and U45559 (N_45559,N_44693,N_44044);
or U45560 (N_45560,N_44723,N_44670);
and U45561 (N_45561,N_44243,N_44757);
or U45562 (N_45562,N_44758,N_44772);
nand U45563 (N_45563,N_44705,N_44542);
nand U45564 (N_45564,N_44075,N_44478);
nand U45565 (N_45565,N_44493,N_44793);
and U45566 (N_45566,N_44232,N_44041);
and U45567 (N_45567,N_44305,N_44666);
nand U45568 (N_45568,N_44254,N_44060);
nor U45569 (N_45569,N_44518,N_44468);
nand U45570 (N_45570,N_44041,N_44401);
and U45571 (N_45571,N_44535,N_44308);
or U45572 (N_45572,N_44689,N_44568);
xor U45573 (N_45573,N_44077,N_44189);
nand U45574 (N_45574,N_44915,N_44066);
nand U45575 (N_45575,N_44911,N_44252);
nand U45576 (N_45576,N_44410,N_44920);
nor U45577 (N_45577,N_44805,N_44578);
nand U45578 (N_45578,N_44287,N_44892);
nor U45579 (N_45579,N_44711,N_44543);
nor U45580 (N_45580,N_44257,N_44836);
xor U45581 (N_45581,N_44850,N_44769);
nor U45582 (N_45582,N_44475,N_44122);
xnor U45583 (N_45583,N_44910,N_44449);
and U45584 (N_45584,N_44292,N_44947);
or U45585 (N_45585,N_44505,N_44718);
xor U45586 (N_45586,N_44399,N_44034);
and U45587 (N_45587,N_44523,N_44014);
nor U45588 (N_45588,N_44799,N_44416);
nand U45589 (N_45589,N_44867,N_44202);
nand U45590 (N_45590,N_44085,N_44626);
nand U45591 (N_45591,N_44434,N_44204);
or U45592 (N_45592,N_44019,N_44795);
xnor U45593 (N_45593,N_44495,N_44936);
or U45594 (N_45594,N_44887,N_44099);
xor U45595 (N_45595,N_44757,N_44028);
and U45596 (N_45596,N_44493,N_44473);
nand U45597 (N_45597,N_44135,N_44881);
and U45598 (N_45598,N_44585,N_44793);
nand U45599 (N_45599,N_44959,N_44361);
or U45600 (N_45600,N_44195,N_44855);
nor U45601 (N_45601,N_44012,N_44726);
or U45602 (N_45602,N_44488,N_44698);
or U45603 (N_45603,N_44981,N_44983);
nor U45604 (N_45604,N_44804,N_44506);
nor U45605 (N_45605,N_44942,N_44961);
xnor U45606 (N_45606,N_44007,N_44686);
nor U45607 (N_45607,N_44433,N_44985);
and U45608 (N_45608,N_44844,N_44678);
nor U45609 (N_45609,N_44484,N_44336);
or U45610 (N_45610,N_44910,N_44644);
and U45611 (N_45611,N_44094,N_44680);
and U45612 (N_45612,N_44609,N_44486);
xnor U45613 (N_45613,N_44683,N_44794);
nand U45614 (N_45614,N_44515,N_44383);
xnor U45615 (N_45615,N_44847,N_44556);
nor U45616 (N_45616,N_44431,N_44276);
nor U45617 (N_45617,N_44166,N_44768);
xnor U45618 (N_45618,N_44822,N_44273);
nor U45619 (N_45619,N_44650,N_44585);
nor U45620 (N_45620,N_44576,N_44988);
xnor U45621 (N_45621,N_44014,N_44471);
nor U45622 (N_45622,N_44633,N_44995);
nor U45623 (N_45623,N_44916,N_44390);
nor U45624 (N_45624,N_44151,N_44562);
nor U45625 (N_45625,N_44527,N_44908);
and U45626 (N_45626,N_44951,N_44132);
xor U45627 (N_45627,N_44565,N_44708);
or U45628 (N_45628,N_44357,N_44945);
xor U45629 (N_45629,N_44054,N_44194);
nand U45630 (N_45630,N_44699,N_44563);
and U45631 (N_45631,N_44417,N_44330);
and U45632 (N_45632,N_44534,N_44509);
and U45633 (N_45633,N_44232,N_44751);
or U45634 (N_45634,N_44900,N_44676);
xnor U45635 (N_45635,N_44413,N_44174);
nand U45636 (N_45636,N_44241,N_44703);
or U45637 (N_45637,N_44382,N_44515);
nand U45638 (N_45638,N_44321,N_44447);
or U45639 (N_45639,N_44762,N_44014);
xnor U45640 (N_45640,N_44273,N_44261);
nor U45641 (N_45641,N_44028,N_44393);
nor U45642 (N_45642,N_44167,N_44805);
xor U45643 (N_45643,N_44548,N_44805);
and U45644 (N_45644,N_44134,N_44961);
xnor U45645 (N_45645,N_44578,N_44726);
or U45646 (N_45646,N_44797,N_44986);
nand U45647 (N_45647,N_44870,N_44671);
or U45648 (N_45648,N_44622,N_44132);
or U45649 (N_45649,N_44261,N_44200);
xor U45650 (N_45650,N_44523,N_44695);
xor U45651 (N_45651,N_44338,N_44428);
nand U45652 (N_45652,N_44956,N_44526);
or U45653 (N_45653,N_44334,N_44294);
nor U45654 (N_45654,N_44186,N_44218);
or U45655 (N_45655,N_44261,N_44745);
nor U45656 (N_45656,N_44546,N_44301);
nand U45657 (N_45657,N_44318,N_44426);
nor U45658 (N_45658,N_44889,N_44562);
and U45659 (N_45659,N_44258,N_44720);
nor U45660 (N_45660,N_44551,N_44320);
nor U45661 (N_45661,N_44261,N_44090);
xnor U45662 (N_45662,N_44658,N_44214);
or U45663 (N_45663,N_44831,N_44326);
nand U45664 (N_45664,N_44639,N_44241);
nor U45665 (N_45665,N_44847,N_44800);
or U45666 (N_45666,N_44910,N_44169);
and U45667 (N_45667,N_44331,N_44588);
xor U45668 (N_45668,N_44558,N_44612);
or U45669 (N_45669,N_44814,N_44784);
nand U45670 (N_45670,N_44303,N_44673);
or U45671 (N_45671,N_44110,N_44214);
nor U45672 (N_45672,N_44213,N_44804);
nor U45673 (N_45673,N_44966,N_44547);
xnor U45674 (N_45674,N_44177,N_44060);
xnor U45675 (N_45675,N_44632,N_44054);
xnor U45676 (N_45676,N_44354,N_44757);
and U45677 (N_45677,N_44503,N_44372);
xor U45678 (N_45678,N_44125,N_44513);
nor U45679 (N_45679,N_44484,N_44488);
nor U45680 (N_45680,N_44502,N_44147);
xnor U45681 (N_45681,N_44660,N_44481);
and U45682 (N_45682,N_44812,N_44043);
or U45683 (N_45683,N_44049,N_44501);
and U45684 (N_45684,N_44522,N_44225);
nand U45685 (N_45685,N_44792,N_44581);
xor U45686 (N_45686,N_44663,N_44664);
xor U45687 (N_45687,N_44805,N_44754);
or U45688 (N_45688,N_44391,N_44080);
and U45689 (N_45689,N_44949,N_44482);
xor U45690 (N_45690,N_44741,N_44671);
or U45691 (N_45691,N_44794,N_44029);
nand U45692 (N_45692,N_44931,N_44713);
nor U45693 (N_45693,N_44218,N_44822);
and U45694 (N_45694,N_44729,N_44567);
nor U45695 (N_45695,N_44097,N_44398);
and U45696 (N_45696,N_44374,N_44507);
nor U45697 (N_45697,N_44654,N_44058);
nor U45698 (N_45698,N_44509,N_44786);
and U45699 (N_45699,N_44678,N_44049);
and U45700 (N_45700,N_44669,N_44648);
xnor U45701 (N_45701,N_44642,N_44418);
or U45702 (N_45702,N_44273,N_44657);
xnor U45703 (N_45703,N_44626,N_44019);
or U45704 (N_45704,N_44868,N_44090);
xor U45705 (N_45705,N_44636,N_44853);
nand U45706 (N_45706,N_44490,N_44010);
nor U45707 (N_45707,N_44291,N_44203);
or U45708 (N_45708,N_44409,N_44541);
nand U45709 (N_45709,N_44229,N_44826);
nor U45710 (N_45710,N_44102,N_44770);
and U45711 (N_45711,N_44425,N_44541);
and U45712 (N_45712,N_44363,N_44973);
nand U45713 (N_45713,N_44079,N_44475);
nand U45714 (N_45714,N_44887,N_44946);
xnor U45715 (N_45715,N_44797,N_44008);
nand U45716 (N_45716,N_44567,N_44115);
nor U45717 (N_45717,N_44430,N_44918);
and U45718 (N_45718,N_44465,N_44374);
nor U45719 (N_45719,N_44913,N_44429);
or U45720 (N_45720,N_44544,N_44817);
nand U45721 (N_45721,N_44577,N_44410);
nor U45722 (N_45722,N_44977,N_44311);
and U45723 (N_45723,N_44129,N_44458);
nor U45724 (N_45724,N_44160,N_44237);
nor U45725 (N_45725,N_44154,N_44259);
or U45726 (N_45726,N_44395,N_44721);
nor U45727 (N_45727,N_44454,N_44272);
nand U45728 (N_45728,N_44981,N_44215);
and U45729 (N_45729,N_44523,N_44030);
nor U45730 (N_45730,N_44942,N_44025);
xor U45731 (N_45731,N_44993,N_44892);
and U45732 (N_45732,N_44731,N_44923);
xnor U45733 (N_45733,N_44884,N_44153);
nor U45734 (N_45734,N_44812,N_44553);
and U45735 (N_45735,N_44756,N_44937);
or U45736 (N_45736,N_44227,N_44301);
nand U45737 (N_45737,N_44655,N_44375);
or U45738 (N_45738,N_44758,N_44318);
xnor U45739 (N_45739,N_44443,N_44425);
xnor U45740 (N_45740,N_44281,N_44974);
nor U45741 (N_45741,N_44042,N_44510);
xnor U45742 (N_45742,N_44659,N_44812);
nor U45743 (N_45743,N_44102,N_44493);
nor U45744 (N_45744,N_44354,N_44210);
nand U45745 (N_45745,N_44245,N_44406);
xnor U45746 (N_45746,N_44330,N_44277);
or U45747 (N_45747,N_44885,N_44425);
or U45748 (N_45748,N_44511,N_44410);
nand U45749 (N_45749,N_44738,N_44215);
nor U45750 (N_45750,N_44066,N_44616);
or U45751 (N_45751,N_44657,N_44962);
xor U45752 (N_45752,N_44022,N_44564);
and U45753 (N_45753,N_44630,N_44837);
nor U45754 (N_45754,N_44886,N_44035);
nand U45755 (N_45755,N_44340,N_44841);
and U45756 (N_45756,N_44462,N_44154);
and U45757 (N_45757,N_44303,N_44931);
nand U45758 (N_45758,N_44054,N_44497);
nor U45759 (N_45759,N_44033,N_44346);
nand U45760 (N_45760,N_44874,N_44290);
nand U45761 (N_45761,N_44698,N_44956);
nand U45762 (N_45762,N_44044,N_44344);
xnor U45763 (N_45763,N_44857,N_44109);
xor U45764 (N_45764,N_44277,N_44398);
nand U45765 (N_45765,N_44380,N_44849);
or U45766 (N_45766,N_44786,N_44291);
nand U45767 (N_45767,N_44855,N_44947);
or U45768 (N_45768,N_44036,N_44664);
and U45769 (N_45769,N_44241,N_44566);
or U45770 (N_45770,N_44783,N_44899);
and U45771 (N_45771,N_44483,N_44078);
nand U45772 (N_45772,N_44054,N_44181);
or U45773 (N_45773,N_44899,N_44554);
or U45774 (N_45774,N_44564,N_44557);
or U45775 (N_45775,N_44615,N_44845);
and U45776 (N_45776,N_44218,N_44463);
and U45777 (N_45777,N_44238,N_44413);
nand U45778 (N_45778,N_44860,N_44206);
or U45779 (N_45779,N_44049,N_44936);
nand U45780 (N_45780,N_44878,N_44154);
xor U45781 (N_45781,N_44002,N_44924);
or U45782 (N_45782,N_44703,N_44355);
nor U45783 (N_45783,N_44160,N_44919);
nor U45784 (N_45784,N_44093,N_44516);
or U45785 (N_45785,N_44250,N_44155);
nor U45786 (N_45786,N_44254,N_44712);
xnor U45787 (N_45787,N_44118,N_44416);
xnor U45788 (N_45788,N_44466,N_44769);
nand U45789 (N_45789,N_44534,N_44956);
and U45790 (N_45790,N_44913,N_44994);
nand U45791 (N_45791,N_44343,N_44878);
nand U45792 (N_45792,N_44392,N_44718);
and U45793 (N_45793,N_44223,N_44497);
and U45794 (N_45794,N_44659,N_44896);
nand U45795 (N_45795,N_44203,N_44257);
nand U45796 (N_45796,N_44027,N_44596);
nand U45797 (N_45797,N_44156,N_44424);
xnor U45798 (N_45798,N_44205,N_44434);
nand U45799 (N_45799,N_44874,N_44011);
or U45800 (N_45800,N_44812,N_44837);
and U45801 (N_45801,N_44843,N_44823);
and U45802 (N_45802,N_44658,N_44536);
and U45803 (N_45803,N_44023,N_44622);
or U45804 (N_45804,N_44654,N_44090);
nor U45805 (N_45805,N_44947,N_44276);
and U45806 (N_45806,N_44646,N_44697);
or U45807 (N_45807,N_44672,N_44608);
and U45808 (N_45808,N_44104,N_44585);
and U45809 (N_45809,N_44262,N_44839);
or U45810 (N_45810,N_44531,N_44396);
nand U45811 (N_45811,N_44141,N_44799);
and U45812 (N_45812,N_44330,N_44121);
nor U45813 (N_45813,N_44948,N_44607);
nand U45814 (N_45814,N_44443,N_44705);
nor U45815 (N_45815,N_44572,N_44969);
xor U45816 (N_45816,N_44395,N_44651);
nor U45817 (N_45817,N_44927,N_44946);
and U45818 (N_45818,N_44435,N_44351);
xnor U45819 (N_45819,N_44933,N_44890);
nand U45820 (N_45820,N_44130,N_44809);
and U45821 (N_45821,N_44985,N_44580);
or U45822 (N_45822,N_44235,N_44482);
or U45823 (N_45823,N_44842,N_44229);
xnor U45824 (N_45824,N_44000,N_44471);
nor U45825 (N_45825,N_44071,N_44703);
xor U45826 (N_45826,N_44774,N_44991);
and U45827 (N_45827,N_44758,N_44297);
or U45828 (N_45828,N_44909,N_44525);
or U45829 (N_45829,N_44584,N_44198);
xor U45830 (N_45830,N_44110,N_44358);
nor U45831 (N_45831,N_44557,N_44630);
nor U45832 (N_45832,N_44252,N_44896);
and U45833 (N_45833,N_44408,N_44109);
or U45834 (N_45834,N_44925,N_44626);
nand U45835 (N_45835,N_44484,N_44578);
nor U45836 (N_45836,N_44786,N_44700);
or U45837 (N_45837,N_44681,N_44951);
or U45838 (N_45838,N_44767,N_44196);
nand U45839 (N_45839,N_44059,N_44032);
xnor U45840 (N_45840,N_44884,N_44200);
nor U45841 (N_45841,N_44434,N_44387);
xor U45842 (N_45842,N_44971,N_44590);
nor U45843 (N_45843,N_44236,N_44245);
nor U45844 (N_45844,N_44670,N_44278);
xnor U45845 (N_45845,N_44981,N_44732);
or U45846 (N_45846,N_44897,N_44132);
nand U45847 (N_45847,N_44032,N_44486);
and U45848 (N_45848,N_44456,N_44715);
or U45849 (N_45849,N_44365,N_44174);
and U45850 (N_45850,N_44703,N_44124);
and U45851 (N_45851,N_44242,N_44392);
nand U45852 (N_45852,N_44080,N_44144);
or U45853 (N_45853,N_44237,N_44813);
xnor U45854 (N_45854,N_44862,N_44063);
or U45855 (N_45855,N_44554,N_44537);
nand U45856 (N_45856,N_44391,N_44605);
nor U45857 (N_45857,N_44715,N_44554);
or U45858 (N_45858,N_44801,N_44045);
and U45859 (N_45859,N_44987,N_44855);
xor U45860 (N_45860,N_44674,N_44598);
xor U45861 (N_45861,N_44556,N_44397);
nor U45862 (N_45862,N_44959,N_44894);
xnor U45863 (N_45863,N_44284,N_44800);
nand U45864 (N_45864,N_44042,N_44861);
and U45865 (N_45865,N_44417,N_44137);
nand U45866 (N_45866,N_44399,N_44423);
nor U45867 (N_45867,N_44386,N_44894);
or U45868 (N_45868,N_44857,N_44685);
or U45869 (N_45869,N_44449,N_44867);
xor U45870 (N_45870,N_44624,N_44745);
and U45871 (N_45871,N_44882,N_44226);
or U45872 (N_45872,N_44602,N_44769);
nor U45873 (N_45873,N_44013,N_44620);
or U45874 (N_45874,N_44455,N_44181);
or U45875 (N_45875,N_44353,N_44211);
or U45876 (N_45876,N_44754,N_44389);
and U45877 (N_45877,N_44845,N_44130);
xnor U45878 (N_45878,N_44687,N_44943);
and U45879 (N_45879,N_44625,N_44996);
nor U45880 (N_45880,N_44521,N_44380);
nand U45881 (N_45881,N_44139,N_44387);
nand U45882 (N_45882,N_44341,N_44654);
and U45883 (N_45883,N_44300,N_44180);
nor U45884 (N_45884,N_44679,N_44859);
or U45885 (N_45885,N_44097,N_44863);
nor U45886 (N_45886,N_44396,N_44076);
nand U45887 (N_45887,N_44145,N_44924);
xor U45888 (N_45888,N_44791,N_44679);
nand U45889 (N_45889,N_44668,N_44264);
and U45890 (N_45890,N_44219,N_44210);
nor U45891 (N_45891,N_44328,N_44300);
and U45892 (N_45892,N_44875,N_44388);
nand U45893 (N_45893,N_44613,N_44911);
or U45894 (N_45894,N_44205,N_44533);
nand U45895 (N_45895,N_44807,N_44936);
and U45896 (N_45896,N_44241,N_44494);
xor U45897 (N_45897,N_44572,N_44551);
and U45898 (N_45898,N_44425,N_44762);
xnor U45899 (N_45899,N_44640,N_44043);
and U45900 (N_45900,N_44623,N_44340);
nor U45901 (N_45901,N_44308,N_44893);
nand U45902 (N_45902,N_44188,N_44108);
and U45903 (N_45903,N_44246,N_44234);
and U45904 (N_45904,N_44242,N_44525);
nor U45905 (N_45905,N_44128,N_44286);
or U45906 (N_45906,N_44240,N_44189);
nor U45907 (N_45907,N_44766,N_44064);
and U45908 (N_45908,N_44589,N_44026);
and U45909 (N_45909,N_44779,N_44132);
nand U45910 (N_45910,N_44776,N_44579);
nor U45911 (N_45911,N_44302,N_44759);
and U45912 (N_45912,N_44178,N_44797);
xor U45913 (N_45913,N_44313,N_44509);
xor U45914 (N_45914,N_44961,N_44026);
or U45915 (N_45915,N_44653,N_44311);
or U45916 (N_45916,N_44798,N_44036);
xor U45917 (N_45917,N_44729,N_44190);
nand U45918 (N_45918,N_44184,N_44583);
xnor U45919 (N_45919,N_44166,N_44967);
nor U45920 (N_45920,N_44776,N_44742);
and U45921 (N_45921,N_44715,N_44698);
nand U45922 (N_45922,N_44396,N_44460);
and U45923 (N_45923,N_44505,N_44298);
xor U45924 (N_45924,N_44916,N_44994);
or U45925 (N_45925,N_44489,N_44823);
or U45926 (N_45926,N_44451,N_44879);
or U45927 (N_45927,N_44609,N_44564);
xor U45928 (N_45928,N_44918,N_44519);
and U45929 (N_45929,N_44625,N_44051);
xor U45930 (N_45930,N_44784,N_44021);
xor U45931 (N_45931,N_44509,N_44608);
and U45932 (N_45932,N_44347,N_44008);
xnor U45933 (N_45933,N_44978,N_44327);
xor U45934 (N_45934,N_44924,N_44540);
or U45935 (N_45935,N_44370,N_44761);
xnor U45936 (N_45936,N_44831,N_44292);
or U45937 (N_45937,N_44319,N_44226);
nand U45938 (N_45938,N_44231,N_44633);
nand U45939 (N_45939,N_44918,N_44062);
or U45940 (N_45940,N_44062,N_44523);
or U45941 (N_45941,N_44338,N_44889);
or U45942 (N_45942,N_44882,N_44020);
or U45943 (N_45943,N_44060,N_44173);
and U45944 (N_45944,N_44484,N_44592);
and U45945 (N_45945,N_44490,N_44556);
xnor U45946 (N_45946,N_44945,N_44073);
and U45947 (N_45947,N_44380,N_44921);
or U45948 (N_45948,N_44489,N_44267);
nor U45949 (N_45949,N_44236,N_44582);
or U45950 (N_45950,N_44305,N_44076);
or U45951 (N_45951,N_44721,N_44499);
xor U45952 (N_45952,N_44547,N_44510);
and U45953 (N_45953,N_44149,N_44729);
nand U45954 (N_45954,N_44637,N_44510);
and U45955 (N_45955,N_44778,N_44941);
nand U45956 (N_45956,N_44133,N_44990);
nand U45957 (N_45957,N_44395,N_44303);
and U45958 (N_45958,N_44973,N_44795);
nand U45959 (N_45959,N_44023,N_44772);
and U45960 (N_45960,N_44776,N_44267);
and U45961 (N_45961,N_44217,N_44858);
and U45962 (N_45962,N_44621,N_44469);
and U45963 (N_45963,N_44693,N_44649);
or U45964 (N_45964,N_44571,N_44330);
or U45965 (N_45965,N_44515,N_44715);
or U45966 (N_45966,N_44994,N_44241);
or U45967 (N_45967,N_44901,N_44184);
xor U45968 (N_45968,N_44927,N_44286);
nand U45969 (N_45969,N_44537,N_44697);
nand U45970 (N_45970,N_44523,N_44297);
nor U45971 (N_45971,N_44043,N_44163);
and U45972 (N_45972,N_44548,N_44205);
or U45973 (N_45973,N_44444,N_44594);
nand U45974 (N_45974,N_44049,N_44844);
and U45975 (N_45975,N_44592,N_44316);
nor U45976 (N_45976,N_44974,N_44534);
xor U45977 (N_45977,N_44480,N_44977);
and U45978 (N_45978,N_44661,N_44536);
and U45979 (N_45979,N_44191,N_44307);
xnor U45980 (N_45980,N_44398,N_44480);
nor U45981 (N_45981,N_44733,N_44753);
nor U45982 (N_45982,N_44594,N_44254);
and U45983 (N_45983,N_44572,N_44913);
xnor U45984 (N_45984,N_44180,N_44581);
xor U45985 (N_45985,N_44060,N_44847);
xnor U45986 (N_45986,N_44980,N_44853);
and U45987 (N_45987,N_44170,N_44472);
or U45988 (N_45988,N_44285,N_44034);
xnor U45989 (N_45989,N_44783,N_44791);
xor U45990 (N_45990,N_44172,N_44630);
nor U45991 (N_45991,N_44363,N_44436);
xor U45992 (N_45992,N_44287,N_44524);
and U45993 (N_45993,N_44288,N_44779);
nand U45994 (N_45994,N_44376,N_44137);
xor U45995 (N_45995,N_44336,N_44841);
xor U45996 (N_45996,N_44773,N_44743);
nor U45997 (N_45997,N_44737,N_44458);
xnor U45998 (N_45998,N_44462,N_44085);
xnor U45999 (N_45999,N_44225,N_44734);
or U46000 (N_46000,N_45366,N_45641);
or U46001 (N_46001,N_45777,N_45483);
or U46002 (N_46002,N_45530,N_45557);
nand U46003 (N_46003,N_45767,N_45762);
and U46004 (N_46004,N_45805,N_45093);
nor U46005 (N_46005,N_45968,N_45194);
or U46006 (N_46006,N_45311,N_45395);
nand U46007 (N_46007,N_45427,N_45669);
and U46008 (N_46008,N_45826,N_45345);
or U46009 (N_46009,N_45255,N_45109);
or U46010 (N_46010,N_45458,N_45516);
nor U46011 (N_46011,N_45682,N_45745);
xor U46012 (N_46012,N_45763,N_45084);
xor U46013 (N_46013,N_45390,N_45631);
nand U46014 (N_46014,N_45640,N_45121);
xor U46015 (N_46015,N_45620,N_45567);
nor U46016 (N_46016,N_45166,N_45170);
nand U46017 (N_46017,N_45987,N_45754);
nor U46018 (N_46018,N_45794,N_45058);
nor U46019 (N_46019,N_45611,N_45949);
xor U46020 (N_46020,N_45268,N_45560);
or U46021 (N_46021,N_45274,N_45228);
nor U46022 (N_46022,N_45145,N_45279);
nor U46023 (N_46023,N_45482,N_45350);
or U46024 (N_46024,N_45210,N_45385);
nor U46025 (N_46025,N_45764,N_45786);
and U46026 (N_46026,N_45928,N_45793);
nor U46027 (N_46027,N_45585,N_45479);
or U46028 (N_46028,N_45966,N_45893);
and U46029 (N_46029,N_45080,N_45334);
or U46030 (N_46030,N_45413,N_45549);
nor U46031 (N_46031,N_45832,N_45984);
nor U46032 (N_46032,N_45846,N_45357);
and U46033 (N_46033,N_45773,N_45340);
nor U46034 (N_46034,N_45378,N_45509);
and U46035 (N_46035,N_45705,N_45320);
nor U46036 (N_46036,N_45937,N_45975);
and U46037 (N_46037,N_45329,N_45811);
nand U46038 (N_46038,N_45223,N_45184);
and U46039 (N_46039,N_45533,N_45437);
xor U46040 (N_46040,N_45871,N_45591);
xnor U46041 (N_46041,N_45445,N_45040);
xnor U46042 (N_46042,N_45843,N_45717);
or U46043 (N_46043,N_45468,N_45330);
xnor U46044 (N_46044,N_45959,N_45208);
nor U46045 (N_46045,N_45162,N_45045);
and U46046 (N_46046,N_45603,N_45607);
or U46047 (N_46047,N_45995,N_45917);
and U46048 (N_46048,N_45033,N_45195);
and U46049 (N_46049,N_45853,N_45635);
nor U46050 (N_46050,N_45552,N_45790);
or U46051 (N_46051,N_45089,N_45155);
nand U46052 (N_46052,N_45851,N_45113);
or U46053 (N_46053,N_45450,N_45368);
xnor U46054 (N_46054,N_45683,N_45289);
nor U46055 (N_46055,N_45911,N_45012);
nand U46056 (N_46056,N_45880,N_45169);
xnor U46057 (N_46057,N_45182,N_45090);
xnor U46058 (N_46058,N_45868,N_45783);
or U46059 (N_46059,N_45927,N_45066);
and U46060 (N_46060,N_45087,N_45931);
nor U46061 (N_46061,N_45116,N_45018);
or U46062 (N_46062,N_45590,N_45602);
xor U46063 (N_46063,N_45784,N_45356);
and U46064 (N_46064,N_45092,N_45636);
xnor U46065 (N_46065,N_45349,N_45251);
nand U46066 (N_46066,N_45142,N_45081);
and U46067 (N_46067,N_45068,N_45808);
xor U46068 (N_46068,N_45220,N_45978);
nor U46069 (N_46069,N_45912,N_45840);
nor U46070 (N_46070,N_45028,N_45086);
and U46071 (N_46071,N_45726,N_45032);
or U46072 (N_46072,N_45095,N_45231);
or U46073 (N_46073,N_45367,N_45643);
nand U46074 (N_46074,N_45406,N_45855);
xor U46075 (N_46075,N_45555,N_45600);
xnor U46076 (N_46076,N_45875,N_45524);
xor U46077 (N_46077,N_45477,N_45891);
nand U46078 (N_46078,N_45275,N_45462);
nor U46079 (N_46079,N_45108,N_45377);
xor U46080 (N_46080,N_45577,N_45565);
or U46081 (N_46081,N_45532,N_45011);
xnor U46082 (N_46082,N_45670,N_45991);
and U46083 (N_46083,N_45594,N_45003);
nand U46084 (N_46084,N_45381,N_45394);
and U46085 (N_46085,N_45077,N_45860);
or U46086 (N_46086,N_45280,N_45302);
nand U46087 (N_46087,N_45229,N_45078);
nor U46088 (N_46088,N_45014,N_45921);
xnor U46089 (N_46089,N_45548,N_45709);
nor U46090 (N_46090,N_45490,N_45955);
xor U46091 (N_46091,N_45434,N_45006);
or U46092 (N_46092,N_45541,N_45511);
nor U46093 (N_46093,N_45624,N_45504);
nor U46094 (N_46094,N_45656,N_45206);
nand U46095 (N_46095,N_45866,N_45934);
xnor U46096 (N_46096,N_45785,N_45105);
nand U46097 (N_46097,N_45862,N_45114);
or U46098 (N_46098,N_45676,N_45134);
and U46099 (N_46099,N_45665,N_45465);
nor U46100 (N_46100,N_45969,N_45212);
or U46101 (N_46101,N_45430,N_45998);
and U46102 (N_46102,N_45841,N_45980);
nor U46103 (N_46103,N_45976,N_45159);
xnor U46104 (N_46104,N_45056,N_45568);
xnor U46105 (N_46105,N_45146,N_45503);
xor U46106 (N_46106,N_45130,N_45382);
and U46107 (N_46107,N_45307,N_45408);
and U46108 (N_46108,N_45753,N_45310);
nor U46109 (N_46109,N_45616,N_45833);
nand U46110 (N_46110,N_45236,N_45671);
xnor U46111 (N_46111,N_45123,N_45967);
nor U46112 (N_46112,N_45688,N_45495);
nor U46113 (N_46113,N_45667,N_45572);
and U46114 (N_46114,N_45262,N_45387);
xnor U46115 (N_46115,N_45375,N_45297);
or U46116 (N_46116,N_45443,N_45147);
and U46117 (N_46117,N_45501,N_45193);
or U46118 (N_46118,N_45749,N_45885);
nand U46119 (N_46119,N_45444,N_45813);
nand U46120 (N_46120,N_45192,N_45818);
nand U46121 (N_46121,N_45822,N_45454);
nor U46122 (N_46122,N_45303,N_45645);
and U46123 (N_46123,N_45471,N_45401);
xor U46124 (N_46124,N_45951,N_45812);
xor U46125 (N_46125,N_45321,N_45913);
or U46126 (N_46126,N_45935,N_45903);
or U46127 (N_46127,N_45569,N_45526);
nand U46128 (N_46128,N_45360,N_45448);
or U46129 (N_46129,N_45491,N_45772);
nand U46130 (N_46130,N_45988,N_45168);
nand U46131 (N_46131,N_45820,N_45947);
nand U46132 (N_46132,N_45725,N_45094);
and U46133 (N_46133,N_45617,N_45965);
nand U46134 (N_46134,N_45371,N_45718);
nor U46135 (N_46135,N_45070,N_45023);
or U46136 (N_46136,N_45249,N_45601);
xnor U46137 (N_46137,N_45977,N_45707);
and U46138 (N_46138,N_45218,N_45857);
nand U46139 (N_46139,N_45895,N_45496);
nand U46140 (N_46140,N_45514,N_45950);
or U46141 (N_46141,N_45703,N_45874);
or U46142 (N_46142,N_45691,N_45225);
xnor U46143 (N_46143,N_45063,N_45737);
nand U46144 (N_46144,N_45689,N_45901);
nor U46145 (N_46145,N_45447,N_45067);
nand U46146 (N_46146,N_45647,N_45655);
xnor U46147 (N_46147,N_45178,N_45740);
or U46148 (N_46148,N_45057,N_45488);
nand U46149 (N_46149,N_45831,N_45126);
and U46150 (N_46150,N_45803,N_45351);
and U46151 (N_46151,N_45799,N_45789);
xor U46152 (N_46152,N_45398,N_45886);
xor U46153 (N_46153,N_45022,N_45136);
nor U46154 (N_46154,N_45242,N_45191);
and U46155 (N_46155,N_45946,N_45456);
or U46156 (N_46156,N_45639,N_45838);
and U46157 (N_46157,N_45002,N_45579);
or U46158 (N_46158,N_45686,N_45884);
xnor U46159 (N_46159,N_45729,N_45796);
xnor U46160 (N_46160,N_45452,N_45628);
and U46161 (N_46161,N_45446,N_45453);
nor U46162 (N_46162,N_45051,N_45219);
nand U46163 (N_46163,N_45954,N_45128);
xor U46164 (N_46164,N_45677,N_45044);
xnor U46165 (N_46165,N_45285,N_45650);
and U46166 (N_46166,N_45088,N_45119);
or U46167 (N_46167,N_45404,N_45770);
or U46168 (N_46168,N_45111,N_45494);
nor U46169 (N_46169,N_45920,N_45905);
or U46170 (N_46170,N_45747,N_45979);
xnor U46171 (N_46171,N_45563,N_45042);
nand U46172 (N_46172,N_45957,N_45738);
nor U46173 (N_46173,N_45308,N_45981);
and U46174 (N_46174,N_45432,N_45273);
and U46175 (N_46175,N_45870,N_45420);
nand U46176 (N_46176,N_45863,N_45963);
and U46177 (N_46177,N_45700,N_45233);
nor U46178 (N_46178,N_45217,N_45806);
xor U46179 (N_46179,N_45464,N_45538);
xnor U46180 (N_46180,N_45389,N_45085);
nor U46181 (N_46181,N_45919,N_45484);
and U46182 (N_46182,N_45540,N_45055);
nor U46183 (N_46183,N_45199,N_45695);
nand U46184 (N_46184,N_45197,N_45227);
and U46185 (N_46185,N_45091,N_45347);
nand U46186 (N_46186,N_45414,N_45898);
xor U46187 (N_46187,N_45774,N_45005);
nand U46188 (N_46188,N_45506,N_45363);
xor U46189 (N_46189,N_45306,N_45160);
xnor U46190 (N_46190,N_45362,N_45889);
xnor U46191 (N_46191,N_45892,N_45266);
or U46192 (N_46192,N_45466,N_45507);
nand U46193 (N_46193,N_45623,N_45486);
or U46194 (N_46194,N_45732,N_45041);
nand U46195 (N_46195,N_45139,N_45668);
nand U46196 (N_46196,N_45721,N_45939);
nand U46197 (N_46197,N_45918,N_45396);
xor U46198 (N_46198,N_45276,N_45035);
nand U46199 (N_46199,N_45926,N_45888);
xnor U46200 (N_46200,N_45250,N_45151);
xnor U46201 (N_46201,N_45286,N_45010);
and U46202 (N_46202,N_45365,N_45263);
and U46203 (N_46203,N_45587,N_45060);
nor U46204 (N_46204,N_45828,N_45867);
or U46205 (N_46205,N_45554,N_45241);
xnor U46206 (N_46206,N_45188,N_45499);
nor U46207 (N_46207,N_45300,N_45036);
xnor U46208 (N_46208,N_45629,N_45632);
nand U46209 (N_46209,N_45973,N_45048);
nor U46210 (N_46210,N_45054,N_45714);
xnor U46211 (N_46211,N_45200,N_45776);
nor U46212 (N_46212,N_45314,N_45386);
and U46213 (N_46213,N_45296,N_45358);
nor U46214 (N_46214,N_45107,N_45025);
nand U46215 (N_46215,N_45269,N_45287);
and U46216 (N_46216,N_45883,N_45960);
nand U46217 (N_46217,N_45982,N_45301);
nor U46218 (N_46218,N_45834,N_45706);
nand U46219 (N_46219,N_45293,N_45797);
and U46220 (N_46220,N_45502,N_45174);
xor U46221 (N_46221,N_45110,N_45017);
nand U46222 (N_46222,N_45065,N_45369);
xnor U46223 (N_46223,N_45932,N_45138);
nand U46224 (N_46224,N_45693,N_45372);
nand U46225 (N_46225,N_45681,N_45472);
xor U46226 (N_46226,N_45692,N_45481);
xnor U46227 (N_46227,N_45167,N_45581);
nor U46228 (N_46228,N_45768,N_45710);
nand U46229 (N_46229,N_45171,N_45425);
nand U46230 (N_46230,N_45411,N_45312);
or U46231 (N_46231,N_45072,N_45062);
xnor U46232 (N_46232,N_45380,N_45124);
xor U46233 (N_46233,N_45235,N_45534);
nand U46234 (N_46234,N_45053,N_45735);
nand U46235 (N_46235,N_45202,N_45254);
nand U46236 (N_46236,N_45216,N_45144);
xnor U46237 (N_46237,N_45451,N_45324);
or U46238 (N_46238,N_45079,N_45364);
and U46239 (N_46239,N_45739,N_45264);
xor U46240 (N_46240,N_45476,N_45539);
and U46241 (N_46241,N_45234,N_45221);
nor U46242 (N_46242,N_45723,N_45614);
or U46243 (N_46243,N_45104,N_45335);
xnor U46244 (N_46244,N_45651,N_45659);
nor U46245 (N_46245,N_45131,N_45043);
xnor U46246 (N_46246,N_45583,N_45117);
or U46247 (N_46247,N_45457,N_45403);
xnor U46248 (N_46248,N_45315,N_45801);
nor U46249 (N_46249,N_45354,N_45150);
and U46250 (N_46250,N_45082,N_45802);
nand U46251 (N_46251,N_45734,N_45546);
and U46252 (N_46252,N_45712,N_45974);
nand U46253 (N_46253,N_45253,N_45240);
and U46254 (N_46254,N_45412,N_45589);
and U46255 (N_46255,N_45433,N_45282);
nand U46256 (N_46256,N_45837,N_45122);
nand U46257 (N_46257,N_45896,N_45948);
nor U46258 (N_46258,N_45698,N_45391);
nor U46259 (N_46259,N_45751,N_45115);
or U46260 (N_46260,N_45050,N_45654);
nor U46261 (N_46261,N_45943,N_45440);
and U46262 (N_46262,N_45983,N_45775);
nand U46263 (N_46263,N_45388,N_45239);
xnor U46264 (N_46264,N_45929,N_45810);
nand U46265 (N_46265,N_45759,N_45596);
xnor U46266 (N_46266,N_45525,N_45835);
nand U46267 (N_46267,N_45515,N_45519);
or U46268 (N_46268,N_45149,N_45076);
or U46269 (N_46269,N_45508,N_45244);
and U46270 (N_46270,N_45788,N_45933);
or U46271 (N_46271,N_45687,N_45597);
nor U46272 (N_46272,N_45845,N_45261);
nor U46273 (N_46273,N_45325,N_45646);
xor U46274 (N_46274,N_45630,N_45232);
xor U46275 (N_46275,N_45187,N_45708);
and U46276 (N_46276,N_45771,N_45945);
or U46277 (N_46277,N_45890,N_45696);
and U46278 (N_46278,N_45230,N_45711);
nor U46279 (N_46279,N_45848,N_45333);
or U46280 (N_46280,N_45971,N_45746);
or U46281 (N_46281,N_45103,N_45795);
nand U46282 (N_46282,N_45852,N_45102);
or U46283 (N_46283,N_45207,N_45816);
and U46284 (N_46284,N_45736,N_45319);
nand U46285 (N_46285,N_45719,N_45798);
nand U46286 (N_46286,N_45399,N_45148);
and U46287 (N_46287,N_45861,N_45172);
and U46288 (N_46288,N_45627,N_45346);
xnor U46289 (N_46289,N_45854,N_45267);
nand U46290 (N_46290,N_45694,N_45348);
xnor U46291 (N_46291,N_45608,N_45819);
xnor U46292 (N_46292,N_45899,N_45566);
nor U46293 (N_46293,N_45438,N_45397);
nor U46294 (N_46294,N_45101,N_45528);
nand U46295 (N_46295,N_45000,N_45498);
xnor U46296 (N_46296,N_45961,N_45634);
nor U46297 (N_46297,N_45165,N_45865);
nor U46298 (N_46298,N_45844,N_45426);
nand U46299 (N_46299,N_45814,N_45383);
nand U46300 (N_46300,N_45908,N_45485);
or U46301 (N_46301,N_45435,N_45294);
xnor U46302 (N_46302,N_45625,N_45588);
xor U46303 (N_46303,N_45823,N_45137);
or U46304 (N_46304,N_45742,N_45564);
nand U46305 (N_46305,N_45183,N_45545);
or U46306 (N_46306,N_45970,N_45100);
or U46307 (N_46307,N_45415,N_45638);
and U46308 (N_46308,N_45661,N_45850);
xnor U46309 (N_46309,N_45140,N_45914);
or U46310 (N_46310,N_45897,N_45859);
nand U46311 (N_46311,N_45480,N_45281);
nor U46312 (N_46312,N_45291,N_45370);
xnor U46313 (N_46313,N_45163,N_45904);
nor U46314 (N_46314,N_45407,N_45153);
nor U46315 (N_46315,N_45052,N_45141);
and U46316 (N_46316,N_45864,N_45522);
nand U46317 (N_46317,N_45653,N_45584);
or U46318 (N_46318,N_45922,N_45270);
and U46319 (N_46319,N_45361,N_45529);
or U46320 (N_46320,N_45295,N_45353);
xor U46321 (N_46321,N_45118,N_45283);
or U46322 (N_46322,N_45175,N_45298);
and U46323 (N_46323,N_45132,N_45059);
nand U46324 (N_46324,N_45675,N_45531);
nand U46325 (N_46325,N_45882,N_45180);
xnor U46326 (N_46326,N_45317,N_45644);
nand U46327 (N_46327,N_45909,N_45699);
or U46328 (N_46328,N_45400,N_45004);
nor U46329 (N_46329,N_45598,N_45605);
nand U46330 (N_46330,N_45143,N_45164);
or U46331 (N_46331,N_45026,N_45743);
nor U46332 (N_46332,N_45940,N_45173);
nand U46333 (N_46333,N_45326,N_45410);
or U46334 (N_46334,N_45599,N_45125);
or U46335 (N_46335,N_45550,N_45008);
nor U46336 (N_46336,N_45573,N_45021);
and U46337 (N_46337,N_45649,N_45064);
or U46338 (N_46338,N_45782,N_45642);
nand U46339 (N_46339,N_45684,N_45925);
or U46340 (N_46340,N_45209,N_45923);
xor U46341 (N_46341,N_45756,N_45500);
xor U46342 (N_46342,N_45313,N_45997);
nor U46343 (N_46343,N_45551,N_45907);
xor U46344 (N_46344,N_45439,N_45881);
xor U46345 (N_46345,N_45741,N_45527);
nand U46346 (N_46346,N_45757,N_45621);
and U46347 (N_46347,N_45074,N_45352);
and U46348 (N_46348,N_45520,N_45720);
xor U46349 (N_46349,N_45460,N_45277);
or U46350 (N_46350,N_45556,N_45730);
and U46351 (N_46351,N_45226,N_45990);
and U46352 (N_46352,N_45821,N_45536);
nand U46353 (N_46353,N_45373,N_45343);
nand U46354 (N_46354,N_45487,N_45030);
nand U46355 (N_46355,N_45936,N_45800);
xor U46356 (N_46356,N_45780,N_45384);
xor U46357 (N_46357,N_45817,N_45513);
or U46358 (N_46358,N_45994,N_45580);
nand U46359 (N_46359,N_45020,N_45576);
nor U46360 (N_46360,N_45697,N_45247);
nand U46361 (N_46361,N_45856,N_45039);
nor U46362 (N_46362,N_45133,N_45612);
xor U46363 (N_46363,N_45402,N_45129);
or U46364 (N_46364,N_45673,N_45878);
or U46365 (N_46365,N_45292,N_45455);
or U46366 (N_46366,N_45827,N_45423);
nor U46367 (N_46367,N_45727,N_45038);
xor U46368 (N_46368,N_45323,N_45222);
and U46369 (N_46369,N_45609,N_45941);
and U46370 (N_46370,N_45037,N_45493);
nor U46371 (N_46371,N_45544,N_45924);
and U46372 (N_46372,N_45179,N_45769);
nand U46373 (N_46373,N_45750,N_45678);
and U46374 (N_46374,N_45731,N_45309);
xor U46375 (N_46375,N_45213,N_45073);
or U46376 (N_46376,N_45258,N_45606);
nor U46377 (N_46377,N_45781,N_45672);
and U46378 (N_46378,N_45265,N_45964);
nand U46379 (N_46379,N_45290,N_45355);
and U46380 (N_46380,N_45374,N_45662);
nor U46381 (N_46381,N_45993,N_45766);
or U46382 (N_46382,N_45205,N_45574);
and U46383 (N_46383,N_45824,N_45553);
nand U46384 (N_46384,N_45761,N_45952);
or U46385 (N_46385,N_45953,N_45622);
nor U46386 (N_46386,N_45666,N_45648);
nor U46387 (N_46387,N_45046,N_45342);
nor U46388 (N_46388,N_45299,N_45492);
and U46389 (N_46389,N_45713,N_45724);
and U46390 (N_46390,N_45825,N_45318);
xor U46391 (N_46391,N_45099,N_45428);
nand U46392 (N_46392,N_45271,N_45475);
nand U46393 (N_46393,N_45702,N_45610);
xor U46394 (N_46394,N_45478,N_45535);
and U46395 (N_46395,N_45429,N_45009);
or U46396 (N_46396,N_45203,N_45422);
or U46397 (N_46397,N_45013,N_45256);
and U46398 (N_46398,N_45461,N_45956);
and U46399 (N_46399,N_45332,N_45186);
nor U46400 (N_46400,N_45047,N_45517);
and U46401 (N_46401,N_45778,N_45595);
xnor U46402 (N_46402,N_45996,N_45615);
nor U46403 (N_46403,N_45424,N_45523);
nand U46404 (N_46404,N_45019,N_45618);
and U46405 (N_46405,N_45792,N_45547);
or U46406 (N_46406,N_45196,N_45211);
nor U46407 (N_46407,N_45604,N_45327);
xor U46408 (N_46408,N_45586,N_45190);
and U46409 (N_46409,N_45071,N_45419);
and U46410 (N_46410,N_45685,N_45787);
and U46411 (N_46411,N_45663,N_45449);
xnor U46412 (N_46412,N_45906,N_45660);
and U46413 (N_46413,N_45379,N_45521);
or U46414 (N_46414,N_45257,N_45106);
xor U46415 (N_46415,N_45015,N_45942);
and U46416 (N_46416,N_45467,N_45376);
and U46417 (N_46417,N_45441,N_45189);
and U46418 (N_46418,N_45542,N_45652);
and U46419 (N_46419,N_45836,N_45999);
or U46420 (N_46420,N_45633,N_45930);
xnor U46421 (N_46421,N_45469,N_45972);
nand U46422 (N_46422,N_45181,N_45658);
nand U46423 (N_46423,N_45436,N_45879);
nor U46424 (N_46424,N_45260,N_45405);
nand U46425 (N_46425,N_45259,N_45755);
and U46426 (N_46426,N_45518,N_45944);
nand U46427 (N_46427,N_45034,N_45701);
and U46428 (N_46428,N_45992,N_45619);
nand U46429 (N_46429,N_45098,N_45765);
xnor U46430 (N_46430,N_45278,N_45716);
nand U46431 (N_46431,N_45284,N_45869);
nand U46432 (N_46432,N_45910,N_45127);
nand U46433 (N_46433,N_45578,N_45657);
or U46434 (N_46434,N_45198,N_45007);
xor U46435 (N_46435,N_45728,N_45593);
nor U46436 (N_46436,N_45872,N_45902);
nand U46437 (N_46437,N_45112,N_45680);
nor U46438 (N_46438,N_45152,N_45031);
or U46439 (N_46439,N_45049,N_45442);
or U46440 (N_46440,N_45061,N_45421);
and U46441 (N_46441,N_45418,N_45001);
or U46442 (N_46442,N_45842,N_45815);
or U46443 (N_46443,N_45679,N_45336);
xnor U46444 (N_46444,N_45473,N_45157);
nor U46445 (N_46445,N_45873,N_45915);
and U46446 (N_46446,N_45459,N_45431);
nand U46447 (N_46447,N_45704,N_45393);
or U46448 (N_46448,N_45339,N_45316);
nor U46449 (N_46449,N_45024,N_45204);
nand U46450 (N_46450,N_45887,N_45733);
or U46451 (N_46451,N_45288,N_45505);
or U46452 (N_46452,N_45075,N_45858);
and U46453 (N_46453,N_45744,N_45637);
or U46454 (N_46454,N_45154,N_45252);
xnor U46455 (N_46455,N_45849,N_45338);
nand U46456 (N_46456,N_45985,N_45246);
nand U46457 (N_46457,N_45416,N_45185);
or U46458 (N_46458,N_45029,N_45748);
nor U46459 (N_46459,N_45839,N_45916);
and U46460 (N_46460,N_45417,N_45986);
or U46461 (N_46461,N_45510,N_45409);
or U46462 (N_46462,N_45537,N_45359);
or U46463 (N_46463,N_45582,N_45674);
and U46464 (N_46464,N_45156,N_45592);
nand U46465 (N_46465,N_45807,N_45237);
nand U46466 (N_46466,N_45238,N_45120);
or U46467 (N_46467,N_45304,N_45664);
nor U46468 (N_46468,N_45248,N_45069);
and U46469 (N_46469,N_45135,N_45224);
nor U46470 (N_46470,N_45830,N_45847);
and U46471 (N_46471,N_45561,N_45331);
xor U46472 (N_46472,N_45328,N_45337);
or U46473 (N_46473,N_45690,N_45176);
nor U46474 (N_46474,N_45760,N_45272);
xor U46475 (N_46475,N_45245,N_45779);
nand U46476 (N_46476,N_45558,N_45305);
and U46477 (N_46477,N_45463,N_45243);
nand U46478 (N_46478,N_45626,N_45962);
or U46479 (N_46479,N_45177,N_45344);
xnor U46480 (N_46480,N_45894,N_45715);
nand U46481 (N_46481,N_45027,N_45083);
nand U46482 (N_46482,N_45322,N_45958);
nor U46483 (N_46483,N_45722,N_45470);
nand U46484 (N_46484,N_45791,N_45158);
nor U46485 (N_46485,N_45752,N_45214);
xor U46486 (N_46486,N_45559,N_45829);
or U46487 (N_46487,N_45877,N_45900);
nor U46488 (N_46488,N_45809,N_45938);
nand U46489 (N_46489,N_45489,N_45215);
nand U46490 (N_46490,N_45096,N_45571);
nor U46491 (N_46491,N_45497,N_45097);
or U46492 (N_46492,N_45758,N_45804);
or U46493 (N_46493,N_45201,N_45016);
nor U46494 (N_46494,N_45512,N_45570);
or U46495 (N_46495,N_45562,N_45341);
nor U46496 (N_46496,N_45543,N_45876);
nor U46497 (N_46497,N_45989,N_45392);
or U46498 (N_46498,N_45575,N_45474);
nand U46499 (N_46499,N_45613,N_45161);
and U46500 (N_46500,N_45881,N_45284);
xor U46501 (N_46501,N_45466,N_45655);
nand U46502 (N_46502,N_45959,N_45630);
xor U46503 (N_46503,N_45651,N_45477);
nand U46504 (N_46504,N_45121,N_45102);
nand U46505 (N_46505,N_45535,N_45738);
xor U46506 (N_46506,N_45182,N_45654);
and U46507 (N_46507,N_45470,N_45543);
nand U46508 (N_46508,N_45109,N_45163);
nand U46509 (N_46509,N_45923,N_45082);
nand U46510 (N_46510,N_45394,N_45094);
nand U46511 (N_46511,N_45806,N_45746);
xor U46512 (N_46512,N_45321,N_45552);
nand U46513 (N_46513,N_45439,N_45788);
and U46514 (N_46514,N_45912,N_45662);
nand U46515 (N_46515,N_45626,N_45015);
nand U46516 (N_46516,N_45679,N_45726);
nand U46517 (N_46517,N_45734,N_45399);
xnor U46518 (N_46518,N_45091,N_45987);
xnor U46519 (N_46519,N_45687,N_45050);
nor U46520 (N_46520,N_45466,N_45560);
and U46521 (N_46521,N_45682,N_45512);
nand U46522 (N_46522,N_45554,N_45330);
nor U46523 (N_46523,N_45065,N_45859);
nor U46524 (N_46524,N_45874,N_45239);
xor U46525 (N_46525,N_45389,N_45014);
xor U46526 (N_46526,N_45646,N_45884);
nor U46527 (N_46527,N_45940,N_45410);
or U46528 (N_46528,N_45844,N_45072);
xnor U46529 (N_46529,N_45773,N_45653);
nand U46530 (N_46530,N_45502,N_45129);
or U46531 (N_46531,N_45121,N_45355);
xor U46532 (N_46532,N_45951,N_45216);
xnor U46533 (N_46533,N_45482,N_45612);
xnor U46534 (N_46534,N_45301,N_45121);
xnor U46535 (N_46535,N_45587,N_45868);
or U46536 (N_46536,N_45658,N_45080);
nor U46537 (N_46537,N_45225,N_45014);
nor U46538 (N_46538,N_45414,N_45463);
and U46539 (N_46539,N_45537,N_45232);
and U46540 (N_46540,N_45343,N_45208);
nor U46541 (N_46541,N_45590,N_45701);
and U46542 (N_46542,N_45000,N_45373);
xnor U46543 (N_46543,N_45859,N_45683);
xnor U46544 (N_46544,N_45535,N_45204);
and U46545 (N_46545,N_45436,N_45272);
nor U46546 (N_46546,N_45370,N_45165);
or U46547 (N_46547,N_45816,N_45167);
nand U46548 (N_46548,N_45981,N_45485);
or U46549 (N_46549,N_45285,N_45535);
nor U46550 (N_46550,N_45852,N_45497);
nor U46551 (N_46551,N_45258,N_45203);
and U46552 (N_46552,N_45984,N_45724);
or U46553 (N_46553,N_45378,N_45818);
and U46554 (N_46554,N_45578,N_45551);
and U46555 (N_46555,N_45159,N_45002);
nor U46556 (N_46556,N_45344,N_45283);
nand U46557 (N_46557,N_45385,N_45083);
and U46558 (N_46558,N_45702,N_45191);
xnor U46559 (N_46559,N_45507,N_45868);
nand U46560 (N_46560,N_45105,N_45349);
nor U46561 (N_46561,N_45207,N_45668);
nor U46562 (N_46562,N_45729,N_45248);
or U46563 (N_46563,N_45438,N_45682);
nand U46564 (N_46564,N_45288,N_45355);
xnor U46565 (N_46565,N_45524,N_45372);
or U46566 (N_46566,N_45458,N_45932);
xor U46567 (N_46567,N_45833,N_45886);
nor U46568 (N_46568,N_45782,N_45309);
xnor U46569 (N_46569,N_45221,N_45795);
xor U46570 (N_46570,N_45150,N_45782);
nor U46571 (N_46571,N_45760,N_45374);
or U46572 (N_46572,N_45688,N_45897);
and U46573 (N_46573,N_45724,N_45828);
or U46574 (N_46574,N_45618,N_45226);
xor U46575 (N_46575,N_45963,N_45012);
nor U46576 (N_46576,N_45986,N_45344);
nand U46577 (N_46577,N_45601,N_45461);
nand U46578 (N_46578,N_45271,N_45620);
and U46579 (N_46579,N_45535,N_45556);
nand U46580 (N_46580,N_45631,N_45728);
nand U46581 (N_46581,N_45324,N_45617);
and U46582 (N_46582,N_45356,N_45231);
or U46583 (N_46583,N_45034,N_45399);
nor U46584 (N_46584,N_45411,N_45080);
nor U46585 (N_46585,N_45530,N_45202);
and U46586 (N_46586,N_45790,N_45279);
or U46587 (N_46587,N_45624,N_45193);
nor U46588 (N_46588,N_45304,N_45964);
xor U46589 (N_46589,N_45069,N_45638);
or U46590 (N_46590,N_45719,N_45371);
xor U46591 (N_46591,N_45906,N_45805);
nor U46592 (N_46592,N_45015,N_45380);
nand U46593 (N_46593,N_45080,N_45753);
nand U46594 (N_46594,N_45706,N_45531);
nand U46595 (N_46595,N_45049,N_45633);
nand U46596 (N_46596,N_45365,N_45130);
nand U46597 (N_46597,N_45495,N_45310);
nand U46598 (N_46598,N_45861,N_45710);
and U46599 (N_46599,N_45125,N_45119);
or U46600 (N_46600,N_45591,N_45848);
or U46601 (N_46601,N_45012,N_45370);
nor U46602 (N_46602,N_45935,N_45005);
and U46603 (N_46603,N_45444,N_45670);
nor U46604 (N_46604,N_45393,N_45561);
xor U46605 (N_46605,N_45052,N_45297);
xor U46606 (N_46606,N_45894,N_45244);
or U46607 (N_46607,N_45543,N_45322);
xnor U46608 (N_46608,N_45078,N_45944);
xnor U46609 (N_46609,N_45463,N_45992);
nor U46610 (N_46610,N_45087,N_45101);
and U46611 (N_46611,N_45572,N_45302);
nand U46612 (N_46612,N_45608,N_45211);
nand U46613 (N_46613,N_45761,N_45677);
xnor U46614 (N_46614,N_45791,N_45362);
xnor U46615 (N_46615,N_45567,N_45401);
and U46616 (N_46616,N_45318,N_45047);
nor U46617 (N_46617,N_45763,N_45002);
nor U46618 (N_46618,N_45389,N_45586);
or U46619 (N_46619,N_45873,N_45576);
nand U46620 (N_46620,N_45245,N_45961);
nor U46621 (N_46621,N_45656,N_45017);
xnor U46622 (N_46622,N_45752,N_45758);
and U46623 (N_46623,N_45143,N_45858);
xor U46624 (N_46624,N_45143,N_45928);
or U46625 (N_46625,N_45147,N_45696);
nor U46626 (N_46626,N_45699,N_45043);
xor U46627 (N_46627,N_45423,N_45738);
and U46628 (N_46628,N_45774,N_45155);
or U46629 (N_46629,N_45817,N_45347);
or U46630 (N_46630,N_45822,N_45937);
nand U46631 (N_46631,N_45966,N_45162);
nor U46632 (N_46632,N_45221,N_45197);
nor U46633 (N_46633,N_45809,N_45754);
nand U46634 (N_46634,N_45790,N_45455);
nor U46635 (N_46635,N_45714,N_45742);
or U46636 (N_46636,N_45720,N_45100);
or U46637 (N_46637,N_45830,N_45808);
nand U46638 (N_46638,N_45482,N_45004);
and U46639 (N_46639,N_45335,N_45492);
nand U46640 (N_46640,N_45474,N_45158);
nor U46641 (N_46641,N_45639,N_45269);
nor U46642 (N_46642,N_45102,N_45747);
or U46643 (N_46643,N_45011,N_45475);
and U46644 (N_46644,N_45362,N_45938);
nor U46645 (N_46645,N_45280,N_45042);
nor U46646 (N_46646,N_45703,N_45953);
nand U46647 (N_46647,N_45716,N_45297);
nand U46648 (N_46648,N_45724,N_45091);
and U46649 (N_46649,N_45772,N_45116);
or U46650 (N_46650,N_45408,N_45147);
nand U46651 (N_46651,N_45057,N_45944);
nand U46652 (N_46652,N_45006,N_45645);
and U46653 (N_46653,N_45918,N_45014);
and U46654 (N_46654,N_45496,N_45698);
xnor U46655 (N_46655,N_45402,N_45893);
nor U46656 (N_46656,N_45444,N_45682);
or U46657 (N_46657,N_45791,N_45658);
nand U46658 (N_46658,N_45730,N_45456);
nand U46659 (N_46659,N_45378,N_45813);
or U46660 (N_46660,N_45564,N_45928);
and U46661 (N_46661,N_45342,N_45709);
and U46662 (N_46662,N_45977,N_45319);
nor U46663 (N_46663,N_45345,N_45668);
nand U46664 (N_46664,N_45298,N_45389);
or U46665 (N_46665,N_45266,N_45234);
nor U46666 (N_46666,N_45956,N_45219);
or U46667 (N_46667,N_45096,N_45364);
nor U46668 (N_46668,N_45424,N_45467);
nor U46669 (N_46669,N_45846,N_45848);
and U46670 (N_46670,N_45302,N_45474);
nand U46671 (N_46671,N_45302,N_45455);
or U46672 (N_46672,N_45959,N_45573);
and U46673 (N_46673,N_45136,N_45040);
nor U46674 (N_46674,N_45356,N_45747);
nand U46675 (N_46675,N_45911,N_45023);
or U46676 (N_46676,N_45615,N_45051);
and U46677 (N_46677,N_45243,N_45762);
and U46678 (N_46678,N_45939,N_45081);
and U46679 (N_46679,N_45047,N_45307);
nand U46680 (N_46680,N_45190,N_45815);
or U46681 (N_46681,N_45264,N_45969);
and U46682 (N_46682,N_45201,N_45883);
nand U46683 (N_46683,N_45975,N_45463);
and U46684 (N_46684,N_45385,N_45976);
or U46685 (N_46685,N_45637,N_45026);
xnor U46686 (N_46686,N_45935,N_45741);
nor U46687 (N_46687,N_45389,N_45327);
or U46688 (N_46688,N_45847,N_45838);
nor U46689 (N_46689,N_45116,N_45103);
and U46690 (N_46690,N_45246,N_45915);
or U46691 (N_46691,N_45054,N_45619);
and U46692 (N_46692,N_45179,N_45503);
nand U46693 (N_46693,N_45577,N_45276);
nor U46694 (N_46694,N_45691,N_45834);
and U46695 (N_46695,N_45017,N_45131);
nand U46696 (N_46696,N_45091,N_45016);
nor U46697 (N_46697,N_45704,N_45069);
or U46698 (N_46698,N_45895,N_45029);
or U46699 (N_46699,N_45632,N_45045);
and U46700 (N_46700,N_45228,N_45466);
nor U46701 (N_46701,N_45678,N_45708);
nand U46702 (N_46702,N_45873,N_45953);
xor U46703 (N_46703,N_45472,N_45152);
nor U46704 (N_46704,N_45370,N_45844);
and U46705 (N_46705,N_45484,N_45850);
nor U46706 (N_46706,N_45653,N_45288);
nand U46707 (N_46707,N_45974,N_45993);
nand U46708 (N_46708,N_45584,N_45733);
nand U46709 (N_46709,N_45185,N_45700);
xor U46710 (N_46710,N_45341,N_45110);
nand U46711 (N_46711,N_45914,N_45010);
or U46712 (N_46712,N_45404,N_45860);
xor U46713 (N_46713,N_45528,N_45984);
xnor U46714 (N_46714,N_45637,N_45204);
or U46715 (N_46715,N_45194,N_45524);
and U46716 (N_46716,N_45851,N_45286);
nand U46717 (N_46717,N_45709,N_45094);
or U46718 (N_46718,N_45235,N_45392);
and U46719 (N_46719,N_45081,N_45811);
and U46720 (N_46720,N_45294,N_45683);
or U46721 (N_46721,N_45714,N_45234);
and U46722 (N_46722,N_45905,N_45518);
xor U46723 (N_46723,N_45999,N_45467);
xnor U46724 (N_46724,N_45604,N_45230);
nand U46725 (N_46725,N_45012,N_45537);
xnor U46726 (N_46726,N_45539,N_45286);
nand U46727 (N_46727,N_45194,N_45132);
nand U46728 (N_46728,N_45733,N_45180);
and U46729 (N_46729,N_45235,N_45817);
xnor U46730 (N_46730,N_45859,N_45163);
and U46731 (N_46731,N_45593,N_45092);
or U46732 (N_46732,N_45478,N_45509);
or U46733 (N_46733,N_45668,N_45331);
nand U46734 (N_46734,N_45056,N_45478);
nand U46735 (N_46735,N_45264,N_45234);
nor U46736 (N_46736,N_45042,N_45097);
nor U46737 (N_46737,N_45188,N_45562);
or U46738 (N_46738,N_45543,N_45775);
nand U46739 (N_46739,N_45268,N_45862);
and U46740 (N_46740,N_45718,N_45839);
and U46741 (N_46741,N_45937,N_45510);
or U46742 (N_46742,N_45971,N_45803);
or U46743 (N_46743,N_45437,N_45493);
nor U46744 (N_46744,N_45408,N_45981);
nand U46745 (N_46745,N_45904,N_45614);
xnor U46746 (N_46746,N_45904,N_45805);
xor U46747 (N_46747,N_45198,N_45357);
xnor U46748 (N_46748,N_45587,N_45627);
xnor U46749 (N_46749,N_45081,N_45779);
xor U46750 (N_46750,N_45319,N_45416);
or U46751 (N_46751,N_45422,N_45140);
nand U46752 (N_46752,N_45394,N_45314);
nand U46753 (N_46753,N_45257,N_45892);
xor U46754 (N_46754,N_45911,N_45974);
nand U46755 (N_46755,N_45577,N_45096);
xnor U46756 (N_46756,N_45076,N_45058);
nand U46757 (N_46757,N_45076,N_45862);
or U46758 (N_46758,N_45055,N_45347);
nand U46759 (N_46759,N_45466,N_45291);
or U46760 (N_46760,N_45471,N_45969);
and U46761 (N_46761,N_45479,N_45114);
or U46762 (N_46762,N_45476,N_45726);
nor U46763 (N_46763,N_45364,N_45513);
xor U46764 (N_46764,N_45065,N_45986);
nor U46765 (N_46765,N_45687,N_45861);
xnor U46766 (N_46766,N_45964,N_45902);
and U46767 (N_46767,N_45541,N_45009);
xor U46768 (N_46768,N_45700,N_45168);
nand U46769 (N_46769,N_45662,N_45539);
or U46770 (N_46770,N_45356,N_45701);
and U46771 (N_46771,N_45253,N_45248);
and U46772 (N_46772,N_45028,N_45914);
or U46773 (N_46773,N_45266,N_45742);
xnor U46774 (N_46774,N_45062,N_45314);
nand U46775 (N_46775,N_45859,N_45313);
xor U46776 (N_46776,N_45327,N_45048);
and U46777 (N_46777,N_45440,N_45690);
and U46778 (N_46778,N_45956,N_45725);
and U46779 (N_46779,N_45394,N_45203);
and U46780 (N_46780,N_45081,N_45010);
xor U46781 (N_46781,N_45564,N_45046);
or U46782 (N_46782,N_45331,N_45679);
xnor U46783 (N_46783,N_45419,N_45860);
nor U46784 (N_46784,N_45807,N_45574);
or U46785 (N_46785,N_45639,N_45499);
and U46786 (N_46786,N_45916,N_45266);
and U46787 (N_46787,N_45176,N_45519);
nor U46788 (N_46788,N_45517,N_45487);
nand U46789 (N_46789,N_45925,N_45793);
and U46790 (N_46790,N_45379,N_45904);
and U46791 (N_46791,N_45620,N_45021);
nand U46792 (N_46792,N_45701,N_45750);
nor U46793 (N_46793,N_45080,N_45864);
xnor U46794 (N_46794,N_45449,N_45066);
nor U46795 (N_46795,N_45754,N_45705);
nor U46796 (N_46796,N_45379,N_45253);
nor U46797 (N_46797,N_45220,N_45779);
and U46798 (N_46798,N_45780,N_45862);
nor U46799 (N_46799,N_45885,N_45665);
nor U46800 (N_46800,N_45302,N_45271);
xor U46801 (N_46801,N_45085,N_45125);
and U46802 (N_46802,N_45514,N_45016);
nand U46803 (N_46803,N_45582,N_45647);
nor U46804 (N_46804,N_45317,N_45503);
nand U46805 (N_46805,N_45569,N_45001);
and U46806 (N_46806,N_45767,N_45110);
nor U46807 (N_46807,N_45115,N_45463);
or U46808 (N_46808,N_45480,N_45089);
xnor U46809 (N_46809,N_45218,N_45450);
or U46810 (N_46810,N_45108,N_45150);
and U46811 (N_46811,N_45284,N_45777);
and U46812 (N_46812,N_45108,N_45429);
xnor U46813 (N_46813,N_45857,N_45337);
or U46814 (N_46814,N_45055,N_45976);
xnor U46815 (N_46815,N_45503,N_45782);
nor U46816 (N_46816,N_45892,N_45733);
or U46817 (N_46817,N_45007,N_45837);
or U46818 (N_46818,N_45222,N_45127);
or U46819 (N_46819,N_45051,N_45050);
nand U46820 (N_46820,N_45237,N_45388);
nand U46821 (N_46821,N_45979,N_45360);
nor U46822 (N_46822,N_45392,N_45101);
xnor U46823 (N_46823,N_45524,N_45074);
and U46824 (N_46824,N_45125,N_45123);
or U46825 (N_46825,N_45993,N_45787);
or U46826 (N_46826,N_45975,N_45788);
or U46827 (N_46827,N_45437,N_45670);
and U46828 (N_46828,N_45674,N_45678);
or U46829 (N_46829,N_45104,N_45899);
and U46830 (N_46830,N_45069,N_45424);
or U46831 (N_46831,N_45326,N_45882);
xnor U46832 (N_46832,N_45790,N_45833);
nor U46833 (N_46833,N_45743,N_45578);
or U46834 (N_46834,N_45379,N_45547);
and U46835 (N_46835,N_45214,N_45164);
nand U46836 (N_46836,N_45916,N_45110);
nor U46837 (N_46837,N_45614,N_45243);
nor U46838 (N_46838,N_45621,N_45162);
nand U46839 (N_46839,N_45561,N_45778);
nand U46840 (N_46840,N_45609,N_45931);
nor U46841 (N_46841,N_45855,N_45580);
nor U46842 (N_46842,N_45102,N_45340);
nor U46843 (N_46843,N_45567,N_45586);
xor U46844 (N_46844,N_45019,N_45524);
and U46845 (N_46845,N_45007,N_45015);
xor U46846 (N_46846,N_45788,N_45397);
nand U46847 (N_46847,N_45324,N_45327);
nand U46848 (N_46848,N_45360,N_45994);
and U46849 (N_46849,N_45729,N_45388);
nand U46850 (N_46850,N_45014,N_45062);
nor U46851 (N_46851,N_45822,N_45452);
nand U46852 (N_46852,N_45524,N_45932);
or U46853 (N_46853,N_45185,N_45121);
nor U46854 (N_46854,N_45813,N_45279);
or U46855 (N_46855,N_45327,N_45740);
or U46856 (N_46856,N_45704,N_45514);
xor U46857 (N_46857,N_45164,N_45571);
nor U46858 (N_46858,N_45235,N_45507);
and U46859 (N_46859,N_45518,N_45539);
xnor U46860 (N_46860,N_45620,N_45765);
xnor U46861 (N_46861,N_45250,N_45917);
nor U46862 (N_46862,N_45265,N_45850);
or U46863 (N_46863,N_45096,N_45952);
nand U46864 (N_46864,N_45565,N_45642);
or U46865 (N_46865,N_45469,N_45279);
nand U46866 (N_46866,N_45645,N_45848);
nand U46867 (N_46867,N_45031,N_45101);
and U46868 (N_46868,N_45799,N_45743);
or U46869 (N_46869,N_45736,N_45040);
nand U46870 (N_46870,N_45100,N_45633);
xnor U46871 (N_46871,N_45003,N_45966);
xnor U46872 (N_46872,N_45385,N_45211);
xnor U46873 (N_46873,N_45037,N_45517);
xor U46874 (N_46874,N_45152,N_45288);
nor U46875 (N_46875,N_45397,N_45970);
nor U46876 (N_46876,N_45675,N_45288);
and U46877 (N_46877,N_45332,N_45189);
nand U46878 (N_46878,N_45950,N_45674);
nor U46879 (N_46879,N_45105,N_45846);
and U46880 (N_46880,N_45563,N_45498);
nand U46881 (N_46881,N_45673,N_45083);
and U46882 (N_46882,N_45936,N_45323);
xor U46883 (N_46883,N_45499,N_45061);
nand U46884 (N_46884,N_45567,N_45528);
nand U46885 (N_46885,N_45144,N_45571);
and U46886 (N_46886,N_45642,N_45277);
nor U46887 (N_46887,N_45487,N_45922);
nand U46888 (N_46888,N_45749,N_45553);
nand U46889 (N_46889,N_45948,N_45172);
or U46890 (N_46890,N_45031,N_45328);
or U46891 (N_46891,N_45370,N_45053);
xnor U46892 (N_46892,N_45732,N_45794);
and U46893 (N_46893,N_45817,N_45090);
xnor U46894 (N_46894,N_45632,N_45283);
nor U46895 (N_46895,N_45905,N_45452);
nand U46896 (N_46896,N_45463,N_45916);
and U46897 (N_46897,N_45082,N_45728);
and U46898 (N_46898,N_45922,N_45124);
nand U46899 (N_46899,N_45311,N_45713);
xnor U46900 (N_46900,N_45185,N_45292);
or U46901 (N_46901,N_45124,N_45289);
nand U46902 (N_46902,N_45302,N_45016);
and U46903 (N_46903,N_45520,N_45442);
nand U46904 (N_46904,N_45272,N_45792);
nor U46905 (N_46905,N_45576,N_45846);
nor U46906 (N_46906,N_45779,N_45591);
or U46907 (N_46907,N_45700,N_45061);
nand U46908 (N_46908,N_45968,N_45128);
nand U46909 (N_46909,N_45708,N_45263);
or U46910 (N_46910,N_45825,N_45066);
and U46911 (N_46911,N_45064,N_45296);
xor U46912 (N_46912,N_45889,N_45409);
nor U46913 (N_46913,N_45623,N_45822);
xnor U46914 (N_46914,N_45386,N_45473);
nand U46915 (N_46915,N_45603,N_45977);
and U46916 (N_46916,N_45184,N_45366);
or U46917 (N_46917,N_45683,N_45178);
or U46918 (N_46918,N_45497,N_45502);
xor U46919 (N_46919,N_45162,N_45820);
nor U46920 (N_46920,N_45481,N_45845);
nor U46921 (N_46921,N_45726,N_45079);
and U46922 (N_46922,N_45777,N_45052);
or U46923 (N_46923,N_45549,N_45056);
nand U46924 (N_46924,N_45121,N_45174);
nand U46925 (N_46925,N_45213,N_45805);
nand U46926 (N_46926,N_45394,N_45794);
nor U46927 (N_46927,N_45737,N_45566);
nor U46928 (N_46928,N_45693,N_45033);
nor U46929 (N_46929,N_45900,N_45761);
xnor U46930 (N_46930,N_45078,N_45806);
nor U46931 (N_46931,N_45777,N_45062);
or U46932 (N_46932,N_45149,N_45234);
xnor U46933 (N_46933,N_45449,N_45474);
xor U46934 (N_46934,N_45966,N_45953);
xnor U46935 (N_46935,N_45888,N_45066);
xor U46936 (N_46936,N_45085,N_45836);
nor U46937 (N_46937,N_45724,N_45814);
nor U46938 (N_46938,N_45466,N_45630);
or U46939 (N_46939,N_45124,N_45713);
nor U46940 (N_46940,N_45442,N_45274);
nor U46941 (N_46941,N_45725,N_45327);
nor U46942 (N_46942,N_45788,N_45686);
nor U46943 (N_46943,N_45776,N_45036);
nor U46944 (N_46944,N_45371,N_45411);
xnor U46945 (N_46945,N_45550,N_45289);
nand U46946 (N_46946,N_45913,N_45757);
xnor U46947 (N_46947,N_45005,N_45811);
and U46948 (N_46948,N_45102,N_45305);
nand U46949 (N_46949,N_45195,N_45902);
and U46950 (N_46950,N_45888,N_45674);
and U46951 (N_46951,N_45519,N_45415);
nand U46952 (N_46952,N_45184,N_45560);
xnor U46953 (N_46953,N_45557,N_45213);
nor U46954 (N_46954,N_45105,N_45959);
xor U46955 (N_46955,N_45682,N_45717);
nand U46956 (N_46956,N_45061,N_45143);
xnor U46957 (N_46957,N_45838,N_45004);
nor U46958 (N_46958,N_45212,N_45058);
nor U46959 (N_46959,N_45306,N_45466);
nand U46960 (N_46960,N_45739,N_45821);
or U46961 (N_46961,N_45895,N_45840);
nand U46962 (N_46962,N_45413,N_45943);
and U46963 (N_46963,N_45540,N_45670);
nor U46964 (N_46964,N_45317,N_45851);
nand U46965 (N_46965,N_45581,N_45447);
nor U46966 (N_46966,N_45878,N_45466);
xor U46967 (N_46967,N_45057,N_45312);
or U46968 (N_46968,N_45227,N_45921);
and U46969 (N_46969,N_45097,N_45253);
nand U46970 (N_46970,N_45061,N_45221);
and U46971 (N_46971,N_45418,N_45502);
nor U46972 (N_46972,N_45741,N_45954);
xor U46973 (N_46973,N_45226,N_45680);
and U46974 (N_46974,N_45462,N_45126);
nor U46975 (N_46975,N_45894,N_45960);
or U46976 (N_46976,N_45945,N_45127);
and U46977 (N_46977,N_45916,N_45745);
and U46978 (N_46978,N_45576,N_45337);
or U46979 (N_46979,N_45143,N_45870);
or U46980 (N_46980,N_45670,N_45259);
nor U46981 (N_46981,N_45848,N_45987);
or U46982 (N_46982,N_45349,N_45919);
nand U46983 (N_46983,N_45634,N_45157);
xor U46984 (N_46984,N_45901,N_45219);
nand U46985 (N_46985,N_45211,N_45658);
nand U46986 (N_46986,N_45207,N_45659);
xnor U46987 (N_46987,N_45936,N_45715);
or U46988 (N_46988,N_45151,N_45650);
and U46989 (N_46989,N_45499,N_45575);
and U46990 (N_46990,N_45677,N_45753);
nor U46991 (N_46991,N_45920,N_45676);
or U46992 (N_46992,N_45698,N_45511);
or U46993 (N_46993,N_45948,N_45816);
and U46994 (N_46994,N_45596,N_45920);
nand U46995 (N_46995,N_45571,N_45614);
or U46996 (N_46996,N_45826,N_45399);
and U46997 (N_46997,N_45717,N_45407);
and U46998 (N_46998,N_45429,N_45662);
xor U46999 (N_46999,N_45651,N_45711);
and U47000 (N_47000,N_46672,N_46302);
xnor U47001 (N_47001,N_46195,N_46210);
and U47002 (N_47002,N_46814,N_46006);
xor U47003 (N_47003,N_46886,N_46413);
and U47004 (N_47004,N_46965,N_46240);
nand U47005 (N_47005,N_46534,N_46407);
nor U47006 (N_47006,N_46930,N_46744);
xor U47007 (N_47007,N_46802,N_46219);
or U47008 (N_47008,N_46949,N_46855);
xor U47009 (N_47009,N_46258,N_46308);
nand U47010 (N_47010,N_46472,N_46818);
and U47011 (N_47011,N_46858,N_46435);
and U47012 (N_47012,N_46446,N_46840);
and U47013 (N_47013,N_46135,N_46951);
nor U47014 (N_47014,N_46616,N_46755);
nand U47015 (N_47015,N_46944,N_46562);
nor U47016 (N_47016,N_46244,N_46971);
nand U47017 (N_47017,N_46202,N_46106);
nand U47018 (N_47018,N_46058,N_46664);
nor U47019 (N_47019,N_46297,N_46735);
xnor U47020 (N_47020,N_46265,N_46163);
xor U47021 (N_47021,N_46272,N_46552);
or U47022 (N_47022,N_46402,N_46774);
and U47023 (N_47023,N_46715,N_46498);
nand U47024 (N_47024,N_46507,N_46206);
or U47025 (N_47025,N_46686,N_46259);
nand U47026 (N_47026,N_46282,N_46129);
xnor U47027 (N_47027,N_46845,N_46980);
xor U47028 (N_47028,N_46540,N_46662);
nor U47029 (N_47029,N_46076,N_46403);
and U47030 (N_47030,N_46139,N_46758);
xor U47031 (N_47031,N_46303,N_46532);
nor U47032 (N_47032,N_46600,N_46409);
xnor U47033 (N_47033,N_46416,N_46669);
nand U47034 (N_47034,N_46471,N_46494);
nor U47035 (N_47035,N_46008,N_46271);
xnor U47036 (N_47036,N_46362,N_46717);
nor U47037 (N_47037,N_46236,N_46518);
and U47038 (N_47038,N_46025,N_46536);
or U47039 (N_47039,N_46701,N_46889);
and U47040 (N_47040,N_46681,N_46398);
xnor U47041 (N_47041,N_46942,N_46036);
or U47042 (N_47042,N_46826,N_46350);
and U47043 (N_47043,N_46527,N_46964);
nand U47044 (N_47044,N_46997,N_46181);
xor U47045 (N_47045,N_46795,N_46477);
nand U47046 (N_47046,N_46974,N_46671);
nor U47047 (N_47047,N_46174,N_46637);
and U47048 (N_47048,N_46685,N_46380);
xnor U47049 (N_47049,N_46233,N_46473);
nand U47050 (N_47050,N_46328,N_46411);
nand U47051 (N_47051,N_46267,N_46724);
and U47052 (N_47052,N_46449,N_46952);
and U47053 (N_47053,N_46079,N_46738);
nor U47054 (N_47054,N_46491,N_46687);
or U47055 (N_47055,N_46234,N_46332);
xnor U47056 (N_47056,N_46970,N_46682);
nor U47057 (N_47057,N_46955,N_46270);
nand U47058 (N_47058,N_46074,N_46617);
or U47059 (N_47059,N_46392,N_46882);
nor U47060 (N_47060,N_46393,N_46582);
nor U47061 (N_47061,N_46389,N_46920);
nor U47062 (N_47062,N_46620,N_46847);
nand U47063 (N_47063,N_46316,N_46199);
nor U47064 (N_47064,N_46209,N_46038);
or U47065 (N_47065,N_46182,N_46089);
nand U47066 (N_47066,N_46512,N_46431);
xor U47067 (N_47067,N_46556,N_46447);
and U47068 (N_47068,N_46545,N_46529);
or U47069 (N_47069,N_46485,N_46732);
nand U47070 (N_47070,N_46301,N_46595);
nor U47071 (N_47071,N_46243,N_46313);
and U47072 (N_47072,N_46461,N_46465);
and U47073 (N_47073,N_46678,N_46694);
and U47074 (N_47074,N_46417,N_46126);
xor U47075 (N_47075,N_46024,N_46923);
nor U47076 (N_47076,N_46223,N_46330);
nand U47077 (N_47077,N_46780,N_46849);
nor U47078 (N_47078,N_46130,N_46204);
or U47079 (N_47079,N_46810,N_46456);
nor U47080 (N_47080,N_46081,N_46549);
or U47081 (N_47081,N_46629,N_46364);
nand U47082 (N_47082,N_46722,N_46880);
nand U47083 (N_47083,N_46224,N_46357);
or U47084 (N_47084,N_46056,N_46570);
and U47085 (N_47085,N_46028,N_46142);
xnor U47086 (N_47086,N_46844,N_46731);
xor U47087 (N_47087,N_46155,N_46022);
xnor U47088 (N_47088,N_46464,N_46688);
xor U47089 (N_47089,N_46913,N_46490);
xor U47090 (N_47090,N_46092,N_46828);
or U47091 (N_47091,N_46111,N_46019);
nand U47092 (N_47092,N_46116,N_46679);
or U47093 (N_47093,N_46586,N_46021);
and U47094 (N_47094,N_46467,N_46231);
nor U47095 (N_47095,N_46706,N_46596);
xnor U47096 (N_47096,N_46597,N_46053);
nand U47097 (N_47097,N_46711,N_46304);
xor U47098 (N_47098,N_46221,N_46439);
and U47099 (N_47099,N_46991,N_46378);
nand U47100 (N_47100,N_46692,N_46911);
or U47101 (N_47101,N_46091,N_46228);
xor U47102 (N_47102,N_46768,N_46311);
nor U47103 (N_47103,N_46026,N_46329);
nand U47104 (N_47104,N_46254,N_46343);
xnor U47105 (N_47105,N_46697,N_46804);
and U47106 (N_47106,N_46245,N_46599);
and U47107 (N_47107,N_46482,N_46852);
xor U47108 (N_47108,N_46300,N_46385);
or U47109 (N_47109,N_46932,N_46422);
xnor U47110 (N_47110,N_46030,N_46784);
xor U47111 (N_47111,N_46086,N_46203);
nand U47112 (N_47112,N_46788,N_46843);
nand U47113 (N_47113,N_46314,N_46631);
or U47114 (N_47114,N_46754,N_46376);
nand U47115 (N_47115,N_46906,N_46121);
xor U47116 (N_47116,N_46587,N_46544);
nor U47117 (N_47117,N_46215,N_46041);
or U47118 (N_47118,N_46198,N_46785);
and U47119 (N_47119,N_46418,N_46381);
nand U47120 (N_47120,N_46729,N_46993);
nor U47121 (N_47121,N_46741,N_46830);
nor U47122 (N_47122,N_46339,N_46324);
and U47123 (N_47123,N_46757,N_46640);
nor U47124 (N_47124,N_46972,N_46288);
nand U47125 (N_47125,N_46745,N_46521);
nor U47126 (N_47126,N_46000,N_46226);
and U47127 (N_47127,N_46611,N_46766);
or U47128 (N_47128,N_46255,N_46211);
nor U47129 (N_47129,N_46504,N_46014);
or U47130 (N_47130,N_46348,N_46391);
nand U47131 (N_47131,N_46172,N_46702);
and U47132 (N_47132,N_46800,N_46190);
nand U47133 (N_47133,N_46138,N_46306);
and U47134 (N_47134,N_46317,N_46957);
nand U47135 (N_47135,N_46811,N_46607);
nor U47136 (N_47136,N_46767,N_46763);
xnor U47137 (N_47137,N_46150,N_46977);
nor U47138 (N_47138,N_46289,N_46644);
or U47139 (N_47139,N_46740,N_46815);
nand U47140 (N_47140,N_46157,N_46619);
nand U47141 (N_47141,N_46356,N_46775);
or U47142 (N_47142,N_46105,N_46824);
and U47143 (N_47143,N_46425,N_46872);
xor U47144 (N_47144,N_46854,N_46127);
and U47145 (N_47145,N_46821,N_46564);
and U47146 (N_47146,N_46382,N_46469);
nand U47147 (N_47147,N_46069,N_46051);
or U47148 (N_47148,N_46037,N_46414);
xnor U47149 (N_47149,N_46333,N_46273);
or U47150 (N_47150,N_46720,N_46756);
or U47151 (N_47151,N_46394,N_46630);
or U47152 (N_47152,N_46865,N_46778);
nand U47153 (N_47153,N_46693,N_46175);
or U47154 (N_47154,N_46238,N_46819);
and U47155 (N_47155,N_46261,N_46430);
or U47156 (N_47156,N_46633,N_46487);
xor U47157 (N_47157,N_46113,N_46003);
nand U47158 (N_47158,N_46230,N_46191);
nand U47159 (N_47159,N_46299,N_46445);
nor U47160 (N_47160,N_46514,N_46695);
or U47161 (N_47161,N_46420,N_46760);
or U47162 (N_47162,N_46836,N_46613);
or U47163 (N_47163,N_46408,N_46039);
nand U47164 (N_47164,N_46438,N_46569);
nand U47165 (N_47165,N_46989,N_46506);
nor U47166 (N_47166,N_46716,N_46460);
or U47167 (N_47167,N_46383,N_46601);
xor U47168 (N_47168,N_46268,N_46145);
and U47169 (N_47169,N_46825,N_46981);
nand U47170 (N_47170,N_46603,N_46887);
and U47171 (N_47171,N_46978,N_46007);
or U47172 (N_47172,N_46747,N_46718);
or U47173 (N_47173,N_46577,N_46759);
or U47174 (N_47174,N_46023,N_46530);
nand U47175 (N_47175,N_46433,N_46165);
nor U47176 (N_47176,N_46752,N_46167);
or U47177 (N_47177,N_46765,N_46178);
nor U47178 (N_47178,N_46123,N_46667);
and U47179 (N_47179,N_46873,N_46018);
nor U47180 (N_47180,N_46112,N_46428);
nor U47181 (N_47181,N_46698,N_46166);
or U47182 (N_47182,N_46598,N_46782);
and U47183 (N_47183,N_46884,N_46876);
nand U47184 (N_47184,N_46415,N_46188);
or U47185 (N_47185,N_46340,N_46612);
xnor U47186 (N_47186,N_46798,N_46922);
nor U47187 (N_47187,N_46973,N_46327);
xnor U47188 (N_47188,N_46010,N_46483);
nor U47189 (N_47189,N_46152,N_46961);
or U47190 (N_47190,N_46859,N_46095);
nor U47191 (N_47191,N_46946,N_46635);
nand U47192 (N_47192,N_46052,N_46065);
nor U47193 (N_47193,N_46550,N_46345);
or U47194 (N_47194,N_46160,N_46256);
xnor U47195 (N_47195,N_46220,N_46526);
or U47196 (N_47196,N_46158,N_46059);
nor U47197 (N_47197,N_46032,N_46813);
and U47198 (N_47198,N_46929,N_46714);
and U47199 (N_47199,N_46277,N_46325);
and U47200 (N_47200,N_46820,N_46434);
and U47201 (N_47201,N_46673,N_46676);
nor U47202 (N_47202,N_46962,N_46251);
or U47203 (N_47203,N_46823,N_46733);
and U47204 (N_47204,N_46419,N_46563);
nand U47205 (N_47205,N_46636,N_46185);
xor U47206 (N_47206,N_46794,N_46846);
or U47207 (N_47207,N_46388,N_46149);
or U47208 (N_47208,N_46996,N_46384);
or U47209 (N_47209,N_46309,N_46594);
and U47210 (N_47210,N_46968,N_46869);
nor U47211 (N_47211,N_46368,N_46558);
and U47212 (N_47212,N_46294,N_46960);
nor U47213 (N_47213,N_46864,N_46634);
or U47214 (N_47214,N_46454,N_46806);
xor U47215 (N_47215,N_46786,N_46031);
or U47216 (N_47216,N_46822,N_46371);
nor U47217 (N_47217,N_46591,N_46837);
and U47218 (N_47218,N_46196,N_46797);
nand U47219 (N_47219,N_46073,N_46541);
and U47220 (N_47220,N_46279,N_46197);
nand U47221 (N_47221,N_46568,N_46901);
nor U47222 (N_47222,N_46040,N_46513);
nand U47223 (N_47223,N_46359,N_46264);
nand U47224 (N_47224,N_46621,N_46857);
nand U47225 (N_47225,N_46638,N_46119);
xnor U47226 (N_47226,N_46066,N_46958);
and U47227 (N_47227,N_46781,N_46280);
xnor U47228 (N_47228,N_46100,N_46812);
nor U47229 (N_47229,N_46665,N_46169);
and U47230 (N_47230,N_46683,N_46015);
nor U47231 (N_47231,N_46444,N_46777);
nand U47232 (N_47232,N_46432,N_46147);
nor U47233 (N_47233,N_46331,N_46290);
nor U47234 (N_47234,N_46475,N_46184);
or U47235 (N_47235,N_46914,N_46684);
xor U47236 (N_47236,N_46011,N_46235);
nand U47237 (N_47237,N_46805,N_46248);
nor U47238 (N_47238,N_46832,N_46423);
nand U47239 (N_47239,N_46538,N_46358);
nor U47240 (N_47240,N_46450,N_46842);
and U47241 (N_47241,N_46173,N_46250);
nand U47242 (N_47242,N_46346,N_46013);
and U47243 (N_47243,N_46275,N_46278);
nand U47244 (N_47244,N_46124,N_46020);
nor U47245 (N_47245,N_46218,N_46510);
xnor U47246 (N_47246,N_46817,N_46286);
nor U47247 (N_47247,N_46925,N_46001);
xor U47248 (N_47248,N_46892,N_46164);
nand U47249 (N_47249,N_46296,N_46917);
and U47250 (N_47250,N_46480,N_46187);
and U47251 (N_47251,N_46560,N_46421);
and U47252 (N_47252,N_46808,N_46452);
and U47253 (N_47253,N_46468,N_46557);
nand U47254 (N_47254,N_46347,N_46749);
or U47255 (N_47255,N_46373,N_46652);
and U47256 (N_47256,N_46322,N_46940);
or U47257 (N_47257,N_46883,N_46336);
xnor U47258 (N_47258,N_46956,N_46533);
or U47259 (N_47259,N_46606,N_46535);
xor U47260 (N_47260,N_46796,N_46156);
nor U47261 (N_47261,N_46426,N_46751);
nand U47262 (N_47262,N_46728,N_46748);
or U47263 (N_47263,N_46943,N_46877);
nor U47264 (N_47264,N_46950,N_46710);
nor U47265 (N_47265,N_46554,N_46581);
and U47266 (N_47266,N_46707,N_46829);
nor U47267 (N_47267,N_46252,N_46353);
and U47268 (N_47268,N_46084,N_46799);
nor U47269 (N_47269,N_46068,N_46372);
xnor U47270 (N_47270,N_46519,N_46213);
xor U47271 (N_47271,N_46650,N_46994);
xor U47272 (N_47272,N_46436,N_46517);
xor U47273 (N_47273,N_46651,N_46400);
or U47274 (N_47274,N_46017,N_46609);
nand U47275 (N_47275,N_46374,N_46488);
nand U47276 (N_47276,N_46938,N_46761);
nor U47277 (N_47277,N_46576,N_46140);
nand U47278 (N_47278,N_46131,N_46674);
or U47279 (N_47279,N_46548,N_46237);
nor U47280 (N_47280,N_46632,N_46624);
nor U47281 (N_47281,N_46072,N_46988);
nand U47282 (N_47282,N_46208,N_46476);
nor U47283 (N_47283,N_46110,N_46916);
and U47284 (N_47284,N_46390,N_46338);
nand U47285 (N_47285,N_46967,N_46976);
nand U47286 (N_47286,N_46508,N_46143);
nand U47287 (N_47287,N_46457,N_46704);
nor U47288 (N_47288,N_46666,N_46623);
xnor U47289 (N_47289,N_46492,N_46451);
and U47290 (N_47290,N_46941,N_46263);
xor U47291 (N_47291,N_46424,N_46497);
or U47292 (N_47292,N_46257,N_46625);
nand U47293 (N_47293,N_46982,N_46262);
nand U47294 (N_47294,N_46719,N_46983);
and U47295 (N_47295,N_46566,N_46764);
nor U47296 (N_47296,N_46241,N_46985);
nand U47297 (N_47297,N_46342,N_46055);
nand U47298 (N_47298,N_46578,N_46910);
nor U47299 (N_47299,N_46907,N_46361);
nor U47300 (N_47300,N_46660,N_46878);
or U47301 (N_47301,N_46016,N_46034);
or U47302 (N_47302,N_46903,N_46397);
nand U47303 (N_47303,N_46405,N_46712);
and U47304 (N_47304,N_46648,N_46680);
nor U47305 (N_47305,N_46212,N_46816);
xor U47306 (N_47306,N_46459,N_46875);
nor U47307 (N_47307,N_46850,N_46101);
and U47308 (N_47308,N_46939,N_46699);
xor U47309 (N_47309,N_46762,N_46723);
xor U47310 (N_47310,N_46305,N_46108);
nor U47311 (N_47311,N_46522,N_46075);
or U47312 (N_47312,N_46194,N_46148);
nor U47313 (N_47313,N_46049,N_46628);
nor U47314 (N_47314,N_46885,N_46269);
nor U47315 (N_47315,N_46060,N_46159);
or U47316 (N_47316,N_46335,N_46260);
xnor U47317 (N_47317,N_46354,N_46363);
nor U47318 (N_47318,N_46659,N_46501);
nand U47319 (N_47319,N_46122,N_46936);
nor U47320 (N_47320,N_46900,N_46984);
nor U47321 (N_47321,N_46310,N_46750);
nor U47322 (N_47322,N_46730,N_46183);
nand U47323 (N_47323,N_46897,N_46365);
or U47324 (N_47324,N_46689,N_46312);
and U47325 (N_47325,N_46908,N_46239);
nand U47326 (N_47326,N_46713,N_46050);
or U47327 (N_47327,N_46746,N_46427);
or U47328 (N_47328,N_46912,N_46047);
xor U47329 (N_47329,N_46180,N_46489);
nand U47330 (N_47330,N_46429,N_46990);
nand U47331 (N_47331,N_46888,N_46344);
xnor U47332 (N_47332,N_46406,N_46789);
nor U47333 (N_47333,N_46769,N_46565);
xnor U47334 (N_47334,N_46690,N_46954);
nor U47335 (N_47335,N_46663,N_46721);
nor U47336 (N_47336,N_46440,N_46868);
nand U47337 (N_47337,N_46899,N_46743);
and U47338 (N_47338,N_46109,N_46103);
xor U47339 (N_47339,N_46098,N_46229);
nor U47340 (N_47340,N_46904,N_46396);
xor U47341 (N_47341,N_46862,N_46179);
or U47342 (N_47342,N_46283,N_46734);
and U47343 (N_47343,N_46367,N_46249);
nand U47344 (N_47344,N_46851,N_46608);
or U47345 (N_47345,N_46064,N_46493);
and U47346 (N_47346,N_46045,N_46531);
and U47347 (N_47347,N_46216,N_46463);
nor U47348 (N_47348,N_46584,N_46057);
or U47349 (N_47349,N_46905,N_46120);
and U47350 (N_47350,N_46931,N_46453);
and U47351 (N_47351,N_46386,N_46499);
xnor U47352 (N_47352,N_46622,N_46177);
xor U47353 (N_47353,N_46863,N_46838);
and U47354 (N_47354,N_46547,N_46352);
or U47355 (N_47355,N_46894,N_46002);
and U47356 (N_47356,N_46736,N_46442);
and U47357 (N_47357,N_46470,N_46004);
xnor U47358 (N_47358,N_46959,N_46088);
and U47359 (N_47359,N_46515,N_46890);
or U47360 (N_47360,N_46661,N_46592);
and U47361 (N_47361,N_46835,N_46627);
and U47362 (N_47362,N_46062,N_46044);
or U47363 (N_47363,N_46771,N_46067);
nor U47364 (N_47364,N_46144,N_46319);
nand U47365 (N_47365,N_46242,N_46999);
nand U47366 (N_47366,N_46189,N_46926);
or U47367 (N_47367,N_46496,N_46227);
nor U47368 (N_47368,N_46827,N_46902);
xor U47369 (N_47369,N_46998,N_46500);
and U47370 (N_47370,N_46874,N_46085);
nand U47371 (N_47371,N_46455,N_46675);
nor U47372 (N_47372,N_46610,N_46104);
nor U47373 (N_47373,N_46787,N_46953);
nand U47374 (N_47374,N_46793,N_46321);
xor U47375 (N_47375,N_46776,N_46404);
xor U47376 (N_47376,N_46575,N_46292);
nand U47377 (N_47377,N_46895,N_46870);
and U47378 (N_47378,N_46969,N_46573);
xor U47379 (N_47379,N_46042,N_46035);
xor U47380 (N_47380,N_46834,N_46207);
nor U47381 (N_47381,N_46839,N_46726);
nor U47382 (N_47382,N_46871,N_46503);
xor U47383 (N_47383,N_46979,N_46520);
xnor U47384 (N_47384,N_46856,N_46162);
and U47385 (N_47385,N_46080,N_46479);
and U47386 (N_47386,N_46571,N_46029);
nor U47387 (N_47387,N_46315,N_46090);
nor U47388 (N_47388,N_46898,N_46928);
nand U47389 (N_47389,N_46247,N_46341);
and U47390 (N_47390,N_46337,N_46070);
xor U47391 (N_47391,N_46287,N_46186);
xor U47392 (N_47392,N_46645,N_46511);
nand U47393 (N_47393,N_46580,N_46474);
or U47394 (N_47394,N_46809,N_46643);
nor U47395 (N_47395,N_46168,N_46546);
nor U47396 (N_47396,N_46077,N_46918);
or U47397 (N_47397,N_46274,N_46935);
nand U47398 (N_47398,N_46656,N_46551);
xnor U47399 (N_47399,N_46653,N_46739);
nand U47400 (N_47400,N_46448,N_46118);
nor U47401 (N_47401,N_46861,N_46909);
nand U47402 (N_47402,N_46083,N_46590);
and U47403 (N_47403,N_46443,N_46934);
and U47404 (N_47404,N_46604,N_46132);
and U47405 (N_47405,N_46246,N_46395);
xor U47406 (N_47406,N_46133,N_46915);
nor U47407 (N_47407,N_46176,N_46700);
and U47408 (N_47408,N_46375,N_46355);
nor U47409 (N_47409,N_46919,N_46696);
and U47410 (N_47410,N_46360,N_46867);
xor U47411 (N_47411,N_46136,N_46703);
nor U47412 (N_47412,N_46987,N_46366);
xnor U47413 (N_47413,N_46641,N_46523);
or U47414 (N_47414,N_46803,N_46525);
nand U47415 (N_47415,N_46567,N_46141);
nor U47416 (N_47416,N_46285,N_46945);
and U47417 (N_47417,N_46896,N_46102);
and U47418 (N_47418,N_46772,N_46071);
xor U47419 (N_47419,N_46553,N_46585);
nor U47420 (N_47420,N_46096,N_46655);
nand U47421 (N_47421,N_46893,N_46537);
xor U47422 (N_47422,N_46539,N_46705);
and U47423 (N_47423,N_46379,N_46561);
or U47424 (N_47424,N_46054,N_46377);
nand U47425 (N_47425,N_46351,N_46589);
and U47426 (N_47426,N_46853,N_46481);
and U47427 (N_47427,N_46170,N_46437);
or U47428 (N_47428,N_46253,N_46048);
and U47429 (N_47429,N_46307,N_46125);
nand U47430 (N_47430,N_46012,N_46115);
nor U47431 (N_47431,N_46323,N_46921);
and U47432 (N_47432,N_46043,N_46266);
xor U47433 (N_47433,N_46284,N_46293);
or U47434 (N_47434,N_46369,N_46107);
xnor U47435 (N_47435,N_46458,N_46214);
nand U47436 (N_47436,N_46975,N_46128);
nand U47437 (N_47437,N_46543,N_46320);
or U47438 (N_47438,N_46927,N_46232);
or U47439 (N_47439,N_46937,N_46318);
nand U47440 (N_47440,N_46281,N_46790);
nor U47441 (N_47441,N_46879,N_46615);
or U47442 (N_47442,N_46725,N_46401);
nor U47443 (N_47443,N_46027,N_46201);
and U47444 (N_47444,N_46502,N_46555);
or U47445 (N_47445,N_46791,N_46947);
and U47446 (N_47446,N_46779,N_46657);
nand U47447 (N_47447,N_46205,N_46154);
nor U47448 (N_47448,N_46495,N_46559);
and U47449 (N_47449,N_46099,N_46061);
xnor U47450 (N_47450,N_46093,N_46117);
or U47451 (N_47451,N_46370,N_46677);
nor U47452 (N_47452,N_46792,N_46114);
xnor U47453 (N_47453,N_46963,N_46833);
nand U47454 (N_47454,N_46524,N_46626);
or U47455 (N_47455,N_46509,N_46866);
xor U47456 (N_47456,N_46146,N_46670);
nor U47457 (N_47457,N_46992,N_46222);
nand U47458 (N_47458,N_46412,N_46737);
or U47459 (N_47459,N_46528,N_46082);
and U47460 (N_47460,N_46484,N_46995);
or U47461 (N_47461,N_46078,N_46753);
and U47462 (N_47462,N_46891,N_46614);
nor U47463 (N_47463,N_46924,N_46691);
nor U47464 (N_47464,N_46593,N_46848);
nor U47465 (N_47465,N_46334,N_46046);
xor U47466 (N_47466,N_46807,N_46709);
or U47467 (N_47467,N_46986,N_46727);
nor U47468 (N_47468,N_46646,N_46579);
nor U47469 (N_47469,N_46387,N_46572);
nand U47470 (N_47470,N_46276,N_46642);
or U47471 (N_47471,N_46192,N_46295);
nand U47472 (N_47472,N_46708,N_46200);
nor U47473 (N_47473,N_46618,N_46161);
xnor U47474 (N_47474,N_46583,N_46639);
and U47475 (N_47475,N_46466,N_46574);
nand U47476 (N_47476,N_46063,N_46087);
or U47477 (N_47477,N_46349,N_46881);
nor U47478 (N_47478,N_46933,N_46668);
nor U47479 (N_47479,N_46505,N_46097);
and U47480 (N_47480,N_46151,N_46486);
and U47481 (N_47481,N_46948,N_46225);
or U47482 (N_47482,N_46217,N_46742);
xor U47483 (N_47483,N_46478,N_46860);
and U47484 (N_47484,N_46542,N_46009);
xnor U47485 (N_47485,N_46649,N_46094);
and U47486 (N_47486,N_46193,N_46291);
nor U47487 (N_47487,N_46783,N_46770);
or U47488 (N_47488,N_46658,N_46966);
nor U47489 (N_47489,N_46171,N_46831);
nor U47490 (N_47490,N_46137,N_46647);
and U47491 (N_47491,N_46462,N_46033);
nand U47492 (N_47492,N_46841,N_46602);
nand U47493 (N_47493,N_46134,N_46399);
and U47494 (N_47494,N_46516,N_46801);
nor U47495 (N_47495,N_46410,N_46773);
xnor U47496 (N_47496,N_46654,N_46298);
nor U47497 (N_47497,N_46153,N_46588);
nand U47498 (N_47498,N_46005,N_46441);
nand U47499 (N_47499,N_46326,N_46605);
or U47500 (N_47500,N_46553,N_46800);
xnor U47501 (N_47501,N_46836,N_46755);
nand U47502 (N_47502,N_46747,N_46727);
or U47503 (N_47503,N_46911,N_46056);
xnor U47504 (N_47504,N_46357,N_46863);
xor U47505 (N_47505,N_46028,N_46760);
nand U47506 (N_47506,N_46680,N_46164);
xnor U47507 (N_47507,N_46249,N_46555);
nand U47508 (N_47508,N_46655,N_46796);
nand U47509 (N_47509,N_46516,N_46921);
nand U47510 (N_47510,N_46287,N_46204);
and U47511 (N_47511,N_46259,N_46952);
xor U47512 (N_47512,N_46625,N_46608);
nor U47513 (N_47513,N_46670,N_46960);
or U47514 (N_47514,N_46873,N_46811);
nand U47515 (N_47515,N_46099,N_46313);
or U47516 (N_47516,N_46205,N_46649);
nor U47517 (N_47517,N_46254,N_46567);
and U47518 (N_47518,N_46380,N_46952);
or U47519 (N_47519,N_46243,N_46098);
and U47520 (N_47520,N_46466,N_46192);
and U47521 (N_47521,N_46177,N_46499);
nand U47522 (N_47522,N_46132,N_46554);
xnor U47523 (N_47523,N_46347,N_46013);
nor U47524 (N_47524,N_46707,N_46663);
nor U47525 (N_47525,N_46096,N_46900);
xor U47526 (N_47526,N_46973,N_46312);
and U47527 (N_47527,N_46868,N_46109);
or U47528 (N_47528,N_46567,N_46811);
and U47529 (N_47529,N_46229,N_46270);
or U47530 (N_47530,N_46698,N_46603);
and U47531 (N_47531,N_46680,N_46555);
nand U47532 (N_47532,N_46272,N_46613);
nand U47533 (N_47533,N_46836,N_46366);
xor U47534 (N_47534,N_46745,N_46269);
nand U47535 (N_47535,N_46307,N_46272);
and U47536 (N_47536,N_46863,N_46151);
or U47537 (N_47537,N_46131,N_46156);
nor U47538 (N_47538,N_46201,N_46753);
and U47539 (N_47539,N_46493,N_46591);
and U47540 (N_47540,N_46934,N_46148);
nand U47541 (N_47541,N_46152,N_46344);
xnor U47542 (N_47542,N_46047,N_46277);
xnor U47543 (N_47543,N_46993,N_46724);
nor U47544 (N_47544,N_46631,N_46876);
nor U47545 (N_47545,N_46665,N_46317);
nor U47546 (N_47546,N_46159,N_46901);
nor U47547 (N_47547,N_46774,N_46792);
nand U47548 (N_47548,N_46640,N_46843);
and U47549 (N_47549,N_46663,N_46411);
and U47550 (N_47550,N_46558,N_46153);
nand U47551 (N_47551,N_46763,N_46668);
nor U47552 (N_47552,N_46921,N_46047);
xor U47553 (N_47553,N_46923,N_46065);
xor U47554 (N_47554,N_46192,N_46078);
xor U47555 (N_47555,N_46777,N_46234);
xnor U47556 (N_47556,N_46055,N_46174);
nor U47557 (N_47557,N_46224,N_46776);
or U47558 (N_47558,N_46959,N_46702);
or U47559 (N_47559,N_46870,N_46102);
and U47560 (N_47560,N_46034,N_46341);
nand U47561 (N_47561,N_46222,N_46397);
or U47562 (N_47562,N_46693,N_46231);
nor U47563 (N_47563,N_46354,N_46644);
and U47564 (N_47564,N_46356,N_46079);
xor U47565 (N_47565,N_46252,N_46727);
or U47566 (N_47566,N_46050,N_46004);
xnor U47567 (N_47567,N_46084,N_46544);
xnor U47568 (N_47568,N_46317,N_46906);
xnor U47569 (N_47569,N_46529,N_46337);
or U47570 (N_47570,N_46855,N_46337);
xnor U47571 (N_47571,N_46190,N_46804);
nand U47572 (N_47572,N_46160,N_46321);
and U47573 (N_47573,N_46659,N_46816);
nor U47574 (N_47574,N_46941,N_46464);
or U47575 (N_47575,N_46038,N_46258);
or U47576 (N_47576,N_46545,N_46514);
nor U47577 (N_47577,N_46349,N_46173);
nand U47578 (N_47578,N_46833,N_46870);
xor U47579 (N_47579,N_46271,N_46833);
xnor U47580 (N_47580,N_46283,N_46758);
xor U47581 (N_47581,N_46267,N_46567);
or U47582 (N_47582,N_46463,N_46486);
nor U47583 (N_47583,N_46610,N_46027);
or U47584 (N_47584,N_46129,N_46559);
nor U47585 (N_47585,N_46443,N_46907);
nand U47586 (N_47586,N_46473,N_46397);
xor U47587 (N_47587,N_46288,N_46629);
and U47588 (N_47588,N_46737,N_46832);
and U47589 (N_47589,N_46034,N_46190);
xnor U47590 (N_47590,N_46147,N_46904);
and U47591 (N_47591,N_46041,N_46522);
nor U47592 (N_47592,N_46870,N_46123);
or U47593 (N_47593,N_46940,N_46738);
or U47594 (N_47594,N_46298,N_46954);
and U47595 (N_47595,N_46486,N_46445);
xnor U47596 (N_47596,N_46964,N_46569);
nand U47597 (N_47597,N_46237,N_46670);
or U47598 (N_47598,N_46868,N_46025);
xnor U47599 (N_47599,N_46144,N_46590);
or U47600 (N_47600,N_46633,N_46841);
nand U47601 (N_47601,N_46605,N_46016);
nand U47602 (N_47602,N_46692,N_46009);
nor U47603 (N_47603,N_46397,N_46731);
and U47604 (N_47604,N_46361,N_46122);
or U47605 (N_47605,N_46836,N_46523);
or U47606 (N_47606,N_46659,N_46209);
nor U47607 (N_47607,N_46814,N_46510);
xor U47608 (N_47608,N_46896,N_46313);
nor U47609 (N_47609,N_46397,N_46486);
nand U47610 (N_47610,N_46994,N_46992);
or U47611 (N_47611,N_46694,N_46114);
or U47612 (N_47612,N_46710,N_46025);
xnor U47613 (N_47613,N_46253,N_46511);
xor U47614 (N_47614,N_46327,N_46296);
or U47615 (N_47615,N_46893,N_46760);
nand U47616 (N_47616,N_46802,N_46679);
xor U47617 (N_47617,N_46956,N_46710);
xnor U47618 (N_47618,N_46221,N_46118);
and U47619 (N_47619,N_46171,N_46906);
nor U47620 (N_47620,N_46266,N_46841);
xor U47621 (N_47621,N_46379,N_46131);
or U47622 (N_47622,N_46933,N_46783);
nor U47623 (N_47623,N_46957,N_46024);
or U47624 (N_47624,N_46213,N_46390);
xor U47625 (N_47625,N_46839,N_46915);
or U47626 (N_47626,N_46282,N_46922);
nand U47627 (N_47627,N_46668,N_46021);
xnor U47628 (N_47628,N_46399,N_46366);
xnor U47629 (N_47629,N_46832,N_46647);
or U47630 (N_47630,N_46341,N_46023);
xor U47631 (N_47631,N_46842,N_46876);
nand U47632 (N_47632,N_46172,N_46917);
xor U47633 (N_47633,N_46839,N_46842);
xor U47634 (N_47634,N_46416,N_46084);
and U47635 (N_47635,N_46487,N_46039);
xnor U47636 (N_47636,N_46803,N_46548);
and U47637 (N_47637,N_46126,N_46331);
nand U47638 (N_47638,N_46507,N_46212);
or U47639 (N_47639,N_46232,N_46349);
or U47640 (N_47640,N_46797,N_46311);
or U47641 (N_47641,N_46588,N_46932);
or U47642 (N_47642,N_46155,N_46903);
nand U47643 (N_47643,N_46260,N_46395);
xnor U47644 (N_47644,N_46564,N_46039);
nand U47645 (N_47645,N_46025,N_46951);
and U47646 (N_47646,N_46804,N_46775);
nand U47647 (N_47647,N_46077,N_46126);
and U47648 (N_47648,N_46712,N_46104);
nor U47649 (N_47649,N_46305,N_46176);
nand U47650 (N_47650,N_46014,N_46465);
nor U47651 (N_47651,N_46733,N_46975);
nand U47652 (N_47652,N_46183,N_46221);
xnor U47653 (N_47653,N_46162,N_46442);
or U47654 (N_47654,N_46939,N_46401);
nand U47655 (N_47655,N_46790,N_46522);
xnor U47656 (N_47656,N_46997,N_46628);
xor U47657 (N_47657,N_46469,N_46668);
nand U47658 (N_47658,N_46802,N_46376);
and U47659 (N_47659,N_46089,N_46773);
nor U47660 (N_47660,N_46534,N_46320);
nor U47661 (N_47661,N_46093,N_46636);
nor U47662 (N_47662,N_46528,N_46110);
xor U47663 (N_47663,N_46458,N_46837);
xor U47664 (N_47664,N_46488,N_46258);
or U47665 (N_47665,N_46036,N_46228);
nand U47666 (N_47666,N_46933,N_46551);
nand U47667 (N_47667,N_46744,N_46025);
nor U47668 (N_47668,N_46991,N_46835);
and U47669 (N_47669,N_46337,N_46631);
and U47670 (N_47670,N_46867,N_46531);
or U47671 (N_47671,N_46076,N_46941);
or U47672 (N_47672,N_46548,N_46635);
nor U47673 (N_47673,N_46631,N_46515);
xnor U47674 (N_47674,N_46713,N_46449);
nor U47675 (N_47675,N_46706,N_46337);
and U47676 (N_47676,N_46033,N_46964);
and U47677 (N_47677,N_46587,N_46806);
nand U47678 (N_47678,N_46846,N_46757);
and U47679 (N_47679,N_46869,N_46531);
and U47680 (N_47680,N_46550,N_46266);
and U47681 (N_47681,N_46038,N_46046);
or U47682 (N_47682,N_46965,N_46330);
nor U47683 (N_47683,N_46916,N_46729);
xor U47684 (N_47684,N_46661,N_46329);
or U47685 (N_47685,N_46530,N_46418);
xor U47686 (N_47686,N_46698,N_46345);
and U47687 (N_47687,N_46060,N_46736);
or U47688 (N_47688,N_46467,N_46803);
nor U47689 (N_47689,N_46226,N_46517);
and U47690 (N_47690,N_46792,N_46606);
and U47691 (N_47691,N_46465,N_46299);
or U47692 (N_47692,N_46755,N_46792);
and U47693 (N_47693,N_46003,N_46027);
and U47694 (N_47694,N_46077,N_46983);
and U47695 (N_47695,N_46148,N_46696);
and U47696 (N_47696,N_46565,N_46548);
or U47697 (N_47697,N_46433,N_46267);
nor U47698 (N_47698,N_46501,N_46561);
nor U47699 (N_47699,N_46304,N_46020);
nand U47700 (N_47700,N_46165,N_46875);
nor U47701 (N_47701,N_46008,N_46087);
nor U47702 (N_47702,N_46514,N_46078);
nor U47703 (N_47703,N_46147,N_46912);
xnor U47704 (N_47704,N_46405,N_46305);
or U47705 (N_47705,N_46478,N_46799);
nor U47706 (N_47706,N_46250,N_46119);
nor U47707 (N_47707,N_46625,N_46995);
nand U47708 (N_47708,N_46628,N_46120);
and U47709 (N_47709,N_46685,N_46026);
nor U47710 (N_47710,N_46533,N_46020);
and U47711 (N_47711,N_46620,N_46496);
nand U47712 (N_47712,N_46940,N_46740);
nor U47713 (N_47713,N_46785,N_46529);
or U47714 (N_47714,N_46264,N_46427);
xnor U47715 (N_47715,N_46074,N_46298);
or U47716 (N_47716,N_46889,N_46909);
and U47717 (N_47717,N_46403,N_46952);
nor U47718 (N_47718,N_46538,N_46509);
and U47719 (N_47719,N_46071,N_46220);
or U47720 (N_47720,N_46899,N_46470);
or U47721 (N_47721,N_46427,N_46887);
nor U47722 (N_47722,N_46667,N_46197);
nand U47723 (N_47723,N_46671,N_46152);
or U47724 (N_47724,N_46958,N_46924);
or U47725 (N_47725,N_46669,N_46012);
or U47726 (N_47726,N_46322,N_46284);
nand U47727 (N_47727,N_46156,N_46106);
nand U47728 (N_47728,N_46889,N_46375);
or U47729 (N_47729,N_46176,N_46278);
nand U47730 (N_47730,N_46905,N_46948);
and U47731 (N_47731,N_46560,N_46386);
or U47732 (N_47732,N_46726,N_46401);
and U47733 (N_47733,N_46794,N_46864);
and U47734 (N_47734,N_46593,N_46234);
nand U47735 (N_47735,N_46298,N_46032);
xor U47736 (N_47736,N_46110,N_46565);
and U47737 (N_47737,N_46564,N_46614);
or U47738 (N_47738,N_46437,N_46525);
xnor U47739 (N_47739,N_46951,N_46685);
nand U47740 (N_47740,N_46494,N_46966);
or U47741 (N_47741,N_46352,N_46157);
nand U47742 (N_47742,N_46526,N_46774);
xor U47743 (N_47743,N_46249,N_46043);
xnor U47744 (N_47744,N_46642,N_46000);
xor U47745 (N_47745,N_46379,N_46827);
and U47746 (N_47746,N_46122,N_46684);
nand U47747 (N_47747,N_46151,N_46886);
nand U47748 (N_47748,N_46150,N_46339);
nor U47749 (N_47749,N_46097,N_46636);
or U47750 (N_47750,N_46281,N_46669);
nand U47751 (N_47751,N_46589,N_46291);
and U47752 (N_47752,N_46290,N_46889);
and U47753 (N_47753,N_46551,N_46739);
and U47754 (N_47754,N_46885,N_46342);
xor U47755 (N_47755,N_46061,N_46414);
xnor U47756 (N_47756,N_46653,N_46754);
and U47757 (N_47757,N_46579,N_46859);
and U47758 (N_47758,N_46770,N_46706);
nor U47759 (N_47759,N_46239,N_46104);
nand U47760 (N_47760,N_46211,N_46163);
or U47761 (N_47761,N_46760,N_46530);
xor U47762 (N_47762,N_46277,N_46268);
nand U47763 (N_47763,N_46148,N_46608);
nor U47764 (N_47764,N_46695,N_46671);
xnor U47765 (N_47765,N_46996,N_46185);
nor U47766 (N_47766,N_46476,N_46066);
xor U47767 (N_47767,N_46189,N_46980);
xnor U47768 (N_47768,N_46832,N_46731);
nand U47769 (N_47769,N_46037,N_46864);
xnor U47770 (N_47770,N_46148,N_46478);
nor U47771 (N_47771,N_46375,N_46790);
nor U47772 (N_47772,N_46081,N_46537);
xor U47773 (N_47773,N_46507,N_46429);
nor U47774 (N_47774,N_46062,N_46600);
xnor U47775 (N_47775,N_46536,N_46979);
and U47776 (N_47776,N_46678,N_46704);
or U47777 (N_47777,N_46629,N_46102);
nand U47778 (N_47778,N_46094,N_46446);
xnor U47779 (N_47779,N_46925,N_46013);
and U47780 (N_47780,N_46183,N_46820);
nand U47781 (N_47781,N_46379,N_46437);
nand U47782 (N_47782,N_46168,N_46694);
xnor U47783 (N_47783,N_46301,N_46857);
nand U47784 (N_47784,N_46134,N_46711);
nand U47785 (N_47785,N_46144,N_46923);
or U47786 (N_47786,N_46578,N_46737);
nor U47787 (N_47787,N_46939,N_46270);
nand U47788 (N_47788,N_46235,N_46556);
nand U47789 (N_47789,N_46309,N_46206);
xor U47790 (N_47790,N_46919,N_46827);
nor U47791 (N_47791,N_46497,N_46268);
xnor U47792 (N_47792,N_46581,N_46388);
xnor U47793 (N_47793,N_46124,N_46951);
or U47794 (N_47794,N_46230,N_46036);
nand U47795 (N_47795,N_46911,N_46810);
xnor U47796 (N_47796,N_46683,N_46701);
nor U47797 (N_47797,N_46200,N_46372);
nand U47798 (N_47798,N_46062,N_46357);
and U47799 (N_47799,N_46038,N_46344);
xor U47800 (N_47800,N_46328,N_46710);
nor U47801 (N_47801,N_46233,N_46190);
or U47802 (N_47802,N_46056,N_46767);
nor U47803 (N_47803,N_46367,N_46241);
nor U47804 (N_47804,N_46085,N_46707);
or U47805 (N_47805,N_46846,N_46686);
nand U47806 (N_47806,N_46381,N_46514);
nor U47807 (N_47807,N_46438,N_46697);
or U47808 (N_47808,N_46827,N_46265);
xor U47809 (N_47809,N_46391,N_46521);
or U47810 (N_47810,N_46676,N_46949);
or U47811 (N_47811,N_46170,N_46652);
nor U47812 (N_47812,N_46473,N_46631);
and U47813 (N_47813,N_46794,N_46947);
nor U47814 (N_47814,N_46087,N_46888);
nand U47815 (N_47815,N_46200,N_46733);
or U47816 (N_47816,N_46059,N_46460);
or U47817 (N_47817,N_46481,N_46260);
xnor U47818 (N_47818,N_46701,N_46559);
nand U47819 (N_47819,N_46265,N_46303);
and U47820 (N_47820,N_46155,N_46006);
and U47821 (N_47821,N_46789,N_46808);
nand U47822 (N_47822,N_46445,N_46012);
xnor U47823 (N_47823,N_46458,N_46595);
xor U47824 (N_47824,N_46759,N_46457);
nand U47825 (N_47825,N_46644,N_46146);
xor U47826 (N_47826,N_46279,N_46169);
or U47827 (N_47827,N_46508,N_46712);
and U47828 (N_47828,N_46448,N_46117);
nand U47829 (N_47829,N_46081,N_46484);
xnor U47830 (N_47830,N_46192,N_46919);
xor U47831 (N_47831,N_46763,N_46794);
nand U47832 (N_47832,N_46716,N_46588);
xor U47833 (N_47833,N_46305,N_46157);
nor U47834 (N_47834,N_46567,N_46723);
or U47835 (N_47835,N_46005,N_46921);
nand U47836 (N_47836,N_46622,N_46606);
nor U47837 (N_47837,N_46482,N_46283);
nand U47838 (N_47838,N_46801,N_46316);
and U47839 (N_47839,N_46703,N_46673);
xnor U47840 (N_47840,N_46350,N_46907);
and U47841 (N_47841,N_46921,N_46726);
xor U47842 (N_47842,N_46117,N_46377);
and U47843 (N_47843,N_46044,N_46543);
nor U47844 (N_47844,N_46088,N_46305);
xor U47845 (N_47845,N_46839,N_46551);
or U47846 (N_47846,N_46501,N_46431);
xnor U47847 (N_47847,N_46264,N_46669);
nand U47848 (N_47848,N_46481,N_46557);
xnor U47849 (N_47849,N_46711,N_46096);
nor U47850 (N_47850,N_46267,N_46098);
nand U47851 (N_47851,N_46235,N_46983);
nand U47852 (N_47852,N_46120,N_46641);
nor U47853 (N_47853,N_46171,N_46395);
xor U47854 (N_47854,N_46541,N_46080);
nand U47855 (N_47855,N_46352,N_46687);
and U47856 (N_47856,N_46039,N_46786);
nand U47857 (N_47857,N_46058,N_46825);
or U47858 (N_47858,N_46661,N_46251);
and U47859 (N_47859,N_46958,N_46737);
nor U47860 (N_47860,N_46819,N_46883);
xnor U47861 (N_47861,N_46133,N_46383);
nand U47862 (N_47862,N_46141,N_46749);
xor U47863 (N_47863,N_46320,N_46378);
nand U47864 (N_47864,N_46919,N_46378);
xnor U47865 (N_47865,N_46368,N_46427);
nor U47866 (N_47866,N_46941,N_46506);
xor U47867 (N_47867,N_46024,N_46471);
and U47868 (N_47868,N_46619,N_46096);
nand U47869 (N_47869,N_46500,N_46682);
nand U47870 (N_47870,N_46227,N_46109);
and U47871 (N_47871,N_46644,N_46760);
and U47872 (N_47872,N_46623,N_46252);
nor U47873 (N_47873,N_46961,N_46212);
or U47874 (N_47874,N_46894,N_46386);
xnor U47875 (N_47875,N_46329,N_46054);
xnor U47876 (N_47876,N_46231,N_46456);
and U47877 (N_47877,N_46317,N_46151);
nand U47878 (N_47878,N_46648,N_46690);
or U47879 (N_47879,N_46482,N_46820);
or U47880 (N_47880,N_46834,N_46106);
and U47881 (N_47881,N_46178,N_46320);
xor U47882 (N_47882,N_46879,N_46268);
or U47883 (N_47883,N_46189,N_46881);
or U47884 (N_47884,N_46628,N_46772);
nor U47885 (N_47885,N_46853,N_46167);
nand U47886 (N_47886,N_46542,N_46372);
or U47887 (N_47887,N_46769,N_46970);
or U47888 (N_47888,N_46092,N_46613);
or U47889 (N_47889,N_46440,N_46202);
nor U47890 (N_47890,N_46973,N_46802);
nand U47891 (N_47891,N_46980,N_46145);
xnor U47892 (N_47892,N_46968,N_46576);
xor U47893 (N_47893,N_46357,N_46532);
xnor U47894 (N_47894,N_46289,N_46233);
nor U47895 (N_47895,N_46076,N_46823);
nand U47896 (N_47896,N_46923,N_46619);
nor U47897 (N_47897,N_46887,N_46566);
and U47898 (N_47898,N_46135,N_46595);
nand U47899 (N_47899,N_46018,N_46516);
or U47900 (N_47900,N_46993,N_46306);
or U47901 (N_47901,N_46134,N_46119);
or U47902 (N_47902,N_46868,N_46546);
or U47903 (N_47903,N_46808,N_46317);
nand U47904 (N_47904,N_46946,N_46717);
nor U47905 (N_47905,N_46852,N_46484);
nand U47906 (N_47906,N_46325,N_46173);
xor U47907 (N_47907,N_46138,N_46287);
and U47908 (N_47908,N_46167,N_46897);
or U47909 (N_47909,N_46205,N_46025);
xnor U47910 (N_47910,N_46411,N_46684);
xor U47911 (N_47911,N_46028,N_46093);
xor U47912 (N_47912,N_46956,N_46492);
nand U47913 (N_47913,N_46073,N_46078);
nor U47914 (N_47914,N_46424,N_46470);
nor U47915 (N_47915,N_46483,N_46976);
xor U47916 (N_47916,N_46600,N_46336);
nor U47917 (N_47917,N_46428,N_46891);
and U47918 (N_47918,N_46344,N_46841);
and U47919 (N_47919,N_46981,N_46757);
and U47920 (N_47920,N_46724,N_46953);
nor U47921 (N_47921,N_46946,N_46281);
nor U47922 (N_47922,N_46906,N_46945);
nor U47923 (N_47923,N_46107,N_46358);
or U47924 (N_47924,N_46773,N_46671);
xor U47925 (N_47925,N_46561,N_46075);
and U47926 (N_47926,N_46365,N_46786);
or U47927 (N_47927,N_46065,N_46554);
nor U47928 (N_47928,N_46566,N_46662);
nand U47929 (N_47929,N_46740,N_46418);
nand U47930 (N_47930,N_46152,N_46608);
nor U47931 (N_47931,N_46416,N_46201);
nor U47932 (N_47932,N_46665,N_46354);
nand U47933 (N_47933,N_46638,N_46059);
and U47934 (N_47934,N_46753,N_46868);
nand U47935 (N_47935,N_46475,N_46743);
or U47936 (N_47936,N_46837,N_46096);
or U47937 (N_47937,N_46377,N_46601);
nand U47938 (N_47938,N_46030,N_46121);
nor U47939 (N_47939,N_46128,N_46148);
nor U47940 (N_47940,N_46574,N_46328);
xor U47941 (N_47941,N_46739,N_46408);
nand U47942 (N_47942,N_46346,N_46599);
nand U47943 (N_47943,N_46421,N_46768);
xnor U47944 (N_47944,N_46648,N_46229);
xor U47945 (N_47945,N_46719,N_46250);
nor U47946 (N_47946,N_46425,N_46575);
and U47947 (N_47947,N_46856,N_46028);
nor U47948 (N_47948,N_46185,N_46369);
nor U47949 (N_47949,N_46032,N_46500);
or U47950 (N_47950,N_46508,N_46226);
and U47951 (N_47951,N_46707,N_46886);
nor U47952 (N_47952,N_46004,N_46088);
or U47953 (N_47953,N_46130,N_46939);
and U47954 (N_47954,N_46477,N_46676);
or U47955 (N_47955,N_46704,N_46227);
nand U47956 (N_47956,N_46238,N_46644);
nand U47957 (N_47957,N_46006,N_46356);
xor U47958 (N_47958,N_46052,N_46277);
or U47959 (N_47959,N_46184,N_46271);
or U47960 (N_47960,N_46943,N_46435);
and U47961 (N_47961,N_46271,N_46461);
nand U47962 (N_47962,N_46820,N_46565);
or U47963 (N_47963,N_46401,N_46367);
nor U47964 (N_47964,N_46059,N_46726);
and U47965 (N_47965,N_46866,N_46984);
xor U47966 (N_47966,N_46699,N_46316);
xnor U47967 (N_47967,N_46595,N_46519);
nand U47968 (N_47968,N_46000,N_46497);
and U47969 (N_47969,N_46193,N_46272);
or U47970 (N_47970,N_46420,N_46234);
or U47971 (N_47971,N_46665,N_46634);
xor U47972 (N_47972,N_46008,N_46861);
or U47973 (N_47973,N_46858,N_46716);
xnor U47974 (N_47974,N_46682,N_46756);
nand U47975 (N_47975,N_46431,N_46222);
and U47976 (N_47976,N_46339,N_46074);
nand U47977 (N_47977,N_46661,N_46574);
xor U47978 (N_47978,N_46545,N_46975);
nand U47979 (N_47979,N_46452,N_46291);
or U47980 (N_47980,N_46649,N_46890);
nand U47981 (N_47981,N_46818,N_46826);
or U47982 (N_47982,N_46750,N_46110);
nor U47983 (N_47983,N_46996,N_46570);
nand U47984 (N_47984,N_46984,N_46499);
nand U47985 (N_47985,N_46904,N_46297);
nand U47986 (N_47986,N_46788,N_46705);
nand U47987 (N_47987,N_46821,N_46989);
and U47988 (N_47988,N_46622,N_46467);
nor U47989 (N_47989,N_46759,N_46767);
or U47990 (N_47990,N_46128,N_46399);
nor U47991 (N_47991,N_46165,N_46981);
and U47992 (N_47992,N_46753,N_46993);
nand U47993 (N_47993,N_46825,N_46464);
and U47994 (N_47994,N_46459,N_46929);
nor U47995 (N_47995,N_46274,N_46913);
nand U47996 (N_47996,N_46150,N_46006);
xor U47997 (N_47997,N_46232,N_46083);
and U47998 (N_47998,N_46117,N_46536);
or U47999 (N_47999,N_46419,N_46712);
or U48000 (N_48000,N_47539,N_47011);
and U48001 (N_48001,N_47739,N_47996);
and U48002 (N_48002,N_47917,N_47017);
or U48003 (N_48003,N_47741,N_47546);
and U48004 (N_48004,N_47212,N_47753);
xnor U48005 (N_48005,N_47640,N_47173);
or U48006 (N_48006,N_47157,N_47332);
nor U48007 (N_48007,N_47374,N_47163);
and U48008 (N_48008,N_47660,N_47644);
xnor U48009 (N_48009,N_47284,N_47036);
xor U48010 (N_48010,N_47750,N_47975);
nor U48011 (N_48011,N_47732,N_47665);
nand U48012 (N_48012,N_47902,N_47442);
xnor U48013 (N_48013,N_47675,N_47051);
xnor U48014 (N_48014,N_47662,N_47877);
xnor U48015 (N_48015,N_47179,N_47200);
nor U48016 (N_48016,N_47736,N_47758);
and U48017 (N_48017,N_47700,N_47420);
nand U48018 (N_48018,N_47116,N_47010);
or U48019 (N_48019,N_47103,N_47194);
xnor U48020 (N_48020,N_47446,N_47401);
nor U48021 (N_48021,N_47931,N_47386);
and U48022 (N_48022,N_47743,N_47467);
nand U48023 (N_48023,N_47137,N_47629);
or U48024 (N_48024,N_47564,N_47243);
or U48025 (N_48025,N_47319,N_47974);
xor U48026 (N_48026,N_47712,N_47087);
xor U48027 (N_48027,N_47953,N_47285);
nand U48028 (N_48028,N_47238,N_47027);
and U48029 (N_48029,N_47500,N_47257);
nand U48030 (N_48030,N_47561,N_47296);
nand U48031 (N_48031,N_47914,N_47574);
nand U48032 (N_48032,N_47612,N_47349);
xnor U48033 (N_48033,N_47936,N_47868);
or U48034 (N_48034,N_47961,N_47343);
xnor U48035 (N_48035,N_47844,N_47393);
xor U48036 (N_48036,N_47049,N_47493);
nand U48037 (N_48037,N_47714,N_47300);
xnor U48038 (N_48038,N_47715,N_47202);
or U48039 (N_48039,N_47253,N_47033);
nor U48040 (N_48040,N_47705,N_47636);
nand U48041 (N_48041,N_47192,N_47971);
and U48042 (N_48042,N_47853,N_47820);
nand U48043 (N_48043,N_47683,N_47759);
nand U48044 (N_48044,N_47836,N_47117);
and U48045 (N_48045,N_47874,N_47622);
xor U48046 (N_48046,N_47314,N_47217);
nand U48047 (N_48047,N_47389,N_47376);
nor U48048 (N_48048,N_47143,N_47638);
nor U48049 (N_48049,N_47102,N_47799);
or U48050 (N_48050,N_47663,N_47538);
nand U48051 (N_48051,N_47244,N_47692);
or U48052 (N_48052,N_47196,N_47141);
nand U48053 (N_48053,N_47220,N_47585);
or U48054 (N_48054,N_47248,N_47086);
nand U48055 (N_48055,N_47562,N_47998);
or U48056 (N_48056,N_47501,N_47726);
xor U48057 (N_48057,N_47068,N_47004);
and U48058 (N_48058,N_47568,N_47527);
nand U48059 (N_48059,N_47160,N_47135);
nand U48060 (N_48060,N_47092,N_47954);
and U48061 (N_48061,N_47579,N_47508);
xor U48062 (N_48062,N_47236,N_47709);
or U48063 (N_48063,N_47789,N_47066);
nand U48064 (N_48064,N_47361,N_47573);
nand U48065 (N_48065,N_47774,N_47840);
xnor U48066 (N_48066,N_47383,N_47843);
nor U48067 (N_48067,N_47762,N_47139);
nor U48068 (N_48068,N_47822,N_47333);
nor U48069 (N_48069,N_47536,N_47312);
nor U48070 (N_48070,N_47835,N_47551);
and U48071 (N_48071,N_47277,N_47183);
xnor U48072 (N_48072,N_47965,N_47364);
xnor U48073 (N_48073,N_47979,N_47384);
or U48074 (N_48074,N_47802,N_47819);
or U48075 (N_48075,N_47846,N_47666);
nand U48076 (N_48076,N_47474,N_47431);
or U48077 (N_48077,N_47825,N_47580);
or U48078 (N_48078,N_47528,N_47293);
nor U48079 (N_48079,N_47997,N_47289);
and U48080 (N_48080,N_47083,N_47871);
nor U48081 (N_48081,N_47186,N_47731);
or U48082 (N_48082,N_47462,N_47991);
xor U48083 (N_48083,N_47617,N_47341);
or U48084 (N_48084,N_47209,N_47335);
xor U48085 (N_48085,N_47667,N_47353);
nor U48086 (N_48086,N_47215,N_47969);
or U48087 (N_48087,N_47777,N_47441);
xnor U48088 (N_48088,N_47531,N_47311);
or U48089 (N_48089,N_47827,N_47413);
or U48090 (N_48090,N_47045,N_47447);
xor U48091 (N_48091,N_47618,N_47177);
and U48092 (N_48092,N_47266,N_47565);
or U48093 (N_48093,N_47856,N_47746);
or U48094 (N_48094,N_47903,N_47077);
nand U48095 (N_48095,N_47656,N_47694);
nor U48096 (N_48096,N_47064,N_47081);
and U48097 (N_48097,N_47717,N_47816);
nor U48098 (N_48098,N_47513,N_47752);
and U48099 (N_48099,N_47125,N_47698);
or U48100 (N_48100,N_47713,N_47166);
xnor U48101 (N_48101,N_47398,N_47309);
or U48102 (N_48102,N_47499,N_47873);
or U48103 (N_48103,N_47532,N_47023);
and U48104 (N_48104,N_47379,N_47515);
nand U48105 (N_48105,N_47788,N_47659);
xor U48106 (N_48106,N_47473,N_47338);
xor U48107 (N_48107,N_47616,N_47110);
or U48108 (N_48108,N_47688,N_47411);
nand U48109 (N_48109,N_47208,N_47778);
or U48110 (N_48110,N_47972,N_47911);
or U48111 (N_48111,N_47830,N_47938);
or U48112 (N_48112,N_47634,N_47610);
xnor U48113 (N_48113,N_47422,N_47523);
xor U48114 (N_48114,N_47794,N_47070);
nor U48115 (N_48115,N_47303,N_47892);
nor U48116 (N_48116,N_47188,N_47283);
nor U48117 (N_48117,N_47557,N_47860);
and U48118 (N_48118,N_47414,N_47721);
or U48119 (N_48119,N_47934,N_47614);
nand U48120 (N_48120,N_47121,N_47605);
or U48121 (N_48121,N_47124,N_47246);
nor U48122 (N_48122,N_47866,N_47833);
and U48123 (N_48123,N_47633,N_47405);
xor U48124 (N_48124,N_47182,N_47482);
nor U48125 (N_48125,N_47534,N_47581);
xnor U48126 (N_48126,N_47061,N_47589);
nor U48127 (N_48127,N_47609,N_47005);
and U48128 (N_48128,N_47304,N_47942);
xor U48129 (N_48129,N_47480,N_47432);
nor U48130 (N_48130,N_47985,N_47318);
xnor U48131 (N_48131,N_47242,N_47187);
xor U48132 (N_48132,N_47899,N_47809);
nand U48133 (N_48133,N_47520,N_47755);
and U48134 (N_48134,N_47488,N_47347);
or U48135 (N_48135,N_47195,N_47098);
xor U48136 (N_48136,N_47075,N_47922);
nor U48137 (N_48137,N_47987,N_47158);
nand U48138 (N_48138,N_47823,N_47362);
nand U48139 (N_48139,N_47403,N_47542);
nand U48140 (N_48140,N_47260,N_47904);
nand U48141 (N_48141,N_47572,N_47521);
or U48142 (N_48142,N_47711,N_47448);
xor U48143 (N_48143,N_47740,N_47486);
xor U48144 (N_48144,N_47438,N_47218);
or U48145 (N_48145,N_47535,N_47437);
nor U48146 (N_48146,N_47963,N_47716);
or U48147 (N_48147,N_47297,N_47131);
or U48148 (N_48148,N_47989,N_47783);
xnor U48149 (N_48149,N_47818,N_47230);
nor U48150 (N_48150,N_47278,N_47838);
nor U48151 (N_48151,N_47054,N_47735);
nand U48152 (N_48152,N_47653,N_47708);
and U48153 (N_48153,N_47136,N_47577);
xnor U48154 (N_48154,N_47962,N_47689);
xor U48155 (N_48155,N_47724,N_47354);
and U48156 (N_48156,N_47648,N_47639);
and U48157 (N_48157,N_47344,N_47901);
or U48158 (N_48158,N_47951,N_47334);
and U48159 (N_48159,N_47592,N_47995);
xnor U48160 (N_48160,N_47152,N_47408);
and U48161 (N_48161,N_47487,N_47053);
and U48162 (N_48162,N_47357,N_47745);
or U48163 (N_48163,N_47980,N_47146);
xnor U48164 (N_48164,N_47664,N_47854);
or U48165 (N_48165,N_47391,N_47138);
and U48166 (N_48166,N_47427,N_47258);
and U48167 (N_48167,N_47001,N_47367);
and U48168 (N_48168,N_47159,N_47031);
xnor U48169 (N_48169,N_47943,N_47720);
and U48170 (N_48170,N_47022,N_47810);
or U48171 (N_48171,N_47986,N_47878);
xnor U48172 (N_48172,N_47063,N_47233);
or U48173 (N_48173,N_47475,N_47882);
xnor U48174 (N_48174,N_47749,N_47381);
nand U48175 (N_48175,N_47894,N_47907);
xnor U48176 (N_48176,N_47576,N_47642);
nand U48177 (N_48177,N_47811,N_47702);
nor U48178 (N_48178,N_47030,N_47728);
and U48179 (N_48179,N_47525,N_47461);
or U48180 (N_48180,N_47505,N_47029);
nand U48181 (N_48181,N_47180,N_47926);
xor U48182 (N_48182,N_47041,N_47071);
nor U48183 (N_48183,N_47729,N_47418);
and U48184 (N_48184,N_47028,N_47178);
nor U48185 (N_48185,N_47540,N_47590);
or U48186 (N_48186,N_47817,N_47142);
nand U48187 (N_48187,N_47324,N_47404);
or U48188 (N_48188,N_47781,N_47761);
nor U48189 (N_48189,N_47869,N_47803);
or U48190 (N_48190,N_47673,N_47945);
and U48191 (N_48191,N_47958,N_47394);
or U48192 (N_48192,N_47197,N_47128);
nor U48193 (N_48193,N_47983,N_47796);
and U48194 (N_48194,N_47966,N_47647);
nor U48195 (N_48195,N_47625,N_47423);
and U48196 (N_48196,N_47425,N_47925);
nand U48197 (N_48197,N_47993,N_47582);
and U48198 (N_48198,N_47459,N_47744);
xnor U48199 (N_48199,N_47575,N_47466);
nand U48200 (N_48200,N_47876,N_47676);
xnor U48201 (N_48201,N_47134,N_47043);
nand U48202 (N_48202,N_47831,N_47804);
xnor U48203 (N_48203,N_47497,N_47250);
xnor U48204 (N_48204,N_47380,N_47850);
nand U48205 (N_48205,N_47725,N_47078);
nand U48206 (N_48206,N_47603,N_47631);
nor U48207 (N_48207,N_47275,N_47757);
xnor U48208 (N_48208,N_47602,N_47537);
xnor U48209 (N_48209,N_47992,N_47814);
or U48210 (N_48210,N_47321,N_47009);
nor U48211 (N_48211,N_47057,N_47928);
and U48212 (N_48212,N_47560,N_47775);
or U48213 (N_48213,N_47176,N_47512);
and U48214 (N_48214,N_47368,N_47346);
or U48215 (N_48215,N_47214,N_47994);
and U48216 (N_48216,N_47913,N_47751);
nand U48217 (N_48217,N_47415,N_47108);
nand U48218 (N_48218,N_47637,N_47893);
xnor U48219 (N_48219,N_47271,N_47879);
xor U48220 (N_48220,N_47905,N_47235);
nor U48221 (N_48221,N_47039,N_47859);
nor U48222 (N_48222,N_47396,N_47498);
or U48223 (N_48223,N_47485,N_47140);
xor U48224 (N_48224,N_47685,N_47923);
and U48225 (N_48225,N_47090,N_47681);
nand U48226 (N_48226,N_47872,N_47672);
nor U48227 (N_48227,N_47455,N_47211);
and U48228 (N_48228,N_47088,N_47037);
and U48229 (N_48229,N_47988,N_47699);
and U48230 (N_48230,N_47084,N_47052);
nand U48231 (N_48231,N_47848,N_47503);
and U48232 (N_48232,N_47012,N_47331);
or U48233 (N_48233,N_47679,N_47502);
xnor U48234 (N_48234,N_47205,N_47748);
nor U48235 (N_48235,N_47530,N_47395);
nand U48236 (N_48236,N_47600,N_47924);
and U48237 (N_48237,N_47552,N_47571);
xor U48238 (N_48238,N_47032,N_47481);
nor U48239 (N_48239,N_47896,N_47276);
nand U48240 (N_48240,N_47419,N_47604);
and U48241 (N_48241,N_47870,N_47933);
nor U48242 (N_48242,N_47337,N_47327);
and U48243 (N_48243,N_47272,N_47147);
nor U48244 (N_48244,N_47627,N_47780);
nor U48245 (N_48245,N_47766,N_47655);
or U48246 (N_48246,N_47787,N_47399);
nand U48247 (N_48247,N_47517,N_47548);
nand U48248 (N_48248,N_47950,N_47821);
nand U48249 (N_48249,N_47932,N_47981);
or U48250 (N_48250,N_47454,N_47308);
nand U48251 (N_48251,N_47509,N_47430);
nor U48252 (N_48252,N_47013,N_47252);
nand U48253 (N_48253,N_47255,N_47007);
xnor U48254 (N_48254,N_47067,N_47615);
nor U48255 (N_48255,N_47623,N_47566);
nor U48256 (N_48256,N_47130,N_47458);
nand U48257 (N_48257,N_47658,N_47939);
nor U48258 (N_48258,N_47489,N_47378);
and U48259 (N_48259,N_47545,N_47185);
and U48260 (N_48260,N_47014,N_47927);
nor U48261 (N_48261,N_47015,N_47153);
nand U48262 (N_48262,N_47829,N_47421);
nor U48263 (N_48263,N_47885,N_47583);
nand U48264 (N_48264,N_47649,N_47767);
nand U48265 (N_48265,N_47101,N_47674);
xor U48266 (N_48266,N_47624,N_47668);
xnor U48267 (N_48267,N_47718,N_47201);
and U48268 (N_48268,N_47567,N_47169);
nor U48269 (N_48269,N_47516,N_47691);
nor U48270 (N_48270,N_47112,N_47231);
nand U48271 (N_48271,N_47558,N_47443);
nor U48272 (N_48272,N_47145,N_47506);
and U48273 (N_48273,N_47707,N_47865);
nor U48274 (N_48274,N_47317,N_47940);
nand U48275 (N_48275,N_47237,N_47193);
nand U48276 (N_48276,N_47678,N_47686);
xor U48277 (N_48277,N_47114,N_47198);
xnor U48278 (N_48278,N_47909,N_47062);
xor U48279 (N_48279,N_47722,N_47792);
nor U48280 (N_48280,N_47042,N_47358);
xor U48281 (N_48281,N_47834,N_47956);
and U48282 (N_48282,N_47510,N_47946);
nor U48283 (N_48283,N_47861,N_47452);
xnor U48284 (N_48284,N_47955,N_47719);
and U48285 (N_48285,N_47213,N_47165);
or U48286 (N_48286,N_47937,N_47120);
or U48287 (N_48287,N_47330,N_47670);
nor U48288 (N_48288,N_47400,N_47111);
nor U48289 (N_48289,N_47779,N_47898);
or U48290 (N_48290,N_47279,N_47360);
xnor U48291 (N_48291,N_47710,N_47072);
xor U48292 (N_48292,N_47598,N_47224);
xnor U48293 (N_48293,N_47763,N_47059);
xnor U48294 (N_48294,N_47687,N_47684);
xor U48295 (N_48295,N_47091,N_47294);
nor U48296 (N_48296,N_47800,N_47181);
nand U48297 (N_48297,N_47407,N_47654);
nand U48298 (N_48298,N_47204,N_47265);
nor U48299 (N_48299,N_47606,N_47305);
nand U48300 (N_48300,N_47490,N_47234);
xnor U48301 (N_48301,N_47232,N_47106);
nand U48302 (N_48302,N_47620,N_47249);
nor U48303 (N_48303,N_47786,N_47984);
and U48304 (N_48304,N_47864,N_47221);
or U48305 (N_48305,N_47329,N_47587);
or U48306 (N_48306,N_47097,N_47776);
nor U48307 (N_48307,N_47782,N_47897);
nand U48308 (N_48308,N_47760,N_47857);
or U48309 (N_48309,N_47290,N_47941);
xor U48310 (N_48310,N_47203,N_47301);
nor U48311 (N_48311,N_47174,N_47348);
or U48312 (N_48312,N_47171,N_47274);
nand U48313 (N_48313,N_47269,N_47514);
nor U48314 (N_48314,N_47471,N_47340);
xor U48315 (N_48315,N_47356,N_47929);
xnor U48316 (N_48316,N_47553,N_47003);
and U48317 (N_48317,N_47578,N_47047);
nand U48318 (N_48318,N_47880,N_47434);
or U48319 (N_48319,N_47967,N_47397);
xor U48320 (N_48320,N_47190,N_47251);
or U48321 (N_48321,N_47315,N_47154);
nand U48322 (N_48322,N_47547,N_47613);
xnor U48323 (N_48323,N_47172,N_47690);
and U48324 (N_48324,N_47162,N_47533);
nor U48325 (N_48325,N_47559,N_47210);
and U48326 (N_48326,N_47355,N_47323);
nand U48327 (N_48327,N_47025,N_47263);
xnor U48328 (N_48328,N_47366,N_47020);
xor U48329 (N_48329,N_47867,N_47842);
nand U48330 (N_48330,N_47504,N_47417);
nor U48331 (N_48331,N_47477,N_47089);
nor U48332 (N_48332,N_47082,N_47646);
or U48333 (N_48333,N_47118,N_47964);
and U48334 (N_48334,N_47035,N_47282);
nor U48335 (N_48335,N_47433,N_47588);
xor U48336 (N_48336,N_47264,N_47768);
nor U48337 (N_48337,N_47550,N_47256);
and U48338 (N_48338,N_47021,N_47149);
or U48339 (N_48339,N_47526,N_47852);
nor U48340 (N_48340,N_47206,N_47365);
nor U48341 (N_48341,N_47930,N_47556);
or U48342 (N_48342,N_47915,N_47921);
nor U48343 (N_48343,N_47677,N_47286);
nand U48344 (N_48344,N_47104,N_47370);
and U48345 (N_48345,N_47507,N_47730);
and U48346 (N_48346,N_47669,N_47635);
xor U48347 (N_48347,N_47544,N_47388);
xnor U48348 (N_48348,N_47093,N_47770);
nor U48349 (N_48349,N_47463,N_47858);
nand U48350 (N_48350,N_47597,N_47591);
xnor U48351 (N_48351,N_47948,N_47109);
and U48352 (N_48352,N_47935,N_47144);
nand U48353 (N_48353,N_47630,N_47148);
nor U48354 (N_48354,N_47765,N_47990);
nand U48355 (N_48355,N_47040,N_47392);
and U48356 (N_48356,N_47280,N_47738);
nand U48357 (N_48357,N_47977,N_47695);
or U48358 (N_48358,N_47460,N_47245);
and U48359 (N_48359,N_47436,N_47608);
and U48360 (N_48360,N_47465,N_47737);
xnor U48361 (N_48361,N_47444,N_47495);
nand U48362 (N_48362,N_47065,N_47519);
or U48363 (N_48363,N_47387,N_47326);
and U48364 (N_48364,N_47594,N_47034);
or U48365 (N_48365,N_47322,N_47626);
nor U48366 (N_48366,N_47416,N_47435);
and U48367 (N_48367,N_47957,N_47259);
nand U48368 (N_48368,N_47080,N_47292);
nand U48369 (N_48369,N_47887,N_47801);
and U48370 (N_48370,N_47601,N_47000);
nor U48371 (N_48371,N_47795,N_47970);
nand U48372 (N_48372,N_47073,N_47813);
nand U48373 (N_48373,N_47484,N_47302);
nor U48374 (N_48374,N_47107,N_47076);
or U48375 (N_48375,N_47372,N_47268);
nor U48376 (N_48376,N_47815,N_47164);
or U48377 (N_48377,N_47628,N_47976);
and U48378 (N_48378,N_47156,N_47476);
nor U48379 (N_48379,N_47797,N_47772);
or U48380 (N_48380,N_47704,N_47593);
or U48381 (N_48381,N_47468,N_47450);
and U48382 (N_48382,N_47095,N_47056);
and U48383 (N_48383,N_47273,N_47478);
nor U48384 (N_48384,N_47069,N_47784);
nor U48385 (N_48385,N_47807,N_47906);
xor U48386 (N_48386,N_47189,N_47227);
or U48387 (N_48387,N_47024,N_47491);
nand U48388 (N_48388,N_47541,N_47058);
or U48389 (N_48389,N_47225,N_47949);
or U48390 (N_48390,N_47440,N_47886);
xnor U48391 (N_48391,N_47390,N_47464);
nand U48392 (N_48392,N_47918,N_47409);
nor U48393 (N_48393,N_47168,N_47944);
xnor U48394 (N_48394,N_47701,N_47191);
and U48395 (N_48395,N_47661,N_47773);
or U48396 (N_48396,N_47320,N_47798);
or U48397 (N_48397,N_47596,N_47469);
nor U48398 (N_48398,N_47960,N_47790);
and U48399 (N_48399,N_47920,N_47999);
nand U48400 (N_48400,N_47947,N_47808);
xor U48401 (N_48401,N_47518,N_47096);
or U48402 (N_48402,N_47207,N_47891);
and U48403 (N_48403,N_47492,N_47428);
xnor U48404 (N_48404,N_47734,N_47254);
or U48405 (N_48405,N_47229,N_47044);
xnor U48406 (N_48406,N_47849,N_47241);
and U48407 (N_48407,N_47599,N_47563);
or U48408 (N_48408,N_47155,N_47170);
nand U48409 (N_48409,N_47050,N_47641);
nand U48410 (N_48410,N_47919,N_47055);
and U48411 (N_48411,N_47115,N_47038);
xnor U48412 (N_48412,N_47262,N_47150);
nor U48413 (N_48413,N_47298,N_47845);
or U48414 (N_48414,N_47412,N_47805);
nor U48415 (N_48415,N_47456,N_47875);
or U48416 (N_48416,N_47046,N_47288);
nand U48417 (N_48417,N_47270,N_47339);
nand U48418 (N_48418,N_47727,N_47912);
xnor U48419 (N_48419,N_47359,N_47812);
nand U48420 (N_48420,N_47832,N_47048);
xnor U48421 (N_48421,N_47385,N_47611);
nor U48422 (N_48422,N_47342,N_47764);
nand U48423 (N_48423,N_47890,N_47099);
xnor U48424 (N_48424,N_47793,N_47828);
nor U48425 (N_48425,N_47851,N_47222);
and U48426 (N_48426,N_47806,N_47281);
xor U48427 (N_48427,N_47369,N_47494);
nor U48428 (N_48428,N_47978,N_47228);
xor U48429 (N_48429,N_47855,N_47016);
nor U48430 (N_48430,N_47952,N_47621);
nor U48431 (N_48431,N_47426,N_47769);
and U48432 (N_48432,N_47439,N_47472);
xnor U48433 (N_48433,N_47643,N_47313);
nand U48434 (N_48434,N_47008,N_47837);
xnor U48435 (N_48435,N_47184,N_47549);
and U48436 (N_48436,N_47129,N_47723);
nor U48437 (N_48437,N_47240,N_47883);
or U48438 (N_48438,N_47652,N_47451);
or U48439 (N_48439,N_47595,N_47375);
nand U48440 (N_48440,N_47570,N_47026);
and U48441 (N_48441,N_47429,N_47316);
and U48442 (N_48442,N_47671,N_47307);
xnor U48443 (N_48443,N_47019,N_47167);
xnor U48444 (N_48444,N_47406,N_47350);
xnor U48445 (N_48445,N_47982,N_47345);
xor U48446 (N_48446,N_47771,N_47453);
or U48447 (N_48447,N_47002,N_47151);
or U48448 (N_48448,N_47100,N_47733);
nand U48449 (N_48449,N_47824,N_47457);
nand U48450 (N_48450,N_47126,N_47410);
nor U48451 (N_48451,N_47569,N_47085);
nor U48452 (N_48452,N_47863,N_47529);
and U48453 (N_48453,N_47584,N_47133);
xnor U48454 (N_48454,N_47373,N_47402);
and U48455 (N_48455,N_47884,N_47650);
nand U48456 (N_48456,N_47619,N_47449);
nand U48457 (N_48457,N_47219,N_47123);
or U48458 (N_48458,N_47839,N_47094);
nor U48459 (N_48459,N_47959,N_47445);
nand U48460 (N_48460,N_47554,N_47881);
or U48461 (N_48461,N_47119,N_47239);
or U48462 (N_48462,N_47363,N_47889);
xnor U48463 (N_48463,N_47522,N_47306);
nor U48464 (N_48464,N_47555,N_47074);
or U48465 (N_48465,N_47291,N_47295);
xnor U48466 (N_48466,N_47199,N_47632);
or U48467 (N_48467,N_47261,N_47696);
xnor U48468 (N_48468,N_47791,N_47122);
and U48469 (N_48469,N_47371,N_47352);
nand U48470 (N_48470,N_47747,N_47113);
nor U48471 (N_48471,N_47483,N_47018);
and U48472 (N_48472,N_47586,N_47847);
xor U48473 (N_48473,N_47006,N_47299);
or U48474 (N_48474,N_47310,N_47132);
nor U48475 (N_48475,N_47841,N_47908);
or U48476 (N_48476,N_47382,N_47226);
or U48477 (N_48477,N_47223,N_47161);
or U48478 (N_48478,N_47607,N_47336);
nand U48479 (N_48479,N_47862,N_47826);
and U48480 (N_48480,N_47785,N_47377);
and U48481 (N_48481,N_47703,N_47524);
and U48482 (N_48482,N_47693,N_47754);
and U48483 (N_48483,N_47756,N_47175);
nand U48484 (N_48484,N_47697,N_47916);
nand U48485 (N_48485,N_47680,N_47127);
nor U48486 (N_48486,N_47543,N_47895);
or U48487 (N_48487,N_47470,N_47105);
or U48488 (N_48488,N_47496,N_47968);
or U48489 (N_48489,N_47351,N_47328);
or U48490 (N_48490,N_47424,N_47742);
or U48491 (N_48491,N_47910,N_47325);
nand U48492 (N_48492,N_47973,N_47706);
nor U48493 (N_48493,N_47216,N_47267);
or U48494 (N_48494,N_47651,N_47247);
nor U48495 (N_48495,N_47682,N_47287);
and U48496 (N_48496,N_47060,N_47479);
nor U48497 (N_48497,N_47888,N_47657);
or U48498 (N_48498,N_47645,N_47900);
and U48499 (N_48499,N_47079,N_47511);
or U48500 (N_48500,N_47298,N_47911);
xnor U48501 (N_48501,N_47201,N_47772);
or U48502 (N_48502,N_47688,N_47818);
xnor U48503 (N_48503,N_47527,N_47287);
and U48504 (N_48504,N_47785,N_47026);
xnor U48505 (N_48505,N_47597,N_47427);
nor U48506 (N_48506,N_47400,N_47262);
nor U48507 (N_48507,N_47996,N_47904);
xor U48508 (N_48508,N_47007,N_47461);
nor U48509 (N_48509,N_47094,N_47446);
xnor U48510 (N_48510,N_47187,N_47557);
nor U48511 (N_48511,N_47564,N_47780);
and U48512 (N_48512,N_47191,N_47016);
nor U48513 (N_48513,N_47767,N_47953);
and U48514 (N_48514,N_47188,N_47126);
or U48515 (N_48515,N_47073,N_47689);
or U48516 (N_48516,N_47785,N_47703);
nor U48517 (N_48517,N_47591,N_47701);
and U48518 (N_48518,N_47022,N_47905);
and U48519 (N_48519,N_47927,N_47215);
nand U48520 (N_48520,N_47258,N_47535);
xor U48521 (N_48521,N_47509,N_47343);
nand U48522 (N_48522,N_47106,N_47493);
or U48523 (N_48523,N_47389,N_47374);
nor U48524 (N_48524,N_47726,N_47654);
nor U48525 (N_48525,N_47010,N_47527);
nor U48526 (N_48526,N_47952,N_47467);
or U48527 (N_48527,N_47842,N_47902);
or U48528 (N_48528,N_47044,N_47547);
and U48529 (N_48529,N_47139,N_47553);
nor U48530 (N_48530,N_47149,N_47257);
and U48531 (N_48531,N_47078,N_47251);
nor U48532 (N_48532,N_47199,N_47250);
and U48533 (N_48533,N_47532,N_47988);
xnor U48534 (N_48534,N_47528,N_47058);
nor U48535 (N_48535,N_47786,N_47774);
nand U48536 (N_48536,N_47261,N_47330);
xnor U48537 (N_48537,N_47532,N_47370);
and U48538 (N_48538,N_47798,N_47489);
or U48539 (N_48539,N_47478,N_47566);
nor U48540 (N_48540,N_47912,N_47963);
and U48541 (N_48541,N_47424,N_47939);
xor U48542 (N_48542,N_47928,N_47160);
nor U48543 (N_48543,N_47891,N_47572);
xor U48544 (N_48544,N_47165,N_47125);
nand U48545 (N_48545,N_47572,N_47719);
nor U48546 (N_48546,N_47801,N_47704);
and U48547 (N_48547,N_47247,N_47675);
xor U48548 (N_48548,N_47243,N_47234);
nand U48549 (N_48549,N_47425,N_47996);
nand U48550 (N_48550,N_47991,N_47803);
xor U48551 (N_48551,N_47511,N_47892);
or U48552 (N_48552,N_47383,N_47822);
xnor U48553 (N_48553,N_47314,N_47275);
nor U48554 (N_48554,N_47278,N_47579);
nand U48555 (N_48555,N_47172,N_47728);
and U48556 (N_48556,N_47040,N_47847);
nor U48557 (N_48557,N_47347,N_47441);
xor U48558 (N_48558,N_47534,N_47397);
nor U48559 (N_48559,N_47803,N_47197);
or U48560 (N_48560,N_47097,N_47712);
or U48561 (N_48561,N_47912,N_47555);
nand U48562 (N_48562,N_47231,N_47440);
nor U48563 (N_48563,N_47176,N_47449);
or U48564 (N_48564,N_47216,N_47812);
or U48565 (N_48565,N_47499,N_47033);
or U48566 (N_48566,N_47448,N_47160);
nand U48567 (N_48567,N_47131,N_47601);
nor U48568 (N_48568,N_47121,N_47535);
and U48569 (N_48569,N_47051,N_47933);
nand U48570 (N_48570,N_47551,N_47862);
and U48571 (N_48571,N_47826,N_47175);
xor U48572 (N_48572,N_47452,N_47512);
or U48573 (N_48573,N_47925,N_47569);
and U48574 (N_48574,N_47660,N_47634);
nand U48575 (N_48575,N_47507,N_47950);
or U48576 (N_48576,N_47791,N_47185);
nor U48577 (N_48577,N_47364,N_47803);
xor U48578 (N_48578,N_47347,N_47214);
xnor U48579 (N_48579,N_47918,N_47889);
xor U48580 (N_48580,N_47319,N_47833);
and U48581 (N_48581,N_47516,N_47803);
xnor U48582 (N_48582,N_47939,N_47820);
nand U48583 (N_48583,N_47068,N_47322);
nand U48584 (N_48584,N_47563,N_47488);
nand U48585 (N_48585,N_47383,N_47066);
nand U48586 (N_48586,N_47283,N_47539);
xor U48587 (N_48587,N_47269,N_47841);
or U48588 (N_48588,N_47826,N_47165);
nor U48589 (N_48589,N_47009,N_47230);
nand U48590 (N_48590,N_47451,N_47865);
xor U48591 (N_48591,N_47599,N_47190);
xor U48592 (N_48592,N_47621,N_47628);
and U48593 (N_48593,N_47055,N_47468);
nand U48594 (N_48594,N_47756,N_47097);
nand U48595 (N_48595,N_47313,N_47480);
nand U48596 (N_48596,N_47302,N_47332);
xor U48597 (N_48597,N_47400,N_47018);
and U48598 (N_48598,N_47375,N_47573);
nor U48599 (N_48599,N_47345,N_47186);
nor U48600 (N_48600,N_47712,N_47698);
nor U48601 (N_48601,N_47192,N_47801);
xor U48602 (N_48602,N_47128,N_47514);
nor U48603 (N_48603,N_47916,N_47726);
and U48604 (N_48604,N_47935,N_47392);
nand U48605 (N_48605,N_47169,N_47236);
nand U48606 (N_48606,N_47245,N_47801);
xnor U48607 (N_48607,N_47929,N_47945);
or U48608 (N_48608,N_47112,N_47522);
nand U48609 (N_48609,N_47866,N_47669);
or U48610 (N_48610,N_47901,N_47371);
nand U48611 (N_48611,N_47067,N_47315);
nand U48612 (N_48612,N_47715,N_47548);
or U48613 (N_48613,N_47372,N_47298);
nor U48614 (N_48614,N_47997,N_47176);
xnor U48615 (N_48615,N_47117,N_47371);
xnor U48616 (N_48616,N_47038,N_47940);
nand U48617 (N_48617,N_47163,N_47894);
and U48618 (N_48618,N_47010,N_47977);
nand U48619 (N_48619,N_47232,N_47035);
nand U48620 (N_48620,N_47560,N_47331);
or U48621 (N_48621,N_47177,N_47315);
and U48622 (N_48622,N_47251,N_47658);
or U48623 (N_48623,N_47078,N_47762);
xor U48624 (N_48624,N_47368,N_47606);
and U48625 (N_48625,N_47737,N_47305);
and U48626 (N_48626,N_47731,N_47542);
and U48627 (N_48627,N_47657,N_47569);
xor U48628 (N_48628,N_47428,N_47238);
or U48629 (N_48629,N_47981,N_47946);
xnor U48630 (N_48630,N_47532,N_47903);
or U48631 (N_48631,N_47539,N_47715);
nor U48632 (N_48632,N_47947,N_47936);
nand U48633 (N_48633,N_47701,N_47755);
and U48634 (N_48634,N_47932,N_47046);
nor U48635 (N_48635,N_47471,N_47798);
nor U48636 (N_48636,N_47315,N_47443);
nand U48637 (N_48637,N_47309,N_47996);
or U48638 (N_48638,N_47175,N_47067);
nand U48639 (N_48639,N_47589,N_47400);
nor U48640 (N_48640,N_47668,N_47951);
nand U48641 (N_48641,N_47066,N_47631);
and U48642 (N_48642,N_47336,N_47816);
xnor U48643 (N_48643,N_47349,N_47476);
and U48644 (N_48644,N_47406,N_47683);
and U48645 (N_48645,N_47249,N_47723);
nand U48646 (N_48646,N_47786,N_47409);
nor U48647 (N_48647,N_47617,N_47970);
nand U48648 (N_48648,N_47225,N_47799);
xor U48649 (N_48649,N_47801,N_47696);
and U48650 (N_48650,N_47699,N_47636);
nand U48651 (N_48651,N_47521,N_47080);
nand U48652 (N_48652,N_47392,N_47498);
and U48653 (N_48653,N_47486,N_47224);
xor U48654 (N_48654,N_47687,N_47612);
nand U48655 (N_48655,N_47747,N_47930);
xnor U48656 (N_48656,N_47517,N_47268);
nor U48657 (N_48657,N_47060,N_47004);
and U48658 (N_48658,N_47045,N_47510);
nand U48659 (N_48659,N_47753,N_47372);
nand U48660 (N_48660,N_47723,N_47721);
nor U48661 (N_48661,N_47348,N_47661);
or U48662 (N_48662,N_47756,N_47170);
or U48663 (N_48663,N_47231,N_47618);
nand U48664 (N_48664,N_47978,N_47910);
and U48665 (N_48665,N_47376,N_47417);
xnor U48666 (N_48666,N_47217,N_47850);
and U48667 (N_48667,N_47389,N_47583);
or U48668 (N_48668,N_47556,N_47017);
nor U48669 (N_48669,N_47719,N_47588);
and U48670 (N_48670,N_47866,N_47432);
nand U48671 (N_48671,N_47883,N_47915);
or U48672 (N_48672,N_47303,N_47799);
or U48673 (N_48673,N_47636,N_47113);
or U48674 (N_48674,N_47007,N_47039);
nand U48675 (N_48675,N_47362,N_47311);
xnor U48676 (N_48676,N_47651,N_47675);
nor U48677 (N_48677,N_47274,N_47348);
and U48678 (N_48678,N_47868,N_47254);
nand U48679 (N_48679,N_47615,N_47095);
nor U48680 (N_48680,N_47523,N_47357);
nor U48681 (N_48681,N_47681,N_47088);
xnor U48682 (N_48682,N_47488,N_47870);
or U48683 (N_48683,N_47212,N_47861);
nand U48684 (N_48684,N_47484,N_47941);
xor U48685 (N_48685,N_47895,N_47002);
or U48686 (N_48686,N_47084,N_47483);
xor U48687 (N_48687,N_47291,N_47093);
or U48688 (N_48688,N_47727,N_47665);
nand U48689 (N_48689,N_47319,N_47560);
nor U48690 (N_48690,N_47140,N_47634);
and U48691 (N_48691,N_47959,N_47882);
and U48692 (N_48692,N_47873,N_47681);
and U48693 (N_48693,N_47565,N_47388);
nand U48694 (N_48694,N_47148,N_47887);
and U48695 (N_48695,N_47977,N_47997);
nand U48696 (N_48696,N_47721,N_47317);
nor U48697 (N_48697,N_47061,N_47887);
xor U48698 (N_48698,N_47242,N_47778);
and U48699 (N_48699,N_47892,N_47552);
or U48700 (N_48700,N_47477,N_47605);
and U48701 (N_48701,N_47906,N_47791);
nor U48702 (N_48702,N_47234,N_47918);
nor U48703 (N_48703,N_47409,N_47248);
and U48704 (N_48704,N_47054,N_47544);
xor U48705 (N_48705,N_47553,N_47615);
and U48706 (N_48706,N_47625,N_47951);
and U48707 (N_48707,N_47847,N_47898);
nor U48708 (N_48708,N_47135,N_47921);
nor U48709 (N_48709,N_47065,N_47118);
or U48710 (N_48710,N_47384,N_47459);
nand U48711 (N_48711,N_47547,N_47641);
nand U48712 (N_48712,N_47904,N_47668);
xnor U48713 (N_48713,N_47344,N_47740);
xor U48714 (N_48714,N_47436,N_47772);
and U48715 (N_48715,N_47238,N_47914);
xnor U48716 (N_48716,N_47025,N_47254);
or U48717 (N_48717,N_47210,N_47973);
and U48718 (N_48718,N_47149,N_47920);
and U48719 (N_48719,N_47684,N_47597);
xor U48720 (N_48720,N_47851,N_47874);
nand U48721 (N_48721,N_47018,N_47728);
nand U48722 (N_48722,N_47790,N_47447);
and U48723 (N_48723,N_47920,N_47840);
xnor U48724 (N_48724,N_47789,N_47517);
or U48725 (N_48725,N_47480,N_47739);
xor U48726 (N_48726,N_47590,N_47716);
and U48727 (N_48727,N_47645,N_47624);
and U48728 (N_48728,N_47140,N_47133);
or U48729 (N_48729,N_47066,N_47343);
nand U48730 (N_48730,N_47289,N_47442);
nor U48731 (N_48731,N_47291,N_47655);
nand U48732 (N_48732,N_47953,N_47188);
or U48733 (N_48733,N_47989,N_47430);
nor U48734 (N_48734,N_47653,N_47039);
nor U48735 (N_48735,N_47511,N_47992);
xor U48736 (N_48736,N_47915,N_47820);
nand U48737 (N_48737,N_47282,N_47084);
nor U48738 (N_48738,N_47189,N_47241);
or U48739 (N_48739,N_47408,N_47610);
xnor U48740 (N_48740,N_47234,N_47233);
nand U48741 (N_48741,N_47358,N_47212);
xnor U48742 (N_48742,N_47087,N_47996);
and U48743 (N_48743,N_47985,N_47876);
nor U48744 (N_48744,N_47766,N_47449);
nand U48745 (N_48745,N_47606,N_47895);
nor U48746 (N_48746,N_47036,N_47317);
nor U48747 (N_48747,N_47281,N_47348);
and U48748 (N_48748,N_47480,N_47695);
and U48749 (N_48749,N_47001,N_47889);
nor U48750 (N_48750,N_47288,N_47159);
nor U48751 (N_48751,N_47552,N_47345);
and U48752 (N_48752,N_47016,N_47620);
nor U48753 (N_48753,N_47841,N_47322);
nor U48754 (N_48754,N_47852,N_47407);
nand U48755 (N_48755,N_47025,N_47293);
xnor U48756 (N_48756,N_47249,N_47882);
nand U48757 (N_48757,N_47972,N_47103);
and U48758 (N_48758,N_47203,N_47123);
xor U48759 (N_48759,N_47857,N_47002);
xor U48760 (N_48760,N_47557,N_47992);
nand U48761 (N_48761,N_47390,N_47773);
nand U48762 (N_48762,N_47426,N_47433);
xor U48763 (N_48763,N_47359,N_47483);
or U48764 (N_48764,N_47764,N_47347);
nor U48765 (N_48765,N_47694,N_47010);
xor U48766 (N_48766,N_47986,N_47868);
or U48767 (N_48767,N_47759,N_47168);
or U48768 (N_48768,N_47372,N_47754);
nor U48769 (N_48769,N_47089,N_47733);
nand U48770 (N_48770,N_47847,N_47987);
nand U48771 (N_48771,N_47468,N_47041);
xnor U48772 (N_48772,N_47158,N_47619);
and U48773 (N_48773,N_47325,N_47435);
or U48774 (N_48774,N_47660,N_47889);
or U48775 (N_48775,N_47626,N_47337);
xnor U48776 (N_48776,N_47836,N_47590);
xnor U48777 (N_48777,N_47796,N_47818);
nand U48778 (N_48778,N_47564,N_47127);
nand U48779 (N_48779,N_47142,N_47643);
nand U48780 (N_48780,N_47067,N_47540);
nor U48781 (N_48781,N_47911,N_47699);
nor U48782 (N_48782,N_47484,N_47963);
or U48783 (N_48783,N_47285,N_47472);
nand U48784 (N_48784,N_47606,N_47658);
xor U48785 (N_48785,N_47262,N_47529);
nand U48786 (N_48786,N_47800,N_47440);
or U48787 (N_48787,N_47032,N_47235);
or U48788 (N_48788,N_47866,N_47099);
or U48789 (N_48789,N_47843,N_47627);
and U48790 (N_48790,N_47535,N_47069);
xor U48791 (N_48791,N_47843,N_47345);
or U48792 (N_48792,N_47007,N_47497);
xnor U48793 (N_48793,N_47647,N_47189);
nor U48794 (N_48794,N_47057,N_47251);
nor U48795 (N_48795,N_47978,N_47621);
xor U48796 (N_48796,N_47104,N_47928);
and U48797 (N_48797,N_47512,N_47433);
nand U48798 (N_48798,N_47599,N_47582);
nor U48799 (N_48799,N_47600,N_47849);
and U48800 (N_48800,N_47159,N_47008);
nor U48801 (N_48801,N_47627,N_47933);
nor U48802 (N_48802,N_47366,N_47614);
nand U48803 (N_48803,N_47911,N_47599);
nor U48804 (N_48804,N_47745,N_47478);
xor U48805 (N_48805,N_47832,N_47031);
or U48806 (N_48806,N_47736,N_47821);
and U48807 (N_48807,N_47555,N_47099);
xor U48808 (N_48808,N_47998,N_47725);
or U48809 (N_48809,N_47168,N_47634);
nand U48810 (N_48810,N_47998,N_47820);
nor U48811 (N_48811,N_47625,N_47101);
and U48812 (N_48812,N_47653,N_47783);
xnor U48813 (N_48813,N_47023,N_47045);
and U48814 (N_48814,N_47845,N_47472);
or U48815 (N_48815,N_47557,N_47321);
nor U48816 (N_48816,N_47355,N_47615);
and U48817 (N_48817,N_47216,N_47927);
and U48818 (N_48818,N_47713,N_47785);
and U48819 (N_48819,N_47230,N_47753);
and U48820 (N_48820,N_47262,N_47582);
and U48821 (N_48821,N_47302,N_47632);
and U48822 (N_48822,N_47015,N_47071);
nand U48823 (N_48823,N_47080,N_47821);
or U48824 (N_48824,N_47834,N_47607);
and U48825 (N_48825,N_47569,N_47706);
nor U48826 (N_48826,N_47812,N_47364);
or U48827 (N_48827,N_47760,N_47746);
or U48828 (N_48828,N_47535,N_47262);
and U48829 (N_48829,N_47926,N_47901);
or U48830 (N_48830,N_47832,N_47809);
nor U48831 (N_48831,N_47267,N_47102);
and U48832 (N_48832,N_47022,N_47362);
or U48833 (N_48833,N_47104,N_47255);
nor U48834 (N_48834,N_47826,N_47273);
or U48835 (N_48835,N_47009,N_47804);
or U48836 (N_48836,N_47872,N_47349);
or U48837 (N_48837,N_47540,N_47704);
nor U48838 (N_48838,N_47740,N_47626);
nor U48839 (N_48839,N_47316,N_47545);
xor U48840 (N_48840,N_47966,N_47913);
xnor U48841 (N_48841,N_47268,N_47036);
nor U48842 (N_48842,N_47937,N_47898);
nor U48843 (N_48843,N_47015,N_47615);
nand U48844 (N_48844,N_47526,N_47966);
or U48845 (N_48845,N_47999,N_47134);
and U48846 (N_48846,N_47196,N_47696);
or U48847 (N_48847,N_47766,N_47447);
and U48848 (N_48848,N_47255,N_47497);
nand U48849 (N_48849,N_47563,N_47022);
xor U48850 (N_48850,N_47662,N_47307);
xnor U48851 (N_48851,N_47502,N_47212);
nand U48852 (N_48852,N_47379,N_47456);
nand U48853 (N_48853,N_47565,N_47862);
or U48854 (N_48854,N_47719,N_47084);
nand U48855 (N_48855,N_47195,N_47872);
or U48856 (N_48856,N_47942,N_47240);
xnor U48857 (N_48857,N_47713,N_47223);
and U48858 (N_48858,N_47959,N_47265);
nor U48859 (N_48859,N_47899,N_47040);
and U48860 (N_48860,N_47643,N_47348);
xnor U48861 (N_48861,N_47611,N_47230);
nor U48862 (N_48862,N_47997,N_47381);
nor U48863 (N_48863,N_47426,N_47152);
or U48864 (N_48864,N_47259,N_47768);
nor U48865 (N_48865,N_47680,N_47697);
xnor U48866 (N_48866,N_47221,N_47088);
nor U48867 (N_48867,N_47943,N_47995);
and U48868 (N_48868,N_47223,N_47448);
xor U48869 (N_48869,N_47982,N_47056);
nand U48870 (N_48870,N_47954,N_47345);
and U48871 (N_48871,N_47070,N_47817);
nand U48872 (N_48872,N_47721,N_47149);
or U48873 (N_48873,N_47673,N_47105);
nor U48874 (N_48874,N_47304,N_47647);
or U48875 (N_48875,N_47827,N_47770);
nor U48876 (N_48876,N_47654,N_47008);
xnor U48877 (N_48877,N_47812,N_47731);
xor U48878 (N_48878,N_47275,N_47166);
and U48879 (N_48879,N_47022,N_47891);
or U48880 (N_48880,N_47580,N_47099);
xnor U48881 (N_48881,N_47311,N_47777);
or U48882 (N_48882,N_47710,N_47423);
nand U48883 (N_48883,N_47854,N_47021);
xor U48884 (N_48884,N_47471,N_47866);
and U48885 (N_48885,N_47321,N_47808);
xor U48886 (N_48886,N_47081,N_47181);
nand U48887 (N_48887,N_47501,N_47516);
and U48888 (N_48888,N_47026,N_47872);
and U48889 (N_48889,N_47239,N_47415);
or U48890 (N_48890,N_47752,N_47020);
and U48891 (N_48891,N_47377,N_47047);
or U48892 (N_48892,N_47242,N_47786);
xnor U48893 (N_48893,N_47839,N_47425);
nand U48894 (N_48894,N_47175,N_47613);
nor U48895 (N_48895,N_47529,N_47667);
nand U48896 (N_48896,N_47883,N_47167);
or U48897 (N_48897,N_47510,N_47306);
and U48898 (N_48898,N_47773,N_47088);
or U48899 (N_48899,N_47841,N_47504);
or U48900 (N_48900,N_47496,N_47939);
or U48901 (N_48901,N_47675,N_47883);
nand U48902 (N_48902,N_47384,N_47365);
nand U48903 (N_48903,N_47292,N_47283);
xor U48904 (N_48904,N_47760,N_47422);
nand U48905 (N_48905,N_47528,N_47157);
or U48906 (N_48906,N_47403,N_47087);
and U48907 (N_48907,N_47328,N_47054);
and U48908 (N_48908,N_47122,N_47491);
nand U48909 (N_48909,N_47412,N_47880);
nor U48910 (N_48910,N_47436,N_47309);
nand U48911 (N_48911,N_47729,N_47522);
nand U48912 (N_48912,N_47394,N_47749);
xor U48913 (N_48913,N_47899,N_47561);
xnor U48914 (N_48914,N_47428,N_47714);
xor U48915 (N_48915,N_47144,N_47032);
nand U48916 (N_48916,N_47463,N_47113);
xnor U48917 (N_48917,N_47146,N_47938);
or U48918 (N_48918,N_47815,N_47315);
and U48919 (N_48919,N_47658,N_47643);
nor U48920 (N_48920,N_47437,N_47645);
or U48921 (N_48921,N_47715,N_47329);
xnor U48922 (N_48922,N_47925,N_47675);
xor U48923 (N_48923,N_47413,N_47667);
nor U48924 (N_48924,N_47707,N_47987);
and U48925 (N_48925,N_47986,N_47562);
nand U48926 (N_48926,N_47868,N_47682);
or U48927 (N_48927,N_47832,N_47257);
nor U48928 (N_48928,N_47427,N_47273);
xnor U48929 (N_48929,N_47814,N_47089);
nand U48930 (N_48930,N_47872,N_47123);
xnor U48931 (N_48931,N_47114,N_47462);
and U48932 (N_48932,N_47352,N_47341);
nor U48933 (N_48933,N_47303,N_47278);
nand U48934 (N_48934,N_47825,N_47258);
xnor U48935 (N_48935,N_47505,N_47455);
nand U48936 (N_48936,N_47929,N_47293);
xor U48937 (N_48937,N_47717,N_47293);
and U48938 (N_48938,N_47600,N_47186);
nand U48939 (N_48939,N_47878,N_47790);
or U48940 (N_48940,N_47314,N_47771);
nor U48941 (N_48941,N_47560,N_47067);
nor U48942 (N_48942,N_47087,N_47035);
or U48943 (N_48943,N_47739,N_47076);
nand U48944 (N_48944,N_47071,N_47857);
xor U48945 (N_48945,N_47056,N_47975);
and U48946 (N_48946,N_47106,N_47801);
nor U48947 (N_48947,N_47658,N_47695);
nor U48948 (N_48948,N_47139,N_47592);
or U48949 (N_48949,N_47500,N_47352);
and U48950 (N_48950,N_47012,N_47792);
nand U48951 (N_48951,N_47647,N_47387);
and U48952 (N_48952,N_47686,N_47781);
and U48953 (N_48953,N_47461,N_47322);
nor U48954 (N_48954,N_47133,N_47989);
and U48955 (N_48955,N_47969,N_47235);
nor U48956 (N_48956,N_47769,N_47665);
nand U48957 (N_48957,N_47754,N_47642);
or U48958 (N_48958,N_47695,N_47910);
xnor U48959 (N_48959,N_47478,N_47419);
nand U48960 (N_48960,N_47346,N_47256);
and U48961 (N_48961,N_47797,N_47557);
nor U48962 (N_48962,N_47272,N_47199);
xor U48963 (N_48963,N_47976,N_47686);
nor U48964 (N_48964,N_47947,N_47886);
xnor U48965 (N_48965,N_47495,N_47859);
nand U48966 (N_48966,N_47478,N_47692);
or U48967 (N_48967,N_47089,N_47537);
or U48968 (N_48968,N_47299,N_47201);
and U48969 (N_48969,N_47782,N_47263);
xnor U48970 (N_48970,N_47658,N_47290);
nand U48971 (N_48971,N_47323,N_47388);
xor U48972 (N_48972,N_47836,N_47524);
and U48973 (N_48973,N_47397,N_47206);
and U48974 (N_48974,N_47513,N_47293);
or U48975 (N_48975,N_47818,N_47897);
or U48976 (N_48976,N_47012,N_47440);
nor U48977 (N_48977,N_47308,N_47460);
nor U48978 (N_48978,N_47087,N_47974);
and U48979 (N_48979,N_47122,N_47666);
or U48980 (N_48980,N_47055,N_47858);
and U48981 (N_48981,N_47620,N_47968);
xnor U48982 (N_48982,N_47887,N_47650);
nand U48983 (N_48983,N_47976,N_47740);
or U48984 (N_48984,N_47787,N_47208);
nor U48985 (N_48985,N_47125,N_47105);
nand U48986 (N_48986,N_47585,N_47570);
xor U48987 (N_48987,N_47341,N_47649);
nand U48988 (N_48988,N_47372,N_47060);
xor U48989 (N_48989,N_47409,N_47217);
or U48990 (N_48990,N_47036,N_47132);
and U48991 (N_48991,N_47177,N_47587);
nand U48992 (N_48992,N_47022,N_47892);
xor U48993 (N_48993,N_47682,N_47634);
nor U48994 (N_48994,N_47836,N_47608);
or U48995 (N_48995,N_47615,N_47619);
nor U48996 (N_48996,N_47008,N_47634);
xnor U48997 (N_48997,N_47745,N_47235);
nand U48998 (N_48998,N_47774,N_47027);
nor U48999 (N_48999,N_47049,N_47276);
xnor U49000 (N_49000,N_48254,N_48568);
or U49001 (N_49001,N_48566,N_48554);
or U49002 (N_49002,N_48418,N_48351);
and U49003 (N_49003,N_48592,N_48315);
nand U49004 (N_49004,N_48694,N_48402);
nor U49005 (N_49005,N_48074,N_48953);
xnor U49006 (N_49006,N_48437,N_48835);
or U49007 (N_49007,N_48628,N_48029);
nor U49008 (N_49008,N_48815,N_48938);
xnor U49009 (N_49009,N_48456,N_48041);
nand U49010 (N_49010,N_48278,N_48421);
nand U49011 (N_49011,N_48441,N_48809);
xor U49012 (N_49012,N_48075,N_48934);
or U49013 (N_49013,N_48546,N_48831);
and U49014 (N_49014,N_48625,N_48914);
xnor U49015 (N_49015,N_48868,N_48367);
or U49016 (N_49016,N_48436,N_48538);
nor U49017 (N_49017,N_48413,N_48755);
nand U49018 (N_49018,N_48655,N_48746);
and U49019 (N_49019,N_48607,N_48140);
and U49020 (N_49020,N_48739,N_48501);
nor U49021 (N_49021,N_48781,N_48676);
xor U49022 (N_49022,N_48925,N_48445);
nand U49023 (N_49023,N_48577,N_48811);
nor U49024 (N_49024,N_48508,N_48558);
xnor U49025 (N_49025,N_48492,N_48915);
xnor U49026 (N_49026,N_48232,N_48180);
xor U49027 (N_49027,N_48939,N_48826);
and U49028 (N_49028,N_48206,N_48887);
xor U49029 (N_49029,N_48740,N_48260);
or U49030 (N_49030,N_48670,N_48957);
xor U49031 (N_49031,N_48082,N_48886);
xor U49032 (N_49032,N_48010,N_48626);
xnor U49033 (N_49033,N_48369,N_48744);
nand U49034 (N_49034,N_48580,N_48808);
nand U49035 (N_49035,N_48723,N_48223);
nand U49036 (N_49036,N_48401,N_48641);
nand U49037 (N_49037,N_48702,N_48742);
xor U49038 (N_49038,N_48797,N_48872);
nand U49039 (N_49039,N_48446,N_48790);
nand U49040 (N_49040,N_48805,N_48590);
and U49041 (N_49041,N_48490,N_48384);
and U49042 (N_49042,N_48926,N_48185);
nand U49043 (N_49043,N_48018,N_48217);
or U49044 (N_49044,N_48770,N_48521);
nand U49045 (N_49045,N_48161,N_48220);
xor U49046 (N_49046,N_48017,N_48012);
nor U49047 (N_49047,N_48160,N_48366);
nor U49048 (N_49048,N_48171,N_48627);
or U49049 (N_49049,N_48997,N_48292);
or U49050 (N_49050,N_48430,N_48803);
nand U49051 (N_49051,N_48523,N_48020);
and U49052 (N_49052,N_48203,N_48178);
nor U49053 (N_49053,N_48272,N_48672);
and U49054 (N_49054,N_48055,N_48488);
nor U49055 (N_49055,N_48856,N_48602);
nor U49056 (N_49056,N_48334,N_48098);
nor U49057 (N_49057,N_48194,N_48861);
and U49058 (N_49058,N_48816,N_48423);
or U49059 (N_49059,N_48116,N_48309);
or U49060 (N_49060,N_48846,N_48720);
nor U49061 (N_49061,N_48349,N_48595);
or U49062 (N_49062,N_48647,N_48724);
nor U49063 (N_49063,N_48467,N_48143);
xnor U49064 (N_49064,N_48393,N_48543);
or U49065 (N_49065,N_48474,N_48903);
nor U49066 (N_49066,N_48230,N_48150);
nor U49067 (N_49067,N_48251,N_48005);
nor U49068 (N_49068,N_48221,N_48434);
nor U49069 (N_49069,N_48611,N_48355);
nor U49070 (N_49070,N_48164,N_48725);
xor U49071 (N_49071,N_48092,N_48202);
or U49072 (N_49072,N_48454,N_48907);
and U49073 (N_49073,N_48191,N_48930);
xor U49074 (N_49074,N_48037,N_48470);
nand U49075 (N_49075,N_48901,N_48606);
nand U49076 (N_49076,N_48473,N_48944);
or U49077 (N_49077,N_48560,N_48310);
xnor U49078 (N_49078,N_48428,N_48866);
and U49079 (N_49079,N_48163,N_48084);
nand U49080 (N_49080,N_48897,N_48978);
or U49081 (N_49081,N_48451,N_48968);
xor U49082 (N_49082,N_48593,N_48485);
nor U49083 (N_49083,N_48524,N_48536);
and U49084 (N_49084,N_48506,N_48553);
and U49085 (N_49085,N_48280,N_48398);
or U49086 (N_49086,N_48295,N_48357);
xor U49087 (N_49087,N_48954,N_48452);
nor U49088 (N_49088,N_48255,N_48646);
or U49089 (N_49089,N_48604,N_48644);
nor U49090 (N_49090,N_48618,N_48412);
nor U49091 (N_49091,N_48051,N_48813);
or U49092 (N_49092,N_48181,N_48064);
nor U49093 (N_49093,N_48124,N_48574);
and U49094 (N_49094,N_48489,N_48963);
xor U49095 (N_49095,N_48537,N_48006);
xnor U49096 (N_49096,N_48136,N_48865);
xnor U49097 (N_49097,N_48305,N_48187);
and U49098 (N_49098,N_48166,N_48209);
and U49099 (N_49099,N_48529,N_48857);
and U49100 (N_49100,N_48825,N_48520);
and U49101 (N_49101,N_48208,N_48952);
or U49102 (N_49102,N_48745,N_48756);
or U49103 (N_49103,N_48296,N_48243);
nor U49104 (N_49104,N_48833,N_48507);
and U49105 (N_49105,N_48383,N_48985);
nor U49106 (N_49106,N_48036,N_48500);
and U49107 (N_49107,N_48125,N_48563);
xor U49108 (N_49108,N_48876,N_48684);
and U49109 (N_49109,N_48513,N_48147);
or U49110 (N_49110,N_48482,N_48431);
or U49111 (N_49111,N_48639,N_48687);
xor U49112 (N_49112,N_48822,N_48101);
or U49113 (N_49113,N_48922,N_48878);
nand U49114 (N_49114,N_48395,N_48091);
nor U49115 (N_49115,N_48575,N_48732);
xnor U49116 (N_49116,N_48754,N_48733);
nand U49117 (N_49117,N_48573,N_48316);
xor U49118 (N_49118,N_48484,N_48659);
and U49119 (N_49119,N_48608,N_48863);
nand U49120 (N_49120,N_48080,N_48603);
nor U49121 (N_49121,N_48731,N_48975);
xor U49122 (N_49122,N_48916,N_48090);
nand U49123 (N_49123,N_48823,N_48556);
nor U49124 (N_49124,N_48552,N_48042);
nor U49125 (N_49125,N_48804,N_48333);
nand U49126 (N_49126,N_48757,N_48858);
xor U49127 (N_49127,N_48396,N_48768);
or U49128 (N_49128,N_48093,N_48612);
nand U49129 (N_49129,N_48601,N_48079);
nor U49130 (N_49130,N_48910,N_48287);
nor U49131 (N_49131,N_48961,N_48992);
and U49132 (N_49132,N_48875,N_48640);
or U49133 (N_49133,N_48576,N_48517);
or U49134 (N_49134,N_48559,N_48148);
nand U49135 (N_49135,N_48570,N_48491);
xor U49136 (N_49136,N_48864,N_48761);
and U49137 (N_49137,N_48698,N_48774);
nor U49138 (N_49138,N_48336,N_48548);
xnor U49139 (N_49139,N_48995,N_48767);
nand U49140 (N_49140,N_48319,N_48234);
nor U49141 (N_49141,N_48883,N_48651);
or U49142 (N_49142,N_48806,N_48867);
nor U49143 (N_49143,N_48519,N_48444);
xnor U49144 (N_49144,N_48104,N_48919);
xor U49145 (N_49145,N_48572,N_48195);
and U49146 (N_49146,N_48432,N_48365);
and U49147 (N_49147,N_48495,N_48526);
nor U49148 (N_49148,N_48274,N_48094);
nor U49149 (N_49149,N_48609,N_48541);
or U49150 (N_49150,N_48126,N_48859);
or U49151 (N_49151,N_48324,N_48844);
or U49152 (N_49152,N_48960,N_48668);
xor U49153 (N_49153,N_48120,N_48894);
and U49154 (N_49154,N_48154,N_48721);
or U49155 (N_49155,N_48810,N_48620);
and U49156 (N_49156,N_48214,N_48263);
or U49157 (N_49157,N_48070,N_48450);
xor U49158 (N_49158,N_48661,N_48685);
and U49159 (N_49159,N_48758,N_48048);
or U49160 (N_49160,N_48701,N_48845);
nor U49161 (N_49161,N_48843,N_48636);
nand U49162 (N_49162,N_48019,N_48989);
nor U49163 (N_49163,N_48929,N_48103);
nor U49164 (N_49164,N_48372,N_48289);
nand U49165 (N_49165,N_48433,N_48654);
or U49166 (N_49166,N_48043,N_48946);
xor U49167 (N_49167,N_48184,N_48216);
and U49168 (N_49168,N_48061,N_48947);
and U49169 (N_49169,N_48696,N_48390);
nand U49170 (N_49170,N_48928,N_48337);
nor U49171 (N_49171,N_48072,N_48664);
or U49172 (N_49172,N_48741,N_48932);
nand U49173 (N_49173,N_48067,N_48719);
xor U49174 (N_49174,N_48215,N_48113);
xor U49175 (N_49175,N_48689,N_48110);
and U49176 (N_49176,N_48777,N_48496);
nor U49177 (N_49177,N_48167,N_48314);
or U49178 (N_49178,N_48293,N_48987);
xor U49179 (N_49179,N_48769,N_48138);
and U49180 (N_49180,N_48677,N_48582);
and U49181 (N_49181,N_48304,N_48127);
xnor U49182 (N_49182,N_48531,N_48213);
or U49183 (N_49183,N_48457,N_48077);
nand U49184 (N_49184,N_48149,N_48973);
xnor U49185 (N_49185,N_48873,N_48776);
nand U49186 (N_49186,N_48169,N_48983);
nand U49187 (N_49187,N_48860,N_48198);
xnor U49188 (N_49188,N_48447,N_48442);
or U49189 (N_49189,N_48045,N_48168);
nand U49190 (N_49190,N_48852,N_48129);
and U49191 (N_49191,N_48008,N_48986);
and U49192 (N_49192,N_48904,N_48068);
nor U49193 (N_49193,N_48902,N_48172);
and U49194 (N_49194,N_48550,N_48736);
and U49195 (N_49195,N_48416,N_48471);
or U49196 (N_49196,N_48346,N_48335);
or U49197 (N_49197,N_48242,N_48648);
xnor U49198 (N_49198,N_48708,N_48680);
nor U49199 (N_49199,N_48503,N_48812);
xor U49200 (N_49200,N_48047,N_48906);
xnor U49201 (N_49201,N_48404,N_48515);
nor U49202 (N_49202,N_48131,N_48182);
and U49203 (N_49203,N_48478,N_48512);
xor U49204 (N_49204,N_48145,N_48882);
xnor U49205 (N_49205,N_48591,N_48764);
and U49206 (N_49206,N_48578,N_48504);
xor U49207 (N_49207,N_48269,N_48974);
or U49208 (N_49208,N_48426,N_48132);
nand U49209 (N_49209,N_48238,N_48440);
xnor U49210 (N_49210,N_48834,N_48584);
nand U49211 (N_49211,N_48193,N_48734);
and U49212 (N_49212,N_48021,N_48851);
and U49213 (N_49213,N_48849,N_48759);
and U49214 (N_49214,N_48923,N_48253);
nor U49215 (N_49215,N_48463,N_48320);
xnor U49216 (N_49216,N_48557,N_48998);
or U49217 (N_49217,N_48400,N_48460);
nand U49218 (N_49218,N_48871,N_48486);
nand U49219 (N_49219,N_48307,N_48879);
nand U49220 (N_49220,N_48605,N_48631);
nor U49221 (N_49221,N_48839,N_48078);
or U49222 (N_49222,N_48798,N_48002);
xor U49223 (N_49223,N_48225,N_48435);
or U49224 (N_49224,N_48323,N_48058);
xor U49225 (N_49225,N_48245,N_48081);
nor U49226 (N_49226,N_48891,N_48801);
or U49227 (N_49227,N_48134,N_48197);
nand U49228 (N_49228,N_48089,N_48945);
xor U49229 (N_49229,N_48829,N_48999);
nor U49230 (N_49230,N_48342,N_48949);
nor U49231 (N_49231,N_48792,N_48419);
or U49232 (N_49232,N_48549,N_48361);
nor U49233 (N_49233,N_48224,N_48062);
or U49234 (N_49234,N_48675,N_48240);
nor U49235 (N_49235,N_48381,N_48981);
nand U49236 (N_49236,N_48505,N_48889);
xnor U49237 (N_49237,N_48425,N_48956);
and U49238 (N_49238,N_48108,N_48117);
xor U49239 (N_49239,N_48326,N_48086);
or U49240 (N_49240,N_48265,N_48955);
xnor U49241 (N_49241,N_48408,N_48033);
nand U49242 (N_49242,N_48669,N_48783);
nor U49243 (N_49243,N_48298,N_48933);
nand U49244 (N_49244,N_48762,N_48417);
nor U49245 (N_49245,N_48060,N_48279);
and U49246 (N_49246,N_48892,N_48115);
or U49247 (N_49247,N_48030,N_48597);
and U49248 (N_49248,N_48271,N_48406);
nand U49249 (N_49249,N_48348,N_48297);
or U49250 (N_49250,N_48535,N_48943);
and U49251 (N_49251,N_48237,N_48373);
and U49252 (N_49252,N_48196,N_48869);
or U49253 (N_49253,N_48231,N_48498);
xor U49254 (N_49254,N_48699,N_48414);
xor U49255 (N_49255,N_48667,N_48236);
or U49256 (N_49256,N_48966,N_48266);
xnor U49257 (N_49257,N_48893,N_48599);
nand U49258 (N_49258,N_48780,N_48913);
xor U49259 (N_49259,N_48128,N_48044);
nor U49260 (N_49260,N_48420,N_48258);
xor U49261 (N_49261,N_48711,N_48703);
and U49262 (N_49262,N_48650,N_48338);
nor U49263 (N_49263,N_48862,N_48422);
or U49264 (N_49264,N_48688,N_48969);
and U49265 (N_49265,N_48306,N_48246);
xnor U49266 (N_49266,N_48615,N_48874);
xnor U49267 (N_49267,N_48637,N_48638);
or U49268 (N_49268,N_48112,N_48011);
xor U49269 (N_49269,N_48257,N_48737);
xnor U49270 (N_49270,N_48817,N_48848);
or U49271 (N_49271,N_48895,N_48371);
and U49272 (N_49272,N_48399,N_48941);
or U49273 (N_49273,N_48502,N_48778);
nor U49274 (N_49274,N_48443,N_48705);
xor U49275 (N_49275,N_48158,N_48545);
nor U49276 (N_49276,N_48157,N_48802);
and U49277 (N_49277,N_48007,N_48097);
xor U49278 (N_49278,N_48118,N_48847);
nor U49279 (N_49279,N_48494,N_48382);
or U49280 (N_49280,N_48635,N_48793);
xor U49281 (N_49281,N_48581,N_48107);
nand U49282 (N_49282,N_48686,N_48343);
or U49283 (N_49283,N_48302,N_48350);
nand U49284 (N_49284,N_48458,N_48643);
and U49285 (N_49285,N_48226,N_48141);
or U49286 (N_49286,N_48653,N_48339);
nand U49287 (N_49287,N_48448,N_48634);
nor U49288 (N_49288,N_48964,N_48885);
xor U49289 (N_49289,N_48481,N_48958);
nor U49290 (N_49290,N_48388,N_48114);
or U49291 (N_49291,N_48119,N_48156);
or U49292 (N_49292,N_48329,N_48682);
or U49293 (N_49293,N_48820,N_48466);
and U49294 (N_49294,N_48996,N_48380);
and U49295 (N_49295,N_48294,N_48332);
nor U49296 (N_49296,N_48477,N_48622);
or U49297 (N_49297,N_48707,N_48789);
nand U49298 (N_49298,N_48616,N_48000);
nor U49299 (N_49299,N_48518,N_48972);
and U49300 (N_49300,N_48908,N_48821);
or U49301 (N_49301,N_48424,N_48814);
and U49302 (N_49302,N_48144,N_48053);
and U49303 (N_49303,N_48409,N_48712);
xnor U49304 (N_49304,N_48516,N_48468);
nand U49305 (N_49305,N_48087,N_48153);
or U49306 (N_49306,N_48256,N_48771);
and U49307 (N_49307,N_48722,N_48102);
or U49308 (N_49308,N_48069,N_48356);
and U49309 (N_49309,N_48173,N_48179);
and U49310 (N_49310,N_48912,N_48617);
nand U49311 (N_49311,N_48379,N_48497);
or U49312 (N_49312,N_48407,N_48850);
nand U49313 (N_49313,N_48971,N_48066);
xnor U49314 (N_49314,N_48328,N_48028);
xor U49315 (N_49315,N_48533,N_48152);
nand U49316 (N_49316,N_48674,N_48728);
xnor U49317 (N_49317,N_48765,N_48429);
xor U49318 (N_49318,N_48345,N_48840);
and U49319 (N_49319,N_48341,N_48666);
xor U49320 (N_49320,N_48645,N_48188);
nand U49321 (N_49321,N_48660,N_48009);
nand U49322 (N_49322,N_48937,N_48250);
nor U49323 (N_49323,N_48176,N_48587);
nand U49324 (N_49324,N_48073,N_48775);
nor U49325 (N_49325,N_48842,N_48273);
xor U49326 (N_49326,N_48527,N_48877);
and U49327 (N_49327,N_48555,N_48469);
xor U49328 (N_49328,N_48359,N_48854);
nor U49329 (N_49329,N_48013,N_48291);
nand U49330 (N_49330,N_48658,N_48819);
or U49331 (N_49331,N_48540,N_48514);
or U49332 (N_49332,N_48059,N_48730);
nand U49333 (N_49333,N_48818,N_48547);
and U49334 (N_49334,N_48076,N_48693);
xor U49335 (N_49335,N_48763,N_48511);
nor U49336 (N_49336,N_48729,N_48277);
nand U49337 (N_49337,N_48024,N_48054);
nor U49338 (N_49338,N_48375,N_48262);
or U49339 (N_49339,N_48397,N_48583);
xor U49340 (N_49340,N_48175,N_48227);
nor U49341 (N_49341,N_48522,N_48050);
nor U49342 (N_49342,N_48657,N_48370);
nor U49343 (N_49343,N_48717,N_48353);
xnor U49344 (N_49344,N_48211,N_48799);
and U49345 (N_49345,N_48088,N_48564);
nor U49346 (N_49346,N_48900,N_48376);
xor U49347 (N_49347,N_48567,N_48322);
nand U49348 (N_49348,N_48347,N_48633);
or U49349 (N_49349,N_48979,N_48321);
nand U49350 (N_49350,N_48403,N_48483);
nand U49351 (N_49351,N_48299,N_48942);
xnor U49352 (N_49352,N_48632,N_48189);
nor U49353 (N_49353,N_48713,N_48888);
nand U49354 (N_49354,N_48385,N_48600);
and U49355 (N_49355,N_48252,N_48718);
or U49356 (N_49356,N_48827,N_48853);
nand U49357 (N_49357,N_48233,N_48855);
xnor U49358 (N_49358,N_48965,N_48259);
and U49359 (N_49359,N_48162,N_48786);
and U49360 (N_49360,N_48690,N_48031);
or U49361 (N_49361,N_48619,N_48317);
and U49362 (N_49362,N_48111,N_48311);
nand U49363 (N_49363,N_48931,N_48629);
and U49364 (N_49364,N_48261,N_48649);
nor U49365 (N_49365,N_48032,N_48235);
or U49366 (N_49366,N_48313,N_48327);
or U49367 (N_49367,N_48023,N_48841);
nand U49368 (N_49368,N_48229,N_48530);
nand U49369 (N_49369,N_48427,N_48204);
or U49370 (N_49370,N_48784,N_48905);
and U49371 (N_49371,N_48281,N_48621);
and U49372 (N_49372,N_48772,N_48199);
nor U49373 (N_49373,N_48534,N_48325);
nor U49374 (N_49374,N_48579,N_48035);
nor U49375 (N_49375,N_48832,N_48787);
and U49376 (N_49376,N_48022,N_48264);
nor U49377 (N_49377,N_48300,N_48249);
nand U49378 (N_49378,N_48386,N_48652);
nand U49379 (N_49379,N_48828,N_48880);
and U49380 (N_49380,N_48714,N_48479);
or U49381 (N_49381,N_48461,N_48219);
or U49382 (N_49382,N_48331,N_48991);
nand U49383 (N_49383,N_48285,N_48982);
nor U49384 (N_49384,N_48268,N_48990);
and U49385 (N_49385,N_48354,N_48063);
or U49386 (N_49386,N_48760,N_48630);
or U49387 (N_49387,N_48462,N_48788);
xnor U49388 (N_49388,N_48830,N_48065);
and U49389 (N_49389,N_48935,N_48003);
nand U49390 (N_49390,N_48896,N_48870);
or U49391 (N_49391,N_48027,N_48681);
nand U49392 (N_49392,N_48312,N_48391);
and U49393 (N_49393,N_48190,N_48499);
xor U49394 (N_49394,N_48673,N_48918);
and U49395 (N_49395,N_48267,N_48836);
nand U49396 (N_49396,N_48994,N_48924);
xnor U49397 (N_49397,N_48034,N_48392);
xnor U49398 (N_49398,N_48283,N_48358);
or U49399 (N_49399,N_48344,N_48096);
nor U49400 (N_49400,N_48228,N_48165);
and U49401 (N_49401,N_48665,N_48014);
nor U49402 (N_49402,N_48984,N_48001);
or U49403 (N_49403,N_48679,N_48137);
nor U49404 (N_49404,N_48394,N_48565);
or U49405 (N_49405,N_48706,N_48239);
nand U49406 (N_49406,N_48951,N_48837);
xor U49407 (N_49407,N_48100,N_48025);
nor U49408 (N_49408,N_48340,N_48544);
nand U49409 (N_49409,N_48493,N_48794);
or U49410 (N_49410,N_48095,N_48807);
and U49411 (N_49411,N_48405,N_48151);
nand U49412 (N_49412,N_48303,N_48439);
xnor U49413 (N_49413,N_48671,N_48779);
or U49414 (N_49414,N_48795,N_48539);
nand U49415 (N_49415,N_48697,N_48950);
nand U49416 (N_49416,N_48276,N_48177);
xor U49417 (N_49417,N_48241,N_48360);
or U49418 (N_49418,N_48683,N_48201);
and U49419 (N_49419,N_48750,N_48284);
nand U49420 (N_49420,N_48330,N_48596);
nor U49421 (N_49421,N_48109,N_48248);
and U49422 (N_49422,N_48890,N_48449);
or U49423 (N_49423,N_48715,N_48598);
or U49424 (N_49424,N_48352,N_48748);
and U49425 (N_49425,N_48212,N_48838);
xnor U49426 (N_49426,N_48085,N_48927);
or U49427 (N_49427,N_48135,N_48624);
or U49428 (N_49428,N_48747,N_48709);
or U49429 (N_49429,N_48898,N_48743);
nor U49430 (N_49430,N_48623,N_48749);
nand U49431 (N_49431,N_48155,N_48959);
and U49432 (N_49432,N_48170,N_48004);
xnor U49433 (N_49433,N_48056,N_48704);
nor U49434 (N_49434,N_48275,N_48528);
or U49435 (N_49435,N_48561,N_48038);
xnor U49436 (N_49436,N_48589,N_48121);
and U49437 (N_49437,N_48920,N_48318);
xor U49438 (N_49438,N_48472,N_48363);
xor U49439 (N_49439,N_48200,N_48105);
nand U49440 (N_49440,N_48057,N_48039);
xnor U49441 (N_49441,N_48726,N_48205);
nor U49442 (N_49442,N_48976,N_48921);
or U49443 (N_49443,N_48782,N_48510);
nor U49444 (N_49444,N_48374,N_48387);
or U49445 (N_49445,N_48753,N_48464);
nand U49446 (N_49446,N_48710,N_48270);
xor U49447 (N_49447,N_48146,N_48099);
nand U49448 (N_49448,N_48210,N_48465);
or U49449 (N_49449,N_48791,N_48716);
nand U49450 (N_49450,N_48884,N_48106);
or U49451 (N_49451,N_48980,N_48663);
nor U49452 (N_49452,N_48288,N_48244);
nor U49453 (N_49453,N_48301,N_48967);
or U49454 (N_49454,N_48586,N_48016);
nor U49455 (N_49455,N_48692,N_48476);
and U49456 (N_49456,N_48911,N_48133);
nand U49457 (N_49457,N_48585,N_48183);
nand U49458 (N_49458,N_48480,N_48766);
xor U49459 (N_49459,N_48475,N_48411);
nand U49460 (N_49460,N_48378,N_48594);
or U49461 (N_49461,N_48752,N_48290);
and U49462 (N_49462,N_48738,N_48123);
xnor U49463 (N_49463,N_48571,N_48610);
and U49464 (N_49464,N_48026,N_48691);
nand U49465 (N_49465,N_48881,N_48207);
and U49466 (N_49466,N_48525,N_48542);
nand U49467 (N_49467,N_48192,N_48459);
nor U49468 (N_49468,N_48453,N_48362);
nor U49469 (N_49469,N_48993,N_48785);
nor U49470 (N_49470,N_48122,N_48642);
or U49471 (N_49471,N_48139,N_48218);
or U49472 (N_49472,N_48389,N_48532);
nand U49473 (N_49473,N_48899,N_48415);
nand U49474 (N_49474,N_48049,N_48455);
nand U49475 (N_49475,N_48308,N_48948);
xor U49476 (N_49476,N_48487,N_48071);
and U49477 (N_49477,N_48562,N_48046);
nand U49478 (N_49478,N_48174,N_48695);
or U49479 (N_49479,N_48282,N_48700);
and U49480 (N_49480,N_48678,N_48186);
xor U49481 (N_49481,N_48569,N_48083);
nand U49482 (N_49482,N_48735,N_48015);
nand U49483 (N_49483,N_48410,N_48988);
nor U49484 (N_49484,N_48509,N_48751);
xor U49485 (N_49485,N_48936,N_48377);
nand U49486 (N_49486,N_48796,N_48940);
nor U49487 (N_49487,N_48824,N_48727);
and U49488 (N_49488,N_48977,N_48551);
xnor U49489 (N_49489,N_48800,N_48368);
and U49490 (N_49490,N_48962,N_48040);
and U49491 (N_49491,N_48613,N_48614);
nand U49492 (N_49492,N_48917,N_48247);
or U49493 (N_49493,N_48656,N_48909);
nor U49494 (N_49494,N_48130,N_48142);
nor U49495 (N_49495,N_48970,N_48662);
and U49496 (N_49496,N_48159,N_48364);
or U49497 (N_49497,N_48052,N_48588);
nand U49498 (N_49498,N_48438,N_48773);
nand U49499 (N_49499,N_48222,N_48286);
or U49500 (N_49500,N_48923,N_48599);
or U49501 (N_49501,N_48571,N_48916);
nand U49502 (N_49502,N_48146,N_48255);
nor U49503 (N_49503,N_48385,N_48945);
nand U49504 (N_49504,N_48831,N_48189);
nand U49505 (N_49505,N_48005,N_48006);
nor U49506 (N_49506,N_48833,N_48533);
nor U49507 (N_49507,N_48736,N_48250);
and U49508 (N_49508,N_48147,N_48530);
and U49509 (N_49509,N_48806,N_48556);
xnor U49510 (N_49510,N_48600,N_48189);
xor U49511 (N_49511,N_48839,N_48601);
nor U49512 (N_49512,N_48485,N_48381);
or U49513 (N_49513,N_48280,N_48375);
and U49514 (N_49514,N_48957,N_48506);
nand U49515 (N_49515,N_48315,N_48271);
nor U49516 (N_49516,N_48521,N_48310);
or U49517 (N_49517,N_48896,N_48387);
and U49518 (N_49518,N_48947,N_48607);
xor U49519 (N_49519,N_48419,N_48006);
and U49520 (N_49520,N_48140,N_48487);
and U49521 (N_49521,N_48158,N_48188);
xnor U49522 (N_49522,N_48189,N_48595);
xor U49523 (N_49523,N_48554,N_48726);
xnor U49524 (N_49524,N_48684,N_48295);
xnor U49525 (N_49525,N_48362,N_48859);
nand U49526 (N_49526,N_48417,N_48545);
xnor U49527 (N_49527,N_48872,N_48845);
nor U49528 (N_49528,N_48413,N_48896);
and U49529 (N_49529,N_48253,N_48137);
nor U49530 (N_49530,N_48066,N_48498);
nor U49531 (N_49531,N_48933,N_48408);
and U49532 (N_49532,N_48152,N_48284);
nor U49533 (N_49533,N_48266,N_48282);
and U49534 (N_49534,N_48028,N_48437);
xor U49535 (N_49535,N_48748,N_48842);
and U49536 (N_49536,N_48815,N_48213);
or U49537 (N_49537,N_48165,N_48720);
nor U49538 (N_49538,N_48805,N_48758);
xnor U49539 (N_49539,N_48000,N_48861);
and U49540 (N_49540,N_48957,N_48207);
nor U49541 (N_49541,N_48232,N_48018);
and U49542 (N_49542,N_48578,N_48557);
nand U49543 (N_49543,N_48141,N_48453);
xnor U49544 (N_49544,N_48001,N_48551);
nand U49545 (N_49545,N_48915,N_48665);
or U49546 (N_49546,N_48361,N_48662);
nand U49547 (N_49547,N_48146,N_48867);
nand U49548 (N_49548,N_48922,N_48843);
nand U49549 (N_49549,N_48370,N_48298);
nand U49550 (N_49550,N_48723,N_48221);
xnor U49551 (N_49551,N_48837,N_48972);
nand U49552 (N_49552,N_48952,N_48011);
xnor U49553 (N_49553,N_48646,N_48849);
nand U49554 (N_49554,N_48155,N_48465);
or U49555 (N_49555,N_48307,N_48331);
xor U49556 (N_49556,N_48707,N_48850);
nor U49557 (N_49557,N_48682,N_48184);
xnor U49558 (N_49558,N_48880,N_48934);
nor U49559 (N_49559,N_48021,N_48620);
nand U49560 (N_49560,N_48435,N_48891);
or U49561 (N_49561,N_48528,N_48666);
nand U49562 (N_49562,N_48085,N_48746);
and U49563 (N_49563,N_48714,N_48470);
nand U49564 (N_49564,N_48300,N_48766);
nand U49565 (N_49565,N_48951,N_48499);
nand U49566 (N_49566,N_48785,N_48902);
nand U49567 (N_49567,N_48583,N_48061);
nand U49568 (N_49568,N_48819,N_48900);
nor U49569 (N_49569,N_48019,N_48244);
or U49570 (N_49570,N_48089,N_48398);
and U49571 (N_49571,N_48822,N_48904);
nand U49572 (N_49572,N_48535,N_48027);
nor U49573 (N_49573,N_48587,N_48488);
and U49574 (N_49574,N_48105,N_48197);
nand U49575 (N_49575,N_48733,N_48171);
xor U49576 (N_49576,N_48215,N_48060);
nor U49577 (N_49577,N_48394,N_48763);
nand U49578 (N_49578,N_48110,N_48933);
nand U49579 (N_49579,N_48147,N_48305);
or U49580 (N_49580,N_48427,N_48868);
xnor U49581 (N_49581,N_48015,N_48169);
nor U49582 (N_49582,N_48397,N_48756);
xor U49583 (N_49583,N_48878,N_48918);
or U49584 (N_49584,N_48195,N_48625);
xnor U49585 (N_49585,N_48911,N_48028);
and U49586 (N_49586,N_48615,N_48793);
or U49587 (N_49587,N_48502,N_48662);
or U49588 (N_49588,N_48835,N_48097);
or U49589 (N_49589,N_48207,N_48843);
or U49590 (N_49590,N_48840,N_48936);
or U49591 (N_49591,N_48422,N_48078);
nor U49592 (N_49592,N_48570,N_48373);
and U49593 (N_49593,N_48945,N_48546);
and U49594 (N_49594,N_48504,N_48804);
nor U49595 (N_49595,N_48922,N_48919);
nor U49596 (N_49596,N_48281,N_48052);
nand U49597 (N_49597,N_48977,N_48416);
and U49598 (N_49598,N_48874,N_48435);
and U49599 (N_49599,N_48240,N_48545);
nand U49600 (N_49600,N_48964,N_48272);
nor U49601 (N_49601,N_48827,N_48778);
nor U49602 (N_49602,N_48817,N_48657);
and U49603 (N_49603,N_48796,N_48851);
and U49604 (N_49604,N_48756,N_48232);
xnor U49605 (N_49605,N_48967,N_48582);
or U49606 (N_49606,N_48836,N_48317);
nor U49607 (N_49607,N_48684,N_48123);
nor U49608 (N_49608,N_48702,N_48146);
and U49609 (N_49609,N_48869,N_48742);
nand U49610 (N_49610,N_48357,N_48362);
or U49611 (N_49611,N_48800,N_48179);
nand U49612 (N_49612,N_48899,N_48789);
nor U49613 (N_49613,N_48985,N_48676);
nand U49614 (N_49614,N_48119,N_48763);
xor U49615 (N_49615,N_48958,N_48697);
nand U49616 (N_49616,N_48536,N_48828);
and U49617 (N_49617,N_48799,N_48380);
and U49618 (N_49618,N_48438,N_48110);
or U49619 (N_49619,N_48277,N_48733);
or U49620 (N_49620,N_48757,N_48424);
nor U49621 (N_49621,N_48401,N_48525);
nor U49622 (N_49622,N_48877,N_48892);
nand U49623 (N_49623,N_48096,N_48523);
and U49624 (N_49624,N_48168,N_48197);
and U49625 (N_49625,N_48164,N_48941);
nand U49626 (N_49626,N_48793,N_48997);
and U49627 (N_49627,N_48413,N_48194);
and U49628 (N_49628,N_48751,N_48350);
nor U49629 (N_49629,N_48546,N_48365);
xor U49630 (N_49630,N_48570,N_48581);
xor U49631 (N_49631,N_48708,N_48950);
nor U49632 (N_49632,N_48200,N_48702);
nor U49633 (N_49633,N_48030,N_48000);
or U49634 (N_49634,N_48864,N_48275);
nand U49635 (N_49635,N_48692,N_48638);
and U49636 (N_49636,N_48898,N_48703);
xor U49637 (N_49637,N_48399,N_48337);
or U49638 (N_49638,N_48970,N_48480);
or U49639 (N_49639,N_48637,N_48886);
xnor U49640 (N_49640,N_48669,N_48875);
nor U49641 (N_49641,N_48470,N_48262);
nand U49642 (N_49642,N_48009,N_48060);
and U49643 (N_49643,N_48454,N_48817);
nor U49644 (N_49644,N_48351,N_48848);
and U49645 (N_49645,N_48663,N_48013);
nor U49646 (N_49646,N_48012,N_48440);
xnor U49647 (N_49647,N_48930,N_48653);
nor U49648 (N_49648,N_48702,N_48400);
nor U49649 (N_49649,N_48003,N_48815);
nor U49650 (N_49650,N_48783,N_48866);
nand U49651 (N_49651,N_48427,N_48292);
nor U49652 (N_49652,N_48344,N_48040);
and U49653 (N_49653,N_48564,N_48735);
and U49654 (N_49654,N_48501,N_48409);
or U49655 (N_49655,N_48381,N_48239);
nor U49656 (N_49656,N_48797,N_48331);
or U49657 (N_49657,N_48679,N_48979);
and U49658 (N_49658,N_48907,N_48879);
or U49659 (N_49659,N_48292,N_48068);
and U49660 (N_49660,N_48794,N_48491);
xnor U49661 (N_49661,N_48892,N_48598);
xnor U49662 (N_49662,N_48554,N_48123);
and U49663 (N_49663,N_48953,N_48047);
and U49664 (N_49664,N_48168,N_48340);
nor U49665 (N_49665,N_48519,N_48815);
nand U49666 (N_49666,N_48163,N_48371);
nand U49667 (N_49667,N_48069,N_48472);
nand U49668 (N_49668,N_48927,N_48953);
and U49669 (N_49669,N_48662,N_48210);
nand U49670 (N_49670,N_48977,N_48867);
or U49671 (N_49671,N_48194,N_48924);
nand U49672 (N_49672,N_48522,N_48898);
nand U49673 (N_49673,N_48748,N_48860);
or U49674 (N_49674,N_48337,N_48449);
and U49675 (N_49675,N_48493,N_48856);
nand U49676 (N_49676,N_48497,N_48724);
and U49677 (N_49677,N_48829,N_48027);
nand U49678 (N_49678,N_48142,N_48007);
nor U49679 (N_49679,N_48906,N_48894);
nor U49680 (N_49680,N_48612,N_48738);
or U49681 (N_49681,N_48491,N_48283);
xnor U49682 (N_49682,N_48220,N_48791);
nor U49683 (N_49683,N_48012,N_48514);
xnor U49684 (N_49684,N_48947,N_48282);
or U49685 (N_49685,N_48262,N_48755);
xor U49686 (N_49686,N_48405,N_48772);
nor U49687 (N_49687,N_48179,N_48925);
nor U49688 (N_49688,N_48817,N_48525);
or U49689 (N_49689,N_48904,N_48755);
nor U49690 (N_49690,N_48779,N_48634);
or U49691 (N_49691,N_48454,N_48751);
nand U49692 (N_49692,N_48921,N_48749);
or U49693 (N_49693,N_48477,N_48508);
nand U49694 (N_49694,N_48640,N_48838);
nor U49695 (N_49695,N_48810,N_48552);
nor U49696 (N_49696,N_48427,N_48862);
xnor U49697 (N_49697,N_48999,N_48095);
nand U49698 (N_49698,N_48318,N_48965);
or U49699 (N_49699,N_48238,N_48914);
or U49700 (N_49700,N_48679,N_48562);
nand U49701 (N_49701,N_48251,N_48647);
nand U49702 (N_49702,N_48033,N_48206);
xnor U49703 (N_49703,N_48883,N_48732);
and U49704 (N_49704,N_48488,N_48468);
and U49705 (N_49705,N_48471,N_48213);
xor U49706 (N_49706,N_48777,N_48294);
and U49707 (N_49707,N_48204,N_48166);
or U49708 (N_49708,N_48994,N_48722);
xnor U49709 (N_49709,N_48092,N_48246);
nor U49710 (N_49710,N_48640,N_48161);
xnor U49711 (N_49711,N_48182,N_48536);
and U49712 (N_49712,N_48124,N_48052);
nor U49713 (N_49713,N_48062,N_48866);
and U49714 (N_49714,N_48778,N_48898);
nor U49715 (N_49715,N_48379,N_48484);
and U49716 (N_49716,N_48045,N_48110);
xor U49717 (N_49717,N_48364,N_48331);
or U49718 (N_49718,N_48690,N_48491);
and U49719 (N_49719,N_48487,N_48355);
nor U49720 (N_49720,N_48867,N_48657);
nand U49721 (N_49721,N_48110,N_48615);
nor U49722 (N_49722,N_48651,N_48027);
nand U49723 (N_49723,N_48403,N_48513);
xor U49724 (N_49724,N_48063,N_48307);
nor U49725 (N_49725,N_48589,N_48137);
nand U49726 (N_49726,N_48415,N_48353);
nor U49727 (N_49727,N_48930,N_48387);
nand U49728 (N_49728,N_48342,N_48002);
xor U49729 (N_49729,N_48797,N_48708);
and U49730 (N_49730,N_48732,N_48098);
or U49731 (N_49731,N_48549,N_48801);
xnor U49732 (N_49732,N_48323,N_48012);
xnor U49733 (N_49733,N_48724,N_48969);
and U49734 (N_49734,N_48183,N_48002);
nand U49735 (N_49735,N_48359,N_48274);
or U49736 (N_49736,N_48787,N_48541);
or U49737 (N_49737,N_48378,N_48375);
and U49738 (N_49738,N_48586,N_48782);
or U49739 (N_49739,N_48869,N_48760);
or U49740 (N_49740,N_48657,N_48526);
nor U49741 (N_49741,N_48047,N_48842);
nor U49742 (N_49742,N_48869,N_48959);
xnor U49743 (N_49743,N_48805,N_48728);
nor U49744 (N_49744,N_48944,N_48945);
and U49745 (N_49745,N_48126,N_48402);
or U49746 (N_49746,N_48443,N_48477);
or U49747 (N_49747,N_48810,N_48740);
or U49748 (N_49748,N_48790,N_48104);
xnor U49749 (N_49749,N_48397,N_48652);
nand U49750 (N_49750,N_48174,N_48210);
xnor U49751 (N_49751,N_48492,N_48668);
or U49752 (N_49752,N_48932,N_48211);
and U49753 (N_49753,N_48490,N_48811);
xnor U49754 (N_49754,N_48028,N_48515);
and U49755 (N_49755,N_48284,N_48084);
and U49756 (N_49756,N_48876,N_48745);
xnor U49757 (N_49757,N_48665,N_48937);
xor U49758 (N_49758,N_48045,N_48621);
and U49759 (N_49759,N_48103,N_48912);
xnor U49760 (N_49760,N_48791,N_48150);
nor U49761 (N_49761,N_48116,N_48592);
xnor U49762 (N_49762,N_48972,N_48021);
nor U49763 (N_49763,N_48064,N_48217);
xor U49764 (N_49764,N_48119,N_48454);
xnor U49765 (N_49765,N_48339,N_48711);
xnor U49766 (N_49766,N_48055,N_48203);
nor U49767 (N_49767,N_48636,N_48492);
xnor U49768 (N_49768,N_48377,N_48880);
and U49769 (N_49769,N_48603,N_48404);
nor U49770 (N_49770,N_48533,N_48893);
and U49771 (N_49771,N_48643,N_48026);
and U49772 (N_49772,N_48511,N_48143);
and U49773 (N_49773,N_48255,N_48413);
nor U49774 (N_49774,N_48984,N_48050);
nand U49775 (N_49775,N_48173,N_48396);
xnor U49776 (N_49776,N_48150,N_48727);
xor U49777 (N_49777,N_48943,N_48958);
and U49778 (N_49778,N_48446,N_48351);
xor U49779 (N_49779,N_48531,N_48681);
or U49780 (N_49780,N_48418,N_48451);
xnor U49781 (N_49781,N_48601,N_48677);
nor U49782 (N_49782,N_48843,N_48483);
xnor U49783 (N_49783,N_48807,N_48888);
nor U49784 (N_49784,N_48528,N_48545);
nor U49785 (N_49785,N_48020,N_48806);
nor U49786 (N_49786,N_48433,N_48656);
or U49787 (N_49787,N_48795,N_48617);
nor U49788 (N_49788,N_48058,N_48351);
or U49789 (N_49789,N_48853,N_48578);
or U49790 (N_49790,N_48504,N_48651);
and U49791 (N_49791,N_48451,N_48096);
or U49792 (N_49792,N_48862,N_48431);
nor U49793 (N_49793,N_48349,N_48470);
xor U49794 (N_49794,N_48797,N_48594);
nor U49795 (N_49795,N_48989,N_48864);
nor U49796 (N_49796,N_48071,N_48752);
xnor U49797 (N_49797,N_48438,N_48675);
nand U49798 (N_49798,N_48917,N_48304);
nand U49799 (N_49799,N_48418,N_48981);
and U49800 (N_49800,N_48924,N_48828);
nor U49801 (N_49801,N_48252,N_48408);
nor U49802 (N_49802,N_48878,N_48149);
xor U49803 (N_49803,N_48387,N_48286);
nor U49804 (N_49804,N_48010,N_48902);
xor U49805 (N_49805,N_48538,N_48844);
nand U49806 (N_49806,N_48576,N_48943);
nor U49807 (N_49807,N_48871,N_48316);
nand U49808 (N_49808,N_48383,N_48593);
nand U49809 (N_49809,N_48516,N_48183);
nand U49810 (N_49810,N_48714,N_48318);
or U49811 (N_49811,N_48895,N_48347);
and U49812 (N_49812,N_48510,N_48376);
nand U49813 (N_49813,N_48978,N_48133);
xor U49814 (N_49814,N_48332,N_48318);
xnor U49815 (N_49815,N_48691,N_48887);
and U49816 (N_49816,N_48260,N_48095);
or U49817 (N_49817,N_48316,N_48070);
or U49818 (N_49818,N_48559,N_48457);
or U49819 (N_49819,N_48932,N_48398);
xnor U49820 (N_49820,N_48037,N_48175);
xnor U49821 (N_49821,N_48445,N_48782);
xor U49822 (N_49822,N_48192,N_48800);
and U49823 (N_49823,N_48479,N_48656);
and U49824 (N_49824,N_48418,N_48453);
xnor U49825 (N_49825,N_48364,N_48686);
nand U49826 (N_49826,N_48574,N_48190);
xor U49827 (N_49827,N_48250,N_48887);
xnor U49828 (N_49828,N_48074,N_48999);
or U49829 (N_49829,N_48002,N_48800);
or U49830 (N_49830,N_48595,N_48565);
xnor U49831 (N_49831,N_48210,N_48427);
and U49832 (N_49832,N_48731,N_48524);
nand U49833 (N_49833,N_48266,N_48853);
xnor U49834 (N_49834,N_48798,N_48338);
nor U49835 (N_49835,N_48390,N_48110);
nand U49836 (N_49836,N_48771,N_48157);
nand U49837 (N_49837,N_48418,N_48851);
nand U49838 (N_49838,N_48048,N_48963);
nand U49839 (N_49839,N_48446,N_48814);
nand U49840 (N_49840,N_48645,N_48259);
nor U49841 (N_49841,N_48958,N_48553);
or U49842 (N_49842,N_48638,N_48561);
nor U49843 (N_49843,N_48508,N_48983);
nor U49844 (N_49844,N_48259,N_48299);
nand U49845 (N_49845,N_48978,N_48284);
and U49846 (N_49846,N_48766,N_48305);
nor U49847 (N_49847,N_48871,N_48302);
or U49848 (N_49848,N_48387,N_48401);
or U49849 (N_49849,N_48063,N_48138);
nand U49850 (N_49850,N_48098,N_48541);
nor U49851 (N_49851,N_48046,N_48849);
or U49852 (N_49852,N_48286,N_48293);
nor U49853 (N_49853,N_48608,N_48264);
nand U49854 (N_49854,N_48947,N_48980);
nand U49855 (N_49855,N_48209,N_48420);
nor U49856 (N_49856,N_48246,N_48910);
nor U49857 (N_49857,N_48104,N_48432);
and U49858 (N_49858,N_48609,N_48163);
nor U49859 (N_49859,N_48055,N_48214);
nand U49860 (N_49860,N_48997,N_48949);
xor U49861 (N_49861,N_48465,N_48909);
xor U49862 (N_49862,N_48788,N_48342);
nand U49863 (N_49863,N_48086,N_48174);
or U49864 (N_49864,N_48387,N_48394);
and U49865 (N_49865,N_48406,N_48729);
or U49866 (N_49866,N_48593,N_48027);
or U49867 (N_49867,N_48364,N_48953);
or U49868 (N_49868,N_48450,N_48449);
nand U49869 (N_49869,N_48113,N_48482);
and U49870 (N_49870,N_48701,N_48159);
or U49871 (N_49871,N_48976,N_48199);
and U49872 (N_49872,N_48607,N_48310);
xnor U49873 (N_49873,N_48945,N_48236);
xor U49874 (N_49874,N_48174,N_48813);
nand U49875 (N_49875,N_48896,N_48205);
or U49876 (N_49876,N_48544,N_48782);
nand U49877 (N_49877,N_48166,N_48503);
or U49878 (N_49878,N_48342,N_48235);
or U49879 (N_49879,N_48955,N_48841);
and U49880 (N_49880,N_48154,N_48217);
or U49881 (N_49881,N_48963,N_48815);
nand U49882 (N_49882,N_48007,N_48752);
nand U49883 (N_49883,N_48944,N_48852);
nand U49884 (N_49884,N_48583,N_48830);
or U49885 (N_49885,N_48277,N_48291);
xnor U49886 (N_49886,N_48939,N_48312);
and U49887 (N_49887,N_48518,N_48085);
nand U49888 (N_49888,N_48028,N_48984);
and U49889 (N_49889,N_48050,N_48568);
nand U49890 (N_49890,N_48932,N_48597);
nor U49891 (N_49891,N_48279,N_48919);
nor U49892 (N_49892,N_48228,N_48645);
nor U49893 (N_49893,N_48690,N_48193);
xnor U49894 (N_49894,N_48937,N_48585);
and U49895 (N_49895,N_48526,N_48768);
and U49896 (N_49896,N_48901,N_48739);
or U49897 (N_49897,N_48656,N_48287);
and U49898 (N_49898,N_48511,N_48610);
nor U49899 (N_49899,N_48650,N_48204);
and U49900 (N_49900,N_48782,N_48747);
or U49901 (N_49901,N_48165,N_48750);
nor U49902 (N_49902,N_48460,N_48056);
and U49903 (N_49903,N_48464,N_48082);
nand U49904 (N_49904,N_48666,N_48090);
nor U49905 (N_49905,N_48741,N_48611);
xnor U49906 (N_49906,N_48046,N_48737);
nand U49907 (N_49907,N_48474,N_48788);
nand U49908 (N_49908,N_48194,N_48000);
or U49909 (N_49909,N_48112,N_48447);
nand U49910 (N_49910,N_48210,N_48391);
nor U49911 (N_49911,N_48977,N_48889);
nor U49912 (N_49912,N_48233,N_48561);
and U49913 (N_49913,N_48930,N_48515);
xor U49914 (N_49914,N_48545,N_48547);
xnor U49915 (N_49915,N_48228,N_48622);
or U49916 (N_49916,N_48128,N_48765);
or U49917 (N_49917,N_48353,N_48230);
nor U49918 (N_49918,N_48083,N_48332);
xnor U49919 (N_49919,N_48579,N_48362);
nand U49920 (N_49920,N_48581,N_48903);
or U49921 (N_49921,N_48659,N_48562);
xnor U49922 (N_49922,N_48361,N_48443);
nor U49923 (N_49923,N_48589,N_48931);
and U49924 (N_49924,N_48378,N_48372);
and U49925 (N_49925,N_48372,N_48708);
or U49926 (N_49926,N_48107,N_48750);
nand U49927 (N_49927,N_48047,N_48641);
nor U49928 (N_49928,N_48868,N_48884);
nand U49929 (N_49929,N_48042,N_48938);
or U49930 (N_49930,N_48887,N_48791);
nand U49931 (N_49931,N_48570,N_48107);
or U49932 (N_49932,N_48674,N_48828);
nor U49933 (N_49933,N_48854,N_48057);
nor U49934 (N_49934,N_48393,N_48970);
nor U49935 (N_49935,N_48075,N_48949);
xor U49936 (N_49936,N_48265,N_48542);
nand U49937 (N_49937,N_48266,N_48578);
and U49938 (N_49938,N_48724,N_48127);
nand U49939 (N_49939,N_48473,N_48832);
and U49940 (N_49940,N_48786,N_48825);
nor U49941 (N_49941,N_48786,N_48158);
nor U49942 (N_49942,N_48660,N_48338);
or U49943 (N_49943,N_48848,N_48969);
or U49944 (N_49944,N_48249,N_48722);
nand U49945 (N_49945,N_48135,N_48282);
and U49946 (N_49946,N_48212,N_48841);
xor U49947 (N_49947,N_48230,N_48289);
nor U49948 (N_49948,N_48170,N_48773);
xnor U49949 (N_49949,N_48160,N_48095);
or U49950 (N_49950,N_48461,N_48269);
or U49951 (N_49951,N_48231,N_48089);
nand U49952 (N_49952,N_48359,N_48362);
nand U49953 (N_49953,N_48890,N_48380);
or U49954 (N_49954,N_48387,N_48469);
or U49955 (N_49955,N_48376,N_48249);
nor U49956 (N_49956,N_48633,N_48518);
and U49957 (N_49957,N_48812,N_48717);
nor U49958 (N_49958,N_48956,N_48998);
nand U49959 (N_49959,N_48761,N_48038);
nor U49960 (N_49960,N_48523,N_48725);
nor U49961 (N_49961,N_48291,N_48293);
xnor U49962 (N_49962,N_48124,N_48654);
or U49963 (N_49963,N_48134,N_48001);
nor U49964 (N_49964,N_48337,N_48352);
nand U49965 (N_49965,N_48541,N_48657);
and U49966 (N_49966,N_48563,N_48952);
and U49967 (N_49967,N_48244,N_48494);
xor U49968 (N_49968,N_48949,N_48380);
nand U49969 (N_49969,N_48911,N_48747);
and U49970 (N_49970,N_48195,N_48733);
or U49971 (N_49971,N_48363,N_48428);
nand U49972 (N_49972,N_48207,N_48870);
or U49973 (N_49973,N_48694,N_48701);
nand U49974 (N_49974,N_48369,N_48021);
nand U49975 (N_49975,N_48585,N_48471);
nor U49976 (N_49976,N_48651,N_48025);
xnor U49977 (N_49977,N_48386,N_48357);
or U49978 (N_49978,N_48284,N_48728);
nand U49979 (N_49979,N_48031,N_48313);
or U49980 (N_49980,N_48378,N_48495);
or U49981 (N_49981,N_48661,N_48541);
nor U49982 (N_49982,N_48271,N_48447);
nor U49983 (N_49983,N_48851,N_48603);
or U49984 (N_49984,N_48638,N_48790);
and U49985 (N_49985,N_48856,N_48442);
xnor U49986 (N_49986,N_48570,N_48706);
nor U49987 (N_49987,N_48502,N_48354);
and U49988 (N_49988,N_48563,N_48672);
or U49989 (N_49989,N_48882,N_48089);
and U49990 (N_49990,N_48997,N_48842);
nand U49991 (N_49991,N_48662,N_48494);
nand U49992 (N_49992,N_48201,N_48030);
and U49993 (N_49993,N_48476,N_48374);
and U49994 (N_49994,N_48623,N_48498);
nor U49995 (N_49995,N_48131,N_48445);
or U49996 (N_49996,N_48247,N_48821);
nand U49997 (N_49997,N_48479,N_48978);
or U49998 (N_49998,N_48459,N_48748);
nand U49999 (N_49999,N_48198,N_48132);
nand UO_0 (O_0,N_49827,N_49035);
and UO_1 (O_1,N_49971,N_49613);
xor UO_2 (O_2,N_49418,N_49689);
xnor UO_3 (O_3,N_49978,N_49211);
nand UO_4 (O_4,N_49917,N_49156);
and UO_5 (O_5,N_49215,N_49120);
nand UO_6 (O_6,N_49564,N_49774);
and UO_7 (O_7,N_49737,N_49247);
xor UO_8 (O_8,N_49715,N_49632);
or UO_9 (O_9,N_49262,N_49937);
nor UO_10 (O_10,N_49458,N_49866);
nor UO_11 (O_11,N_49688,N_49697);
nor UO_12 (O_12,N_49029,N_49699);
xor UO_13 (O_13,N_49565,N_49437);
nand UO_14 (O_14,N_49114,N_49017);
nand UO_15 (O_15,N_49043,N_49544);
or UO_16 (O_16,N_49260,N_49097);
or UO_17 (O_17,N_49002,N_49951);
and UO_18 (O_18,N_49930,N_49568);
xnor UO_19 (O_19,N_49850,N_49063);
and UO_20 (O_20,N_49142,N_49611);
and UO_21 (O_21,N_49635,N_49224);
or UO_22 (O_22,N_49925,N_49704);
nor UO_23 (O_23,N_49187,N_49863);
nor UO_24 (O_24,N_49967,N_49435);
nor UO_25 (O_25,N_49077,N_49973);
nor UO_26 (O_26,N_49096,N_49333);
xor UO_27 (O_27,N_49497,N_49181);
or UO_28 (O_28,N_49230,N_49069);
nand UO_29 (O_29,N_49417,N_49048);
and UO_30 (O_30,N_49442,N_49463);
and UO_31 (O_31,N_49674,N_49316);
and UO_32 (O_32,N_49118,N_49042);
xor UO_33 (O_33,N_49678,N_49185);
nor UO_34 (O_34,N_49348,N_49374);
nand UO_35 (O_35,N_49558,N_49892);
and UO_36 (O_36,N_49844,N_49865);
xnor UO_37 (O_37,N_49542,N_49665);
nor UO_38 (O_38,N_49566,N_49111);
nand UO_39 (O_39,N_49398,N_49078);
or UO_40 (O_40,N_49084,N_49349);
or UO_41 (O_41,N_49231,N_49481);
nor UO_42 (O_42,N_49406,N_49412);
nor UO_43 (O_43,N_49893,N_49477);
and UO_44 (O_44,N_49770,N_49221);
nor UO_45 (O_45,N_49071,N_49277);
or UO_46 (O_46,N_49263,N_49296);
nor UO_47 (O_47,N_49436,N_49005);
nor UO_48 (O_48,N_49856,N_49778);
and UO_49 (O_49,N_49714,N_49131);
nor UO_50 (O_50,N_49027,N_49837);
xor UO_51 (O_51,N_49008,N_49815);
nor UO_52 (O_52,N_49001,N_49755);
xor UO_53 (O_53,N_49407,N_49546);
xnor UO_54 (O_54,N_49528,N_49482);
or UO_55 (O_55,N_49629,N_49679);
xor UO_56 (O_56,N_49462,N_49498);
xor UO_57 (O_57,N_49775,N_49425);
xnor UO_58 (O_58,N_49103,N_49431);
xnor UO_59 (O_59,N_49643,N_49824);
nand UO_60 (O_60,N_49534,N_49660);
nor UO_61 (O_61,N_49876,N_49499);
nor UO_62 (O_62,N_49014,N_49113);
nor UO_63 (O_63,N_49199,N_49501);
xor UO_64 (O_64,N_49050,N_49145);
and UO_65 (O_65,N_49479,N_49694);
xor UO_66 (O_66,N_49752,N_49175);
or UO_67 (O_67,N_49154,N_49377);
or UO_68 (O_68,N_49486,N_49299);
nand UO_69 (O_69,N_49556,N_49341);
nand UO_70 (O_70,N_49639,N_49238);
nor UO_71 (O_71,N_49064,N_49343);
nand UO_72 (O_72,N_49147,N_49272);
nand UO_73 (O_73,N_49057,N_49100);
nor UO_74 (O_74,N_49140,N_49276);
nand UO_75 (O_75,N_49738,N_49711);
nand UO_76 (O_76,N_49245,N_49725);
and UO_77 (O_77,N_49567,N_49642);
and UO_78 (O_78,N_49355,N_49692);
nor UO_79 (O_79,N_49781,N_49233);
nand UO_80 (O_80,N_49004,N_49936);
xor UO_81 (O_81,N_49172,N_49950);
nor UO_82 (O_82,N_49817,N_49516);
and UO_83 (O_83,N_49883,N_49091);
or UO_84 (O_84,N_49577,N_49378);
or UO_85 (O_85,N_49405,N_49987);
and UO_86 (O_86,N_49769,N_49779);
and UO_87 (O_87,N_49960,N_49445);
or UO_88 (O_88,N_49541,N_49943);
nor UO_89 (O_89,N_49828,N_49163);
and UO_90 (O_90,N_49659,N_49419);
or UO_91 (O_91,N_49803,N_49015);
nor UO_92 (O_92,N_49696,N_49724);
and UO_93 (O_93,N_49616,N_49321);
nor UO_94 (O_94,N_49439,N_49855);
nand UO_95 (O_95,N_49232,N_49751);
nor UO_96 (O_96,N_49510,N_49243);
nand UO_97 (O_97,N_49746,N_49143);
nand UO_98 (O_98,N_49018,N_49900);
and UO_99 (O_99,N_49133,N_49522);
and UO_100 (O_100,N_49625,N_49508);
nor UO_101 (O_101,N_49488,N_49072);
and UO_102 (O_102,N_49700,N_49790);
or UO_103 (O_103,N_49743,N_49947);
xnor UO_104 (O_104,N_49810,N_49748);
or UO_105 (O_105,N_49076,N_49440);
nor UO_106 (O_106,N_49806,N_49784);
nand UO_107 (O_107,N_49283,N_49535);
nor UO_108 (O_108,N_49288,N_49821);
nand UO_109 (O_109,N_49125,N_49684);
nor UO_110 (O_110,N_49919,N_49257);
or UO_111 (O_111,N_49630,N_49146);
or UO_112 (O_112,N_49836,N_49039);
or UO_113 (O_113,N_49841,N_49912);
xnor UO_114 (O_114,N_49661,N_49101);
xnor UO_115 (O_115,N_49839,N_49605);
or UO_116 (O_116,N_49466,N_49615);
nor UO_117 (O_117,N_49590,N_49222);
or UO_118 (O_118,N_49603,N_49180);
and UO_119 (O_119,N_49033,N_49273);
and UO_120 (O_120,N_49010,N_49640);
and UO_121 (O_121,N_49350,N_49081);
xnor UO_122 (O_122,N_49906,N_49368);
or UO_123 (O_123,N_49213,N_49470);
and UO_124 (O_124,N_49274,N_49177);
nand UO_125 (O_125,N_49673,N_49701);
nand UO_126 (O_126,N_49734,N_49792);
xnor UO_127 (O_127,N_49323,N_49414);
xor UO_128 (O_128,N_49956,N_49052);
xnor UO_129 (O_129,N_49586,N_49771);
or UO_130 (O_130,N_49965,N_49918);
nand UO_131 (O_131,N_49631,N_49484);
nor UO_132 (O_132,N_49090,N_49832);
or UO_133 (O_133,N_49526,N_49351);
and UO_134 (O_134,N_49862,N_49576);
and UO_135 (O_135,N_49990,N_49878);
and UO_136 (O_136,N_49130,N_49203);
nor UO_137 (O_137,N_49754,N_49791);
nor UO_138 (O_138,N_49882,N_49924);
or UO_139 (O_139,N_49223,N_49342);
nor UO_140 (O_140,N_49291,N_49106);
xnor UO_141 (O_141,N_49547,N_49730);
xnor UO_142 (O_142,N_49676,N_49427);
or UO_143 (O_143,N_49514,N_49581);
or UO_144 (O_144,N_49835,N_49713);
nand UO_145 (O_145,N_49195,N_49958);
or UO_146 (O_146,N_49413,N_49552);
nor UO_147 (O_147,N_49339,N_49383);
or UO_148 (O_148,N_49459,N_49135);
xnor UO_149 (O_149,N_49119,N_49996);
nor UO_150 (O_150,N_49986,N_49944);
or UO_151 (O_151,N_49691,N_49898);
nand UO_152 (O_152,N_49788,N_49085);
nand UO_153 (O_153,N_49287,N_49264);
nor UO_154 (O_154,N_49105,N_49468);
or UO_155 (O_155,N_49762,N_49226);
nand UO_156 (O_156,N_49196,N_49595);
and UO_157 (O_157,N_49877,N_49415);
nand UO_158 (O_158,N_49575,N_49957);
and UO_159 (O_159,N_49220,N_49471);
and UO_160 (O_160,N_49229,N_49198);
xnor UO_161 (O_161,N_49067,N_49520);
nor UO_162 (O_162,N_49599,N_49214);
nor UO_163 (O_163,N_49026,N_49244);
nand UO_164 (O_164,N_49046,N_49910);
and UO_165 (O_165,N_49388,N_49313);
nor UO_166 (O_166,N_49741,N_49151);
xnor UO_167 (O_167,N_49401,N_49805);
nor UO_168 (O_168,N_49500,N_49166);
xnor UO_169 (O_169,N_49895,N_49928);
xnor UO_170 (O_170,N_49330,N_49395);
nor UO_171 (O_171,N_49158,N_49749);
nand UO_172 (O_172,N_49776,N_49373);
nand UO_173 (O_173,N_49225,N_49766);
or UO_174 (O_174,N_49032,N_49455);
xnor UO_175 (O_175,N_49804,N_49550);
or UO_176 (O_176,N_49840,N_49563);
nor UO_177 (O_177,N_49517,N_49681);
or UO_178 (O_178,N_49347,N_49150);
or UO_179 (O_179,N_49169,N_49838);
xor UO_180 (O_180,N_49812,N_49980);
or UO_181 (O_181,N_49710,N_49739);
nand UO_182 (O_182,N_49447,N_49527);
or UO_183 (O_183,N_49066,N_49080);
or UO_184 (O_184,N_49235,N_49153);
nor UO_185 (O_185,N_49089,N_49529);
nor UO_186 (O_186,N_49851,N_49476);
nor UO_187 (O_187,N_49116,N_49370);
or UO_188 (O_188,N_49622,N_49829);
nor UO_189 (O_189,N_49456,N_49494);
and UO_190 (O_190,N_49496,N_49104);
nor UO_191 (O_191,N_49144,N_49644);
or UO_192 (O_192,N_49353,N_49310);
xnor UO_193 (O_193,N_49695,N_49795);
nor UO_194 (O_194,N_49843,N_49102);
and UO_195 (O_195,N_49942,N_49555);
nand UO_196 (O_196,N_49858,N_49206);
nor UO_197 (O_197,N_49946,N_49070);
and UO_198 (O_198,N_49049,N_49324);
nor UO_199 (O_199,N_49290,N_49492);
xor UO_200 (O_200,N_49361,N_49000);
nor UO_201 (O_201,N_49178,N_49628);
xor UO_202 (O_202,N_49281,N_49079);
or UO_203 (O_203,N_49627,N_49054);
and UO_204 (O_204,N_49972,N_49300);
nor UO_205 (O_205,N_49217,N_49816);
xor UO_206 (O_206,N_49783,N_49409);
nand UO_207 (O_207,N_49503,N_49578);
or UO_208 (O_208,N_49601,N_49597);
and UO_209 (O_209,N_49450,N_49592);
xor UO_210 (O_210,N_49793,N_49127);
nor UO_211 (O_211,N_49826,N_49813);
xor UO_212 (O_212,N_49410,N_49830);
nand UO_213 (O_213,N_49121,N_49404);
xnor UO_214 (O_214,N_49610,N_49190);
nand UO_215 (O_215,N_49164,N_49391);
nor UO_216 (O_216,N_49712,N_49473);
nand UO_217 (O_217,N_49464,N_49744);
or UO_218 (O_218,N_49016,N_49184);
or UO_219 (O_219,N_49985,N_49205);
nor UO_220 (O_220,N_49997,N_49652);
nand UO_221 (O_221,N_49504,N_49927);
xor UO_222 (O_222,N_49569,N_49524);
xnor UO_223 (O_223,N_49236,N_49201);
or UO_224 (O_224,N_49657,N_49051);
nand UO_225 (O_225,N_49088,N_49656);
nor UO_226 (O_226,N_49219,N_49717);
and UO_227 (O_227,N_49396,N_49637);
nand UO_228 (O_228,N_49891,N_49653);
nor UO_229 (O_229,N_49242,N_49303);
nand UO_230 (O_230,N_49325,N_49914);
or UO_231 (O_231,N_49159,N_49212);
or UO_232 (O_232,N_49871,N_49952);
nand UO_233 (O_233,N_49949,N_49995);
xnor UO_234 (O_234,N_49006,N_49059);
xnor UO_235 (O_235,N_49756,N_49671);
or UO_236 (O_236,N_49512,N_49905);
nand UO_237 (O_237,N_49536,N_49941);
or UO_238 (O_238,N_49358,N_49268);
xor UO_239 (O_239,N_49495,N_49240);
nand UO_240 (O_240,N_49654,N_49802);
or UO_241 (O_241,N_49687,N_49945);
nand UO_242 (O_242,N_49545,N_49908);
nor UO_243 (O_243,N_49626,N_49966);
and UO_244 (O_244,N_49718,N_49598);
xnor UO_245 (O_245,N_49831,N_49525);
and UO_246 (O_246,N_49428,N_49297);
nand UO_247 (O_247,N_49183,N_49399);
and UO_248 (O_248,N_49538,N_49367);
xor UO_249 (O_249,N_49868,N_49385);
or UO_250 (O_250,N_49619,N_49289);
nand UO_251 (O_251,N_49117,N_49709);
or UO_252 (O_252,N_49962,N_49003);
nor UO_253 (O_253,N_49270,N_49561);
and UO_254 (O_254,N_49726,N_49811);
nand UO_255 (O_255,N_49375,N_49636);
and UO_256 (O_256,N_49025,N_49707);
xnor UO_257 (O_257,N_49265,N_49607);
xor UO_258 (O_258,N_49612,N_49068);
nand UO_259 (O_259,N_49963,N_49160);
xnor UO_260 (O_260,N_49092,N_49842);
xnor UO_261 (O_261,N_49573,N_49095);
and UO_262 (O_262,N_49904,N_49761);
and UO_263 (O_263,N_49308,N_49392);
nand UO_264 (O_264,N_49162,N_49873);
nor UO_265 (O_265,N_49009,N_49833);
and UO_266 (O_266,N_49502,N_49278);
xor UO_267 (O_267,N_49115,N_49108);
nand UO_268 (O_268,N_49022,N_49721);
xnor UO_269 (O_269,N_49251,N_49320);
nor UO_270 (O_270,N_49354,N_49663);
nand UO_271 (O_271,N_49279,N_49531);
or UO_272 (O_272,N_49271,N_49808);
nand UO_273 (O_273,N_49571,N_49362);
nor UO_274 (O_274,N_49065,N_49800);
or UO_275 (O_275,N_49041,N_49060);
and UO_276 (O_276,N_49787,N_49490);
xnor UO_277 (O_277,N_49149,N_49940);
xnor UO_278 (O_278,N_49365,N_49706);
and UO_279 (O_279,N_49915,N_49888);
xor UO_280 (O_280,N_49931,N_49719);
and UO_281 (O_281,N_49551,N_49602);
nand UO_282 (O_282,N_49894,N_49328);
xnor UO_283 (O_283,N_49600,N_49294);
or UO_284 (O_284,N_49533,N_49747);
xor UO_285 (O_285,N_49369,N_49825);
or UO_286 (O_286,N_49519,N_49773);
nor UO_287 (O_287,N_49736,N_49200);
nor UO_288 (O_288,N_49782,N_49588);
nor UO_289 (O_289,N_49614,N_49469);
and UO_290 (O_290,N_49735,N_49823);
nor UO_291 (O_291,N_49194,N_49911);
nor UO_292 (O_292,N_49107,N_49921);
nor UO_293 (O_293,N_49887,N_49693);
xnor UO_294 (O_294,N_49028,N_49777);
xnor UO_295 (O_295,N_49173,N_49087);
nor UO_296 (O_296,N_49969,N_49618);
or UO_297 (O_297,N_49193,N_49820);
or UO_298 (O_298,N_49593,N_49620);
nand UO_299 (O_299,N_49847,N_49939);
nand UO_300 (O_300,N_49668,N_49188);
or UO_301 (O_301,N_49444,N_49218);
xnor UO_302 (O_302,N_49454,N_49394);
or UO_303 (O_303,N_49553,N_49979);
nor UO_304 (O_304,N_49591,N_49340);
and UO_305 (O_305,N_49968,N_49138);
and UO_306 (O_306,N_49227,N_49926);
nor UO_307 (O_307,N_49452,N_49255);
or UO_308 (O_308,N_49210,N_49907);
and UO_309 (O_309,N_49305,N_49382);
and UO_310 (O_310,N_49608,N_49861);
and UO_311 (O_311,N_49386,N_49315);
and UO_312 (O_312,N_49650,N_49352);
nor UO_313 (O_313,N_49886,N_49047);
or UO_314 (O_314,N_49849,N_49397);
and UO_315 (O_315,N_49112,N_49532);
or UO_316 (O_316,N_49472,N_49698);
nand UO_317 (O_317,N_49584,N_49543);
and UO_318 (O_318,N_49493,N_49124);
nor UO_319 (O_319,N_49923,N_49870);
or UO_320 (O_320,N_49438,N_49344);
and UO_321 (O_321,N_49768,N_49372);
nor UO_322 (O_322,N_49467,N_49582);
nor UO_323 (O_323,N_49648,N_49253);
and UO_324 (O_324,N_49056,N_49110);
and UO_325 (O_325,N_49982,N_49443);
and UO_326 (O_326,N_49617,N_49171);
nor UO_327 (O_327,N_49301,N_49023);
xnor UO_328 (O_328,N_49539,N_49261);
nand UO_329 (O_329,N_49157,N_49690);
xor UO_330 (O_330,N_49959,N_49794);
and UO_331 (O_331,N_49922,N_49624);
and UO_332 (O_332,N_49916,N_49318);
and UO_333 (O_333,N_49680,N_49745);
nor UO_334 (O_334,N_49583,N_49012);
and UO_335 (O_335,N_49819,N_49682);
xnor UO_336 (O_336,N_49393,N_49433);
and UO_337 (O_337,N_49651,N_49137);
xor UO_338 (O_338,N_49366,N_49729);
xor UO_339 (O_339,N_49909,N_49449);
and UO_340 (O_340,N_49356,N_49662);
and UO_341 (O_341,N_49441,N_49562);
nor UO_342 (O_342,N_49518,N_49322);
or UO_343 (O_343,N_49239,N_49757);
and UO_344 (O_344,N_49649,N_49034);
nor UO_345 (O_345,N_49403,N_49670);
xnor UO_346 (O_346,N_49400,N_49174);
nor UO_347 (O_347,N_49460,N_49875);
nand UO_348 (O_348,N_49345,N_49764);
or UO_349 (O_349,N_49451,N_49515);
and UO_350 (O_350,N_49126,N_49013);
nand UO_351 (O_351,N_49740,N_49275);
or UO_352 (O_352,N_49703,N_49880);
and UO_353 (O_353,N_49993,N_49786);
nor UO_354 (O_354,N_49513,N_49426);
nand UO_355 (O_355,N_49360,N_49030);
nand UO_356 (O_356,N_49929,N_49822);
nand UO_357 (O_357,N_49371,N_49666);
nand UO_358 (O_358,N_49763,N_49363);
nand UO_359 (O_359,N_49753,N_49991);
nor UO_360 (O_360,N_49728,N_49304);
xnor UO_361 (O_361,N_49557,N_49364);
nand UO_362 (O_362,N_49899,N_49634);
and UO_363 (O_363,N_49429,N_49570);
xor UO_364 (O_364,N_49326,N_49667);
xnor UO_365 (O_365,N_49478,N_49981);
xnor UO_366 (O_366,N_49938,N_49334);
nand UO_367 (O_367,N_49974,N_49075);
or UO_368 (O_368,N_49336,N_49548);
or UO_369 (O_369,N_49621,N_49387);
xor UO_370 (O_370,N_49489,N_49411);
nor UO_371 (O_371,N_49675,N_49293);
and UO_372 (O_372,N_49580,N_49953);
and UO_373 (O_373,N_49302,N_49845);
and UO_374 (O_374,N_49983,N_49335);
and UO_375 (O_375,N_49867,N_49772);
nor UO_376 (O_376,N_49186,N_49129);
xor UO_377 (O_377,N_49252,N_49148);
xnor UO_378 (O_378,N_49317,N_49572);
and UO_379 (O_379,N_49606,N_49708);
nand UO_380 (O_380,N_49669,N_49723);
xor UO_381 (O_381,N_49854,N_49881);
nor UO_382 (O_382,N_49457,N_49818);
nand UO_383 (O_383,N_49256,N_49073);
nor UO_384 (O_384,N_49141,N_49246);
nor UO_385 (O_385,N_49860,N_49086);
xor UO_386 (O_386,N_49984,N_49789);
nor UO_387 (O_387,N_49021,N_49337);
nand UO_388 (O_388,N_49579,N_49338);
xnor UO_389 (O_389,N_49037,N_49955);
xnor UO_390 (O_390,N_49430,N_49019);
and UO_391 (O_391,N_49280,N_49170);
and UO_392 (O_392,N_49475,N_49376);
nor UO_393 (O_393,N_49785,N_49731);
nand UO_394 (O_394,N_49448,N_49864);
nor UO_395 (O_395,N_49970,N_49540);
nor UO_396 (O_396,N_49999,N_49633);
nand UO_397 (O_397,N_49976,N_49647);
nand UO_398 (O_398,N_49589,N_49327);
nand UO_399 (O_399,N_49885,N_49062);
nor UO_400 (O_400,N_49474,N_49920);
or UO_401 (O_401,N_49521,N_49530);
and UO_402 (O_402,N_49155,N_49191);
xnor UO_403 (O_403,N_49380,N_49988);
nand UO_404 (O_404,N_49040,N_49020);
nand UO_405 (O_405,N_49872,N_49846);
and UO_406 (O_406,N_49903,N_49058);
and UO_407 (O_407,N_49152,N_49932);
and UO_408 (O_408,N_49128,N_49853);
and UO_409 (O_409,N_49587,N_49241);
nor UO_410 (O_410,N_49286,N_49596);
and UO_411 (O_411,N_49742,N_49207);
or UO_412 (O_412,N_49874,N_49007);
and UO_413 (O_413,N_49765,N_49549);
xnor UO_414 (O_414,N_49269,N_49282);
or UO_415 (O_415,N_49594,N_49480);
and UO_416 (O_416,N_49964,N_49416);
nand UO_417 (O_417,N_49209,N_49852);
nor UO_418 (O_418,N_49897,N_49848);
or UO_419 (O_419,N_49461,N_49053);
and UO_420 (O_420,N_49797,N_49672);
xor UO_421 (O_421,N_49292,N_49685);
nor UO_422 (O_422,N_49798,N_49483);
xor UO_423 (O_423,N_49179,N_49432);
nor UO_424 (O_424,N_49759,N_49182);
and UO_425 (O_425,N_49319,N_49585);
xor UO_426 (O_426,N_49176,N_49359);
nand UO_427 (O_427,N_49249,N_49389);
xor UO_428 (O_428,N_49686,N_49329);
nand UO_429 (O_429,N_49507,N_49312);
and UO_430 (O_430,N_49093,N_49267);
and UO_431 (O_431,N_49560,N_49446);
or UO_432 (O_432,N_49082,N_49408);
xor UO_433 (O_433,N_49574,N_49168);
and UO_434 (O_434,N_49331,N_49031);
or UO_435 (O_435,N_49998,N_49658);
xnor UO_436 (O_436,N_49722,N_49357);
nor UO_437 (O_437,N_49934,N_49055);
and UO_438 (O_438,N_49641,N_49204);
and UO_439 (O_439,N_49857,N_49948);
xor UO_440 (O_440,N_49123,N_49420);
and UO_441 (O_441,N_49801,N_49750);
nor UO_442 (O_442,N_49799,N_49165);
or UO_443 (O_443,N_49859,N_49045);
or UO_444 (O_444,N_49896,N_49537);
nor UO_445 (O_445,N_49705,N_49307);
or UO_446 (O_446,N_49250,N_49884);
nand UO_447 (O_447,N_49677,N_49228);
nand UO_448 (O_448,N_49134,N_49879);
and UO_449 (O_449,N_49098,N_49011);
or UO_450 (O_450,N_49890,N_49202);
and UO_451 (O_451,N_49933,N_49453);
nor UO_452 (O_452,N_49259,N_49796);
nand UO_453 (O_453,N_49234,N_49237);
nand UO_454 (O_454,N_49780,N_49189);
or UO_455 (O_455,N_49609,N_49683);
and UO_456 (O_456,N_49167,N_49381);
and UO_457 (O_457,N_49834,N_49487);
nand UO_458 (O_458,N_49346,N_49758);
or UO_459 (O_459,N_49284,N_49954);
or UO_460 (O_460,N_49132,N_49314);
nor UO_461 (O_461,N_49266,N_49422);
or UO_462 (O_462,N_49311,N_49254);
xor UO_463 (O_463,N_49889,N_49994);
nor UO_464 (O_464,N_49638,N_49094);
nor UO_465 (O_465,N_49109,N_49024);
nor UO_466 (O_466,N_49989,N_49975);
xnor UO_467 (O_467,N_49814,N_49161);
xnor UO_468 (O_468,N_49623,N_49604);
xnor UO_469 (O_469,N_49423,N_49044);
nand UO_470 (O_470,N_49248,N_49309);
or UO_471 (O_471,N_49645,N_49646);
nor UO_472 (O_472,N_49511,N_49807);
nand UO_473 (O_473,N_49424,N_49036);
and UO_474 (O_474,N_49306,N_49122);
nor UO_475 (O_475,N_49197,N_49402);
or UO_476 (O_476,N_49298,N_49216);
nand UO_477 (O_477,N_49139,N_49720);
nor UO_478 (O_478,N_49421,N_49192);
or UO_479 (O_479,N_49136,N_49992);
and UO_480 (O_480,N_49716,N_49379);
xor UO_481 (O_481,N_49902,N_49869);
xor UO_482 (O_482,N_49655,N_49809);
xor UO_483 (O_483,N_49961,N_49767);
xor UO_484 (O_484,N_49913,N_49760);
and UO_485 (O_485,N_49384,N_49258);
or UO_486 (O_486,N_49505,N_49702);
nor UO_487 (O_487,N_49559,N_49390);
xnor UO_488 (O_488,N_49506,N_49038);
and UO_489 (O_489,N_49491,N_49285);
or UO_490 (O_490,N_49434,N_49332);
xor UO_491 (O_491,N_49465,N_49977);
nand UO_492 (O_492,N_49523,N_49727);
nor UO_493 (O_493,N_49074,N_49099);
and UO_494 (O_494,N_49935,N_49554);
and UO_495 (O_495,N_49061,N_49208);
nand UO_496 (O_496,N_49733,N_49732);
and UO_497 (O_497,N_49509,N_49901);
and UO_498 (O_498,N_49295,N_49083);
nand UO_499 (O_499,N_49485,N_49664);
nand UO_500 (O_500,N_49928,N_49378);
xor UO_501 (O_501,N_49069,N_49204);
and UO_502 (O_502,N_49415,N_49946);
xnor UO_503 (O_503,N_49947,N_49763);
or UO_504 (O_504,N_49148,N_49673);
or UO_505 (O_505,N_49545,N_49786);
nor UO_506 (O_506,N_49462,N_49186);
and UO_507 (O_507,N_49033,N_49253);
and UO_508 (O_508,N_49473,N_49732);
and UO_509 (O_509,N_49254,N_49079);
and UO_510 (O_510,N_49235,N_49843);
and UO_511 (O_511,N_49441,N_49507);
nor UO_512 (O_512,N_49415,N_49100);
xor UO_513 (O_513,N_49302,N_49084);
nor UO_514 (O_514,N_49838,N_49689);
or UO_515 (O_515,N_49305,N_49254);
and UO_516 (O_516,N_49877,N_49226);
nand UO_517 (O_517,N_49004,N_49240);
or UO_518 (O_518,N_49604,N_49417);
nor UO_519 (O_519,N_49079,N_49238);
or UO_520 (O_520,N_49155,N_49661);
xor UO_521 (O_521,N_49531,N_49936);
xor UO_522 (O_522,N_49448,N_49134);
nor UO_523 (O_523,N_49423,N_49540);
and UO_524 (O_524,N_49792,N_49056);
and UO_525 (O_525,N_49164,N_49291);
or UO_526 (O_526,N_49289,N_49649);
xnor UO_527 (O_527,N_49817,N_49902);
nor UO_528 (O_528,N_49974,N_49152);
xnor UO_529 (O_529,N_49729,N_49561);
nand UO_530 (O_530,N_49754,N_49092);
nand UO_531 (O_531,N_49982,N_49379);
nor UO_532 (O_532,N_49240,N_49176);
nor UO_533 (O_533,N_49890,N_49662);
or UO_534 (O_534,N_49567,N_49732);
nor UO_535 (O_535,N_49042,N_49487);
nand UO_536 (O_536,N_49614,N_49403);
nor UO_537 (O_537,N_49985,N_49359);
nand UO_538 (O_538,N_49041,N_49635);
nor UO_539 (O_539,N_49159,N_49639);
nor UO_540 (O_540,N_49855,N_49034);
and UO_541 (O_541,N_49749,N_49906);
and UO_542 (O_542,N_49609,N_49387);
nor UO_543 (O_543,N_49694,N_49183);
or UO_544 (O_544,N_49921,N_49110);
and UO_545 (O_545,N_49217,N_49652);
and UO_546 (O_546,N_49284,N_49904);
nand UO_547 (O_547,N_49355,N_49915);
nor UO_548 (O_548,N_49434,N_49526);
or UO_549 (O_549,N_49501,N_49145);
nor UO_550 (O_550,N_49916,N_49107);
xor UO_551 (O_551,N_49110,N_49419);
nor UO_552 (O_552,N_49769,N_49944);
nor UO_553 (O_553,N_49117,N_49870);
nor UO_554 (O_554,N_49868,N_49037);
nand UO_555 (O_555,N_49081,N_49128);
nand UO_556 (O_556,N_49631,N_49807);
and UO_557 (O_557,N_49776,N_49537);
and UO_558 (O_558,N_49621,N_49747);
and UO_559 (O_559,N_49754,N_49668);
nand UO_560 (O_560,N_49935,N_49245);
or UO_561 (O_561,N_49035,N_49350);
nand UO_562 (O_562,N_49425,N_49412);
nor UO_563 (O_563,N_49464,N_49449);
xor UO_564 (O_564,N_49461,N_49649);
and UO_565 (O_565,N_49258,N_49358);
nor UO_566 (O_566,N_49163,N_49798);
xor UO_567 (O_567,N_49138,N_49797);
xor UO_568 (O_568,N_49584,N_49687);
and UO_569 (O_569,N_49967,N_49723);
nand UO_570 (O_570,N_49091,N_49679);
nor UO_571 (O_571,N_49126,N_49020);
or UO_572 (O_572,N_49452,N_49841);
nor UO_573 (O_573,N_49693,N_49826);
or UO_574 (O_574,N_49455,N_49690);
nor UO_575 (O_575,N_49490,N_49791);
and UO_576 (O_576,N_49013,N_49281);
nor UO_577 (O_577,N_49055,N_49456);
nand UO_578 (O_578,N_49577,N_49155);
xor UO_579 (O_579,N_49264,N_49780);
xor UO_580 (O_580,N_49027,N_49455);
nand UO_581 (O_581,N_49196,N_49867);
nor UO_582 (O_582,N_49590,N_49781);
xor UO_583 (O_583,N_49494,N_49132);
or UO_584 (O_584,N_49855,N_49005);
nor UO_585 (O_585,N_49436,N_49632);
nor UO_586 (O_586,N_49755,N_49115);
xnor UO_587 (O_587,N_49337,N_49819);
nand UO_588 (O_588,N_49727,N_49017);
nand UO_589 (O_589,N_49849,N_49832);
nor UO_590 (O_590,N_49075,N_49382);
nor UO_591 (O_591,N_49126,N_49834);
nor UO_592 (O_592,N_49280,N_49923);
nand UO_593 (O_593,N_49945,N_49870);
nor UO_594 (O_594,N_49809,N_49164);
nand UO_595 (O_595,N_49296,N_49107);
and UO_596 (O_596,N_49525,N_49048);
and UO_597 (O_597,N_49610,N_49172);
or UO_598 (O_598,N_49451,N_49404);
and UO_599 (O_599,N_49470,N_49942);
nor UO_600 (O_600,N_49175,N_49015);
xnor UO_601 (O_601,N_49255,N_49863);
and UO_602 (O_602,N_49098,N_49550);
nand UO_603 (O_603,N_49873,N_49523);
xor UO_604 (O_604,N_49277,N_49001);
nand UO_605 (O_605,N_49717,N_49257);
and UO_606 (O_606,N_49354,N_49879);
or UO_607 (O_607,N_49220,N_49167);
xor UO_608 (O_608,N_49839,N_49496);
xor UO_609 (O_609,N_49882,N_49789);
nand UO_610 (O_610,N_49404,N_49842);
or UO_611 (O_611,N_49315,N_49657);
or UO_612 (O_612,N_49743,N_49058);
or UO_613 (O_613,N_49669,N_49377);
or UO_614 (O_614,N_49142,N_49578);
nor UO_615 (O_615,N_49322,N_49881);
and UO_616 (O_616,N_49265,N_49761);
xor UO_617 (O_617,N_49870,N_49226);
and UO_618 (O_618,N_49976,N_49610);
nor UO_619 (O_619,N_49033,N_49284);
or UO_620 (O_620,N_49912,N_49404);
and UO_621 (O_621,N_49861,N_49709);
xor UO_622 (O_622,N_49558,N_49475);
nor UO_623 (O_623,N_49069,N_49080);
or UO_624 (O_624,N_49890,N_49691);
or UO_625 (O_625,N_49001,N_49391);
and UO_626 (O_626,N_49742,N_49100);
nor UO_627 (O_627,N_49628,N_49558);
nor UO_628 (O_628,N_49420,N_49622);
and UO_629 (O_629,N_49066,N_49596);
and UO_630 (O_630,N_49396,N_49335);
nand UO_631 (O_631,N_49407,N_49531);
xor UO_632 (O_632,N_49935,N_49341);
nand UO_633 (O_633,N_49859,N_49520);
nor UO_634 (O_634,N_49399,N_49300);
or UO_635 (O_635,N_49027,N_49461);
xnor UO_636 (O_636,N_49256,N_49910);
xor UO_637 (O_637,N_49413,N_49987);
and UO_638 (O_638,N_49894,N_49341);
or UO_639 (O_639,N_49599,N_49868);
and UO_640 (O_640,N_49545,N_49668);
nor UO_641 (O_641,N_49881,N_49584);
nor UO_642 (O_642,N_49318,N_49015);
and UO_643 (O_643,N_49729,N_49682);
or UO_644 (O_644,N_49153,N_49437);
or UO_645 (O_645,N_49521,N_49355);
xor UO_646 (O_646,N_49961,N_49584);
and UO_647 (O_647,N_49065,N_49487);
nor UO_648 (O_648,N_49564,N_49122);
nand UO_649 (O_649,N_49440,N_49590);
nor UO_650 (O_650,N_49259,N_49983);
and UO_651 (O_651,N_49514,N_49553);
nand UO_652 (O_652,N_49029,N_49675);
and UO_653 (O_653,N_49916,N_49153);
nor UO_654 (O_654,N_49531,N_49578);
nand UO_655 (O_655,N_49164,N_49378);
nor UO_656 (O_656,N_49691,N_49408);
nand UO_657 (O_657,N_49759,N_49194);
or UO_658 (O_658,N_49326,N_49573);
and UO_659 (O_659,N_49321,N_49365);
nand UO_660 (O_660,N_49291,N_49055);
xor UO_661 (O_661,N_49053,N_49029);
nor UO_662 (O_662,N_49049,N_49716);
xnor UO_663 (O_663,N_49401,N_49695);
nand UO_664 (O_664,N_49494,N_49337);
or UO_665 (O_665,N_49769,N_49635);
or UO_666 (O_666,N_49510,N_49577);
or UO_667 (O_667,N_49297,N_49049);
and UO_668 (O_668,N_49550,N_49097);
nand UO_669 (O_669,N_49176,N_49181);
or UO_670 (O_670,N_49944,N_49417);
nand UO_671 (O_671,N_49502,N_49375);
and UO_672 (O_672,N_49676,N_49614);
and UO_673 (O_673,N_49208,N_49941);
xor UO_674 (O_674,N_49283,N_49830);
nand UO_675 (O_675,N_49662,N_49211);
nand UO_676 (O_676,N_49161,N_49560);
or UO_677 (O_677,N_49354,N_49268);
xor UO_678 (O_678,N_49662,N_49945);
nand UO_679 (O_679,N_49628,N_49583);
nor UO_680 (O_680,N_49849,N_49710);
and UO_681 (O_681,N_49642,N_49221);
nor UO_682 (O_682,N_49067,N_49837);
nand UO_683 (O_683,N_49258,N_49972);
or UO_684 (O_684,N_49872,N_49067);
xor UO_685 (O_685,N_49869,N_49417);
nor UO_686 (O_686,N_49472,N_49718);
nor UO_687 (O_687,N_49925,N_49662);
or UO_688 (O_688,N_49678,N_49922);
or UO_689 (O_689,N_49284,N_49052);
nor UO_690 (O_690,N_49907,N_49152);
or UO_691 (O_691,N_49191,N_49470);
xor UO_692 (O_692,N_49524,N_49876);
or UO_693 (O_693,N_49684,N_49576);
and UO_694 (O_694,N_49735,N_49693);
xnor UO_695 (O_695,N_49831,N_49467);
and UO_696 (O_696,N_49723,N_49044);
and UO_697 (O_697,N_49679,N_49165);
or UO_698 (O_698,N_49343,N_49570);
xor UO_699 (O_699,N_49730,N_49513);
nor UO_700 (O_700,N_49295,N_49823);
nor UO_701 (O_701,N_49448,N_49847);
nor UO_702 (O_702,N_49280,N_49661);
or UO_703 (O_703,N_49475,N_49703);
nand UO_704 (O_704,N_49765,N_49016);
nor UO_705 (O_705,N_49347,N_49433);
or UO_706 (O_706,N_49101,N_49701);
nor UO_707 (O_707,N_49099,N_49671);
xnor UO_708 (O_708,N_49694,N_49090);
or UO_709 (O_709,N_49893,N_49886);
and UO_710 (O_710,N_49265,N_49632);
or UO_711 (O_711,N_49764,N_49605);
nand UO_712 (O_712,N_49427,N_49693);
nor UO_713 (O_713,N_49870,N_49787);
nand UO_714 (O_714,N_49381,N_49356);
nor UO_715 (O_715,N_49857,N_49841);
or UO_716 (O_716,N_49217,N_49973);
or UO_717 (O_717,N_49491,N_49334);
and UO_718 (O_718,N_49348,N_49245);
nand UO_719 (O_719,N_49649,N_49384);
xor UO_720 (O_720,N_49318,N_49896);
xnor UO_721 (O_721,N_49800,N_49914);
and UO_722 (O_722,N_49713,N_49384);
or UO_723 (O_723,N_49167,N_49363);
or UO_724 (O_724,N_49375,N_49560);
or UO_725 (O_725,N_49021,N_49764);
xnor UO_726 (O_726,N_49888,N_49292);
or UO_727 (O_727,N_49078,N_49369);
or UO_728 (O_728,N_49034,N_49857);
and UO_729 (O_729,N_49522,N_49232);
xor UO_730 (O_730,N_49539,N_49923);
xnor UO_731 (O_731,N_49325,N_49788);
nor UO_732 (O_732,N_49499,N_49904);
nand UO_733 (O_733,N_49774,N_49699);
xor UO_734 (O_734,N_49819,N_49475);
or UO_735 (O_735,N_49175,N_49324);
nor UO_736 (O_736,N_49231,N_49412);
nand UO_737 (O_737,N_49519,N_49231);
nor UO_738 (O_738,N_49846,N_49887);
xor UO_739 (O_739,N_49575,N_49152);
nor UO_740 (O_740,N_49076,N_49455);
and UO_741 (O_741,N_49783,N_49624);
nand UO_742 (O_742,N_49885,N_49824);
or UO_743 (O_743,N_49370,N_49331);
xnor UO_744 (O_744,N_49698,N_49808);
or UO_745 (O_745,N_49925,N_49581);
xor UO_746 (O_746,N_49535,N_49083);
nand UO_747 (O_747,N_49509,N_49691);
or UO_748 (O_748,N_49667,N_49734);
or UO_749 (O_749,N_49159,N_49665);
nand UO_750 (O_750,N_49321,N_49022);
nand UO_751 (O_751,N_49551,N_49340);
or UO_752 (O_752,N_49384,N_49244);
xnor UO_753 (O_753,N_49052,N_49782);
or UO_754 (O_754,N_49907,N_49277);
or UO_755 (O_755,N_49224,N_49769);
or UO_756 (O_756,N_49491,N_49667);
nor UO_757 (O_757,N_49331,N_49495);
or UO_758 (O_758,N_49921,N_49168);
nor UO_759 (O_759,N_49597,N_49230);
nand UO_760 (O_760,N_49805,N_49385);
nor UO_761 (O_761,N_49141,N_49378);
nand UO_762 (O_762,N_49218,N_49900);
or UO_763 (O_763,N_49293,N_49113);
xor UO_764 (O_764,N_49544,N_49640);
and UO_765 (O_765,N_49620,N_49223);
nand UO_766 (O_766,N_49965,N_49050);
or UO_767 (O_767,N_49638,N_49336);
xnor UO_768 (O_768,N_49177,N_49340);
nand UO_769 (O_769,N_49624,N_49322);
xnor UO_770 (O_770,N_49690,N_49600);
and UO_771 (O_771,N_49164,N_49680);
or UO_772 (O_772,N_49408,N_49444);
xor UO_773 (O_773,N_49114,N_49221);
and UO_774 (O_774,N_49140,N_49957);
or UO_775 (O_775,N_49224,N_49464);
nand UO_776 (O_776,N_49018,N_49390);
xor UO_777 (O_777,N_49074,N_49605);
nor UO_778 (O_778,N_49851,N_49290);
xnor UO_779 (O_779,N_49565,N_49239);
and UO_780 (O_780,N_49543,N_49077);
or UO_781 (O_781,N_49263,N_49082);
xor UO_782 (O_782,N_49183,N_49586);
nand UO_783 (O_783,N_49915,N_49875);
and UO_784 (O_784,N_49844,N_49881);
or UO_785 (O_785,N_49164,N_49450);
or UO_786 (O_786,N_49094,N_49345);
xnor UO_787 (O_787,N_49310,N_49525);
nand UO_788 (O_788,N_49894,N_49604);
xnor UO_789 (O_789,N_49491,N_49555);
xor UO_790 (O_790,N_49898,N_49378);
and UO_791 (O_791,N_49407,N_49079);
nand UO_792 (O_792,N_49781,N_49799);
or UO_793 (O_793,N_49295,N_49357);
or UO_794 (O_794,N_49059,N_49218);
xnor UO_795 (O_795,N_49871,N_49754);
xnor UO_796 (O_796,N_49406,N_49676);
and UO_797 (O_797,N_49264,N_49658);
and UO_798 (O_798,N_49711,N_49525);
nor UO_799 (O_799,N_49337,N_49484);
or UO_800 (O_800,N_49045,N_49351);
nor UO_801 (O_801,N_49123,N_49451);
nand UO_802 (O_802,N_49840,N_49956);
nor UO_803 (O_803,N_49985,N_49538);
nor UO_804 (O_804,N_49339,N_49721);
and UO_805 (O_805,N_49757,N_49231);
nor UO_806 (O_806,N_49836,N_49450);
nor UO_807 (O_807,N_49278,N_49377);
nand UO_808 (O_808,N_49699,N_49282);
and UO_809 (O_809,N_49512,N_49844);
nand UO_810 (O_810,N_49897,N_49685);
nand UO_811 (O_811,N_49086,N_49025);
or UO_812 (O_812,N_49036,N_49988);
nor UO_813 (O_813,N_49480,N_49586);
xor UO_814 (O_814,N_49557,N_49357);
nor UO_815 (O_815,N_49365,N_49810);
or UO_816 (O_816,N_49340,N_49348);
or UO_817 (O_817,N_49618,N_49848);
and UO_818 (O_818,N_49670,N_49680);
nor UO_819 (O_819,N_49645,N_49084);
nor UO_820 (O_820,N_49795,N_49175);
or UO_821 (O_821,N_49799,N_49754);
xor UO_822 (O_822,N_49691,N_49585);
nand UO_823 (O_823,N_49633,N_49891);
nor UO_824 (O_824,N_49772,N_49174);
nand UO_825 (O_825,N_49346,N_49581);
xor UO_826 (O_826,N_49174,N_49824);
and UO_827 (O_827,N_49362,N_49221);
or UO_828 (O_828,N_49298,N_49240);
and UO_829 (O_829,N_49420,N_49112);
or UO_830 (O_830,N_49375,N_49421);
nor UO_831 (O_831,N_49102,N_49729);
or UO_832 (O_832,N_49406,N_49343);
and UO_833 (O_833,N_49059,N_49581);
nor UO_834 (O_834,N_49180,N_49359);
and UO_835 (O_835,N_49702,N_49865);
or UO_836 (O_836,N_49444,N_49946);
xnor UO_837 (O_837,N_49231,N_49561);
nor UO_838 (O_838,N_49567,N_49814);
xnor UO_839 (O_839,N_49224,N_49565);
and UO_840 (O_840,N_49337,N_49526);
xnor UO_841 (O_841,N_49019,N_49477);
nor UO_842 (O_842,N_49531,N_49693);
nand UO_843 (O_843,N_49549,N_49406);
nor UO_844 (O_844,N_49653,N_49640);
or UO_845 (O_845,N_49525,N_49126);
xnor UO_846 (O_846,N_49078,N_49176);
or UO_847 (O_847,N_49101,N_49860);
and UO_848 (O_848,N_49955,N_49775);
nor UO_849 (O_849,N_49099,N_49666);
nor UO_850 (O_850,N_49112,N_49603);
xnor UO_851 (O_851,N_49502,N_49637);
nand UO_852 (O_852,N_49331,N_49476);
nand UO_853 (O_853,N_49471,N_49447);
or UO_854 (O_854,N_49235,N_49403);
xor UO_855 (O_855,N_49126,N_49294);
nor UO_856 (O_856,N_49208,N_49464);
nor UO_857 (O_857,N_49009,N_49382);
nor UO_858 (O_858,N_49277,N_49745);
xnor UO_859 (O_859,N_49750,N_49889);
nand UO_860 (O_860,N_49197,N_49227);
and UO_861 (O_861,N_49475,N_49361);
or UO_862 (O_862,N_49925,N_49615);
nand UO_863 (O_863,N_49308,N_49079);
or UO_864 (O_864,N_49458,N_49171);
or UO_865 (O_865,N_49989,N_49981);
or UO_866 (O_866,N_49580,N_49218);
and UO_867 (O_867,N_49296,N_49535);
and UO_868 (O_868,N_49364,N_49665);
and UO_869 (O_869,N_49782,N_49118);
and UO_870 (O_870,N_49829,N_49018);
and UO_871 (O_871,N_49238,N_49047);
and UO_872 (O_872,N_49155,N_49114);
or UO_873 (O_873,N_49741,N_49192);
xor UO_874 (O_874,N_49303,N_49984);
nand UO_875 (O_875,N_49073,N_49982);
and UO_876 (O_876,N_49848,N_49971);
and UO_877 (O_877,N_49539,N_49434);
nand UO_878 (O_878,N_49396,N_49839);
nor UO_879 (O_879,N_49641,N_49004);
nand UO_880 (O_880,N_49923,N_49751);
nand UO_881 (O_881,N_49657,N_49308);
nor UO_882 (O_882,N_49239,N_49515);
xnor UO_883 (O_883,N_49363,N_49772);
nor UO_884 (O_884,N_49694,N_49786);
xnor UO_885 (O_885,N_49108,N_49855);
xor UO_886 (O_886,N_49974,N_49224);
or UO_887 (O_887,N_49540,N_49252);
nand UO_888 (O_888,N_49146,N_49315);
nor UO_889 (O_889,N_49801,N_49819);
and UO_890 (O_890,N_49838,N_49422);
xor UO_891 (O_891,N_49319,N_49459);
nor UO_892 (O_892,N_49013,N_49986);
nand UO_893 (O_893,N_49476,N_49391);
xor UO_894 (O_894,N_49987,N_49838);
xnor UO_895 (O_895,N_49417,N_49601);
and UO_896 (O_896,N_49727,N_49279);
and UO_897 (O_897,N_49471,N_49540);
nor UO_898 (O_898,N_49973,N_49349);
and UO_899 (O_899,N_49777,N_49628);
nor UO_900 (O_900,N_49202,N_49232);
xor UO_901 (O_901,N_49434,N_49985);
or UO_902 (O_902,N_49850,N_49410);
nand UO_903 (O_903,N_49083,N_49245);
or UO_904 (O_904,N_49794,N_49653);
and UO_905 (O_905,N_49193,N_49709);
nor UO_906 (O_906,N_49192,N_49140);
and UO_907 (O_907,N_49516,N_49068);
nor UO_908 (O_908,N_49824,N_49488);
nor UO_909 (O_909,N_49477,N_49942);
and UO_910 (O_910,N_49425,N_49348);
nand UO_911 (O_911,N_49712,N_49429);
nor UO_912 (O_912,N_49809,N_49552);
or UO_913 (O_913,N_49503,N_49180);
or UO_914 (O_914,N_49943,N_49554);
xnor UO_915 (O_915,N_49640,N_49262);
nor UO_916 (O_916,N_49834,N_49180);
nand UO_917 (O_917,N_49347,N_49092);
xor UO_918 (O_918,N_49234,N_49169);
and UO_919 (O_919,N_49949,N_49470);
or UO_920 (O_920,N_49832,N_49398);
xor UO_921 (O_921,N_49815,N_49205);
xnor UO_922 (O_922,N_49481,N_49268);
nor UO_923 (O_923,N_49379,N_49155);
nand UO_924 (O_924,N_49872,N_49871);
and UO_925 (O_925,N_49418,N_49666);
xor UO_926 (O_926,N_49631,N_49503);
nand UO_927 (O_927,N_49266,N_49256);
nor UO_928 (O_928,N_49021,N_49060);
xor UO_929 (O_929,N_49879,N_49864);
xnor UO_930 (O_930,N_49196,N_49897);
nor UO_931 (O_931,N_49909,N_49919);
nor UO_932 (O_932,N_49509,N_49783);
nor UO_933 (O_933,N_49106,N_49058);
nor UO_934 (O_934,N_49994,N_49562);
xnor UO_935 (O_935,N_49027,N_49460);
and UO_936 (O_936,N_49946,N_49693);
and UO_937 (O_937,N_49023,N_49842);
and UO_938 (O_938,N_49424,N_49044);
xnor UO_939 (O_939,N_49522,N_49173);
and UO_940 (O_940,N_49500,N_49825);
nand UO_941 (O_941,N_49087,N_49284);
or UO_942 (O_942,N_49072,N_49331);
or UO_943 (O_943,N_49467,N_49283);
and UO_944 (O_944,N_49037,N_49111);
or UO_945 (O_945,N_49824,N_49614);
xnor UO_946 (O_946,N_49549,N_49448);
nand UO_947 (O_947,N_49629,N_49937);
nor UO_948 (O_948,N_49571,N_49266);
nand UO_949 (O_949,N_49119,N_49773);
and UO_950 (O_950,N_49999,N_49690);
nand UO_951 (O_951,N_49672,N_49720);
nor UO_952 (O_952,N_49968,N_49980);
xnor UO_953 (O_953,N_49380,N_49337);
nor UO_954 (O_954,N_49962,N_49556);
nor UO_955 (O_955,N_49360,N_49868);
or UO_956 (O_956,N_49991,N_49035);
or UO_957 (O_957,N_49063,N_49287);
and UO_958 (O_958,N_49470,N_49783);
and UO_959 (O_959,N_49624,N_49262);
nand UO_960 (O_960,N_49294,N_49580);
or UO_961 (O_961,N_49313,N_49674);
nand UO_962 (O_962,N_49868,N_49227);
and UO_963 (O_963,N_49912,N_49580);
xor UO_964 (O_964,N_49562,N_49157);
and UO_965 (O_965,N_49287,N_49920);
xor UO_966 (O_966,N_49438,N_49704);
or UO_967 (O_967,N_49401,N_49958);
and UO_968 (O_968,N_49865,N_49550);
nor UO_969 (O_969,N_49773,N_49107);
nor UO_970 (O_970,N_49700,N_49433);
or UO_971 (O_971,N_49367,N_49902);
xor UO_972 (O_972,N_49128,N_49917);
and UO_973 (O_973,N_49350,N_49873);
and UO_974 (O_974,N_49730,N_49348);
nand UO_975 (O_975,N_49311,N_49954);
nor UO_976 (O_976,N_49308,N_49487);
nor UO_977 (O_977,N_49788,N_49912);
nor UO_978 (O_978,N_49705,N_49894);
or UO_979 (O_979,N_49438,N_49618);
nand UO_980 (O_980,N_49826,N_49400);
and UO_981 (O_981,N_49139,N_49491);
nand UO_982 (O_982,N_49452,N_49938);
nor UO_983 (O_983,N_49247,N_49233);
or UO_984 (O_984,N_49910,N_49187);
xor UO_985 (O_985,N_49880,N_49007);
nand UO_986 (O_986,N_49351,N_49831);
or UO_987 (O_987,N_49882,N_49676);
nand UO_988 (O_988,N_49407,N_49824);
nand UO_989 (O_989,N_49100,N_49728);
nor UO_990 (O_990,N_49802,N_49472);
or UO_991 (O_991,N_49314,N_49832);
nor UO_992 (O_992,N_49880,N_49722);
xor UO_993 (O_993,N_49145,N_49656);
xnor UO_994 (O_994,N_49881,N_49208);
or UO_995 (O_995,N_49552,N_49590);
and UO_996 (O_996,N_49740,N_49106);
xor UO_997 (O_997,N_49748,N_49787);
or UO_998 (O_998,N_49185,N_49193);
or UO_999 (O_999,N_49222,N_49584);
nor UO_1000 (O_1000,N_49271,N_49551);
nor UO_1001 (O_1001,N_49046,N_49769);
nor UO_1002 (O_1002,N_49598,N_49744);
nand UO_1003 (O_1003,N_49424,N_49410);
or UO_1004 (O_1004,N_49567,N_49288);
and UO_1005 (O_1005,N_49362,N_49994);
xnor UO_1006 (O_1006,N_49033,N_49838);
and UO_1007 (O_1007,N_49833,N_49495);
nand UO_1008 (O_1008,N_49832,N_49387);
nand UO_1009 (O_1009,N_49870,N_49723);
xor UO_1010 (O_1010,N_49838,N_49710);
xor UO_1011 (O_1011,N_49877,N_49748);
nor UO_1012 (O_1012,N_49480,N_49651);
or UO_1013 (O_1013,N_49560,N_49239);
xor UO_1014 (O_1014,N_49598,N_49933);
and UO_1015 (O_1015,N_49685,N_49560);
nand UO_1016 (O_1016,N_49585,N_49202);
nand UO_1017 (O_1017,N_49562,N_49287);
nand UO_1018 (O_1018,N_49358,N_49433);
nor UO_1019 (O_1019,N_49783,N_49755);
or UO_1020 (O_1020,N_49154,N_49584);
and UO_1021 (O_1021,N_49932,N_49599);
nor UO_1022 (O_1022,N_49402,N_49169);
and UO_1023 (O_1023,N_49543,N_49627);
and UO_1024 (O_1024,N_49020,N_49386);
xor UO_1025 (O_1025,N_49548,N_49192);
and UO_1026 (O_1026,N_49389,N_49111);
or UO_1027 (O_1027,N_49145,N_49372);
xor UO_1028 (O_1028,N_49209,N_49029);
or UO_1029 (O_1029,N_49570,N_49992);
or UO_1030 (O_1030,N_49570,N_49154);
xnor UO_1031 (O_1031,N_49966,N_49935);
nor UO_1032 (O_1032,N_49754,N_49953);
and UO_1033 (O_1033,N_49215,N_49192);
nor UO_1034 (O_1034,N_49142,N_49249);
xnor UO_1035 (O_1035,N_49019,N_49316);
xnor UO_1036 (O_1036,N_49753,N_49124);
or UO_1037 (O_1037,N_49601,N_49141);
nand UO_1038 (O_1038,N_49155,N_49021);
and UO_1039 (O_1039,N_49506,N_49189);
or UO_1040 (O_1040,N_49145,N_49160);
xnor UO_1041 (O_1041,N_49681,N_49814);
or UO_1042 (O_1042,N_49471,N_49183);
xnor UO_1043 (O_1043,N_49456,N_49950);
and UO_1044 (O_1044,N_49544,N_49261);
nor UO_1045 (O_1045,N_49686,N_49673);
nand UO_1046 (O_1046,N_49805,N_49874);
nand UO_1047 (O_1047,N_49198,N_49397);
xor UO_1048 (O_1048,N_49379,N_49287);
or UO_1049 (O_1049,N_49506,N_49332);
xnor UO_1050 (O_1050,N_49034,N_49577);
nor UO_1051 (O_1051,N_49684,N_49824);
and UO_1052 (O_1052,N_49909,N_49535);
nor UO_1053 (O_1053,N_49460,N_49753);
or UO_1054 (O_1054,N_49356,N_49599);
or UO_1055 (O_1055,N_49056,N_49499);
and UO_1056 (O_1056,N_49531,N_49640);
and UO_1057 (O_1057,N_49693,N_49932);
and UO_1058 (O_1058,N_49735,N_49213);
nor UO_1059 (O_1059,N_49474,N_49094);
nor UO_1060 (O_1060,N_49479,N_49404);
or UO_1061 (O_1061,N_49711,N_49718);
or UO_1062 (O_1062,N_49637,N_49190);
or UO_1063 (O_1063,N_49119,N_49581);
xnor UO_1064 (O_1064,N_49216,N_49574);
and UO_1065 (O_1065,N_49984,N_49370);
xnor UO_1066 (O_1066,N_49108,N_49087);
xnor UO_1067 (O_1067,N_49363,N_49844);
or UO_1068 (O_1068,N_49351,N_49296);
or UO_1069 (O_1069,N_49712,N_49825);
or UO_1070 (O_1070,N_49275,N_49995);
or UO_1071 (O_1071,N_49999,N_49330);
nor UO_1072 (O_1072,N_49081,N_49721);
and UO_1073 (O_1073,N_49169,N_49798);
nor UO_1074 (O_1074,N_49759,N_49462);
and UO_1075 (O_1075,N_49014,N_49292);
nand UO_1076 (O_1076,N_49977,N_49044);
nand UO_1077 (O_1077,N_49808,N_49700);
and UO_1078 (O_1078,N_49781,N_49604);
or UO_1079 (O_1079,N_49024,N_49765);
or UO_1080 (O_1080,N_49925,N_49930);
nand UO_1081 (O_1081,N_49879,N_49149);
nand UO_1082 (O_1082,N_49766,N_49677);
nand UO_1083 (O_1083,N_49009,N_49567);
nor UO_1084 (O_1084,N_49551,N_49774);
xor UO_1085 (O_1085,N_49892,N_49422);
nor UO_1086 (O_1086,N_49403,N_49556);
nor UO_1087 (O_1087,N_49494,N_49561);
xnor UO_1088 (O_1088,N_49063,N_49662);
or UO_1089 (O_1089,N_49160,N_49109);
or UO_1090 (O_1090,N_49110,N_49415);
or UO_1091 (O_1091,N_49000,N_49814);
xnor UO_1092 (O_1092,N_49252,N_49565);
nand UO_1093 (O_1093,N_49799,N_49325);
or UO_1094 (O_1094,N_49025,N_49133);
nand UO_1095 (O_1095,N_49039,N_49923);
and UO_1096 (O_1096,N_49475,N_49936);
xor UO_1097 (O_1097,N_49175,N_49701);
xor UO_1098 (O_1098,N_49725,N_49146);
or UO_1099 (O_1099,N_49721,N_49858);
xor UO_1100 (O_1100,N_49519,N_49527);
nor UO_1101 (O_1101,N_49829,N_49778);
and UO_1102 (O_1102,N_49767,N_49320);
nand UO_1103 (O_1103,N_49928,N_49760);
xnor UO_1104 (O_1104,N_49365,N_49548);
xor UO_1105 (O_1105,N_49484,N_49043);
xor UO_1106 (O_1106,N_49657,N_49766);
nand UO_1107 (O_1107,N_49531,N_49119);
xnor UO_1108 (O_1108,N_49951,N_49575);
nor UO_1109 (O_1109,N_49894,N_49485);
nand UO_1110 (O_1110,N_49234,N_49641);
or UO_1111 (O_1111,N_49214,N_49700);
nand UO_1112 (O_1112,N_49570,N_49480);
nand UO_1113 (O_1113,N_49738,N_49736);
xnor UO_1114 (O_1114,N_49332,N_49622);
xor UO_1115 (O_1115,N_49567,N_49264);
or UO_1116 (O_1116,N_49412,N_49899);
or UO_1117 (O_1117,N_49822,N_49545);
xnor UO_1118 (O_1118,N_49860,N_49674);
or UO_1119 (O_1119,N_49037,N_49022);
xor UO_1120 (O_1120,N_49291,N_49667);
nor UO_1121 (O_1121,N_49715,N_49635);
nand UO_1122 (O_1122,N_49787,N_49592);
or UO_1123 (O_1123,N_49214,N_49603);
xor UO_1124 (O_1124,N_49429,N_49909);
or UO_1125 (O_1125,N_49702,N_49185);
nand UO_1126 (O_1126,N_49737,N_49967);
nand UO_1127 (O_1127,N_49406,N_49297);
xnor UO_1128 (O_1128,N_49602,N_49383);
and UO_1129 (O_1129,N_49968,N_49560);
and UO_1130 (O_1130,N_49616,N_49303);
nor UO_1131 (O_1131,N_49599,N_49437);
nand UO_1132 (O_1132,N_49404,N_49622);
or UO_1133 (O_1133,N_49067,N_49224);
nand UO_1134 (O_1134,N_49511,N_49004);
or UO_1135 (O_1135,N_49409,N_49401);
or UO_1136 (O_1136,N_49570,N_49410);
and UO_1137 (O_1137,N_49102,N_49447);
or UO_1138 (O_1138,N_49302,N_49843);
or UO_1139 (O_1139,N_49109,N_49524);
nor UO_1140 (O_1140,N_49517,N_49000);
and UO_1141 (O_1141,N_49288,N_49684);
xor UO_1142 (O_1142,N_49300,N_49699);
nand UO_1143 (O_1143,N_49303,N_49273);
and UO_1144 (O_1144,N_49297,N_49722);
nor UO_1145 (O_1145,N_49476,N_49964);
nand UO_1146 (O_1146,N_49190,N_49788);
and UO_1147 (O_1147,N_49922,N_49458);
or UO_1148 (O_1148,N_49611,N_49191);
nand UO_1149 (O_1149,N_49572,N_49011);
and UO_1150 (O_1150,N_49976,N_49805);
nor UO_1151 (O_1151,N_49256,N_49912);
and UO_1152 (O_1152,N_49330,N_49919);
and UO_1153 (O_1153,N_49521,N_49140);
and UO_1154 (O_1154,N_49418,N_49665);
nor UO_1155 (O_1155,N_49924,N_49476);
and UO_1156 (O_1156,N_49562,N_49698);
xnor UO_1157 (O_1157,N_49939,N_49779);
xnor UO_1158 (O_1158,N_49905,N_49947);
nor UO_1159 (O_1159,N_49852,N_49353);
or UO_1160 (O_1160,N_49431,N_49750);
xor UO_1161 (O_1161,N_49882,N_49955);
or UO_1162 (O_1162,N_49004,N_49087);
and UO_1163 (O_1163,N_49492,N_49801);
nand UO_1164 (O_1164,N_49176,N_49043);
nor UO_1165 (O_1165,N_49490,N_49565);
nor UO_1166 (O_1166,N_49397,N_49297);
xor UO_1167 (O_1167,N_49027,N_49757);
xnor UO_1168 (O_1168,N_49155,N_49796);
nor UO_1169 (O_1169,N_49017,N_49929);
and UO_1170 (O_1170,N_49069,N_49878);
and UO_1171 (O_1171,N_49708,N_49236);
or UO_1172 (O_1172,N_49916,N_49828);
nand UO_1173 (O_1173,N_49904,N_49694);
and UO_1174 (O_1174,N_49246,N_49389);
nand UO_1175 (O_1175,N_49089,N_49986);
nand UO_1176 (O_1176,N_49303,N_49458);
xnor UO_1177 (O_1177,N_49444,N_49551);
and UO_1178 (O_1178,N_49441,N_49609);
nand UO_1179 (O_1179,N_49698,N_49163);
nand UO_1180 (O_1180,N_49785,N_49713);
nand UO_1181 (O_1181,N_49513,N_49305);
and UO_1182 (O_1182,N_49847,N_49324);
nand UO_1183 (O_1183,N_49033,N_49416);
xor UO_1184 (O_1184,N_49661,N_49598);
nand UO_1185 (O_1185,N_49090,N_49414);
xnor UO_1186 (O_1186,N_49161,N_49534);
xnor UO_1187 (O_1187,N_49403,N_49970);
or UO_1188 (O_1188,N_49940,N_49388);
nand UO_1189 (O_1189,N_49052,N_49236);
and UO_1190 (O_1190,N_49466,N_49099);
and UO_1191 (O_1191,N_49455,N_49580);
xor UO_1192 (O_1192,N_49748,N_49318);
and UO_1193 (O_1193,N_49444,N_49291);
or UO_1194 (O_1194,N_49617,N_49504);
nand UO_1195 (O_1195,N_49720,N_49472);
nand UO_1196 (O_1196,N_49713,N_49301);
nand UO_1197 (O_1197,N_49938,N_49810);
nor UO_1198 (O_1198,N_49092,N_49939);
nor UO_1199 (O_1199,N_49378,N_49028);
nand UO_1200 (O_1200,N_49137,N_49889);
nand UO_1201 (O_1201,N_49047,N_49598);
and UO_1202 (O_1202,N_49813,N_49834);
or UO_1203 (O_1203,N_49903,N_49515);
nand UO_1204 (O_1204,N_49888,N_49392);
nand UO_1205 (O_1205,N_49403,N_49826);
nand UO_1206 (O_1206,N_49270,N_49649);
or UO_1207 (O_1207,N_49310,N_49981);
nand UO_1208 (O_1208,N_49261,N_49061);
or UO_1209 (O_1209,N_49001,N_49274);
nor UO_1210 (O_1210,N_49994,N_49286);
nand UO_1211 (O_1211,N_49005,N_49379);
nand UO_1212 (O_1212,N_49219,N_49476);
nor UO_1213 (O_1213,N_49902,N_49928);
xor UO_1214 (O_1214,N_49874,N_49277);
or UO_1215 (O_1215,N_49993,N_49867);
nand UO_1216 (O_1216,N_49951,N_49263);
or UO_1217 (O_1217,N_49807,N_49003);
nor UO_1218 (O_1218,N_49753,N_49970);
or UO_1219 (O_1219,N_49680,N_49052);
or UO_1220 (O_1220,N_49893,N_49204);
and UO_1221 (O_1221,N_49923,N_49269);
or UO_1222 (O_1222,N_49181,N_49579);
nor UO_1223 (O_1223,N_49001,N_49083);
or UO_1224 (O_1224,N_49787,N_49854);
and UO_1225 (O_1225,N_49643,N_49559);
nand UO_1226 (O_1226,N_49825,N_49554);
or UO_1227 (O_1227,N_49252,N_49827);
nand UO_1228 (O_1228,N_49989,N_49416);
xnor UO_1229 (O_1229,N_49262,N_49241);
xnor UO_1230 (O_1230,N_49344,N_49449);
nor UO_1231 (O_1231,N_49885,N_49484);
xor UO_1232 (O_1232,N_49637,N_49950);
and UO_1233 (O_1233,N_49751,N_49698);
nand UO_1234 (O_1234,N_49405,N_49951);
nor UO_1235 (O_1235,N_49932,N_49658);
or UO_1236 (O_1236,N_49063,N_49972);
or UO_1237 (O_1237,N_49418,N_49499);
nand UO_1238 (O_1238,N_49657,N_49921);
and UO_1239 (O_1239,N_49169,N_49334);
nor UO_1240 (O_1240,N_49853,N_49625);
and UO_1241 (O_1241,N_49610,N_49725);
nand UO_1242 (O_1242,N_49692,N_49524);
nor UO_1243 (O_1243,N_49922,N_49900);
xnor UO_1244 (O_1244,N_49905,N_49026);
and UO_1245 (O_1245,N_49781,N_49747);
and UO_1246 (O_1246,N_49221,N_49052);
and UO_1247 (O_1247,N_49119,N_49756);
nor UO_1248 (O_1248,N_49303,N_49056);
and UO_1249 (O_1249,N_49209,N_49622);
nand UO_1250 (O_1250,N_49073,N_49537);
xor UO_1251 (O_1251,N_49086,N_49373);
or UO_1252 (O_1252,N_49034,N_49054);
and UO_1253 (O_1253,N_49837,N_49844);
or UO_1254 (O_1254,N_49717,N_49923);
nand UO_1255 (O_1255,N_49385,N_49335);
nand UO_1256 (O_1256,N_49951,N_49206);
or UO_1257 (O_1257,N_49076,N_49959);
xor UO_1258 (O_1258,N_49134,N_49850);
or UO_1259 (O_1259,N_49546,N_49474);
and UO_1260 (O_1260,N_49409,N_49749);
xnor UO_1261 (O_1261,N_49430,N_49144);
nor UO_1262 (O_1262,N_49924,N_49191);
nor UO_1263 (O_1263,N_49743,N_49893);
xnor UO_1264 (O_1264,N_49933,N_49454);
nand UO_1265 (O_1265,N_49557,N_49898);
nor UO_1266 (O_1266,N_49241,N_49975);
or UO_1267 (O_1267,N_49418,N_49447);
nor UO_1268 (O_1268,N_49990,N_49121);
nor UO_1269 (O_1269,N_49475,N_49476);
and UO_1270 (O_1270,N_49705,N_49616);
xnor UO_1271 (O_1271,N_49827,N_49787);
nand UO_1272 (O_1272,N_49740,N_49828);
and UO_1273 (O_1273,N_49849,N_49830);
xnor UO_1274 (O_1274,N_49530,N_49144);
or UO_1275 (O_1275,N_49348,N_49554);
nand UO_1276 (O_1276,N_49053,N_49452);
or UO_1277 (O_1277,N_49465,N_49068);
xor UO_1278 (O_1278,N_49308,N_49499);
nor UO_1279 (O_1279,N_49872,N_49463);
xor UO_1280 (O_1280,N_49130,N_49813);
nand UO_1281 (O_1281,N_49993,N_49019);
and UO_1282 (O_1282,N_49421,N_49843);
xor UO_1283 (O_1283,N_49866,N_49539);
nor UO_1284 (O_1284,N_49591,N_49085);
or UO_1285 (O_1285,N_49642,N_49022);
nand UO_1286 (O_1286,N_49274,N_49289);
or UO_1287 (O_1287,N_49213,N_49210);
and UO_1288 (O_1288,N_49148,N_49549);
nand UO_1289 (O_1289,N_49568,N_49417);
nor UO_1290 (O_1290,N_49366,N_49423);
xor UO_1291 (O_1291,N_49001,N_49951);
and UO_1292 (O_1292,N_49597,N_49928);
or UO_1293 (O_1293,N_49055,N_49866);
xnor UO_1294 (O_1294,N_49299,N_49431);
or UO_1295 (O_1295,N_49047,N_49200);
and UO_1296 (O_1296,N_49219,N_49887);
nand UO_1297 (O_1297,N_49926,N_49551);
xor UO_1298 (O_1298,N_49339,N_49033);
xnor UO_1299 (O_1299,N_49521,N_49296);
or UO_1300 (O_1300,N_49433,N_49082);
nor UO_1301 (O_1301,N_49132,N_49500);
or UO_1302 (O_1302,N_49729,N_49323);
xnor UO_1303 (O_1303,N_49701,N_49460);
nor UO_1304 (O_1304,N_49593,N_49185);
nor UO_1305 (O_1305,N_49536,N_49000);
xor UO_1306 (O_1306,N_49402,N_49718);
and UO_1307 (O_1307,N_49294,N_49820);
nand UO_1308 (O_1308,N_49164,N_49293);
nor UO_1309 (O_1309,N_49739,N_49772);
or UO_1310 (O_1310,N_49844,N_49940);
nor UO_1311 (O_1311,N_49723,N_49986);
and UO_1312 (O_1312,N_49426,N_49263);
nor UO_1313 (O_1313,N_49541,N_49426);
nand UO_1314 (O_1314,N_49158,N_49298);
or UO_1315 (O_1315,N_49959,N_49085);
or UO_1316 (O_1316,N_49289,N_49757);
and UO_1317 (O_1317,N_49875,N_49873);
and UO_1318 (O_1318,N_49825,N_49935);
nand UO_1319 (O_1319,N_49745,N_49222);
and UO_1320 (O_1320,N_49510,N_49005);
xnor UO_1321 (O_1321,N_49641,N_49040);
or UO_1322 (O_1322,N_49567,N_49560);
or UO_1323 (O_1323,N_49805,N_49898);
nor UO_1324 (O_1324,N_49182,N_49977);
nor UO_1325 (O_1325,N_49075,N_49586);
and UO_1326 (O_1326,N_49623,N_49760);
nor UO_1327 (O_1327,N_49956,N_49883);
and UO_1328 (O_1328,N_49562,N_49442);
nor UO_1329 (O_1329,N_49464,N_49966);
nor UO_1330 (O_1330,N_49963,N_49294);
or UO_1331 (O_1331,N_49283,N_49041);
or UO_1332 (O_1332,N_49517,N_49506);
xor UO_1333 (O_1333,N_49822,N_49290);
or UO_1334 (O_1334,N_49446,N_49241);
xor UO_1335 (O_1335,N_49554,N_49549);
xnor UO_1336 (O_1336,N_49684,N_49307);
nand UO_1337 (O_1337,N_49415,N_49641);
or UO_1338 (O_1338,N_49772,N_49063);
nand UO_1339 (O_1339,N_49232,N_49871);
xor UO_1340 (O_1340,N_49360,N_49463);
xnor UO_1341 (O_1341,N_49853,N_49863);
and UO_1342 (O_1342,N_49928,N_49819);
and UO_1343 (O_1343,N_49656,N_49140);
or UO_1344 (O_1344,N_49597,N_49876);
nor UO_1345 (O_1345,N_49903,N_49372);
xor UO_1346 (O_1346,N_49663,N_49471);
xor UO_1347 (O_1347,N_49530,N_49003);
or UO_1348 (O_1348,N_49443,N_49726);
xor UO_1349 (O_1349,N_49341,N_49269);
or UO_1350 (O_1350,N_49324,N_49849);
nor UO_1351 (O_1351,N_49317,N_49420);
or UO_1352 (O_1352,N_49321,N_49627);
nor UO_1353 (O_1353,N_49912,N_49876);
nand UO_1354 (O_1354,N_49051,N_49780);
nor UO_1355 (O_1355,N_49070,N_49563);
nor UO_1356 (O_1356,N_49521,N_49697);
xnor UO_1357 (O_1357,N_49057,N_49078);
and UO_1358 (O_1358,N_49409,N_49717);
nand UO_1359 (O_1359,N_49186,N_49851);
and UO_1360 (O_1360,N_49214,N_49488);
nand UO_1361 (O_1361,N_49614,N_49346);
xor UO_1362 (O_1362,N_49435,N_49228);
nor UO_1363 (O_1363,N_49764,N_49963);
nor UO_1364 (O_1364,N_49627,N_49643);
nor UO_1365 (O_1365,N_49994,N_49096);
and UO_1366 (O_1366,N_49479,N_49630);
or UO_1367 (O_1367,N_49397,N_49725);
nand UO_1368 (O_1368,N_49615,N_49019);
and UO_1369 (O_1369,N_49105,N_49349);
or UO_1370 (O_1370,N_49890,N_49065);
nor UO_1371 (O_1371,N_49069,N_49148);
nor UO_1372 (O_1372,N_49289,N_49893);
and UO_1373 (O_1373,N_49233,N_49206);
xor UO_1374 (O_1374,N_49168,N_49617);
xnor UO_1375 (O_1375,N_49791,N_49278);
xnor UO_1376 (O_1376,N_49461,N_49394);
xnor UO_1377 (O_1377,N_49215,N_49824);
and UO_1378 (O_1378,N_49451,N_49637);
xor UO_1379 (O_1379,N_49800,N_49144);
xnor UO_1380 (O_1380,N_49451,N_49391);
and UO_1381 (O_1381,N_49991,N_49928);
nor UO_1382 (O_1382,N_49793,N_49675);
nor UO_1383 (O_1383,N_49456,N_49825);
and UO_1384 (O_1384,N_49035,N_49665);
or UO_1385 (O_1385,N_49093,N_49481);
or UO_1386 (O_1386,N_49416,N_49599);
xnor UO_1387 (O_1387,N_49992,N_49034);
or UO_1388 (O_1388,N_49772,N_49562);
xor UO_1389 (O_1389,N_49750,N_49722);
or UO_1390 (O_1390,N_49352,N_49303);
xor UO_1391 (O_1391,N_49944,N_49262);
nand UO_1392 (O_1392,N_49562,N_49742);
xnor UO_1393 (O_1393,N_49563,N_49424);
and UO_1394 (O_1394,N_49766,N_49940);
xor UO_1395 (O_1395,N_49426,N_49813);
or UO_1396 (O_1396,N_49855,N_49561);
and UO_1397 (O_1397,N_49595,N_49311);
xnor UO_1398 (O_1398,N_49416,N_49287);
or UO_1399 (O_1399,N_49005,N_49513);
and UO_1400 (O_1400,N_49046,N_49809);
or UO_1401 (O_1401,N_49897,N_49445);
and UO_1402 (O_1402,N_49041,N_49185);
xnor UO_1403 (O_1403,N_49196,N_49727);
or UO_1404 (O_1404,N_49882,N_49700);
xor UO_1405 (O_1405,N_49855,N_49132);
nor UO_1406 (O_1406,N_49485,N_49249);
xor UO_1407 (O_1407,N_49619,N_49442);
or UO_1408 (O_1408,N_49359,N_49312);
xnor UO_1409 (O_1409,N_49439,N_49676);
xnor UO_1410 (O_1410,N_49596,N_49379);
xor UO_1411 (O_1411,N_49312,N_49357);
xor UO_1412 (O_1412,N_49123,N_49124);
xor UO_1413 (O_1413,N_49493,N_49211);
and UO_1414 (O_1414,N_49131,N_49476);
and UO_1415 (O_1415,N_49650,N_49969);
nand UO_1416 (O_1416,N_49237,N_49275);
or UO_1417 (O_1417,N_49170,N_49256);
xnor UO_1418 (O_1418,N_49895,N_49474);
nor UO_1419 (O_1419,N_49170,N_49974);
and UO_1420 (O_1420,N_49751,N_49747);
and UO_1421 (O_1421,N_49352,N_49085);
or UO_1422 (O_1422,N_49997,N_49915);
nand UO_1423 (O_1423,N_49112,N_49298);
nand UO_1424 (O_1424,N_49042,N_49205);
and UO_1425 (O_1425,N_49546,N_49460);
xnor UO_1426 (O_1426,N_49098,N_49993);
or UO_1427 (O_1427,N_49809,N_49724);
or UO_1428 (O_1428,N_49657,N_49895);
nand UO_1429 (O_1429,N_49847,N_49976);
nand UO_1430 (O_1430,N_49267,N_49556);
or UO_1431 (O_1431,N_49965,N_49194);
and UO_1432 (O_1432,N_49016,N_49857);
xor UO_1433 (O_1433,N_49096,N_49116);
nand UO_1434 (O_1434,N_49769,N_49778);
and UO_1435 (O_1435,N_49696,N_49626);
xor UO_1436 (O_1436,N_49145,N_49865);
nand UO_1437 (O_1437,N_49592,N_49648);
nand UO_1438 (O_1438,N_49372,N_49234);
and UO_1439 (O_1439,N_49977,N_49597);
nand UO_1440 (O_1440,N_49956,N_49103);
nor UO_1441 (O_1441,N_49593,N_49192);
or UO_1442 (O_1442,N_49137,N_49491);
xor UO_1443 (O_1443,N_49935,N_49080);
and UO_1444 (O_1444,N_49409,N_49996);
nor UO_1445 (O_1445,N_49796,N_49464);
nand UO_1446 (O_1446,N_49077,N_49668);
nor UO_1447 (O_1447,N_49882,N_49330);
nor UO_1448 (O_1448,N_49562,N_49855);
or UO_1449 (O_1449,N_49244,N_49369);
or UO_1450 (O_1450,N_49301,N_49904);
and UO_1451 (O_1451,N_49365,N_49024);
xnor UO_1452 (O_1452,N_49925,N_49373);
nand UO_1453 (O_1453,N_49423,N_49900);
xnor UO_1454 (O_1454,N_49218,N_49651);
and UO_1455 (O_1455,N_49831,N_49173);
xnor UO_1456 (O_1456,N_49979,N_49837);
or UO_1457 (O_1457,N_49652,N_49169);
and UO_1458 (O_1458,N_49519,N_49784);
or UO_1459 (O_1459,N_49851,N_49374);
nand UO_1460 (O_1460,N_49657,N_49065);
or UO_1461 (O_1461,N_49972,N_49888);
nand UO_1462 (O_1462,N_49557,N_49704);
and UO_1463 (O_1463,N_49876,N_49672);
or UO_1464 (O_1464,N_49397,N_49323);
nand UO_1465 (O_1465,N_49146,N_49168);
nor UO_1466 (O_1466,N_49215,N_49172);
or UO_1467 (O_1467,N_49218,N_49560);
nand UO_1468 (O_1468,N_49589,N_49609);
nor UO_1469 (O_1469,N_49796,N_49613);
and UO_1470 (O_1470,N_49100,N_49829);
and UO_1471 (O_1471,N_49158,N_49525);
or UO_1472 (O_1472,N_49158,N_49035);
nand UO_1473 (O_1473,N_49586,N_49449);
nor UO_1474 (O_1474,N_49209,N_49474);
and UO_1475 (O_1475,N_49097,N_49085);
nand UO_1476 (O_1476,N_49955,N_49956);
and UO_1477 (O_1477,N_49875,N_49151);
nand UO_1478 (O_1478,N_49343,N_49329);
nor UO_1479 (O_1479,N_49596,N_49207);
xnor UO_1480 (O_1480,N_49242,N_49566);
nor UO_1481 (O_1481,N_49301,N_49710);
nor UO_1482 (O_1482,N_49251,N_49044);
and UO_1483 (O_1483,N_49194,N_49778);
nor UO_1484 (O_1484,N_49384,N_49071);
xnor UO_1485 (O_1485,N_49743,N_49261);
xnor UO_1486 (O_1486,N_49209,N_49752);
nor UO_1487 (O_1487,N_49672,N_49080);
nor UO_1488 (O_1488,N_49585,N_49580);
nor UO_1489 (O_1489,N_49719,N_49906);
and UO_1490 (O_1490,N_49492,N_49104);
or UO_1491 (O_1491,N_49452,N_49453);
xnor UO_1492 (O_1492,N_49871,N_49281);
nor UO_1493 (O_1493,N_49995,N_49056);
nor UO_1494 (O_1494,N_49373,N_49922);
and UO_1495 (O_1495,N_49211,N_49285);
nor UO_1496 (O_1496,N_49033,N_49834);
nor UO_1497 (O_1497,N_49410,N_49812);
nor UO_1498 (O_1498,N_49294,N_49596);
and UO_1499 (O_1499,N_49424,N_49734);
xor UO_1500 (O_1500,N_49802,N_49946);
or UO_1501 (O_1501,N_49521,N_49082);
or UO_1502 (O_1502,N_49057,N_49298);
nand UO_1503 (O_1503,N_49974,N_49377);
and UO_1504 (O_1504,N_49151,N_49806);
and UO_1505 (O_1505,N_49531,N_49608);
nand UO_1506 (O_1506,N_49533,N_49940);
nand UO_1507 (O_1507,N_49668,N_49570);
or UO_1508 (O_1508,N_49931,N_49294);
or UO_1509 (O_1509,N_49355,N_49541);
nand UO_1510 (O_1510,N_49585,N_49722);
or UO_1511 (O_1511,N_49329,N_49165);
and UO_1512 (O_1512,N_49559,N_49635);
and UO_1513 (O_1513,N_49582,N_49006);
and UO_1514 (O_1514,N_49250,N_49196);
nor UO_1515 (O_1515,N_49787,N_49045);
and UO_1516 (O_1516,N_49628,N_49556);
and UO_1517 (O_1517,N_49462,N_49360);
nor UO_1518 (O_1518,N_49181,N_49381);
and UO_1519 (O_1519,N_49612,N_49276);
or UO_1520 (O_1520,N_49776,N_49289);
xnor UO_1521 (O_1521,N_49522,N_49321);
and UO_1522 (O_1522,N_49670,N_49004);
or UO_1523 (O_1523,N_49284,N_49923);
xor UO_1524 (O_1524,N_49928,N_49507);
and UO_1525 (O_1525,N_49901,N_49528);
nand UO_1526 (O_1526,N_49478,N_49360);
xnor UO_1527 (O_1527,N_49521,N_49547);
nand UO_1528 (O_1528,N_49493,N_49391);
nor UO_1529 (O_1529,N_49192,N_49805);
xor UO_1530 (O_1530,N_49773,N_49917);
nand UO_1531 (O_1531,N_49527,N_49392);
nor UO_1532 (O_1532,N_49287,N_49186);
and UO_1533 (O_1533,N_49874,N_49141);
nand UO_1534 (O_1534,N_49885,N_49328);
nand UO_1535 (O_1535,N_49913,N_49463);
or UO_1536 (O_1536,N_49978,N_49892);
nor UO_1537 (O_1537,N_49810,N_49054);
xor UO_1538 (O_1538,N_49676,N_49616);
xnor UO_1539 (O_1539,N_49438,N_49182);
or UO_1540 (O_1540,N_49163,N_49379);
or UO_1541 (O_1541,N_49479,N_49090);
nor UO_1542 (O_1542,N_49514,N_49912);
or UO_1543 (O_1543,N_49072,N_49631);
nor UO_1544 (O_1544,N_49211,N_49844);
nand UO_1545 (O_1545,N_49483,N_49846);
nand UO_1546 (O_1546,N_49325,N_49805);
and UO_1547 (O_1547,N_49607,N_49736);
nor UO_1548 (O_1548,N_49406,N_49775);
nor UO_1549 (O_1549,N_49712,N_49094);
or UO_1550 (O_1550,N_49699,N_49786);
nor UO_1551 (O_1551,N_49428,N_49892);
xor UO_1552 (O_1552,N_49892,N_49777);
or UO_1553 (O_1553,N_49583,N_49569);
or UO_1554 (O_1554,N_49270,N_49983);
nand UO_1555 (O_1555,N_49649,N_49444);
and UO_1556 (O_1556,N_49874,N_49628);
and UO_1557 (O_1557,N_49444,N_49199);
or UO_1558 (O_1558,N_49086,N_49663);
xnor UO_1559 (O_1559,N_49762,N_49094);
xnor UO_1560 (O_1560,N_49681,N_49195);
nor UO_1561 (O_1561,N_49508,N_49487);
or UO_1562 (O_1562,N_49108,N_49549);
xor UO_1563 (O_1563,N_49019,N_49566);
nand UO_1564 (O_1564,N_49645,N_49333);
and UO_1565 (O_1565,N_49123,N_49569);
nand UO_1566 (O_1566,N_49040,N_49959);
or UO_1567 (O_1567,N_49894,N_49294);
nor UO_1568 (O_1568,N_49097,N_49719);
or UO_1569 (O_1569,N_49885,N_49931);
or UO_1570 (O_1570,N_49590,N_49064);
and UO_1571 (O_1571,N_49281,N_49674);
or UO_1572 (O_1572,N_49863,N_49802);
xor UO_1573 (O_1573,N_49719,N_49371);
nand UO_1574 (O_1574,N_49333,N_49093);
xnor UO_1575 (O_1575,N_49019,N_49126);
and UO_1576 (O_1576,N_49973,N_49335);
nand UO_1577 (O_1577,N_49329,N_49727);
nor UO_1578 (O_1578,N_49968,N_49173);
or UO_1579 (O_1579,N_49523,N_49408);
and UO_1580 (O_1580,N_49533,N_49253);
or UO_1581 (O_1581,N_49541,N_49199);
nand UO_1582 (O_1582,N_49597,N_49493);
or UO_1583 (O_1583,N_49487,N_49420);
nand UO_1584 (O_1584,N_49786,N_49429);
nand UO_1585 (O_1585,N_49645,N_49897);
and UO_1586 (O_1586,N_49965,N_49705);
and UO_1587 (O_1587,N_49670,N_49597);
nor UO_1588 (O_1588,N_49402,N_49850);
nand UO_1589 (O_1589,N_49659,N_49155);
or UO_1590 (O_1590,N_49510,N_49025);
xnor UO_1591 (O_1591,N_49644,N_49978);
nor UO_1592 (O_1592,N_49271,N_49043);
or UO_1593 (O_1593,N_49171,N_49593);
nand UO_1594 (O_1594,N_49761,N_49499);
or UO_1595 (O_1595,N_49848,N_49302);
nor UO_1596 (O_1596,N_49613,N_49805);
nand UO_1597 (O_1597,N_49690,N_49233);
nor UO_1598 (O_1598,N_49717,N_49201);
or UO_1599 (O_1599,N_49322,N_49855);
nor UO_1600 (O_1600,N_49652,N_49139);
nand UO_1601 (O_1601,N_49258,N_49690);
nor UO_1602 (O_1602,N_49426,N_49290);
nor UO_1603 (O_1603,N_49772,N_49910);
or UO_1604 (O_1604,N_49563,N_49912);
xor UO_1605 (O_1605,N_49174,N_49685);
and UO_1606 (O_1606,N_49507,N_49496);
nand UO_1607 (O_1607,N_49750,N_49402);
or UO_1608 (O_1608,N_49693,N_49240);
xor UO_1609 (O_1609,N_49597,N_49771);
or UO_1610 (O_1610,N_49022,N_49922);
or UO_1611 (O_1611,N_49047,N_49345);
xnor UO_1612 (O_1612,N_49048,N_49743);
nor UO_1613 (O_1613,N_49186,N_49084);
or UO_1614 (O_1614,N_49378,N_49700);
nor UO_1615 (O_1615,N_49696,N_49079);
or UO_1616 (O_1616,N_49453,N_49384);
nand UO_1617 (O_1617,N_49946,N_49539);
and UO_1618 (O_1618,N_49070,N_49229);
nor UO_1619 (O_1619,N_49392,N_49971);
or UO_1620 (O_1620,N_49595,N_49236);
or UO_1621 (O_1621,N_49692,N_49070);
nor UO_1622 (O_1622,N_49087,N_49964);
or UO_1623 (O_1623,N_49744,N_49538);
nand UO_1624 (O_1624,N_49948,N_49802);
xor UO_1625 (O_1625,N_49418,N_49022);
nor UO_1626 (O_1626,N_49395,N_49290);
nand UO_1627 (O_1627,N_49358,N_49482);
xor UO_1628 (O_1628,N_49173,N_49323);
nor UO_1629 (O_1629,N_49288,N_49031);
xor UO_1630 (O_1630,N_49773,N_49273);
or UO_1631 (O_1631,N_49029,N_49538);
and UO_1632 (O_1632,N_49417,N_49027);
or UO_1633 (O_1633,N_49413,N_49706);
nand UO_1634 (O_1634,N_49138,N_49179);
xnor UO_1635 (O_1635,N_49337,N_49349);
and UO_1636 (O_1636,N_49977,N_49719);
xor UO_1637 (O_1637,N_49473,N_49075);
or UO_1638 (O_1638,N_49908,N_49988);
and UO_1639 (O_1639,N_49567,N_49955);
xor UO_1640 (O_1640,N_49906,N_49712);
xor UO_1641 (O_1641,N_49728,N_49256);
and UO_1642 (O_1642,N_49453,N_49331);
nor UO_1643 (O_1643,N_49236,N_49969);
nor UO_1644 (O_1644,N_49060,N_49819);
nand UO_1645 (O_1645,N_49800,N_49325);
nand UO_1646 (O_1646,N_49227,N_49906);
xor UO_1647 (O_1647,N_49397,N_49887);
and UO_1648 (O_1648,N_49955,N_49487);
and UO_1649 (O_1649,N_49544,N_49739);
nand UO_1650 (O_1650,N_49774,N_49028);
and UO_1651 (O_1651,N_49499,N_49076);
nand UO_1652 (O_1652,N_49791,N_49472);
nand UO_1653 (O_1653,N_49767,N_49831);
nor UO_1654 (O_1654,N_49275,N_49160);
nor UO_1655 (O_1655,N_49765,N_49659);
nand UO_1656 (O_1656,N_49688,N_49531);
nor UO_1657 (O_1657,N_49081,N_49148);
and UO_1658 (O_1658,N_49438,N_49461);
and UO_1659 (O_1659,N_49596,N_49310);
and UO_1660 (O_1660,N_49196,N_49688);
or UO_1661 (O_1661,N_49253,N_49148);
nand UO_1662 (O_1662,N_49521,N_49827);
and UO_1663 (O_1663,N_49103,N_49638);
nor UO_1664 (O_1664,N_49486,N_49130);
and UO_1665 (O_1665,N_49336,N_49090);
or UO_1666 (O_1666,N_49321,N_49137);
nand UO_1667 (O_1667,N_49761,N_49926);
nor UO_1668 (O_1668,N_49822,N_49793);
nor UO_1669 (O_1669,N_49811,N_49587);
xor UO_1670 (O_1670,N_49516,N_49774);
nor UO_1671 (O_1671,N_49549,N_49029);
nand UO_1672 (O_1672,N_49613,N_49677);
xor UO_1673 (O_1673,N_49734,N_49965);
or UO_1674 (O_1674,N_49208,N_49503);
nor UO_1675 (O_1675,N_49855,N_49483);
or UO_1676 (O_1676,N_49823,N_49134);
xnor UO_1677 (O_1677,N_49972,N_49146);
nor UO_1678 (O_1678,N_49491,N_49772);
or UO_1679 (O_1679,N_49287,N_49627);
xnor UO_1680 (O_1680,N_49986,N_49810);
or UO_1681 (O_1681,N_49555,N_49387);
or UO_1682 (O_1682,N_49083,N_49420);
xnor UO_1683 (O_1683,N_49208,N_49144);
nand UO_1684 (O_1684,N_49087,N_49310);
nand UO_1685 (O_1685,N_49772,N_49849);
nand UO_1686 (O_1686,N_49282,N_49549);
nor UO_1687 (O_1687,N_49858,N_49724);
nor UO_1688 (O_1688,N_49529,N_49356);
or UO_1689 (O_1689,N_49438,N_49305);
nor UO_1690 (O_1690,N_49931,N_49445);
xor UO_1691 (O_1691,N_49937,N_49163);
or UO_1692 (O_1692,N_49395,N_49348);
or UO_1693 (O_1693,N_49504,N_49871);
or UO_1694 (O_1694,N_49033,N_49327);
and UO_1695 (O_1695,N_49690,N_49165);
and UO_1696 (O_1696,N_49715,N_49291);
or UO_1697 (O_1697,N_49102,N_49463);
and UO_1698 (O_1698,N_49566,N_49069);
nor UO_1699 (O_1699,N_49561,N_49206);
nor UO_1700 (O_1700,N_49260,N_49406);
xor UO_1701 (O_1701,N_49877,N_49573);
xnor UO_1702 (O_1702,N_49273,N_49715);
nand UO_1703 (O_1703,N_49941,N_49673);
and UO_1704 (O_1704,N_49153,N_49966);
or UO_1705 (O_1705,N_49691,N_49952);
and UO_1706 (O_1706,N_49982,N_49984);
nand UO_1707 (O_1707,N_49998,N_49687);
nor UO_1708 (O_1708,N_49827,N_49032);
and UO_1709 (O_1709,N_49139,N_49205);
nor UO_1710 (O_1710,N_49351,N_49901);
and UO_1711 (O_1711,N_49636,N_49176);
nand UO_1712 (O_1712,N_49449,N_49699);
and UO_1713 (O_1713,N_49423,N_49870);
nor UO_1714 (O_1714,N_49914,N_49574);
nor UO_1715 (O_1715,N_49665,N_49198);
and UO_1716 (O_1716,N_49646,N_49187);
nand UO_1717 (O_1717,N_49841,N_49888);
and UO_1718 (O_1718,N_49483,N_49269);
and UO_1719 (O_1719,N_49215,N_49008);
xnor UO_1720 (O_1720,N_49156,N_49442);
nor UO_1721 (O_1721,N_49732,N_49120);
nand UO_1722 (O_1722,N_49971,N_49619);
nor UO_1723 (O_1723,N_49289,N_49783);
and UO_1724 (O_1724,N_49843,N_49269);
nor UO_1725 (O_1725,N_49351,N_49414);
or UO_1726 (O_1726,N_49183,N_49289);
nand UO_1727 (O_1727,N_49479,N_49553);
or UO_1728 (O_1728,N_49250,N_49461);
xnor UO_1729 (O_1729,N_49632,N_49230);
nor UO_1730 (O_1730,N_49312,N_49899);
nor UO_1731 (O_1731,N_49618,N_49381);
xnor UO_1732 (O_1732,N_49558,N_49645);
or UO_1733 (O_1733,N_49448,N_49160);
xor UO_1734 (O_1734,N_49927,N_49716);
nand UO_1735 (O_1735,N_49496,N_49971);
nand UO_1736 (O_1736,N_49399,N_49544);
xor UO_1737 (O_1737,N_49989,N_49315);
nor UO_1738 (O_1738,N_49993,N_49155);
xor UO_1739 (O_1739,N_49145,N_49354);
nor UO_1740 (O_1740,N_49824,N_49631);
nand UO_1741 (O_1741,N_49360,N_49258);
or UO_1742 (O_1742,N_49364,N_49959);
nor UO_1743 (O_1743,N_49341,N_49095);
or UO_1744 (O_1744,N_49341,N_49604);
nand UO_1745 (O_1745,N_49645,N_49059);
and UO_1746 (O_1746,N_49431,N_49781);
nand UO_1747 (O_1747,N_49461,N_49686);
or UO_1748 (O_1748,N_49904,N_49952);
nor UO_1749 (O_1749,N_49762,N_49662);
and UO_1750 (O_1750,N_49129,N_49765);
or UO_1751 (O_1751,N_49939,N_49727);
xnor UO_1752 (O_1752,N_49099,N_49255);
or UO_1753 (O_1753,N_49231,N_49863);
or UO_1754 (O_1754,N_49903,N_49234);
xor UO_1755 (O_1755,N_49903,N_49376);
or UO_1756 (O_1756,N_49273,N_49146);
and UO_1757 (O_1757,N_49052,N_49379);
nor UO_1758 (O_1758,N_49871,N_49307);
xor UO_1759 (O_1759,N_49601,N_49883);
nor UO_1760 (O_1760,N_49260,N_49367);
or UO_1761 (O_1761,N_49447,N_49467);
nand UO_1762 (O_1762,N_49421,N_49521);
or UO_1763 (O_1763,N_49958,N_49449);
and UO_1764 (O_1764,N_49522,N_49606);
or UO_1765 (O_1765,N_49974,N_49762);
nand UO_1766 (O_1766,N_49707,N_49585);
or UO_1767 (O_1767,N_49942,N_49886);
or UO_1768 (O_1768,N_49753,N_49536);
or UO_1769 (O_1769,N_49462,N_49995);
nor UO_1770 (O_1770,N_49338,N_49236);
or UO_1771 (O_1771,N_49618,N_49363);
nor UO_1772 (O_1772,N_49409,N_49391);
or UO_1773 (O_1773,N_49233,N_49041);
nand UO_1774 (O_1774,N_49593,N_49912);
nor UO_1775 (O_1775,N_49904,N_49938);
and UO_1776 (O_1776,N_49412,N_49400);
nand UO_1777 (O_1777,N_49724,N_49175);
or UO_1778 (O_1778,N_49753,N_49229);
and UO_1779 (O_1779,N_49794,N_49695);
xor UO_1780 (O_1780,N_49420,N_49992);
or UO_1781 (O_1781,N_49406,N_49548);
nor UO_1782 (O_1782,N_49502,N_49486);
nor UO_1783 (O_1783,N_49527,N_49157);
nor UO_1784 (O_1784,N_49375,N_49212);
nand UO_1785 (O_1785,N_49945,N_49068);
nor UO_1786 (O_1786,N_49249,N_49088);
or UO_1787 (O_1787,N_49379,N_49745);
xnor UO_1788 (O_1788,N_49227,N_49223);
nand UO_1789 (O_1789,N_49823,N_49625);
and UO_1790 (O_1790,N_49843,N_49771);
and UO_1791 (O_1791,N_49057,N_49329);
or UO_1792 (O_1792,N_49592,N_49060);
xnor UO_1793 (O_1793,N_49583,N_49670);
or UO_1794 (O_1794,N_49050,N_49588);
xor UO_1795 (O_1795,N_49405,N_49535);
and UO_1796 (O_1796,N_49025,N_49741);
or UO_1797 (O_1797,N_49667,N_49342);
or UO_1798 (O_1798,N_49525,N_49229);
and UO_1799 (O_1799,N_49984,N_49763);
xor UO_1800 (O_1800,N_49570,N_49327);
nand UO_1801 (O_1801,N_49862,N_49856);
nor UO_1802 (O_1802,N_49441,N_49020);
and UO_1803 (O_1803,N_49071,N_49902);
or UO_1804 (O_1804,N_49925,N_49165);
nand UO_1805 (O_1805,N_49442,N_49009);
nor UO_1806 (O_1806,N_49653,N_49168);
nand UO_1807 (O_1807,N_49298,N_49704);
xnor UO_1808 (O_1808,N_49306,N_49704);
or UO_1809 (O_1809,N_49185,N_49642);
and UO_1810 (O_1810,N_49479,N_49374);
xor UO_1811 (O_1811,N_49973,N_49182);
or UO_1812 (O_1812,N_49855,N_49548);
and UO_1813 (O_1813,N_49197,N_49916);
xor UO_1814 (O_1814,N_49098,N_49770);
or UO_1815 (O_1815,N_49899,N_49104);
and UO_1816 (O_1816,N_49831,N_49764);
nor UO_1817 (O_1817,N_49352,N_49451);
xnor UO_1818 (O_1818,N_49529,N_49905);
or UO_1819 (O_1819,N_49939,N_49716);
nand UO_1820 (O_1820,N_49415,N_49029);
and UO_1821 (O_1821,N_49133,N_49573);
xor UO_1822 (O_1822,N_49740,N_49328);
xnor UO_1823 (O_1823,N_49540,N_49561);
nor UO_1824 (O_1824,N_49721,N_49068);
xnor UO_1825 (O_1825,N_49928,N_49731);
and UO_1826 (O_1826,N_49961,N_49325);
nor UO_1827 (O_1827,N_49312,N_49716);
and UO_1828 (O_1828,N_49879,N_49443);
and UO_1829 (O_1829,N_49050,N_49699);
and UO_1830 (O_1830,N_49687,N_49159);
nand UO_1831 (O_1831,N_49368,N_49365);
nor UO_1832 (O_1832,N_49993,N_49506);
or UO_1833 (O_1833,N_49976,N_49418);
and UO_1834 (O_1834,N_49899,N_49064);
or UO_1835 (O_1835,N_49431,N_49416);
and UO_1836 (O_1836,N_49156,N_49527);
xor UO_1837 (O_1837,N_49654,N_49549);
nand UO_1838 (O_1838,N_49491,N_49473);
nor UO_1839 (O_1839,N_49166,N_49663);
or UO_1840 (O_1840,N_49057,N_49188);
xor UO_1841 (O_1841,N_49966,N_49288);
xnor UO_1842 (O_1842,N_49690,N_49666);
or UO_1843 (O_1843,N_49249,N_49070);
xor UO_1844 (O_1844,N_49762,N_49307);
and UO_1845 (O_1845,N_49897,N_49098);
nor UO_1846 (O_1846,N_49590,N_49134);
and UO_1847 (O_1847,N_49949,N_49619);
and UO_1848 (O_1848,N_49728,N_49243);
nor UO_1849 (O_1849,N_49769,N_49406);
and UO_1850 (O_1850,N_49373,N_49718);
nor UO_1851 (O_1851,N_49359,N_49551);
or UO_1852 (O_1852,N_49856,N_49545);
or UO_1853 (O_1853,N_49898,N_49985);
xor UO_1854 (O_1854,N_49290,N_49792);
nand UO_1855 (O_1855,N_49185,N_49823);
or UO_1856 (O_1856,N_49871,N_49446);
nor UO_1857 (O_1857,N_49084,N_49163);
xnor UO_1858 (O_1858,N_49393,N_49163);
nor UO_1859 (O_1859,N_49951,N_49119);
nor UO_1860 (O_1860,N_49963,N_49037);
or UO_1861 (O_1861,N_49580,N_49676);
or UO_1862 (O_1862,N_49323,N_49675);
nand UO_1863 (O_1863,N_49962,N_49230);
xor UO_1864 (O_1864,N_49894,N_49321);
and UO_1865 (O_1865,N_49549,N_49379);
nand UO_1866 (O_1866,N_49681,N_49755);
xnor UO_1867 (O_1867,N_49405,N_49087);
nor UO_1868 (O_1868,N_49426,N_49456);
or UO_1869 (O_1869,N_49105,N_49297);
nand UO_1870 (O_1870,N_49533,N_49218);
xor UO_1871 (O_1871,N_49539,N_49175);
xor UO_1872 (O_1872,N_49050,N_49744);
xor UO_1873 (O_1873,N_49810,N_49410);
nand UO_1874 (O_1874,N_49816,N_49666);
nand UO_1875 (O_1875,N_49761,N_49850);
nand UO_1876 (O_1876,N_49643,N_49404);
nand UO_1877 (O_1877,N_49175,N_49561);
nand UO_1878 (O_1878,N_49145,N_49727);
nor UO_1879 (O_1879,N_49882,N_49821);
xnor UO_1880 (O_1880,N_49362,N_49402);
and UO_1881 (O_1881,N_49714,N_49215);
and UO_1882 (O_1882,N_49696,N_49588);
nand UO_1883 (O_1883,N_49504,N_49578);
or UO_1884 (O_1884,N_49428,N_49317);
nor UO_1885 (O_1885,N_49983,N_49151);
nor UO_1886 (O_1886,N_49031,N_49752);
xnor UO_1887 (O_1887,N_49055,N_49674);
nor UO_1888 (O_1888,N_49726,N_49696);
xor UO_1889 (O_1889,N_49194,N_49935);
nand UO_1890 (O_1890,N_49321,N_49593);
and UO_1891 (O_1891,N_49055,N_49108);
nor UO_1892 (O_1892,N_49999,N_49063);
or UO_1893 (O_1893,N_49272,N_49898);
or UO_1894 (O_1894,N_49891,N_49166);
xor UO_1895 (O_1895,N_49557,N_49607);
and UO_1896 (O_1896,N_49691,N_49507);
xnor UO_1897 (O_1897,N_49248,N_49112);
nand UO_1898 (O_1898,N_49589,N_49008);
and UO_1899 (O_1899,N_49298,N_49432);
nand UO_1900 (O_1900,N_49244,N_49409);
nor UO_1901 (O_1901,N_49834,N_49381);
or UO_1902 (O_1902,N_49985,N_49559);
nor UO_1903 (O_1903,N_49216,N_49343);
or UO_1904 (O_1904,N_49100,N_49802);
nand UO_1905 (O_1905,N_49331,N_49533);
nand UO_1906 (O_1906,N_49414,N_49042);
nor UO_1907 (O_1907,N_49808,N_49446);
xnor UO_1908 (O_1908,N_49757,N_49252);
xnor UO_1909 (O_1909,N_49879,N_49945);
or UO_1910 (O_1910,N_49598,N_49328);
xor UO_1911 (O_1911,N_49309,N_49915);
nor UO_1912 (O_1912,N_49783,N_49192);
nand UO_1913 (O_1913,N_49500,N_49797);
xor UO_1914 (O_1914,N_49163,N_49353);
nand UO_1915 (O_1915,N_49493,N_49928);
xnor UO_1916 (O_1916,N_49873,N_49572);
xnor UO_1917 (O_1917,N_49011,N_49118);
nand UO_1918 (O_1918,N_49372,N_49248);
nor UO_1919 (O_1919,N_49951,N_49893);
xor UO_1920 (O_1920,N_49533,N_49130);
nand UO_1921 (O_1921,N_49329,N_49050);
or UO_1922 (O_1922,N_49217,N_49297);
xor UO_1923 (O_1923,N_49912,N_49629);
nor UO_1924 (O_1924,N_49580,N_49678);
nor UO_1925 (O_1925,N_49986,N_49027);
nand UO_1926 (O_1926,N_49805,N_49962);
or UO_1927 (O_1927,N_49316,N_49273);
nor UO_1928 (O_1928,N_49954,N_49869);
and UO_1929 (O_1929,N_49508,N_49517);
nand UO_1930 (O_1930,N_49062,N_49095);
and UO_1931 (O_1931,N_49294,N_49667);
nor UO_1932 (O_1932,N_49544,N_49947);
or UO_1933 (O_1933,N_49593,N_49488);
and UO_1934 (O_1934,N_49454,N_49364);
xnor UO_1935 (O_1935,N_49825,N_49211);
xnor UO_1936 (O_1936,N_49045,N_49219);
or UO_1937 (O_1937,N_49972,N_49376);
and UO_1938 (O_1938,N_49272,N_49089);
nand UO_1939 (O_1939,N_49986,N_49140);
nor UO_1940 (O_1940,N_49058,N_49637);
or UO_1941 (O_1941,N_49731,N_49192);
or UO_1942 (O_1942,N_49295,N_49826);
xor UO_1943 (O_1943,N_49111,N_49699);
xor UO_1944 (O_1944,N_49029,N_49790);
nand UO_1945 (O_1945,N_49980,N_49361);
and UO_1946 (O_1946,N_49095,N_49843);
or UO_1947 (O_1947,N_49071,N_49745);
or UO_1948 (O_1948,N_49123,N_49580);
or UO_1949 (O_1949,N_49639,N_49385);
xor UO_1950 (O_1950,N_49086,N_49080);
nand UO_1951 (O_1951,N_49978,N_49656);
nor UO_1952 (O_1952,N_49430,N_49526);
and UO_1953 (O_1953,N_49244,N_49258);
and UO_1954 (O_1954,N_49816,N_49607);
nor UO_1955 (O_1955,N_49665,N_49924);
or UO_1956 (O_1956,N_49736,N_49438);
xor UO_1957 (O_1957,N_49589,N_49245);
or UO_1958 (O_1958,N_49880,N_49335);
xor UO_1959 (O_1959,N_49539,N_49396);
xor UO_1960 (O_1960,N_49984,N_49527);
or UO_1961 (O_1961,N_49672,N_49950);
nor UO_1962 (O_1962,N_49172,N_49539);
xnor UO_1963 (O_1963,N_49124,N_49892);
nand UO_1964 (O_1964,N_49460,N_49255);
xor UO_1965 (O_1965,N_49526,N_49058);
or UO_1966 (O_1966,N_49735,N_49601);
and UO_1967 (O_1967,N_49261,N_49382);
and UO_1968 (O_1968,N_49975,N_49868);
or UO_1969 (O_1969,N_49364,N_49826);
nor UO_1970 (O_1970,N_49195,N_49499);
or UO_1971 (O_1971,N_49337,N_49789);
nor UO_1972 (O_1972,N_49115,N_49347);
nor UO_1973 (O_1973,N_49693,N_49825);
nor UO_1974 (O_1974,N_49463,N_49348);
or UO_1975 (O_1975,N_49303,N_49516);
and UO_1976 (O_1976,N_49876,N_49112);
nor UO_1977 (O_1977,N_49603,N_49712);
xnor UO_1978 (O_1978,N_49846,N_49954);
and UO_1979 (O_1979,N_49819,N_49993);
and UO_1980 (O_1980,N_49308,N_49969);
nand UO_1981 (O_1981,N_49877,N_49462);
and UO_1982 (O_1982,N_49087,N_49558);
xnor UO_1983 (O_1983,N_49072,N_49137);
or UO_1984 (O_1984,N_49262,N_49154);
nand UO_1985 (O_1985,N_49327,N_49286);
or UO_1986 (O_1986,N_49411,N_49684);
nand UO_1987 (O_1987,N_49257,N_49097);
and UO_1988 (O_1988,N_49467,N_49656);
nand UO_1989 (O_1989,N_49827,N_49900);
nor UO_1990 (O_1990,N_49800,N_49008);
and UO_1991 (O_1991,N_49691,N_49003);
or UO_1992 (O_1992,N_49108,N_49619);
xor UO_1993 (O_1993,N_49117,N_49070);
xor UO_1994 (O_1994,N_49743,N_49418);
nor UO_1995 (O_1995,N_49862,N_49506);
or UO_1996 (O_1996,N_49584,N_49005);
nor UO_1997 (O_1997,N_49515,N_49288);
and UO_1998 (O_1998,N_49317,N_49907);
and UO_1999 (O_1999,N_49283,N_49703);
nor UO_2000 (O_2000,N_49299,N_49738);
or UO_2001 (O_2001,N_49119,N_49793);
or UO_2002 (O_2002,N_49130,N_49234);
nand UO_2003 (O_2003,N_49742,N_49854);
and UO_2004 (O_2004,N_49706,N_49490);
nand UO_2005 (O_2005,N_49733,N_49003);
nand UO_2006 (O_2006,N_49945,N_49632);
or UO_2007 (O_2007,N_49357,N_49251);
and UO_2008 (O_2008,N_49784,N_49542);
nand UO_2009 (O_2009,N_49639,N_49399);
xor UO_2010 (O_2010,N_49204,N_49316);
xor UO_2011 (O_2011,N_49246,N_49993);
nor UO_2012 (O_2012,N_49986,N_49531);
and UO_2013 (O_2013,N_49320,N_49009);
and UO_2014 (O_2014,N_49650,N_49783);
or UO_2015 (O_2015,N_49737,N_49014);
xor UO_2016 (O_2016,N_49589,N_49544);
or UO_2017 (O_2017,N_49278,N_49945);
nand UO_2018 (O_2018,N_49460,N_49976);
and UO_2019 (O_2019,N_49702,N_49791);
and UO_2020 (O_2020,N_49279,N_49545);
and UO_2021 (O_2021,N_49696,N_49830);
nor UO_2022 (O_2022,N_49573,N_49200);
nand UO_2023 (O_2023,N_49604,N_49837);
nor UO_2024 (O_2024,N_49002,N_49871);
nor UO_2025 (O_2025,N_49036,N_49481);
nand UO_2026 (O_2026,N_49521,N_49081);
and UO_2027 (O_2027,N_49348,N_49458);
or UO_2028 (O_2028,N_49178,N_49899);
or UO_2029 (O_2029,N_49908,N_49121);
or UO_2030 (O_2030,N_49661,N_49976);
nand UO_2031 (O_2031,N_49019,N_49461);
or UO_2032 (O_2032,N_49848,N_49361);
xor UO_2033 (O_2033,N_49369,N_49192);
or UO_2034 (O_2034,N_49179,N_49624);
nor UO_2035 (O_2035,N_49044,N_49584);
nand UO_2036 (O_2036,N_49751,N_49342);
nor UO_2037 (O_2037,N_49585,N_49951);
and UO_2038 (O_2038,N_49483,N_49333);
nor UO_2039 (O_2039,N_49806,N_49249);
xnor UO_2040 (O_2040,N_49487,N_49322);
and UO_2041 (O_2041,N_49147,N_49743);
xnor UO_2042 (O_2042,N_49516,N_49573);
nor UO_2043 (O_2043,N_49817,N_49293);
nor UO_2044 (O_2044,N_49347,N_49026);
nand UO_2045 (O_2045,N_49053,N_49898);
or UO_2046 (O_2046,N_49613,N_49004);
xnor UO_2047 (O_2047,N_49203,N_49824);
nand UO_2048 (O_2048,N_49186,N_49638);
or UO_2049 (O_2049,N_49012,N_49456);
nand UO_2050 (O_2050,N_49986,N_49724);
xor UO_2051 (O_2051,N_49667,N_49512);
and UO_2052 (O_2052,N_49307,N_49176);
nor UO_2053 (O_2053,N_49971,N_49096);
nand UO_2054 (O_2054,N_49095,N_49953);
and UO_2055 (O_2055,N_49508,N_49433);
nor UO_2056 (O_2056,N_49170,N_49864);
and UO_2057 (O_2057,N_49006,N_49892);
xnor UO_2058 (O_2058,N_49670,N_49076);
or UO_2059 (O_2059,N_49937,N_49861);
nand UO_2060 (O_2060,N_49242,N_49571);
nand UO_2061 (O_2061,N_49879,N_49808);
nor UO_2062 (O_2062,N_49436,N_49869);
xnor UO_2063 (O_2063,N_49382,N_49600);
nor UO_2064 (O_2064,N_49950,N_49098);
xor UO_2065 (O_2065,N_49970,N_49674);
and UO_2066 (O_2066,N_49016,N_49411);
xnor UO_2067 (O_2067,N_49243,N_49420);
nor UO_2068 (O_2068,N_49343,N_49454);
nor UO_2069 (O_2069,N_49612,N_49168);
and UO_2070 (O_2070,N_49548,N_49615);
xnor UO_2071 (O_2071,N_49201,N_49328);
nor UO_2072 (O_2072,N_49196,N_49400);
nand UO_2073 (O_2073,N_49665,N_49627);
nand UO_2074 (O_2074,N_49340,N_49183);
xor UO_2075 (O_2075,N_49594,N_49736);
nor UO_2076 (O_2076,N_49728,N_49777);
nor UO_2077 (O_2077,N_49100,N_49915);
nor UO_2078 (O_2078,N_49973,N_49797);
nor UO_2079 (O_2079,N_49977,N_49971);
and UO_2080 (O_2080,N_49262,N_49857);
and UO_2081 (O_2081,N_49765,N_49945);
nor UO_2082 (O_2082,N_49029,N_49800);
nand UO_2083 (O_2083,N_49591,N_49856);
xnor UO_2084 (O_2084,N_49135,N_49520);
xor UO_2085 (O_2085,N_49291,N_49413);
or UO_2086 (O_2086,N_49055,N_49286);
nand UO_2087 (O_2087,N_49219,N_49146);
nor UO_2088 (O_2088,N_49206,N_49537);
and UO_2089 (O_2089,N_49107,N_49845);
and UO_2090 (O_2090,N_49431,N_49346);
or UO_2091 (O_2091,N_49157,N_49219);
and UO_2092 (O_2092,N_49697,N_49899);
or UO_2093 (O_2093,N_49999,N_49336);
and UO_2094 (O_2094,N_49794,N_49702);
xor UO_2095 (O_2095,N_49348,N_49270);
nand UO_2096 (O_2096,N_49450,N_49508);
xor UO_2097 (O_2097,N_49621,N_49039);
nand UO_2098 (O_2098,N_49631,N_49422);
nand UO_2099 (O_2099,N_49898,N_49650);
or UO_2100 (O_2100,N_49344,N_49595);
or UO_2101 (O_2101,N_49156,N_49383);
xnor UO_2102 (O_2102,N_49817,N_49469);
nor UO_2103 (O_2103,N_49793,N_49137);
nand UO_2104 (O_2104,N_49003,N_49746);
and UO_2105 (O_2105,N_49269,N_49708);
nand UO_2106 (O_2106,N_49055,N_49677);
or UO_2107 (O_2107,N_49267,N_49112);
nand UO_2108 (O_2108,N_49361,N_49104);
xnor UO_2109 (O_2109,N_49295,N_49046);
nand UO_2110 (O_2110,N_49158,N_49629);
nor UO_2111 (O_2111,N_49669,N_49053);
or UO_2112 (O_2112,N_49668,N_49164);
xor UO_2113 (O_2113,N_49380,N_49075);
nand UO_2114 (O_2114,N_49465,N_49144);
nor UO_2115 (O_2115,N_49087,N_49131);
nor UO_2116 (O_2116,N_49131,N_49611);
nand UO_2117 (O_2117,N_49131,N_49118);
or UO_2118 (O_2118,N_49523,N_49864);
or UO_2119 (O_2119,N_49450,N_49993);
nand UO_2120 (O_2120,N_49546,N_49741);
nor UO_2121 (O_2121,N_49132,N_49786);
xor UO_2122 (O_2122,N_49177,N_49736);
nor UO_2123 (O_2123,N_49056,N_49591);
nor UO_2124 (O_2124,N_49405,N_49917);
xnor UO_2125 (O_2125,N_49762,N_49322);
xor UO_2126 (O_2126,N_49855,N_49566);
and UO_2127 (O_2127,N_49953,N_49311);
nand UO_2128 (O_2128,N_49652,N_49690);
xnor UO_2129 (O_2129,N_49739,N_49765);
nand UO_2130 (O_2130,N_49968,N_49676);
or UO_2131 (O_2131,N_49674,N_49432);
xor UO_2132 (O_2132,N_49354,N_49166);
nor UO_2133 (O_2133,N_49814,N_49418);
or UO_2134 (O_2134,N_49837,N_49281);
nor UO_2135 (O_2135,N_49723,N_49156);
xnor UO_2136 (O_2136,N_49071,N_49789);
and UO_2137 (O_2137,N_49540,N_49736);
or UO_2138 (O_2138,N_49496,N_49529);
or UO_2139 (O_2139,N_49086,N_49431);
or UO_2140 (O_2140,N_49119,N_49712);
nor UO_2141 (O_2141,N_49232,N_49072);
and UO_2142 (O_2142,N_49886,N_49370);
and UO_2143 (O_2143,N_49942,N_49347);
nor UO_2144 (O_2144,N_49991,N_49722);
and UO_2145 (O_2145,N_49570,N_49801);
nor UO_2146 (O_2146,N_49690,N_49421);
nor UO_2147 (O_2147,N_49716,N_49025);
nand UO_2148 (O_2148,N_49069,N_49512);
nor UO_2149 (O_2149,N_49451,N_49931);
nor UO_2150 (O_2150,N_49913,N_49322);
or UO_2151 (O_2151,N_49966,N_49833);
or UO_2152 (O_2152,N_49767,N_49015);
or UO_2153 (O_2153,N_49180,N_49316);
and UO_2154 (O_2154,N_49073,N_49012);
or UO_2155 (O_2155,N_49695,N_49470);
nand UO_2156 (O_2156,N_49744,N_49451);
and UO_2157 (O_2157,N_49507,N_49663);
and UO_2158 (O_2158,N_49852,N_49001);
nand UO_2159 (O_2159,N_49622,N_49202);
xor UO_2160 (O_2160,N_49087,N_49258);
or UO_2161 (O_2161,N_49638,N_49677);
nand UO_2162 (O_2162,N_49857,N_49509);
nand UO_2163 (O_2163,N_49850,N_49832);
or UO_2164 (O_2164,N_49884,N_49255);
nor UO_2165 (O_2165,N_49096,N_49248);
xor UO_2166 (O_2166,N_49815,N_49249);
xor UO_2167 (O_2167,N_49049,N_49622);
or UO_2168 (O_2168,N_49650,N_49455);
xnor UO_2169 (O_2169,N_49467,N_49094);
and UO_2170 (O_2170,N_49732,N_49020);
nand UO_2171 (O_2171,N_49572,N_49018);
and UO_2172 (O_2172,N_49522,N_49247);
nor UO_2173 (O_2173,N_49026,N_49611);
nand UO_2174 (O_2174,N_49502,N_49213);
and UO_2175 (O_2175,N_49625,N_49063);
nand UO_2176 (O_2176,N_49803,N_49026);
or UO_2177 (O_2177,N_49074,N_49425);
xor UO_2178 (O_2178,N_49460,N_49385);
and UO_2179 (O_2179,N_49922,N_49778);
nand UO_2180 (O_2180,N_49615,N_49600);
or UO_2181 (O_2181,N_49829,N_49104);
xnor UO_2182 (O_2182,N_49392,N_49514);
and UO_2183 (O_2183,N_49967,N_49875);
nand UO_2184 (O_2184,N_49602,N_49277);
or UO_2185 (O_2185,N_49527,N_49847);
xnor UO_2186 (O_2186,N_49333,N_49459);
or UO_2187 (O_2187,N_49902,N_49380);
nor UO_2188 (O_2188,N_49346,N_49843);
xnor UO_2189 (O_2189,N_49694,N_49627);
and UO_2190 (O_2190,N_49653,N_49481);
nor UO_2191 (O_2191,N_49016,N_49050);
and UO_2192 (O_2192,N_49791,N_49917);
nor UO_2193 (O_2193,N_49740,N_49515);
and UO_2194 (O_2194,N_49488,N_49175);
nand UO_2195 (O_2195,N_49347,N_49608);
xnor UO_2196 (O_2196,N_49913,N_49894);
nor UO_2197 (O_2197,N_49589,N_49971);
and UO_2198 (O_2198,N_49190,N_49524);
nor UO_2199 (O_2199,N_49557,N_49747);
and UO_2200 (O_2200,N_49078,N_49551);
or UO_2201 (O_2201,N_49270,N_49786);
or UO_2202 (O_2202,N_49439,N_49834);
xor UO_2203 (O_2203,N_49503,N_49518);
nand UO_2204 (O_2204,N_49521,N_49618);
xor UO_2205 (O_2205,N_49997,N_49050);
nand UO_2206 (O_2206,N_49816,N_49468);
xnor UO_2207 (O_2207,N_49002,N_49195);
nor UO_2208 (O_2208,N_49715,N_49359);
nand UO_2209 (O_2209,N_49199,N_49037);
nor UO_2210 (O_2210,N_49254,N_49790);
or UO_2211 (O_2211,N_49978,N_49439);
nand UO_2212 (O_2212,N_49802,N_49348);
and UO_2213 (O_2213,N_49629,N_49370);
or UO_2214 (O_2214,N_49508,N_49961);
nand UO_2215 (O_2215,N_49196,N_49392);
and UO_2216 (O_2216,N_49512,N_49663);
xor UO_2217 (O_2217,N_49727,N_49777);
or UO_2218 (O_2218,N_49807,N_49236);
and UO_2219 (O_2219,N_49156,N_49375);
and UO_2220 (O_2220,N_49771,N_49978);
nor UO_2221 (O_2221,N_49680,N_49399);
nor UO_2222 (O_2222,N_49100,N_49406);
and UO_2223 (O_2223,N_49697,N_49731);
nand UO_2224 (O_2224,N_49858,N_49748);
xnor UO_2225 (O_2225,N_49562,N_49116);
or UO_2226 (O_2226,N_49140,N_49252);
nand UO_2227 (O_2227,N_49439,N_49940);
and UO_2228 (O_2228,N_49185,N_49206);
xnor UO_2229 (O_2229,N_49769,N_49557);
nand UO_2230 (O_2230,N_49399,N_49281);
and UO_2231 (O_2231,N_49379,N_49959);
nor UO_2232 (O_2232,N_49894,N_49821);
nand UO_2233 (O_2233,N_49977,N_49266);
nor UO_2234 (O_2234,N_49013,N_49193);
xor UO_2235 (O_2235,N_49850,N_49933);
or UO_2236 (O_2236,N_49191,N_49627);
xnor UO_2237 (O_2237,N_49520,N_49628);
and UO_2238 (O_2238,N_49926,N_49528);
and UO_2239 (O_2239,N_49949,N_49187);
and UO_2240 (O_2240,N_49668,N_49795);
xor UO_2241 (O_2241,N_49668,N_49041);
nor UO_2242 (O_2242,N_49467,N_49334);
and UO_2243 (O_2243,N_49657,N_49529);
or UO_2244 (O_2244,N_49984,N_49162);
and UO_2245 (O_2245,N_49139,N_49297);
and UO_2246 (O_2246,N_49820,N_49630);
nand UO_2247 (O_2247,N_49245,N_49106);
nand UO_2248 (O_2248,N_49292,N_49838);
nor UO_2249 (O_2249,N_49343,N_49729);
and UO_2250 (O_2250,N_49175,N_49847);
nor UO_2251 (O_2251,N_49850,N_49171);
and UO_2252 (O_2252,N_49381,N_49471);
xnor UO_2253 (O_2253,N_49813,N_49058);
xnor UO_2254 (O_2254,N_49391,N_49483);
and UO_2255 (O_2255,N_49106,N_49055);
nor UO_2256 (O_2256,N_49584,N_49511);
xnor UO_2257 (O_2257,N_49212,N_49098);
or UO_2258 (O_2258,N_49123,N_49063);
or UO_2259 (O_2259,N_49890,N_49739);
and UO_2260 (O_2260,N_49458,N_49695);
or UO_2261 (O_2261,N_49566,N_49606);
nand UO_2262 (O_2262,N_49321,N_49820);
nand UO_2263 (O_2263,N_49563,N_49294);
and UO_2264 (O_2264,N_49680,N_49925);
and UO_2265 (O_2265,N_49337,N_49017);
nand UO_2266 (O_2266,N_49277,N_49359);
or UO_2267 (O_2267,N_49224,N_49495);
and UO_2268 (O_2268,N_49576,N_49008);
xor UO_2269 (O_2269,N_49610,N_49203);
or UO_2270 (O_2270,N_49364,N_49750);
and UO_2271 (O_2271,N_49079,N_49870);
xor UO_2272 (O_2272,N_49163,N_49814);
nor UO_2273 (O_2273,N_49434,N_49407);
and UO_2274 (O_2274,N_49294,N_49242);
and UO_2275 (O_2275,N_49413,N_49934);
nor UO_2276 (O_2276,N_49345,N_49791);
nor UO_2277 (O_2277,N_49355,N_49636);
nand UO_2278 (O_2278,N_49529,N_49582);
and UO_2279 (O_2279,N_49781,N_49033);
and UO_2280 (O_2280,N_49116,N_49208);
xor UO_2281 (O_2281,N_49080,N_49834);
xor UO_2282 (O_2282,N_49968,N_49966);
nand UO_2283 (O_2283,N_49244,N_49503);
nor UO_2284 (O_2284,N_49434,N_49088);
nand UO_2285 (O_2285,N_49686,N_49546);
nand UO_2286 (O_2286,N_49048,N_49017);
or UO_2287 (O_2287,N_49154,N_49937);
nor UO_2288 (O_2288,N_49800,N_49936);
and UO_2289 (O_2289,N_49203,N_49617);
and UO_2290 (O_2290,N_49170,N_49642);
nor UO_2291 (O_2291,N_49248,N_49180);
nor UO_2292 (O_2292,N_49720,N_49501);
or UO_2293 (O_2293,N_49570,N_49201);
and UO_2294 (O_2294,N_49014,N_49562);
or UO_2295 (O_2295,N_49881,N_49025);
nand UO_2296 (O_2296,N_49953,N_49218);
xor UO_2297 (O_2297,N_49265,N_49164);
or UO_2298 (O_2298,N_49743,N_49914);
and UO_2299 (O_2299,N_49088,N_49537);
nand UO_2300 (O_2300,N_49829,N_49559);
nor UO_2301 (O_2301,N_49310,N_49314);
or UO_2302 (O_2302,N_49738,N_49072);
and UO_2303 (O_2303,N_49209,N_49739);
xnor UO_2304 (O_2304,N_49308,N_49745);
or UO_2305 (O_2305,N_49008,N_49810);
or UO_2306 (O_2306,N_49333,N_49236);
nor UO_2307 (O_2307,N_49424,N_49389);
nor UO_2308 (O_2308,N_49680,N_49081);
nand UO_2309 (O_2309,N_49408,N_49808);
or UO_2310 (O_2310,N_49134,N_49829);
or UO_2311 (O_2311,N_49471,N_49649);
or UO_2312 (O_2312,N_49898,N_49092);
nand UO_2313 (O_2313,N_49542,N_49229);
nor UO_2314 (O_2314,N_49988,N_49409);
and UO_2315 (O_2315,N_49512,N_49890);
nor UO_2316 (O_2316,N_49668,N_49191);
nor UO_2317 (O_2317,N_49366,N_49455);
nor UO_2318 (O_2318,N_49033,N_49999);
xor UO_2319 (O_2319,N_49173,N_49336);
and UO_2320 (O_2320,N_49341,N_49193);
and UO_2321 (O_2321,N_49051,N_49899);
and UO_2322 (O_2322,N_49531,N_49875);
xnor UO_2323 (O_2323,N_49152,N_49472);
and UO_2324 (O_2324,N_49265,N_49505);
or UO_2325 (O_2325,N_49276,N_49674);
and UO_2326 (O_2326,N_49049,N_49772);
xor UO_2327 (O_2327,N_49166,N_49448);
nand UO_2328 (O_2328,N_49725,N_49135);
xnor UO_2329 (O_2329,N_49013,N_49820);
and UO_2330 (O_2330,N_49128,N_49095);
nand UO_2331 (O_2331,N_49624,N_49156);
or UO_2332 (O_2332,N_49837,N_49260);
or UO_2333 (O_2333,N_49606,N_49421);
nor UO_2334 (O_2334,N_49078,N_49216);
nor UO_2335 (O_2335,N_49718,N_49995);
nor UO_2336 (O_2336,N_49217,N_49675);
nor UO_2337 (O_2337,N_49239,N_49697);
xnor UO_2338 (O_2338,N_49565,N_49554);
nor UO_2339 (O_2339,N_49174,N_49099);
nor UO_2340 (O_2340,N_49353,N_49991);
nand UO_2341 (O_2341,N_49756,N_49112);
nor UO_2342 (O_2342,N_49787,N_49098);
nor UO_2343 (O_2343,N_49960,N_49756);
or UO_2344 (O_2344,N_49383,N_49044);
or UO_2345 (O_2345,N_49874,N_49772);
nor UO_2346 (O_2346,N_49493,N_49289);
nor UO_2347 (O_2347,N_49983,N_49735);
and UO_2348 (O_2348,N_49262,N_49644);
xnor UO_2349 (O_2349,N_49808,N_49897);
and UO_2350 (O_2350,N_49126,N_49732);
or UO_2351 (O_2351,N_49205,N_49123);
nand UO_2352 (O_2352,N_49536,N_49609);
nor UO_2353 (O_2353,N_49642,N_49318);
and UO_2354 (O_2354,N_49976,N_49720);
xor UO_2355 (O_2355,N_49715,N_49964);
xor UO_2356 (O_2356,N_49139,N_49322);
nand UO_2357 (O_2357,N_49205,N_49564);
nor UO_2358 (O_2358,N_49431,N_49114);
and UO_2359 (O_2359,N_49525,N_49055);
or UO_2360 (O_2360,N_49250,N_49495);
and UO_2361 (O_2361,N_49626,N_49296);
nor UO_2362 (O_2362,N_49043,N_49915);
and UO_2363 (O_2363,N_49775,N_49132);
xnor UO_2364 (O_2364,N_49760,N_49978);
nor UO_2365 (O_2365,N_49512,N_49099);
and UO_2366 (O_2366,N_49836,N_49813);
xnor UO_2367 (O_2367,N_49677,N_49963);
and UO_2368 (O_2368,N_49560,N_49952);
nor UO_2369 (O_2369,N_49974,N_49858);
nor UO_2370 (O_2370,N_49973,N_49972);
xor UO_2371 (O_2371,N_49193,N_49558);
or UO_2372 (O_2372,N_49515,N_49672);
and UO_2373 (O_2373,N_49435,N_49061);
and UO_2374 (O_2374,N_49658,N_49876);
nand UO_2375 (O_2375,N_49420,N_49995);
xor UO_2376 (O_2376,N_49621,N_49445);
nand UO_2377 (O_2377,N_49775,N_49365);
xor UO_2378 (O_2378,N_49601,N_49915);
and UO_2379 (O_2379,N_49609,N_49436);
nand UO_2380 (O_2380,N_49764,N_49127);
or UO_2381 (O_2381,N_49631,N_49997);
and UO_2382 (O_2382,N_49749,N_49718);
and UO_2383 (O_2383,N_49987,N_49520);
and UO_2384 (O_2384,N_49943,N_49673);
and UO_2385 (O_2385,N_49674,N_49831);
nor UO_2386 (O_2386,N_49991,N_49316);
nand UO_2387 (O_2387,N_49361,N_49083);
and UO_2388 (O_2388,N_49824,N_49815);
nand UO_2389 (O_2389,N_49342,N_49633);
nand UO_2390 (O_2390,N_49026,N_49454);
nor UO_2391 (O_2391,N_49263,N_49813);
nand UO_2392 (O_2392,N_49764,N_49627);
nor UO_2393 (O_2393,N_49646,N_49247);
nor UO_2394 (O_2394,N_49169,N_49166);
xnor UO_2395 (O_2395,N_49569,N_49618);
nand UO_2396 (O_2396,N_49210,N_49851);
or UO_2397 (O_2397,N_49423,N_49969);
nand UO_2398 (O_2398,N_49664,N_49952);
nand UO_2399 (O_2399,N_49594,N_49791);
xnor UO_2400 (O_2400,N_49803,N_49895);
xnor UO_2401 (O_2401,N_49439,N_49812);
nand UO_2402 (O_2402,N_49102,N_49272);
and UO_2403 (O_2403,N_49249,N_49509);
xor UO_2404 (O_2404,N_49333,N_49962);
and UO_2405 (O_2405,N_49774,N_49726);
xnor UO_2406 (O_2406,N_49017,N_49664);
nor UO_2407 (O_2407,N_49597,N_49311);
nor UO_2408 (O_2408,N_49568,N_49898);
xnor UO_2409 (O_2409,N_49188,N_49454);
xnor UO_2410 (O_2410,N_49402,N_49953);
nor UO_2411 (O_2411,N_49910,N_49785);
nand UO_2412 (O_2412,N_49733,N_49752);
nor UO_2413 (O_2413,N_49926,N_49348);
nor UO_2414 (O_2414,N_49881,N_49923);
or UO_2415 (O_2415,N_49904,N_49163);
nand UO_2416 (O_2416,N_49472,N_49900);
nor UO_2417 (O_2417,N_49153,N_49528);
and UO_2418 (O_2418,N_49268,N_49246);
xor UO_2419 (O_2419,N_49866,N_49291);
and UO_2420 (O_2420,N_49034,N_49498);
nand UO_2421 (O_2421,N_49821,N_49107);
or UO_2422 (O_2422,N_49352,N_49672);
nor UO_2423 (O_2423,N_49386,N_49697);
xnor UO_2424 (O_2424,N_49294,N_49353);
and UO_2425 (O_2425,N_49344,N_49260);
or UO_2426 (O_2426,N_49323,N_49856);
xor UO_2427 (O_2427,N_49089,N_49256);
and UO_2428 (O_2428,N_49925,N_49452);
or UO_2429 (O_2429,N_49421,N_49314);
and UO_2430 (O_2430,N_49069,N_49039);
xnor UO_2431 (O_2431,N_49128,N_49560);
xor UO_2432 (O_2432,N_49958,N_49179);
nor UO_2433 (O_2433,N_49753,N_49567);
nand UO_2434 (O_2434,N_49485,N_49259);
xnor UO_2435 (O_2435,N_49057,N_49505);
nor UO_2436 (O_2436,N_49328,N_49702);
and UO_2437 (O_2437,N_49747,N_49953);
xor UO_2438 (O_2438,N_49463,N_49741);
nand UO_2439 (O_2439,N_49838,N_49303);
nand UO_2440 (O_2440,N_49961,N_49888);
and UO_2441 (O_2441,N_49112,N_49982);
nor UO_2442 (O_2442,N_49116,N_49034);
nand UO_2443 (O_2443,N_49851,N_49099);
nor UO_2444 (O_2444,N_49893,N_49482);
xnor UO_2445 (O_2445,N_49065,N_49270);
and UO_2446 (O_2446,N_49373,N_49103);
nor UO_2447 (O_2447,N_49112,N_49521);
xnor UO_2448 (O_2448,N_49560,N_49806);
and UO_2449 (O_2449,N_49092,N_49164);
xnor UO_2450 (O_2450,N_49083,N_49347);
nand UO_2451 (O_2451,N_49284,N_49973);
or UO_2452 (O_2452,N_49501,N_49041);
xnor UO_2453 (O_2453,N_49990,N_49229);
or UO_2454 (O_2454,N_49103,N_49855);
nand UO_2455 (O_2455,N_49237,N_49557);
and UO_2456 (O_2456,N_49967,N_49176);
and UO_2457 (O_2457,N_49021,N_49377);
and UO_2458 (O_2458,N_49540,N_49510);
or UO_2459 (O_2459,N_49690,N_49352);
and UO_2460 (O_2460,N_49641,N_49646);
and UO_2461 (O_2461,N_49935,N_49425);
and UO_2462 (O_2462,N_49508,N_49266);
nor UO_2463 (O_2463,N_49828,N_49646);
or UO_2464 (O_2464,N_49887,N_49514);
and UO_2465 (O_2465,N_49572,N_49130);
nand UO_2466 (O_2466,N_49256,N_49940);
xor UO_2467 (O_2467,N_49171,N_49782);
nor UO_2468 (O_2468,N_49937,N_49882);
or UO_2469 (O_2469,N_49371,N_49493);
nor UO_2470 (O_2470,N_49257,N_49156);
or UO_2471 (O_2471,N_49642,N_49091);
and UO_2472 (O_2472,N_49111,N_49131);
and UO_2473 (O_2473,N_49550,N_49949);
and UO_2474 (O_2474,N_49528,N_49603);
nand UO_2475 (O_2475,N_49681,N_49293);
nor UO_2476 (O_2476,N_49625,N_49213);
nor UO_2477 (O_2477,N_49468,N_49884);
xor UO_2478 (O_2478,N_49753,N_49130);
xor UO_2479 (O_2479,N_49290,N_49475);
nand UO_2480 (O_2480,N_49425,N_49739);
nand UO_2481 (O_2481,N_49430,N_49842);
nor UO_2482 (O_2482,N_49193,N_49391);
and UO_2483 (O_2483,N_49421,N_49554);
xor UO_2484 (O_2484,N_49630,N_49645);
or UO_2485 (O_2485,N_49591,N_49920);
xnor UO_2486 (O_2486,N_49957,N_49318);
nor UO_2487 (O_2487,N_49694,N_49193);
and UO_2488 (O_2488,N_49368,N_49062);
nand UO_2489 (O_2489,N_49714,N_49202);
and UO_2490 (O_2490,N_49770,N_49194);
xnor UO_2491 (O_2491,N_49093,N_49122);
xnor UO_2492 (O_2492,N_49717,N_49784);
or UO_2493 (O_2493,N_49468,N_49829);
nor UO_2494 (O_2494,N_49334,N_49258);
or UO_2495 (O_2495,N_49715,N_49193);
xnor UO_2496 (O_2496,N_49979,N_49642);
nand UO_2497 (O_2497,N_49907,N_49588);
xnor UO_2498 (O_2498,N_49517,N_49928);
nor UO_2499 (O_2499,N_49853,N_49359);
nor UO_2500 (O_2500,N_49096,N_49856);
or UO_2501 (O_2501,N_49698,N_49610);
xnor UO_2502 (O_2502,N_49881,N_49653);
nand UO_2503 (O_2503,N_49332,N_49426);
nor UO_2504 (O_2504,N_49587,N_49955);
nor UO_2505 (O_2505,N_49506,N_49375);
or UO_2506 (O_2506,N_49401,N_49676);
and UO_2507 (O_2507,N_49457,N_49946);
or UO_2508 (O_2508,N_49141,N_49444);
xor UO_2509 (O_2509,N_49498,N_49527);
and UO_2510 (O_2510,N_49185,N_49715);
and UO_2511 (O_2511,N_49179,N_49746);
nor UO_2512 (O_2512,N_49851,N_49746);
nor UO_2513 (O_2513,N_49426,N_49148);
and UO_2514 (O_2514,N_49253,N_49666);
xnor UO_2515 (O_2515,N_49436,N_49174);
and UO_2516 (O_2516,N_49839,N_49976);
nor UO_2517 (O_2517,N_49355,N_49130);
and UO_2518 (O_2518,N_49082,N_49811);
nand UO_2519 (O_2519,N_49820,N_49514);
nor UO_2520 (O_2520,N_49758,N_49819);
or UO_2521 (O_2521,N_49204,N_49755);
nand UO_2522 (O_2522,N_49068,N_49872);
or UO_2523 (O_2523,N_49903,N_49782);
and UO_2524 (O_2524,N_49481,N_49817);
nor UO_2525 (O_2525,N_49638,N_49927);
nand UO_2526 (O_2526,N_49191,N_49296);
nor UO_2527 (O_2527,N_49099,N_49331);
nor UO_2528 (O_2528,N_49805,N_49203);
or UO_2529 (O_2529,N_49911,N_49320);
xor UO_2530 (O_2530,N_49684,N_49276);
or UO_2531 (O_2531,N_49821,N_49248);
nor UO_2532 (O_2532,N_49388,N_49533);
or UO_2533 (O_2533,N_49000,N_49657);
nor UO_2534 (O_2534,N_49725,N_49398);
nor UO_2535 (O_2535,N_49629,N_49095);
nand UO_2536 (O_2536,N_49606,N_49239);
nand UO_2537 (O_2537,N_49315,N_49301);
or UO_2538 (O_2538,N_49671,N_49044);
or UO_2539 (O_2539,N_49511,N_49969);
and UO_2540 (O_2540,N_49794,N_49799);
and UO_2541 (O_2541,N_49069,N_49586);
nand UO_2542 (O_2542,N_49144,N_49881);
nand UO_2543 (O_2543,N_49150,N_49235);
or UO_2544 (O_2544,N_49393,N_49691);
nor UO_2545 (O_2545,N_49431,N_49902);
xnor UO_2546 (O_2546,N_49316,N_49386);
nor UO_2547 (O_2547,N_49610,N_49832);
and UO_2548 (O_2548,N_49456,N_49629);
xnor UO_2549 (O_2549,N_49037,N_49466);
or UO_2550 (O_2550,N_49154,N_49716);
and UO_2551 (O_2551,N_49292,N_49608);
nand UO_2552 (O_2552,N_49161,N_49287);
nor UO_2553 (O_2553,N_49525,N_49081);
or UO_2554 (O_2554,N_49715,N_49691);
xor UO_2555 (O_2555,N_49662,N_49157);
xnor UO_2556 (O_2556,N_49782,N_49813);
xor UO_2557 (O_2557,N_49879,N_49265);
nand UO_2558 (O_2558,N_49915,N_49871);
xnor UO_2559 (O_2559,N_49362,N_49126);
nand UO_2560 (O_2560,N_49827,N_49392);
or UO_2561 (O_2561,N_49226,N_49360);
nand UO_2562 (O_2562,N_49066,N_49875);
and UO_2563 (O_2563,N_49695,N_49123);
and UO_2564 (O_2564,N_49919,N_49192);
nand UO_2565 (O_2565,N_49759,N_49760);
nand UO_2566 (O_2566,N_49540,N_49264);
and UO_2567 (O_2567,N_49789,N_49830);
nand UO_2568 (O_2568,N_49603,N_49500);
nand UO_2569 (O_2569,N_49125,N_49754);
nor UO_2570 (O_2570,N_49846,N_49349);
xnor UO_2571 (O_2571,N_49008,N_49268);
xor UO_2572 (O_2572,N_49772,N_49427);
nor UO_2573 (O_2573,N_49385,N_49979);
nand UO_2574 (O_2574,N_49338,N_49909);
or UO_2575 (O_2575,N_49020,N_49736);
and UO_2576 (O_2576,N_49705,N_49308);
or UO_2577 (O_2577,N_49851,N_49492);
nor UO_2578 (O_2578,N_49220,N_49600);
and UO_2579 (O_2579,N_49963,N_49341);
xor UO_2580 (O_2580,N_49906,N_49000);
and UO_2581 (O_2581,N_49293,N_49921);
or UO_2582 (O_2582,N_49609,N_49807);
nand UO_2583 (O_2583,N_49904,N_49193);
and UO_2584 (O_2584,N_49816,N_49972);
and UO_2585 (O_2585,N_49082,N_49080);
nor UO_2586 (O_2586,N_49829,N_49798);
nor UO_2587 (O_2587,N_49074,N_49077);
or UO_2588 (O_2588,N_49096,N_49572);
xnor UO_2589 (O_2589,N_49027,N_49623);
nand UO_2590 (O_2590,N_49773,N_49144);
and UO_2591 (O_2591,N_49490,N_49470);
or UO_2592 (O_2592,N_49022,N_49369);
nor UO_2593 (O_2593,N_49044,N_49862);
nand UO_2594 (O_2594,N_49822,N_49199);
nand UO_2595 (O_2595,N_49371,N_49781);
nor UO_2596 (O_2596,N_49344,N_49990);
or UO_2597 (O_2597,N_49734,N_49925);
xor UO_2598 (O_2598,N_49310,N_49916);
xnor UO_2599 (O_2599,N_49286,N_49402);
nor UO_2600 (O_2600,N_49453,N_49726);
and UO_2601 (O_2601,N_49556,N_49364);
xnor UO_2602 (O_2602,N_49090,N_49463);
and UO_2603 (O_2603,N_49743,N_49066);
nand UO_2604 (O_2604,N_49996,N_49732);
nand UO_2605 (O_2605,N_49191,N_49076);
or UO_2606 (O_2606,N_49802,N_49723);
nand UO_2607 (O_2607,N_49094,N_49281);
nand UO_2608 (O_2608,N_49290,N_49253);
nand UO_2609 (O_2609,N_49718,N_49873);
nand UO_2610 (O_2610,N_49224,N_49135);
xor UO_2611 (O_2611,N_49315,N_49037);
xor UO_2612 (O_2612,N_49702,N_49067);
or UO_2613 (O_2613,N_49918,N_49409);
nand UO_2614 (O_2614,N_49258,N_49819);
and UO_2615 (O_2615,N_49822,N_49884);
and UO_2616 (O_2616,N_49622,N_49067);
or UO_2617 (O_2617,N_49801,N_49968);
xor UO_2618 (O_2618,N_49284,N_49165);
xor UO_2619 (O_2619,N_49384,N_49346);
and UO_2620 (O_2620,N_49757,N_49101);
xnor UO_2621 (O_2621,N_49679,N_49922);
or UO_2622 (O_2622,N_49734,N_49998);
nand UO_2623 (O_2623,N_49017,N_49467);
nand UO_2624 (O_2624,N_49978,N_49969);
or UO_2625 (O_2625,N_49024,N_49713);
and UO_2626 (O_2626,N_49083,N_49986);
or UO_2627 (O_2627,N_49342,N_49976);
and UO_2628 (O_2628,N_49483,N_49430);
or UO_2629 (O_2629,N_49381,N_49399);
and UO_2630 (O_2630,N_49050,N_49988);
xor UO_2631 (O_2631,N_49466,N_49652);
nor UO_2632 (O_2632,N_49107,N_49554);
or UO_2633 (O_2633,N_49315,N_49835);
xnor UO_2634 (O_2634,N_49858,N_49742);
and UO_2635 (O_2635,N_49477,N_49068);
and UO_2636 (O_2636,N_49706,N_49055);
nand UO_2637 (O_2637,N_49804,N_49871);
nand UO_2638 (O_2638,N_49994,N_49732);
nand UO_2639 (O_2639,N_49309,N_49929);
or UO_2640 (O_2640,N_49407,N_49525);
nand UO_2641 (O_2641,N_49387,N_49245);
xnor UO_2642 (O_2642,N_49256,N_49622);
xnor UO_2643 (O_2643,N_49803,N_49133);
xnor UO_2644 (O_2644,N_49100,N_49862);
xnor UO_2645 (O_2645,N_49480,N_49627);
nor UO_2646 (O_2646,N_49255,N_49407);
and UO_2647 (O_2647,N_49354,N_49936);
nor UO_2648 (O_2648,N_49820,N_49270);
and UO_2649 (O_2649,N_49130,N_49131);
xnor UO_2650 (O_2650,N_49680,N_49090);
nor UO_2651 (O_2651,N_49077,N_49949);
nand UO_2652 (O_2652,N_49617,N_49500);
nor UO_2653 (O_2653,N_49459,N_49782);
nor UO_2654 (O_2654,N_49564,N_49397);
nor UO_2655 (O_2655,N_49480,N_49589);
nand UO_2656 (O_2656,N_49172,N_49328);
or UO_2657 (O_2657,N_49800,N_49782);
and UO_2658 (O_2658,N_49318,N_49344);
nand UO_2659 (O_2659,N_49856,N_49781);
nor UO_2660 (O_2660,N_49479,N_49171);
and UO_2661 (O_2661,N_49617,N_49961);
nor UO_2662 (O_2662,N_49448,N_49117);
and UO_2663 (O_2663,N_49091,N_49362);
nand UO_2664 (O_2664,N_49913,N_49671);
nor UO_2665 (O_2665,N_49013,N_49030);
nor UO_2666 (O_2666,N_49933,N_49413);
nor UO_2667 (O_2667,N_49879,N_49001);
nand UO_2668 (O_2668,N_49910,N_49685);
nor UO_2669 (O_2669,N_49518,N_49132);
nor UO_2670 (O_2670,N_49627,N_49580);
and UO_2671 (O_2671,N_49624,N_49814);
and UO_2672 (O_2672,N_49678,N_49151);
and UO_2673 (O_2673,N_49370,N_49104);
nor UO_2674 (O_2674,N_49786,N_49478);
xor UO_2675 (O_2675,N_49311,N_49862);
and UO_2676 (O_2676,N_49111,N_49941);
or UO_2677 (O_2677,N_49726,N_49793);
and UO_2678 (O_2678,N_49468,N_49451);
or UO_2679 (O_2679,N_49535,N_49703);
nor UO_2680 (O_2680,N_49637,N_49380);
nor UO_2681 (O_2681,N_49067,N_49798);
nand UO_2682 (O_2682,N_49435,N_49310);
or UO_2683 (O_2683,N_49387,N_49338);
xnor UO_2684 (O_2684,N_49632,N_49420);
and UO_2685 (O_2685,N_49952,N_49574);
or UO_2686 (O_2686,N_49242,N_49543);
and UO_2687 (O_2687,N_49855,N_49032);
nand UO_2688 (O_2688,N_49466,N_49601);
or UO_2689 (O_2689,N_49175,N_49996);
or UO_2690 (O_2690,N_49481,N_49418);
nor UO_2691 (O_2691,N_49558,N_49849);
or UO_2692 (O_2692,N_49850,N_49362);
and UO_2693 (O_2693,N_49335,N_49972);
and UO_2694 (O_2694,N_49049,N_49456);
nor UO_2695 (O_2695,N_49023,N_49521);
xor UO_2696 (O_2696,N_49734,N_49579);
xor UO_2697 (O_2697,N_49697,N_49159);
and UO_2698 (O_2698,N_49609,N_49970);
xor UO_2699 (O_2699,N_49258,N_49321);
xor UO_2700 (O_2700,N_49935,N_49538);
nand UO_2701 (O_2701,N_49493,N_49117);
nor UO_2702 (O_2702,N_49717,N_49268);
or UO_2703 (O_2703,N_49408,N_49438);
xor UO_2704 (O_2704,N_49680,N_49200);
xor UO_2705 (O_2705,N_49204,N_49367);
nand UO_2706 (O_2706,N_49127,N_49331);
nand UO_2707 (O_2707,N_49887,N_49237);
or UO_2708 (O_2708,N_49275,N_49069);
nand UO_2709 (O_2709,N_49764,N_49071);
nand UO_2710 (O_2710,N_49013,N_49166);
nor UO_2711 (O_2711,N_49868,N_49254);
xnor UO_2712 (O_2712,N_49604,N_49041);
or UO_2713 (O_2713,N_49154,N_49495);
xnor UO_2714 (O_2714,N_49432,N_49106);
nor UO_2715 (O_2715,N_49838,N_49242);
and UO_2716 (O_2716,N_49613,N_49075);
or UO_2717 (O_2717,N_49686,N_49999);
xor UO_2718 (O_2718,N_49729,N_49249);
xor UO_2719 (O_2719,N_49522,N_49769);
nand UO_2720 (O_2720,N_49591,N_49686);
or UO_2721 (O_2721,N_49932,N_49168);
and UO_2722 (O_2722,N_49925,N_49347);
xnor UO_2723 (O_2723,N_49517,N_49359);
or UO_2724 (O_2724,N_49044,N_49692);
nor UO_2725 (O_2725,N_49530,N_49325);
or UO_2726 (O_2726,N_49963,N_49758);
and UO_2727 (O_2727,N_49613,N_49916);
nand UO_2728 (O_2728,N_49478,N_49429);
nand UO_2729 (O_2729,N_49865,N_49744);
xnor UO_2730 (O_2730,N_49467,N_49940);
or UO_2731 (O_2731,N_49206,N_49572);
nand UO_2732 (O_2732,N_49409,N_49971);
or UO_2733 (O_2733,N_49091,N_49116);
and UO_2734 (O_2734,N_49957,N_49101);
xor UO_2735 (O_2735,N_49072,N_49956);
xor UO_2736 (O_2736,N_49483,N_49216);
nand UO_2737 (O_2737,N_49867,N_49948);
nor UO_2738 (O_2738,N_49006,N_49831);
xnor UO_2739 (O_2739,N_49899,N_49250);
xnor UO_2740 (O_2740,N_49781,N_49211);
nand UO_2741 (O_2741,N_49879,N_49960);
nor UO_2742 (O_2742,N_49526,N_49593);
nor UO_2743 (O_2743,N_49421,N_49810);
and UO_2744 (O_2744,N_49255,N_49573);
nor UO_2745 (O_2745,N_49821,N_49452);
and UO_2746 (O_2746,N_49668,N_49740);
nand UO_2747 (O_2747,N_49491,N_49111);
and UO_2748 (O_2748,N_49165,N_49821);
and UO_2749 (O_2749,N_49985,N_49035);
xor UO_2750 (O_2750,N_49979,N_49630);
nand UO_2751 (O_2751,N_49188,N_49087);
nor UO_2752 (O_2752,N_49400,N_49991);
or UO_2753 (O_2753,N_49097,N_49427);
and UO_2754 (O_2754,N_49242,N_49019);
nand UO_2755 (O_2755,N_49000,N_49636);
or UO_2756 (O_2756,N_49949,N_49952);
and UO_2757 (O_2757,N_49862,N_49033);
and UO_2758 (O_2758,N_49114,N_49979);
or UO_2759 (O_2759,N_49854,N_49905);
and UO_2760 (O_2760,N_49425,N_49084);
xor UO_2761 (O_2761,N_49462,N_49091);
xor UO_2762 (O_2762,N_49385,N_49644);
nor UO_2763 (O_2763,N_49230,N_49783);
nor UO_2764 (O_2764,N_49395,N_49709);
xor UO_2765 (O_2765,N_49956,N_49947);
xor UO_2766 (O_2766,N_49725,N_49280);
xnor UO_2767 (O_2767,N_49466,N_49648);
and UO_2768 (O_2768,N_49716,N_49325);
nand UO_2769 (O_2769,N_49416,N_49364);
nor UO_2770 (O_2770,N_49364,N_49408);
or UO_2771 (O_2771,N_49197,N_49117);
or UO_2772 (O_2772,N_49646,N_49669);
xnor UO_2773 (O_2773,N_49939,N_49319);
xnor UO_2774 (O_2774,N_49855,N_49401);
or UO_2775 (O_2775,N_49473,N_49286);
xnor UO_2776 (O_2776,N_49684,N_49250);
or UO_2777 (O_2777,N_49126,N_49856);
xnor UO_2778 (O_2778,N_49828,N_49472);
or UO_2779 (O_2779,N_49688,N_49771);
xor UO_2780 (O_2780,N_49104,N_49794);
or UO_2781 (O_2781,N_49900,N_49209);
or UO_2782 (O_2782,N_49027,N_49083);
or UO_2783 (O_2783,N_49364,N_49027);
or UO_2784 (O_2784,N_49986,N_49428);
or UO_2785 (O_2785,N_49970,N_49349);
nand UO_2786 (O_2786,N_49978,N_49276);
or UO_2787 (O_2787,N_49723,N_49907);
nor UO_2788 (O_2788,N_49807,N_49394);
and UO_2789 (O_2789,N_49003,N_49432);
nand UO_2790 (O_2790,N_49688,N_49973);
nor UO_2791 (O_2791,N_49927,N_49748);
nor UO_2792 (O_2792,N_49372,N_49776);
or UO_2793 (O_2793,N_49450,N_49506);
nand UO_2794 (O_2794,N_49248,N_49030);
or UO_2795 (O_2795,N_49929,N_49343);
xnor UO_2796 (O_2796,N_49593,N_49786);
nor UO_2797 (O_2797,N_49968,N_49285);
or UO_2798 (O_2798,N_49396,N_49471);
xor UO_2799 (O_2799,N_49223,N_49215);
nand UO_2800 (O_2800,N_49455,N_49393);
or UO_2801 (O_2801,N_49581,N_49088);
and UO_2802 (O_2802,N_49956,N_49289);
or UO_2803 (O_2803,N_49859,N_49244);
nand UO_2804 (O_2804,N_49460,N_49915);
and UO_2805 (O_2805,N_49878,N_49603);
and UO_2806 (O_2806,N_49677,N_49825);
or UO_2807 (O_2807,N_49027,N_49694);
nand UO_2808 (O_2808,N_49930,N_49805);
nand UO_2809 (O_2809,N_49570,N_49016);
nand UO_2810 (O_2810,N_49751,N_49561);
or UO_2811 (O_2811,N_49703,N_49450);
xnor UO_2812 (O_2812,N_49106,N_49717);
nand UO_2813 (O_2813,N_49185,N_49124);
nand UO_2814 (O_2814,N_49213,N_49595);
or UO_2815 (O_2815,N_49957,N_49689);
and UO_2816 (O_2816,N_49799,N_49181);
nand UO_2817 (O_2817,N_49734,N_49828);
and UO_2818 (O_2818,N_49049,N_49691);
and UO_2819 (O_2819,N_49784,N_49945);
or UO_2820 (O_2820,N_49693,N_49308);
nor UO_2821 (O_2821,N_49435,N_49085);
xor UO_2822 (O_2822,N_49399,N_49428);
and UO_2823 (O_2823,N_49279,N_49710);
and UO_2824 (O_2824,N_49866,N_49966);
nand UO_2825 (O_2825,N_49021,N_49536);
and UO_2826 (O_2826,N_49598,N_49796);
nor UO_2827 (O_2827,N_49975,N_49663);
or UO_2828 (O_2828,N_49970,N_49804);
or UO_2829 (O_2829,N_49922,N_49570);
nor UO_2830 (O_2830,N_49645,N_49381);
or UO_2831 (O_2831,N_49865,N_49832);
and UO_2832 (O_2832,N_49701,N_49672);
or UO_2833 (O_2833,N_49035,N_49175);
or UO_2834 (O_2834,N_49018,N_49062);
or UO_2835 (O_2835,N_49654,N_49698);
nand UO_2836 (O_2836,N_49138,N_49653);
nor UO_2837 (O_2837,N_49484,N_49719);
or UO_2838 (O_2838,N_49342,N_49424);
xnor UO_2839 (O_2839,N_49388,N_49059);
or UO_2840 (O_2840,N_49622,N_49212);
or UO_2841 (O_2841,N_49216,N_49634);
xor UO_2842 (O_2842,N_49379,N_49519);
nand UO_2843 (O_2843,N_49307,N_49178);
or UO_2844 (O_2844,N_49793,N_49266);
xnor UO_2845 (O_2845,N_49177,N_49516);
xnor UO_2846 (O_2846,N_49683,N_49429);
or UO_2847 (O_2847,N_49773,N_49379);
or UO_2848 (O_2848,N_49261,N_49255);
or UO_2849 (O_2849,N_49988,N_49806);
xnor UO_2850 (O_2850,N_49424,N_49660);
nand UO_2851 (O_2851,N_49885,N_49003);
nor UO_2852 (O_2852,N_49411,N_49802);
nand UO_2853 (O_2853,N_49303,N_49452);
nor UO_2854 (O_2854,N_49235,N_49073);
and UO_2855 (O_2855,N_49560,N_49642);
nand UO_2856 (O_2856,N_49430,N_49220);
nor UO_2857 (O_2857,N_49163,N_49903);
nor UO_2858 (O_2858,N_49644,N_49257);
nand UO_2859 (O_2859,N_49724,N_49896);
nand UO_2860 (O_2860,N_49193,N_49154);
and UO_2861 (O_2861,N_49860,N_49706);
and UO_2862 (O_2862,N_49343,N_49404);
xnor UO_2863 (O_2863,N_49788,N_49987);
nand UO_2864 (O_2864,N_49730,N_49444);
and UO_2865 (O_2865,N_49246,N_49437);
and UO_2866 (O_2866,N_49495,N_49881);
or UO_2867 (O_2867,N_49521,N_49970);
or UO_2868 (O_2868,N_49264,N_49879);
xnor UO_2869 (O_2869,N_49171,N_49887);
nand UO_2870 (O_2870,N_49614,N_49200);
xnor UO_2871 (O_2871,N_49907,N_49295);
xnor UO_2872 (O_2872,N_49156,N_49812);
nand UO_2873 (O_2873,N_49773,N_49302);
nand UO_2874 (O_2874,N_49223,N_49420);
nor UO_2875 (O_2875,N_49335,N_49399);
xor UO_2876 (O_2876,N_49415,N_49889);
xor UO_2877 (O_2877,N_49022,N_49126);
nand UO_2878 (O_2878,N_49120,N_49861);
nor UO_2879 (O_2879,N_49663,N_49818);
nand UO_2880 (O_2880,N_49722,N_49134);
nor UO_2881 (O_2881,N_49674,N_49448);
nor UO_2882 (O_2882,N_49650,N_49043);
and UO_2883 (O_2883,N_49846,N_49348);
nor UO_2884 (O_2884,N_49108,N_49251);
xnor UO_2885 (O_2885,N_49612,N_49007);
nand UO_2886 (O_2886,N_49956,N_49086);
xor UO_2887 (O_2887,N_49212,N_49089);
or UO_2888 (O_2888,N_49163,N_49967);
and UO_2889 (O_2889,N_49680,N_49297);
nor UO_2890 (O_2890,N_49793,N_49013);
nand UO_2891 (O_2891,N_49481,N_49230);
nand UO_2892 (O_2892,N_49855,N_49537);
xor UO_2893 (O_2893,N_49638,N_49944);
and UO_2894 (O_2894,N_49200,N_49440);
nand UO_2895 (O_2895,N_49951,N_49165);
nand UO_2896 (O_2896,N_49483,N_49634);
and UO_2897 (O_2897,N_49416,N_49986);
nand UO_2898 (O_2898,N_49910,N_49065);
and UO_2899 (O_2899,N_49906,N_49417);
or UO_2900 (O_2900,N_49742,N_49058);
xnor UO_2901 (O_2901,N_49551,N_49267);
xor UO_2902 (O_2902,N_49639,N_49873);
nor UO_2903 (O_2903,N_49153,N_49315);
or UO_2904 (O_2904,N_49069,N_49948);
and UO_2905 (O_2905,N_49199,N_49803);
and UO_2906 (O_2906,N_49776,N_49301);
nand UO_2907 (O_2907,N_49693,N_49044);
xor UO_2908 (O_2908,N_49307,N_49227);
and UO_2909 (O_2909,N_49115,N_49051);
nor UO_2910 (O_2910,N_49821,N_49760);
xnor UO_2911 (O_2911,N_49811,N_49855);
or UO_2912 (O_2912,N_49880,N_49798);
or UO_2913 (O_2913,N_49764,N_49433);
xor UO_2914 (O_2914,N_49843,N_49978);
nor UO_2915 (O_2915,N_49844,N_49976);
nand UO_2916 (O_2916,N_49138,N_49833);
xnor UO_2917 (O_2917,N_49592,N_49209);
xor UO_2918 (O_2918,N_49195,N_49804);
or UO_2919 (O_2919,N_49104,N_49459);
xor UO_2920 (O_2920,N_49542,N_49364);
or UO_2921 (O_2921,N_49284,N_49340);
or UO_2922 (O_2922,N_49693,N_49920);
and UO_2923 (O_2923,N_49581,N_49519);
and UO_2924 (O_2924,N_49071,N_49336);
xnor UO_2925 (O_2925,N_49052,N_49903);
nand UO_2926 (O_2926,N_49074,N_49364);
xnor UO_2927 (O_2927,N_49558,N_49840);
xnor UO_2928 (O_2928,N_49819,N_49332);
or UO_2929 (O_2929,N_49991,N_49723);
nor UO_2930 (O_2930,N_49377,N_49678);
nor UO_2931 (O_2931,N_49478,N_49379);
nand UO_2932 (O_2932,N_49572,N_49184);
nor UO_2933 (O_2933,N_49898,N_49277);
nand UO_2934 (O_2934,N_49090,N_49877);
and UO_2935 (O_2935,N_49202,N_49839);
nor UO_2936 (O_2936,N_49321,N_49051);
xor UO_2937 (O_2937,N_49408,N_49246);
nand UO_2938 (O_2938,N_49938,N_49120);
or UO_2939 (O_2939,N_49569,N_49431);
and UO_2940 (O_2940,N_49670,N_49009);
nand UO_2941 (O_2941,N_49821,N_49646);
nand UO_2942 (O_2942,N_49984,N_49741);
nor UO_2943 (O_2943,N_49567,N_49249);
nand UO_2944 (O_2944,N_49311,N_49785);
nand UO_2945 (O_2945,N_49562,N_49470);
or UO_2946 (O_2946,N_49363,N_49572);
nand UO_2947 (O_2947,N_49743,N_49027);
nor UO_2948 (O_2948,N_49510,N_49088);
xor UO_2949 (O_2949,N_49199,N_49191);
nor UO_2950 (O_2950,N_49650,N_49289);
nand UO_2951 (O_2951,N_49410,N_49613);
and UO_2952 (O_2952,N_49251,N_49577);
nor UO_2953 (O_2953,N_49352,N_49811);
nor UO_2954 (O_2954,N_49734,N_49687);
or UO_2955 (O_2955,N_49195,N_49734);
or UO_2956 (O_2956,N_49972,N_49792);
nor UO_2957 (O_2957,N_49695,N_49248);
or UO_2958 (O_2958,N_49249,N_49449);
and UO_2959 (O_2959,N_49663,N_49127);
nand UO_2960 (O_2960,N_49930,N_49278);
xor UO_2961 (O_2961,N_49649,N_49379);
xor UO_2962 (O_2962,N_49553,N_49084);
xor UO_2963 (O_2963,N_49035,N_49149);
nor UO_2964 (O_2964,N_49322,N_49097);
and UO_2965 (O_2965,N_49082,N_49619);
nand UO_2966 (O_2966,N_49790,N_49848);
nand UO_2967 (O_2967,N_49835,N_49870);
nand UO_2968 (O_2968,N_49985,N_49582);
nor UO_2969 (O_2969,N_49639,N_49255);
nor UO_2970 (O_2970,N_49827,N_49129);
or UO_2971 (O_2971,N_49328,N_49611);
and UO_2972 (O_2972,N_49502,N_49385);
xnor UO_2973 (O_2973,N_49385,N_49187);
xnor UO_2974 (O_2974,N_49965,N_49076);
or UO_2975 (O_2975,N_49581,N_49135);
nor UO_2976 (O_2976,N_49339,N_49478);
and UO_2977 (O_2977,N_49625,N_49624);
nand UO_2978 (O_2978,N_49426,N_49348);
nand UO_2979 (O_2979,N_49866,N_49804);
or UO_2980 (O_2980,N_49402,N_49874);
xor UO_2981 (O_2981,N_49627,N_49409);
and UO_2982 (O_2982,N_49184,N_49535);
or UO_2983 (O_2983,N_49449,N_49962);
and UO_2984 (O_2984,N_49839,N_49747);
nor UO_2985 (O_2985,N_49918,N_49580);
and UO_2986 (O_2986,N_49700,N_49134);
nand UO_2987 (O_2987,N_49818,N_49774);
nand UO_2988 (O_2988,N_49877,N_49432);
nand UO_2989 (O_2989,N_49588,N_49609);
and UO_2990 (O_2990,N_49129,N_49894);
xor UO_2991 (O_2991,N_49390,N_49712);
or UO_2992 (O_2992,N_49467,N_49203);
or UO_2993 (O_2993,N_49340,N_49665);
xor UO_2994 (O_2994,N_49028,N_49619);
or UO_2995 (O_2995,N_49867,N_49641);
xor UO_2996 (O_2996,N_49593,N_49422);
and UO_2997 (O_2997,N_49719,N_49597);
nor UO_2998 (O_2998,N_49981,N_49565);
nor UO_2999 (O_2999,N_49450,N_49756);
or UO_3000 (O_3000,N_49046,N_49436);
or UO_3001 (O_3001,N_49271,N_49767);
nor UO_3002 (O_3002,N_49479,N_49886);
xor UO_3003 (O_3003,N_49929,N_49958);
and UO_3004 (O_3004,N_49769,N_49275);
xor UO_3005 (O_3005,N_49619,N_49499);
xor UO_3006 (O_3006,N_49472,N_49440);
nor UO_3007 (O_3007,N_49525,N_49611);
or UO_3008 (O_3008,N_49598,N_49283);
or UO_3009 (O_3009,N_49456,N_49382);
or UO_3010 (O_3010,N_49140,N_49023);
nand UO_3011 (O_3011,N_49558,N_49128);
nand UO_3012 (O_3012,N_49993,N_49331);
and UO_3013 (O_3013,N_49116,N_49628);
or UO_3014 (O_3014,N_49724,N_49194);
nand UO_3015 (O_3015,N_49763,N_49494);
and UO_3016 (O_3016,N_49407,N_49794);
or UO_3017 (O_3017,N_49358,N_49450);
and UO_3018 (O_3018,N_49395,N_49325);
and UO_3019 (O_3019,N_49251,N_49339);
xnor UO_3020 (O_3020,N_49651,N_49707);
or UO_3021 (O_3021,N_49949,N_49929);
xor UO_3022 (O_3022,N_49183,N_49904);
nand UO_3023 (O_3023,N_49946,N_49845);
nand UO_3024 (O_3024,N_49038,N_49949);
xor UO_3025 (O_3025,N_49087,N_49220);
and UO_3026 (O_3026,N_49620,N_49802);
nand UO_3027 (O_3027,N_49950,N_49960);
xnor UO_3028 (O_3028,N_49687,N_49686);
xor UO_3029 (O_3029,N_49283,N_49878);
and UO_3030 (O_3030,N_49734,N_49759);
or UO_3031 (O_3031,N_49340,N_49530);
and UO_3032 (O_3032,N_49698,N_49568);
and UO_3033 (O_3033,N_49933,N_49880);
nand UO_3034 (O_3034,N_49615,N_49837);
or UO_3035 (O_3035,N_49317,N_49408);
xor UO_3036 (O_3036,N_49187,N_49887);
and UO_3037 (O_3037,N_49000,N_49749);
nor UO_3038 (O_3038,N_49584,N_49589);
nand UO_3039 (O_3039,N_49083,N_49708);
or UO_3040 (O_3040,N_49000,N_49405);
nand UO_3041 (O_3041,N_49531,N_49872);
and UO_3042 (O_3042,N_49153,N_49757);
nor UO_3043 (O_3043,N_49161,N_49776);
xnor UO_3044 (O_3044,N_49191,N_49129);
nor UO_3045 (O_3045,N_49399,N_49077);
xnor UO_3046 (O_3046,N_49370,N_49471);
xnor UO_3047 (O_3047,N_49144,N_49178);
and UO_3048 (O_3048,N_49030,N_49535);
or UO_3049 (O_3049,N_49383,N_49241);
nor UO_3050 (O_3050,N_49608,N_49191);
nand UO_3051 (O_3051,N_49778,N_49276);
xnor UO_3052 (O_3052,N_49310,N_49757);
and UO_3053 (O_3053,N_49967,N_49226);
nor UO_3054 (O_3054,N_49166,N_49640);
or UO_3055 (O_3055,N_49142,N_49926);
nand UO_3056 (O_3056,N_49209,N_49687);
and UO_3057 (O_3057,N_49253,N_49508);
nor UO_3058 (O_3058,N_49610,N_49068);
nand UO_3059 (O_3059,N_49275,N_49431);
nor UO_3060 (O_3060,N_49232,N_49322);
and UO_3061 (O_3061,N_49687,N_49731);
nor UO_3062 (O_3062,N_49050,N_49729);
xor UO_3063 (O_3063,N_49917,N_49611);
nand UO_3064 (O_3064,N_49990,N_49177);
nor UO_3065 (O_3065,N_49508,N_49803);
or UO_3066 (O_3066,N_49687,N_49966);
xnor UO_3067 (O_3067,N_49434,N_49411);
xnor UO_3068 (O_3068,N_49919,N_49582);
nand UO_3069 (O_3069,N_49528,N_49966);
xor UO_3070 (O_3070,N_49578,N_49273);
nand UO_3071 (O_3071,N_49046,N_49077);
nand UO_3072 (O_3072,N_49895,N_49609);
or UO_3073 (O_3073,N_49274,N_49356);
xnor UO_3074 (O_3074,N_49146,N_49983);
or UO_3075 (O_3075,N_49847,N_49046);
xnor UO_3076 (O_3076,N_49964,N_49837);
xnor UO_3077 (O_3077,N_49350,N_49432);
nor UO_3078 (O_3078,N_49025,N_49399);
nand UO_3079 (O_3079,N_49004,N_49560);
or UO_3080 (O_3080,N_49838,N_49516);
xor UO_3081 (O_3081,N_49406,N_49980);
nor UO_3082 (O_3082,N_49801,N_49511);
xor UO_3083 (O_3083,N_49938,N_49532);
or UO_3084 (O_3084,N_49643,N_49157);
and UO_3085 (O_3085,N_49491,N_49057);
nor UO_3086 (O_3086,N_49718,N_49362);
and UO_3087 (O_3087,N_49320,N_49897);
nand UO_3088 (O_3088,N_49965,N_49667);
nand UO_3089 (O_3089,N_49469,N_49377);
or UO_3090 (O_3090,N_49667,N_49034);
or UO_3091 (O_3091,N_49874,N_49810);
nor UO_3092 (O_3092,N_49353,N_49570);
nand UO_3093 (O_3093,N_49807,N_49260);
nor UO_3094 (O_3094,N_49587,N_49502);
nor UO_3095 (O_3095,N_49609,N_49316);
xnor UO_3096 (O_3096,N_49653,N_49945);
nand UO_3097 (O_3097,N_49441,N_49088);
nand UO_3098 (O_3098,N_49692,N_49883);
or UO_3099 (O_3099,N_49071,N_49993);
nor UO_3100 (O_3100,N_49675,N_49993);
nand UO_3101 (O_3101,N_49025,N_49569);
nand UO_3102 (O_3102,N_49895,N_49024);
or UO_3103 (O_3103,N_49649,N_49234);
xnor UO_3104 (O_3104,N_49560,N_49305);
and UO_3105 (O_3105,N_49070,N_49223);
and UO_3106 (O_3106,N_49791,N_49583);
nor UO_3107 (O_3107,N_49177,N_49301);
or UO_3108 (O_3108,N_49955,N_49990);
nor UO_3109 (O_3109,N_49043,N_49405);
nor UO_3110 (O_3110,N_49709,N_49023);
and UO_3111 (O_3111,N_49660,N_49303);
nor UO_3112 (O_3112,N_49307,N_49879);
nor UO_3113 (O_3113,N_49437,N_49774);
or UO_3114 (O_3114,N_49059,N_49944);
nor UO_3115 (O_3115,N_49939,N_49110);
and UO_3116 (O_3116,N_49391,N_49955);
xnor UO_3117 (O_3117,N_49393,N_49817);
nor UO_3118 (O_3118,N_49360,N_49529);
xnor UO_3119 (O_3119,N_49554,N_49167);
xor UO_3120 (O_3120,N_49264,N_49414);
and UO_3121 (O_3121,N_49605,N_49814);
or UO_3122 (O_3122,N_49492,N_49850);
nand UO_3123 (O_3123,N_49055,N_49627);
xor UO_3124 (O_3124,N_49478,N_49418);
xor UO_3125 (O_3125,N_49871,N_49651);
nor UO_3126 (O_3126,N_49500,N_49186);
nor UO_3127 (O_3127,N_49833,N_49346);
and UO_3128 (O_3128,N_49096,N_49568);
nor UO_3129 (O_3129,N_49509,N_49046);
or UO_3130 (O_3130,N_49610,N_49346);
or UO_3131 (O_3131,N_49659,N_49870);
nor UO_3132 (O_3132,N_49682,N_49042);
or UO_3133 (O_3133,N_49997,N_49860);
nand UO_3134 (O_3134,N_49728,N_49001);
or UO_3135 (O_3135,N_49909,N_49744);
nor UO_3136 (O_3136,N_49603,N_49617);
or UO_3137 (O_3137,N_49937,N_49756);
xnor UO_3138 (O_3138,N_49430,N_49611);
nand UO_3139 (O_3139,N_49960,N_49251);
nand UO_3140 (O_3140,N_49779,N_49541);
or UO_3141 (O_3141,N_49231,N_49805);
xnor UO_3142 (O_3142,N_49454,N_49341);
and UO_3143 (O_3143,N_49947,N_49777);
nor UO_3144 (O_3144,N_49410,N_49390);
nor UO_3145 (O_3145,N_49107,N_49796);
nor UO_3146 (O_3146,N_49793,N_49583);
nor UO_3147 (O_3147,N_49307,N_49501);
and UO_3148 (O_3148,N_49264,N_49024);
nand UO_3149 (O_3149,N_49207,N_49681);
or UO_3150 (O_3150,N_49755,N_49485);
and UO_3151 (O_3151,N_49104,N_49139);
xor UO_3152 (O_3152,N_49255,N_49548);
or UO_3153 (O_3153,N_49525,N_49968);
and UO_3154 (O_3154,N_49373,N_49267);
nand UO_3155 (O_3155,N_49991,N_49587);
xnor UO_3156 (O_3156,N_49275,N_49394);
or UO_3157 (O_3157,N_49601,N_49497);
xor UO_3158 (O_3158,N_49690,N_49199);
xor UO_3159 (O_3159,N_49175,N_49213);
xnor UO_3160 (O_3160,N_49020,N_49055);
and UO_3161 (O_3161,N_49714,N_49544);
or UO_3162 (O_3162,N_49946,N_49804);
xor UO_3163 (O_3163,N_49189,N_49310);
nor UO_3164 (O_3164,N_49823,N_49230);
nor UO_3165 (O_3165,N_49152,N_49967);
nand UO_3166 (O_3166,N_49454,N_49869);
or UO_3167 (O_3167,N_49862,N_49458);
nand UO_3168 (O_3168,N_49275,N_49761);
and UO_3169 (O_3169,N_49417,N_49603);
nand UO_3170 (O_3170,N_49686,N_49751);
or UO_3171 (O_3171,N_49782,N_49560);
and UO_3172 (O_3172,N_49840,N_49898);
nor UO_3173 (O_3173,N_49399,N_49692);
and UO_3174 (O_3174,N_49200,N_49689);
and UO_3175 (O_3175,N_49605,N_49319);
or UO_3176 (O_3176,N_49081,N_49029);
or UO_3177 (O_3177,N_49129,N_49027);
nor UO_3178 (O_3178,N_49081,N_49050);
nor UO_3179 (O_3179,N_49768,N_49248);
nand UO_3180 (O_3180,N_49303,N_49817);
nor UO_3181 (O_3181,N_49503,N_49376);
nand UO_3182 (O_3182,N_49629,N_49853);
and UO_3183 (O_3183,N_49145,N_49450);
or UO_3184 (O_3184,N_49326,N_49930);
and UO_3185 (O_3185,N_49472,N_49523);
nand UO_3186 (O_3186,N_49762,N_49127);
and UO_3187 (O_3187,N_49215,N_49567);
or UO_3188 (O_3188,N_49121,N_49980);
and UO_3189 (O_3189,N_49479,N_49540);
nand UO_3190 (O_3190,N_49310,N_49312);
xor UO_3191 (O_3191,N_49633,N_49604);
nor UO_3192 (O_3192,N_49402,N_49440);
and UO_3193 (O_3193,N_49820,N_49928);
nand UO_3194 (O_3194,N_49567,N_49388);
nor UO_3195 (O_3195,N_49693,N_49541);
nor UO_3196 (O_3196,N_49799,N_49925);
xor UO_3197 (O_3197,N_49765,N_49401);
xnor UO_3198 (O_3198,N_49239,N_49747);
or UO_3199 (O_3199,N_49309,N_49384);
nor UO_3200 (O_3200,N_49536,N_49384);
and UO_3201 (O_3201,N_49276,N_49512);
and UO_3202 (O_3202,N_49500,N_49374);
or UO_3203 (O_3203,N_49237,N_49116);
and UO_3204 (O_3204,N_49749,N_49363);
nand UO_3205 (O_3205,N_49858,N_49134);
xor UO_3206 (O_3206,N_49065,N_49966);
nor UO_3207 (O_3207,N_49932,N_49097);
or UO_3208 (O_3208,N_49675,N_49062);
or UO_3209 (O_3209,N_49665,N_49451);
or UO_3210 (O_3210,N_49277,N_49979);
or UO_3211 (O_3211,N_49381,N_49248);
and UO_3212 (O_3212,N_49249,N_49320);
or UO_3213 (O_3213,N_49242,N_49808);
and UO_3214 (O_3214,N_49169,N_49855);
nand UO_3215 (O_3215,N_49991,N_49182);
or UO_3216 (O_3216,N_49821,N_49041);
nor UO_3217 (O_3217,N_49100,N_49637);
nor UO_3218 (O_3218,N_49165,N_49181);
nor UO_3219 (O_3219,N_49447,N_49832);
or UO_3220 (O_3220,N_49221,N_49834);
or UO_3221 (O_3221,N_49914,N_49920);
or UO_3222 (O_3222,N_49607,N_49113);
xnor UO_3223 (O_3223,N_49419,N_49727);
or UO_3224 (O_3224,N_49639,N_49844);
xnor UO_3225 (O_3225,N_49926,N_49725);
or UO_3226 (O_3226,N_49160,N_49951);
xor UO_3227 (O_3227,N_49145,N_49138);
nand UO_3228 (O_3228,N_49129,N_49648);
nor UO_3229 (O_3229,N_49052,N_49814);
nand UO_3230 (O_3230,N_49920,N_49922);
xnor UO_3231 (O_3231,N_49121,N_49366);
xor UO_3232 (O_3232,N_49923,N_49559);
nor UO_3233 (O_3233,N_49173,N_49157);
and UO_3234 (O_3234,N_49141,N_49827);
nand UO_3235 (O_3235,N_49090,N_49476);
xor UO_3236 (O_3236,N_49985,N_49534);
and UO_3237 (O_3237,N_49452,N_49592);
and UO_3238 (O_3238,N_49306,N_49143);
or UO_3239 (O_3239,N_49785,N_49845);
nor UO_3240 (O_3240,N_49604,N_49731);
and UO_3241 (O_3241,N_49316,N_49378);
or UO_3242 (O_3242,N_49832,N_49738);
xnor UO_3243 (O_3243,N_49524,N_49183);
nand UO_3244 (O_3244,N_49975,N_49265);
xnor UO_3245 (O_3245,N_49797,N_49084);
or UO_3246 (O_3246,N_49627,N_49640);
and UO_3247 (O_3247,N_49155,N_49204);
xnor UO_3248 (O_3248,N_49963,N_49615);
and UO_3249 (O_3249,N_49023,N_49262);
nor UO_3250 (O_3250,N_49369,N_49659);
nand UO_3251 (O_3251,N_49256,N_49619);
and UO_3252 (O_3252,N_49916,N_49896);
nand UO_3253 (O_3253,N_49497,N_49763);
xor UO_3254 (O_3254,N_49023,N_49904);
and UO_3255 (O_3255,N_49537,N_49950);
xnor UO_3256 (O_3256,N_49173,N_49236);
nor UO_3257 (O_3257,N_49751,N_49045);
nand UO_3258 (O_3258,N_49160,N_49170);
nor UO_3259 (O_3259,N_49343,N_49288);
nor UO_3260 (O_3260,N_49709,N_49028);
nand UO_3261 (O_3261,N_49611,N_49303);
nor UO_3262 (O_3262,N_49947,N_49172);
xor UO_3263 (O_3263,N_49537,N_49251);
or UO_3264 (O_3264,N_49755,N_49564);
xor UO_3265 (O_3265,N_49751,N_49007);
nand UO_3266 (O_3266,N_49685,N_49391);
and UO_3267 (O_3267,N_49019,N_49527);
xor UO_3268 (O_3268,N_49659,N_49028);
nor UO_3269 (O_3269,N_49412,N_49784);
xnor UO_3270 (O_3270,N_49219,N_49245);
or UO_3271 (O_3271,N_49372,N_49774);
xor UO_3272 (O_3272,N_49480,N_49948);
nor UO_3273 (O_3273,N_49947,N_49374);
xnor UO_3274 (O_3274,N_49960,N_49367);
nand UO_3275 (O_3275,N_49344,N_49851);
and UO_3276 (O_3276,N_49214,N_49210);
nor UO_3277 (O_3277,N_49539,N_49111);
xor UO_3278 (O_3278,N_49060,N_49966);
nor UO_3279 (O_3279,N_49428,N_49661);
nand UO_3280 (O_3280,N_49532,N_49680);
nand UO_3281 (O_3281,N_49028,N_49117);
xor UO_3282 (O_3282,N_49594,N_49170);
nor UO_3283 (O_3283,N_49516,N_49758);
nor UO_3284 (O_3284,N_49106,N_49130);
nand UO_3285 (O_3285,N_49467,N_49024);
nor UO_3286 (O_3286,N_49276,N_49906);
xnor UO_3287 (O_3287,N_49670,N_49985);
nand UO_3288 (O_3288,N_49168,N_49563);
nand UO_3289 (O_3289,N_49049,N_49123);
xnor UO_3290 (O_3290,N_49526,N_49528);
xnor UO_3291 (O_3291,N_49911,N_49725);
and UO_3292 (O_3292,N_49208,N_49072);
xnor UO_3293 (O_3293,N_49202,N_49236);
nor UO_3294 (O_3294,N_49741,N_49792);
and UO_3295 (O_3295,N_49420,N_49567);
nor UO_3296 (O_3296,N_49048,N_49853);
and UO_3297 (O_3297,N_49215,N_49253);
xnor UO_3298 (O_3298,N_49504,N_49900);
xor UO_3299 (O_3299,N_49529,N_49771);
and UO_3300 (O_3300,N_49109,N_49055);
xnor UO_3301 (O_3301,N_49882,N_49859);
and UO_3302 (O_3302,N_49754,N_49706);
nor UO_3303 (O_3303,N_49508,N_49052);
or UO_3304 (O_3304,N_49118,N_49830);
nand UO_3305 (O_3305,N_49366,N_49018);
nand UO_3306 (O_3306,N_49309,N_49450);
or UO_3307 (O_3307,N_49055,N_49307);
nand UO_3308 (O_3308,N_49595,N_49552);
and UO_3309 (O_3309,N_49886,N_49665);
and UO_3310 (O_3310,N_49417,N_49501);
and UO_3311 (O_3311,N_49728,N_49651);
nand UO_3312 (O_3312,N_49281,N_49875);
xor UO_3313 (O_3313,N_49266,N_49901);
and UO_3314 (O_3314,N_49844,N_49662);
nand UO_3315 (O_3315,N_49026,N_49930);
nand UO_3316 (O_3316,N_49833,N_49491);
nor UO_3317 (O_3317,N_49321,N_49006);
nor UO_3318 (O_3318,N_49744,N_49273);
nand UO_3319 (O_3319,N_49565,N_49713);
nand UO_3320 (O_3320,N_49637,N_49633);
or UO_3321 (O_3321,N_49005,N_49216);
and UO_3322 (O_3322,N_49353,N_49625);
or UO_3323 (O_3323,N_49415,N_49143);
xor UO_3324 (O_3324,N_49708,N_49666);
xor UO_3325 (O_3325,N_49690,N_49123);
or UO_3326 (O_3326,N_49589,N_49941);
and UO_3327 (O_3327,N_49196,N_49019);
or UO_3328 (O_3328,N_49233,N_49504);
xnor UO_3329 (O_3329,N_49933,N_49048);
and UO_3330 (O_3330,N_49277,N_49680);
xnor UO_3331 (O_3331,N_49873,N_49277);
or UO_3332 (O_3332,N_49787,N_49848);
nand UO_3333 (O_3333,N_49425,N_49612);
or UO_3334 (O_3334,N_49494,N_49547);
or UO_3335 (O_3335,N_49961,N_49836);
nand UO_3336 (O_3336,N_49739,N_49021);
nand UO_3337 (O_3337,N_49186,N_49901);
xnor UO_3338 (O_3338,N_49305,N_49024);
nor UO_3339 (O_3339,N_49128,N_49650);
nand UO_3340 (O_3340,N_49728,N_49574);
xnor UO_3341 (O_3341,N_49468,N_49172);
nand UO_3342 (O_3342,N_49767,N_49685);
and UO_3343 (O_3343,N_49515,N_49762);
xnor UO_3344 (O_3344,N_49312,N_49898);
and UO_3345 (O_3345,N_49807,N_49106);
nor UO_3346 (O_3346,N_49544,N_49343);
nand UO_3347 (O_3347,N_49290,N_49816);
and UO_3348 (O_3348,N_49648,N_49394);
nand UO_3349 (O_3349,N_49714,N_49996);
nand UO_3350 (O_3350,N_49054,N_49615);
and UO_3351 (O_3351,N_49493,N_49555);
nor UO_3352 (O_3352,N_49240,N_49629);
nand UO_3353 (O_3353,N_49047,N_49893);
nor UO_3354 (O_3354,N_49406,N_49069);
nor UO_3355 (O_3355,N_49095,N_49962);
or UO_3356 (O_3356,N_49814,N_49635);
and UO_3357 (O_3357,N_49985,N_49717);
and UO_3358 (O_3358,N_49638,N_49487);
nor UO_3359 (O_3359,N_49208,N_49657);
nand UO_3360 (O_3360,N_49370,N_49198);
xor UO_3361 (O_3361,N_49931,N_49008);
xor UO_3362 (O_3362,N_49502,N_49507);
xor UO_3363 (O_3363,N_49618,N_49993);
xor UO_3364 (O_3364,N_49796,N_49142);
xnor UO_3365 (O_3365,N_49842,N_49602);
nand UO_3366 (O_3366,N_49311,N_49246);
nand UO_3367 (O_3367,N_49239,N_49678);
or UO_3368 (O_3368,N_49949,N_49690);
xor UO_3369 (O_3369,N_49926,N_49509);
nand UO_3370 (O_3370,N_49168,N_49275);
and UO_3371 (O_3371,N_49693,N_49994);
nor UO_3372 (O_3372,N_49200,N_49252);
or UO_3373 (O_3373,N_49936,N_49126);
nor UO_3374 (O_3374,N_49216,N_49353);
nand UO_3375 (O_3375,N_49888,N_49210);
and UO_3376 (O_3376,N_49778,N_49131);
nor UO_3377 (O_3377,N_49247,N_49806);
nand UO_3378 (O_3378,N_49339,N_49017);
or UO_3379 (O_3379,N_49656,N_49452);
xnor UO_3380 (O_3380,N_49708,N_49570);
or UO_3381 (O_3381,N_49737,N_49152);
or UO_3382 (O_3382,N_49500,N_49528);
nor UO_3383 (O_3383,N_49904,N_49601);
nand UO_3384 (O_3384,N_49290,N_49490);
or UO_3385 (O_3385,N_49922,N_49581);
and UO_3386 (O_3386,N_49130,N_49496);
and UO_3387 (O_3387,N_49767,N_49782);
nand UO_3388 (O_3388,N_49575,N_49215);
xor UO_3389 (O_3389,N_49213,N_49246);
nand UO_3390 (O_3390,N_49788,N_49726);
and UO_3391 (O_3391,N_49520,N_49125);
nor UO_3392 (O_3392,N_49999,N_49654);
or UO_3393 (O_3393,N_49644,N_49264);
nor UO_3394 (O_3394,N_49473,N_49861);
nand UO_3395 (O_3395,N_49992,N_49949);
or UO_3396 (O_3396,N_49588,N_49223);
or UO_3397 (O_3397,N_49355,N_49121);
or UO_3398 (O_3398,N_49984,N_49681);
nor UO_3399 (O_3399,N_49363,N_49404);
nor UO_3400 (O_3400,N_49381,N_49737);
nor UO_3401 (O_3401,N_49846,N_49134);
nand UO_3402 (O_3402,N_49080,N_49380);
nor UO_3403 (O_3403,N_49212,N_49658);
and UO_3404 (O_3404,N_49099,N_49960);
and UO_3405 (O_3405,N_49561,N_49134);
xor UO_3406 (O_3406,N_49682,N_49397);
nand UO_3407 (O_3407,N_49667,N_49843);
xnor UO_3408 (O_3408,N_49673,N_49119);
or UO_3409 (O_3409,N_49090,N_49192);
and UO_3410 (O_3410,N_49234,N_49553);
nor UO_3411 (O_3411,N_49905,N_49956);
nand UO_3412 (O_3412,N_49742,N_49060);
nor UO_3413 (O_3413,N_49053,N_49647);
or UO_3414 (O_3414,N_49299,N_49085);
nor UO_3415 (O_3415,N_49973,N_49524);
or UO_3416 (O_3416,N_49495,N_49729);
or UO_3417 (O_3417,N_49510,N_49580);
or UO_3418 (O_3418,N_49424,N_49682);
and UO_3419 (O_3419,N_49371,N_49974);
nor UO_3420 (O_3420,N_49767,N_49495);
and UO_3421 (O_3421,N_49492,N_49387);
xor UO_3422 (O_3422,N_49557,N_49520);
nand UO_3423 (O_3423,N_49421,N_49808);
xnor UO_3424 (O_3424,N_49938,N_49082);
nor UO_3425 (O_3425,N_49012,N_49191);
xnor UO_3426 (O_3426,N_49373,N_49030);
and UO_3427 (O_3427,N_49798,N_49594);
nor UO_3428 (O_3428,N_49343,N_49384);
and UO_3429 (O_3429,N_49509,N_49786);
or UO_3430 (O_3430,N_49026,N_49342);
nand UO_3431 (O_3431,N_49869,N_49623);
nor UO_3432 (O_3432,N_49372,N_49344);
xor UO_3433 (O_3433,N_49227,N_49016);
or UO_3434 (O_3434,N_49211,N_49748);
and UO_3435 (O_3435,N_49748,N_49347);
or UO_3436 (O_3436,N_49165,N_49881);
nand UO_3437 (O_3437,N_49638,N_49561);
nor UO_3438 (O_3438,N_49666,N_49359);
xnor UO_3439 (O_3439,N_49637,N_49285);
nand UO_3440 (O_3440,N_49355,N_49103);
nor UO_3441 (O_3441,N_49728,N_49122);
or UO_3442 (O_3442,N_49259,N_49905);
or UO_3443 (O_3443,N_49476,N_49773);
xor UO_3444 (O_3444,N_49920,N_49694);
or UO_3445 (O_3445,N_49123,N_49130);
xnor UO_3446 (O_3446,N_49251,N_49694);
xor UO_3447 (O_3447,N_49636,N_49348);
nand UO_3448 (O_3448,N_49329,N_49959);
or UO_3449 (O_3449,N_49403,N_49001);
xnor UO_3450 (O_3450,N_49357,N_49609);
or UO_3451 (O_3451,N_49540,N_49633);
or UO_3452 (O_3452,N_49709,N_49562);
nor UO_3453 (O_3453,N_49167,N_49533);
xor UO_3454 (O_3454,N_49073,N_49015);
and UO_3455 (O_3455,N_49471,N_49030);
or UO_3456 (O_3456,N_49715,N_49227);
xor UO_3457 (O_3457,N_49824,N_49111);
or UO_3458 (O_3458,N_49066,N_49718);
xnor UO_3459 (O_3459,N_49588,N_49859);
xor UO_3460 (O_3460,N_49365,N_49423);
or UO_3461 (O_3461,N_49639,N_49013);
nand UO_3462 (O_3462,N_49599,N_49705);
and UO_3463 (O_3463,N_49849,N_49938);
nand UO_3464 (O_3464,N_49944,N_49261);
and UO_3465 (O_3465,N_49792,N_49324);
nor UO_3466 (O_3466,N_49434,N_49289);
and UO_3467 (O_3467,N_49877,N_49567);
nand UO_3468 (O_3468,N_49184,N_49531);
or UO_3469 (O_3469,N_49047,N_49806);
and UO_3470 (O_3470,N_49360,N_49069);
and UO_3471 (O_3471,N_49760,N_49799);
and UO_3472 (O_3472,N_49433,N_49368);
or UO_3473 (O_3473,N_49817,N_49517);
xnor UO_3474 (O_3474,N_49403,N_49920);
or UO_3475 (O_3475,N_49669,N_49280);
nor UO_3476 (O_3476,N_49717,N_49536);
and UO_3477 (O_3477,N_49286,N_49497);
or UO_3478 (O_3478,N_49092,N_49491);
nor UO_3479 (O_3479,N_49747,N_49730);
xnor UO_3480 (O_3480,N_49846,N_49041);
nand UO_3481 (O_3481,N_49432,N_49944);
and UO_3482 (O_3482,N_49546,N_49623);
nand UO_3483 (O_3483,N_49100,N_49950);
and UO_3484 (O_3484,N_49050,N_49438);
or UO_3485 (O_3485,N_49090,N_49886);
or UO_3486 (O_3486,N_49816,N_49701);
and UO_3487 (O_3487,N_49345,N_49100);
and UO_3488 (O_3488,N_49050,N_49129);
xnor UO_3489 (O_3489,N_49363,N_49038);
xor UO_3490 (O_3490,N_49260,N_49783);
nand UO_3491 (O_3491,N_49163,N_49589);
or UO_3492 (O_3492,N_49144,N_49140);
or UO_3493 (O_3493,N_49813,N_49206);
or UO_3494 (O_3494,N_49959,N_49104);
nor UO_3495 (O_3495,N_49034,N_49357);
nand UO_3496 (O_3496,N_49155,N_49911);
and UO_3497 (O_3497,N_49865,N_49984);
or UO_3498 (O_3498,N_49277,N_49018);
and UO_3499 (O_3499,N_49261,N_49953);
nor UO_3500 (O_3500,N_49211,N_49666);
or UO_3501 (O_3501,N_49341,N_49469);
and UO_3502 (O_3502,N_49285,N_49068);
and UO_3503 (O_3503,N_49006,N_49746);
nor UO_3504 (O_3504,N_49226,N_49831);
or UO_3505 (O_3505,N_49787,N_49293);
or UO_3506 (O_3506,N_49905,N_49926);
xor UO_3507 (O_3507,N_49982,N_49463);
nor UO_3508 (O_3508,N_49009,N_49506);
nor UO_3509 (O_3509,N_49478,N_49621);
nand UO_3510 (O_3510,N_49416,N_49853);
nor UO_3511 (O_3511,N_49354,N_49029);
nand UO_3512 (O_3512,N_49775,N_49026);
nand UO_3513 (O_3513,N_49118,N_49435);
nand UO_3514 (O_3514,N_49019,N_49681);
nor UO_3515 (O_3515,N_49839,N_49832);
xnor UO_3516 (O_3516,N_49982,N_49867);
or UO_3517 (O_3517,N_49142,N_49654);
nor UO_3518 (O_3518,N_49116,N_49310);
xor UO_3519 (O_3519,N_49092,N_49742);
xnor UO_3520 (O_3520,N_49274,N_49780);
and UO_3521 (O_3521,N_49129,N_49630);
or UO_3522 (O_3522,N_49400,N_49528);
and UO_3523 (O_3523,N_49662,N_49591);
nand UO_3524 (O_3524,N_49074,N_49432);
xor UO_3525 (O_3525,N_49952,N_49484);
xor UO_3526 (O_3526,N_49682,N_49307);
or UO_3527 (O_3527,N_49415,N_49492);
nand UO_3528 (O_3528,N_49548,N_49667);
or UO_3529 (O_3529,N_49687,N_49809);
xor UO_3530 (O_3530,N_49450,N_49391);
and UO_3531 (O_3531,N_49032,N_49059);
xor UO_3532 (O_3532,N_49885,N_49362);
xnor UO_3533 (O_3533,N_49904,N_49009);
or UO_3534 (O_3534,N_49606,N_49542);
nor UO_3535 (O_3535,N_49534,N_49948);
and UO_3536 (O_3536,N_49100,N_49601);
nor UO_3537 (O_3537,N_49945,N_49774);
nor UO_3538 (O_3538,N_49704,N_49661);
xor UO_3539 (O_3539,N_49874,N_49258);
nor UO_3540 (O_3540,N_49558,N_49638);
xnor UO_3541 (O_3541,N_49385,N_49555);
nor UO_3542 (O_3542,N_49788,N_49305);
and UO_3543 (O_3543,N_49778,N_49006);
nand UO_3544 (O_3544,N_49570,N_49720);
or UO_3545 (O_3545,N_49216,N_49803);
xnor UO_3546 (O_3546,N_49489,N_49079);
and UO_3547 (O_3547,N_49424,N_49533);
nor UO_3548 (O_3548,N_49638,N_49216);
or UO_3549 (O_3549,N_49388,N_49082);
xor UO_3550 (O_3550,N_49466,N_49929);
and UO_3551 (O_3551,N_49836,N_49551);
or UO_3552 (O_3552,N_49182,N_49317);
or UO_3553 (O_3553,N_49179,N_49671);
nor UO_3554 (O_3554,N_49134,N_49613);
xnor UO_3555 (O_3555,N_49483,N_49281);
or UO_3556 (O_3556,N_49447,N_49121);
and UO_3557 (O_3557,N_49472,N_49950);
and UO_3558 (O_3558,N_49897,N_49184);
nand UO_3559 (O_3559,N_49422,N_49561);
xnor UO_3560 (O_3560,N_49548,N_49516);
and UO_3561 (O_3561,N_49875,N_49216);
nor UO_3562 (O_3562,N_49064,N_49089);
or UO_3563 (O_3563,N_49369,N_49364);
nand UO_3564 (O_3564,N_49380,N_49476);
xor UO_3565 (O_3565,N_49506,N_49128);
or UO_3566 (O_3566,N_49849,N_49233);
xnor UO_3567 (O_3567,N_49400,N_49001);
or UO_3568 (O_3568,N_49576,N_49152);
or UO_3569 (O_3569,N_49801,N_49772);
xor UO_3570 (O_3570,N_49221,N_49423);
nor UO_3571 (O_3571,N_49065,N_49688);
or UO_3572 (O_3572,N_49326,N_49378);
and UO_3573 (O_3573,N_49895,N_49386);
nand UO_3574 (O_3574,N_49024,N_49426);
nand UO_3575 (O_3575,N_49177,N_49951);
and UO_3576 (O_3576,N_49293,N_49698);
nor UO_3577 (O_3577,N_49635,N_49761);
xnor UO_3578 (O_3578,N_49829,N_49777);
and UO_3579 (O_3579,N_49043,N_49924);
or UO_3580 (O_3580,N_49050,N_49660);
nand UO_3581 (O_3581,N_49548,N_49817);
and UO_3582 (O_3582,N_49635,N_49874);
nand UO_3583 (O_3583,N_49821,N_49544);
xnor UO_3584 (O_3584,N_49059,N_49183);
nand UO_3585 (O_3585,N_49864,N_49367);
nand UO_3586 (O_3586,N_49247,N_49589);
and UO_3587 (O_3587,N_49843,N_49401);
nor UO_3588 (O_3588,N_49175,N_49202);
xor UO_3589 (O_3589,N_49943,N_49575);
and UO_3590 (O_3590,N_49792,N_49620);
and UO_3591 (O_3591,N_49541,N_49430);
and UO_3592 (O_3592,N_49787,N_49415);
nand UO_3593 (O_3593,N_49450,N_49767);
nor UO_3594 (O_3594,N_49301,N_49143);
xnor UO_3595 (O_3595,N_49930,N_49205);
and UO_3596 (O_3596,N_49020,N_49995);
nor UO_3597 (O_3597,N_49684,N_49211);
nand UO_3598 (O_3598,N_49759,N_49780);
nor UO_3599 (O_3599,N_49727,N_49322);
nor UO_3600 (O_3600,N_49185,N_49756);
nor UO_3601 (O_3601,N_49258,N_49729);
nand UO_3602 (O_3602,N_49498,N_49987);
and UO_3603 (O_3603,N_49250,N_49310);
nor UO_3604 (O_3604,N_49252,N_49764);
and UO_3605 (O_3605,N_49414,N_49383);
and UO_3606 (O_3606,N_49557,N_49707);
xnor UO_3607 (O_3607,N_49381,N_49332);
nor UO_3608 (O_3608,N_49640,N_49323);
nor UO_3609 (O_3609,N_49361,N_49089);
and UO_3610 (O_3610,N_49471,N_49297);
and UO_3611 (O_3611,N_49344,N_49339);
xnor UO_3612 (O_3612,N_49691,N_49197);
xor UO_3613 (O_3613,N_49594,N_49878);
and UO_3614 (O_3614,N_49746,N_49531);
nand UO_3615 (O_3615,N_49885,N_49657);
nor UO_3616 (O_3616,N_49911,N_49004);
nand UO_3617 (O_3617,N_49748,N_49518);
or UO_3618 (O_3618,N_49643,N_49417);
nand UO_3619 (O_3619,N_49923,N_49165);
and UO_3620 (O_3620,N_49928,N_49188);
xnor UO_3621 (O_3621,N_49816,N_49162);
or UO_3622 (O_3622,N_49617,N_49800);
nand UO_3623 (O_3623,N_49444,N_49844);
or UO_3624 (O_3624,N_49750,N_49994);
or UO_3625 (O_3625,N_49828,N_49488);
xor UO_3626 (O_3626,N_49735,N_49299);
xnor UO_3627 (O_3627,N_49126,N_49861);
nand UO_3628 (O_3628,N_49635,N_49577);
nand UO_3629 (O_3629,N_49136,N_49864);
and UO_3630 (O_3630,N_49221,N_49710);
and UO_3631 (O_3631,N_49741,N_49129);
nand UO_3632 (O_3632,N_49568,N_49199);
nor UO_3633 (O_3633,N_49772,N_49837);
nor UO_3634 (O_3634,N_49843,N_49716);
nand UO_3635 (O_3635,N_49024,N_49477);
nor UO_3636 (O_3636,N_49266,N_49424);
xor UO_3637 (O_3637,N_49427,N_49550);
nor UO_3638 (O_3638,N_49515,N_49348);
or UO_3639 (O_3639,N_49270,N_49876);
nor UO_3640 (O_3640,N_49236,N_49107);
or UO_3641 (O_3641,N_49454,N_49993);
nand UO_3642 (O_3642,N_49903,N_49124);
xnor UO_3643 (O_3643,N_49623,N_49659);
nand UO_3644 (O_3644,N_49296,N_49827);
nand UO_3645 (O_3645,N_49159,N_49289);
and UO_3646 (O_3646,N_49923,N_49018);
or UO_3647 (O_3647,N_49060,N_49167);
or UO_3648 (O_3648,N_49088,N_49009);
nand UO_3649 (O_3649,N_49754,N_49979);
and UO_3650 (O_3650,N_49084,N_49012);
or UO_3651 (O_3651,N_49816,N_49559);
or UO_3652 (O_3652,N_49986,N_49049);
nand UO_3653 (O_3653,N_49061,N_49168);
and UO_3654 (O_3654,N_49171,N_49615);
nor UO_3655 (O_3655,N_49530,N_49624);
or UO_3656 (O_3656,N_49694,N_49067);
and UO_3657 (O_3657,N_49749,N_49529);
or UO_3658 (O_3658,N_49827,N_49910);
or UO_3659 (O_3659,N_49849,N_49674);
or UO_3660 (O_3660,N_49425,N_49749);
or UO_3661 (O_3661,N_49306,N_49252);
xnor UO_3662 (O_3662,N_49793,N_49610);
nor UO_3663 (O_3663,N_49517,N_49105);
xor UO_3664 (O_3664,N_49388,N_49328);
nand UO_3665 (O_3665,N_49639,N_49815);
xnor UO_3666 (O_3666,N_49881,N_49949);
or UO_3667 (O_3667,N_49762,N_49774);
nand UO_3668 (O_3668,N_49307,N_49415);
and UO_3669 (O_3669,N_49869,N_49865);
nor UO_3670 (O_3670,N_49183,N_49587);
or UO_3671 (O_3671,N_49466,N_49594);
or UO_3672 (O_3672,N_49383,N_49582);
and UO_3673 (O_3673,N_49045,N_49470);
or UO_3674 (O_3674,N_49953,N_49705);
xor UO_3675 (O_3675,N_49554,N_49631);
nor UO_3676 (O_3676,N_49192,N_49528);
xnor UO_3677 (O_3677,N_49742,N_49592);
xnor UO_3678 (O_3678,N_49026,N_49646);
nor UO_3679 (O_3679,N_49814,N_49184);
or UO_3680 (O_3680,N_49008,N_49465);
and UO_3681 (O_3681,N_49162,N_49270);
nand UO_3682 (O_3682,N_49036,N_49888);
or UO_3683 (O_3683,N_49479,N_49366);
or UO_3684 (O_3684,N_49396,N_49751);
nand UO_3685 (O_3685,N_49157,N_49312);
nand UO_3686 (O_3686,N_49150,N_49141);
or UO_3687 (O_3687,N_49443,N_49686);
or UO_3688 (O_3688,N_49242,N_49593);
nor UO_3689 (O_3689,N_49348,N_49650);
nor UO_3690 (O_3690,N_49317,N_49114);
xnor UO_3691 (O_3691,N_49147,N_49537);
nor UO_3692 (O_3692,N_49270,N_49444);
xnor UO_3693 (O_3693,N_49079,N_49845);
nand UO_3694 (O_3694,N_49220,N_49117);
and UO_3695 (O_3695,N_49215,N_49735);
nand UO_3696 (O_3696,N_49229,N_49662);
and UO_3697 (O_3697,N_49908,N_49587);
nand UO_3698 (O_3698,N_49264,N_49586);
xnor UO_3699 (O_3699,N_49210,N_49084);
nand UO_3700 (O_3700,N_49298,N_49819);
nor UO_3701 (O_3701,N_49084,N_49150);
nor UO_3702 (O_3702,N_49770,N_49525);
or UO_3703 (O_3703,N_49104,N_49363);
and UO_3704 (O_3704,N_49653,N_49410);
nand UO_3705 (O_3705,N_49421,N_49162);
nor UO_3706 (O_3706,N_49383,N_49502);
nor UO_3707 (O_3707,N_49819,N_49080);
and UO_3708 (O_3708,N_49786,N_49777);
or UO_3709 (O_3709,N_49808,N_49103);
nand UO_3710 (O_3710,N_49589,N_49800);
xnor UO_3711 (O_3711,N_49422,N_49069);
or UO_3712 (O_3712,N_49243,N_49794);
nand UO_3713 (O_3713,N_49053,N_49883);
or UO_3714 (O_3714,N_49011,N_49551);
xnor UO_3715 (O_3715,N_49253,N_49583);
and UO_3716 (O_3716,N_49279,N_49905);
nand UO_3717 (O_3717,N_49948,N_49637);
or UO_3718 (O_3718,N_49220,N_49829);
or UO_3719 (O_3719,N_49181,N_49189);
xor UO_3720 (O_3720,N_49137,N_49431);
or UO_3721 (O_3721,N_49414,N_49389);
or UO_3722 (O_3722,N_49808,N_49078);
nand UO_3723 (O_3723,N_49610,N_49171);
xor UO_3724 (O_3724,N_49397,N_49615);
nor UO_3725 (O_3725,N_49863,N_49272);
nand UO_3726 (O_3726,N_49349,N_49795);
xor UO_3727 (O_3727,N_49657,N_49087);
nor UO_3728 (O_3728,N_49670,N_49974);
nand UO_3729 (O_3729,N_49237,N_49211);
nand UO_3730 (O_3730,N_49109,N_49959);
nand UO_3731 (O_3731,N_49071,N_49937);
xnor UO_3732 (O_3732,N_49273,N_49213);
nand UO_3733 (O_3733,N_49353,N_49705);
or UO_3734 (O_3734,N_49459,N_49695);
and UO_3735 (O_3735,N_49488,N_49151);
or UO_3736 (O_3736,N_49187,N_49174);
and UO_3737 (O_3737,N_49004,N_49425);
xor UO_3738 (O_3738,N_49330,N_49241);
and UO_3739 (O_3739,N_49722,N_49564);
nand UO_3740 (O_3740,N_49364,N_49745);
xnor UO_3741 (O_3741,N_49394,N_49674);
xor UO_3742 (O_3742,N_49625,N_49387);
xor UO_3743 (O_3743,N_49505,N_49504);
xor UO_3744 (O_3744,N_49102,N_49726);
or UO_3745 (O_3745,N_49208,N_49186);
nor UO_3746 (O_3746,N_49042,N_49636);
and UO_3747 (O_3747,N_49970,N_49643);
xor UO_3748 (O_3748,N_49978,N_49477);
or UO_3749 (O_3749,N_49623,N_49998);
or UO_3750 (O_3750,N_49279,N_49215);
or UO_3751 (O_3751,N_49285,N_49274);
nor UO_3752 (O_3752,N_49564,N_49103);
xor UO_3753 (O_3753,N_49375,N_49652);
xnor UO_3754 (O_3754,N_49894,N_49454);
and UO_3755 (O_3755,N_49456,N_49164);
or UO_3756 (O_3756,N_49777,N_49601);
xor UO_3757 (O_3757,N_49869,N_49296);
nor UO_3758 (O_3758,N_49731,N_49111);
nor UO_3759 (O_3759,N_49524,N_49678);
xor UO_3760 (O_3760,N_49259,N_49545);
nor UO_3761 (O_3761,N_49831,N_49204);
xnor UO_3762 (O_3762,N_49169,N_49952);
nor UO_3763 (O_3763,N_49700,N_49727);
xnor UO_3764 (O_3764,N_49878,N_49165);
nand UO_3765 (O_3765,N_49763,N_49270);
or UO_3766 (O_3766,N_49973,N_49941);
or UO_3767 (O_3767,N_49927,N_49961);
nor UO_3768 (O_3768,N_49389,N_49163);
nor UO_3769 (O_3769,N_49618,N_49874);
xnor UO_3770 (O_3770,N_49507,N_49381);
or UO_3771 (O_3771,N_49735,N_49494);
xor UO_3772 (O_3772,N_49173,N_49663);
and UO_3773 (O_3773,N_49589,N_49741);
xnor UO_3774 (O_3774,N_49222,N_49295);
or UO_3775 (O_3775,N_49262,N_49430);
nor UO_3776 (O_3776,N_49551,N_49809);
xnor UO_3777 (O_3777,N_49400,N_49016);
nor UO_3778 (O_3778,N_49767,N_49198);
xor UO_3779 (O_3779,N_49285,N_49469);
and UO_3780 (O_3780,N_49974,N_49225);
or UO_3781 (O_3781,N_49618,N_49807);
nand UO_3782 (O_3782,N_49408,N_49369);
nor UO_3783 (O_3783,N_49218,N_49022);
nor UO_3784 (O_3784,N_49529,N_49873);
xor UO_3785 (O_3785,N_49823,N_49476);
and UO_3786 (O_3786,N_49489,N_49512);
or UO_3787 (O_3787,N_49102,N_49099);
xnor UO_3788 (O_3788,N_49392,N_49396);
and UO_3789 (O_3789,N_49920,N_49883);
and UO_3790 (O_3790,N_49448,N_49309);
and UO_3791 (O_3791,N_49957,N_49378);
nor UO_3792 (O_3792,N_49160,N_49620);
nand UO_3793 (O_3793,N_49910,N_49027);
nand UO_3794 (O_3794,N_49929,N_49493);
and UO_3795 (O_3795,N_49318,N_49756);
and UO_3796 (O_3796,N_49052,N_49386);
nor UO_3797 (O_3797,N_49236,N_49949);
and UO_3798 (O_3798,N_49959,N_49225);
or UO_3799 (O_3799,N_49841,N_49782);
nand UO_3800 (O_3800,N_49487,N_49854);
xor UO_3801 (O_3801,N_49768,N_49986);
nand UO_3802 (O_3802,N_49145,N_49900);
or UO_3803 (O_3803,N_49676,N_49144);
or UO_3804 (O_3804,N_49023,N_49477);
xnor UO_3805 (O_3805,N_49471,N_49077);
or UO_3806 (O_3806,N_49705,N_49684);
and UO_3807 (O_3807,N_49174,N_49475);
xor UO_3808 (O_3808,N_49905,N_49616);
and UO_3809 (O_3809,N_49401,N_49428);
and UO_3810 (O_3810,N_49824,N_49391);
or UO_3811 (O_3811,N_49065,N_49556);
and UO_3812 (O_3812,N_49875,N_49749);
xnor UO_3813 (O_3813,N_49425,N_49598);
nor UO_3814 (O_3814,N_49654,N_49428);
xor UO_3815 (O_3815,N_49798,N_49043);
and UO_3816 (O_3816,N_49208,N_49412);
nor UO_3817 (O_3817,N_49429,N_49387);
nor UO_3818 (O_3818,N_49115,N_49734);
nor UO_3819 (O_3819,N_49457,N_49507);
or UO_3820 (O_3820,N_49904,N_49798);
xor UO_3821 (O_3821,N_49865,N_49666);
nand UO_3822 (O_3822,N_49513,N_49552);
nand UO_3823 (O_3823,N_49032,N_49533);
or UO_3824 (O_3824,N_49978,N_49679);
xnor UO_3825 (O_3825,N_49616,N_49026);
nand UO_3826 (O_3826,N_49277,N_49651);
xor UO_3827 (O_3827,N_49757,N_49835);
xor UO_3828 (O_3828,N_49473,N_49808);
or UO_3829 (O_3829,N_49276,N_49032);
nand UO_3830 (O_3830,N_49038,N_49756);
nand UO_3831 (O_3831,N_49524,N_49345);
nand UO_3832 (O_3832,N_49612,N_49284);
nor UO_3833 (O_3833,N_49617,N_49299);
xnor UO_3834 (O_3834,N_49045,N_49754);
xor UO_3835 (O_3835,N_49146,N_49413);
and UO_3836 (O_3836,N_49499,N_49212);
or UO_3837 (O_3837,N_49034,N_49584);
and UO_3838 (O_3838,N_49594,N_49137);
and UO_3839 (O_3839,N_49387,N_49317);
or UO_3840 (O_3840,N_49712,N_49816);
nor UO_3841 (O_3841,N_49375,N_49645);
nor UO_3842 (O_3842,N_49300,N_49889);
nand UO_3843 (O_3843,N_49180,N_49651);
and UO_3844 (O_3844,N_49552,N_49990);
xor UO_3845 (O_3845,N_49131,N_49102);
xor UO_3846 (O_3846,N_49072,N_49377);
or UO_3847 (O_3847,N_49548,N_49981);
nor UO_3848 (O_3848,N_49897,N_49295);
and UO_3849 (O_3849,N_49727,N_49935);
nor UO_3850 (O_3850,N_49278,N_49447);
or UO_3851 (O_3851,N_49189,N_49667);
or UO_3852 (O_3852,N_49431,N_49060);
or UO_3853 (O_3853,N_49993,N_49544);
and UO_3854 (O_3854,N_49064,N_49096);
or UO_3855 (O_3855,N_49880,N_49295);
nand UO_3856 (O_3856,N_49977,N_49453);
and UO_3857 (O_3857,N_49897,N_49398);
and UO_3858 (O_3858,N_49847,N_49028);
nor UO_3859 (O_3859,N_49995,N_49830);
xnor UO_3860 (O_3860,N_49275,N_49542);
nand UO_3861 (O_3861,N_49124,N_49686);
or UO_3862 (O_3862,N_49969,N_49889);
nand UO_3863 (O_3863,N_49646,N_49538);
nor UO_3864 (O_3864,N_49092,N_49432);
and UO_3865 (O_3865,N_49074,N_49886);
nand UO_3866 (O_3866,N_49699,N_49315);
or UO_3867 (O_3867,N_49906,N_49755);
or UO_3868 (O_3868,N_49063,N_49167);
or UO_3869 (O_3869,N_49505,N_49689);
xnor UO_3870 (O_3870,N_49812,N_49694);
nor UO_3871 (O_3871,N_49750,N_49081);
nor UO_3872 (O_3872,N_49911,N_49845);
and UO_3873 (O_3873,N_49307,N_49731);
nor UO_3874 (O_3874,N_49825,N_49601);
nand UO_3875 (O_3875,N_49337,N_49452);
xor UO_3876 (O_3876,N_49209,N_49708);
and UO_3877 (O_3877,N_49021,N_49761);
nor UO_3878 (O_3878,N_49016,N_49878);
or UO_3879 (O_3879,N_49966,N_49547);
nor UO_3880 (O_3880,N_49524,N_49341);
xnor UO_3881 (O_3881,N_49689,N_49888);
nor UO_3882 (O_3882,N_49826,N_49618);
or UO_3883 (O_3883,N_49867,N_49163);
and UO_3884 (O_3884,N_49046,N_49825);
nand UO_3885 (O_3885,N_49738,N_49535);
xnor UO_3886 (O_3886,N_49661,N_49022);
nand UO_3887 (O_3887,N_49339,N_49781);
nor UO_3888 (O_3888,N_49519,N_49637);
xnor UO_3889 (O_3889,N_49887,N_49404);
or UO_3890 (O_3890,N_49062,N_49169);
nand UO_3891 (O_3891,N_49751,N_49731);
and UO_3892 (O_3892,N_49282,N_49500);
nand UO_3893 (O_3893,N_49652,N_49538);
or UO_3894 (O_3894,N_49865,N_49628);
nand UO_3895 (O_3895,N_49781,N_49300);
xor UO_3896 (O_3896,N_49536,N_49751);
xor UO_3897 (O_3897,N_49438,N_49605);
nor UO_3898 (O_3898,N_49218,N_49597);
and UO_3899 (O_3899,N_49636,N_49217);
nand UO_3900 (O_3900,N_49595,N_49947);
nand UO_3901 (O_3901,N_49390,N_49087);
xnor UO_3902 (O_3902,N_49142,N_49696);
and UO_3903 (O_3903,N_49506,N_49788);
xnor UO_3904 (O_3904,N_49011,N_49104);
nand UO_3905 (O_3905,N_49532,N_49050);
xnor UO_3906 (O_3906,N_49215,N_49006);
xnor UO_3907 (O_3907,N_49762,N_49637);
and UO_3908 (O_3908,N_49999,N_49838);
nand UO_3909 (O_3909,N_49212,N_49081);
or UO_3910 (O_3910,N_49798,N_49238);
xnor UO_3911 (O_3911,N_49390,N_49655);
nand UO_3912 (O_3912,N_49147,N_49768);
nand UO_3913 (O_3913,N_49885,N_49738);
xnor UO_3914 (O_3914,N_49370,N_49352);
xor UO_3915 (O_3915,N_49042,N_49718);
and UO_3916 (O_3916,N_49858,N_49600);
or UO_3917 (O_3917,N_49049,N_49023);
xor UO_3918 (O_3918,N_49475,N_49689);
or UO_3919 (O_3919,N_49871,N_49090);
or UO_3920 (O_3920,N_49121,N_49443);
or UO_3921 (O_3921,N_49119,N_49514);
and UO_3922 (O_3922,N_49470,N_49776);
xor UO_3923 (O_3923,N_49284,N_49502);
and UO_3924 (O_3924,N_49237,N_49253);
and UO_3925 (O_3925,N_49207,N_49266);
or UO_3926 (O_3926,N_49646,N_49866);
nor UO_3927 (O_3927,N_49790,N_49450);
or UO_3928 (O_3928,N_49299,N_49238);
or UO_3929 (O_3929,N_49205,N_49422);
nand UO_3930 (O_3930,N_49550,N_49029);
xor UO_3931 (O_3931,N_49934,N_49181);
nor UO_3932 (O_3932,N_49278,N_49428);
or UO_3933 (O_3933,N_49498,N_49471);
nand UO_3934 (O_3934,N_49380,N_49370);
nand UO_3935 (O_3935,N_49881,N_49586);
and UO_3936 (O_3936,N_49345,N_49302);
and UO_3937 (O_3937,N_49232,N_49444);
nor UO_3938 (O_3938,N_49482,N_49359);
nor UO_3939 (O_3939,N_49747,N_49884);
or UO_3940 (O_3940,N_49636,N_49560);
and UO_3941 (O_3941,N_49221,N_49496);
nand UO_3942 (O_3942,N_49666,N_49018);
xnor UO_3943 (O_3943,N_49114,N_49118);
and UO_3944 (O_3944,N_49847,N_49946);
nor UO_3945 (O_3945,N_49342,N_49915);
xnor UO_3946 (O_3946,N_49474,N_49711);
or UO_3947 (O_3947,N_49653,N_49433);
nor UO_3948 (O_3948,N_49042,N_49719);
nand UO_3949 (O_3949,N_49645,N_49907);
nand UO_3950 (O_3950,N_49559,N_49069);
nand UO_3951 (O_3951,N_49555,N_49146);
xnor UO_3952 (O_3952,N_49594,N_49201);
nand UO_3953 (O_3953,N_49574,N_49074);
nor UO_3954 (O_3954,N_49813,N_49744);
and UO_3955 (O_3955,N_49125,N_49293);
xor UO_3956 (O_3956,N_49593,N_49495);
and UO_3957 (O_3957,N_49553,N_49750);
nor UO_3958 (O_3958,N_49098,N_49425);
nand UO_3959 (O_3959,N_49509,N_49702);
nor UO_3960 (O_3960,N_49925,N_49350);
xnor UO_3961 (O_3961,N_49390,N_49853);
or UO_3962 (O_3962,N_49171,N_49879);
xor UO_3963 (O_3963,N_49646,N_49757);
nor UO_3964 (O_3964,N_49521,N_49844);
nor UO_3965 (O_3965,N_49676,N_49536);
nor UO_3966 (O_3966,N_49509,N_49848);
nor UO_3967 (O_3967,N_49944,N_49635);
and UO_3968 (O_3968,N_49495,N_49172);
nor UO_3969 (O_3969,N_49961,N_49232);
or UO_3970 (O_3970,N_49517,N_49192);
xor UO_3971 (O_3971,N_49514,N_49059);
nor UO_3972 (O_3972,N_49927,N_49632);
and UO_3973 (O_3973,N_49520,N_49488);
nand UO_3974 (O_3974,N_49156,N_49145);
nor UO_3975 (O_3975,N_49436,N_49145);
nor UO_3976 (O_3976,N_49037,N_49838);
xnor UO_3977 (O_3977,N_49882,N_49376);
or UO_3978 (O_3978,N_49299,N_49067);
nor UO_3979 (O_3979,N_49472,N_49117);
nor UO_3980 (O_3980,N_49100,N_49701);
nand UO_3981 (O_3981,N_49237,N_49516);
xor UO_3982 (O_3982,N_49819,N_49216);
and UO_3983 (O_3983,N_49088,N_49570);
or UO_3984 (O_3984,N_49227,N_49638);
or UO_3985 (O_3985,N_49044,N_49416);
nand UO_3986 (O_3986,N_49653,N_49458);
nand UO_3987 (O_3987,N_49165,N_49877);
xor UO_3988 (O_3988,N_49835,N_49673);
and UO_3989 (O_3989,N_49480,N_49982);
xor UO_3990 (O_3990,N_49711,N_49443);
or UO_3991 (O_3991,N_49542,N_49214);
and UO_3992 (O_3992,N_49903,N_49891);
nor UO_3993 (O_3993,N_49202,N_49698);
nor UO_3994 (O_3994,N_49658,N_49101);
nor UO_3995 (O_3995,N_49986,N_49171);
and UO_3996 (O_3996,N_49759,N_49945);
xor UO_3997 (O_3997,N_49220,N_49809);
and UO_3998 (O_3998,N_49432,N_49937);
or UO_3999 (O_3999,N_49613,N_49792);
nand UO_4000 (O_4000,N_49865,N_49224);
nor UO_4001 (O_4001,N_49405,N_49790);
and UO_4002 (O_4002,N_49283,N_49117);
nand UO_4003 (O_4003,N_49863,N_49413);
nand UO_4004 (O_4004,N_49161,N_49998);
or UO_4005 (O_4005,N_49085,N_49285);
nand UO_4006 (O_4006,N_49184,N_49499);
nand UO_4007 (O_4007,N_49107,N_49085);
and UO_4008 (O_4008,N_49130,N_49388);
and UO_4009 (O_4009,N_49435,N_49433);
xnor UO_4010 (O_4010,N_49926,N_49877);
and UO_4011 (O_4011,N_49737,N_49301);
nand UO_4012 (O_4012,N_49193,N_49359);
and UO_4013 (O_4013,N_49712,N_49891);
nor UO_4014 (O_4014,N_49787,N_49505);
nand UO_4015 (O_4015,N_49908,N_49420);
xnor UO_4016 (O_4016,N_49171,N_49219);
or UO_4017 (O_4017,N_49842,N_49924);
and UO_4018 (O_4018,N_49468,N_49311);
and UO_4019 (O_4019,N_49211,N_49103);
nand UO_4020 (O_4020,N_49958,N_49396);
nor UO_4021 (O_4021,N_49640,N_49558);
xnor UO_4022 (O_4022,N_49195,N_49987);
or UO_4023 (O_4023,N_49639,N_49111);
or UO_4024 (O_4024,N_49958,N_49909);
xnor UO_4025 (O_4025,N_49719,N_49424);
and UO_4026 (O_4026,N_49093,N_49550);
xor UO_4027 (O_4027,N_49192,N_49613);
xor UO_4028 (O_4028,N_49061,N_49560);
or UO_4029 (O_4029,N_49126,N_49273);
nand UO_4030 (O_4030,N_49747,N_49408);
or UO_4031 (O_4031,N_49028,N_49804);
and UO_4032 (O_4032,N_49386,N_49519);
nand UO_4033 (O_4033,N_49590,N_49947);
or UO_4034 (O_4034,N_49337,N_49308);
and UO_4035 (O_4035,N_49196,N_49026);
nand UO_4036 (O_4036,N_49336,N_49769);
and UO_4037 (O_4037,N_49219,N_49803);
nor UO_4038 (O_4038,N_49026,N_49982);
and UO_4039 (O_4039,N_49085,N_49485);
or UO_4040 (O_4040,N_49628,N_49402);
and UO_4041 (O_4041,N_49766,N_49708);
or UO_4042 (O_4042,N_49672,N_49361);
and UO_4043 (O_4043,N_49485,N_49374);
nor UO_4044 (O_4044,N_49766,N_49412);
xor UO_4045 (O_4045,N_49961,N_49814);
nor UO_4046 (O_4046,N_49528,N_49354);
nor UO_4047 (O_4047,N_49070,N_49838);
xor UO_4048 (O_4048,N_49098,N_49582);
or UO_4049 (O_4049,N_49009,N_49745);
nor UO_4050 (O_4050,N_49844,N_49278);
nor UO_4051 (O_4051,N_49298,N_49144);
nand UO_4052 (O_4052,N_49634,N_49278);
or UO_4053 (O_4053,N_49449,N_49176);
nand UO_4054 (O_4054,N_49291,N_49003);
xor UO_4055 (O_4055,N_49855,N_49522);
and UO_4056 (O_4056,N_49642,N_49690);
and UO_4057 (O_4057,N_49757,N_49778);
nor UO_4058 (O_4058,N_49116,N_49739);
or UO_4059 (O_4059,N_49976,N_49698);
nand UO_4060 (O_4060,N_49957,N_49914);
and UO_4061 (O_4061,N_49563,N_49282);
or UO_4062 (O_4062,N_49122,N_49455);
xnor UO_4063 (O_4063,N_49385,N_49956);
xnor UO_4064 (O_4064,N_49925,N_49248);
or UO_4065 (O_4065,N_49460,N_49962);
or UO_4066 (O_4066,N_49488,N_49786);
nor UO_4067 (O_4067,N_49025,N_49688);
nand UO_4068 (O_4068,N_49169,N_49209);
and UO_4069 (O_4069,N_49879,N_49398);
nor UO_4070 (O_4070,N_49857,N_49649);
or UO_4071 (O_4071,N_49811,N_49649);
or UO_4072 (O_4072,N_49501,N_49477);
nand UO_4073 (O_4073,N_49575,N_49081);
nand UO_4074 (O_4074,N_49064,N_49168);
or UO_4075 (O_4075,N_49059,N_49787);
or UO_4076 (O_4076,N_49413,N_49433);
nor UO_4077 (O_4077,N_49558,N_49275);
and UO_4078 (O_4078,N_49643,N_49848);
and UO_4079 (O_4079,N_49407,N_49585);
xnor UO_4080 (O_4080,N_49013,N_49285);
xnor UO_4081 (O_4081,N_49197,N_49258);
nor UO_4082 (O_4082,N_49191,N_49341);
and UO_4083 (O_4083,N_49850,N_49950);
and UO_4084 (O_4084,N_49172,N_49152);
xnor UO_4085 (O_4085,N_49140,N_49308);
xnor UO_4086 (O_4086,N_49540,N_49197);
nor UO_4087 (O_4087,N_49151,N_49567);
xnor UO_4088 (O_4088,N_49387,N_49061);
or UO_4089 (O_4089,N_49054,N_49678);
and UO_4090 (O_4090,N_49785,N_49953);
nand UO_4091 (O_4091,N_49549,N_49908);
xnor UO_4092 (O_4092,N_49508,N_49673);
or UO_4093 (O_4093,N_49836,N_49869);
nand UO_4094 (O_4094,N_49931,N_49322);
and UO_4095 (O_4095,N_49695,N_49777);
nand UO_4096 (O_4096,N_49579,N_49702);
nor UO_4097 (O_4097,N_49842,N_49038);
or UO_4098 (O_4098,N_49506,N_49455);
xnor UO_4099 (O_4099,N_49722,N_49861);
and UO_4100 (O_4100,N_49704,N_49601);
nor UO_4101 (O_4101,N_49488,N_49433);
xor UO_4102 (O_4102,N_49335,N_49410);
or UO_4103 (O_4103,N_49119,N_49780);
xor UO_4104 (O_4104,N_49888,N_49431);
or UO_4105 (O_4105,N_49024,N_49350);
xnor UO_4106 (O_4106,N_49918,N_49723);
nand UO_4107 (O_4107,N_49238,N_49066);
xor UO_4108 (O_4108,N_49424,N_49312);
and UO_4109 (O_4109,N_49552,N_49832);
xnor UO_4110 (O_4110,N_49345,N_49227);
nor UO_4111 (O_4111,N_49820,N_49035);
and UO_4112 (O_4112,N_49066,N_49454);
nand UO_4113 (O_4113,N_49549,N_49147);
or UO_4114 (O_4114,N_49468,N_49719);
or UO_4115 (O_4115,N_49555,N_49850);
nand UO_4116 (O_4116,N_49528,N_49610);
nand UO_4117 (O_4117,N_49660,N_49613);
or UO_4118 (O_4118,N_49083,N_49382);
or UO_4119 (O_4119,N_49543,N_49266);
or UO_4120 (O_4120,N_49167,N_49273);
nor UO_4121 (O_4121,N_49095,N_49606);
and UO_4122 (O_4122,N_49327,N_49255);
xnor UO_4123 (O_4123,N_49493,N_49189);
xnor UO_4124 (O_4124,N_49215,N_49704);
nand UO_4125 (O_4125,N_49093,N_49322);
and UO_4126 (O_4126,N_49107,N_49034);
nand UO_4127 (O_4127,N_49373,N_49818);
nand UO_4128 (O_4128,N_49185,N_49096);
or UO_4129 (O_4129,N_49149,N_49965);
nand UO_4130 (O_4130,N_49526,N_49200);
and UO_4131 (O_4131,N_49590,N_49741);
and UO_4132 (O_4132,N_49405,N_49725);
and UO_4133 (O_4133,N_49024,N_49460);
and UO_4134 (O_4134,N_49793,N_49110);
nand UO_4135 (O_4135,N_49321,N_49762);
nand UO_4136 (O_4136,N_49516,N_49720);
nor UO_4137 (O_4137,N_49925,N_49785);
or UO_4138 (O_4138,N_49516,N_49575);
and UO_4139 (O_4139,N_49258,N_49436);
xnor UO_4140 (O_4140,N_49028,N_49685);
nand UO_4141 (O_4141,N_49554,N_49175);
and UO_4142 (O_4142,N_49926,N_49835);
nand UO_4143 (O_4143,N_49068,N_49318);
or UO_4144 (O_4144,N_49232,N_49537);
nor UO_4145 (O_4145,N_49986,N_49054);
and UO_4146 (O_4146,N_49860,N_49917);
or UO_4147 (O_4147,N_49115,N_49899);
xor UO_4148 (O_4148,N_49458,N_49320);
xor UO_4149 (O_4149,N_49403,N_49386);
xor UO_4150 (O_4150,N_49472,N_49475);
xnor UO_4151 (O_4151,N_49339,N_49217);
nand UO_4152 (O_4152,N_49581,N_49566);
xnor UO_4153 (O_4153,N_49899,N_49426);
nor UO_4154 (O_4154,N_49233,N_49827);
and UO_4155 (O_4155,N_49128,N_49388);
nor UO_4156 (O_4156,N_49488,N_49225);
nor UO_4157 (O_4157,N_49960,N_49127);
and UO_4158 (O_4158,N_49087,N_49242);
and UO_4159 (O_4159,N_49262,N_49072);
or UO_4160 (O_4160,N_49336,N_49008);
nand UO_4161 (O_4161,N_49703,N_49575);
nand UO_4162 (O_4162,N_49555,N_49652);
and UO_4163 (O_4163,N_49860,N_49212);
nor UO_4164 (O_4164,N_49187,N_49339);
nor UO_4165 (O_4165,N_49143,N_49223);
xor UO_4166 (O_4166,N_49186,N_49487);
nand UO_4167 (O_4167,N_49084,N_49316);
and UO_4168 (O_4168,N_49408,N_49924);
nand UO_4169 (O_4169,N_49724,N_49993);
nor UO_4170 (O_4170,N_49930,N_49107);
nor UO_4171 (O_4171,N_49511,N_49410);
nand UO_4172 (O_4172,N_49048,N_49949);
nor UO_4173 (O_4173,N_49152,N_49662);
nand UO_4174 (O_4174,N_49072,N_49398);
or UO_4175 (O_4175,N_49820,N_49749);
nand UO_4176 (O_4176,N_49666,N_49781);
and UO_4177 (O_4177,N_49883,N_49251);
or UO_4178 (O_4178,N_49752,N_49602);
and UO_4179 (O_4179,N_49818,N_49029);
or UO_4180 (O_4180,N_49340,N_49946);
xor UO_4181 (O_4181,N_49594,N_49033);
xnor UO_4182 (O_4182,N_49220,N_49610);
nor UO_4183 (O_4183,N_49864,N_49107);
nand UO_4184 (O_4184,N_49148,N_49070);
or UO_4185 (O_4185,N_49360,N_49005);
nor UO_4186 (O_4186,N_49125,N_49863);
nor UO_4187 (O_4187,N_49709,N_49557);
or UO_4188 (O_4188,N_49307,N_49368);
and UO_4189 (O_4189,N_49597,N_49119);
nand UO_4190 (O_4190,N_49244,N_49110);
and UO_4191 (O_4191,N_49450,N_49682);
or UO_4192 (O_4192,N_49455,N_49420);
and UO_4193 (O_4193,N_49395,N_49632);
and UO_4194 (O_4194,N_49019,N_49797);
and UO_4195 (O_4195,N_49722,N_49478);
and UO_4196 (O_4196,N_49964,N_49884);
nor UO_4197 (O_4197,N_49623,N_49194);
xnor UO_4198 (O_4198,N_49445,N_49287);
nor UO_4199 (O_4199,N_49470,N_49496);
nor UO_4200 (O_4200,N_49317,N_49597);
and UO_4201 (O_4201,N_49039,N_49984);
xnor UO_4202 (O_4202,N_49313,N_49661);
or UO_4203 (O_4203,N_49901,N_49497);
nand UO_4204 (O_4204,N_49577,N_49531);
or UO_4205 (O_4205,N_49057,N_49670);
nor UO_4206 (O_4206,N_49608,N_49288);
nor UO_4207 (O_4207,N_49250,N_49179);
nor UO_4208 (O_4208,N_49934,N_49293);
and UO_4209 (O_4209,N_49136,N_49721);
nor UO_4210 (O_4210,N_49705,N_49605);
and UO_4211 (O_4211,N_49911,N_49380);
or UO_4212 (O_4212,N_49107,N_49848);
nand UO_4213 (O_4213,N_49763,N_49589);
nand UO_4214 (O_4214,N_49856,N_49872);
nor UO_4215 (O_4215,N_49985,N_49397);
nand UO_4216 (O_4216,N_49736,N_49205);
xor UO_4217 (O_4217,N_49191,N_49825);
xnor UO_4218 (O_4218,N_49145,N_49567);
or UO_4219 (O_4219,N_49053,N_49502);
or UO_4220 (O_4220,N_49037,N_49345);
nand UO_4221 (O_4221,N_49766,N_49245);
and UO_4222 (O_4222,N_49201,N_49084);
and UO_4223 (O_4223,N_49913,N_49364);
nand UO_4224 (O_4224,N_49305,N_49831);
xor UO_4225 (O_4225,N_49555,N_49291);
and UO_4226 (O_4226,N_49704,N_49194);
and UO_4227 (O_4227,N_49274,N_49295);
and UO_4228 (O_4228,N_49726,N_49634);
and UO_4229 (O_4229,N_49944,N_49456);
nand UO_4230 (O_4230,N_49502,N_49249);
nand UO_4231 (O_4231,N_49148,N_49663);
or UO_4232 (O_4232,N_49427,N_49470);
nor UO_4233 (O_4233,N_49191,N_49913);
nand UO_4234 (O_4234,N_49368,N_49650);
nor UO_4235 (O_4235,N_49282,N_49617);
and UO_4236 (O_4236,N_49220,N_49741);
nor UO_4237 (O_4237,N_49597,N_49861);
or UO_4238 (O_4238,N_49338,N_49233);
nor UO_4239 (O_4239,N_49916,N_49331);
xnor UO_4240 (O_4240,N_49357,N_49696);
nand UO_4241 (O_4241,N_49529,N_49730);
nand UO_4242 (O_4242,N_49696,N_49102);
xnor UO_4243 (O_4243,N_49743,N_49790);
nor UO_4244 (O_4244,N_49293,N_49989);
nand UO_4245 (O_4245,N_49691,N_49864);
nand UO_4246 (O_4246,N_49805,N_49860);
xnor UO_4247 (O_4247,N_49819,N_49265);
xor UO_4248 (O_4248,N_49468,N_49768);
or UO_4249 (O_4249,N_49469,N_49943);
and UO_4250 (O_4250,N_49231,N_49831);
xnor UO_4251 (O_4251,N_49525,N_49805);
or UO_4252 (O_4252,N_49906,N_49122);
xnor UO_4253 (O_4253,N_49400,N_49440);
nand UO_4254 (O_4254,N_49139,N_49414);
xnor UO_4255 (O_4255,N_49655,N_49778);
nand UO_4256 (O_4256,N_49759,N_49127);
nand UO_4257 (O_4257,N_49737,N_49009);
xnor UO_4258 (O_4258,N_49307,N_49373);
xnor UO_4259 (O_4259,N_49409,N_49090);
nor UO_4260 (O_4260,N_49212,N_49464);
xnor UO_4261 (O_4261,N_49224,N_49156);
or UO_4262 (O_4262,N_49642,N_49355);
nand UO_4263 (O_4263,N_49346,N_49048);
or UO_4264 (O_4264,N_49148,N_49762);
xor UO_4265 (O_4265,N_49389,N_49474);
nand UO_4266 (O_4266,N_49940,N_49927);
and UO_4267 (O_4267,N_49607,N_49408);
and UO_4268 (O_4268,N_49041,N_49977);
nand UO_4269 (O_4269,N_49092,N_49659);
or UO_4270 (O_4270,N_49705,N_49227);
or UO_4271 (O_4271,N_49490,N_49559);
or UO_4272 (O_4272,N_49750,N_49637);
and UO_4273 (O_4273,N_49605,N_49124);
and UO_4274 (O_4274,N_49285,N_49151);
and UO_4275 (O_4275,N_49707,N_49588);
and UO_4276 (O_4276,N_49347,N_49979);
nor UO_4277 (O_4277,N_49183,N_49517);
nand UO_4278 (O_4278,N_49149,N_49651);
or UO_4279 (O_4279,N_49546,N_49917);
xor UO_4280 (O_4280,N_49482,N_49396);
nor UO_4281 (O_4281,N_49596,N_49914);
xor UO_4282 (O_4282,N_49230,N_49949);
and UO_4283 (O_4283,N_49025,N_49796);
and UO_4284 (O_4284,N_49067,N_49473);
and UO_4285 (O_4285,N_49099,N_49847);
nor UO_4286 (O_4286,N_49567,N_49234);
nor UO_4287 (O_4287,N_49815,N_49331);
nor UO_4288 (O_4288,N_49730,N_49604);
or UO_4289 (O_4289,N_49679,N_49746);
nor UO_4290 (O_4290,N_49821,N_49113);
and UO_4291 (O_4291,N_49707,N_49419);
or UO_4292 (O_4292,N_49026,N_49814);
or UO_4293 (O_4293,N_49851,N_49291);
and UO_4294 (O_4294,N_49736,N_49252);
nand UO_4295 (O_4295,N_49406,N_49567);
and UO_4296 (O_4296,N_49505,N_49914);
nor UO_4297 (O_4297,N_49832,N_49487);
and UO_4298 (O_4298,N_49627,N_49897);
and UO_4299 (O_4299,N_49206,N_49963);
nor UO_4300 (O_4300,N_49236,N_49274);
or UO_4301 (O_4301,N_49382,N_49577);
nand UO_4302 (O_4302,N_49378,N_49562);
nor UO_4303 (O_4303,N_49644,N_49249);
xnor UO_4304 (O_4304,N_49512,N_49011);
nor UO_4305 (O_4305,N_49205,N_49181);
nand UO_4306 (O_4306,N_49721,N_49085);
nor UO_4307 (O_4307,N_49182,N_49542);
and UO_4308 (O_4308,N_49125,N_49871);
nand UO_4309 (O_4309,N_49109,N_49742);
nand UO_4310 (O_4310,N_49331,N_49243);
nor UO_4311 (O_4311,N_49075,N_49628);
nor UO_4312 (O_4312,N_49885,N_49572);
or UO_4313 (O_4313,N_49031,N_49530);
nand UO_4314 (O_4314,N_49916,N_49275);
and UO_4315 (O_4315,N_49537,N_49014);
nand UO_4316 (O_4316,N_49562,N_49896);
and UO_4317 (O_4317,N_49996,N_49062);
or UO_4318 (O_4318,N_49087,N_49732);
nor UO_4319 (O_4319,N_49072,N_49934);
or UO_4320 (O_4320,N_49021,N_49660);
nor UO_4321 (O_4321,N_49960,N_49405);
xnor UO_4322 (O_4322,N_49812,N_49535);
nand UO_4323 (O_4323,N_49308,N_49063);
or UO_4324 (O_4324,N_49704,N_49176);
and UO_4325 (O_4325,N_49853,N_49354);
or UO_4326 (O_4326,N_49680,N_49485);
or UO_4327 (O_4327,N_49810,N_49709);
or UO_4328 (O_4328,N_49280,N_49253);
and UO_4329 (O_4329,N_49150,N_49228);
and UO_4330 (O_4330,N_49578,N_49067);
xor UO_4331 (O_4331,N_49982,N_49470);
or UO_4332 (O_4332,N_49616,N_49483);
xnor UO_4333 (O_4333,N_49987,N_49071);
nor UO_4334 (O_4334,N_49758,N_49207);
or UO_4335 (O_4335,N_49172,N_49095);
or UO_4336 (O_4336,N_49374,N_49392);
or UO_4337 (O_4337,N_49519,N_49688);
and UO_4338 (O_4338,N_49376,N_49951);
or UO_4339 (O_4339,N_49943,N_49812);
xnor UO_4340 (O_4340,N_49730,N_49046);
nand UO_4341 (O_4341,N_49713,N_49966);
nand UO_4342 (O_4342,N_49115,N_49021);
and UO_4343 (O_4343,N_49203,N_49557);
or UO_4344 (O_4344,N_49544,N_49195);
or UO_4345 (O_4345,N_49876,N_49981);
and UO_4346 (O_4346,N_49072,N_49549);
xor UO_4347 (O_4347,N_49969,N_49395);
and UO_4348 (O_4348,N_49660,N_49558);
and UO_4349 (O_4349,N_49305,N_49572);
xnor UO_4350 (O_4350,N_49055,N_49024);
or UO_4351 (O_4351,N_49161,N_49243);
nand UO_4352 (O_4352,N_49919,N_49924);
or UO_4353 (O_4353,N_49637,N_49333);
nor UO_4354 (O_4354,N_49459,N_49399);
and UO_4355 (O_4355,N_49599,N_49326);
nand UO_4356 (O_4356,N_49806,N_49451);
nor UO_4357 (O_4357,N_49566,N_49077);
nand UO_4358 (O_4358,N_49538,N_49562);
or UO_4359 (O_4359,N_49362,N_49320);
nand UO_4360 (O_4360,N_49409,N_49441);
xnor UO_4361 (O_4361,N_49004,N_49685);
nand UO_4362 (O_4362,N_49415,N_49645);
nand UO_4363 (O_4363,N_49474,N_49766);
nor UO_4364 (O_4364,N_49401,N_49036);
or UO_4365 (O_4365,N_49411,N_49854);
and UO_4366 (O_4366,N_49215,N_49617);
nand UO_4367 (O_4367,N_49449,N_49008);
and UO_4368 (O_4368,N_49271,N_49455);
and UO_4369 (O_4369,N_49685,N_49814);
or UO_4370 (O_4370,N_49024,N_49377);
and UO_4371 (O_4371,N_49075,N_49881);
xnor UO_4372 (O_4372,N_49142,N_49137);
or UO_4373 (O_4373,N_49695,N_49999);
xnor UO_4374 (O_4374,N_49982,N_49066);
nand UO_4375 (O_4375,N_49908,N_49574);
nand UO_4376 (O_4376,N_49013,N_49573);
xor UO_4377 (O_4377,N_49106,N_49190);
nand UO_4378 (O_4378,N_49841,N_49784);
nand UO_4379 (O_4379,N_49591,N_49303);
and UO_4380 (O_4380,N_49701,N_49428);
nand UO_4381 (O_4381,N_49452,N_49845);
and UO_4382 (O_4382,N_49395,N_49210);
or UO_4383 (O_4383,N_49052,N_49377);
xor UO_4384 (O_4384,N_49487,N_49229);
nor UO_4385 (O_4385,N_49221,N_49768);
nand UO_4386 (O_4386,N_49998,N_49115);
and UO_4387 (O_4387,N_49160,N_49206);
nor UO_4388 (O_4388,N_49928,N_49313);
and UO_4389 (O_4389,N_49908,N_49302);
xnor UO_4390 (O_4390,N_49283,N_49275);
nand UO_4391 (O_4391,N_49605,N_49916);
xor UO_4392 (O_4392,N_49939,N_49970);
xor UO_4393 (O_4393,N_49660,N_49301);
or UO_4394 (O_4394,N_49320,N_49901);
or UO_4395 (O_4395,N_49825,N_49536);
nor UO_4396 (O_4396,N_49005,N_49458);
xnor UO_4397 (O_4397,N_49562,N_49419);
nand UO_4398 (O_4398,N_49308,N_49028);
xor UO_4399 (O_4399,N_49738,N_49670);
or UO_4400 (O_4400,N_49175,N_49485);
xnor UO_4401 (O_4401,N_49509,N_49013);
nor UO_4402 (O_4402,N_49085,N_49775);
xnor UO_4403 (O_4403,N_49955,N_49042);
nor UO_4404 (O_4404,N_49006,N_49821);
and UO_4405 (O_4405,N_49182,N_49802);
or UO_4406 (O_4406,N_49912,N_49545);
and UO_4407 (O_4407,N_49834,N_49217);
nor UO_4408 (O_4408,N_49161,N_49595);
nand UO_4409 (O_4409,N_49831,N_49595);
and UO_4410 (O_4410,N_49896,N_49875);
or UO_4411 (O_4411,N_49588,N_49470);
and UO_4412 (O_4412,N_49752,N_49466);
nor UO_4413 (O_4413,N_49109,N_49462);
xnor UO_4414 (O_4414,N_49637,N_49243);
nand UO_4415 (O_4415,N_49334,N_49413);
nand UO_4416 (O_4416,N_49069,N_49554);
and UO_4417 (O_4417,N_49221,N_49935);
nor UO_4418 (O_4418,N_49220,N_49706);
nand UO_4419 (O_4419,N_49685,N_49778);
nand UO_4420 (O_4420,N_49480,N_49799);
and UO_4421 (O_4421,N_49966,N_49529);
nor UO_4422 (O_4422,N_49602,N_49247);
or UO_4423 (O_4423,N_49583,N_49915);
and UO_4424 (O_4424,N_49777,N_49447);
xor UO_4425 (O_4425,N_49875,N_49290);
xnor UO_4426 (O_4426,N_49427,N_49649);
nor UO_4427 (O_4427,N_49184,N_49903);
xor UO_4428 (O_4428,N_49470,N_49959);
nand UO_4429 (O_4429,N_49742,N_49676);
xor UO_4430 (O_4430,N_49992,N_49486);
or UO_4431 (O_4431,N_49504,N_49859);
and UO_4432 (O_4432,N_49485,N_49229);
or UO_4433 (O_4433,N_49509,N_49785);
nand UO_4434 (O_4434,N_49449,N_49490);
xor UO_4435 (O_4435,N_49364,N_49423);
xnor UO_4436 (O_4436,N_49241,N_49069);
or UO_4437 (O_4437,N_49061,N_49693);
nor UO_4438 (O_4438,N_49733,N_49120);
nor UO_4439 (O_4439,N_49837,N_49639);
nand UO_4440 (O_4440,N_49853,N_49081);
or UO_4441 (O_4441,N_49386,N_49905);
nand UO_4442 (O_4442,N_49684,N_49882);
or UO_4443 (O_4443,N_49574,N_49957);
or UO_4444 (O_4444,N_49324,N_49805);
xnor UO_4445 (O_4445,N_49916,N_49472);
nor UO_4446 (O_4446,N_49075,N_49712);
nand UO_4447 (O_4447,N_49265,N_49339);
nand UO_4448 (O_4448,N_49338,N_49550);
or UO_4449 (O_4449,N_49975,N_49775);
or UO_4450 (O_4450,N_49465,N_49984);
nand UO_4451 (O_4451,N_49425,N_49212);
nand UO_4452 (O_4452,N_49151,N_49098);
and UO_4453 (O_4453,N_49612,N_49972);
or UO_4454 (O_4454,N_49946,N_49234);
nor UO_4455 (O_4455,N_49286,N_49256);
and UO_4456 (O_4456,N_49800,N_49946);
xor UO_4457 (O_4457,N_49933,N_49039);
and UO_4458 (O_4458,N_49068,N_49126);
nand UO_4459 (O_4459,N_49386,N_49580);
nor UO_4460 (O_4460,N_49731,N_49958);
or UO_4461 (O_4461,N_49937,N_49170);
nand UO_4462 (O_4462,N_49762,N_49065);
nand UO_4463 (O_4463,N_49947,N_49372);
and UO_4464 (O_4464,N_49750,N_49030);
nor UO_4465 (O_4465,N_49256,N_49155);
and UO_4466 (O_4466,N_49166,N_49920);
or UO_4467 (O_4467,N_49432,N_49292);
nor UO_4468 (O_4468,N_49138,N_49127);
or UO_4469 (O_4469,N_49969,N_49940);
nor UO_4470 (O_4470,N_49465,N_49339);
or UO_4471 (O_4471,N_49285,N_49503);
and UO_4472 (O_4472,N_49493,N_49344);
nand UO_4473 (O_4473,N_49449,N_49778);
nor UO_4474 (O_4474,N_49618,N_49576);
nand UO_4475 (O_4475,N_49803,N_49043);
nand UO_4476 (O_4476,N_49471,N_49380);
nand UO_4477 (O_4477,N_49595,N_49265);
nand UO_4478 (O_4478,N_49102,N_49172);
or UO_4479 (O_4479,N_49530,N_49728);
xnor UO_4480 (O_4480,N_49454,N_49206);
or UO_4481 (O_4481,N_49008,N_49580);
xor UO_4482 (O_4482,N_49174,N_49104);
or UO_4483 (O_4483,N_49713,N_49735);
nor UO_4484 (O_4484,N_49044,N_49284);
nand UO_4485 (O_4485,N_49657,N_49210);
or UO_4486 (O_4486,N_49198,N_49648);
xor UO_4487 (O_4487,N_49053,N_49097);
nor UO_4488 (O_4488,N_49520,N_49243);
nor UO_4489 (O_4489,N_49733,N_49074);
nand UO_4490 (O_4490,N_49822,N_49824);
nor UO_4491 (O_4491,N_49307,N_49961);
or UO_4492 (O_4492,N_49651,N_49373);
nor UO_4493 (O_4493,N_49200,N_49708);
or UO_4494 (O_4494,N_49441,N_49304);
nor UO_4495 (O_4495,N_49422,N_49919);
nor UO_4496 (O_4496,N_49011,N_49067);
xor UO_4497 (O_4497,N_49960,N_49363);
xor UO_4498 (O_4498,N_49403,N_49668);
xor UO_4499 (O_4499,N_49762,N_49918);
and UO_4500 (O_4500,N_49594,N_49342);
and UO_4501 (O_4501,N_49669,N_49678);
nand UO_4502 (O_4502,N_49805,N_49144);
nor UO_4503 (O_4503,N_49211,N_49436);
xnor UO_4504 (O_4504,N_49219,N_49537);
and UO_4505 (O_4505,N_49556,N_49691);
xor UO_4506 (O_4506,N_49318,N_49873);
and UO_4507 (O_4507,N_49738,N_49106);
nor UO_4508 (O_4508,N_49297,N_49534);
or UO_4509 (O_4509,N_49913,N_49230);
and UO_4510 (O_4510,N_49491,N_49908);
nor UO_4511 (O_4511,N_49686,N_49299);
nand UO_4512 (O_4512,N_49108,N_49493);
xnor UO_4513 (O_4513,N_49269,N_49159);
or UO_4514 (O_4514,N_49773,N_49211);
or UO_4515 (O_4515,N_49205,N_49548);
nand UO_4516 (O_4516,N_49053,N_49076);
and UO_4517 (O_4517,N_49317,N_49991);
or UO_4518 (O_4518,N_49007,N_49809);
or UO_4519 (O_4519,N_49850,N_49300);
and UO_4520 (O_4520,N_49252,N_49594);
nand UO_4521 (O_4521,N_49807,N_49833);
nor UO_4522 (O_4522,N_49201,N_49820);
xnor UO_4523 (O_4523,N_49763,N_49997);
nor UO_4524 (O_4524,N_49572,N_49324);
and UO_4525 (O_4525,N_49196,N_49056);
nand UO_4526 (O_4526,N_49801,N_49974);
nor UO_4527 (O_4527,N_49312,N_49005);
nand UO_4528 (O_4528,N_49858,N_49081);
nand UO_4529 (O_4529,N_49730,N_49169);
nand UO_4530 (O_4530,N_49731,N_49851);
nand UO_4531 (O_4531,N_49741,N_49578);
nand UO_4532 (O_4532,N_49589,N_49099);
nand UO_4533 (O_4533,N_49309,N_49352);
xor UO_4534 (O_4534,N_49741,N_49675);
nand UO_4535 (O_4535,N_49943,N_49605);
xnor UO_4536 (O_4536,N_49607,N_49108);
nor UO_4537 (O_4537,N_49108,N_49763);
or UO_4538 (O_4538,N_49051,N_49149);
xnor UO_4539 (O_4539,N_49747,N_49880);
nand UO_4540 (O_4540,N_49060,N_49016);
xnor UO_4541 (O_4541,N_49673,N_49202);
or UO_4542 (O_4542,N_49089,N_49220);
nor UO_4543 (O_4543,N_49240,N_49386);
nand UO_4544 (O_4544,N_49101,N_49288);
nor UO_4545 (O_4545,N_49650,N_49172);
xnor UO_4546 (O_4546,N_49153,N_49921);
nand UO_4547 (O_4547,N_49089,N_49820);
or UO_4548 (O_4548,N_49826,N_49912);
and UO_4549 (O_4549,N_49208,N_49891);
xor UO_4550 (O_4550,N_49706,N_49502);
xnor UO_4551 (O_4551,N_49371,N_49035);
xor UO_4552 (O_4552,N_49360,N_49056);
or UO_4553 (O_4553,N_49561,N_49763);
or UO_4554 (O_4554,N_49648,N_49427);
xnor UO_4555 (O_4555,N_49865,N_49379);
or UO_4556 (O_4556,N_49990,N_49560);
nor UO_4557 (O_4557,N_49113,N_49775);
nor UO_4558 (O_4558,N_49718,N_49318);
or UO_4559 (O_4559,N_49842,N_49063);
or UO_4560 (O_4560,N_49781,N_49502);
and UO_4561 (O_4561,N_49311,N_49626);
xor UO_4562 (O_4562,N_49698,N_49761);
nor UO_4563 (O_4563,N_49729,N_49224);
and UO_4564 (O_4564,N_49423,N_49407);
or UO_4565 (O_4565,N_49475,N_49100);
or UO_4566 (O_4566,N_49425,N_49141);
xor UO_4567 (O_4567,N_49986,N_49813);
nand UO_4568 (O_4568,N_49159,N_49441);
and UO_4569 (O_4569,N_49574,N_49509);
nor UO_4570 (O_4570,N_49570,N_49132);
and UO_4571 (O_4571,N_49056,N_49577);
nor UO_4572 (O_4572,N_49026,N_49563);
and UO_4573 (O_4573,N_49316,N_49634);
nand UO_4574 (O_4574,N_49263,N_49707);
or UO_4575 (O_4575,N_49539,N_49020);
or UO_4576 (O_4576,N_49197,N_49092);
nor UO_4577 (O_4577,N_49150,N_49391);
or UO_4578 (O_4578,N_49486,N_49079);
nor UO_4579 (O_4579,N_49164,N_49061);
and UO_4580 (O_4580,N_49960,N_49956);
xor UO_4581 (O_4581,N_49607,N_49203);
nand UO_4582 (O_4582,N_49739,N_49076);
or UO_4583 (O_4583,N_49918,N_49964);
nand UO_4584 (O_4584,N_49106,N_49293);
and UO_4585 (O_4585,N_49392,N_49781);
xnor UO_4586 (O_4586,N_49265,N_49685);
and UO_4587 (O_4587,N_49844,N_49738);
nor UO_4588 (O_4588,N_49407,N_49086);
nand UO_4589 (O_4589,N_49074,N_49841);
and UO_4590 (O_4590,N_49768,N_49852);
nand UO_4591 (O_4591,N_49765,N_49309);
nor UO_4592 (O_4592,N_49406,N_49704);
xor UO_4593 (O_4593,N_49565,N_49482);
or UO_4594 (O_4594,N_49319,N_49688);
nor UO_4595 (O_4595,N_49917,N_49368);
nand UO_4596 (O_4596,N_49883,N_49734);
and UO_4597 (O_4597,N_49592,N_49355);
xnor UO_4598 (O_4598,N_49952,N_49684);
or UO_4599 (O_4599,N_49678,N_49084);
nor UO_4600 (O_4600,N_49337,N_49105);
nand UO_4601 (O_4601,N_49032,N_49425);
xnor UO_4602 (O_4602,N_49940,N_49912);
or UO_4603 (O_4603,N_49771,N_49427);
nand UO_4604 (O_4604,N_49439,N_49076);
or UO_4605 (O_4605,N_49473,N_49585);
nor UO_4606 (O_4606,N_49428,N_49457);
or UO_4607 (O_4607,N_49695,N_49783);
xnor UO_4608 (O_4608,N_49896,N_49081);
and UO_4609 (O_4609,N_49303,N_49948);
or UO_4610 (O_4610,N_49445,N_49673);
or UO_4611 (O_4611,N_49703,N_49384);
and UO_4612 (O_4612,N_49397,N_49712);
xor UO_4613 (O_4613,N_49552,N_49488);
or UO_4614 (O_4614,N_49310,N_49601);
nor UO_4615 (O_4615,N_49149,N_49052);
nor UO_4616 (O_4616,N_49887,N_49845);
nor UO_4617 (O_4617,N_49001,N_49151);
and UO_4618 (O_4618,N_49096,N_49706);
and UO_4619 (O_4619,N_49434,N_49639);
or UO_4620 (O_4620,N_49167,N_49475);
nor UO_4621 (O_4621,N_49910,N_49984);
xor UO_4622 (O_4622,N_49465,N_49835);
or UO_4623 (O_4623,N_49381,N_49825);
xor UO_4624 (O_4624,N_49867,N_49325);
nand UO_4625 (O_4625,N_49304,N_49769);
xnor UO_4626 (O_4626,N_49282,N_49959);
or UO_4627 (O_4627,N_49441,N_49235);
or UO_4628 (O_4628,N_49104,N_49931);
nand UO_4629 (O_4629,N_49234,N_49230);
xor UO_4630 (O_4630,N_49060,N_49080);
and UO_4631 (O_4631,N_49252,N_49553);
nand UO_4632 (O_4632,N_49099,N_49700);
xnor UO_4633 (O_4633,N_49454,N_49591);
nor UO_4634 (O_4634,N_49680,N_49930);
nand UO_4635 (O_4635,N_49565,N_49452);
or UO_4636 (O_4636,N_49526,N_49616);
xor UO_4637 (O_4637,N_49485,N_49959);
or UO_4638 (O_4638,N_49382,N_49686);
and UO_4639 (O_4639,N_49950,N_49633);
nand UO_4640 (O_4640,N_49804,N_49509);
or UO_4641 (O_4641,N_49178,N_49448);
xnor UO_4642 (O_4642,N_49291,N_49739);
and UO_4643 (O_4643,N_49781,N_49587);
and UO_4644 (O_4644,N_49711,N_49526);
or UO_4645 (O_4645,N_49993,N_49329);
and UO_4646 (O_4646,N_49119,N_49680);
and UO_4647 (O_4647,N_49182,N_49981);
or UO_4648 (O_4648,N_49124,N_49403);
nor UO_4649 (O_4649,N_49027,N_49510);
nand UO_4650 (O_4650,N_49673,N_49027);
nand UO_4651 (O_4651,N_49261,N_49532);
or UO_4652 (O_4652,N_49820,N_49845);
or UO_4653 (O_4653,N_49801,N_49494);
and UO_4654 (O_4654,N_49263,N_49298);
nor UO_4655 (O_4655,N_49489,N_49162);
nand UO_4656 (O_4656,N_49938,N_49832);
xnor UO_4657 (O_4657,N_49938,N_49416);
xnor UO_4658 (O_4658,N_49986,N_49902);
and UO_4659 (O_4659,N_49804,N_49776);
nor UO_4660 (O_4660,N_49821,N_49057);
or UO_4661 (O_4661,N_49391,N_49782);
nand UO_4662 (O_4662,N_49468,N_49689);
xnor UO_4663 (O_4663,N_49838,N_49531);
nand UO_4664 (O_4664,N_49255,N_49318);
xnor UO_4665 (O_4665,N_49862,N_49999);
nor UO_4666 (O_4666,N_49897,N_49079);
and UO_4667 (O_4667,N_49984,N_49395);
and UO_4668 (O_4668,N_49970,N_49392);
nand UO_4669 (O_4669,N_49642,N_49986);
and UO_4670 (O_4670,N_49470,N_49051);
nor UO_4671 (O_4671,N_49015,N_49192);
xnor UO_4672 (O_4672,N_49818,N_49295);
and UO_4673 (O_4673,N_49765,N_49769);
nor UO_4674 (O_4674,N_49347,N_49505);
xor UO_4675 (O_4675,N_49211,N_49753);
xnor UO_4676 (O_4676,N_49662,N_49391);
and UO_4677 (O_4677,N_49394,N_49926);
nor UO_4678 (O_4678,N_49721,N_49338);
xor UO_4679 (O_4679,N_49547,N_49074);
or UO_4680 (O_4680,N_49820,N_49279);
nor UO_4681 (O_4681,N_49522,N_49011);
nand UO_4682 (O_4682,N_49858,N_49449);
xnor UO_4683 (O_4683,N_49274,N_49794);
or UO_4684 (O_4684,N_49004,N_49994);
xor UO_4685 (O_4685,N_49571,N_49529);
and UO_4686 (O_4686,N_49394,N_49603);
nor UO_4687 (O_4687,N_49639,N_49603);
nand UO_4688 (O_4688,N_49071,N_49396);
or UO_4689 (O_4689,N_49928,N_49956);
and UO_4690 (O_4690,N_49485,N_49413);
nor UO_4691 (O_4691,N_49647,N_49615);
or UO_4692 (O_4692,N_49994,N_49707);
and UO_4693 (O_4693,N_49499,N_49823);
or UO_4694 (O_4694,N_49335,N_49729);
or UO_4695 (O_4695,N_49426,N_49032);
or UO_4696 (O_4696,N_49124,N_49706);
xnor UO_4697 (O_4697,N_49197,N_49240);
xnor UO_4698 (O_4698,N_49239,N_49623);
or UO_4699 (O_4699,N_49215,N_49999);
nor UO_4700 (O_4700,N_49724,N_49423);
or UO_4701 (O_4701,N_49755,N_49369);
nor UO_4702 (O_4702,N_49422,N_49657);
nand UO_4703 (O_4703,N_49860,N_49346);
nor UO_4704 (O_4704,N_49275,N_49594);
or UO_4705 (O_4705,N_49339,N_49565);
nor UO_4706 (O_4706,N_49723,N_49397);
and UO_4707 (O_4707,N_49389,N_49274);
nor UO_4708 (O_4708,N_49322,N_49653);
nand UO_4709 (O_4709,N_49090,N_49616);
nand UO_4710 (O_4710,N_49197,N_49532);
and UO_4711 (O_4711,N_49506,N_49510);
xnor UO_4712 (O_4712,N_49400,N_49921);
and UO_4713 (O_4713,N_49386,N_49523);
nand UO_4714 (O_4714,N_49751,N_49074);
or UO_4715 (O_4715,N_49654,N_49047);
and UO_4716 (O_4716,N_49675,N_49426);
nand UO_4717 (O_4717,N_49324,N_49670);
or UO_4718 (O_4718,N_49766,N_49814);
xnor UO_4719 (O_4719,N_49440,N_49485);
and UO_4720 (O_4720,N_49538,N_49697);
and UO_4721 (O_4721,N_49548,N_49623);
xnor UO_4722 (O_4722,N_49420,N_49647);
nand UO_4723 (O_4723,N_49032,N_49984);
and UO_4724 (O_4724,N_49007,N_49158);
nand UO_4725 (O_4725,N_49195,N_49686);
nand UO_4726 (O_4726,N_49365,N_49182);
xnor UO_4727 (O_4727,N_49692,N_49581);
xor UO_4728 (O_4728,N_49109,N_49728);
xor UO_4729 (O_4729,N_49622,N_49564);
and UO_4730 (O_4730,N_49912,N_49385);
or UO_4731 (O_4731,N_49888,N_49351);
or UO_4732 (O_4732,N_49297,N_49243);
nor UO_4733 (O_4733,N_49304,N_49179);
and UO_4734 (O_4734,N_49384,N_49503);
nand UO_4735 (O_4735,N_49548,N_49147);
xnor UO_4736 (O_4736,N_49758,N_49240);
xnor UO_4737 (O_4737,N_49265,N_49169);
nor UO_4738 (O_4738,N_49740,N_49798);
or UO_4739 (O_4739,N_49786,N_49515);
nor UO_4740 (O_4740,N_49408,N_49590);
xnor UO_4741 (O_4741,N_49037,N_49451);
or UO_4742 (O_4742,N_49573,N_49183);
nand UO_4743 (O_4743,N_49125,N_49428);
xnor UO_4744 (O_4744,N_49331,N_49604);
xnor UO_4745 (O_4745,N_49631,N_49720);
and UO_4746 (O_4746,N_49510,N_49190);
and UO_4747 (O_4747,N_49620,N_49766);
or UO_4748 (O_4748,N_49668,N_49676);
or UO_4749 (O_4749,N_49992,N_49740);
nor UO_4750 (O_4750,N_49057,N_49504);
nand UO_4751 (O_4751,N_49995,N_49742);
and UO_4752 (O_4752,N_49539,N_49809);
nand UO_4753 (O_4753,N_49078,N_49226);
xor UO_4754 (O_4754,N_49178,N_49085);
and UO_4755 (O_4755,N_49784,N_49907);
nand UO_4756 (O_4756,N_49949,N_49367);
nand UO_4757 (O_4757,N_49097,N_49603);
or UO_4758 (O_4758,N_49198,N_49345);
xor UO_4759 (O_4759,N_49878,N_49155);
xnor UO_4760 (O_4760,N_49502,N_49935);
and UO_4761 (O_4761,N_49475,N_49564);
and UO_4762 (O_4762,N_49435,N_49670);
nand UO_4763 (O_4763,N_49284,N_49056);
or UO_4764 (O_4764,N_49417,N_49158);
nand UO_4765 (O_4765,N_49767,N_49193);
nand UO_4766 (O_4766,N_49037,N_49425);
nor UO_4767 (O_4767,N_49517,N_49532);
and UO_4768 (O_4768,N_49755,N_49569);
nand UO_4769 (O_4769,N_49046,N_49238);
xor UO_4770 (O_4770,N_49781,N_49184);
or UO_4771 (O_4771,N_49109,N_49783);
nor UO_4772 (O_4772,N_49145,N_49223);
xor UO_4773 (O_4773,N_49442,N_49380);
nand UO_4774 (O_4774,N_49845,N_49803);
xnor UO_4775 (O_4775,N_49680,N_49103);
or UO_4776 (O_4776,N_49173,N_49119);
and UO_4777 (O_4777,N_49104,N_49393);
xnor UO_4778 (O_4778,N_49764,N_49026);
or UO_4779 (O_4779,N_49557,N_49621);
or UO_4780 (O_4780,N_49053,N_49208);
or UO_4781 (O_4781,N_49125,N_49035);
xor UO_4782 (O_4782,N_49676,N_49892);
nand UO_4783 (O_4783,N_49502,N_49277);
xnor UO_4784 (O_4784,N_49980,N_49961);
nor UO_4785 (O_4785,N_49894,N_49224);
nand UO_4786 (O_4786,N_49523,N_49415);
nand UO_4787 (O_4787,N_49866,N_49624);
nor UO_4788 (O_4788,N_49505,N_49738);
or UO_4789 (O_4789,N_49639,N_49235);
and UO_4790 (O_4790,N_49249,N_49652);
xor UO_4791 (O_4791,N_49638,N_49276);
or UO_4792 (O_4792,N_49899,N_49419);
nor UO_4793 (O_4793,N_49593,N_49143);
and UO_4794 (O_4794,N_49175,N_49987);
nand UO_4795 (O_4795,N_49476,N_49729);
xor UO_4796 (O_4796,N_49160,N_49465);
xor UO_4797 (O_4797,N_49102,N_49834);
or UO_4798 (O_4798,N_49849,N_49372);
and UO_4799 (O_4799,N_49683,N_49093);
xnor UO_4800 (O_4800,N_49220,N_49283);
and UO_4801 (O_4801,N_49243,N_49948);
xor UO_4802 (O_4802,N_49358,N_49345);
nand UO_4803 (O_4803,N_49686,N_49886);
nor UO_4804 (O_4804,N_49137,N_49525);
nand UO_4805 (O_4805,N_49151,N_49391);
nand UO_4806 (O_4806,N_49951,N_49239);
nand UO_4807 (O_4807,N_49064,N_49372);
nor UO_4808 (O_4808,N_49391,N_49979);
or UO_4809 (O_4809,N_49040,N_49869);
or UO_4810 (O_4810,N_49684,N_49945);
and UO_4811 (O_4811,N_49728,N_49080);
nand UO_4812 (O_4812,N_49467,N_49217);
xnor UO_4813 (O_4813,N_49881,N_49824);
nor UO_4814 (O_4814,N_49277,N_49689);
or UO_4815 (O_4815,N_49062,N_49782);
nand UO_4816 (O_4816,N_49303,N_49021);
nand UO_4817 (O_4817,N_49184,N_49700);
and UO_4818 (O_4818,N_49153,N_49674);
and UO_4819 (O_4819,N_49307,N_49774);
or UO_4820 (O_4820,N_49996,N_49950);
and UO_4821 (O_4821,N_49163,N_49511);
and UO_4822 (O_4822,N_49929,N_49041);
or UO_4823 (O_4823,N_49315,N_49450);
nor UO_4824 (O_4824,N_49697,N_49101);
xnor UO_4825 (O_4825,N_49181,N_49844);
xnor UO_4826 (O_4826,N_49521,N_49335);
and UO_4827 (O_4827,N_49360,N_49870);
or UO_4828 (O_4828,N_49134,N_49895);
and UO_4829 (O_4829,N_49432,N_49807);
or UO_4830 (O_4830,N_49492,N_49420);
xnor UO_4831 (O_4831,N_49366,N_49408);
nand UO_4832 (O_4832,N_49428,N_49336);
or UO_4833 (O_4833,N_49536,N_49288);
nand UO_4834 (O_4834,N_49074,N_49963);
nor UO_4835 (O_4835,N_49830,N_49713);
xor UO_4836 (O_4836,N_49026,N_49076);
or UO_4837 (O_4837,N_49701,N_49458);
xnor UO_4838 (O_4838,N_49227,N_49681);
xnor UO_4839 (O_4839,N_49676,N_49624);
or UO_4840 (O_4840,N_49943,N_49993);
nor UO_4841 (O_4841,N_49807,N_49036);
and UO_4842 (O_4842,N_49644,N_49103);
nor UO_4843 (O_4843,N_49704,N_49241);
and UO_4844 (O_4844,N_49136,N_49684);
xnor UO_4845 (O_4845,N_49290,N_49873);
nand UO_4846 (O_4846,N_49256,N_49891);
xor UO_4847 (O_4847,N_49349,N_49461);
xor UO_4848 (O_4848,N_49825,N_49748);
xnor UO_4849 (O_4849,N_49875,N_49269);
nand UO_4850 (O_4850,N_49152,N_49298);
xnor UO_4851 (O_4851,N_49078,N_49465);
and UO_4852 (O_4852,N_49922,N_49902);
nor UO_4853 (O_4853,N_49686,N_49490);
nand UO_4854 (O_4854,N_49451,N_49173);
and UO_4855 (O_4855,N_49163,N_49461);
nand UO_4856 (O_4856,N_49563,N_49005);
xor UO_4857 (O_4857,N_49707,N_49979);
nand UO_4858 (O_4858,N_49774,N_49835);
or UO_4859 (O_4859,N_49645,N_49617);
xor UO_4860 (O_4860,N_49779,N_49144);
and UO_4861 (O_4861,N_49207,N_49460);
nand UO_4862 (O_4862,N_49789,N_49723);
and UO_4863 (O_4863,N_49426,N_49439);
or UO_4864 (O_4864,N_49129,N_49135);
nand UO_4865 (O_4865,N_49275,N_49281);
and UO_4866 (O_4866,N_49475,N_49087);
and UO_4867 (O_4867,N_49078,N_49267);
xnor UO_4868 (O_4868,N_49584,N_49813);
nor UO_4869 (O_4869,N_49251,N_49218);
nor UO_4870 (O_4870,N_49950,N_49943);
xor UO_4871 (O_4871,N_49097,N_49854);
xor UO_4872 (O_4872,N_49508,N_49556);
nand UO_4873 (O_4873,N_49353,N_49011);
xor UO_4874 (O_4874,N_49925,N_49428);
and UO_4875 (O_4875,N_49135,N_49987);
and UO_4876 (O_4876,N_49207,N_49696);
nand UO_4877 (O_4877,N_49008,N_49909);
nor UO_4878 (O_4878,N_49873,N_49758);
or UO_4879 (O_4879,N_49625,N_49583);
or UO_4880 (O_4880,N_49029,N_49441);
or UO_4881 (O_4881,N_49835,N_49530);
or UO_4882 (O_4882,N_49938,N_49211);
nor UO_4883 (O_4883,N_49312,N_49621);
nor UO_4884 (O_4884,N_49468,N_49993);
and UO_4885 (O_4885,N_49407,N_49046);
nand UO_4886 (O_4886,N_49112,N_49641);
nor UO_4887 (O_4887,N_49199,N_49888);
nor UO_4888 (O_4888,N_49259,N_49364);
and UO_4889 (O_4889,N_49271,N_49017);
nand UO_4890 (O_4890,N_49157,N_49514);
or UO_4891 (O_4891,N_49801,N_49190);
xnor UO_4892 (O_4892,N_49605,N_49451);
and UO_4893 (O_4893,N_49528,N_49464);
or UO_4894 (O_4894,N_49550,N_49883);
nor UO_4895 (O_4895,N_49176,N_49108);
and UO_4896 (O_4896,N_49244,N_49252);
xor UO_4897 (O_4897,N_49662,N_49968);
nor UO_4898 (O_4898,N_49343,N_49766);
and UO_4899 (O_4899,N_49173,N_49609);
and UO_4900 (O_4900,N_49634,N_49448);
nor UO_4901 (O_4901,N_49378,N_49454);
and UO_4902 (O_4902,N_49936,N_49733);
xnor UO_4903 (O_4903,N_49364,N_49870);
xnor UO_4904 (O_4904,N_49053,N_49566);
xor UO_4905 (O_4905,N_49920,N_49635);
and UO_4906 (O_4906,N_49437,N_49807);
nor UO_4907 (O_4907,N_49871,N_49567);
xor UO_4908 (O_4908,N_49713,N_49013);
or UO_4909 (O_4909,N_49975,N_49018);
and UO_4910 (O_4910,N_49373,N_49203);
or UO_4911 (O_4911,N_49790,N_49230);
and UO_4912 (O_4912,N_49895,N_49751);
nor UO_4913 (O_4913,N_49940,N_49231);
or UO_4914 (O_4914,N_49199,N_49749);
nand UO_4915 (O_4915,N_49635,N_49787);
nor UO_4916 (O_4916,N_49550,N_49152);
nor UO_4917 (O_4917,N_49444,N_49012);
or UO_4918 (O_4918,N_49523,N_49334);
nor UO_4919 (O_4919,N_49647,N_49611);
or UO_4920 (O_4920,N_49313,N_49357);
or UO_4921 (O_4921,N_49322,N_49109);
xor UO_4922 (O_4922,N_49101,N_49037);
xor UO_4923 (O_4923,N_49897,N_49597);
or UO_4924 (O_4924,N_49463,N_49039);
or UO_4925 (O_4925,N_49037,N_49415);
and UO_4926 (O_4926,N_49778,N_49542);
nor UO_4927 (O_4927,N_49456,N_49638);
nand UO_4928 (O_4928,N_49429,N_49349);
xnor UO_4929 (O_4929,N_49822,N_49969);
nand UO_4930 (O_4930,N_49815,N_49661);
or UO_4931 (O_4931,N_49820,N_49140);
xnor UO_4932 (O_4932,N_49165,N_49254);
xor UO_4933 (O_4933,N_49804,N_49212);
nand UO_4934 (O_4934,N_49391,N_49189);
or UO_4935 (O_4935,N_49803,N_49167);
or UO_4936 (O_4936,N_49192,N_49329);
nor UO_4937 (O_4937,N_49592,N_49260);
nor UO_4938 (O_4938,N_49597,N_49306);
or UO_4939 (O_4939,N_49701,N_49142);
nand UO_4940 (O_4940,N_49552,N_49958);
xnor UO_4941 (O_4941,N_49330,N_49402);
or UO_4942 (O_4942,N_49402,N_49199);
or UO_4943 (O_4943,N_49291,N_49849);
and UO_4944 (O_4944,N_49277,N_49011);
and UO_4945 (O_4945,N_49374,N_49621);
and UO_4946 (O_4946,N_49150,N_49599);
nand UO_4947 (O_4947,N_49597,N_49746);
xnor UO_4948 (O_4948,N_49981,N_49474);
and UO_4949 (O_4949,N_49728,N_49555);
xor UO_4950 (O_4950,N_49208,N_49864);
nor UO_4951 (O_4951,N_49545,N_49649);
and UO_4952 (O_4952,N_49242,N_49055);
nand UO_4953 (O_4953,N_49245,N_49273);
or UO_4954 (O_4954,N_49195,N_49437);
or UO_4955 (O_4955,N_49088,N_49594);
or UO_4956 (O_4956,N_49202,N_49194);
xnor UO_4957 (O_4957,N_49908,N_49756);
and UO_4958 (O_4958,N_49355,N_49613);
xnor UO_4959 (O_4959,N_49490,N_49383);
nand UO_4960 (O_4960,N_49827,N_49526);
or UO_4961 (O_4961,N_49509,N_49607);
nand UO_4962 (O_4962,N_49233,N_49406);
nor UO_4963 (O_4963,N_49967,N_49497);
and UO_4964 (O_4964,N_49136,N_49708);
nor UO_4965 (O_4965,N_49908,N_49897);
and UO_4966 (O_4966,N_49159,N_49541);
nor UO_4967 (O_4967,N_49148,N_49091);
or UO_4968 (O_4968,N_49176,N_49887);
and UO_4969 (O_4969,N_49624,N_49498);
nor UO_4970 (O_4970,N_49629,N_49439);
and UO_4971 (O_4971,N_49783,N_49898);
xnor UO_4972 (O_4972,N_49552,N_49356);
and UO_4973 (O_4973,N_49202,N_49325);
nor UO_4974 (O_4974,N_49155,N_49477);
and UO_4975 (O_4975,N_49588,N_49185);
nor UO_4976 (O_4976,N_49622,N_49136);
nand UO_4977 (O_4977,N_49008,N_49448);
or UO_4978 (O_4978,N_49041,N_49023);
nor UO_4979 (O_4979,N_49054,N_49778);
nor UO_4980 (O_4980,N_49400,N_49536);
and UO_4981 (O_4981,N_49834,N_49416);
xnor UO_4982 (O_4982,N_49379,N_49590);
nand UO_4983 (O_4983,N_49956,N_49025);
and UO_4984 (O_4984,N_49482,N_49367);
nand UO_4985 (O_4985,N_49035,N_49163);
nor UO_4986 (O_4986,N_49017,N_49043);
xnor UO_4987 (O_4987,N_49607,N_49766);
and UO_4988 (O_4988,N_49361,N_49270);
nand UO_4989 (O_4989,N_49523,N_49380);
nor UO_4990 (O_4990,N_49644,N_49253);
or UO_4991 (O_4991,N_49957,N_49084);
nor UO_4992 (O_4992,N_49055,N_49835);
nand UO_4993 (O_4993,N_49180,N_49364);
nor UO_4994 (O_4994,N_49338,N_49595);
xor UO_4995 (O_4995,N_49830,N_49136);
nand UO_4996 (O_4996,N_49084,N_49649);
nand UO_4997 (O_4997,N_49678,N_49767);
xor UO_4998 (O_4998,N_49174,N_49745);
and UO_4999 (O_4999,N_49462,N_49931);
endmodule