module basic_1500_15000_2000_10_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_845,In_101);
or U1 (N_1,In_751,In_205);
and U2 (N_2,In_283,In_1199);
and U3 (N_3,In_674,In_916);
and U4 (N_4,In_1408,In_1054);
and U5 (N_5,In_1205,In_970);
nand U6 (N_6,In_1089,In_601);
xnor U7 (N_7,In_943,In_321);
nand U8 (N_8,In_14,In_322);
xnor U9 (N_9,In_724,In_491);
or U10 (N_10,In_1092,In_841);
nand U11 (N_11,In_42,In_85);
nand U12 (N_12,In_1325,In_722);
xor U13 (N_13,In_1260,In_1178);
and U14 (N_14,In_887,In_1273);
nand U15 (N_15,In_1381,In_1167);
nor U16 (N_16,In_1316,In_22);
nor U17 (N_17,In_1341,In_740);
xnor U18 (N_18,In_1338,In_517);
nand U19 (N_19,In_363,In_796);
and U20 (N_20,In_410,In_655);
xor U21 (N_21,In_1490,In_12);
or U22 (N_22,In_155,In_1418);
and U23 (N_23,In_832,In_256);
nand U24 (N_24,In_1377,In_1051);
or U25 (N_25,In_1176,In_711);
xnor U26 (N_26,In_170,In_1286);
or U27 (N_27,In_1101,In_697);
xnor U28 (N_28,In_2,In_492);
and U29 (N_29,In_1188,In_825);
or U30 (N_30,In_501,In_1407);
and U31 (N_31,In_168,In_1467);
or U32 (N_32,In_1011,In_1242);
or U33 (N_33,In_1072,In_1264);
or U34 (N_34,In_1098,In_53);
nand U35 (N_35,In_1062,In_1077);
nand U36 (N_36,In_843,In_965);
and U37 (N_37,In_511,In_461);
and U38 (N_38,In_561,In_474);
or U39 (N_39,In_641,In_355);
or U40 (N_40,In_465,In_787);
and U41 (N_41,In_550,In_190);
nand U42 (N_42,In_922,In_166);
and U43 (N_43,In_254,In_948);
nand U44 (N_44,In_1268,In_135);
and U45 (N_45,In_804,In_1008);
or U46 (N_46,In_1061,In_177);
nor U47 (N_47,In_750,In_1030);
nand U48 (N_48,In_704,In_1454);
nor U49 (N_49,In_1102,In_273);
nand U50 (N_50,In_1150,In_1296);
xor U51 (N_51,In_701,In_624);
and U52 (N_52,In_638,In_1324);
and U53 (N_53,In_771,In_149);
or U54 (N_54,In_672,In_536);
or U55 (N_55,In_274,In_762);
and U56 (N_56,In_946,In_230);
and U57 (N_57,In_667,In_17);
and U58 (N_58,In_1481,In_1228);
nor U59 (N_59,In_164,In_147);
nor U60 (N_60,In_23,In_596);
nand U61 (N_61,In_666,In_829);
and U62 (N_62,In_241,In_1125);
nand U63 (N_63,In_107,In_1103);
nor U64 (N_64,In_1451,In_1184);
or U65 (N_65,In_1255,In_1015);
or U66 (N_66,In_124,In_1350);
and U67 (N_67,In_1081,In_897);
nand U68 (N_68,In_585,In_1269);
or U69 (N_69,In_734,In_1060);
and U70 (N_70,In_1311,In_702);
xor U71 (N_71,In_376,In_560);
or U72 (N_72,In_860,In_1174);
or U73 (N_73,In_982,In_86);
and U74 (N_74,In_464,In_478);
nor U75 (N_75,In_289,In_68);
or U76 (N_76,In_746,In_113);
and U77 (N_77,In_1074,In_1220);
and U78 (N_78,In_1497,In_873);
xnor U79 (N_79,In_633,In_1032);
and U80 (N_80,In_1148,In_422);
nor U81 (N_81,In_20,In_764);
nor U82 (N_82,In_47,In_304);
nand U83 (N_83,In_419,In_444);
or U84 (N_84,In_1227,In_800);
nand U85 (N_85,In_368,In_526);
nand U86 (N_86,In_104,In_1195);
nand U87 (N_87,In_330,In_1327);
nand U88 (N_88,In_0,In_815);
nand U89 (N_89,In_944,In_1342);
or U90 (N_90,In_1013,In_116);
nand U91 (N_91,In_665,In_670);
xor U92 (N_92,In_581,In_628);
nand U93 (N_93,In_936,In_502);
or U94 (N_94,In_1275,In_529);
nor U95 (N_95,In_906,In_1096);
and U96 (N_96,In_212,In_1486);
or U97 (N_97,In_699,In_677);
or U98 (N_98,In_950,In_1035);
nor U99 (N_99,In_1000,In_1285);
and U100 (N_100,In_275,In_772);
or U101 (N_101,In_980,In_1024);
nand U102 (N_102,In_807,In_1443);
nor U103 (N_103,In_853,In_455);
and U104 (N_104,In_436,In_611);
and U105 (N_105,In_221,In_657);
xnor U106 (N_106,In_610,In_1254);
nand U107 (N_107,In_1231,In_973);
nand U108 (N_108,In_213,In_1361);
nand U109 (N_109,In_954,In_1389);
xor U110 (N_110,In_442,In_453);
or U111 (N_111,In_1427,In_317);
and U112 (N_112,In_987,In_854);
xor U113 (N_113,In_938,In_584);
and U114 (N_114,In_1189,In_671);
or U115 (N_115,In_365,In_604);
nor U116 (N_116,In_857,In_579);
or U117 (N_117,In_310,In_700);
and U118 (N_118,In_341,In_1014);
nand U119 (N_119,In_1244,In_488);
and U120 (N_120,In_358,In_1320);
nand U121 (N_121,In_393,In_708);
xnor U122 (N_122,In_1073,In_281);
nand U123 (N_123,In_1403,In_1033);
nor U124 (N_124,In_544,In_174);
nand U125 (N_125,In_486,In_1290);
or U126 (N_126,In_542,In_430);
xnor U127 (N_127,In_114,In_319);
nand U128 (N_128,In_1281,In_730);
nor U129 (N_129,In_783,In_1139);
and U130 (N_130,In_400,In_1247);
nor U131 (N_131,In_731,In_882);
and U132 (N_132,In_588,In_423);
nand U133 (N_133,In_1163,In_139);
or U134 (N_134,In_745,In_695);
or U135 (N_135,In_1141,In_1357);
nor U136 (N_136,In_9,In_364);
nand U137 (N_137,In_569,In_131);
nand U138 (N_138,In_255,In_1134);
nand U139 (N_139,In_1160,In_271);
and U140 (N_140,In_901,In_990);
and U141 (N_141,In_564,In_1289);
and U142 (N_142,In_1238,In_1005);
or U143 (N_143,In_1235,In_1043);
nand U144 (N_144,In_237,In_1322);
and U145 (N_145,In_359,In_1469);
or U146 (N_146,In_1455,In_685);
nor U147 (N_147,In_573,In_661);
nor U148 (N_148,In_997,In_1293);
nor U149 (N_149,In_951,In_1373);
or U150 (N_150,In_1055,In_52);
nor U151 (N_151,In_328,In_975);
nor U152 (N_152,In_480,In_36);
nor U153 (N_153,In_1065,In_910);
nand U154 (N_154,In_490,In_947);
nor U155 (N_155,In_1262,In_597);
or U156 (N_156,In_599,In_425);
xor U157 (N_157,In_144,In_1007);
or U158 (N_158,In_1374,In_129);
nand U159 (N_159,In_810,In_818);
or U160 (N_160,In_1230,In_466);
nor U161 (N_161,In_993,In_758);
nor U162 (N_162,In_559,In_1474);
nor U163 (N_163,In_1113,In_713);
and U164 (N_164,In_1371,In_890);
xor U165 (N_165,In_774,In_379);
nand U166 (N_166,In_881,In_407);
and U167 (N_167,In_216,In_1162);
xor U168 (N_168,In_862,In_1378);
and U169 (N_169,In_875,In_755);
and U170 (N_170,In_1356,In_658);
nor U171 (N_171,In_138,In_361);
or U172 (N_172,In_928,In_1211);
and U173 (N_173,In_1217,In_505);
nand U174 (N_174,In_871,In_180);
and U175 (N_175,In_1223,In_345);
nor U176 (N_176,In_1093,In_75);
nor U177 (N_177,In_752,In_749);
nor U178 (N_178,In_1314,In_962);
nor U179 (N_179,In_662,In_1240);
nand U180 (N_180,In_1450,In_399);
xor U181 (N_181,In_272,In_90);
nand U182 (N_182,In_777,In_903);
or U183 (N_183,In_207,In_782);
nor U184 (N_184,In_864,In_248);
xnor U185 (N_185,In_959,In_1364);
xnor U186 (N_186,In_958,In_1456);
nand U187 (N_187,In_404,In_156);
or U188 (N_188,In_1334,In_316);
and U189 (N_189,In_1154,In_13);
and U190 (N_190,In_996,In_1222);
nand U191 (N_191,In_925,In_899);
and U192 (N_192,In_26,In_1473);
and U193 (N_193,In_1022,In_443);
and U194 (N_194,In_1018,In_117);
nand U195 (N_195,In_888,In_1442);
nor U196 (N_196,In_202,In_985);
or U197 (N_197,In_554,In_1441);
and U198 (N_198,In_32,In_199);
nor U199 (N_199,In_305,In_28);
or U200 (N_200,In_1124,In_1470);
nand U201 (N_201,In_504,In_314);
and U202 (N_202,In_214,In_1353);
nand U203 (N_203,In_1294,In_198);
nor U204 (N_204,In_719,In_522);
xor U205 (N_205,In_974,In_1464);
or U206 (N_206,In_932,In_720);
nand U207 (N_207,In_1336,In_495);
and U208 (N_208,In_1483,In_95);
nand U209 (N_209,In_176,In_1232);
xnor U210 (N_210,In_439,In_1012);
nor U211 (N_211,In_65,In_484);
or U212 (N_212,In_960,In_757);
or U213 (N_213,In_595,In_1498);
xor U214 (N_214,In_684,In_1169);
nor U215 (N_215,In_88,In_433);
or U216 (N_216,In_318,In_836);
and U217 (N_217,In_150,In_1375);
nand U218 (N_218,In_300,In_868);
nand U219 (N_219,In_767,In_420);
nor U220 (N_220,In_1354,In_8);
nor U221 (N_221,In_1419,In_1224);
or U222 (N_222,In_130,In_243);
nor U223 (N_223,In_528,In_696);
nand U224 (N_224,In_1291,In_983);
nor U225 (N_225,In_1395,In_683);
and U226 (N_226,In_1433,In_776);
nor U227 (N_227,In_952,In_127);
and U228 (N_228,In_942,In_1376);
nor U229 (N_229,In_162,In_178);
nand U230 (N_230,In_929,In_1239);
and U231 (N_231,In_386,In_335);
nand U232 (N_232,In_1006,In_1145);
nand U233 (N_233,In_703,In_840);
nand U234 (N_234,In_1352,In_848);
and U235 (N_235,In_440,In_1121);
and U236 (N_236,In_1380,In_593);
xnor U237 (N_237,In_828,In_1057);
or U238 (N_238,In_877,In_209);
xnor U239 (N_239,In_1059,In_842);
nor U240 (N_240,In_521,In_540);
xor U241 (N_241,In_1406,In_1432);
nand U242 (N_242,In_591,In_1144);
nor U243 (N_243,In_642,In_592);
nand U244 (N_244,In_1156,In_885);
nand U245 (N_245,In_817,In_999);
and U246 (N_246,In_1094,In_370);
and U247 (N_247,In_1095,In_191);
nor U248 (N_248,In_298,In_351);
nand U249 (N_249,In_1248,In_353);
or U250 (N_250,In_19,In_1108);
nand U251 (N_251,In_506,In_184);
nand U252 (N_252,In_986,In_1187);
or U253 (N_253,In_535,In_570);
and U254 (N_254,In_1204,In_51);
nand U255 (N_255,In_100,In_756);
nor U256 (N_256,In_367,In_238);
and U257 (N_257,In_435,In_1137);
and U258 (N_258,In_438,In_193);
xor U259 (N_259,In_1344,In_531);
nor U260 (N_260,In_781,In_1253);
xor U261 (N_261,In_913,In_228);
and U262 (N_262,In_813,In_543);
or U263 (N_263,In_240,In_729);
and U264 (N_264,In_1112,In_390);
nor U265 (N_265,In_659,In_481);
nand U266 (N_266,In_879,In_968);
and U267 (N_267,In_904,In_1114);
xor U268 (N_268,In_1328,In_1409);
or U269 (N_269,In_768,In_1368);
and U270 (N_270,In_615,In_878);
nor U271 (N_271,In_737,In_148);
nor U272 (N_272,In_1164,In_1360);
xor U273 (N_273,In_1277,In_1460);
xnor U274 (N_274,In_57,In_1129);
xor U275 (N_275,In_99,In_1272);
nand U276 (N_276,In_1123,In_1111);
and U277 (N_277,In_1346,In_1476);
or U278 (N_278,In_446,In_865);
nor U279 (N_279,In_354,In_134);
or U280 (N_280,In_485,In_77);
and U281 (N_281,In_1106,In_891);
nand U282 (N_282,In_1050,In_1090);
or U283 (N_283,In_552,In_995);
nor U284 (N_284,In_11,In_680);
and U285 (N_285,In_374,In_87);
xnor U286 (N_286,In_1430,In_861);
or U287 (N_287,In_1313,In_1391);
nor U288 (N_288,In_824,In_471);
xor U289 (N_289,In_892,In_627);
xor U290 (N_290,In_1034,In_1405);
xnor U291 (N_291,In_1383,In_1207);
or U292 (N_292,In_636,In_80);
or U293 (N_293,In_197,In_1063);
or U294 (N_294,In_1142,In_372);
or U295 (N_295,In_826,In_664);
and U296 (N_296,In_833,In_132);
and U297 (N_297,In_647,In_1166);
nand U298 (N_298,In_172,In_921);
xnor U299 (N_299,In_1362,In_1122);
or U300 (N_300,In_143,In_278);
or U301 (N_301,In_447,In_126);
nand U302 (N_302,In_336,In_189);
or U303 (N_303,In_524,In_1412);
and U304 (N_304,In_673,In_565);
nor U305 (N_305,In_280,In_409);
nand U306 (N_306,In_1306,In_509);
nor U307 (N_307,In_1039,In_1143);
nor U308 (N_308,In_378,In_525);
nand U309 (N_309,In_362,In_1283);
xnor U310 (N_310,In_902,In_911);
or U311 (N_311,In_739,In_277);
or U312 (N_312,In_500,In_935);
nor U313 (N_313,In_270,In_21);
nand U314 (N_314,In_219,In_792);
and U315 (N_315,In_1267,In_1318);
nand U316 (N_316,In_726,In_1126);
nand U317 (N_317,In_431,In_369);
nand U318 (N_318,In_94,In_852);
xor U319 (N_319,In_1351,In_794);
and U320 (N_320,In_58,In_1028);
nand U321 (N_321,In_4,In_246);
nand U322 (N_322,In_991,In_681);
nor U323 (N_323,In_69,In_508);
nor U324 (N_324,In_618,In_884);
or U325 (N_325,In_360,In_515);
xor U326 (N_326,In_231,In_1308);
nor U327 (N_327,In_1333,In_898);
or U328 (N_328,In_242,In_1069);
xnor U329 (N_329,In_1251,In_859);
or U330 (N_330,In_778,In_606);
and U331 (N_331,In_686,In_953);
and U332 (N_332,In_476,In_646);
nor U333 (N_333,In_1100,In_1127);
nand U334 (N_334,In_333,In_118);
nand U335 (N_335,In_741,In_121);
nor U336 (N_336,In_806,In_366);
nor U337 (N_337,In_437,In_1196);
or U338 (N_338,In_1263,In_1031);
or U339 (N_339,In_309,In_1170);
and U340 (N_340,In_837,In_346);
nor U341 (N_341,In_926,In_924);
and U342 (N_342,In_1171,In_161);
or U343 (N_343,In_556,In_918);
and U344 (N_344,In_1044,In_1250);
nand U345 (N_345,In_217,In_153);
and U346 (N_346,In_115,In_1146);
nand U347 (N_347,In_1379,In_222);
nor U348 (N_348,In_223,In_110);
nor U349 (N_349,In_1394,In_252);
nand U350 (N_350,In_1386,In_1261);
nand U351 (N_351,In_1052,In_1117);
nand U352 (N_352,In_41,In_226);
or U353 (N_353,In_1457,In_1023);
and U354 (N_354,In_1038,In_1440);
and U355 (N_355,In_608,In_454);
and U356 (N_356,In_414,In_1482);
and U357 (N_357,In_429,In_640);
nand U358 (N_358,In_1449,In_558);
nand U359 (N_359,In_1084,In_1119);
xor U360 (N_360,In_1215,In_1465);
nor U361 (N_361,In_574,In_1493);
and U362 (N_362,In_417,In_306);
and U363 (N_363,In_621,In_1434);
and U364 (N_364,In_1203,In_770);
and U365 (N_365,In_1168,In_449);
and U366 (N_366,In_1002,In_937);
and U367 (N_367,In_623,In_265);
nand U368 (N_368,In_766,In_743);
or U369 (N_369,In_603,In_1128);
or U370 (N_370,In_102,In_203);
nor U371 (N_371,In_562,In_1274);
nand U372 (N_372,In_1249,In_1037);
xor U373 (N_373,In_523,In_40);
nand U374 (N_374,In_571,In_337);
nand U375 (N_375,In_555,In_786);
nor U376 (N_376,In_392,In_652);
xor U377 (N_377,In_285,In_470);
or U378 (N_378,In_356,In_1214);
nor U379 (N_379,In_577,In_247);
nand U380 (N_380,In_250,In_208);
nor U381 (N_381,In_769,In_387);
or U382 (N_382,In_183,In_789);
and U383 (N_383,In_1071,In_917);
or U384 (N_384,In_259,In_1105);
or U385 (N_385,In_589,In_1151);
nand U386 (N_386,In_1216,In_1179);
nor U387 (N_387,In_450,In_1067);
or U388 (N_388,In_537,In_1083);
or U389 (N_389,In_1452,In_590);
and U390 (N_390,In_1218,In_855);
or U391 (N_391,In_1367,In_428);
nand U392 (N_392,In_204,In_1206);
nor U393 (N_393,In_512,In_1234);
nor U394 (N_394,In_644,In_181);
xnor U395 (N_395,In_693,In_736);
nand U396 (N_396,In_55,In_1444);
nand U397 (N_397,In_691,In_269);
nand U398 (N_398,In_1495,In_790);
xnor U399 (N_399,In_263,In_759);
or U400 (N_400,In_320,In_1068);
or U401 (N_401,In_1003,In_715);
or U402 (N_402,In_296,In_206);
and U403 (N_403,In_656,In_342);
nor U404 (N_404,In_89,In_883);
and U405 (N_405,In_1424,In_1209);
and U406 (N_406,In_940,In_227);
or U407 (N_407,In_451,In_1225);
or U408 (N_408,In_78,In_234);
and U409 (N_409,In_1001,In_1278);
and U410 (N_410,In_424,In_192);
and U411 (N_411,In_344,In_738);
nor U412 (N_412,In_448,In_748);
and U413 (N_413,In_432,In_1107);
or U414 (N_414,In_557,In_1130);
nand U415 (N_415,In_1027,In_1410);
nor U416 (N_416,In_613,In_347);
and U417 (N_417,In_137,In_457);
and U418 (N_418,In_251,In_302);
nor U419 (N_419,In_617,In_827);
or U420 (N_420,In_846,In_648);
nor U421 (N_421,In_175,In_744);
nand U422 (N_422,In_1036,In_1431);
nor U423 (N_423,In_635,In_201);
nor U424 (N_424,In_1042,In_520);
xor U425 (N_425,In_598,In_1202);
and U426 (N_426,In_1016,In_1393);
xnor U427 (N_427,In_1288,In_1229);
and U428 (N_428,In_539,In_63);
or U429 (N_429,In_1080,In_496);
and U430 (N_430,In_714,In_258);
and U431 (N_431,In_629,In_1305);
xnor U432 (N_432,In_1366,In_548);
and U433 (N_433,In_572,In_1226);
nand U434 (N_434,In_25,In_896);
and U435 (N_435,In_1348,In_1133);
xor U436 (N_436,In_185,In_717);
and U437 (N_437,In_357,In_972);
and U438 (N_438,In_377,In_709);
and U439 (N_439,In_1411,In_1303);
nand U440 (N_440,In_286,In_587);
and U441 (N_441,In_1335,In_620);
nand U442 (N_442,In_866,In_388);
xnor U443 (N_443,In_669,In_1301);
and U444 (N_444,In_239,In_1319);
nand U445 (N_445,In_384,In_473);
or U446 (N_446,In_907,In_880);
and U447 (N_447,In_1088,In_489);
and U448 (N_448,In_513,In_1287);
nor U449 (N_449,In_1329,In_1485);
xor U450 (N_450,In_1448,In_299);
nor U451 (N_451,In_630,In_1401);
nand U452 (N_452,In_1414,In_634);
or U453 (N_453,In_742,In_602);
nand U454 (N_454,In_914,In_1173);
nor U455 (N_455,In_992,In_452);
or U456 (N_456,In_293,In_775);
or U457 (N_457,In_716,In_1310);
nand U458 (N_458,In_867,In_1259);
nor U459 (N_459,In_1172,In_1459);
or U460 (N_460,In_838,In_1326);
or U461 (N_461,In_1079,In_260);
and U462 (N_462,In_288,In_67);
nor U463 (N_463,In_325,In_1292);
nand U464 (N_464,In_735,In_195);
or U465 (N_465,In_1307,In_3);
nor U466 (N_466,In_39,In_1026);
nor U467 (N_467,In_773,In_939);
nor U468 (N_468,In_851,In_732);
nand U469 (N_469,In_1478,In_38);
nor U470 (N_470,In_1331,In_956);
and U471 (N_471,In_233,In_83);
nor U472 (N_472,In_1445,In_1140);
and U473 (N_473,In_728,In_1104);
or U474 (N_474,In_619,In_1309);
nand U475 (N_475,In_805,In_791);
nand U476 (N_476,In_519,In_292);
nand U477 (N_477,In_923,In_1347);
nand U478 (N_478,In_1369,In_35);
nor U479 (N_479,In_1219,In_169);
or U480 (N_480,In_313,In_103);
or U481 (N_481,In_567,In_931);
nand U482 (N_482,In_327,In_1477);
or U483 (N_483,In_160,In_1298);
and U484 (N_484,In_1058,In_1177);
or U485 (N_485,In_1256,In_403);
nor U486 (N_486,In_1020,In_1082);
nor U487 (N_487,In_1049,In_847);
or U488 (N_488,In_499,In_839);
or U489 (N_489,In_1438,In_266);
nand U490 (N_490,In_282,In_1479);
nand U491 (N_491,In_799,In_1384);
nor U492 (N_492,In_1337,In_1019);
and U493 (N_493,In_663,In_725);
nand U494 (N_494,In_232,In_831);
nand U495 (N_495,In_1468,In_173);
and U496 (N_496,In_1025,In_721);
nor U497 (N_497,In_385,In_609);
and U498 (N_498,In_1382,In_236);
nor U499 (N_499,In_582,In_830);
nand U500 (N_500,In_889,In_1197);
or U501 (N_501,In_733,In_1241);
nand U502 (N_502,In_919,In_1372);
and U503 (N_503,In_532,In_622);
nor U504 (N_504,In_514,In_811);
nor U505 (N_505,In_391,In_727);
and U506 (N_506,In_1021,In_812);
nor U507 (N_507,In_760,In_1066);
nor U508 (N_508,In_1439,In_1257);
or U509 (N_509,In_445,In_583);
and U510 (N_510,In_820,In_163);
and U511 (N_511,In_76,In_224);
or U512 (N_512,In_780,In_91);
nor U513 (N_513,In_381,In_245);
or U514 (N_514,In_326,In_1200);
or U515 (N_515,In_1297,In_262);
or U516 (N_516,In_415,In_527);
nor U517 (N_517,In_93,In_600);
nor U518 (N_518,In_182,In_1265);
nor U519 (N_519,In_1402,In_546);
and U520 (N_520,In_1115,In_905);
or U521 (N_521,In_1365,In_1110);
or U522 (N_522,In_334,In_754);
or U523 (N_523,In_566,In_1208);
or U524 (N_524,In_984,In_692);
or U525 (N_525,In_798,In_1157);
nand U526 (N_526,In_1118,In_405);
and U527 (N_527,In_1400,In_493);
nand U528 (N_528,In_1416,In_689);
nor U529 (N_529,In_941,In_73);
and U530 (N_530,In_331,In_507);
or U531 (N_531,In_105,In_784);
and U532 (N_532,In_1388,In_510);
nor U533 (N_533,In_1009,In_268);
or U534 (N_534,In_1475,In_397);
nand U535 (N_535,In_1461,In_1396);
nor U536 (N_536,In_1420,In_1284);
or U537 (N_537,In_1472,In_797);
or U538 (N_538,In_61,In_834);
xnor U539 (N_539,In_1191,In_1153);
xnor U540 (N_540,In_7,In_50);
xor U541 (N_541,In_261,In_553);
and U542 (N_542,In_1161,In_912);
and U543 (N_543,In_339,In_1138);
or U544 (N_544,In_123,In_303);
and U545 (N_545,In_421,In_284);
nand U546 (N_546,In_688,In_441);
and U547 (N_547,In_779,In_159);
and U548 (N_548,In_1423,In_534);
nor U549 (N_549,In_1422,In_1245);
and U550 (N_550,In_412,In_1149);
nor U551 (N_551,In_1355,In_1132);
and U552 (N_552,In_1295,In_332);
nor U553 (N_553,In_1330,In_886);
nand U554 (N_554,In_1212,In_133);
nand U555 (N_555,In_1471,In_795);
nor U556 (N_556,In_1004,In_253);
nand U557 (N_557,In_338,In_352);
xnor U558 (N_558,In_971,In_1120);
nand U559 (N_559,In_62,In_413);
xor U560 (N_560,In_1466,In_895);
nand U561 (N_561,In_348,In_687);
and U562 (N_562,In_698,In_1417);
or U563 (N_563,In_235,In_967);
or U564 (N_564,In_477,In_34);
nand U565 (N_565,In_1053,In_70);
or U566 (N_566,In_434,In_276);
and U567 (N_567,In_6,In_312);
nand U568 (N_568,In_395,In_1017);
nand U569 (N_569,In_981,In_616);
and U570 (N_570,In_291,In_1155);
nand U571 (N_571,In_1210,In_761);
and U572 (N_572,In_1458,In_1064);
nor U573 (N_573,In_1186,In_60);
and U574 (N_574,In_1040,In_1421);
and U575 (N_575,In_545,In_125);
xnor U576 (N_576,In_1087,In_66);
or U577 (N_577,In_158,In_1300);
and U578 (N_578,In_1463,In_483);
nand U579 (N_579,In_863,In_1415);
or U580 (N_580,In_533,In_653);
xor U581 (N_581,In_1192,In_297);
nand U582 (N_582,In_290,In_1091);
nand U583 (N_583,In_72,In_179);
and U584 (N_584,In_632,In_349);
xor U585 (N_585,In_1413,In_79);
and U586 (N_586,In_30,In_816);
xor U587 (N_587,In_1302,In_1499);
xnor U588 (N_588,In_614,In_814);
nand U589 (N_589,In_1029,In_92);
and U590 (N_590,In_154,In_858);
nor U591 (N_591,In_876,In_998);
and U592 (N_592,In_1135,In_530);
or U593 (N_593,In_955,In_1236);
or U594 (N_594,In_712,In_822);
nand U595 (N_595,In_870,In_37);
and U596 (N_596,In_1246,In_1494);
or U597 (N_597,In_97,In_16);
and U598 (N_598,In_690,In_401);
or U599 (N_599,In_1099,In_463);
nor U600 (N_600,In_612,In_74);
and U601 (N_601,In_1279,In_1116);
xnor U602 (N_602,In_1086,In_675);
nand U603 (N_603,In_989,In_1252);
nand U604 (N_604,In_109,In_626);
and U605 (N_605,In_287,In_607);
nand U606 (N_606,In_340,In_398);
nand U607 (N_607,In_1056,In_1390);
xnor U608 (N_608,In_1,In_1243);
nand U609 (N_609,In_343,In_497);
or U610 (N_610,In_1221,In_111);
or U611 (N_611,In_396,In_563);
nand U612 (N_612,In_5,In_1304);
and U613 (N_613,In_56,In_188);
xor U614 (N_614,In_1385,In_1194);
or U615 (N_615,In_225,In_788);
or U616 (N_616,In_141,In_978);
or U617 (N_617,In_893,In_1258);
nand U618 (N_618,In_1201,In_1048);
nor U619 (N_619,In_718,In_1462);
nor U620 (N_620,In_994,In_963);
nand U621 (N_621,In_152,In_1147);
or U622 (N_622,In_1312,In_650);
nand U623 (N_623,In_1339,In_1436);
and U624 (N_624,In_29,In_707);
nand U625 (N_625,In_1387,In_538);
nor U626 (N_626,In_145,In_1392);
nand U627 (N_627,In_1198,In_835);
nand U628 (N_628,In_668,In_908);
or U629 (N_629,In_605,In_187);
nand U630 (N_630,In_1041,In_324);
nand U631 (N_631,In_964,In_1398);
and U632 (N_632,In_1321,In_945);
and U633 (N_633,In_1276,In_1271);
and U634 (N_634,In_171,In_122);
nor U635 (N_635,In_10,In_1447);
or U636 (N_636,In_1317,In_518);
nor U637 (N_637,In_301,In_631);
nor U638 (N_638,In_1270,In_244);
or U639 (N_639,In_1190,In_988);
nor U640 (N_640,In_165,In_637);
and U641 (N_641,In_64,In_679);
nor U642 (N_642,In_541,In_45);
nor U643 (N_643,In_900,In_753);
and U644 (N_644,In_112,In_874);
nand U645 (N_645,In_311,In_462);
and U646 (N_646,In_763,In_1488);
or U647 (N_647,In_1045,In_819);
or U648 (N_648,In_869,In_406);
nor U649 (N_649,In_568,In_1359);
and U650 (N_650,In_1185,In_18);
nand U651 (N_651,In_1399,In_682);
nand U652 (N_652,In_142,In_383);
and U653 (N_653,In_157,In_1489);
and U654 (N_654,In_594,In_1349);
xnor U655 (N_655,In_249,In_257);
and U656 (N_656,In_27,In_427);
and U657 (N_657,In_1159,In_308);
and U658 (N_658,In_1180,In_1446);
and U659 (N_659,In_850,In_549);
nand U660 (N_660,In_196,In_1193);
or U661 (N_661,In_31,In_894);
nor U662 (N_662,In_872,In_458);
or U663 (N_663,In_1437,In_654);
or U664 (N_664,In_1315,In_676);
nor U665 (N_665,In_933,In_1131);
nand U666 (N_666,In_801,In_949);
nor U667 (N_667,In_1097,In_81);
xor U668 (N_668,In_71,In_1492);
nand U669 (N_669,In_279,In_15);
nand U670 (N_670,In_639,In_108);
and U671 (N_671,In_747,In_979);
and U672 (N_672,In_1183,In_625);
nor U673 (N_673,In_660,In_380);
or U674 (N_674,In_1175,In_849);
and U675 (N_675,In_803,In_1404);
and U676 (N_676,In_785,In_844);
or U677 (N_677,In_649,In_48);
nand U678 (N_678,In_809,In_586);
nand U679 (N_679,In_1340,In_1046);
nand U680 (N_680,In_140,In_146);
nand U681 (N_681,In_373,In_1233);
or U682 (N_682,In_1010,In_264);
nand U683 (N_683,In_371,In_961);
nor U684 (N_684,In_389,In_1237);
and U685 (N_685,In_220,In_823);
nand U686 (N_686,In_482,In_516);
nand U687 (N_687,In_210,In_307);
or U688 (N_688,In_408,In_678);
or U689 (N_689,In_551,In_969);
xor U690 (N_690,In_167,In_96);
nor U691 (N_691,In_1429,In_793);
and U692 (N_692,In_416,In_1182);
and U693 (N_693,In_200,In_418);
nand U694 (N_694,In_186,In_1453);
nand U695 (N_695,In_580,In_706);
or U696 (N_696,In_645,In_498);
nand U697 (N_697,In_1213,In_43);
nor U698 (N_698,In_1491,In_44);
or U699 (N_699,In_426,In_487);
xnor U700 (N_700,In_375,In_1078);
nor U701 (N_701,In_1299,In_1484);
and U702 (N_702,In_411,In_494);
nand U703 (N_703,In_315,In_211);
and U704 (N_704,In_84,In_1282);
and U705 (N_705,In_976,In_1435);
or U706 (N_706,In_1047,In_1266);
xor U707 (N_707,In_1343,In_267);
xnor U708 (N_708,In_930,In_475);
and U709 (N_709,In_120,In_1345);
nand U710 (N_710,In_1152,In_468);
nand U711 (N_711,In_977,In_295);
or U712 (N_712,In_765,In_1181);
nand U713 (N_713,In_350,In_909);
nand U714 (N_714,In_1075,In_1480);
and U715 (N_715,In_1332,In_1136);
and U716 (N_716,In_920,In_54);
nor U717 (N_717,In_469,In_576);
nand U718 (N_718,In_467,In_503);
xor U719 (N_719,In_1165,In_651);
and U720 (N_720,In_119,In_460);
xor U721 (N_721,In_1323,In_1397);
nand U722 (N_722,In_1085,In_456);
or U723 (N_723,In_479,In_821);
nor U724 (N_724,In_46,In_705);
and U725 (N_725,In_323,In_802);
nand U726 (N_726,In_1070,In_723);
and U727 (N_727,In_229,In_1426);
and U728 (N_728,In_1358,In_1280);
nand U729 (N_729,In_151,In_472);
or U730 (N_730,In_329,In_59);
and U731 (N_731,In_215,In_402);
nand U732 (N_732,In_98,In_1425);
and U733 (N_733,In_856,In_49);
or U734 (N_734,In_694,In_106);
nand U735 (N_735,In_1428,In_294);
and U736 (N_736,In_1370,In_33);
nand U737 (N_737,In_394,In_934);
xor U738 (N_738,In_194,In_1076);
or U739 (N_739,In_927,In_1487);
nor U740 (N_740,In_575,In_643);
or U741 (N_741,In_915,In_1158);
nand U742 (N_742,In_957,In_1363);
or U743 (N_743,In_382,In_1109);
or U744 (N_744,In_128,In_1496);
nand U745 (N_745,In_578,In_710);
nor U746 (N_746,In_82,In_24);
or U747 (N_747,In_966,In_547);
nor U748 (N_748,In_136,In_808);
nand U749 (N_749,In_459,In_218);
nor U750 (N_750,In_1196,In_926);
nor U751 (N_751,In_18,In_1158);
and U752 (N_752,In_298,In_486);
and U753 (N_753,In_424,In_561);
nand U754 (N_754,In_1386,In_493);
nand U755 (N_755,In_1197,In_553);
or U756 (N_756,In_158,In_745);
or U757 (N_757,In_1179,In_1359);
nor U758 (N_758,In_86,In_1442);
nand U759 (N_759,In_1315,In_1150);
xor U760 (N_760,In_1024,In_1490);
xor U761 (N_761,In_352,In_1372);
nor U762 (N_762,In_408,In_810);
and U763 (N_763,In_336,In_360);
nand U764 (N_764,In_130,In_1314);
or U765 (N_765,In_290,In_506);
or U766 (N_766,In_1360,In_1175);
nor U767 (N_767,In_200,In_465);
and U768 (N_768,In_576,In_143);
nor U769 (N_769,In_203,In_210);
nand U770 (N_770,In_229,In_1197);
or U771 (N_771,In_578,In_896);
nor U772 (N_772,In_467,In_202);
or U773 (N_773,In_1270,In_826);
nand U774 (N_774,In_343,In_1274);
nor U775 (N_775,In_183,In_660);
nor U776 (N_776,In_952,In_683);
nor U777 (N_777,In_670,In_1216);
or U778 (N_778,In_1054,In_550);
nand U779 (N_779,In_809,In_332);
nand U780 (N_780,In_1257,In_317);
and U781 (N_781,In_1388,In_511);
xnor U782 (N_782,In_470,In_1119);
and U783 (N_783,In_1394,In_142);
or U784 (N_784,In_1496,In_1346);
nor U785 (N_785,In_522,In_1041);
and U786 (N_786,In_236,In_1443);
nand U787 (N_787,In_1260,In_1189);
or U788 (N_788,In_167,In_356);
or U789 (N_789,In_836,In_46);
and U790 (N_790,In_568,In_390);
and U791 (N_791,In_1115,In_1146);
nor U792 (N_792,In_898,In_1139);
xnor U793 (N_793,In_872,In_276);
xor U794 (N_794,In_1436,In_1330);
xnor U795 (N_795,In_562,In_235);
nand U796 (N_796,In_796,In_681);
or U797 (N_797,In_770,In_474);
nor U798 (N_798,In_219,In_269);
and U799 (N_799,In_1355,In_301);
nor U800 (N_800,In_1205,In_927);
or U801 (N_801,In_28,In_1159);
or U802 (N_802,In_1347,In_228);
or U803 (N_803,In_687,In_67);
or U804 (N_804,In_719,In_1436);
nor U805 (N_805,In_1095,In_1306);
or U806 (N_806,In_969,In_984);
and U807 (N_807,In_532,In_1236);
nand U808 (N_808,In_637,In_50);
or U809 (N_809,In_932,In_182);
nor U810 (N_810,In_1235,In_959);
nor U811 (N_811,In_415,In_833);
and U812 (N_812,In_915,In_212);
nand U813 (N_813,In_113,In_149);
or U814 (N_814,In_1437,In_1248);
xnor U815 (N_815,In_1396,In_1034);
or U816 (N_816,In_314,In_1395);
nor U817 (N_817,In_1300,In_961);
and U818 (N_818,In_931,In_1302);
or U819 (N_819,In_136,In_1229);
xor U820 (N_820,In_1171,In_335);
or U821 (N_821,In_180,In_1190);
and U822 (N_822,In_1301,In_1220);
xnor U823 (N_823,In_896,In_347);
or U824 (N_824,In_980,In_433);
or U825 (N_825,In_12,In_1118);
nand U826 (N_826,In_413,In_244);
nor U827 (N_827,In_831,In_939);
and U828 (N_828,In_1077,In_451);
or U829 (N_829,In_978,In_1240);
or U830 (N_830,In_608,In_1334);
and U831 (N_831,In_19,In_565);
or U832 (N_832,In_699,In_393);
nor U833 (N_833,In_235,In_1372);
xnor U834 (N_834,In_445,In_1155);
nand U835 (N_835,In_881,In_601);
or U836 (N_836,In_1017,In_581);
nand U837 (N_837,In_1055,In_1253);
or U838 (N_838,In_995,In_1200);
and U839 (N_839,In_18,In_356);
xor U840 (N_840,In_129,In_32);
and U841 (N_841,In_626,In_445);
nand U842 (N_842,In_140,In_403);
nor U843 (N_843,In_1245,In_261);
and U844 (N_844,In_1119,In_218);
or U845 (N_845,In_1067,In_758);
nor U846 (N_846,In_705,In_789);
and U847 (N_847,In_687,In_1295);
nand U848 (N_848,In_1197,In_109);
xnor U849 (N_849,In_72,In_396);
nor U850 (N_850,In_1279,In_1355);
and U851 (N_851,In_100,In_614);
xnor U852 (N_852,In_513,In_337);
nand U853 (N_853,In_1389,In_908);
nand U854 (N_854,In_664,In_1321);
nand U855 (N_855,In_229,In_1190);
and U856 (N_856,In_1274,In_330);
and U857 (N_857,In_109,In_906);
or U858 (N_858,In_796,In_1328);
and U859 (N_859,In_1065,In_1323);
or U860 (N_860,In_546,In_62);
nand U861 (N_861,In_477,In_1191);
nand U862 (N_862,In_1448,In_230);
nand U863 (N_863,In_704,In_1174);
or U864 (N_864,In_795,In_828);
nand U865 (N_865,In_778,In_677);
nor U866 (N_866,In_879,In_334);
nor U867 (N_867,In_1030,In_1488);
nor U868 (N_868,In_910,In_709);
nor U869 (N_869,In_158,In_1221);
or U870 (N_870,In_420,In_522);
nor U871 (N_871,In_296,In_438);
nand U872 (N_872,In_570,In_1320);
or U873 (N_873,In_526,In_1430);
or U874 (N_874,In_1399,In_1018);
and U875 (N_875,In_443,In_879);
nand U876 (N_876,In_833,In_1000);
nor U877 (N_877,In_1444,In_422);
nand U878 (N_878,In_1426,In_526);
or U879 (N_879,In_1266,In_29);
and U880 (N_880,In_568,In_1200);
or U881 (N_881,In_1112,In_416);
or U882 (N_882,In_268,In_390);
or U883 (N_883,In_1356,In_467);
nor U884 (N_884,In_1072,In_564);
nand U885 (N_885,In_1113,In_1271);
and U886 (N_886,In_1199,In_1003);
and U887 (N_887,In_537,In_1402);
and U888 (N_888,In_698,In_1452);
nand U889 (N_889,In_1106,In_327);
nor U890 (N_890,In_23,In_307);
nor U891 (N_891,In_576,In_768);
nor U892 (N_892,In_605,In_877);
nand U893 (N_893,In_807,In_783);
nor U894 (N_894,In_1448,In_986);
nand U895 (N_895,In_1376,In_952);
and U896 (N_896,In_235,In_1259);
or U897 (N_897,In_122,In_1465);
or U898 (N_898,In_144,In_306);
or U899 (N_899,In_229,In_673);
nor U900 (N_900,In_501,In_1307);
nor U901 (N_901,In_25,In_1059);
or U902 (N_902,In_139,In_1462);
and U903 (N_903,In_1156,In_281);
xnor U904 (N_904,In_1051,In_1358);
nand U905 (N_905,In_660,In_300);
nand U906 (N_906,In_1303,In_858);
nand U907 (N_907,In_378,In_765);
or U908 (N_908,In_618,In_1131);
and U909 (N_909,In_902,In_723);
xnor U910 (N_910,In_1005,In_515);
xnor U911 (N_911,In_585,In_159);
or U912 (N_912,In_1138,In_959);
and U913 (N_913,In_399,In_183);
and U914 (N_914,In_1461,In_1129);
and U915 (N_915,In_402,In_1347);
or U916 (N_916,In_606,In_590);
or U917 (N_917,In_316,In_123);
xor U918 (N_918,In_38,In_784);
nand U919 (N_919,In_70,In_1411);
nand U920 (N_920,In_91,In_5);
nand U921 (N_921,In_889,In_4);
or U922 (N_922,In_1263,In_1128);
and U923 (N_923,In_252,In_1180);
and U924 (N_924,In_1104,In_1422);
nand U925 (N_925,In_1066,In_1316);
and U926 (N_926,In_964,In_1422);
nand U927 (N_927,In_1348,In_1019);
or U928 (N_928,In_1018,In_921);
nand U929 (N_929,In_1284,In_435);
or U930 (N_930,In_1000,In_961);
xor U931 (N_931,In_316,In_1319);
xnor U932 (N_932,In_266,In_86);
nor U933 (N_933,In_894,In_91);
and U934 (N_934,In_924,In_1027);
nand U935 (N_935,In_1332,In_1111);
or U936 (N_936,In_1270,In_1398);
xnor U937 (N_937,In_18,In_249);
and U938 (N_938,In_789,In_464);
nor U939 (N_939,In_314,In_1406);
and U940 (N_940,In_1446,In_837);
nor U941 (N_941,In_1181,In_65);
and U942 (N_942,In_952,In_420);
and U943 (N_943,In_580,In_642);
xor U944 (N_944,In_1068,In_260);
nor U945 (N_945,In_221,In_43);
or U946 (N_946,In_1325,In_1457);
or U947 (N_947,In_854,In_1094);
and U948 (N_948,In_767,In_1424);
xor U949 (N_949,In_1226,In_6);
nand U950 (N_950,In_337,In_1472);
and U951 (N_951,In_886,In_179);
and U952 (N_952,In_341,In_706);
and U953 (N_953,In_1255,In_573);
and U954 (N_954,In_229,In_1230);
or U955 (N_955,In_67,In_823);
nand U956 (N_956,In_153,In_1382);
or U957 (N_957,In_336,In_1085);
xor U958 (N_958,In_958,In_635);
or U959 (N_959,In_368,In_90);
or U960 (N_960,In_1243,In_850);
and U961 (N_961,In_770,In_322);
nand U962 (N_962,In_61,In_1067);
nand U963 (N_963,In_322,In_1364);
or U964 (N_964,In_169,In_1235);
and U965 (N_965,In_1247,In_532);
and U966 (N_966,In_175,In_38);
or U967 (N_967,In_875,In_21);
and U968 (N_968,In_1084,In_467);
nand U969 (N_969,In_1257,In_550);
or U970 (N_970,In_488,In_821);
nor U971 (N_971,In_762,In_1319);
or U972 (N_972,In_902,In_166);
xnor U973 (N_973,In_1325,In_32);
or U974 (N_974,In_221,In_1469);
nand U975 (N_975,In_938,In_1323);
and U976 (N_976,In_768,In_425);
nor U977 (N_977,In_650,In_612);
and U978 (N_978,In_40,In_936);
and U979 (N_979,In_1479,In_737);
nand U980 (N_980,In_1093,In_1047);
and U981 (N_981,In_865,In_911);
xnor U982 (N_982,In_145,In_263);
or U983 (N_983,In_335,In_1462);
nor U984 (N_984,In_22,In_1172);
nand U985 (N_985,In_321,In_1152);
xnor U986 (N_986,In_1021,In_533);
nor U987 (N_987,In_875,In_328);
xnor U988 (N_988,In_1425,In_773);
nand U989 (N_989,In_1085,In_651);
and U990 (N_990,In_988,In_1191);
or U991 (N_991,In_825,In_384);
xor U992 (N_992,In_102,In_197);
nor U993 (N_993,In_498,In_1096);
nand U994 (N_994,In_1289,In_1194);
and U995 (N_995,In_1084,In_1464);
nor U996 (N_996,In_1473,In_389);
nor U997 (N_997,In_992,In_166);
xor U998 (N_998,In_832,In_200);
and U999 (N_999,In_20,In_921);
and U1000 (N_1000,In_700,In_911);
or U1001 (N_1001,In_662,In_733);
nand U1002 (N_1002,In_205,In_613);
nand U1003 (N_1003,In_1103,In_415);
and U1004 (N_1004,In_1032,In_674);
nand U1005 (N_1005,In_192,In_39);
nor U1006 (N_1006,In_469,In_947);
and U1007 (N_1007,In_1290,In_408);
nor U1008 (N_1008,In_1010,In_96);
nor U1009 (N_1009,In_977,In_1288);
nor U1010 (N_1010,In_1393,In_1185);
nand U1011 (N_1011,In_288,In_1110);
nor U1012 (N_1012,In_1147,In_377);
nand U1013 (N_1013,In_1397,In_1298);
nor U1014 (N_1014,In_883,In_26);
nand U1015 (N_1015,In_1298,In_109);
nor U1016 (N_1016,In_599,In_764);
nor U1017 (N_1017,In_262,In_14);
or U1018 (N_1018,In_1185,In_1152);
xor U1019 (N_1019,In_776,In_687);
or U1020 (N_1020,In_1313,In_1030);
nor U1021 (N_1021,In_604,In_853);
and U1022 (N_1022,In_8,In_770);
nor U1023 (N_1023,In_99,In_1118);
or U1024 (N_1024,In_24,In_672);
xnor U1025 (N_1025,In_36,In_1322);
nand U1026 (N_1026,In_1443,In_1487);
xnor U1027 (N_1027,In_308,In_824);
nand U1028 (N_1028,In_281,In_566);
or U1029 (N_1029,In_686,In_835);
nor U1030 (N_1030,In_48,In_305);
nand U1031 (N_1031,In_1097,In_1239);
or U1032 (N_1032,In_68,In_1380);
and U1033 (N_1033,In_929,In_219);
nand U1034 (N_1034,In_1323,In_1489);
or U1035 (N_1035,In_394,In_1082);
and U1036 (N_1036,In_469,In_568);
and U1037 (N_1037,In_859,In_1408);
nand U1038 (N_1038,In_1273,In_1405);
nand U1039 (N_1039,In_328,In_621);
xor U1040 (N_1040,In_548,In_414);
and U1041 (N_1041,In_1241,In_9);
nand U1042 (N_1042,In_1026,In_1186);
nand U1043 (N_1043,In_1099,In_883);
or U1044 (N_1044,In_730,In_1464);
nor U1045 (N_1045,In_144,In_436);
nand U1046 (N_1046,In_60,In_1360);
nor U1047 (N_1047,In_1240,In_244);
nor U1048 (N_1048,In_1374,In_1142);
nor U1049 (N_1049,In_661,In_94);
xor U1050 (N_1050,In_376,In_922);
or U1051 (N_1051,In_1284,In_1150);
nor U1052 (N_1052,In_100,In_1325);
and U1053 (N_1053,In_1114,In_1118);
nor U1054 (N_1054,In_620,In_667);
and U1055 (N_1055,In_977,In_1341);
nand U1056 (N_1056,In_1363,In_849);
nor U1057 (N_1057,In_1189,In_752);
xnor U1058 (N_1058,In_1347,In_96);
xnor U1059 (N_1059,In_2,In_1211);
and U1060 (N_1060,In_391,In_434);
nand U1061 (N_1061,In_706,In_982);
or U1062 (N_1062,In_22,In_803);
xnor U1063 (N_1063,In_542,In_897);
or U1064 (N_1064,In_973,In_409);
or U1065 (N_1065,In_258,In_489);
or U1066 (N_1066,In_214,In_932);
and U1067 (N_1067,In_999,In_1105);
xnor U1068 (N_1068,In_232,In_1379);
nand U1069 (N_1069,In_516,In_283);
and U1070 (N_1070,In_697,In_1262);
and U1071 (N_1071,In_211,In_735);
xor U1072 (N_1072,In_1465,In_540);
nand U1073 (N_1073,In_27,In_1297);
nand U1074 (N_1074,In_467,In_799);
xor U1075 (N_1075,In_1238,In_750);
nor U1076 (N_1076,In_1131,In_0);
or U1077 (N_1077,In_736,In_1088);
and U1078 (N_1078,In_224,In_154);
and U1079 (N_1079,In_954,In_692);
and U1080 (N_1080,In_203,In_435);
nand U1081 (N_1081,In_317,In_1197);
and U1082 (N_1082,In_1125,In_217);
or U1083 (N_1083,In_1424,In_1262);
nand U1084 (N_1084,In_1250,In_1222);
or U1085 (N_1085,In_1065,In_834);
nor U1086 (N_1086,In_1180,In_869);
nor U1087 (N_1087,In_765,In_793);
nor U1088 (N_1088,In_558,In_224);
nor U1089 (N_1089,In_453,In_1435);
and U1090 (N_1090,In_1457,In_1308);
nor U1091 (N_1091,In_876,In_263);
and U1092 (N_1092,In_261,In_1316);
nor U1093 (N_1093,In_591,In_186);
nand U1094 (N_1094,In_78,In_144);
nor U1095 (N_1095,In_227,In_1218);
nor U1096 (N_1096,In_1144,In_89);
nand U1097 (N_1097,In_528,In_673);
nand U1098 (N_1098,In_796,In_455);
and U1099 (N_1099,In_1411,In_90);
nor U1100 (N_1100,In_703,In_1361);
or U1101 (N_1101,In_327,In_1408);
or U1102 (N_1102,In_1274,In_257);
or U1103 (N_1103,In_871,In_1133);
nor U1104 (N_1104,In_958,In_184);
nor U1105 (N_1105,In_211,In_297);
nor U1106 (N_1106,In_1015,In_547);
or U1107 (N_1107,In_435,In_60);
nand U1108 (N_1108,In_285,In_1289);
nor U1109 (N_1109,In_695,In_1107);
nand U1110 (N_1110,In_676,In_242);
and U1111 (N_1111,In_635,In_213);
or U1112 (N_1112,In_432,In_377);
xor U1113 (N_1113,In_900,In_616);
nand U1114 (N_1114,In_69,In_1148);
nand U1115 (N_1115,In_914,In_828);
and U1116 (N_1116,In_484,In_1038);
nor U1117 (N_1117,In_1249,In_1063);
or U1118 (N_1118,In_911,In_536);
and U1119 (N_1119,In_211,In_1319);
nand U1120 (N_1120,In_257,In_1130);
and U1121 (N_1121,In_1375,In_309);
nor U1122 (N_1122,In_882,In_823);
and U1123 (N_1123,In_1021,In_193);
nand U1124 (N_1124,In_886,In_973);
nand U1125 (N_1125,In_510,In_571);
or U1126 (N_1126,In_1364,In_837);
nand U1127 (N_1127,In_881,In_950);
nand U1128 (N_1128,In_871,In_96);
nor U1129 (N_1129,In_1423,In_249);
or U1130 (N_1130,In_1073,In_1452);
nand U1131 (N_1131,In_837,In_696);
or U1132 (N_1132,In_241,In_966);
nor U1133 (N_1133,In_957,In_660);
nor U1134 (N_1134,In_154,In_238);
nor U1135 (N_1135,In_1389,In_325);
or U1136 (N_1136,In_636,In_253);
or U1137 (N_1137,In_193,In_853);
and U1138 (N_1138,In_1444,In_553);
nor U1139 (N_1139,In_462,In_731);
nand U1140 (N_1140,In_432,In_832);
and U1141 (N_1141,In_663,In_445);
or U1142 (N_1142,In_1295,In_568);
nor U1143 (N_1143,In_125,In_15);
or U1144 (N_1144,In_649,In_1406);
nand U1145 (N_1145,In_118,In_146);
or U1146 (N_1146,In_1048,In_1335);
and U1147 (N_1147,In_431,In_373);
nor U1148 (N_1148,In_1004,In_189);
and U1149 (N_1149,In_321,In_911);
nor U1150 (N_1150,In_618,In_240);
nor U1151 (N_1151,In_34,In_929);
nand U1152 (N_1152,In_930,In_838);
nand U1153 (N_1153,In_1032,In_1112);
and U1154 (N_1154,In_840,In_637);
or U1155 (N_1155,In_1389,In_1259);
or U1156 (N_1156,In_1338,In_370);
or U1157 (N_1157,In_842,In_276);
nand U1158 (N_1158,In_350,In_867);
nor U1159 (N_1159,In_86,In_1424);
and U1160 (N_1160,In_873,In_305);
nand U1161 (N_1161,In_716,In_1025);
xnor U1162 (N_1162,In_1011,In_1424);
or U1163 (N_1163,In_260,In_983);
or U1164 (N_1164,In_1204,In_1321);
nand U1165 (N_1165,In_1281,In_590);
xor U1166 (N_1166,In_1312,In_515);
nor U1167 (N_1167,In_684,In_1357);
and U1168 (N_1168,In_1080,In_140);
or U1169 (N_1169,In_745,In_472);
or U1170 (N_1170,In_1123,In_317);
or U1171 (N_1171,In_834,In_230);
nand U1172 (N_1172,In_529,In_1464);
and U1173 (N_1173,In_350,In_1096);
nand U1174 (N_1174,In_751,In_183);
nor U1175 (N_1175,In_92,In_1325);
and U1176 (N_1176,In_1036,In_222);
xnor U1177 (N_1177,In_675,In_228);
xnor U1178 (N_1178,In_1258,In_131);
and U1179 (N_1179,In_1118,In_1090);
nor U1180 (N_1180,In_1445,In_949);
nand U1181 (N_1181,In_1267,In_543);
xor U1182 (N_1182,In_398,In_506);
and U1183 (N_1183,In_687,In_628);
and U1184 (N_1184,In_1218,In_529);
nor U1185 (N_1185,In_979,In_1449);
nor U1186 (N_1186,In_657,In_293);
or U1187 (N_1187,In_279,In_1412);
nand U1188 (N_1188,In_210,In_1376);
nor U1189 (N_1189,In_522,In_1465);
xor U1190 (N_1190,In_243,In_220);
nor U1191 (N_1191,In_273,In_107);
nor U1192 (N_1192,In_872,In_173);
and U1193 (N_1193,In_185,In_473);
nand U1194 (N_1194,In_1464,In_278);
nand U1195 (N_1195,In_1453,In_223);
nor U1196 (N_1196,In_1116,In_1157);
and U1197 (N_1197,In_1125,In_167);
nand U1198 (N_1198,In_467,In_28);
and U1199 (N_1199,In_1450,In_598);
and U1200 (N_1200,In_206,In_1012);
nand U1201 (N_1201,In_796,In_638);
or U1202 (N_1202,In_1061,In_1280);
nand U1203 (N_1203,In_1433,In_57);
nand U1204 (N_1204,In_1327,In_191);
nor U1205 (N_1205,In_1220,In_364);
and U1206 (N_1206,In_1224,In_563);
or U1207 (N_1207,In_1291,In_1028);
xnor U1208 (N_1208,In_1056,In_152);
and U1209 (N_1209,In_1359,In_333);
nor U1210 (N_1210,In_1336,In_116);
and U1211 (N_1211,In_1425,In_420);
nand U1212 (N_1212,In_194,In_37);
or U1213 (N_1213,In_913,In_855);
and U1214 (N_1214,In_833,In_659);
or U1215 (N_1215,In_334,In_827);
nand U1216 (N_1216,In_425,In_679);
nand U1217 (N_1217,In_1268,In_513);
or U1218 (N_1218,In_133,In_1408);
or U1219 (N_1219,In_144,In_1191);
xnor U1220 (N_1220,In_963,In_68);
xnor U1221 (N_1221,In_946,In_1171);
or U1222 (N_1222,In_816,In_830);
nand U1223 (N_1223,In_1124,In_559);
nand U1224 (N_1224,In_532,In_493);
and U1225 (N_1225,In_1265,In_975);
nor U1226 (N_1226,In_191,In_159);
and U1227 (N_1227,In_432,In_778);
xor U1228 (N_1228,In_343,In_51);
and U1229 (N_1229,In_374,In_53);
and U1230 (N_1230,In_228,In_1187);
xnor U1231 (N_1231,In_865,In_1245);
and U1232 (N_1232,In_870,In_715);
nand U1233 (N_1233,In_344,In_518);
or U1234 (N_1234,In_371,In_1375);
nor U1235 (N_1235,In_926,In_249);
nand U1236 (N_1236,In_1106,In_658);
or U1237 (N_1237,In_1113,In_967);
nor U1238 (N_1238,In_1321,In_217);
and U1239 (N_1239,In_276,In_1424);
nor U1240 (N_1240,In_402,In_147);
nor U1241 (N_1241,In_1491,In_263);
and U1242 (N_1242,In_1226,In_1216);
nor U1243 (N_1243,In_341,In_651);
nor U1244 (N_1244,In_552,In_1264);
nand U1245 (N_1245,In_1338,In_1266);
xnor U1246 (N_1246,In_120,In_565);
nand U1247 (N_1247,In_897,In_195);
nor U1248 (N_1248,In_1269,In_111);
nand U1249 (N_1249,In_49,In_1432);
or U1250 (N_1250,In_450,In_174);
nor U1251 (N_1251,In_1132,In_519);
and U1252 (N_1252,In_724,In_137);
or U1253 (N_1253,In_319,In_496);
or U1254 (N_1254,In_1180,In_1287);
nor U1255 (N_1255,In_1481,In_1023);
nand U1256 (N_1256,In_249,In_684);
nor U1257 (N_1257,In_1267,In_897);
or U1258 (N_1258,In_1235,In_1393);
xor U1259 (N_1259,In_809,In_746);
and U1260 (N_1260,In_248,In_650);
xor U1261 (N_1261,In_1467,In_1353);
nor U1262 (N_1262,In_499,In_607);
nand U1263 (N_1263,In_178,In_540);
nand U1264 (N_1264,In_1125,In_1399);
and U1265 (N_1265,In_756,In_1092);
and U1266 (N_1266,In_655,In_641);
nor U1267 (N_1267,In_1433,In_555);
nor U1268 (N_1268,In_439,In_221);
or U1269 (N_1269,In_1092,In_1277);
or U1270 (N_1270,In_208,In_679);
nor U1271 (N_1271,In_1093,In_503);
and U1272 (N_1272,In_894,In_666);
or U1273 (N_1273,In_1056,In_996);
or U1274 (N_1274,In_1206,In_585);
or U1275 (N_1275,In_283,In_561);
and U1276 (N_1276,In_758,In_908);
nor U1277 (N_1277,In_670,In_722);
and U1278 (N_1278,In_875,In_1200);
nand U1279 (N_1279,In_871,In_161);
nor U1280 (N_1280,In_1482,In_540);
and U1281 (N_1281,In_695,In_1131);
and U1282 (N_1282,In_334,In_1286);
and U1283 (N_1283,In_1466,In_1031);
nor U1284 (N_1284,In_746,In_267);
and U1285 (N_1285,In_722,In_521);
and U1286 (N_1286,In_1047,In_163);
nand U1287 (N_1287,In_1387,In_878);
xor U1288 (N_1288,In_1205,In_555);
and U1289 (N_1289,In_825,In_744);
nor U1290 (N_1290,In_490,In_477);
or U1291 (N_1291,In_443,In_490);
and U1292 (N_1292,In_1208,In_34);
and U1293 (N_1293,In_910,In_267);
nand U1294 (N_1294,In_714,In_1455);
nor U1295 (N_1295,In_1093,In_708);
nor U1296 (N_1296,In_967,In_489);
nand U1297 (N_1297,In_245,In_364);
and U1298 (N_1298,In_1148,In_543);
nor U1299 (N_1299,In_401,In_972);
nor U1300 (N_1300,In_1072,In_358);
and U1301 (N_1301,In_758,In_728);
nand U1302 (N_1302,In_1496,In_474);
nand U1303 (N_1303,In_408,In_185);
and U1304 (N_1304,In_1096,In_592);
and U1305 (N_1305,In_313,In_147);
nor U1306 (N_1306,In_1298,In_1361);
nand U1307 (N_1307,In_513,In_990);
nor U1308 (N_1308,In_742,In_944);
nand U1309 (N_1309,In_432,In_604);
or U1310 (N_1310,In_548,In_1057);
or U1311 (N_1311,In_619,In_865);
and U1312 (N_1312,In_456,In_1306);
nor U1313 (N_1313,In_620,In_1230);
and U1314 (N_1314,In_923,In_1355);
nor U1315 (N_1315,In_311,In_904);
nand U1316 (N_1316,In_1347,In_1242);
or U1317 (N_1317,In_1297,In_1463);
xor U1318 (N_1318,In_683,In_887);
nand U1319 (N_1319,In_689,In_312);
xor U1320 (N_1320,In_428,In_681);
nand U1321 (N_1321,In_1451,In_430);
nor U1322 (N_1322,In_1146,In_662);
xor U1323 (N_1323,In_1297,In_238);
nor U1324 (N_1324,In_350,In_266);
or U1325 (N_1325,In_8,In_1475);
nand U1326 (N_1326,In_1273,In_1022);
or U1327 (N_1327,In_862,In_1496);
nand U1328 (N_1328,In_244,In_159);
nor U1329 (N_1329,In_1228,In_663);
nor U1330 (N_1330,In_700,In_447);
nor U1331 (N_1331,In_442,In_779);
nand U1332 (N_1332,In_815,In_824);
nor U1333 (N_1333,In_241,In_490);
nor U1334 (N_1334,In_636,In_1282);
and U1335 (N_1335,In_1465,In_1);
nand U1336 (N_1336,In_1250,In_734);
and U1337 (N_1337,In_1421,In_64);
nand U1338 (N_1338,In_811,In_193);
and U1339 (N_1339,In_1165,In_156);
nor U1340 (N_1340,In_806,In_824);
and U1341 (N_1341,In_520,In_1267);
nand U1342 (N_1342,In_206,In_1060);
nor U1343 (N_1343,In_714,In_1138);
nor U1344 (N_1344,In_19,In_815);
nand U1345 (N_1345,In_584,In_778);
and U1346 (N_1346,In_14,In_764);
and U1347 (N_1347,In_863,In_64);
or U1348 (N_1348,In_1024,In_45);
nor U1349 (N_1349,In_167,In_40);
nand U1350 (N_1350,In_711,In_580);
nor U1351 (N_1351,In_65,In_276);
and U1352 (N_1352,In_754,In_506);
or U1353 (N_1353,In_75,In_1202);
nand U1354 (N_1354,In_1318,In_569);
and U1355 (N_1355,In_866,In_1279);
and U1356 (N_1356,In_643,In_121);
nand U1357 (N_1357,In_1321,In_1019);
nor U1358 (N_1358,In_416,In_926);
nand U1359 (N_1359,In_177,In_1431);
and U1360 (N_1360,In_915,In_352);
nand U1361 (N_1361,In_1066,In_257);
or U1362 (N_1362,In_235,In_1493);
nand U1363 (N_1363,In_782,In_315);
or U1364 (N_1364,In_251,In_879);
and U1365 (N_1365,In_1397,In_708);
and U1366 (N_1366,In_139,In_862);
nand U1367 (N_1367,In_681,In_611);
or U1368 (N_1368,In_1465,In_1066);
nand U1369 (N_1369,In_956,In_1109);
nand U1370 (N_1370,In_889,In_107);
nor U1371 (N_1371,In_912,In_1267);
nor U1372 (N_1372,In_762,In_35);
nand U1373 (N_1373,In_828,In_1409);
nand U1374 (N_1374,In_259,In_1286);
and U1375 (N_1375,In_644,In_164);
nand U1376 (N_1376,In_35,In_512);
nand U1377 (N_1377,In_111,In_906);
nand U1378 (N_1378,In_1447,In_337);
and U1379 (N_1379,In_179,In_374);
and U1380 (N_1380,In_1109,In_0);
and U1381 (N_1381,In_528,In_186);
nand U1382 (N_1382,In_1219,In_689);
or U1383 (N_1383,In_37,In_95);
nand U1384 (N_1384,In_623,In_1057);
nor U1385 (N_1385,In_1312,In_1154);
xnor U1386 (N_1386,In_89,In_641);
and U1387 (N_1387,In_1358,In_953);
or U1388 (N_1388,In_337,In_210);
or U1389 (N_1389,In_743,In_52);
and U1390 (N_1390,In_147,In_874);
and U1391 (N_1391,In_1007,In_975);
nor U1392 (N_1392,In_1153,In_149);
nand U1393 (N_1393,In_345,In_787);
and U1394 (N_1394,In_574,In_733);
xor U1395 (N_1395,In_1421,In_1252);
nand U1396 (N_1396,In_1122,In_198);
nand U1397 (N_1397,In_376,In_1441);
and U1398 (N_1398,In_477,In_1092);
xnor U1399 (N_1399,In_279,In_552);
nand U1400 (N_1400,In_733,In_444);
nand U1401 (N_1401,In_120,In_169);
or U1402 (N_1402,In_127,In_237);
nand U1403 (N_1403,In_426,In_1185);
or U1404 (N_1404,In_231,In_1047);
nand U1405 (N_1405,In_478,In_1017);
or U1406 (N_1406,In_749,In_621);
nor U1407 (N_1407,In_1006,In_1067);
nor U1408 (N_1408,In_846,In_803);
or U1409 (N_1409,In_705,In_270);
nor U1410 (N_1410,In_794,In_293);
nor U1411 (N_1411,In_1394,In_1210);
or U1412 (N_1412,In_785,In_1052);
nand U1413 (N_1413,In_842,In_1049);
nor U1414 (N_1414,In_1002,In_362);
and U1415 (N_1415,In_1214,In_1375);
xor U1416 (N_1416,In_1194,In_367);
or U1417 (N_1417,In_669,In_873);
nor U1418 (N_1418,In_559,In_389);
xnor U1419 (N_1419,In_267,In_462);
or U1420 (N_1420,In_1246,In_980);
nand U1421 (N_1421,In_721,In_819);
xnor U1422 (N_1422,In_1403,In_1178);
nand U1423 (N_1423,In_714,In_429);
and U1424 (N_1424,In_1399,In_745);
nand U1425 (N_1425,In_618,In_539);
nand U1426 (N_1426,In_1044,In_1323);
or U1427 (N_1427,In_924,In_1322);
and U1428 (N_1428,In_1272,In_1197);
and U1429 (N_1429,In_253,In_1280);
nand U1430 (N_1430,In_1454,In_455);
or U1431 (N_1431,In_623,In_34);
and U1432 (N_1432,In_892,In_1405);
and U1433 (N_1433,In_577,In_190);
nand U1434 (N_1434,In_117,In_679);
xnor U1435 (N_1435,In_204,In_1202);
nand U1436 (N_1436,In_795,In_49);
and U1437 (N_1437,In_622,In_225);
nor U1438 (N_1438,In_1387,In_1428);
or U1439 (N_1439,In_565,In_229);
and U1440 (N_1440,In_947,In_94);
or U1441 (N_1441,In_381,In_428);
or U1442 (N_1442,In_700,In_1021);
or U1443 (N_1443,In_856,In_932);
nor U1444 (N_1444,In_317,In_207);
nor U1445 (N_1445,In_1255,In_1221);
nand U1446 (N_1446,In_39,In_757);
and U1447 (N_1447,In_304,In_554);
and U1448 (N_1448,In_110,In_376);
nand U1449 (N_1449,In_1151,In_1202);
nand U1450 (N_1450,In_1350,In_1113);
or U1451 (N_1451,In_15,In_383);
nor U1452 (N_1452,In_818,In_507);
nor U1453 (N_1453,In_1236,In_547);
or U1454 (N_1454,In_456,In_1087);
and U1455 (N_1455,In_132,In_776);
and U1456 (N_1456,In_1055,In_755);
nor U1457 (N_1457,In_1433,In_229);
nand U1458 (N_1458,In_253,In_996);
or U1459 (N_1459,In_644,In_1450);
or U1460 (N_1460,In_537,In_301);
nor U1461 (N_1461,In_1018,In_88);
and U1462 (N_1462,In_1488,In_289);
nor U1463 (N_1463,In_1414,In_208);
nor U1464 (N_1464,In_898,In_867);
or U1465 (N_1465,In_860,In_289);
and U1466 (N_1466,In_573,In_1281);
nand U1467 (N_1467,In_468,In_1127);
or U1468 (N_1468,In_783,In_1042);
and U1469 (N_1469,In_695,In_1427);
nor U1470 (N_1470,In_79,In_92);
nand U1471 (N_1471,In_12,In_753);
or U1472 (N_1472,In_1418,In_203);
and U1473 (N_1473,In_430,In_1336);
nor U1474 (N_1474,In_68,In_948);
nor U1475 (N_1475,In_1025,In_653);
nand U1476 (N_1476,In_1385,In_399);
or U1477 (N_1477,In_698,In_217);
nor U1478 (N_1478,In_390,In_771);
nand U1479 (N_1479,In_50,In_1431);
or U1480 (N_1480,In_1315,In_96);
nor U1481 (N_1481,In_1181,In_1030);
and U1482 (N_1482,In_418,In_1389);
and U1483 (N_1483,In_500,In_772);
nor U1484 (N_1484,In_767,In_1415);
xnor U1485 (N_1485,In_335,In_686);
nand U1486 (N_1486,In_860,In_845);
and U1487 (N_1487,In_704,In_316);
nand U1488 (N_1488,In_303,In_95);
xnor U1489 (N_1489,In_918,In_1081);
or U1490 (N_1490,In_999,In_209);
xnor U1491 (N_1491,In_1125,In_805);
and U1492 (N_1492,In_1258,In_945);
nand U1493 (N_1493,In_257,In_1323);
nand U1494 (N_1494,In_855,In_1337);
xnor U1495 (N_1495,In_1136,In_150);
and U1496 (N_1496,In_997,In_946);
or U1497 (N_1497,In_1115,In_356);
nor U1498 (N_1498,In_698,In_549);
or U1499 (N_1499,In_277,In_346);
and U1500 (N_1500,N_561,N_689);
nor U1501 (N_1501,N_894,N_570);
nor U1502 (N_1502,N_695,N_1299);
xnor U1503 (N_1503,N_152,N_1328);
nor U1504 (N_1504,N_1158,N_1449);
and U1505 (N_1505,N_338,N_273);
or U1506 (N_1506,N_66,N_1488);
and U1507 (N_1507,N_390,N_451);
xor U1508 (N_1508,N_721,N_912);
nand U1509 (N_1509,N_1373,N_1453);
nor U1510 (N_1510,N_168,N_357);
nand U1511 (N_1511,N_190,N_95);
nor U1512 (N_1512,N_491,N_1413);
nor U1513 (N_1513,N_995,N_481);
and U1514 (N_1514,N_1211,N_910);
nand U1515 (N_1515,N_517,N_895);
nor U1516 (N_1516,N_196,N_1232);
xnor U1517 (N_1517,N_205,N_512);
and U1518 (N_1518,N_239,N_226);
nand U1519 (N_1519,N_666,N_128);
nand U1520 (N_1520,N_1244,N_1274);
or U1521 (N_1521,N_1452,N_313);
nor U1522 (N_1522,N_1256,N_576);
or U1523 (N_1523,N_90,N_39);
or U1524 (N_1524,N_796,N_137);
nand U1525 (N_1525,N_307,N_443);
or U1526 (N_1526,N_597,N_891);
and U1527 (N_1527,N_899,N_765);
or U1528 (N_1528,N_464,N_1147);
or U1529 (N_1529,N_1041,N_636);
nor U1530 (N_1530,N_474,N_377);
nor U1531 (N_1531,N_658,N_672);
nor U1532 (N_1532,N_1411,N_601);
and U1533 (N_1533,N_1149,N_106);
nand U1534 (N_1534,N_497,N_1255);
nor U1535 (N_1535,N_642,N_982);
nor U1536 (N_1536,N_777,N_203);
and U1537 (N_1537,N_678,N_20);
nor U1538 (N_1538,N_957,N_1166);
and U1539 (N_1539,N_1354,N_109);
nor U1540 (N_1540,N_1026,N_865);
xnor U1541 (N_1541,N_1098,N_583);
and U1542 (N_1542,N_424,N_1151);
nor U1543 (N_1543,N_1050,N_581);
nor U1544 (N_1544,N_732,N_1421);
nand U1545 (N_1545,N_355,N_855);
nand U1546 (N_1546,N_10,N_1068);
nor U1547 (N_1547,N_404,N_696);
nand U1548 (N_1548,N_1367,N_644);
and U1549 (N_1549,N_124,N_1187);
or U1550 (N_1550,N_905,N_1125);
nor U1551 (N_1551,N_857,N_734);
or U1552 (N_1552,N_402,N_316);
or U1553 (N_1553,N_1227,N_235);
xor U1554 (N_1554,N_192,N_122);
and U1555 (N_1555,N_225,N_1445);
or U1556 (N_1556,N_1215,N_242);
xnor U1557 (N_1557,N_690,N_64);
or U1558 (N_1558,N_94,N_155);
nor U1559 (N_1559,N_674,N_448);
and U1560 (N_1560,N_646,N_484);
and U1561 (N_1561,N_923,N_426);
nand U1562 (N_1562,N_574,N_963);
nor U1563 (N_1563,N_897,N_6);
and U1564 (N_1564,N_1303,N_1217);
nor U1565 (N_1565,N_1469,N_573);
nor U1566 (N_1566,N_1218,N_766);
nor U1567 (N_1567,N_1014,N_80);
nand U1568 (N_1568,N_1330,N_1038);
nand U1569 (N_1569,N_29,N_1353);
and U1570 (N_1570,N_476,N_1175);
nor U1571 (N_1571,N_121,N_111);
and U1572 (N_1572,N_1203,N_300);
nand U1573 (N_1573,N_548,N_1495);
xnor U1574 (N_1574,N_379,N_1356);
nor U1575 (N_1575,N_293,N_7);
nand U1576 (N_1576,N_826,N_255);
nor U1577 (N_1577,N_544,N_340);
or U1578 (N_1578,N_1403,N_57);
nor U1579 (N_1579,N_1333,N_420);
and U1580 (N_1580,N_1129,N_904);
and U1581 (N_1581,N_858,N_578);
nand U1582 (N_1582,N_1262,N_1365);
and U1583 (N_1583,N_1165,N_913);
xor U1584 (N_1584,N_656,N_1432);
and U1585 (N_1585,N_1182,N_840);
nor U1586 (N_1586,N_483,N_643);
or U1587 (N_1587,N_233,N_50);
and U1588 (N_1588,N_639,N_1221);
or U1589 (N_1589,N_1079,N_1347);
nor U1590 (N_1590,N_1318,N_1275);
or U1591 (N_1591,N_1065,N_1295);
nand U1592 (N_1592,N_1200,N_728);
nor U1593 (N_1593,N_44,N_538);
or U1594 (N_1594,N_279,N_286);
nor U1595 (N_1595,N_392,N_1118);
and U1596 (N_1596,N_565,N_413);
nor U1597 (N_1597,N_489,N_798);
and U1598 (N_1598,N_1185,N_1020);
nor U1599 (N_1599,N_475,N_388);
or U1600 (N_1600,N_405,N_385);
and U1601 (N_1601,N_1342,N_793);
or U1602 (N_1602,N_1241,N_113);
nor U1603 (N_1603,N_353,N_669);
nor U1604 (N_1604,N_1131,N_1039);
or U1605 (N_1605,N_968,N_1101);
and U1606 (N_1606,N_993,N_622);
nand U1607 (N_1607,N_188,N_148);
xnor U1608 (N_1608,N_1315,N_169);
xnor U1609 (N_1609,N_82,N_958);
nand U1610 (N_1610,N_909,N_318);
nand U1611 (N_1611,N_1176,N_709);
nand U1612 (N_1612,N_815,N_1183);
or U1613 (N_1613,N_825,N_1460);
or U1614 (N_1614,N_432,N_1035);
nor U1615 (N_1615,N_36,N_181);
and U1616 (N_1616,N_1458,N_1338);
nor U1617 (N_1617,N_584,N_72);
or U1618 (N_1618,N_1252,N_976);
or U1619 (N_1619,N_1097,N_753);
nor U1620 (N_1620,N_372,N_979);
and U1621 (N_1621,N_662,N_860);
and U1622 (N_1622,N_408,N_737);
or U1623 (N_1623,N_65,N_1385);
nand U1624 (N_1624,N_810,N_1459);
or U1625 (N_1625,N_668,N_911);
and U1626 (N_1626,N_1376,N_1161);
and U1627 (N_1627,N_505,N_216);
nor U1628 (N_1628,N_1340,N_795);
nor U1629 (N_1629,N_150,N_527);
nand U1630 (N_1630,N_1181,N_592);
nor U1631 (N_1631,N_247,N_705);
nor U1632 (N_1632,N_1369,N_454);
and U1633 (N_1633,N_240,N_692);
nor U1634 (N_1634,N_711,N_1420);
xnor U1635 (N_1635,N_49,N_1194);
and U1636 (N_1636,N_944,N_149);
or U1637 (N_1637,N_163,N_1423);
or U1638 (N_1638,N_32,N_492);
nand U1639 (N_1639,N_362,N_16);
nand U1640 (N_1640,N_579,N_783);
and U1641 (N_1641,N_1424,N_381);
xnor U1642 (N_1642,N_1384,N_1132);
nor U1643 (N_1643,N_934,N_369);
or U1644 (N_1644,N_1427,N_302);
nor U1645 (N_1645,N_1372,N_1243);
and U1646 (N_1646,N_1152,N_319);
and U1647 (N_1647,N_321,N_829);
or U1648 (N_1648,N_530,N_496);
nand U1649 (N_1649,N_540,N_482);
nor U1650 (N_1650,N_1063,N_760);
or U1651 (N_1651,N_789,N_972);
or U1652 (N_1652,N_68,N_1293);
nand U1653 (N_1653,N_470,N_1276);
or U1654 (N_1654,N_959,N_174);
or U1655 (N_1655,N_844,N_43);
nand U1656 (N_1656,N_81,N_661);
and U1657 (N_1657,N_1091,N_1085);
and U1658 (N_1658,N_1408,N_136);
or U1659 (N_1659,N_193,N_1378);
xnor U1660 (N_1660,N_359,N_1419);
nor U1661 (N_1661,N_553,N_845);
xnor U1662 (N_1662,N_564,N_232);
and U1663 (N_1663,N_344,N_1444);
nor U1664 (N_1664,N_613,N_1350);
and U1665 (N_1665,N_277,N_23);
nand U1666 (N_1666,N_585,N_699);
and U1667 (N_1667,N_189,N_1220);
nor U1668 (N_1668,N_1280,N_433);
nand U1669 (N_1669,N_1180,N_1261);
or U1670 (N_1670,N_722,N_473);
and U1671 (N_1671,N_1455,N_1226);
nand U1672 (N_1672,N_983,N_294);
nor U1673 (N_1673,N_182,N_373);
or U1674 (N_1674,N_851,N_875);
and U1675 (N_1675,N_918,N_1381);
and U1676 (N_1676,N_1389,N_1489);
and U1677 (N_1677,N_490,N_363);
and U1678 (N_1678,N_1134,N_998);
and U1679 (N_1679,N_237,N_389);
nand U1680 (N_1680,N_202,N_1172);
nor U1681 (N_1681,N_973,N_871);
nor U1682 (N_1682,N_1382,N_1164);
or U1683 (N_1683,N_1402,N_38);
xnor U1684 (N_1684,N_1466,N_364);
and U1685 (N_1685,N_422,N_114);
and U1686 (N_1686,N_807,N_477);
nor U1687 (N_1687,N_323,N_1162);
or U1688 (N_1688,N_403,N_1437);
xnor U1689 (N_1689,N_681,N_738);
nor U1690 (N_1690,N_281,N_507);
nor U1691 (N_1691,N_1012,N_542);
nand U1692 (N_1692,N_1179,N_160);
or U1693 (N_1693,N_41,N_515);
and U1694 (N_1694,N_394,N_1105);
and U1695 (N_1695,N_42,N_442);
xor U1696 (N_1696,N_261,N_1054);
and U1697 (N_1697,N_595,N_1407);
nand U1698 (N_1698,N_593,N_882);
nand U1699 (N_1699,N_817,N_856);
and U1700 (N_1700,N_556,N_466);
xnor U1701 (N_1701,N_1298,N_980);
and U1702 (N_1702,N_1268,N_499);
and U1703 (N_1703,N_741,N_267);
xnor U1704 (N_1704,N_134,N_92);
and U1705 (N_1705,N_1249,N_1112);
or U1706 (N_1706,N_125,N_673);
xnor U1707 (N_1707,N_1399,N_1492);
or U1708 (N_1708,N_932,N_1474);
nor U1709 (N_1709,N_1076,N_1145);
and U1710 (N_1710,N_179,N_1345);
nor U1711 (N_1711,N_131,N_735);
nor U1712 (N_1712,N_212,N_532);
or U1713 (N_1713,N_487,N_1092);
nand U1714 (N_1714,N_914,N_521);
nor U1715 (N_1715,N_986,N_511);
nand U1716 (N_1716,N_1009,N_230);
or U1717 (N_1717,N_1248,N_652);
nor U1718 (N_1718,N_1394,N_1360);
or U1719 (N_1719,N_435,N_693);
nor U1720 (N_1720,N_218,N_606);
nor U1721 (N_1721,N_291,N_764);
nand U1722 (N_1722,N_902,N_272);
or U1723 (N_1723,N_145,N_1425);
nor U1724 (N_1724,N_609,N_749);
and U1725 (N_1725,N_602,N_407);
or U1726 (N_1726,N_98,N_587);
xnor U1727 (N_1727,N_1102,N_1059);
or U1728 (N_1728,N_621,N_616);
and U1729 (N_1729,N_206,N_378);
and U1730 (N_1730,N_1374,N_1106);
and U1731 (N_1731,N_784,N_1088);
or U1732 (N_1732,N_1370,N_869);
and U1733 (N_1733,N_1480,N_221);
and U1734 (N_1734,N_841,N_854);
and U1735 (N_1735,N_770,N_1081);
and U1736 (N_1736,N_526,N_1084);
nand U1737 (N_1737,N_727,N_701);
and U1738 (N_1738,N_522,N_370);
nor U1739 (N_1739,N_356,N_309);
or U1740 (N_1740,N_289,N_920);
xor U1741 (N_1741,N_1406,N_271);
xor U1742 (N_1742,N_623,N_717);
nor U1743 (N_1743,N_1017,N_4);
or U1744 (N_1744,N_867,N_1349);
nor U1745 (N_1745,N_813,N_71);
xor U1746 (N_1746,N_335,N_520);
xor U1747 (N_1747,N_410,N_518);
or U1748 (N_1748,N_686,N_1380);
and U1749 (N_1749,N_1077,N_423);
xor U1750 (N_1750,N_224,N_1311);
nor U1751 (N_1751,N_447,N_1351);
and U1752 (N_1752,N_933,N_1301);
and U1753 (N_1753,N_1148,N_663);
xnor U1754 (N_1754,N_414,N_1337);
nor U1755 (N_1755,N_115,N_22);
and U1756 (N_1756,N_679,N_478);
nor U1757 (N_1757,N_1143,N_1410);
and U1758 (N_1758,N_1484,N_1352);
nor U1759 (N_1759,N_525,N_1302);
and U1760 (N_1760,N_384,N_627);
nand U1761 (N_1761,N_371,N_768);
nor U1762 (N_1762,N_37,N_393);
and U1763 (N_1763,N_791,N_682);
nand U1764 (N_1764,N_1082,N_396);
nand U1765 (N_1765,N_1485,N_450);
xnor U1766 (N_1766,N_926,N_901);
nand U1767 (N_1767,N_698,N_1477);
nor U1768 (N_1768,N_1048,N_758);
or U1769 (N_1769,N_142,N_74);
and U1770 (N_1770,N_214,N_468);
nor U1771 (N_1771,N_295,N_987);
nand U1772 (N_1772,N_1156,N_870);
nor U1773 (N_1773,N_931,N_614);
nand U1774 (N_1774,N_1364,N_415);
or U1775 (N_1775,N_1053,N_89);
nor U1776 (N_1776,N_346,N_1289);
xnor U1777 (N_1777,N_1387,N_645);
nand U1778 (N_1778,N_1,N_61);
and U1779 (N_1779,N_594,N_996);
or U1780 (N_1780,N_1168,N_440);
and U1781 (N_1781,N_251,N_219);
and U1782 (N_1782,N_11,N_1023);
or U1783 (N_1783,N_1154,N_781);
and U1784 (N_1784,N_397,N_1032);
nand U1785 (N_1785,N_848,N_731);
or U1786 (N_1786,N_519,N_1309);
xnor U1787 (N_1787,N_619,N_1201);
and U1788 (N_1788,N_1117,N_898);
nor U1789 (N_1789,N_1095,N_776);
xor U1790 (N_1790,N_461,N_266);
xor U1791 (N_1791,N_1324,N_1319);
and U1792 (N_1792,N_685,N_1003);
and U1793 (N_1793,N_1358,N_697);
and U1794 (N_1794,N_480,N_937);
and U1795 (N_1795,N_1044,N_400);
nor U1796 (N_1796,N_655,N_1078);
and U1797 (N_1797,N_108,N_366);
and U1798 (N_1798,N_861,N_1133);
nand U1799 (N_1799,N_1290,N_183);
nand U1800 (N_1800,N_651,N_1173);
and U1801 (N_1801,N_157,N_588);
nor U1802 (N_1802,N_624,N_284);
or U1803 (N_1803,N_1006,N_533);
or U1804 (N_1804,N_332,N_751);
nand U1805 (N_1805,N_767,N_649);
nand U1806 (N_1806,N_387,N_1482);
and U1807 (N_1807,N_195,N_812);
nand U1808 (N_1808,N_1171,N_1135);
nand U1809 (N_1809,N_243,N_1368);
or U1810 (N_1810,N_1391,N_1074);
nor U1811 (N_1811,N_437,N_774);
xor U1812 (N_1812,N_1481,N_1283);
and U1813 (N_1813,N_637,N_1198);
xnor U1814 (N_1814,N_1110,N_514);
nor U1815 (N_1815,N_462,N_1379);
or U1816 (N_1816,N_165,N_1062);
nand U1817 (N_1817,N_536,N_27);
nor U1818 (N_1818,N_329,N_199);
or U1819 (N_1819,N_1027,N_740);
nor U1820 (N_1820,N_1467,N_969);
nor U1821 (N_1821,N_63,N_1028);
nand U1822 (N_1822,N_1121,N_215);
nor U1823 (N_1823,N_809,N_1308);
xor U1824 (N_1824,N_305,N_1208);
nor U1825 (N_1825,N_1069,N_175);
xnor U1826 (N_1826,N_1314,N_1470);
nor U1827 (N_1827,N_1055,N_1216);
or U1828 (N_1828,N_1426,N_978);
xnor U1829 (N_1829,N_1089,N_962);
nand U1830 (N_1830,N_1417,N_974);
nor U1831 (N_1831,N_187,N_504);
or U1832 (N_1832,N_151,N_33);
and U1833 (N_1833,N_792,N_463);
xor U1834 (N_1834,N_1355,N_1439);
nor U1835 (N_1835,N_1184,N_269);
and U1836 (N_1836,N_772,N_1253);
nor U1837 (N_1837,N_782,N_1259);
and U1838 (N_1838,N_1321,N_1199);
and U1839 (N_1839,N_1416,N_494);
or U1840 (N_1840,N_778,N_427);
or U1841 (N_1841,N_874,N_1479);
xor U1842 (N_1842,N_1235,N_1435);
and U1843 (N_1843,N_949,N_757);
or U1844 (N_1844,N_2,N_984);
nand U1845 (N_1845,N_1343,N_850);
xor U1846 (N_1846,N_1433,N_887);
nand U1847 (N_1847,N_950,N_118);
nand U1848 (N_1848,N_406,N_1212);
nand U1849 (N_1849,N_660,N_391);
or U1850 (N_1850,N_900,N_1291);
and U1851 (N_1851,N_1103,N_859);
and U1852 (N_1852,N_1093,N_325);
nand U1853 (N_1853,N_945,N_1113);
or U1854 (N_1854,N_752,N_47);
and U1855 (N_1855,N_285,N_785);
or U1856 (N_1856,N_105,N_469);
and U1857 (N_1857,N_1031,N_1177);
and U1858 (N_1858,N_452,N_209);
or U1859 (N_1859,N_297,N_939);
and U1860 (N_1860,N_1141,N_186);
nand U1861 (N_1861,N_715,N_1042);
and U1862 (N_1862,N_971,N_58);
and U1863 (N_1863,N_927,N_1163);
or U1864 (N_1864,N_317,N_201);
and U1865 (N_1865,N_418,N_1300);
nand U1866 (N_1866,N_331,N_811);
nor U1867 (N_1867,N_1230,N_31);
nand U1868 (N_1868,N_1285,N_1204);
xor U1869 (N_1869,N_822,N_1155);
and U1870 (N_1870,N_311,N_46);
and U1871 (N_1871,N_797,N_683);
nor U1872 (N_1872,N_398,N_1499);
xor U1873 (N_1873,N_1206,N_264);
or U1874 (N_1874,N_1107,N_1128);
nor U1875 (N_1875,N_358,N_546);
nand U1876 (N_1876,N_1071,N_723);
nor U1877 (N_1877,N_558,N_970);
nand U1878 (N_1878,N_582,N_431);
nor U1879 (N_1879,N_110,N_453);
or U1880 (N_1880,N_1116,N_167);
or U1881 (N_1881,N_940,N_893);
or U1882 (N_1882,N_234,N_1294);
xnor U1883 (N_1883,N_1130,N_1266);
xor U1884 (N_1884,N_290,N_936);
nor U1885 (N_1885,N_953,N_1386);
and U1886 (N_1886,N_176,N_327);
nand U1887 (N_1887,N_560,N_287);
nor U1888 (N_1888,N_127,N_720);
nand U1889 (N_1889,N_1094,N_298);
xor U1890 (N_1890,N_162,N_1336);
and U1891 (N_1891,N_523,N_703);
nand U1892 (N_1892,N_77,N_180);
and U1893 (N_1893,N_1418,N_1224);
and U1894 (N_1894,N_1144,N_1451);
xor U1895 (N_1895,N_460,N_383);
nand U1896 (N_1896,N_1405,N_1138);
or U1897 (N_1897,N_952,N_743);
and U1898 (N_1898,N_1316,N_1277);
nor U1899 (N_1899,N_1335,N_177);
or U1900 (N_1900,N_399,N_1346);
nand U1901 (N_1901,N_754,N_629);
or U1902 (N_1902,N_70,N_827);
or U1903 (N_1903,N_547,N_1496);
nand U1904 (N_1904,N_1011,N_191);
or U1905 (N_1905,N_830,N_19);
nand U1906 (N_1906,N_376,N_677);
or U1907 (N_1907,N_630,N_742);
or U1908 (N_1908,N_129,N_1339);
nand U1909 (N_1909,N_991,N_253);
or U1910 (N_1910,N_270,N_528);
and U1911 (N_1911,N_563,N_550);
or U1912 (N_1912,N_535,N_1051);
nand U1913 (N_1913,N_710,N_541);
xnor U1914 (N_1914,N_278,N_946);
and U1915 (N_1915,N_1153,N_1442);
nand U1916 (N_1916,N_608,N_615);
nand U1917 (N_1917,N_1440,N_641);
or U1918 (N_1918,N_1398,N_586);
nand U1919 (N_1919,N_1334,N_184);
nand U1920 (N_1920,N_1075,N_1272);
nor U1921 (N_1921,N_1238,N_634);
nand U1922 (N_1922,N_35,N_412);
nor U1923 (N_1923,N_1279,N_1450);
nand U1924 (N_1924,N_965,N_828);
nor U1925 (N_1925,N_1305,N_343);
and U1926 (N_1926,N_1196,N_361);
nand U1927 (N_1927,N_1001,N_688);
nor U1928 (N_1928,N_884,N_1428);
nand U1929 (N_1929,N_632,N_91);
xnor U1930 (N_1930,N_401,N_1265);
nand U1931 (N_1931,N_1066,N_1273);
or U1932 (N_1932,N_375,N_1322);
nor U1933 (N_1933,N_1197,N_600);
xor U1934 (N_1934,N_1229,N_471);
and U1935 (N_1935,N_260,N_1468);
and U1936 (N_1936,N_1447,N_5);
xor U1937 (N_1937,N_1287,N_1064);
and U1938 (N_1938,N_211,N_126);
nand U1939 (N_1939,N_194,N_707);
nand U1940 (N_1940,N_138,N_1472);
or U1941 (N_1941,N_1393,N_1160);
or U1942 (N_1942,N_17,N_154);
nor U1943 (N_1943,N_509,N_954);
nand U1944 (N_1944,N_1325,N_1237);
and U1945 (N_1945,N_292,N_773);
xor U1946 (N_1946,N_324,N_14);
nor U1947 (N_1947,N_862,N_1331);
and U1948 (N_1948,N_1002,N_999);
nand U1949 (N_1949,N_429,N_1412);
nor U1950 (N_1950,N_883,N_498);
or U1951 (N_1951,N_1233,N_1278);
nand U1952 (N_1952,N_83,N_835);
nor U1953 (N_1953,N_769,N_1361);
or U1954 (N_1954,N_1126,N_409);
or U1955 (N_1955,N_938,N_258);
and U1956 (N_1956,N_780,N_1250);
xor U1957 (N_1957,N_76,N_102);
xor U1958 (N_1958,N_787,N_348);
and U1959 (N_1959,N_992,N_274);
nand U1960 (N_1960,N_1024,N_1371);
nand U1961 (N_1961,N_1438,N_657);
or U1962 (N_1962,N_1231,N_360);
nand U1963 (N_1963,N_1396,N_1013);
nand U1964 (N_1964,N_638,N_786);
nand U1965 (N_1965,N_330,N_628);
xnor U1966 (N_1966,N_744,N_419);
nor U1967 (N_1967,N_69,N_141);
nor U1968 (N_1968,N_1214,N_1475);
or U1969 (N_1969,N_761,N_1159);
xor U1970 (N_1970,N_640,N_1476);
nand U1971 (N_1971,N_417,N_248);
or U1972 (N_1972,N_382,N_888);
nand U1973 (N_1973,N_1251,N_552);
nand U1974 (N_1974,N_589,N_411);
and U1975 (N_1975,N_889,N_488);
or U1976 (N_1976,N_97,N_1120);
or U1977 (N_1977,N_1448,N_1288);
or U1978 (N_1978,N_173,N_172);
nor U1979 (N_1979,N_928,N_596);
or U1980 (N_1980,N_925,N_878);
nand U1981 (N_1981,N_745,N_1269);
and U1982 (N_1982,N_1357,N_164);
nor U1983 (N_1983,N_1083,N_1483);
and U1984 (N_1984,N_495,N_1111);
nor U1985 (N_1985,N_864,N_99);
and U1986 (N_1986,N_207,N_101);
or U1987 (N_1987,N_892,N_877);
nor U1988 (N_1988,N_1004,N_929);
nor U1989 (N_1989,N_566,N_529);
xor U1990 (N_1990,N_8,N_1326);
nor U1991 (N_1991,N_153,N_756);
and U1992 (N_1992,N_1086,N_238);
nor U1993 (N_1993,N_326,N_837);
and U1994 (N_1994,N_1015,N_374);
xor U1995 (N_1995,N_1067,N_555);
or U1996 (N_1996,N_119,N_1292);
and U1997 (N_1997,N_53,N_771);
or U1998 (N_1998,N_365,N_312);
or U1999 (N_1999,N_1429,N_706);
and U2000 (N_2000,N_1463,N_161);
and U2001 (N_2001,N_964,N_763);
and U2002 (N_2002,N_1056,N_1090);
nor U2003 (N_2003,N_1375,N_434);
xnor U2004 (N_2004,N_1323,N_367);
nor U2005 (N_2005,N_569,N_680);
xor U2006 (N_2006,N_200,N_667);
and U2007 (N_2007,N_549,N_303);
and U2008 (N_2008,N_1016,N_103);
or U2009 (N_2009,N_1073,N_185);
nor U2010 (N_2010,N_625,N_84);
or U2011 (N_2011,N_1123,N_48);
nor U2012 (N_2012,N_1007,N_1119);
nor U2013 (N_2013,N_1043,N_1236);
or U2014 (N_2014,N_1127,N_1037);
nor U2015 (N_2015,N_607,N_59);
nand U2016 (N_2016,N_951,N_368);
nor U2017 (N_2017,N_257,N_506);
nor U2018 (N_2018,N_967,N_352);
nand U2019 (N_2019,N_1246,N_1465);
nand U2020 (N_2020,N_1240,N_1025);
and U2021 (N_2021,N_612,N_107);
xnor U2022 (N_2022,N_263,N_846);
nor U2023 (N_2023,N_87,N_1058);
nor U2024 (N_2024,N_1049,N_222);
nand U2025 (N_2025,N_1320,N_675);
and U2026 (N_2026,N_320,N_805);
nand U2027 (N_2027,N_1270,N_868);
nor U2028 (N_2028,N_220,N_617);
nand U2029 (N_2029,N_665,N_956);
nand U2030 (N_2030,N_1142,N_345);
nand U2031 (N_2031,N_339,N_1207);
and U2032 (N_2032,N_322,N_198);
xor U2033 (N_2033,N_9,N_762);
and U2034 (N_2034,N_997,N_120);
or U2035 (N_2035,N_631,N_1186);
nor U2036 (N_2036,N_915,N_1099);
and U2037 (N_2037,N_256,N_961);
nor U2038 (N_2038,N_1146,N_941);
nand U2039 (N_2039,N_441,N_906);
and U2040 (N_2040,N_40,N_1307);
and U2041 (N_2041,N_534,N_18);
nand U2042 (N_2042,N_733,N_1498);
nor U2043 (N_2043,N_739,N_1124);
or U2044 (N_2044,N_853,N_575);
nand U2045 (N_2045,N_486,N_1195);
nor U2046 (N_2046,N_26,N_143);
nand U2047 (N_2047,N_1030,N_54);
nor U2048 (N_2048,N_1257,N_671);
nor U2049 (N_2049,N_551,N_228);
or U2050 (N_2050,N_1036,N_849);
or U2051 (N_2051,N_1312,N_1473);
nor U2052 (N_2052,N_684,N_1188);
and U2053 (N_2053,N_635,N_465);
nand U2054 (N_2054,N_1264,N_839);
xnor U2055 (N_2055,N_459,N_1494);
or U2056 (N_2056,N_687,N_876);
or U2057 (N_2057,N_806,N_259);
nand U2058 (N_2058,N_748,N_1430);
nor U2059 (N_2059,N_1190,N_975);
and U2060 (N_2060,N_500,N_1018);
or U2061 (N_2061,N_133,N_159);
nand U2062 (N_2062,N_543,N_268);
nor U2063 (N_2063,N_1045,N_30);
nor U2064 (N_2064,N_1390,N_12);
or U2065 (N_2065,N_1456,N_568);
and U2066 (N_2066,N_994,N_246);
and U2067 (N_2067,N_790,N_304);
or U2068 (N_2068,N_341,N_907);
nand U2069 (N_2069,N_620,N_1061);
and U2070 (N_2070,N_1137,N_229);
and U2071 (N_2071,N_299,N_966);
or U2072 (N_2072,N_836,N_691);
or U2073 (N_2073,N_1359,N_166);
and U2074 (N_2074,N_314,N_1000);
nand U2075 (N_2075,N_123,N_1169);
and U2076 (N_2076,N_1441,N_702);
or U2077 (N_2077,N_890,N_833);
nand U2078 (N_2078,N_45,N_1258);
nand U2079 (N_2079,N_252,N_1392);
xor U2080 (N_2080,N_283,N_831);
or U2081 (N_2081,N_55,N_916);
nand U2082 (N_2082,N_981,N_342);
and U2083 (N_2083,N_873,N_1491);
or U2084 (N_2084,N_516,N_819);
nand U2085 (N_2085,N_814,N_100);
and U2086 (N_2086,N_989,N_1260);
nor U2087 (N_2087,N_988,N_605);
nor U2088 (N_2088,N_1115,N_85);
or U2089 (N_2089,N_510,N_704);
or U2090 (N_2090,N_421,N_863);
nor U2091 (N_2091,N_852,N_571);
nand U2092 (N_2092,N_88,N_1209);
and U2093 (N_2093,N_310,N_296);
or U2094 (N_2094,N_1446,N_921);
and U2095 (N_2095,N_1219,N_960);
nor U2096 (N_2096,N_537,N_1178);
xnor U2097 (N_2097,N_333,N_1454);
nor U2098 (N_2098,N_262,N_610);
and U2099 (N_2099,N_130,N_1461);
or U2100 (N_2100,N_425,N_1087);
or U2101 (N_2101,N_712,N_73);
nand U2102 (N_2102,N_158,N_664);
or U2103 (N_2103,N_3,N_436);
nor U2104 (N_2104,N_1415,N_838);
nor U2105 (N_2105,N_1242,N_485);
nand U2106 (N_2106,N_1239,N_1202);
and U2107 (N_2107,N_1210,N_178);
and U2108 (N_2108,N_1327,N_832);
nand U2109 (N_2109,N_1034,N_140);
nand U2110 (N_2110,N_117,N_501);
and U2111 (N_2111,N_750,N_531);
xnor U2112 (N_2112,N_801,N_1114);
nand U2113 (N_2113,N_472,N_1397);
or U2114 (N_2114,N_93,N_1486);
or U2115 (N_2115,N_554,N_503);
and U2116 (N_2116,N_1404,N_479);
and U2117 (N_2117,N_794,N_455);
and U2118 (N_2118,N_79,N_650);
and U2119 (N_2119,N_598,N_430);
and U2120 (N_2120,N_1471,N_823);
nand U2121 (N_2121,N_908,N_1189);
nand U2122 (N_2122,N_948,N_223);
and U2123 (N_2123,N_1296,N_204);
and U2124 (N_2124,N_1497,N_337);
and U2125 (N_2125,N_834,N_1493);
and U2126 (N_2126,N_919,N_820);
xnor U2127 (N_2127,N_280,N_416);
or U2128 (N_2128,N_1057,N_1422);
or U2129 (N_2129,N_990,N_903);
nor U2130 (N_2130,N_670,N_804);
or U2131 (N_2131,N_545,N_1150);
or U2132 (N_2132,N_439,N_265);
or U2133 (N_2133,N_135,N_924);
nor U2134 (N_2134,N_438,N_1464);
or U2135 (N_2135,N_1140,N_208);
and U2136 (N_2136,N_866,N_1286);
or U2137 (N_2137,N_347,N_241);
nor U2138 (N_2138,N_654,N_170);
or U2139 (N_2139,N_947,N_1362);
nor U2140 (N_2140,N_729,N_308);
and U2141 (N_2141,N_62,N_799);
or U2142 (N_2142,N_611,N_1122);
or U2143 (N_2143,N_112,N_1271);
or U2144 (N_2144,N_524,N_1400);
nand U2145 (N_2145,N_1228,N_1281);
nor U2146 (N_2146,N_719,N_1344);
and U2147 (N_2147,N_116,N_428);
nand U2148 (N_2148,N_315,N_881);
and U2149 (N_2149,N_197,N_590);
nor U2150 (N_2150,N_34,N_306);
nor U2151 (N_2151,N_1008,N_213);
nand U2152 (N_2152,N_0,N_676);
and U2153 (N_2153,N_718,N_1383);
and U2154 (N_2154,N_802,N_1436);
nand U2155 (N_2155,N_493,N_1100);
nor U2156 (N_2156,N_885,N_1040);
xor U2157 (N_2157,N_96,N_249);
nand U2158 (N_2158,N_139,N_1157);
and U2159 (N_2159,N_334,N_1304);
nor U2160 (N_2160,N_276,N_1191);
and U2161 (N_2161,N_1193,N_386);
nor U2162 (N_2162,N_502,N_1070);
and U2163 (N_2163,N_577,N_816);
nand U2164 (N_2164,N_572,N_15);
nand U2165 (N_2165,N_1096,N_351);
nand U2166 (N_2166,N_1317,N_1205);
and U2167 (N_2167,N_896,N_354);
and U2168 (N_2168,N_288,N_1487);
or U2169 (N_2169,N_275,N_67);
or U2170 (N_2170,N_599,N_824);
or U2171 (N_2171,N_1409,N_1052);
and U2172 (N_2172,N_1282,N_25);
or U2173 (N_2173,N_716,N_755);
and U2174 (N_2174,N_380,N_1478);
and U2175 (N_2175,N_1431,N_1174);
nor U2176 (N_2176,N_227,N_935);
and U2177 (N_2177,N_1297,N_156);
or U2178 (N_2178,N_1443,N_254);
nand U2179 (N_2179,N_445,N_653);
and U2180 (N_2180,N_457,N_1225);
nand U2181 (N_2181,N_1401,N_847);
and U2182 (N_2182,N_51,N_21);
xor U2183 (N_2183,N_604,N_449);
xor U2184 (N_2184,N_922,N_1366);
and U2185 (N_2185,N_1139,N_942);
xor U2186 (N_2186,N_659,N_245);
and U2187 (N_2187,N_943,N_985);
or U2188 (N_2188,N_1060,N_513);
nand U2189 (N_2189,N_539,N_562);
nor U2190 (N_2190,N_880,N_350);
or U2191 (N_2191,N_1136,N_803);
and U2192 (N_2192,N_1263,N_713);
and U2193 (N_2193,N_872,N_1377);
or U2194 (N_2194,N_1254,N_955);
nor U2195 (N_2195,N_726,N_1213);
nor U2196 (N_2196,N_1332,N_132);
and U2197 (N_2197,N_775,N_1192);
nor U2198 (N_2198,N_56,N_328);
or U2199 (N_2199,N_1033,N_700);
or U2200 (N_2200,N_1223,N_446);
and U2201 (N_2201,N_1245,N_626);
or U2202 (N_2202,N_1029,N_788);
xor U2203 (N_2203,N_1167,N_648);
nand U2204 (N_2204,N_1104,N_1010);
nand U2205 (N_2205,N_618,N_747);
or U2206 (N_2206,N_842,N_725);
or U2207 (N_2207,N_467,N_821);
nand U2208 (N_2208,N_746,N_1313);
and U2209 (N_2209,N_60,N_818);
and U2210 (N_2210,N_800,N_171);
nor U2211 (N_2211,N_1046,N_1310);
xor U2212 (N_2212,N_28,N_886);
or U2213 (N_2213,N_458,N_24);
xor U2214 (N_2214,N_843,N_1247);
nand U2215 (N_2215,N_567,N_1022);
or U2216 (N_2216,N_75,N_250);
nor U2217 (N_2217,N_395,N_13);
or U2218 (N_2218,N_1341,N_1388);
nand U2219 (N_2219,N_879,N_244);
nand U2220 (N_2220,N_282,N_647);
and U2221 (N_2221,N_694,N_217);
and U2222 (N_2222,N_336,N_1348);
or U2223 (N_2223,N_301,N_808);
nor U2224 (N_2224,N_508,N_930);
nand U2225 (N_2225,N_1005,N_1434);
and U2226 (N_2226,N_730,N_977);
xor U2227 (N_2227,N_559,N_104);
or U2228 (N_2228,N_580,N_917);
or U2229 (N_2229,N_603,N_1457);
and U2230 (N_2230,N_1395,N_231);
nor U2231 (N_2231,N_591,N_456);
xnor U2232 (N_2232,N_1080,N_1234);
and U2233 (N_2233,N_708,N_759);
and U2234 (N_2234,N_1109,N_210);
nor U2235 (N_2235,N_779,N_1490);
and U2236 (N_2236,N_1019,N_714);
and U2237 (N_2237,N_1170,N_1047);
nor U2238 (N_2238,N_78,N_1363);
or U2239 (N_2239,N_349,N_736);
or U2240 (N_2240,N_1306,N_146);
xor U2241 (N_2241,N_1108,N_1222);
nand U2242 (N_2242,N_1414,N_144);
nor U2243 (N_2243,N_86,N_724);
nand U2244 (N_2244,N_633,N_1267);
and U2245 (N_2245,N_1462,N_557);
or U2246 (N_2246,N_236,N_147);
and U2247 (N_2247,N_1284,N_444);
and U2248 (N_2248,N_1329,N_1021);
nor U2249 (N_2249,N_52,N_1072);
and U2250 (N_2250,N_1314,N_1212);
nor U2251 (N_2251,N_1344,N_509);
and U2252 (N_2252,N_1179,N_577);
nor U2253 (N_2253,N_1067,N_601);
or U2254 (N_2254,N_869,N_1075);
nor U2255 (N_2255,N_472,N_1325);
nand U2256 (N_2256,N_806,N_252);
nand U2257 (N_2257,N_779,N_437);
or U2258 (N_2258,N_449,N_110);
nand U2259 (N_2259,N_837,N_1336);
or U2260 (N_2260,N_1145,N_1422);
nor U2261 (N_2261,N_1338,N_998);
nor U2262 (N_2262,N_160,N_1234);
xnor U2263 (N_2263,N_919,N_1099);
and U2264 (N_2264,N_477,N_1323);
and U2265 (N_2265,N_311,N_815);
nand U2266 (N_2266,N_81,N_1030);
nand U2267 (N_2267,N_340,N_791);
or U2268 (N_2268,N_634,N_1184);
and U2269 (N_2269,N_560,N_106);
or U2270 (N_2270,N_68,N_710);
or U2271 (N_2271,N_81,N_765);
and U2272 (N_2272,N_202,N_1178);
and U2273 (N_2273,N_1288,N_214);
or U2274 (N_2274,N_177,N_288);
xnor U2275 (N_2275,N_982,N_438);
and U2276 (N_2276,N_284,N_303);
and U2277 (N_2277,N_313,N_1383);
nor U2278 (N_2278,N_43,N_633);
and U2279 (N_2279,N_1029,N_141);
and U2280 (N_2280,N_1379,N_132);
nor U2281 (N_2281,N_593,N_26);
nor U2282 (N_2282,N_1284,N_1141);
or U2283 (N_2283,N_365,N_878);
nand U2284 (N_2284,N_1252,N_1129);
nor U2285 (N_2285,N_151,N_426);
and U2286 (N_2286,N_206,N_510);
or U2287 (N_2287,N_1156,N_1071);
xnor U2288 (N_2288,N_951,N_1479);
nand U2289 (N_2289,N_528,N_216);
nand U2290 (N_2290,N_244,N_272);
nor U2291 (N_2291,N_429,N_884);
nor U2292 (N_2292,N_1361,N_1095);
nor U2293 (N_2293,N_179,N_1132);
or U2294 (N_2294,N_467,N_323);
nor U2295 (N_2295,N_741,N_894);
nand U2296 (N_2296,N_90,N_211);
or U2297 (N_2297,N_329,N_1045);
xor U2298 (N_2298,N_535,N_492);
nand U2299 (N_2299,N_812,N_644);
and U2300 (N_2300,N_248,N_941);
xor U2301 (N_2301,N_28,N_320);
nand U2302 (N_2302,N_207,N_1001);
xnor U2303 (N_2303,N_75,N_135);
nor U2304 (N_2304,N_624,N_1156);
and U2305 (N_2305,N_1186,N_674);
nor U2306 (N_2306,N_460,N_972);
xor U2307 (N_2307,N_411,N_860);
nand U2308 (N_2308,N_1206,N_1244);
or U2309 (N_2309,N_1058,N_1497);
nor U2310 (N_2310,N_1477,N_192);
xnor U2311 (N_2311,N_1292,N_6);
nor U2312 (N_2312,N_818,N_887);
nor U2313 (N_2313,N_1418,N_1067);
and U2314 (N_2314,N_353,N_889);
nand U2315 (N_2315,N_476,N_1452);
and U2316 (N_2316,N_1214,N_1273);
nor U2317 (N_2317,N_34,N_1210);
xor U2318 (N_2318,N_728,N_303);
nand U2319 (N_2319,N_594,N_703);
nand U2320 (N_2320,N_578,N_1253);
nor U2321 (N_2321,N_28,N_1104);
nor U2322 (N_2322,N_1346,N_286);
nand U2323 (N_2323,N_49,N_452);
or U2324 (N_2324,N_536,N_21);
and U2325 (N_2325,N_822,N_1142);
nand U2326 (N_2326,N_41,N_1136);
nor U2327 (N_2327,N_1254,N_815);
nand U2328 (N_2328,N_585,N_726);
nor U2329 (N_2329,N_761,N_1290);
or U2330 (N_2330,N_7,N_1481);
and U2331 (N_2331,N_1048,N_1282);
or U2332 (N_2332,N_1404,N_498);
xnor U2333 (N_2333,N_72,N_321);
nor U2334 (N_2334,N_635,N_205);
nor U2335 (N_2335,N_668,N_1209);
or U2336 (N_2336,N_15,N_315);
nand U2337 (N_2337,N_292,N_1058);
nor U2338 (N_2338,N_1091,N_100);
or U2339 (N_2339,N_1291,N_1144);
and U2340 (N_2340,N_1267,N_802);
xnor U2341 (N_2341,N_121,N_1277);
nor U2342 (N_2342,N_1119,N_1359);
and U2343 (N_2343,N_1259,N_1357);
and U2344 (N_2344,N_366,N_28);
nor U2345 (N_2345,N_784,N_246);
or U2346 (N_2346,N_67,N_760);
nor U2347 (N_2347,N_515,N_306);
xor U2348 (N_2348,N_782,N_1049);
nand U2349 (N_2349,N_755,N_381);
or U2350 (N_2350,N_168,N_575);
nand U2351 (N_2351,N_633,N_69);
nor U2352 (N_2352,N_112,N_1334);
or U2353 (N_2353,N_1207,N_178);
or U2354 (N_2354,N_688,N_284);
nor U2355 (N_2355,N_89,N_308);
xnor U2356 (N_2356,N_529,N_835);
nand U2357 (N_2357,N_786,N_636);
xor U2358 (N_2358,N_1014,N_313);
nor U2359 (N_2359,N_816,N_943);
and U2360 (N_2360,N_134,N_1201);
nand U2361 (N_2361,N_1318,N_898);
nor U2362 (N_2362,N_143,N_1207);
or U2363 (N_2363,N_103,N_1477);
and U2364 (N_2364,N_981,N_327);
nand U2365 (N_2365,N_250,N_1022);
xnor U2366 (N_2366,N_473,N_586);
or U2367 (N_2367,N_441,N_1372);
nor U2368 (N_2368,N_1398,N_1343);
or U2369 (N_2369,N_278,N_480);
nor U2370 (N_2370,N_1345,N_35);
nor U2371 (N_2371,N_1222,N_1349);
and U2372 (N_2372,N_1175,N_622);
and U2373 (N_2373,N_1418,N_1112);
nor U2374 (N_2374,N_594,N_1236);
or U2375 (N_2375,N_851,N_27);
and U2376 (N_2376,N_1189,N_784);
nand U2377 (N_2377,N_1027,N_851);
nand U2378 (N_2378,N_1027,N_271);
and U2379 (N_2379,N_1396,N_375);
and U2380 (N_2380,N_240,N_1128);
nand U2381 (N_2381,N_546,N_332);
nor U2382 (N_2382,N_842,N_1079);
or U2383 (N_2383,N_1127,N_1373);
and U2384 (N_2384,N_668,N_1442);
nand U2385 (N_2385,N_212,N_1339);
nor U2386 (N_2386,N_1200,N_620);
xor U2387 (N_2387,N_668,N_2);
nand U2388 (N_2388,N_950,N_1110);
or U2389 (N_2389,N_170,N_448);
nand U2390 (N_2390,N_885,N_878);
or U2391 (N_2391,N_667,N_940);
and U2392 (N_2392,N_725,N_1307);
or U2393 (N_2393,N_1066,N_386);
and U2394 (N_2394,N_202,N_281);
nor U2395 (N_2395,N_155,N_1225);
nor U2396 (N_2396,N_200,N_937);
and U2397 (N_2397,N_825,N_310);
nand U2398 (N_2398,N_1203,N_978);
or U2399 (N_2399,N_151,N_1415);
xor U2400 (N_2400,N_916,N_381);
and U2401 (N_2401,N_404,N_1044);
and U2402 (N_2402,N_490,N_607);
or U2403 (N_2403,N_893,N_219);
nor U2404 (N_2404,N_1441,N_853);
and U2405 (N_2405,N_1446,N_495);
and U2406 (N_2406,N_928,N_366);
nor U2407 (N_2407,N_1062,N_356);
nand U2408 (N_2408,N_1063,N_1491);
nand U2409 (N_2409,N_1075,N_270);
and U2410 (N_2410,N_876,N_840);
or U2411 (N_2411,N_1295,N_619);
nor U2412 (N_2412,N_602,N_186);
xnor U2413 (N_2413,N_432,N_911);
or U2414 (N_2414,N_892,N_781);
nand U2415 (N_2415,N_477,N_263);
nor U2416 (N_2416,N_709,N_433);
nor U2417 (N_2417,N_59,N_510);
nand U2418 (N_2418,N_401,N_1254);
and U2419 (N_2419,N_1172,N_325);
or U2420 (N_2420,N_394,N_707);
nor U2421 (N_2421,N_734,N_398);
nand U2422 (N_2422,N_905,N_903);
nor U2423 (N_2423,N_606,N_757);
or U2424 (N_2424,N_1328,N_1104);
and U2425 (N_2425,N_878,N_1317);
or U2426 (N_2426,N_846,N_1390);
nand U2427 (N_2427,N_1423,N_102);
or U2428 (N_2428,N_471,N_1171);
nand U2429 (N_2429,N_789,N_126);
or U2430 (N_2430,N_90,N_213);
nand U2431 (N_2431,N_659,N_119);
xnor U2432 (N_2432,N_585,N_526);
nand U2433 (N_2433,N_977,N_1196);
and U2434 (N_2434,N_1395,N_99);
nor U2435 (N_2435,N_20,N_1299);
nor U2436 (N_2436,N_586,N_636);
and U2437 (N_2437,N_504,N_858);
and U2438 (N_2438,N_519,N_1101);
xnor U2439 (N_2439,N_811,N_578);
or U2440 (N_2440,N_1365,N_1229);
and U2441 (N_2441,N_1285,N_253);
nor U2442 (N_2442,N_1070,N_985);
nor U2443 (N_2443,N_1253,N_368);
nor U2444 (N_2444,N_1408,N_247);
nand U2445 (N_2445,N_148,N_531);
nor U2446 (N_2446,N_61,N_505);
and U2447 (N_2447,N_619,N_1382);
xnor U2448 (N_2448,N_708,N_57);
or U2449 (N_2449,N_1002,N_1109);
nand U2450 (N_2450,N_377,N_1177);
and U2451 (N_2451,N_62,N_733);
nor U2452 (N_2452,N_571,N_395);
and U2453 (N_2453,N_1090,N_92);
xnor U2454 (N_2454,N_1095,N_139);
nor U2455 (N_2455,N_1123,N_354);
nand U2456 (N_2456,N_274,N_723);
nor U2457 (N_2457,N_1471,N_1357);
and U2458 (N_2458,N_1419,N_29);
nand U2459 (N_2459,N_1098,N_1050);
or U2460 (N_2460,N_420,N_167);
and U2461 (N_2461,N_1051,N_1222);
nand U2462 (N_2462,N_1187,N_811);
or U2463 (N_2463,N_761,N_1339);
xor U2464 (N_2464,N_1485,N_259);
nor U2465 (N_2465,N_391,N_318);
xnor U2466 (N_2466,N_1059,N_486);
and U2467 (N_2467,N_413,N_391);
nor U2468 (N_2468,N_487,N_1404);
and U2469 (N_2469,N_15,N_553);
nand U2470 (N_2470,N_297,N_282);
or U2471 (N_2471,N_573,N_1103);
and U2472 (N_2472,N_532,N_1203);
or U2473 (N_2473,N_776,N_1495);
nand U2474 (N_2474,N_435,N_46);
or U2475 (N_2475,N_701,N_44);
nor U2476 (N_2476,N_403,N_28);
or U2477 (N_2477,N_1139,N_950);
nor U2478 (N_2478,N_1106,N_783);
nor U2479 (N_2479,N_765,N_1119);
nand U2480 (N_2480,N_759,N_672);
xnor U2481 (N_2481,N_475,N_891);
and U2482 (N_2482,N_772,N_851);
nor U2483 (N_2483,N_859,N_231);
nand U2484 (N_2484,N_19,N_1270);
nor U2485 (N_2485,N_347,N_337);
nand U2486 (N_2486,N_1216,N_978);
nand U2487 (N_2487,N_1413,N_395);
or U2488 (N_2488,N_833,N_820);
and U2489 (N_2489,N_1048,N_102);
or U2490 (N_2490,N_1336,N_1288);
and U2491 (N_2491,N_807,N_814);
or U2492 (N_2492,N_202,N_442);
and U2493 (N_2493,N_1240,N_489);
and U2494 (N_2494,N_968,N_1367);
nand U2495 (N_2495,N_355,N_1065);
or U2496 (N_2496,N_720,N_1482);
nor U2497 (N_2497,N_1171,N_1213);
nand U2498 (N_2498,N_161,N_1215);
and U2499 (N_2499,N_116,N_135);
nor U2500 (N_2500,N_1347,N_807);
or U2501 (N_2501,N_1486,N_773);
nand U2502 (N_2502,N_1197,N_926);
nand U2503 (N_2503,N_456,N_709);
nand U2504 (N_2504,N_1306,N_1243);
or U2505 (N_2505,N_1172,N_1462);
or U2506 (N_2506,N_939,N_850);
nand U2507 (N_2507,N_1235,N_537);
or U2508 (N_2508,N_1164,N_402);
and U2509 (N_2509,N_432,N_243);
nand U2510 (N_2510,N_1490,N_1469);
nor U2511 (N_2511,N_742,N_253);
and U2512 (N_2512,N_1014,N_896);
nor U2513 (N_2513,N_423,N_1450);
or U2514 (N_2514,N_1373,N_584);
and U2515 (N_2515,N_324,N_1246);
and U2516 (N_2516,N_220,N_1385);
nand U2517 (N_2517,N_542,N_789);
nand U2518 (N_2518,N_1201,N_1495);
or U2519 (N_2519,N_668,N_429);
xor U2520 (N_2520,N_901,N_785);
nand U2521 (N_2521,N_916,N_1310);
or U2522 (N_2522,N_877,N_1217);
nor U2523 (N_2523,N_390,N_127);
nand U2524 (N_2524,N_1042,N_382);
nand U2525 (N_2525,N_1016,N_1435);
nand U2526 (N_2526,N_743,N_493);
nand U2527 (N_2527,N_1423,N_366);
xor U2528 (N_2528,N_429,N_823);
and U2529 (N_2529,N_661,N_33);
nor U2530 (N_2530,N_123,N_990);
and U2531 (N_2531,N_478,N_1062);
and U2532 (N_2532,N_909,N_366);
nand U2533 (N_2533,N_288,N_872);
and U2534 (N_2534,N_1237,N_74);
nor U2535 (N_2535,N_757,N_590);
or U2536 (N_2536,N_1384,N_1154);
nor U2537 (N_2537,N_620,N_222);
nor U2538 (N_2538,N_282,N_105);
and U2539 (N_2539,N_13,N_500);
nand U2540 (N_2540,N_924,N_130);
or U2541 (N_2541,N_911,N_945);
nand U2542 (N_2542,N_237,N_859);
xnor U2543 (N_2543,N_1185,N_191);
nand U2544 (N_2544,N_1039,N_66);
nand U2545 (N_2545,N_44,N_458);
and U2546 (N_2546,N_804,N_85);
xnor U2547 (N_2547,N_613,N_285);
nand U2548 (N_2548,N_596,N_535);
or U2549 (N_2549,N_1017,N_961);
and U2550 (N_2550,N_780,N_903);
nand U2551 (N_2551,N_636,N_1086);
nand U2552 (N_2552,N_241,N_200);
nand U2553 (N_2553,N_445,N_727);
nor U2554 (N_2554,N_9,N_1019);
and U2555 (N_2555,N_929,N_186);
nor U2556 (N_2556,N_380,N_899);
or U2557 (N_2557,N_325,N_646);
nor U2558 (N_2558,N_605,N_550);
nor U2559 (N_2559,N_815,N_543);
or U2560 (N_2560,N_337,N_1495);
and U2561 (N_2561,N_368,N_215);
xor U2562 (N_2562,N_1321,N_960);
or U2563 (N_2563,N_1204,N_1002);
and U2564 (N_2564,N_1023,N_1028);
xnor U2565 (N_2565,N_1100,N_226);
and U2566 (N_2566,N_843,N_1407);
or U2567 (N_2567,N_520,N_1319);
xor U2568 (N_2568,N_556,N_407);
and U2569 (N_2569,N_406,N_783);
nor U2570 (N_2570,N_895,N_1490);
or U2571 (N_2571,N_766,N_1237);
and U2572 (N_2572,N_605,N_1194);
nor U2573 (N_2573,N_1202,N_1172);
or U2574 (N_2574,N_746,N_21);
nor U2575 (N_2575,N_851,N_1373);
and U2576 (N_2576,N_17,N_177);
or U2577 (N_2577,N_175,N_701);
nand U2578 (N_2578,N_382,N_159);
and U2579 (N_2579,N_1379,N_752);
nor U2580 (N_2580,N_951,N_493);
nand U2581 (N_2581,N_413,N_1063);
nor U2582 (N_2582,N_633,N_534);
and U2583 (N_2583,N_555,N_1364);
xnor U2584 (N_2584,N_1463,N_781);
and U2585 (N_2585,N_496,N_255);
and U2586 (N_2586,N_704,N_537);
nand U2587 (N_2587,N_1463,N_1272);
or U2588 (N_2588,N_1379,N_1216);
nand U2589 (N_2589,N_46,N_467);
nand U2590 (N_2590,N_720,N_610);
nor U2591 (N_2591,N_940,N_1424);
and U2592 (N_2592,N_1160,N_65);
and U2593 (N_2593,N_1012,N_897);
or U2594 (N_2594,N_299,N_282);
and U2595 (N_2595,N_621,N_863);
and U2596 (N_2596,N_876,N_1326);
nand U2597 (N_2597,N_88,N_1314);
xnor U2598 (N_2598,N_112,N_1131);
or U2599 (N_2599,N_1006,N_490);
or U2600 (N_2600,N_1114,N_480);
nand U2601 (N_2601,N_1192,N_266);
nand U2602 (N_2602,N_1209,N_1203);
or U2603 (N_2603,N_734,N_322);
or U2604 (N_2604,N_926,N_1203);
nand U2605 (N_2605,N_1235,N_1381);
or U2606 (N_2606,N_1229,N_933);
and U2607 (N_2607,N_549,N_72);
nor U2608 (N_2608,N_40,N_993);
or U2609 (N_2609,N_443,N_521);
or U2610 (N_2610,N_1066,N_632);
xnor U2611 (N_2611,N_775,N_123);
or U2612 (N_2612,N_972,N_336);
or U2613 (N_2613,N_1128,N_1266);
nor U2614 (N_2614,N_445,N_666);
nand U2615 (N_2615,N_207,N_701);
nor U2616 (N_2616,N_414,N_374);
nor U2617 (N_2617,N_251,N_109);
nor U2618 (N_2618,N_1215,N_601);
nor U2619 (N_2619,N_1232,N_1125);
nor U2620 (N_2620,N_714,N_1366);
or U2621 (N_2621,N_358,N_248);
nor U2622 (N_2622,N_976,N_65);
nand U2623 (N_2623,N_236,N_146);
xor U2624 (N_2624,N_465,N_105);
or U2625 (N_2625,N_860,N_424);
and U2626 (N_2626,N_259,N_967);
nor U2627 (N_2627,N_48,N_391);
or U2628 (N_2628,N_36,N_771);
or U2629 (N_2629,N_334,N_447);
nor U2630 (N_2630,N_1426,N_797);
or U2631 (N_2631,N_1422,N_194);
or U2632 (N_2632,N_458,N_1097);
xor U2633 (N_2633,N_387,N_972);
xor U2634 (N_2634,N_1298,N_1012);
nand U2635 (N_2635,N_381,N_29);
xnor U2636 (N_2636,N_426,N_844);
and U2637 (N_2637,N_1135,N_764);
or U2638 (N_2638,N_870,N_1073);
or U2639 (N_2639,N_472,N_378);
or U2640 (N_2640,N_927,N_1296);
nor U2641 (N_2641,N_1411,N_1478);
or U2642 (N_2642,N_107,N_832);
nand U2643 (N_2643,N_262,N_777);
nand U2644 (N_2644,N_264,N_581);
or U2645 (N_2645,N_680,N_190);
or U2646 (N_2646,N_683,N_283);
nand U2647 (N_2647,N_107,N_1012);
and U2648 (N_2648,N_346,N_418);
or U2649 (N_2649,N_1198,N_52);
nor U2650 (N_2650,N_140,N_40);
nor U2651 (N_2651,N_961,N_281);
xnor U2652 (N_2652,N_1493,N_362);
nor U2653 (N_2653,N_69,N_985);
or U2654 (N_2654,N_71,N_820);
nand U2655 (N_2655,N_256,N_365);
nor U2656 (N_2656,N_980,N_919);
nand U2657 (N_2657,N_366,N_286);
nand U2658 (N_2658,N_751,N_500);
xor U2659 (N_2659,N_1029,N_119);
nand U2660 (N_2660,N_164,N_305);
xnor U2661 (N_2661,N_1030,N_141);
nor U2662 (N_2662,N_753,N_956);
nor U2663 (N_2663,N_1060,N_86);
nand U2664 (N_2664,N_342,N_912);
nor U2665 (N_2665,N_348,N_273);
xnor U2666 (N_2666,N_19,N_1214);
nor U2667 (N_2667,N_415,N_1226);
nand U2668 (N_2668,N_788,N_801);
or U2669 (N_2669,N_190,N_1048);
nand U2670 (N_2670,N_1230,N_658);
or U2671 (N_2671,N_104,N_1380);
and U2672 (N_2672,N_417,N_1365);
nand U2673 (N_2673,N_307,N_225);
nand U2674 (N_2674,N_899,N_86);
nand U2675 (N_2675,N_1050,N_648);
or U2676 (N_2676,N_131,N_1003);
and U2677 (N_2677,N_200,N_1339);
or U2678 (N_2678,N_1239,N_248);
nand U2679 (N_2679,N_770,N_355);
nor U2680 (N_2680,N_1279,N_391);
nor U2681 (N_2681,N_376,N_938);
xor U2682 (N_2682,N_1135,N_460);
nor U2683 (N_2683,N_1356,N_212);
nand U2684 (N_2684,N_601,N_273);
nor U2685 (N_2685,N_1008,N_611);
xnor U2686 (N_2686,N_1346,N_452);
or U2687 (N_2687,N_980,N_1398);
or U2688 (N_2688,N_1218,N_97);
and U2689 (N_2689,N_1029,N_1004);
xnor U2690 (N_2690,N_140,N_1413);
nor U2691 (N_2691,N_1285,N_1200);
nand U2692 (N_2692,N_587,N_689);
nor U2693 (N_2693,N_1404,N_1275);
nor U2694 (N_2694,N_81,N_18);
and U2695 (N_2695,N_865,N_783);
and U2696 (N_2696,N_364,N_1256);
and U2697 (N_2697,N_1074,N_1448);
and U2698 (N_2698,N_1288,N_1321);
nand U2699 (N_2699,N_1287,N_812);
nor U2700 (N_2700,N_315,N_596);
nand U2701 (N_2701,N_660,N_451);
xor U2702 (N_2702,N_1174,N_310);
nand U2703 (N_2703,N_809,N_905);
nand U2704 (N_2704,N_62,N_492);
xnor U2705 (N_2705,N_560,N_802);
and U2706 (N_2706,N_1374,N_219);
xnor U2707 (N_2707,N_1305,N_974);
nand U2708 (N_2708,N_990,N_1104);
nand U2709 (N_2709,N_1145,N_783);
or U2710 (N_2710,N_1463,N_626);
nand U2711 (N_2711,N_986,N_712);
and U2712 (N_2712,N_992,N_1021);
nor U2713 (N_2713,N_336,N_992);
and U2714 (N_2714,N_1343,N_1087);
nor U2715 (N_2715,N_196,N_371);
nand U2716 (N_2716,N_1007,N_414);
or U2717 (N_2717,N_1370,N_1053);
nor U2718 (N_2718,N_146,N_631);
or U2719 (N_2719,N_559,N_1175);
nor U2720 (N_2720,N_988,N_122);
nor U2721 (N_2721,N_1263,N_525);
and U2722 (N_2722,N_1068,N_401);
nor U2723 (N_2723,N_1230,N_1118);
nor U2724 (N_2724,N_998,N_777);
and U2725 (N_2725,N_760,N_730);
xor U2726 (N_2726,N_1242,N_341);
or U2727 (N_2727,N_107,N_303);
nand U2728 (N_2728,N_1112,N_865);
xor U2729 (N_2729,N_488,N_849);
and U2730 (N_2730,N_1404,N_797);
and U2731 (N_2731,N_411,N_664);
xnor U2732 (N_2732,N_1224,N_15);
nor U2733 (N_2733,N_1219,N_1155);
and U2734 (N_2734,N_866,N_782);
nand U2735 (N_2735,N_97,N_616);
and U2736 (N_2736,N_426,N_1122);
or U2737 (N_2737,N_1230,N_1299);
nand U2738 (N_2738,N_112,N_849);
or U2739 (N_2739,N_392,N_199);
nor U2740 (N_2740,N_1003,N_772);
or U2741 (N_2741,N_1121,N_291);
and U2742 (N_2742,N_1247,N_336);
nor U2743 (N_2743,N_194,N_746);
nor U2744 (N_2744,N_945,N_1096);
or U2745 (N_2745,N_1047,N_793);
nand U2746 (N_2746,N_1224,N_1168);
xnor U2747 (N_2747,N_674,N_550);
and U2748 (N_2748,N_167,N_206);
and U2749 (N_2749,N_346,N_1328);
or U2750 (N_2750,N_5,N_699);
and U2751 (N_2751,N_126,N_659);
nor U2752 (N_2752,N_1438,N_169);
and U2753 (N_2753,N_1320,N_1062);
xor U2754 (N_2754,N_868,N_314);
xor U2755 (N_2755,N_223,N_1491);
xnor U2756 (N_2756,N_1471,N_759);
or U2757 (N_2757,N_1124,N_452);
and U2758 (N_2758,N_1331,N_1332);
nor U2759 (N_2759,N_881,N_471);
or U2760 (N_2760,N_602,N_1409);
and U2761 (N_2761,N_892,N_695);
xor U2762 (N_2762,N_1049,N_1367);
or U2763 (N_2763,N_1309,N_395);
nand U2764 (N_2764,N_1037,N_370);
or U2765 (N_2765,N_1294,N_843);
and U2766 (N_2766,N_598,N_709);
or U2767 (N_2767,N_36,N_333);
nand U2768 (N_2768,N_711,N_674);
nand U2769 (N_2769,N_1191,N_1327);
or U2770 (N_2770,N_1402,N_1266);
nand U2771 (N_2771,N_340,N_483);
and U2772 (N_2772,N_1492,N_1465);
nor U2773 (N_2773,N_643,N_58);
or U2774 (N_2774,N_1259,N_675);
or U2775 (N_2775,N_379,N_344);
and U2776 (N_2776,N_578,N_1377);
nand U2777 (N_2777,N_1490,N_880);
nand U2778 (N_2778,N_441,N_740);
and U2779 (N_2779,N_490,N_520);
xor U2780 (N_2780,N_1301,N_703);
or U2781 (N_2781,N_359,N_71);
or U2782 (N_2782,N_726,N_10);
nor U2783 (N_2783,N_397,N_793);
and U2784 (N_2784,N_1252,N_258);
nand U2785 (N_2785,N_123,N_61);
nand U2786 (N_2786,N_1321,N_1474);
or U2787 (N_2787,N_311,N_462);
and U2788 (N_2788,N_378,N_429);
nand U2789 (N_2789,N_601,N_1161);
nor U2790 (N_2790,N_446,N_853);
nand U2791 (N_2791,N_654,N_546);
nor U2792 (N_2792,N_920,N_1318);
or U2793 (N_2793,N_981,N_662);
xnor U2794 (N_2794,N_1031,N_698);
or U2795 (N_2795,N_1049,N_829);
nor U2796 (N_2796,N_963,N_111);
nor U2797 (N_2797,N_1405,N_1237);
xnor U2798 (N_2798,N_1232,N_1113);
nor U2799 (N_2799,N_987,N_284);
nor U2800 (N_2800,N_107,N_713);
or U2801 (N_2801,N_980,N_1051);
nor U2802 (N_2802,N_568,N_922);
nor U2803 (N_2803,N_1309,N_1422);
or U2804 (N_2804,N_710,N_817);
xnor U2805 (N_2805,N_837,N_999);
or U2806 (N_2806,N_1154,N_872);
or U2807 (N_2807,N_1494,N_891);
or U2808 (N_2808,N_426,N_1410);
or U2809 (N_2809,N_530,N_587);
or U2810 (N_2810,N_115,N_181);
and U2811 (N_2811,N_377,N_78);
xor U2812 (N_2812,N_949,N_687);
xnor U2813 (N_2813,N_984,N_1128);
and U2814 (N_2814,N_574,N_446);
and U2815 (N_2815,N_922,N_1244);
nor U2816 (N_2816,N_302,N_700);
or U2817 (N_2817,N_49,N_155);
and U2818 (N_2818,N_640,N_886);
nand U2819 (N_2819,N_1291,N_429);
nand U2820 (N_2820,N_514,N_36);
or U2821 (N_2821,N_1111,N_424);
and U2822 (N_2822,N_1419,N_656);
nor U2823 (N_2823,N_225,N_1399);
and U2824 (N_2824,N_462,N_41);
nor U2825 (N_2825,N_768,N_324);
and U2826 (N_2826,N_580,N_1362);
nand U2827 (N_2827,N_1357,N_245);
nor U2828 (N_2828,N_1077,N_996);
xor U2829 (N_2829,N_1226,N_848);
or U2830 (N_2830,N_1002,N_806);
nor U2831 (N_2831,N_120,N_916);
and U2832 (N_2832,N_760,N_1481);
or U2833 (N_2833,N_125,N_367);
nand U2834 (N_2834,N_945,N_863);
or U2835 (N_2835,N_1338,N_1325);
nand U2836 (N_2836,N_867,N_16);
nor U2837 (N_2837,N_1433,N_173);
nand U2838 (N_2838,N_773,N_525);
nand U2839 (N_2839,N_792,N_1178);
or U2840 (N_2840,N_7,N_1014);
or U2841 (N_2841,N_43,N_58);
nor U2842 (N_2842,N_596,N_559);
nor U2843 (N_2843,N_1417,N_3);
and U2844 (N_2844,N_1115,N_1379);
and U2845 (N_2845,N_1330,N_807);
xnor U2846 (N_2846,N_185,N_809);
or U2847 (N_2847,N_996,N_748);
nor U2848 (N_2848,N_674,N_546);
nand U2849 (N_2849,N_461,N_1366);
nor U2850 (N_2850,N_663,N_707);
or U2851 (N_2851,N_609,N_1374);
or U2852 (N_2852,N_676,N_759);
nor U2853 (N_2853,N_522,N_406);
or U2854 (N_2854,N_552,N_1388);
nand U2855 (N_2855,N_363,N_1251);
and U2856 (N_2856,N_1243,N_714);
nand U2857 (N_2857,N_503,N_1407);
nand U2858 (N_2858,N_613,N_969);
or U2859 (N_2859,N_757,N_158);
nand U2860 (N_2860,N_1236,N_1305);
or U2861 (N_2861,N_828,N_519);
and U2862 (N_2862,N_473,N_658);
xnor U2863 (N_2863,N_190,N_1424);
and U2864 (N_2864,N_1275,N_1388);
or U2865 (N_2865,N_1179,N_557);
and U2866 (N_2866,N_557,N_554);
xnor U2867 (N_2867,N_227,N_245);
and U2868 (N_2868,N_960,N_1298);
and U2869 (N_2869,N_261,N_234);
nand U2870 (N_2870,N_1499,N_868);
or U2871 (N_2871,N_259,N_489);
and U2872 (N_2872,N_267,N_1499);
and U2873 (N_2873,N_1275,N_160);
and U2874 (N_2874,N_595,N_417);
nor U2875 (N_2875,N_964,N_46);
xnor U2876 (N_2876,N_47,N_313);
nor U2877 (N_2877,N_774,N_186);
and U2878 (N_2878,N_1375,N_356);
and U2879 (N_2879,N_989,N_82);
and U2880 (N_2880,N_798,N_1095);
or U2881 (N_2881,N_436,N_1390);
nand U2882 (N_2882,N_1073,N_1120);
nor U2883 (N_2883,N_125,N_236);
nand U2884 (N_2884,N_437,N_497);
and U2885 (N_2885,N_548,N_149);
or U2886 (N_2886,N_855,N_422);
or U2887 (N_2887,N_23,N_1385);
nand U2888 (N_2888,N_335,N_910);
nor U2889 (N_2889,N_167,N_562);
nor U2890 (N_2890,N_358,N_498);
nor U2891 (N_2891,N_1179,N_502);
and U2892 (N_2892,N_574,N_773);
or U2893 (N_2893,N_357,N_1188);
nor U2894 (N_2894,N_1075,N_836);
nor U2895 (N_2895,N_747,N_203);
and U2896 (N_2896,N_265,N_21);
nand U2897 (N_2897,N_353,N_209);
xnor U2898 (N_2898,N_1459,N_546);
nand U2899 (N_2899,N_786,N_513);
nor U2900 (N_2900,N_642,N_469);
nand U2901 (N_2901,N_703,N_261);
or U2902 (N_2902,N_998,N_1446);
nor U2903 (N_2903,N_562,N_1104);
nand U2904 (N_2904,N_1183,N_810);
nand U2905 (N_2905,N_675,N_444);
nand U2906 (N_2906,N_732,N_1416);
or U2907 (N_2907,N_1177,N_521);
and U2908 (N_2908,N_348,N_555);
or U2909 (N_2909,N_641,N_184);
nor U2910 (N_2910,N_1126,N_872);
nor U2911 (N_2911,N_478,N_656);
nand U2912 (N_2912,N_95,N_1167);
xnor U2913 (N_2913,N_258,N_353);
or U2914 (N_2914,N_713,N_750);
and U2915 (N_2915,N_804,N_717);
nand U2916 (N_2916,N_962,N_270);
nor U2917 (N_2917,N_615,N_410);
nand U2918 (N_2918,N_701,N_1273);
nand U2919 (N_2919,N_768,N_922);
and U2920 (N_2920,N_723,N_1405);
or U2921 (N_2921,N_477,N_959);
xnor U2922 (N_2922,N_1034,N_1136);
nor U2923 (N_2923,N_1317,N_99);
xor U2924 (N_2924,N_1373,N_274);
or U2925 (N_2925,N_498,N_622);
and U2926 (N_2926,N_1248,N_1041);
and U2927 (N_2927,N_1385,N_1028);
xor U2928 (N_2928,N_497,N_1141);
nor U2929 (N_2929,N_1242,N_131);
nor U2930 (N_2930,N_995,N_311);
and U2931 (N_2931,N_974,N_1373);
and U2932 (N_2932,N_1360,N_1420);
or U2933 (N_2933,N_745,N_403);
or U2934 (N_2934,N_847,N_699);
nor U2935 (N_2935,N_424,N_230);
nor U2936 (N_2936,N_559,N_622);
and U2937 (N_2937,N_1450,N_727);
nand U2938 (N_2938,N_941,N_983);
or U2939 (N_2939,N_312,N_1069);
and U2940 (N_2940,N_1412,N_166);
or U2941 (N_2941,N_749,N_659);
or U2942 (N_2942,N_1288,N_269);
nand U2943 (N_2943,N_1013,N_1447);
or U2944 (N_2944,N_189,N_1346);
xnor U2945 (N_2945,N_727,N_1078);
and U2946 (N_2946,N_204,N_1434);
nand U2947 (N_2947,N_409,N_623);
nand U2948 (N_2948,N_588,N_494);
or U2949 (N_2949,N_1385,N_91);
nand U2950 (N_2950,N_570,N_929);
nand U2951 (N_2951,N_410,N_1377);
nor U2952 (N_2952,N_702,N_359);
or U2953 (N_2953,N_1052,N_769);
nor U2954 (N_2954,N_405,N_1062);
and U2955 (N_2955,N_1027,N_1299);
or U2956 (N_2956,N_216,N_1378);
or U2957 (N_2957,N_321,N_1180);
nand U2958 (N_2958,N_1212,N_511);
nand U2959 (N_2959,N_621,N_1429);
and U2960 (N_2960,N_1085,N_763);
nand U2961 (N_2961,N_1352,N_1493);
or U2962 (N_2962,N_380,N_1015);
and U2963 (N_2963,N_1143,N_277);
nor U2964 (N_2964,N_1438,N_1094);
or U2965 (N_2965,N_792,N_858);
and U2966 (N_2966,N_1233,N_47);
or U2967 (N_2967,N_1453,N_150);
nand U2968 (N_2968,N_962,N_1073);
and U2969 (N_2969,N_1010,N_633);
or U2970 (N_2970,N_1276,N_379);
or U2971 (N_2971,N_115,N_1218);
nand U2972 (N_2972,N_787,N_1006);
xnor U2973 (N_2973,N_82,N_47);
and U2974 (N_2974,N_1291,N_42);
xor U2975 (N_2975,N_207,N_808);
nand U2976 (N_2976,N_920,N_501);
and U2977 (N_2977,N_1130,N_840);
nand U2978 (N_2978,N_591,N_669);
xnor U2979 (N_2979,N_752,N_425);
nand U2980 (N_2980,N_158,N_348);
nor U2981 (N_2981,N_299,N_796);
or U2982 (N_2982,N_404,N_930);
xnor U2983 (N_2983,N_46,N_935);
nor U2984 (N_2984,N_168,N_422);
and U2985 (N_2985,N_122,N_1465);
xor U2986 (N_2986,N_1189,N_791);
nand U2987 (N_2987,N_1,N_39);
xnor U2988 (N_2988,N_35,N_1079);
or U2989 (N_2989,N_416,N_1004);
xnor U2990 (N_2990,N_81,N_133);
or U2991 (N_2991,N_1253,N_721);
nand U2992 (N_2992,N_224,N_1159);
or U2993 (N_2993,N_730,N_610);
or U2994 (N_2994,N_924,N_730);
nor U2995 (N_2995,N_612,N_980);
nand U2996 (N_2996,N_327,N_828);
nand U2997 (N_2997,N_935,N_1258);
nand U2998 (N_2998,N_604,N_107);
or U2999 (N_2999,N_1329,N_427);
or U3000 (N_3000,N_1763,N_2445);
or U3001 (N_3001,N_2868,N_1739);
xor U3002 (N_3002,N_2751,N_2558);
and U3003 (N_3003,N_1578,N_2974);
and U3004 (N_3004,N_2297,N_1889);
or U3005 (N_3005,N_1841,N_2225);
and U3006 (N_3006,N_1667,N_1997);
nand U3007 (N_3007,N_2412,N_2264);
and U3008 (N_3008,N_2941,N_2118);
or U3009 (N_3009,N_1781,N_2496);
or U3010 (N_3010,N_1757,N_2083);
and U3011 (N_3011,N_1947,N_1777);
and U3012 (N_3012,N_1555,N_1719);
or U3013 (N_3013,N_1731,N_2074);
and U3014 (N_3014,N_2457,N_2367);
nor U3015 (N_3015,N_2382,N_2882);
xnor U3016 (N_3016,N_1536,N_1671);
nor U3017 (N_3017,N_2652,N_2580);
xor U3018 (N_3018,N_1694,N_1756);
nor U3019 (N_3019,N_1675,N_1620);
and U3020 (N_3020,N_1524,N_1635);
and U3021 (N_3021,N_1581,N_1506);
nand U3022 (N_3022,N_1897,N_2198);
nor U3023 (N_3023,N_2324,N_1571);
nand U3024 (N_3024,N_2420,N_2177);
nor U3025 (N_3025,N_2998,N_2244);
or U3026 (N_3026,N_2869,N_2912);
or U3027 (N_3027,N_2044,N_1604);
nor U3028 (N_3028,N_2042,N_2729);
and U3029 (N_3029,N_1552,N_1655);
or U3030 (N_3030,N_2062,N_1874);
and U3031 (N_3031,N_1627,N_2229);
nand U3032 (N_3032,N_1669,N_1676);
and U3033 (N_3033,N_2022,N_2502);
nand U3034 (N_3034,N_2529,N_2208);
xor U3035 (N_3035,N_2184,N_2035);
and U3036 (N_3036,N_2576,N_1726);
nand U3037 (N_3037,N_2907,N_2833);
or U3038 (N_3038,N_1745,N_2484);
or U3039 (N_3039,N_2671,N_1804);
nor U3040 (N_3040,N_2552,N_2607);
nand U3041 (N_3041,N_2474,N_2028);
and U3042 (N_3042,N_2634,N_1556);
xor U3043 (N_3043,N_1780,N_2845);
nor U3044 (N_3044,N_2122,N_1943);
nand U3045 (N_3045,N_2435,N_2589);
or U3046 (N_3046,N_1785,N_2338);
and U3047 (N_3047,N_2767,N_2128);
nor U3048 (N_3048,N_1570,N_2973);
nand U3049 (N_3049,N_2965,N_2906);
nand U3050 (N_3050,N_2064,N_1815);
nor U3051 (N_3051,N_2525,N_2646);
nand U3052 (N_3052,N_2187,N_1853);
nor U3053 (N_3053,N_1911,N_2095);
nand U3054 (N_3054,N_1992,N_2760);
or U3055 (N_3055,N_1658,N_1964);
and U3056 (N_3056,N_2395,N_1686);
xnor U3057 (N_3057,N_1865,N_2599);
and U3058 (N_3058,N_1799,N_2790);
and U3059 (N_3059,N_2109,N_1925);
and U3060 (N_3060,N_2391,N_1843);
or U3061 (N_3061,N_1639,N_1586);
and U3062 (N_3062,N_2571,N_1946);
and U3063 (N_3063,N_2092,N_2458);
xor U3064 (N_3064,N_2014,N_1940);
and U3065 (N_3065,N_2460,N_2000);
xnor U3066 (N_3066,N_2029,N_2934);
xnor U3067 (N_3067,N_2428,N_1542);
xor U3068 (N_3068,N_1910,N_2079);
nand U3069 (N_3069,N_2712,N_2718);
and U3070 (N_3070,N_1835,N_2146);
or U3071 (N_3071,N_2066,N_2213);
nor U3072 (N_3072,N_2050,N_2344);
nand U3073 (N_3073,N_2449,N_2057);
nand U3074 (N_3074,N_2308,N_2535);
nand U3075 (N_3075,N_2768,N_2656);
nand U3076 (N_3076,N_1993,N_2590);
and U3077 (N_3077,N_2037,N_2695);
nor U3078 (N_3078,N_2158,N_2688);
or U3079 (N_3079,N_1613,N_2415);
xnor U3080 (N_3080,N_2844,N_1965);
nand U3081 (N_3081,N_2299,N_2280);
nor U3082 (N_3082,N_2155,N_2997);
nor U3083 (N_3083,N_2903,N_2045);
nand U3084 (N_3084,N_2181,N_1858);
nor U3085 (N_3085,N_1568,N_2740);
nor U3086 (N_3086,N_2834,N_2808);
or U3087 (N_3087,N_1605,N_1818);
nor U3088 (N_3088,N_1806,N_2026);
nand U3089 (N_3089,N_1896,N_2317);
and U3090 (N_3090,N_1831,N_2931);
or U3091 (N_3091,N_2696,N_2375);
or U3092 (N_3092,N_2333,N_2419);
and U3093 (N_3093,N_1827,N_2777);
and U3094 (N_3094,N_2314,N_2786);
nor U3095 (N_3095,N_2292,N_2475);
nand U3096 (N_3096,N_2832,N_1684);
and U3097 (N_3097,N_2052,N_2896);
or U3098 (N_3098,N_2318,N_2549);
or U3099 (N_3099,N_1699,N_2734);
and U3100 (N_3100,N_2809,N_2967);
and U3101 (N_3101,N_2792,N_1982);
nand U3102 (N_3102,N_1820,N_2798);
nand U3103 (N_3103,N_1913,N_2481);
and U3104 (N_3104,N_2032,N_2309);
nand U3105 (N_3105,N_1950,N_1798);
and U3106 (N_3106,N_1930,N_2569);
or U3107 (N_3107,N_1936,N_2946);
nor U3108 (N_3108,N_1862,N_2454);
and U3109 (N_3109,N_2255,N_2469);
and U3110 (N_3110,N_1673,N_2743);
xnor U3111 (N_3111,N_1530,N_1645);
nand U3112 (N_3112,N_2877,N_2061);
and U3113 (N_3113,N_2495,N_2937);
nor U3114 (N_3114,N_2852,N_1918);
nor U3115 (N_3115,N_1904,N_2924);
nor U3116 (N_3116,N_2408,N_1657);
nor U3117 (N_3117,N_2156,N_1888);
xnor U3118 (N_3118,N_2392,N_2409);
and U3119 (N_3119,N_2618,N_2103);
and U3120 (N_3120,N_1616,N_2568);
xor U3121 (N_3121,N_1984,N_2168);
nand U3122 (N_3122,N_2609,N_2096);
xnor U3123 (N_3123,N_2979,N_2041);
and U3124 (N_3124,N_2977,N_2519);
and U3125 (N_3125,N_2254,N_1519);
nand U3126 (N_3126,N_1634,N_2228);
nand U3127 (N_3127,N_2724,N_1702);
or U3128 (N_3128,N_2628,N_1535);
or U3129 (N_3129,N_2547,N_1576);
nand U3130 (N_3130,N_2285,N_2645);
or U3131 (N_3131,N_2094,N_2144);
and U3132 (N_3132,N_1750,N_2873);
or U3133 (N_3133,N_2070,N_1725);
and U3134 (N_3134,N_2102,N_2648);
and U3135 (N_3135,N_2653,N_2494);
nand U3136 (N_3136,N_2883,N_2744);
xnor U3137 (N_3137,N_2219,N_2835);
or U3138 (N_3138,N_2771,N_2049);
nor U3139 (N_3139,N_2658,N_2206);
nor U3140 (N_3140,N_2828,N_2350);
nor U3141 (N_3141,N_2537,N_2346);
nor U3142 (N_3142,N_2795,N_1705);
nor U3143 (N_3143,N_2216,N_2204);
and U3144 (N_3144,N_2614,N_2301);
or U3145 (N_3145,N_1560,N_1845);
or U3146 (N_3146,N_2217,N_2429);
and U3147 (N_3147,N_2018,N_2259);
or U3148 (N_3148,N_2247,N_2627);
or U3149 (N_3149,N_2253,N_2551);
and U3150 (N_3150,N_2030,N_2200);
or U3151 (N_3151,N_2955,N_1527);
or U3152 (N_3152,N_1764,N_2433);
and U3153 (N_3153,N_1929,N_1622);
or U3154 (N_3154,N_2672,N_2315);
or U3155 (N_3155,N_1855,N_2179);
nand U3156 (N_3156,N_2680,N_1958);
nor U3157 (N_3157,N_2436,N_2266);
nand U3158 (N_3158,N_2141,N_1842);
xor U3159 (N_3159,N_1901,N_2754);
and U3160 (N_3160,N_1584,N_2823);
and U3161 (N_3161,N_2157,N_1707);
nand U3162 (N_3162,N_1975,N_1534);
xor U3163 (N_3163,N_2651,N_2875);
xnor U3164 (N_3164,N_1680,N_2610);
and U3165 (N_3165,N_2690,N_2195);
nand U3166 (N_3166,N_2647,N_1974);
nand U3167 (N_3167,N_1987,N_2133);
or U3168 (N_3168,N_2170,N_1908);
and U3169 (N_3169,N_1718,N_2557);
xor U3170 (N_3170,N_2283,N_2060);
or U3171 (N_3171,N_2175,N_2386);
nand U3172 (N_3172,N_2267,N_1744);
and U3173 (N_3173,N_2132,N_2788);
nor U3174 (N_3174,N_2006,N_1952);
nand U3175 (N_3175,N_1618,N_1572);
xnor U3176 (N_3176,N_2838,N_2593);
nand U3177 (N_3177,N_2686,N_1955);
or U3178 (N_3178,N_2766,N_2613);
and U3179 (N_3179,N_2622,N_1662);
nor U3180 (N_3180,N_2670,N_2523);
and U3181 (N_3181,N_2082,N_2359);
xor U3182 (N_3182,N_1860,N_2769);
and U3183 (N_3183,N_2929,N_1588);
or U3184 (N_3184,N_2954,N_2027);
and U3185 (N_3185,N_1751,N_2491);
nor U3186 (N_3186,N_1994,N_1832);
nor U3187 (N_3187,N_1792,N_1838);
or U3188 (N_3188,N_1828,N_2281);
nor U3189 (N_3189,N_1749,N_2240);
xor U3190 (N_3190,N_2504,N_2234);
xor U3191 (N_3191,N_2348,N_1670);
nand U3192 (N_3192,N_2526,N_2555);
and U3193 (N_3193,N_2108,N_2007);
xnor U3194 (N_3194,N_2706,N_2192);
and U3195 (N_3195,N_1549,N_2236);
and U3196 (N_3196,N_2098,N_2840);
and U3197 (N_3197,N_2666,N_2483);
and U3198 (N_3198,N_2129,N_1767);
nand U3199 (N_3199,N_2802,N_2649);
nand U3200 (N_3200,N_1935,N_2400);
or U3201 (N_3201,N_1601,N_2689);
and U3202 (N_3202,N_2515,N_1771);
or U3203 (N_3203,N_2124,N_2490);
xor U3204 (N_3204,N_2363,N_2963);
nor U3205 (N_3205,N_2960,N_2335);
or U3206 (N_3206,N_2635,N_2075);
nand U3207 (N_3207,N_2939,N_2813);
nand U3208 (N_3208,N_2910,N_1778);
and U3209 (N_3209,N_2013,N_1922);
and U3210 (N_3210,N_2885,N_2665);
nand U3211 (N_3211,N_2661,N_2764);
and U3212 (N_3212,N_1633,N_2737);
or U3213 (N_3213,N_2601,N_1837);
and U3214 (N_3214,N_2922,N_1742);
or U3215 (N_3215,N_2858,N_2638);
or U3216 (N_3216,N_1907,N_1649);
or U3217 (N_3217,N_2659,N_2624);
nand U3218 (N_3218,N_1983,N_2295);
or U3219 (N_3219,N_2176,N_1824);
nor U3220 (N_3220,N_2180,N_1839);
xnor U3221 (N_3221,N_1734,N_2619);
nand U3222 (N_3222,N_2294,N_1890);
or U3223 (N_3223,N_2739,N_2721);
or U3224 (N_3224,N_2747,N_2302);
nand U3225 (N_3225,N_2932,N_2938);
or U3226 (N_3226,N_2664,N_2820);
nor U3227 (N_3227,N_2919,N_2510);
nor U3228 (N_3228,N_1668,N_2218);
nand U3229 (N_3229,N_2167,N_1583);
nand U3230 (N_3230,N_2499,N_2422);
or U3231 (N_3231,N_2608,N_2524);
nand U3232 (N_3232,N_2135,N_2498);
nand U3233 (N_3233,N_2692,N_2536);
and U3234 (N_3234,N_2559,N_2072);
nor U3235 (N_3235,N_2376,N_2999);
nor U3236 (N_3236,N_2377,N_2224);
or U3237 (N_3237,N_2759,N_1892);
xor U3238 (N_3238,N_2811,N_1585);
xor U3239 (N_3239,N_2925,N_2418);
or U3240 (N_3240,N_1700,N_2824);
and U3241 (N_3241,N_2864,N_2620);
or U3242 (N_3242,N_1558,N_2186);
nor U3243 (N_3243,N_2456,N_2365);
nand U3244 (N_3244,N_1885,N_2794);
and U3245 (N_3245,N_2394,N_2632);
xor U3246 (N_3246,N_2693,N_1682);
and U3247 (N_3247,N_2856,N_2326);
nand U3248 (N_3248,N_2451,N_2816);
nand U3249 (N_3249,N_1557,N_1573);
or U3250 (N_3250,N_1967,N_2113);
and U3251 (N_3251,N_1927,N_1696);
xnor U3252 (N_3252,N_2334,N_2574);
nor U3253 (N_3253,N_2807,N_2126);
nor U3254 (N_3254,N_2424,N_1612);
or U3255 (N_3255,N_2862,N_1921);
or U3256 (N_3256,N_2165,N_2644);
and U3257 (N_3257,N_1953,N_2839);
nor U3258 (N_3258,N_2166,N_1539);
nand U3259 (N_3259,N_2860,N_2231);
or U3260 (N_3260,N_1912,N_2948);
and U3261 (N_3261,N_2928,N_2370);
nand U3262 (N_3262,N_1900,N_2069);
or U3263 (N_3263,N_1779,N_2237);
nor U3264 (N_3264,N_2423,N_1807);
or U3265 (N_3265,N_1971,N_1577);
xnor U3266 (N_3266,N_2730,N_2406);
nand U3267 (N_3267,N_2316,N_2258);
and U3268 (N_3268,N_2450,N_2543);
nor U3269 (N_3269,N_2034,N_2417);
or U3270 (N_3270,N_2789,N_1500);
xor U3271 (N_3271,N_2514,N_2051);
nor U3272 (N_3272,N_1790,N_2540);
nor U3273 (N_3273,N_2289,N_2780);
or U3274 (N_3274,N_2570,N_2678);
xnor U3275 (N_3275,N_2468,N_1772);
and U3276 (N_3276,N_1978,N_1991);
xor U3277 (N_3277,N_1966,N_1582);
nand U3278 (N_3278,N_1891,N_2921);
nor U3279 (N_3279,N_2637,N_1548);
and U3280 (N_3280,N_2185,N_2398);
nor U3281 (N_3281,N_2448,N_2043);
xnor U3282 (N_3282,N_2591,N_2085);
or U3283 (N_3283,N_1773,N_2818);
nand U3284 (N_3284,N_1698,N_2781);
and U3285 (N_3285,N_1653,N_1532);
or U3286 (N_3286,N_2311,N_2755);
or U3287 (N_3287,N_2709,N_2726);
nand U3288 (N_3288,N_1916,N_1961);
nor U3289 (N_3289,N_2548,N_2587);
nand U3290 (N_3290,N_1879,N_1920);
nand U3291 (N_3291,N_1854,N_1716);
and U3292 (N_3292,N_2261,N_1880);
nor U3293 (N_3293,N_2194,N_2046);
nor U3294 (N_3294,N_2336,N_2303);
nor U3295 (N_3295,N_2164,N_1512);
nand U3296 (N_3296,N_1553,N_2174);
and U3297 (N_3297,N_1643,N_1986);
or U3298 (N_3298,N_2742,N_2917);
nor U3299 (N_3299,N_2011,N_2441);
xnor U3300 (N_3300,N_1803,N_2898);
xor U3301 (N_3301,N_2715,N_2466);
and U3302 (N_3302,N_2667,N_2039);
and U3303 (N_3303,N_2757,N_2151);
or U3304 (N_3304,N_2274,N_2854);
or U3305 (N_3305,N_1753,N_1830);
or U3306 (N_3306,N_1515,N_2982);
nand U3307 (N_3307,N_2863,N_2810);
or U3308 (N_3308,N_1621,N_2899);
and U3309 (N_3309,N_1501,N_2616);
nor U3310 (N_3310,N_1640,N_1509);
xor U3311 (N_3311,N_2775,N_1681);
or U3312 (N_3312,N_2432,N_2633);
nand U3313 (N_3313,N_2089,N_2506);
or U3314 (N_3314,N_1632,N_2770);
nor U3315 (N_3315,N_2354,N_1666);
or U3316 (N_3316,N_1969,N_2477);
and U3317 (N_3317,N_1979,N_1840);
nor U3318 (N_3318,N_2078,N_1939);
nand U3319 (N_3319,N_2968,N_2031);
xnor U3320 (N_3320,N_2298,N_1775);
nand U3321 (N_3321,N_2797,N_1727);
xor U3322 (N_3322,N_2478,N_2595);
nor U3323 (N_3323,N_1985,N_1656);
xor U3324 (N_3324,N_1661,N_2945);
and U3325 (N_3325,N_2290,N_2093);
nand U3326 (N_3326,N_2065,N_2566);
xor U3327 (N_3327,N_2090,N_2849);
and U3328 (N_3328,N_2464,N_2641);
nand U3329 (N_3329,N_1735,N_2268);
and U3330 (N_3330,N_1659,N_2169);
or U3331 (N_3331,N_1747,N_1794);
or U3332 (N_3332,N_1760,N_2888);
and U3333 (N_3333,N_2511,N_2304);
or U3334 (N_3334,N_1516,N_2642);
and U3335 (N_3335,N_2732,N_2630);
or U3336 (N_3336,N_1962,N_1579);
nand U3337 (N_3337,N_2291,N_2446);
nor U3338 (N_3338,N_2956,N_2337);
or U3339 (N_3339,N_2250,N_1608);
and U3340 (N_3340,N_1688,N_2545);
nor U3341 (N_3341,N_1769,N_2533);
and U3342 (N_3342,N_1637,N_2829);
or U3343 (N_3343,N_1728,N_1689);
or U3344 (N_3344,N_2836,N_1505);
nand U3345 (N_3345,N_1826,N_2246);
and U3346 (N_3346,N_2381,N_2147);
and U3347 (N_3347,N_2711,N_2325);
or U3348 (N_3348,N_1521,N_2713);
nor U3349 (N_3349,N_2462,N_1602);
or U3350 (N_3350,N_2611,N_2837);
and U3351 (N_3351,N_2509,N_2241);
or U3352 (N_3352,N_2889,N_2097);
or U3353 (N_3353,N_2162,N_1793);
or U3354 (N_3354,N_1631,N_1945);
or U3355 (N_3355,N_2353,N_2397);
nand U3356 (N_3356,N_1937,N_2220);
nand U3357 (N_3357,N_2343,N_2025);
nand U3358 (N_3358,N_2940,N_1754);
and U3359 (N_3359,N_2091,N_2313);
and U3360 (N_3360,N_2733,N_2145);
nor U3361 (N_3361,N_2668,N_2592);
nand U3362 (N_3362,N_1683,N_2959);
nor U3363 (N_3363,N_2782,N_1902);
nor U3364 (N_3364,N_1981,N_2371);
or U3365 (N_3365,N_2366,N_2805);
nor U3366 (N_3366,N_1796,N_2971);
or U3367 (N_3367,N_2332,N_1619);
or U3368 (N_3368,N_2163,N_2286);
nand U3369 (N_3369,N_2073,N_2183);
nor U3370 (N_3370,N_2579,N_1723);
xor U3371 (N_3371,N_1758,N_2479);
or U3372 (N_3372,N_2305,N_2459);
nand U3373 (N_3373,N_2585,N_2578);
or U3374 (N_3374,N_2077,N_2821);
nand U3375 (N_3375,N_2694,N_1859);
or U3376 (N_3376,N_1919,N_2914);
nand U3377 (N_3377,N_1610,N_2153);
and U3378 (N_3378,N_1973,N_2735);
nand U3379 (N_3379,N_1692,N_2330);
or U3380 (N_3380,N_2473,N_2357);
xnor U3381 (N_3381,N_1599,N_1654);
xnor U3382 (N_3382,N_2235,N_2512);
xnor U3383 (N_3383,N_1648,N_2364);
nand U3384 (N_3384,N_2556,N_2639);
and U3385 (N_3385,N_2612,N_1924);
and U3386 (N_3386,N_1660,N_2866);
or U3387 (N_3387,N_2776,N_2761);
and U3388 (N_3388,N_1672,N_2100);
and U3389 (N_3389,N_2232,N_2895);
xor U3390 (N_3390,N_1596,N_1511);
nor U3391 (N_3391,N_2284,N_2719);
or U3392 (N_3392,N_2437,N_1884);
nor U3393 (N_3393,N_1540,N_2983);
or U3394 (N_3394,N_2379,N_1864);
nand U3395 (N_3395,N_2947,N_1531);
or U3396 (N_3396,N_1867,N_2918);
nor U3397 (N_3397,N_1812,N_1703);
nand U3398 (N_3398,N_2438,N_2892);
and U3399 (N_3399,N_2911,N_2086);
and U3400 (N_3400,N_2943,N_2372);
or U3401 (N_3401,N_1898,N_2339);
nor U3402 (N_3402,N_2752,N_2951);
nand U3403 (N_3403,N_1876,N_2071);
or U3404 (N_3404,N_2038,N_1999);
and U3405 (N_3405,N_2312,N_2773);
or U3406 (N_3406,N_1871,N_2361);
nor U3407 (N_3407,N_2534,N_1537);
and U3408 (N_3408,N_2857,N_2012);
nor U3409 (N_3409,N_1825,N_1651);
and U3410 (N_3410,N_2909,N_2560);
xnor U3411 (N_3411,N_2189,N_2518);
nor U3412 (N_3412,N_1886,N_2842);
nor U3413 (N_3413,N_2594,N_2426);
xor U3414 (N_3414,N_1520,N_1685);
and U3415 (N_3415,N_1730,N_1733);
or U3416 (N_3416,N_2791,N_2431);
or U3417 (N_3417,N_1977,N_2564);
or U3418 (N_3418,N_2399,N_1677);
or U3419 (N_3419,N_2684,N_1595);
nand U3420 (N_3420,N_2362,N_2561);
nor U3421 (N_3421,N_1710,N_2673);
nand U3422 (N_3422,N_1944,N_2565);
or U3423 (N_3423,N_2942,N_1868);
xnor U3424 (N_3424,N_1708,N_2403);
or U3425 (N_3425,N_1507,N_1729);
nor U3426 (N_3426,N_2636,N_2080);
or U3427 (N_3427,N_2342,N_2193);
nor U3428 (N_3428,N_2685,N_2389);
nor U3429 (N_3429,N_2785,N_2401);
and U3430 (N_3430,N_2230,N_1598);
nand U3431 (N_3431,N_2698,N_2248);
nor U3432 (N_3432,N_2150,N_2989);
or U3433 (N_3433,N_1715,N_1543);
or U3434 (N_3434,N_2105,N_2582);
and U3435 (N_3435,N_2276,N_1954);
nand U3436 (N_3436,N_2991,N_2904);
and U3437 (N_3437,N_2282,N_2923);
nor U3438 (N_3438,N_2981,N_1517);
or U3439 (N_3439,N_2871,N_2725);
nand U3440 (N_3440,N_1565,N_2008);
nor U3441 (N_3441,N_2002,N_1895);
or U3442 (N_3442,N_2952,N_2604);
or U3443 (N_3443,N_2830,N_2416);
and U3444 (N_3444,N_1748,N_2104);
nor U3445 (N_3445,N_1988,N_2148);
nor U3446 (N_3446,N_2881,N_2784);
and U3447 (N_3447,N_2756,N_2351);
and U3448 (N_3448,N_2654,N_2452);
nand U3449 (N_3449,N_1990,N_2278);
nor U3450 (N_3450,N_2384,N_2814);
nand U3451 (N_3451,N_2239,N_2887);
nand U3452 (N_3452,N_2211,N_2876);
and U3453 (N_3453,N_2443,N_2125);
nor U3454 (N_3454,N_2682,N_2214);
or U3455 (N_3455,N_2036,N_2476);
and U3456 (N_3456,N_2987,N_2762);
and U3457 (N_3457,N_1712,N_1844);
nand U3458 (N_3458,N_1624,N_2178);
and U3459 (N_3459,N_2139,N_2953);
xnor U3460 (N_3460,N_2890,N_1502);
nor U3461 (N_3461,N_2657,N_2596);
or U3462 (N_3462,N_2826,N_1823);
or U3463 (N_3463,N_2319,N_2439);
or U3464 (N_3464,N_2879,N_2503);
xnor U3465 (N_3465,N_2710,N_2493);
and U3466 (N_3466,N_2210,N_1846);
nor U3467 (N_3467,N_2778,N_2356);
nand U3468 (N_3468,N_2087,N_2427);
nor U3469 (N_3469,N_2763,N_2603);
nor U3470 (N_3470,N_2676,N_2927);
nor U3471 (N_3471,N_1607,N_1510);
and U3472 (N_3472,N_2413,N_2444);
nor U3473 (N_3473,N_1717,N_1679);
and U3474 (N_3474,N_2800,N_2142);
nor U3475 (N_3475,N_1593,N_1630);
xnor U3476 (N_3476,N_1695,N_2501);
or U3477 (N_3477,N_2859,N_2508);
or U3478 (N_3478,N_2115,N_2421);
nor U3479 (N_3479,N_2728,N_2033);
nor U3480 (N_3480,N_1759,N_1550);
nand U3481 (N_3481,N_2660,N_2256);
xor U3482 (N_3482,N_2975,N_2272);
nor U3483 (N_3483,N_2531,N_2597);
and U3484 (N_3484,N_1768,N_1554);
nor U3485 (N_3485,N_2251,N_2279);
nand U3486 (N_3486,N_2470,N_2874);
or U3487 (N_3487,N_2327,N_1872);
nor U3488 (N_3488,N_1877,N_1836);
nand U3489 (N_3489,N_2161,N_2986);
nand U3490 (N_3490,N_2149,N_2583);
nor U3491 (N_3491,N_1822,N_2905);
or U3492 (N_3492,N_1809,N_2787);
nand U3493 (N_3493,N_1609,N_2345);
nor U3494 (N_3494,N_2550,N_2467);
nand U3495 (N_3495,N_1931,N_2016);
xnor U3496 (N_3496,N_2677,N_2222);
nor U3497 (N_3497,N_2380,N_2005);
or U3498 (N_3498,N_1693,N_2112);
nor U3499 (N_3499,N_2741,N_1724);
xor U3500 (N_3500,N_2765,N_2488);
and U3501 (N_3501,N_2750,N_1567);
nand U3502 (N_3502,N_2238,N_2385);
nand U3503 (N_3503,N_2527,N_1587);
and U3504 (N_3504,N_2486,N_1638);
or U3505 (N_3505,N_2993,N_2731);
nand U3506 (N_3506,N_2598,N_1866);
nand U3507 (N_3507,N_1664,N_2723);
nor U3508 (N_3508,N_2964,N_2841);
nor U3509 (N_3509,N_2393,N_1663);
nand U3510 (N_3510,N_2373,N_2870);
nand U3511 (N_3511,N_2390,N_2434);
xnor U3512 (N_3512,N_2621,N_1561);
nor U3513 (N_3513,N_2843,N_2544);
or U3514 (N_3514,N_1852,N_1915);
or U3515 (N_3515,N_2626,N_1770);
or U3516 (N_3516,N_2152,N_2121);
and U3517 (N_3517,N_2949,N_2825);
and U3518 (N_3518,N_1810,N_2817);
nor U3519 (N_3519,N_1523,N_2205);
and U3520 (N_3520,N_2663,N_1547);
and U3521 (N_3521,N_2275,N_1566);
nor U3522 (N_3522,N_2801,N_2374);
nor U3523 (N_3523,N_1575,N_1528);
nand U3524 (N_3524,N_2851,N_2328);
xor U3525 (N_3525,N_2383,N_1644);
and U3526 (N_3526,N_2040,N_2223);
or U3527 (N_3527,N_2846,N_2310);
nand U3528 (N_3528,N_1833,N_2962);
and U3529 (N_3529,N_1851,N_2442);
nor U3530 (N_3530,N_1541,N_2774);
and U3531 (N_3531,N_1873,N_2936);
and U3532 (N_3532,N_2867,N_2819);
nor U3533 (N_3533,N_2847,N_2465);
or U3534 (N_3534,N_2472,N_2068);
or U3535 (N_3535,N_2463,N_2930);
nor U3536 (N_3536,N_2271,N_1665);
nor U3537 (N_3537,N_2471,N_2368);
nand U3538 (N_3538,N_2137,N_2602);
and U3539 (N_3539,N_2662,N_2702);
nor U3540 (N_3540,N_1646,N_1782);
and U3541 (N_3541,N_1861,N_2378);
or U3542 (N_3542,N_1914,N_2402);
nand U3543 (N_3543,N_2119,N_1941);
nor U3544 (N_3544,N_2772,N_2542);
nand U3545 (N_3545,N_2848,N_1546);
nor U3546 (N_3546,N_2160,N_2131);
nor U3547 (N_3547,N_2209,N_2447);
and U3548 (N_3548,N_1791,N_2812);
nor U3549 (N_3549,N_2352,N_2188);
and U3550 (N_3550,N_2957,N_2720);
and U3551 (N_3551,N_2893,N_2207);
and U3552 (N_3552,N_1562,N_2081);
xnor U3553 (N_3553,N_2004,N_1814);
or U3554 (N_3554,N_2154,N_1642);
nor U3555 (N_3555,N_2307,N_1816);
nand U3556 (N_3556,N_2516,N_2492);
or U3557 (N_3557,N_1801,N_2329);
nor U3558 (N_3558,N_1544,N_2683);
xnor U3559 (N_3559,N_2969,N_2260);
nand U3560 (N_3560,N_1522,N_2970);
nand U3561 (N_3561,N_1903,N_1713);
and U3562 (N_3562,N_2655,N_2926);
xor U3563 (N_3563,N_2584,N_2541);
or U3564 (N_3564,N_1606,N_2779);
nand U3565 (N_3565,N_1714,N_1743);
or U3566 (N_3566,N_2528,N_2110);
or U3567 (N_3567,N_2404,N_2196);
or U3568 (N_3568,N_2047,N_1783);
and U3569 (N_3569,N_2130,N_2358);
or U3570 (N_3570,N_2880,N_1623);
xnor U3571 (N_3571,N_2387,N_2992);
nor U3572 (N_3572,N_2573,N_2572);
nand U3573 (N_3573,N_2703,N_2700);
xnor U3574 (N_3574,N_1697,N_2455);
and U3575 (N_3575,N_1706,N_1963);
nand U3576 (N_3576,N_2257,N_1995);
and U3577 (N_3577,N_1942,N_2606);
and U3578 (N_3578,N_1629,N_2978);
nand U3579 (N_3579,N_2749,N_1732);
or U3580 (N_3580,N_2480,N_2405);
nand U3581 (N_3581,N_1765,N_1761);
nand U3582 (N_3582,N_2738,N_2674);
nor U3583 (N_3583,N_1504,N_2306);
and U3584 (N_3584,N_1529,N_2263);
xor U3585 (N_3585,N_2575,N_2293);
and U3586 (N_3586,N_2067,N_1551);
and U3587 (N_3587,N_2058,N_2500);
nor U3588 (N_3588,N_1614,N_1701);
or U3589 (N_3589,N_2553,N_2799);
or U3590 (N_3590,N_2127,N_1849);
or U3591 (N_3591,N_2513,N_2489);
nor U3592 (N_3592,N_2884,N_1875);
nor U3593 (N_3593,N_1949,N_2714);
or U3594 (N_3594,N_2827,N_2017);
and U3595 (N_3595,N_2891,N_2001);
xnor U3596 (N_3596,N_2252,N_2407);
xnor U3597 (N_3597,N_2976,N_1788);
nand U3598 (N_3598,N_2099,N_2581);
nor U3599 (N_3599,N_2212,N_1766);
nand U3600 (N_3600,N_2722,N_2134);
nand U3601 (N_3601,N_2539,N_1674);
xor U3602 (N_3602,N_1980,N_1926);
nor U3603 (N_3603,N_1569,N_2815);
and U3604 (N_3604,N_1752,N_1795);
nor U3605 (N_3605,N_2521,N_2650);
and U3606 (N_3606,N_2520,N_1970);
nor U3607 (N_3607,N_1923,N_1722);
xnor U3608 (N_3608,N_2054,N_1592);
and U3609 (N_3609,N_1508,N_1641);
and U3610 (N_3610,N_2143,N_2485);
nor U3611 (N_3611,N_1589,N_2988);
nand U3612 (N_3612,N_2425,N_2117);
nor U3613 (N_3613,N_2717,N_2758);
and U3614 (N_3614,N_1636,N_2562);
nand U3615 (N_3615,N_2242,N_2396);
nand U3616 (N_3616,N_2640,N_2554);
xnor U3617 (N_3617,N_2872,N_2107);
nand U3618 (N_3618,N_1741,N_2355);
nor U3619 (N_3619,N_2269,N_1737);
and U3620 (N_3620,N_2916,N_1808);
or U3621 (N_3621,N_1784,N_2878);
nor U3622 (N_3622,N_2745,N_2369);
nand U3623 (N_3623,N_1533,N_2886);
or U3624 (N_3624,N_1850,N_1580);
xor U3625 (N_3625,N_1590,N_2320);
nand U3626 (N_3626,N_2300,N_2625);
nand U3627 (N_3627,N_1736,N_1591);
and U3628 (N_3628,N_2522,N_1856);
or U3629 (N_3629,N_1847,N_1538);
nand U3630 (N_3630,N_2221,N_2972);
or U3631 (N_3631,N_1594,N_2265);
and U3632 (N_3632,N_2783,N_1776);
nand U3633 (N_3633,N_1989,N_2287);
and U3634 (N_3634,N_2227,N_1882);
nand U3635 (N_3635,N_2296,N_1932);
nor U3636 (N_3636,N_2461,N_2140);
xnor U3637 (N_3637,N_2623,N_2243);
nand U3638 (N_3638,N_2804,N_2985);
and U3639 (N_3639,N_2679,N_2055);
nand U3640 (N_3640,N_2123,N_1704);
nand U3641 (N_3641,N_2349,N_1829);
nor U3642 (N_3642,N_1972,N_2063);
or U3643 (N_3643,N_1503,N_2600);
nand U3644 (N_3644,N_2120,N_2716);
or U3645 (N_3645,N_1691,N_2933);
or U3646 (N_3646,N_2736,N_1647);
or U3647 (N_3647,N_2203,N_2950);
or U3648 (N_3648,N_1834,N_2487);
nand U3649 (N_3649,N_1878,N_1525);
and U3650 (N_3650,N_2748,N_1956);
or U3651 (N_3651,N_2053,N_1611);
and U3652 (N_3652,N_2831,N_2629);
nand U3653 (N_3653,N_2159,N_2245);
and U3654 (N_3654,N_1887,N_2563);
nand U3655 (N_3655,N_1526,N_2746);
xor U3656 (N_3656,N_2009,N_2056);
or U3657 (N_3657,N_2111,N_2114);
and U3658 (N_3658,N_2643,N_2101);
nor U3659 (N_3659,N_1559,N_2226);
nor U3660 (N_3660,N_1797,N_2822);
nor U3661 (N_3661,N_1821,N_2249);
or U3662 (N_3662,N_2341,N_1800);
and U3663 (N_3663,N_2532,N_2577);
and U3664 (N_3664,N_2996,N_2727);
nand U3665 (N_3665,N_1721,N_2605);
nor U3666 (N_3666,N_1957,N_1563);
nor U3667 (N_3667,N_2687,N_1762);
nand U3668 (N_3668,N_2958,N_2023);
or U3669 (N_3669,N_2708,N_1917);
or U3670 (N_3670,N_2410,N_1899);
and U3671 (N_3671,N_2288,N_2691);
nand U3672 (N_3672,N_1687,N_1863);
nand U3673 (N_3673,N_2806,N_2497);
nor U3674 (N_3674,N_2019,N_2900);
or U3675 (N_3675,N_2704,N_2901);
and U3676 (N_3676,N_1615,N_2530);
nor U3677 (N_3677,N_1709,N_2990);
nand U3678 (N_3678,N_1881,N_2010);
nor U3679 (N_3679,N_1960,N_2482);
xor U3680 (N_3680,N_2201,N_2803);
nand U3681 (N_3681,N_2191,N_2277);
xor U3682 (N_3682,N_2048,N_2088);
nand U3683 (N_3683,N_1906,N_2669);
nor U3684 (N_3684,N_2546,N_2617);
xor U3685 (N_3685,N_2507,N_2106);
nand U3686 (N_3686,N_2414,N_2853);
or U3687 (N_3687,N_1787,N_2675);
xor U3688 (N_3688,N_1996,N_2173);
nand U3689 (N_3689,N_1928,N_1514);
xnor U3690 (N_3690,N_1597,N_2084);
xor U3691 (N_3691,N_2190,N_2517);
or U3692 (N_3692,N_1650,N_2270);
and U3693 (N_3693,N_2262,N_1545);
nand U3694 (N_3694,N_2894,N_1909);
nor U3695 (N_3695,N_1617,N_1786);
and U3696 (N_3696,N_2681,N_2233);
or U3697 (N_3697,N_1746,N_2015);
nand U3698 (N_3698,N_2388,N_2505);
nor U3699 (N_3699,N_2961,N_2915);
nor U3700 (N_3700,N_1626,N_1805);
nor U3701 (N_3701,N_2321,N_2172);
nand U3702 (N_3702,N_2430,N_2171);
and U3703 (N_3703,N_2850,N_2059);
or U3704 (N_3704,N_1720,N_2705);
and U3705 (N_3705,N_2273,N_1774);
and U3706 (N_3706,N_1513,N_1938);
nand U3707 (N_3707,N_1951,N_2331);
nand U3708 (N_3708,N_2865,N_2994);
xor U3709 (N_3709,N_2984,N_2020);
nor U3710 (N_3710,N_2215,N_1817);
and U3711 (N_3711,N_2538,N_1976);
nand U3712 (N_3712,N_2116,N_2411);
or U3713 (N_3713,N_1811,N_2908);
nand U3714 (N_3714,N_1625,N_2340);
nor U3715 (N_3715,N_1603,N_2897);
nand U3716 (N_3716,N_1869,N_2076);
nor U3717 (N_3717,N_1870,N_2021);
or U3718 (N_3718,N_2697,N_2567);
nor U3719 (N_3719,N_2966,N_1998);
xor U3720 (N_3720,N_2588,N_1848);
nor U3721 (N_3721,N_2347,N_2753);
or U3722 (N_3722,N_2796,N_2003);
nand U3723 (N_3723,N_2980,N_1893);
or U3724 (N_3724,N_2935,N_1883);
xnor U3725 (N_3725,N_2920,N_2855);
nor U3726 (N_3726,N_2913,N_1678);
and U3727 (N_3727,N_1740,N_2995);
nand U3728 (N_3728,N_2024,N_1711);
and U3729 (N_3729,N_2202,N_2701);
or U3730 (N_3730,N_2199,N_1600);
and U3731 (N_3731,N_1564,N_2440);
and U3732 (N_3732,N_2707,N_1802);
nor U3733 (N_3733,N_2136,N_1905);
and U3734 (N_3734,N_1755,N_1652);
and U3735 (N_3735,N_2861,N_2699);
nand U3736 (N_3736,N_2944,N_1690);
or U3737 (N_3737,N_1959,N_1738);
or U3738 (N_3738,N_1968,N_1813);
and U3739 (N_3739,N_1934,N_1933);
and U3740 (N_3740,N_2322,N_1789);
nand U3741 (N_3741,N_1819,N_2586);
and U3742 (N_3742,N_2902,N_1518);
or U3743 (N_3743,N_2793,N_2631);
and U3744 (N_3744,N_1628,N_2615);
or U3745 (N_3745,N_2360,N_2138);
xor U3746 (N_3746,N_1894,N_2453);
or U3747 (N_3747,N_2197,N_2182);
nor U3748 (N_3748,N_1574,N_2323);
or U3749 (N_3749,N_1857,N_1948);
or U3750 (N_3750,N_1666,N_1850);
and U3751 (N_3751,N_2474,N_2972);
xor U3752 (N_3752,N_1527,N_2446);
nor U3753 (N_3753,N_1871,N_1903);
nand U3754 (N_3754,N_2383,N_2755);
xnor U3755 (N_3755,N_1799,N_2675);
xnor U3756 (N_3756,N_2019,N_2048);
xnor U3757 (N_3757,N_1711,N_2185);
or U3758 (N_3758,N_2582,N_1967);
and U3759 (N_3759,N_2584,N_2460);
nor U3760 (N_3760,N_1742,N_1931);
nor U3761 (N_3761,N_2138,N_1935);
and U3762 (N_3762,N_2627,N_1659);
nor U3763 (N_3763,N_1650,N_2170);
or U3764 (N_3764,N_2879,N_2206);
nand U3765 (N_3765,N_1512,N_2386);
or U3766 (N_3766,N_2634,N_1509);
and U3767 (N_3767,N_2265,N_2375);
and U3768 (N_3768,N_2788,N_2864);
and U3769 (N_3769,N_2607,N_2433);
and U3770 (N_3770,N_2479,N_1531);
or U3771 (N_3771,N_2265,N_1904);
nor U3772 (N_3772,N_2716,N_2794);
and U3773 (N_3773,N_2251,N_2460);
nor U3774 (N_3774,N_2859,N_2406);
or U3775 (N_3775,N_1898,N_2660);
or U3776 (N_3776,N_2171,N_2818);
nor U3777 (N_3777,N_2727,N_2901);
nand U3778 (N_3778,N_2609,N_2775);
and U3779 (N_3779,N_1768,N_2906);
and U3780 (N_3780,N_2811,N_1791);
nand U3781 (N_3781,N_2566,N_2691);
nor U3782 (N_3782,N_2114,N_1838);
xor U3783 (N_3783,N_1746,N_2486);
and U3784 (N_3784,N_1909,N_1633);
nand U3785 (N_3785,N_2352,N_1975);
nor U3786 (N_3786,N_2754,N_2891);
or U3787 (N_3787,N_2323,N_2304);
and U3788 (N_3788,N_2195,N_1912);
or U3789 (N_3789,N_1966,N_2184);
nor U3790 (N_3790,N_1617,N_1527);
and U3791 (N_3791,N_2086,N_1554);
xor U3792 (N_3792,N_1671,N_2331);
nor U3793 (N_3793,N_1585,N_2583);
nand U3794 (N_3794,N_2301,N_1601);
or U3795 (N_3795,N_1549,N_1748);
nand U3796 (N_3796,N_2293,N_2935);
nand U3797 (N_3797,N_1632,N_1587);
or U3798 (N_3798,N_1849,N_1799);
nand U3799 (N_3799,N_2502,N_2724);
nor U3800 (N_3800,N_2691,N_2539);
nand U3801 (N_3801,N_2039,N_1889);
or U3802 (N_3802,N_2793,N_2034);
nor U3803 (N_3803,N_1654,N_2450);
nor U3804 (N_3804,N_1633,N_2225);
nor U3805 (N_3805,N_2016,N_2005);
nand U3806 (N_3806,N_2319,N_2496);
or U3807 (N_3807,N_1530,N_2697);
xor U3808 (N_3808,N_2362,N_2386);
xor U3809 (N_3809,N_1610,N_1864);
nand U3810 (N_3810,N_2097,N_1734);
nor U3811 (N_3811,N_2630,N_2381);
nor U3812 (N_3812,N_1688,N_1966);
nor U3813 (N_3813,N_1731,N_1850);
and U3814 (N_3814,N_1829,N_1509);
and U3815 (N_3815,N_2847,N_2536);
xnor U3816 (N_3816,N_1549,N_1860);
and U3817 (N_3817,N_2449,N_2221);
or U3818 (N_3818,N_2340,N_1554);
nor U3819 (N_3819,N_2319,N_2580);
nand U3820 (N_3820,N_1924,N_2898);
xnor U3821 (N_3821,N_1848,N_2334);
nand U3822 (N_3822,N_2127,N_2199);
xnor U3823 (N_3823,N_2431,N_1570);
or U3824 (N_3824,N_2846,N_2875);
xor U3825 (N_3825,N_2437,N_1945);
or U3826 (N_3826,N_2830,N_2010);
nand U3827 (N_3827,N_1627,N_2837);
nor U3828 (N_3828,N_1727,N_1711);
and U3829 (N_3829,N_2109,N_1711);
nor U3830 (N_3830,N_1579,N_2953);
and U3831 (N_3831,N_1991,N_2884);
nand U3832 (N_3832,N_2197,N_1547);
nor U3833 (N_3833,N_2302,N_2468);
or U3834 (N_3834,N_2547,N_1762);
nor U3835 (N_3835,N_1532,N_2916);
and U3836 (N_3836,N_2593,N_2996);
and U3837 (N_3837,N_2440,N_1809);
and U3838 (N_3838,N_2675,N_1574);
xnor U3839 (N_3839,N_2608,N_2355);
xor U3840 (N_3840,N_2491,N_2323);
or U3841 (N_3841,N_1980,N_2476);
nand U3842 (N_3842,N_1859,N_2258);
or U3843 (N_3843,N_2468,N_2256);
nand U3844 (N_3844,N_1690,N_2135);
xnor U3845 (N_3845,N_1765,N_2679);
nand U3846 (N_3846,N_2069,N_2584);
nand U3847 (N_3847,N_2880,N_2701);
nand U3848 (N_3848,N_2680,N_2906);
nand U3849 (N_3849,N_2349,N_2029);
and U3850 (N_3850,N_2139,N_1861);
nor U3851 (N_3851,N_2813,N_1533);
or U3852 (N_3852,N_1866,N_2286);
and U3853 (N_3853,N_2008,N_1847);
nor U3854 (N_3854,N_2284,N_2078);
and U3855 (N_3855,N_2499,N_2532);
nor U3856 (N_3856,N_2916,N_1526);
nor U3857 (N_3857,N_1984,N_2821);
xnor U3858 (N_3858,N_1818,N_1704);
nor U3859 (N_3859,N_2509,N_2372);
nor U3860 (N_3860,N_2327,N_2105);
nor U3861 (N_3861,N_2253,N_1566);
or U3862 (N_3862,N_1970,N_2483);
xor U3863 (N_3863,N_1687,N_1859);
and U3864 (N_3864,N_2120,N_2047);
and U3865 (N_3865,N_2826,N_1647);
and U3866 (N_3866,N_1902,N_1951);
xnor U3867 (N_3867,N_2440,N_1677);
or U3868 (N_3868,N_1672,N_2418);
and U3869 (N_3869,N_1965,N_2682);
or U3870 (N_3870,N_2716,N_2915);
nand U3871 (N_3871,N_2560,N_2800);
or U3872 (N_3872,N_1508,N_2445);
xor U3873 (N_3873,N_2603,N_2132);
and U3874 (N_3874,N_2147,N_2982);
xnor U3875 (N_3875,N_1850,N_2278);
nand U3876 (N_3876,N_1798,N_2035);
and U3877 (N_3877,N_1950,N_1946);
or U3878 (N_3878,N_2748,N_2044);
nand U3879 (N_3879,N_2512,N_1777);
nand U3880 (N_3880,N_2260,N_1789);
or U3881 (N_3881,N_2703,N_2082);
xor U3882 (N_3882,N_2103,N_1555);
nand U3883 (N_3883,N_1564,N_2150);
nor U3884 (N_3884,N_1685,N_2102);
or U3885 (N_3885,N_1894,N_2015);
or U3886 (N_3886,N_2221,N_2602);
and U3887 (N_3887,N_1711,N_2762);
nor U3888 (N_3888,N_2596,N_1829);
nor U3889 (N_3889,N_1736,N_1885);
nand U3890 (N_3890,N_2859,N_2088);
or U3891 (N_3891,N_2300,N_2518);
and U3892 (N_3892,N_1645,N_1657);
and U3893 (N_3893,N_2705,N_2888);
or U3894 (N_3894,N_2012,N_1732);
nand U3895 (N_3895,N_2208,N_2949);
and U3896 (N_3896,N_2598,N_1631);
and U3897 (N_3897,N_2058,N_1742);
or U3898 (N_3898,N_1689,N_2370);
and U3899 (N_3899,N_1905,N_2547);
nand U3900 (N_3900,N_1633,N_2933);
or U3901 (N_3901,N_1500,N_2432);
xnor U3902 (N_3902,N_1677,N_2940);
or U3903 (N_3903,N_2904,N_2398);
nand U3904 (N_3904,N_2075,N_1572);
or U3905 (N_3905,N_2005,N_2768);
and U3906 (N_3906,N_2157,N_2394);
and U3907 (N_3907,N_2110,N_1742);
or U3908 (N_3908,N_2618,N_2991);
nand U3909 (N_3909,N_2144,N_2399);
or U3910 (N_3910,N_2843,N_2708);
nand U3911 (N_3911,N_2638,N_2957);
and U3912 (N_3912,N_2318,N_2371);
or U3913 (N_3913,N_2386,N_1527);
and U3914 (N_3914,N_2345,N_1671);
and U3915 (N_3915,N_2247,N_2859);
nand U3916 (N_3916,N_2468,N_2899);
nor U3917 (N_3917,N_2139,N_2707);
xor U3918 (N_3918,N_2824,N_2843);
and U3919 (N_3919,N_2118,N_2549);
and U3920 (N_3920,N_1865,N_1699);
nor U3921 (N_3921,N_1982,N_1870);
xor U3922 (N_3922,N_2147,N_2217);
nor U3923 (N_3923,N_2448,N_2343);
or U3924 (N_3924,N_1837,N_1903);
nor U3925 (N_3925,N_2488,N_2674);
nand U3926 (N_3926,N_2072,N_1617);
xor U3927 (N_3927,N_2182,N_1964);
and U3928 (N_3928,N_1538,N_1830);
nor U3929 (N_3929,N_2270,N_1962);
and U3930 (N_3930,N_2789,N_2180);
nand U3931 (N_3931,N_2043,N_2693);
nor U3932 (N_3932,N_2878,N_2738);
nor U3933 (N_3933,N_2258,N_2691);
or U3934 (N_3934,N_2117,N_1502);
or U3935 (N_3935,N_2465,N_1856);
nor U3936 (N_3936,N_2434,N_2444);
and U3937 (N_3937,N_1624,N_2169);
xnor U3938 (N_3938,N_2124,N_2234);
and U3939 (N_3939,N_2635,N_2122);
or U3940 (N_3940,N_2308,N_2688);
nor U3941 (N_3941,N_1872,N_2052);
and U3942 (N_3942,N_1879,N_1953);
nor U3943 (N_3943,N_2143,N_2293);
nor U3944 (N_3944,N_2254,N_2646);
or U3945 (N_3945,N_1815,N_2726);
and U3946 (N_3946,N_2459,N_2151);
or U3947 (N_3947,N_1754,N_2261);
xnor U3948 (N_3948,N_2826,N_2950);
and U3949 (N_3949,N_2932,N_2291);
nor U3950 (N_3950,N_1591,N_2892);
or U3951 (N_3951,N_2818,N_2670);
and U3952 (N_3952,N_1952,N_1623);
nand U3953 (N_3953,N_2181,N_1839);
nor U3954 (N_3954,N_2611,N_2516);
nand U3955 (N_3955,N_2945,N_2464);
nand U3956 (N_3956,N_2360,N_2538);
or U3957 (N_3957,N_2301,N_1820);
and U3958 (N_3958,N_2495,N_1858);
and U3959 (N_3959,N_2176,N_2709);
or U3960 (N_3960,N_2548,N_1559);
and U3961 (N_3961,N_2957,N_1691);
or U3962 (N_3962,N_2928,N_2759);
nor U3963 (N_3963,N_2136,N_2413);
or U3964 (N_3964,N_2574,N_1667);
nor U3965 (N_3965,N_2175,N_2514);
or U3966 (N_3966,N_2539,N_2477);
and U3967 (N_3967,N_2998,N_2007);
or U3968 (N_3968,N_2901,N_2922);
or U3969 (N_3969,N_2665,N_2026);
or U3970 (N_3970,N_2735,N_2045);
or U3971 (N_3971,N_2528,N_1715);
or U3972 (N_3972,N_2665,N_2006);
or U3973 (N_3973,N_2819,N_2977);
xor U3974 (N_3974,N_2808,N_2830);
nand U3975 (N_3975,N_1942,N_1634);
and U3976 (N_3976,N_1660,N_1820);
and U3977 (N_3977,N_2561,N_2702);
and U3978 (N_3978,N_2404,N_1862);
or U3979 (N_3979,N_2927,N_2077);
nand U3980 (N_3980,N_1629,N_1799);
or U3981 (N_3981,N_1548,N_2079);
nor U3982 (N_3982,N_2207,N_1853);
nor U3983 (N_3983,N_1686,N_2014);
or U3984 (N_3984,N_2910,N_2504);
and U3985 (N_3985,N_2711,N_1516);
and U3986 (N_3986,N_2985,N_2849);
or U3987 (N_3987,N_2297,N_2357);
or U3988 (N_3988,N_2751,N_2358);
or U3989 (N_3989,N_2145,N_2651);
and U3990 (N_3990,N_2683,N_2524);
nor U3991 (N_3991,N_2762,N_1555);
nand U3992 (N_3992,N_2216,N_2529);
nor U3993 (N_3993,N_2416,N_2204);
nand U3994 (N_3994,N_2878,N_2405);
nand U3995 (N_3995,N_2983,N_1868);
xor U3996 (N_3996,N_2359,N_1520);
xnor U3997 (N_3997,N_2692,N_2860);
and U3998 (N_3998,N_2170,N_2863);
nand U3999 (N_3999,N_1843,N_1531);
and U4000 (N_4000,N_2234,N_2033);
nor U4001 (N_4001,N_2646,N_2322);
and U4002 (N_4002,N_2208,N_2783);
xor U4003 (N_4003,N_1510,N_2755);
nand U4004 (N_4004,N_1862,N_2055);
nor U4005 (N_4005,N_1911,N_2005);
or U4006 (N_4006,N_1902,N_1567);
xnor U4007 (N_4007,N_2926,N_2878);
nand U4008 (N_4008,N_2016,N_2834);
or U4009 (N_4009,N_1682,N_1705);
and U4010 (N_4010,N_2160,N_2890);
nor U4011 (N_4011,N_2558,N_2272);
or U4012 (N_4012,N_1666,N_2819);
or U4013 (N_4013,N_1681,N_2050);
or U4014 (N_4014,N_2700,N_2893);
nand U4015 (N_4015,N_1761,N_2173);
xor U4016 (N_4016,N_2578,N_1607);
or U4017 (N_4017,N_2988,N_2227);
nand U4018 (N_4018,N_2340,N_2795);
and U4019 (N_4019,N_2674,N_2967);
nor U4020 (N_4020,N_2942,N_2164);
nand U4021 (N_4021,N_2285,N_1824);
or U4022 (N_4022,N_2334,N_2453);
and U4023 (N_4023,N_2682,N_2295);
nand U4024 (N_4024,N_2008,N_2925);
and U4025 (N_4025,N_2888,N_2287);
nor U4026 (N_4026,N_2291,N_2022);
nor U4027 (N_4027,N_1660,N_2573);
nand U4028 (N_4028,N_1602,N_2805);
nor U4029 (N_4029,N_1700,N_2923);
nor U4030 (N_4030,N_2877,N_1888);
or U4031 (N_4031,N_2303,N_1836);
nor U4032 (N_4032,N_2477,N_2630);
nor U4033 (N_4033,N_2079,N_1972);
or U4034 (N_4034,N_2067,N_2467);
nor U4035 (N_4035,N_1514,N_2824);
or U4036 (N_4036,N_2665,N_2486);
nor U4037 (N_4037,N_1541,N_1744);
nand U4038 (N_4038,N_2359,N_2701);
nor U4039 (N_4039,N_2446,N_1604);
nand U4040 (N_4040,N_2386,N_2479);
nand U4041 (N_4041,N_2899,N_1815);
or U4042 (N_4042,N_2596,N_1926);
xor U4043 (N_4043,N_1502,N_2269);
or U4044 (N_4044,N_2736,N_2347);
nor U4045 (N_4045,N_2262,N_1858);
or U4046 (N_4046,N_2911,N_2018);
or U4047 (N_4047,N_2732,N_2675);
nand U4048 (N_4048,N_2485,N_1879);
nand U4049 (N_4049,N_2016,N_2677);
and U4050 (N_4050,N_2484,N_1776);
or U4051 (N_4051,N_2486,N_1682);
nor U4052 (N_4052,N_2411,N_1600);
or U4053 (N_4053,N_1714,N_2775);
nand U4054 (N_4054,N_2404,N_2308);
and U4055 (N_4055,N_2516,N_2320);
and U4056 (N_4056,N_2079,N_1740);
nand U4057 (N_4057,N_1597,N_2854);
nor U4058 (N_4058,N_2709,N_1644);
nand U4059 (N_4059,N_2494,N_2325);
or U4060 (N_4060,N_2997,N_2952);
and U4061 (N_4061,N_2675,N_2096);
xor U4062 (N_4062,N_1713,N_1781);
nor U4063 (N_4063,N_2167,N_2704);
nand U4064 (N_4064,N_2474,N_2885);
and U4065 (N_4065,N_2123,N_1849);
or U4066 (N_4066,N_2544,N_1981);
xor U4067 (N_4067,N_2144,N_2225);
nand U4068 (N_4068,N_1955,N_1889);
nand U4069 (N_4069,N_1598,N_2103);
and U4070 (N_4070,N_2983,N_2928);
or U4071 (N_4071,N_2036,N_1764);
nor U4072 (N_4072,N_1709,N_1880);
nand U4073 (N_4073,N_2177,N_1544);
nor U4074 (N_4074,N_2086,N_1552);
nor U4075 (N_4075,N_1958,N_1624);
xnor U4076 (N_4076,N_1673,N_1863);
or U4077 (N_4077,N_2625,N_2472);
nor U4078 (N_4078,N_2439,N_1599);
nand U4079 (N_4079,N_2008,N_1663);
or U4080 (N_4080,N_2340,N_2360);
xor U4081 (N_4081,N_2931,N_2379);
and U4082 (N_4082,N_2710,N_1713);
xnor U4083 (N_4083,N_2766,N_2011);
nand U4084 (N_4084,N_2875,N_2897);
nand U4085 (N_4085,N_2476,N_2350);
and U4086 (N_4086,N_2857,N_2896);
nor U4087 (N_4087,N_2505,N_2105);
and U4088 (N_4088,N_2129,N_2498);
or U4089 (N_4089,N_2089,N_2838);
nor U4090 (N_4090,N_2789,N_2200);
nand U4091 (N_4091,N_1611,N_2588);
nor U4092 (N_4092,N_2878,N_2594);
nand U4093 (N_4093,N_1815,N_2197);
and U4094 (N_4094,N_2434,N_2689);
xor U4095 (N_4095,N_1512,N_1883);
xnor U4096 (N_4096,N_2658,N_2438);
and U4097 (N_4097,N_1977,N_1746);
nand U4098 (N_4098,N_1504,N_2138);
and U4099 (N_4099,N_2369,N_2158);
or U4100 (N_4100,N_1709,N_2434);
and U4101 (N_4101,N_2182,N_1991);
nand U4102 (N_4102,N_2483,N_2791);
nand U4103 (N_4103,N_2572,N_2743);
nor U4104 (N_4104,N_1948,N_2003);
or U4105 (N_4105,N_1728,N_2839);
nand U4106 (N_4106,N_2651,N_2319);
nand U4107 (N_4107,N_2035,N_1553);
xnor U4108 (N_4108,N_2581,N_2967);
and U4109 (N_4109,N_1670,N_2878);
and U4110 (N_4110,N_1616,N_2324);
and U4111 (N_4111,N_2610,N_2933);
xor U4112 (N_4112,N_1899,N_2521);
nor U4113 (N_4113,N_2525,N_1802);
nand U4114 (N_4114,N_2892,N_2906);
nor U4115 (N_4115,N_2008,N_1864);
nor U4116 (N_4116,N_1858,N_2642);
or U4117 (N_4117,N_1811,N_2386);
nand U4118 (N_4118,N_2794,N_1988);
nor U4119 (N_4119,N_2858,N_2500);
or U4120 (N_4120,N_2188,N_1624);
nor U4121 (N_4121,N_2562,N_2573);
nand U4122 (N_4122,N_1786,N_2044);
and U4123 (N_4123,N_1748,N_1620);
nor U4124 (N_4124,N_1967,N_2375);
and U4125 (N_4125,N_2696,N_2197);
nand U4126 (N_4126,N_2241,N_2911);
or U4127 (N_4127,N_2828,N_1934);
or U4128 (N_4128,N_2882,N_2968);
and U4129 (N_4129,N_2047,N_2957);
nor U4130 (N_4130,N_2247,N_1681);
and U4131 (N_4131,N_1612,N_2932);
xnor U4132 (N_4132,N_2131,N_2414);
and U4133 (N_4133,N_2089,N_2685);
nand U4134 (N_4134,N_2841,N_2066);
or U4135 (N_4135,N_2921,N_2744);
or U4136 (N_4136,N_2847,N_2462);
or U4137 (N_4137,N_1853,N_2391);
xnor U4138 (N_4138,N_2863,N_2256);
nand U4139 (N_4139,N_2985,N_2268);
nor U4140 (N_4140,N_1824,N_2725);
nand U4141 (N_4141,N_1897,N_1809);
and U4142 (N_4142,N_2781,N_2080);
or U4143 (N_4143,N_2927,N_2835);
nor U4144 (N_4144,N_1777,N_1994);
nor U4145 (N_4145,N_2243,N_2899);
nand U4146 (N_4146,N_2883,N_2786);
nor U4147 (N_4147,N_1716,N_2162);
nor U4148 (N_4148,N_1728,N_2593);
nand U4149 (N_4149,N_2677,N_1701);
and U4150 (N_4150,N_2441,N_1840);
xor U4151 (N_4151,N_1874,N_2846);
or U4152 (N_4152,N_1695,N_2787);
nor U4153 (N_4153,N_1631,N_2165);
and U4154 (N_4154,N_2859,N_1860);
nor U4155 (N_4155,N_2109,N_1933);
or U4156 (N_4156,N_2945,N_2350);
nand U4157 (N_4157,N_2105,N_1592);
nor U4158 (N_4158,N_1692,N_1778);
or U4159 (N_4159,N_1834,N_1935);
or U4160 (N_4160,N_1652,N_1533);
or U4161 (N_4161,N_2480,N_2173);
nor U4162 (N_4162,N_1572,N_2492);
nor U4163 (N_4163,N_2690,N_1677);
nor U4164 (N_4164,N_2369,N_1604);
nor U4165 (N_4165,N_1956,N_2023);
or U4166 (N_4166,N_2292,N_2854);
nor U4167 (N_4167,N_1850,N_1753);
nand U4168 (N_4168,N_1521,N_2917);
nor U4169 (N_4169,N_2142,N_1979);
and U4170 (N_4170,N_1795,N_1739);
nor U4171 (N_4171,N_1881,N_1628);
nand U4172 (N_4172,N_2073,N_2297);
nand U4173 (N_4173,N_2698,N_2649);
or U4174 (N_4174,N_2560,N_2095);
nor U4175 (N_4175,N_2952,N_1849);
nand U4176 (N_4176,N_2876,N_1909);
nor U4177 (N_4177,N_2875,N_2984);
and U4178 (N_4178,N_1973,N_2102);
and U4179 (N_4179,N_1976,N_2392);
or U4180 (N_4180,N_1919,N_2023);
nor U4181 (N_4181,N_1548,N_2768);
and U4182 (N_4182,N_1962,N_1978);
and U4183 (N_4183,N_2788,N_2169);
and U4184 (N_4184,N_2604,N_1696);
nand U4185 (N_4185,N_1882,N_1535);
xnor U4186 (N_4186,N_1859,N_2817);
and U4187 (N_4187,N_2633,N_1602);
and U4188 (N_4188,N_2044,N_1755);
nand U4189 (N_4189,N_1601,N_2795);
nor U4190 (N_4190,N_1520,N_2107);
or U4191 (N_4191,N_2021,N_2342);
xnor U4192 (N_4192,N_2273,N_2587);
nand U4193 (N_4193,N_2711,N_2343);
nor U4194 (N_4194,N_2926,N_2647);
or U4195 (N_4195,N_1947,N_2120);
nor U4196 (N_4196,N_2209,N_1747);
nor U4197 (N_4197,N_2298,N_2115);
xor U4198 (N_4198,N_2526,N_2325);
or U4199 (N_4199,N_1531,N_1673);
and U4200 (N_4200,N_1952,N_2752);
or U4201 (N_4201,N_2077,N_1643);
xor U4202 (N_4202,N_1758,N_2832);
nand U4203 (N_4203,N_1902,N_1738);
nand U4204 (N_4204,N_2613,N_1678);
nor U4205 (N_4205,N_1826,N_2893);
nor U4206 (N_4206,N_2911,N_1828);
or U4207 (N_4207,N_1976,N_2590);
and U4208 (N_4208,N_2658,N_1766);
or U4209 (N_4209,N_1795,N_2600);
nor U4210 (N_4210,N_2355,N_2182);
nor U4211 (N_4211,N_2849,N_2395);
nand U4212 (N_4212,N_2189,N_2855);
xor U4213 (N_4213,N_2145,N_2496);
or U4214 (N_4214,N_1585,N_2008);
nor U4215 (N_4215,N_1697,N_1543);
or U4216 (N_4216,N_2133,N_2432);
or U4217 (N_4217,N_2670,N_2739);
and U4218 (N_4218,N_2297,N_2736);
nand U4219 (N_4219,N_2614,N_1628);
nor U4220 (N_4220,N_2762,N_2641);
nor U4221 (N_4221,N_2736,N_1763);
nor U4222 (N_4222,N_2478,N_2819);
or U4223 (N_4223,N_1516,N_1705);
nand U4224 (N_4224,N_2717,N_2757);
or U4225 (N_4225,N_1619,N_2059);
nand U4226 (N_4226,N_2213,N_2778);
and U4227 (N_4227,N_2031,N_2077);
and U4228 (N_4228,N_2778,N_2965);
and U4229 (N_4229,N_2515,N_2511);
nor U4230 (N_4230,N_2156,N_2700);
nand U4231 (N_4231,N_2193,N_1852);
and U4232 (N_4232,N_1787,N_1989);
and U4233 (N_4233,N_2458,N_2967);
nor U4234 (N_4234,N_2927,N_1514);
or U4235 (N_4235,N_2515,N_1531);
or U4236 (N_4236,N_2223,N_2194);
nor U4237 (N_4237,N_2889,N_2630);
or U4238 (N_4238,N_1699,N_2546);
and U4239 (N_4239,N_1601,N_2667);
or U4240 (N_4240,N_2840,N_2624);
nor U4241 (N_4241,N_1690,N_2481);
nor U4242 (N_4242,N_2957,N_2307);
nor U4243 (N_4243,N_2359,N_2161);
nor U4244 (N_4244,N_2789,N_2656);
and U4245 (N_4245,N_2249,N_2457);
nand U4246 (N_4246,N_2964,N_2591);
and U4247 (N_4247,N_2820,N_2777);
or U4248 (N_4248,N_1790,N_2208);
nand U4249 (N_4249,N_2572,N_1928);
nand U4250 (N_4250,N_2504,N_2215);
and U4251 (N_4251,N_1755,N_1805);
or U4252 (N_4252,N_2831,N_1519);
and U4253 (N_4253,N_2353,N_2527);
nor U4254 (N_4254,N_1729,N_2294);
nand U4255 (N_4255,N_2566,N_2197);
xnor U4256 (N_4256,N_2602,N_2115);
nand U4257 (N_4257,N_2812,N_1962);
or U4258 (N_4258,N_1996,N_2480);
nand U4259 (N_4259,N_2796,N_2768);
or U4260 (N_4260,N_2721,N_2144);
and U4261 (N_4261,N_1509,N_2674);
and U4262 (N_4262,N_2512,N_1597);
nand U4263 (N_4263,N_2293,N_2022);
nand U4264 (N_4264,N_2808,N_2646);
and U4265 (N_4265,N_2183,N_2270);
nor U4266 (N_4266,N_2244,N_1641);
nand U4267 (N_4267,N_1899,N_1569);
xnor U4268 (N_4268,N_2042,N_1573);
nand U4269 (N_4269,N_2461,N_2842);
nand U4270 (N_4270,N_2235,N_2721);
or U4271 (N_4271,N_2179,N_2112);
and U4272 (N_4272,N_1932,N_2227);
nand U4273 (N_4273,N_2888,N_2345);
xor U4274 (N_4274,N_2572,N_1709);
xor U4275 (N_4275,N_1955,N_2082);
nand U4276 (N_4276,N_1807,N_1623);
nand U4277 (N_4277,N_2940,N_2360);
and U4278 (N_4278,N_2610,N_1785);
nand U4279 (N_4279,N_2202,N_1785);
xor U4280 (N_4280,N_2440,N_1619);
nand U4281 (N_4281,N_1594,N_1920);
nor U4282 (N_4282,N_2072,N_1590);
and U4283 (N_4283,N_1846,N_2379);
or U4284 (N_4284,N_2177,N_2051);
and U4285 (N_4285,N_1983,N_1886);
nand U4286 (N_4286,N_2182,N_2360);
or U4287 (N_4287,N_2202,N_2716);
nor U4288 (N_4288,N_2079,N_2373);
nor U4289 (N_4289,N_2520,N_1521);
or U4290 (N_4290,N_2687,N_2719);
and U4291 (N_4291,N_2174,N_1897);
nor U4292 (N_4292,N_1769,N_1783);
and U4293 (N_4293,N_2680,N_2292);
and U4294 (N_4294,N_1733,N_1555);
nand U4295 (N_4295,N_2463,N_1808);
xor U4296 (N_4296,N_1559,N_1720);
or U4297 (N_4297,N_1657,N_2432);
or U4298 (N_4298,N_1986,N_2131);
and U4299 (N_4299,N_2809,N_1635);
and U4300 (N_4300,N_2462,N_2115);
nor U4301 (N_4301,N_1699,N_2803);
nor U4302 (N_4302,N_2052,N_1758);
or U4303 (N_4303,N_1839,N_2397);
and U4304 (N_4304,N_2289,N_2666);
and U4305 (N_4305,N_2179,N_1611);
and U4306 (N_4306,N_1703,N_2219);
nor U4307 (N_4307,N_2588,N_2898);
nor U4308 (N_4308,N_1779,N_2588);
xnor U4309 (N_4309,N_2954,N_2320);
nor U4310 (N_4310,N_2460,N_1885);
and U4311 (N_4311,N_2948,N_1688);
nor U4312 (N_4312,N_1773,N_2480);
and U4313 (N_4313,N_1638,N_2029);
nand U4314 (N_4314,N_1951,N_2086);
nand U4315 (N_4315,N_2851,N_2876);
nor U4316 (N_4316,N_2537,N_1769);
or U4317 (N_4317,N_2416,N_1991);
and U4318 (N_4318,N_1810,N_2082);
nor U4319 (N_4319,N_2925,N_2932);
and U4320 (N_4320,N_1993,N_2034);
or U4321 (N_4321,N_2047,N_2212);
nand U4322 (N_4322,N_2368,N_1652);
or U4323 (N_4323,N_1653,N_2214);
or U4324 (N_4324,N_1833,N_2660);
or U4325 (N_4325,N_2287,N_1566);
or U4326 (N_4326,N_1880,N_2780);
nor U4327 (N_4327,N_2606,N_2004);
or U4328 (N_4328,N_2196,N_1637);
and U4329 (N_4329,N_1686,N_2892);
nand U4330 (N_4330,N_2681,N_1850);
nor U4331 (N_4331,N_2754,N_2968);
or U4332 (N_4332,N_1924,N_1874);
nand U4333 (N_4333,N_1866,N_2816);
nand U4334 (N_4334,N_1768,N_1936);
nand U4335 (N_4335,N_2323,N_2929);
nor U4336 (N_4336,N_2351,N_1722);
nor U4337 (N_4337,N_2302,N_1566);
nor U4338 (N_4338,N_2174,N_2111);
or U4339 (N_4339,N_2703,N_1639);
nand U4340 (N_4340,N_2013,N_2395);
or U4341 (N_4341,N_1547,N_2789);
nand U4342 (N_4342,N_2029,N_2148);
nand U4343 (N_4343,N_2228,N_2678);
or U4344 (N_4344,N_2851,N_1616);
xnor U4345 (N_4345,N_2907,N_2361);
nor U4346 (N_4346,N_1840,N_2493);
xor U4347 (N_4347,N_2576,N_2625);
nand U4348 (N_4348,N_1709,N_1666);
and U4349 (N_4349,N_2215,N_2493);
and U4350 (N_4350,N_2470,N_1942);
and U4351 (N_4351,N_1752,N_1834);
and U4352 (N_4352,N_2389,N_2205);
nand U4353 (N_4353,N_2540,N_2209);
nand U4354 (N_4354,N_1974,N_2166);
nand U4355 (N_4355,N_1533,N_2568);
xor U4356 (N_4356,N_2554,N_2545);
or U4357 (N_4357,N_1882,N_2793);
nand U4358 (N_4358,N_2621,N_2763);
nand U4359 (N_4359,N_1931,N_2615);
nor U4360 (N_4360,N_2324,N_1984);
or U4361 (N_4361,N_2678,N_2645);
and U4362 (N_4362,N_2264,N_1696);
and U4363 (N_4363,N_1604,N_2632);
nor U4364 (N_4364,N_2512,N_2722);
or U4365 (N_4365,N_2717,N_1739);
xor U4366 (N_4366,N_2776,N_2812);
nor U4367 (N_4367,N_2769,N_2987);
nor U4368 (N_4368,N_1627,N_1504);
nand U4369 (N_4369,N_2892,N_1656);
or U4370 (N_4370,N_1830,N_2024);
nor U4371 (N_4371,N_2400,N_2043);
nor U4372 (N_4372,N_1806,N_2918);
and U4373 (N_4373,N_2264,N_1756);
nand U4374 (N_4374,N_2170,N_1846);
xnor U4375 (N_4375,N_2692,N_1862);
nor U4376 (N_4376,N_2720,N_2898);
xnor U4377 (N_4377,N_1749,N_1718);
nand U4378 (N_4378,N_1551,N_2540);
nor U4379 (N_4379,N_2806,N_2316);
and U4380 (N_4380,N_2520,N_2736);
or U4381 (N_4381,N_2544,N_2702);
and U4382 (N_4382,N_2917,N_1920);
nor U4383 (N_4383,N_1577,N_2276);
and U4384 (N_4384,N_2512,N_2207);
nor U4385 (N_4385,N_2298,N_2132);
nand U4386 (N_4386,N_2934,N_1967);
nor U4387 (N_4387,N_2876,N_2384);
nor U4388 (N_4388,N_2479,N_2994);
or U4389 (N_4389,N_2555,N_1835);
nand U4390 (N_4390,N_2213,N_2012);
xnor U4391 (N_4391,N_2250,N_2185);
and U4392 (N_4392,N_2062,N_2928);
nor U4393 (N_4393,N_2212,N_2625);
nand U4394 (N_4394,N_2450,N_2855);
nand U4395 (N_4395,N_2804,N_2428);
xnor U4396 (N_4396,N_2650,N_2516);
nor U4397 (N_4397,N_2247,N_2075);
nor U4398 (N_4398,N_2377,N_2157);
nand U4399 (N_4399,N_2755,N_2457);
nand U4400 (N_4400,N_1984,N_1757);
and U4401 (N_4401,N_2491,N_2774);
nand U4402 (N_4402,N_2782,N_2741);
or U4403 (N_4403,N_2556,N_2806);
or U4404 (N_4404,N_2372,N_2461);
nor U4405 (N_4405,N_2908,N_2961);
and U4406 (N_4406,N_1846,N_2608);
and U4407 (N_4407,N_1932,N_1648);
and U4408 (N_4408,N_2409,N_1513);
or U4409 (N_4409,N_2674,N_2306);
or U4410 (N_4410,N_2167,N_1989);
nor U4411 (N_4411,N_2320,N_2165);
nand U4412 (N_4412,N_2954,N_2774);
nand U4413 (N_4413,N_2604,N_1897);
nand U4414 (N_4414,N_1751,N_2717);
or U4415 (N_4415,N_2970,N_2450);
nor U4416 (N_4416,N_2723,N_2967);
xnor U4417 (N_4417,N_2314,N_2204);
and U4418 (N_4418,N_2188,N_2356);
and U4419 (N_4419,N_2532,N_2177);
nand U4420 (N_4420,N_1614,N_1568);
xnor U4421 (N_4421,N_2054,N_2248);
or U4422 (N_4422,N_2465,N_1606);
nand U4423 (N_4423,N_1845,N_2920);
and U4424 (N_4424,N_2784,N_1502);
nand U4425 (N_4425,N_2727,N_2231);
nor U4426 (N_4426,N_1755,N_2279);
nor U4427 (N_4427,N_2230,N_2278);
and U4428 (N_4428,N_2585,N_2556);
xor U4429 (N_4429,N_1986,N_2783);
xnor U4430 (N_4430,N_2647,N_2315);
nor U4431 (N_4431,N_1897,N_1753);
nand U4432 (N_4432,N_2477,N_1583);
and U4433 (N_4433,N_2850,N_1732);
nand U4434 (N_4434,N_2922,N_2221);
or U4435 (N_4435,N_2132,N_2344);
and U4436 (N_4436,N_2331,N_2429);
nand U4437 (N_4437,N_2724,N_2656);
nor U4438 (N_4438,N_1796,N_2288);
or U4439 (N_4439,N_2487,N_2214);
or U4440 (N_4440,N_1590,N_2118);
nor U4441 (N_4441,N_1859,N_1510);
or U4442 (N_4442,N_2025,N_1513);
nor U4443 (N_4443,N_2524,N_1805);
nor U4444 (N_4444,N_2738,N_1627);
nand U4445 (N_4445,N_2182,N_2935);
and U4446 (N_4446,N_1542,N_2481);
nand U4447 (N_4447,N_2346,N_1919);
or U4448 (N_4448,N_1587,N_2088);
or U4449 (N_4449,N_1729,N_2489);
xor U4450 (N_4450,N_2774,N_2216);
or U4451 (N_4451,N_2438,N_2036);
and U4452 (N_4452,N_2090,N_1714);
or U4453 (N_4453,N_1976,N_1546);
xnor U4454 (N_4454,N_1933,N_2804);
xor U4455 (N_4455,N_1965,N_2709);
or U4456 (N_4456,N_1830,N_2559);
or U4457 (N_4457,N_2621,N_2704);
and U4458 (N_4458,N_2910,N_2107);
and U4459 (N_4459,N_2287,N_1884);
and U4460 (N_4460,N_2351,N_2946);
or U4461 (N_4461,N_2166,N_2051);
nor U4462 (N_4462,N_1590,N_2524);
and U4463 (N_4463,N_2614,N_2779);
and U4464 (N_4464,N_2008,N_2607);
or U4465 (N_4465,N_1547,N_2244);
and U4466 (N_4466,N_2440,N_1526);
or U4467 (N_4467,N_2433,N_2230);
or U4468 (N_4468,N_2254,N_1827);
and U4469 (N_4469,N_1880,N_2031);
nor U4470 (N_4470,N_2000,N_2673);
nand U4471 (N_4471,N_2657,N_2082);
nand U4472 (N_4472,N_2635,N_1859);
nor U4473 (N_4473,N_2282,N_1612);
or U4474 (N_4474,N_1815,N_2738);
nand U4475 (N_4475,N_1975,N_1510);
and U4476 (N_4476,N_1663,N_2588);
or U4477 (N_4477,N_2023,N_2304);
or U4478 (N_4478,N_2737,N_2546);
or U4479 (N_4479,N_2527,N_2150);
and U4480 (N_4480,N_1789,N_1695);
and U4481 (N_4481,N_2860,N_2148);
xor U4482 (N_4482,N_2177,N_2219);
nand U4483 (N_4483,N_2194,N_2670);
or U4484 (N_4484,N_2988,N_1891);
and U4485 (N_4485,N_2357,N_2932);
nor U4486 (N_4486,N_2858,N_2695);
nor U4487 (N_4487,N_2473,N_1641);
nand U4488 (N_4488,N_2683,N_1760);
nor U4489 (N_4489,N_2722,N_1562);
nand U4490 (N_4490,N_2830,N_2762);
and U4491 (N_4491,N_1659,N_2389);
or U4492 (N_4492,N_2806,N_2125);
or U4493 (N_4493,N_2096,N_1928);
and U4494 (N_4494,N_2209,N_1936);
nand U4495 (N_4495,N_2411,N_1505);
nor U4496 (N_4496,N_1676,N_2823);
or U4497 (N_4497,N_2931,N_1656);
or U4498 (N_4498,N_2418,N_1978);
nand U4499 (N_4499,N_1518,N_2275);
or U4500 (N_4500,N_3842,N_4126);
nand U4501 (N_4501,N_3899,N_3986);
nand U4502 (N_4502,N_4187,N_3496);
or U4503 (N_4503,N_4474,N_3069);
and U4504 (N_4504,N_3573,N_4218);
or U4505 (N_4505,N_3850,N_4365);
nor U4506 (N_4506,N_4092,N_3332);
nor U4507 (N_4507,N_3703,N_3979);
or U4508 (N_4508,N_3369,N_4300);
or U4509 (N_4509,N_3556,N_3783);
nor U4510 (N_4510,N_3502,N_4395);
nor U4511 (N_4511,N_4138,N_3622);
xor U4512 (N_4512,N_3233,N_4408);
nor U4513 (N_4513,N_3206,N_4225);
or U4514 (N_4514,N_4392,N_4324);
nor U4515 (N_4515,N_3290,N_3659);
nor U4516 (N_4516,N_3358,N_3023);
nand U4517 (N_4517,N_4032,N_4255);
and U4518 (N_4518,N_3150,N_3539);
nor U4519 (N_4519,N_3221,N_3019);
nor U4520 (N_4520,N_3084,N_3061);
xnor U4521 (N_4521,N_3431,N_4337);
nor U4522 (N_4522,N_4442,N_4253);
and U4523 (N_4523,N_4307,N_4286);
xor U4524 (N_4524,N_4051,N_4322);
nand U4525 (N_4525,N_4409,N_3542);
or U4526 (N_4526,N_4022,N_3507);
nor U4527 (N_4527,N_3082,N_3446);
xnor U4528 (N_4528,N_3232,N_4393);
nand U4529 (N_4529,N_3944,N_4270);
or U4530 (N_4530,N_3643,N_4093);
and U4531 (N_4531,N_4150,N_3626);
and U4532 (N_4532,N_3183,N_3301);
nand U4533 (N_4533,N_3854,N_4122);
nand U4534 (N_4534,N_3879,N_4490);
nor U4535 (N_4535,N_3548,N_4413);
or U4536 (N_4536,N_4193,N_4134);
and U4537 (N_4537,N_3837,N_4151);
or U4538 (N_4538,N_3417,N_3202);
nand U4539 (N_4539,N_3709,N_4443);
and U4540 (N_4540,N_3445,N_3305);
and U4541 (N_4541,N_4407,N_4293);
nand U4542 (N_4542,N_3164,N_3063);
nand U4543 (N_4543,N_4470,N_3972);
or U4544 (N_4544,N_4149,N_3863);
and U4545 (N_4545,N_3179,N_3282);
or U4546 (N_4546,N_3444,N_3744);
xnor U4547 (N_4547,N_4239,N_3825);
or U4548 (N_4548,N_3068,N_3572);
nor U4549 (N_4549,N_3003,N_3043);
or U4550 (N_4550,N_4252,N_3258);
or U4551 (N_4551,N_4353,N_3508);
nor U4552 (N_4552,N_4207,N_4279);
nor U4553 (N_4553,N_3103,N_4476);
nor U4554 (N_4554,N_4308,N_3859);
or U4555 (N_4555,N_3457,N_4236);
nand U4556 (N_4556,N_3326,N_3845);
or U4557 (N_4557,N_3111,N_3857);
nand U4558 (N_4558,N_3581,N_4311);
nor U4559 (N_4559,N_4021,N_3451);
and U4560 (N_4560,N_3480,N_3815);
or U4561 (N_4561,N_4109,N_4387);
or U4562 (N_4562,N_3328,N_4352);
nand U4563 (N_4563,N_3847,N_4347);
and U4564 (N_4564,N_3216,N_3813);
nand U4565 (N_4565,N_3959,N_4176);
or U4566 (N_4566,N_3578,N_4402);
and U4567 (N_4567,N_3130,N_3797);
or U4568 (N_4568,N_3104,N_3177);
or U4569 (N_4569,N_4425,N_3283);
nand U4570 (N_4570,N_3157,N_4073);
or U4571 (N_4571,N_4209,N_3376);
and U4572 (N_4572,N_3566,N_3518);
or U4573 (N_4573,N_3575,N_4131);
and U4574 (N_4574,N_3873,N_4070);
or U4575 (N_4575,N_3561,N_3357);
and U4576 (N_4576,N_3192,N_4201);
nor U4577 (N_4577,N_3218,N_3702);
xnor U4578 (N_4578,N_3375,N_4180);
or U4579 (N_4579,N_4047,N_3299);
and U4580 (N_4580,N_3952,N_3186);
nor U4581 (N_4581,N_3577,N_3368);
nor U4582 (N_4582,N_3246,N_4119);
and U4583 (N_4583,N_3737,N_3292);
or U4584 (N_4584,N_4418,N_3670);
xnor U4585 (N_4585,N_3275,N_4289);
and U4586 (N_4586,N_3361,N_3151);
nand U4587 (N_4587,N_3285,N_3569);
and U4588 (N_4588,N_3470,N_3831);
and U4589 (N_4589,N_3145,N_4383);
and U4590 (N_4590,N_3464,N_3605);
nor U4591 (N_4591,N_4361,N_3435);
or U4592 (N_4592,N_3592,N_3909);
or U4593 (N_4593,N_3491,N_3756);
and U4594 (N_4594,N_3187,N_3726);
or U4595 (N_4595,N_4132,N_3633);
nand U4596 (N_4596,N_3208,N_3591);
nor U4597 (N_4597,N_4057,N_3385);
nor U4598 (N_4598,N_3676,N_3765);
nand U4599 (N_4599,N_4433,N_3963);
nor U4600 (N_4600,N_3038,N_3231);
or U4601 (N_4601,N_3387,N_3379);
nor U4602 (N_4602,N_3681,N_3380);
nor U4603 (N_4603,N_4229,N_4091);
xnor U4604 (N_4604,N_3168,N_4044);
nor U4605 (N_4605,N_3138,N_4344);
nor U4606 (N_4606,N_3012,N_4332);
nor U4607 (N_4607,N_3364,N_3532);
nor U4608 (N_4608,N_4019,N_4053);
or U4609 (N_4609,N_3930,N_3732);
or U4610 (N_4610,N_4364,N_3646);
and U4611 (N_4611,N_3317,N_4463);
nor U4612 (N_4612,N_3096,N_3320);
or U4613 (N_4613,N_3762,N_3757);
and U4614 (N_4614,N_3638,N_4472);
nand U4615 (N_4615,N_4055,N_3897);
or U4616 (N_4616,N_4359,N_3517);
or U4617 (N_4617,N_3399,N_4030);
or U4618 (N_4618,N_3439,N_3109);
nand U4619 (N_4619,N_4056,N_4422);
or U4620 (N_4620,N_3499,N_4196);
xor U4621 (N_4621,N_4449,N_3777);
nor U4622 (N_4622,N_3363,N_3018);
and U4623 (N_4623,N_3447,N_3913);
and U4624 (N_4624,N_4427,N_3429);
nand U4625 (N_4625,N_4245,N_4269);
and U4626 (N_4626,N_4368,N_4283);
and U4627 (N_4627,N_4379,N_3693);
or U4628 (N_4628,N_3587,N_3761);
or U4629 (N_4629,N_3014,N_4033);
nand U4630 (N_4630,N_3776,N_4054);
xnor U4631 (N_4631,N_4356,N_4220);
and U4632 (N_4632,N_4412,N_3459);
nand U4633 (N_4633,N_3461,N_3735);
nor U4634 (N_4634,N_4215,N_3818);
nor U4635 (N_4635,N_4483,N_4240);
nor U4636 (N_4636,N_3147,N_4295);
nand U4637 (N_4637,N_3821,N_3291);
or U4638 (N_4638,N_3201,N_4110);
and U4639 (N_4639,N_3957,N_4144);
or U4640 (N_4640,N_4185,N_3174);
and U4641 (N_4641,N_3475,N_4335);
nand U4642 (N_4642,N_3987,N_3421);
nand U4643 (N_4643,N_3948,N_3936);
nand U4644 (N_4644,N_3161,N_3356);
or U4645 (N_4645,N_3865,N_4204);
or U4646 (N_4646,N_3989,N_3318);
nand U4647 (N_4647,N_3809,N_4224);
or U4648 (N_4648,N_3300,N_3162);
nor U4649 (N_4649,N_3412,N_4278);
nand U4650 (N_4650,N_4008,N_3826);
and U4651 (N_4651,N_3793,N_3625);
xor U4652 (N_4652,N_4350,N_4296);
nand U4653 (N_4653,N_3734,N_3409);
and U4654 (N_4654,N_3642,N_3759);
or U4655 (N_4655,N_3701,N_3982);
and U4656 (N_4656,N_4120,N_4186);
or U4657 (N_4657,N_3214,N_4112);
nand U4658 (N_4658,N_3799,N_4417);
nor U4659 (N_4659,N_3060,N_4231);
and U4660 (N_4660,N_3611,N_3067);
nand U4661 (N_4661,N_3100,N_3665);
or U4662 (N_4662,N_3302,N_4242);
or U4663 (N_4663,N_4029,N_4199);
nand U4664 (N_4664,N_3079,N_3939);
and U4665 (N_4665,N_3105,N_3234);
nand U4666 (N_4666,N_3477,N_3712);
nand U4667 (N_4667,N_3182,N_4023);
or U4668 (N_4668,N_3054,N_3312);
nand U4669 (N_4669,N_4380,N_4128);
nand U4670 (N_4670,N_3892,N_3352);
or U4671 (N_4671,N_4377,N_3816);
xor U4672 (N_4672,N_4330,N_3789);
nor U4673 (N_4673,N_3052,N_3371);
nand U4674 (N_4674,N_4473,N_3691);
and U4675 (N_4675,N_4465,N_3918);
nor U4676 (N_4676,N_3032,N_3741);
nand U4677 (N_4677,N_3031,N_4046);
nor U4678 (N_4678,N_4080,N_4168);
xor U4679 (N_4679,N_3313,N_3306);
nor U4680 (N_4680,N_3296,N_4058);
nor U4681 (N_4681,N_4397,N_3689);
or U4682 (N_4682,N_3666,N_4262);
nand U4683 (N_4683,N_3512,N_3974);
or U4684 (N_4684,N_3133,N_3976);
or U4685 (N_4685,N_3993,N_3910);
and U4686 (N_4686,N_3881,N_3794);
and U4687 (N_4687,N_4020,N_3346);
nand U4688 (N_4688,N_4116,N_3700);
nand U4689 (N_4689,N_4299,N_3048);
nand U4690 (N_4690,N_3534,N_3230);
nor U4691 (N_4691,N_3568,N_4384);
nand U4692 (N_4692,N_3452,N_3123);
nand U4693 (N_4693,N_3880,N_3423);
and U4694 (N_4694,N_3848,N_4237);
and U4695 (N_4695,N_3450,N_3595);
nor U4696 (N_4696,N_3134,N_3335);
and U4697 (N_4697,N_3355,N_3758);
nor U4698 (N_4698,N_3805,N_3981);
or U4699 (N_4699,N_3391,N_4024);
xnor U4700 (N_4700,N_3198,N_3663);
nor U4701 (N_4701,N_3844,N_3710);
and U4702 (N_4702,N_3715,N_4174);
nand U4703 (N_4703,N_4410,N_3672);
xnor U4704 (N_4704,N_4290,N_3624);
and U4705 (N_4705,N_3740,N_3327);
nor U4706 (N_4706,N_3353,N_3339);
or U4707 (N_4707,N_3612,N_3281);
nand U4708 (N_4708,N_3303,N_4461);
nor U4709 (N_4709,N_3872,N_3427);
nor U4710 (N_4710,N_3545,N_3535);
nor U4711 (N_4711,N_3639,N_3751);
or U4712 (N_4712,N_4285,N_4235);
and U4713 (N_4713,N_3547,N_3731);
and U4714 (N_4714,N_4342,N_3253);
and U4715 (N_4715,N_3504,N_3212);
or U4716 (N_4716,N_3076,N_4437);
nor U4717 (N_4717,N_3614,N_3365);
or U4718 (N_4718,N_3754,N_4405);
or U4719 (N_4719,N_3832,N_4411);
and U4720 (N_4720,N_3252,N_3658);
and U4721 (N_4721,N_3692,N_3933);
nand U4722 (N_4722,N_3222,N_4171);
nor U4723 (N_4723,N_3228,N_4489);
or U4724 (N_4724,N_3011,N_4363);
and U4725 (N_4725,N_3268,N_4090);
nor U4726 (N_4726,N_4457,N_4165);
nor U4727 (N_4727,N_3432,N_4406);
nand U4728 (N_4728,N_4381,N_3823);
and U4729 (N_4729,N_3092,N_3466);
nor U4730 (N_4730,N_4205,N_3045);
nand U4731 (N_4731,N_4142,N_3273);
nor U4732 (N_4732,N_3126,N_4145);
or U4733 (N_4733,N_4358,N_3307);
and U4734 (N_4734,N_4447,N_3966);
nor U4735 (N_4735,N_3927,N_3738);
nand U4736 (N_4736,N_4048,N_3030);
xor U4737 (N_4737,N_4428,N_3627);
and U4738 (N_4738,N_4266,N_3645);
nand U4739 (N_4739,N_3648,N_4067);
nor U4740 (N_4740,N_3097,N_3462);
xor U4741 (N_4741,N_4388,N_4179);
nor U4742 (N_4742,N_3215,N_4014);
nand U4743 (N_4743,N_3960,N_3802);
and U4744 (N_4744,N_3264,N_3458);
and U4745 (N_4745,N_3965,N_4315);
nand U4746 (N_4746,N_4081,N_3278);
nand U4747 (N_4747,N_4261,N_3928);
or U4748 (N_4748,N_3277,N_3784);
nand U4749 (N_4749,N_3261,N_3382);
and U4750 (N_4750,N_3558,N_3235);
and U4751 (N_4751,N_4164,N_3849);
or U4752 (N_4752,N_3570,N_4265);
or U4753 (N_4753,N_3449,N_3366);
and U4754 (N_4754,N_3093,N_3634);
and U4755 (N_4755,N_3074,N_3750);
nor U4756 (N_4756,N_3773,N_3649);
nor U4757 (N_4757,N_3276,N_3597);
and U4758 (N_4758,N_3340,N_3999);
nor U4759 (N_4759,N_4336,N_3567);
and U4760 (N_4760,N_3488,N_4499);
or U4761 (N_4761,N_3687,N_3316);
nor U4762 (N_4762,N_3533,N_3425);
or U4763 (N_4763,N_3644,N_3329);
or U4764 (N_4764,N_3437,N_3563);
or U4765 (N_4765,N_3181,N_4140);
nand U4766 (N_4766,N_3184,N_3819);
nand U4767 (N_4767,N_3596,N_4498);
and U4768 (N_4768,N_3180,N_3543);
nor U4769 (N_4769,N_3293,N_3707);
or U4770 (N_4770,N_3144,N_3747);
nand U4771 (N_4771,N_4037,N_4345);
or U4772 (N_4772,N_3372,N_4223);
nor U4773 (N_4773,N_3331,N_3620);
nor U4774 (N_4774,N_3240,N_4075);
nand U4775 (N_4775,N_4370,N_3021);
nor U4776 (N_4776,N_4354,N_4107);
nor U4777 (N_4777,N_4305,N_4031);
or U4778 (N_4778,N_3322,N_3530);
or U4779 (N_4779,N_3055,N_4191);
nor U4780 (N_4780,N_4130,N_4063);
nor U4781 (N_4781,N_3260,N_3402);
and U4782 (N_4782,N_4398,N_3553);
or U4783 (N_4783,N_4163,N_4320);
or U4784 (N_4784,N_4401,N_3146);
xnor U4785 (N_4785,N_3237,N_3404);
or U4786 (N_4786,N_3397,N_3661);
nand U4787 (N_4787,N_3210,N_4233);
xor U4788 (N_4788,N_4034,N_3493);
and U4789 (N_4789,N_3217,N_4039);
nor U4790 (N_4790,N_3448,N_4178);
nor U4791 (N_4791,N_3098,N_3227);
xor U4792 (N_4792,N_3419,N_3197);
or U4793 (N_4793,N_3115,N_3058);
nand U4794 (N_4794,N_3653,N_4121);
or U4795 (N_4795,N_4087,N_3536);
or U4796 (N_4796,N_4221,N_4009);
or U4797 (N_4797,N_4040,N_3975);
nand U4798 (N_4798,N_4230,N_3997);
or U4799 (N_4799,N_4181,N_4488);
or U4800 (N_4800,N_3034,N_3651);
and U4801 (N_4801,N_3280,N_3720);
and U4802 (N_4802,N_3686,N_4202);
nor U4803 (N_4803,N_3711,N_4317);
nand U4804 (N_4804,N_3410,N_3526);
and U4805 (N_4805,N_3244,N_3549);
or U4806 (N_4806,N_3887,N_3852);
nand U4807 (N_4807,N_3698,N_4494);
and U4808 (N_4808,N_3297,N_3962);
nor U4809 (N_4809,N_3039,N_3091);
xnor U4810 (N_4810,N_3263,N_3995);
and U4811 (N_4811,N_3991,N_4195);
and U4812 (N_4812,N_4139,N_3615);
nor U4813 (N_4813,N_3000,N_4434);
nor U4814 (N_4814,N_3855,N_4281);
nand U4815 (N_4815,N_3436,N_3153);
or U4816 (N_4816,N_4183,N_3571);
nand U4817 (N_4817,N_3455,N_3631);
and U4818 (N_4818,N_3119,N_3619);
or U4819 (N_4819,N_3359,N_4329);
nand U4820 (N_4820,N_3882,N_4456);
or U4821 (N_4821,N_3473,N_3647);
nand U4822 (N_4822,N_3489,N_3071);
xnor U4823 (N_4823,N_3107,N_4156);
nand U4824 (N_4824,N_4113,N_4391);
and U4825 (N_4825,N_4303,N_3089);
or U4826 (N_4826,N_3617,N_4228);
nor U4827 (N_4827,N_4043,N_4357);
or U4828 (N_4828,N_3271,N_3623);
nor U4829 (N_4829,N_4477,N_3454);
nor U4830 (N_4830,N_3771,N_3705);
xnor U4831 (N_4831,N_3036,N_3373);
nor U4832 (N_4832,N_4349,N_3072);
and U4833 (N_4833,N_3931,N_3728);
or U4834 (N_4834,N_3652,N_4104);
and U4835 (N_4835,N_3348,N_3800);
nand U4836 (N_4836,N_3514,N_4421);
or U4837 (N_4837,N_3118,N_3868);
or U4838 (N_4838,N_3286,N_4385);
and U4839 (N_4839,N_4129,N_3487);
or U4840 (N_4840,N_3607,N_3853);
or U4841 (N_4841,N_3017,N_4097);
or U4842 (N_4842,N_3500,N_4117);
or U4843 (N_4843,N_3912,N_3416);
nor U4844 (N_4844,N_3817,N_4440);
nand U4845 (N_4845,N_4318,N_4276);
and U4846 (N_4846,N_4376,N_3781);
nand U4847 (N_4847,N_4125,N_3716);
and U4848 (N_4848,N_4026,N_3085);
nand U4849 (N_4849,N_3934,N_4069);
or U4850 (N_4850,N_3139,N_3608);
and U4851 (N_4851,N_3178,N_3890);
nor U4852 (N_4852,N_4079,N_3440);
or U4853 (N_4853,N_3041,N_3238);
nand U4854 (N_4854,N_4094,N_4256);
and U4855 (N_4855,N_4466,N_3323);
nand U4856 (N_4856,N_3010,N_3113);
or U4857 (N_4857,N_3893,N_3628);
xor U4858 (N_4858,N_3527,N_3343);
and U4859 (N_4859,N_3764,N_3158);
or U4860 (N_4860,N_3472,N_4486);
or U4861 (N_4861,N_3876,N_3769);
or U4862 (N_4862,N_3110,N_3673);
nand U4863 (N_4863,N_3945,N_3108);
nand U4864 (N_4864,N_3870,N_4160);
xnor U4865 (N_4865,N_3501,N_3694);
or U4866 (N_4866,N_4078,N_3116);
and U4867 (N_4867,N_4314,N_3977);
nor U4868 (N_4868,N_4272,N_4159);
nand U4869 (N_4869,N_3708,N_4002);
and U4870 (N_4870,N_4136,N_3827);
xnor U4871 (N_4871,N_3274,N_3128);
xor U4872 (N_4872,N_3998,N_3006);
xnor U4873 (N_4873,N_4162,N_4492);
nor U4874 (N_4874,N_4246,N_3907);
and U4875 (N_4875,N_4190,N_4250);
or U4876 (N_4876,N_3225,N_3022);
or U4877 (N_4877,N_3035,N_3603);
nand U4878 (N_4878,N_3242,N_3742);
nand U4879 (N_4879,N_3867,N_3468);
nand U4880 (N_4880,N_3519,N_3257);
or U4881 (N_4881,N_3176,N_3037);
nand U4882 (N_4882,N_4169,N_4018);
nor U4883 (N_4883,N_4103,N_3554);
nand U4884 (N_4884,N_3008,N_3748);
xor U4885 (N_4885,N_3664,N_4082);
and U4886 (N_4886,N_3669,N_3333);
nor U4887 (N_4887,N_3806,N_3262);
or U4888 (N_4888,N_3194,N_3755);
nand U4889 (N_4889,N_3170,N_3095);
and U4890 (N_4890,N_3864,N_3336);
nand U4891 (N_4891,N_3964,N_4400);
and U4892 (N_4892,N_4467,N_3334);
xnor U4893 (N_4893,N_3537,N_3269);
and U4894 (N_4894,N_3550,N_3114);
nor U4895 (N_4895,N_3564,N_3562);
nand U4896 (N_4896,N_3505,N_4025);
nor U4897 (N_4897,N_3441,N_4099);
nor U4898 (N_4898,N_4243,N_3236);
nand U4899 (N_4899,N_3479,N_3641);
or U4900 (N_4900,N_3908,N_3350);
nor U4901 (N_4901,N_3937,N_3791);
nor U4902 (N_4902,N_4212,N_4001);
and U4903 (N_4903,N_3219,N_3050);
xor U4904 (N_4904,N_3051,N_3175);
nor U4905 (N_4905,N_3256,N_3408);
nand U4906 (N_4906,N_3047,N_3398);
nand U4907 (N_4907,N_3400,N_3191);
nand U4908 (N_4908,N_3667,N_3743);
or U4909 (N_4909,N_4366,N_3745);
nor U4910 (N_4910,N_4098,N_3406);
nor U4911 (N_4911,N_3779,N_4275);
or U4912 (N_4912,N_4042,N_3433);
and U4913 (N_4913,N_3586,N_3516);
nor U4914 (N_4914,N_4423,N_3319);
and U4915 (N_4915,N_3778,N_3988);
nor U4916 (N_4916,N_4154,N_3671);
and U4917 (N_4917,N_3121,N_4292);
and U4918 (N_4918,N_3298,N_3557);
nand U4919 (N_4919,N_4462,N_3836);
and U4920 (N_4920,N_3509,N_4479);
or U4921 (N_4921,N_3420,N_3636);
or U4922 (N_4922,N_3973,N_4451);
and U4923 (N_4923,N_4394,N_3405);
and U4924 (N_4924,N_3788,N_4455);
or U4925 (N_4925,N_3985,N_4257);
nand U4926 (N_4926,N_4328,N_3824);
and U4927 (N_4927,N_3351,N_3226);
nor U4928 (N_4928,N_3248,N_3866);
or U4929 (N_4929,N_3886,N_3424);
xor U4930 (N_4930,N_4172,N_3016);
nand U4931 (N_4931,N_4260,N_4077);
nand U4932 (N_4932,N_3056,N_4127);
and U4933 (N_4933,N_4010,N_4167);
nor U4934 (N_4934,N_4334,N_3456);
or U4935 (N_4935,N_3919,N_3494);
nand U4936 (N_4936,N_4475,N_3696);
nand U4937 (N_4937,N_4309,N_3330);
and U4938 (N_4938,N_3656,N_3683);
or U4939 (N_4939,N_3524,N_4007);
xor U4940 (N_4940,N_3254,N_3902);
or U4941 (N_4941,N_3725,N_3163);
or U4942 (N_4942,N_3971,N_3722);
and U4943 (N_4943,N_3718,N_3211);
nand U4944 (N_4944,N_3338,N_3884);
nor U4945 (N_4945,N_3239,N_4182);
or U4946 (N_4946,N_3954,N_4485);
or U4947 (N_4947,N_3983,N_4439);
nor U4948 (N_4948,N_4386,N_3159);
or U4949 (N_4949,N_4282,N_3552);
or U4950 (N_4950,N_3953,N_3403);
and U4951 (N_4951,N_3838,N_3594);
and U4952 (N_4952,N_3040,N_4049);
nor U4953 (N_4953,N_3053,N_3984);
xnor U4954 (N_4954,N_3674,N_4341);
and U4955 (N_4955,N_4027,N_3858);
and U4956 (N_4956,N_4152,N_3127);
and U4957 (N_4957,N_3188,N_4389);
and U4958 (N_4958,N_3807,N_3834);
nand U4959 (N_4959,N_3266,N_3801);
xor U4960 (N_4960,N_3413,N_3888);
nand U4961 (N_4961,N_3349,N_3438);
nand U4962 (N_4962,N_4313,N_3723);
nor U4963 (N_4963,N_3780,N_3894);
nand U4964 (N_4964,N_3635,N_3090);
nor U4965 (N_4965,N_3616,N_3699);
xnor U4966 (N_4966,N_3678,N_3511);
and U4967 (N_4967,N_3044,N_3141);
nand U4968 (N_4968,N_4325,N_3467);
and U4969 (N_4969,N_4419,N_3443);
and U4970 (N_4970,N_4432,N_3407);
nand U4971 (N_4971,N_3916,N_4445);
and U4972 (N_4972,N_4066,N_4017);
and U4973 (N_4973,N_3680,N_3288);
xnor U4974 (N_4974,N_3724,N_3721);
and U4975 (N_4975,N_4390,N_4036);
or U4976 (N_4976,N_3345,N_4271);
or U4977 (N_4977,N_3024,N_4106);
nor U4978 (N_4978,N_3199,N_3830);
and U4979 (N_4979,N_4016,N_4468);
nor U4980 (N_4980,N_3200,N_3808);
nor U4981 (N_4981,N_4115,N_3767);
xnor U4982 (N_4982,N_3970,N_4089);
or U4983 (N_4983,N_4471,N_4105);
xor U4984 (N_4984,N_3310,N_3582);
and U4985 (N_4985,N_3279,N_3484);
nand U4986 (N_4986,N_3760,N_3396);
or U4987 (N_4987,N_3885,N_3682);
nand U4988 (N_4988,N_4192,N_4148);
xnor U4989 (N_4989,N_3584,N_3950);
and U4990 (N_4990,N_3655,N_3898);
nand U4991 (N_4991,N_3921,N_3704);
nand U4992 (N_4992,N_3967,N_4369);
or U4993 (N_4993,N_3083,N_3590);
nor U4994 (N_4994,N_3172,N_4346);
or U4995 (N_4995,N_3497,N_3677);
and U4996 (N_4996,N_3798,N_3020);
or U4997 (N_4997,N_4448,N_3160);
nand U4998 (N_4998,N_3106,N_3871);
nor U4999 (N_4999,N_3321,N_3049);
nor U5000 (N_5000,N_3978,N_4006);
and U5001 (N_5001,N_3422,N_3129);
nor U5002 (N_5002,N_4118,N_3195);
or U5003 (N_5003,N_3510,N_3846);
or U5004 (N_5004,N_4372,N_3002);
and U5005 (N_5005,N_3775,N_3272);
nor U5006 (N_5006,N_3001,N_3101);
or U5007 (N_5007,N_4013,N_3498);
or U5008 (N_5008,N_4326,N_4086);
xor U5009 (N_5009,N_4454,N_3630);
xnor U5010 (N_5010,N_4469,N_3015);
xor U5011 (N_5011,N_4157,N_3684);
and U5012 (N_5012,N_3875,N_4198);
or U5013 (N_5013,N_3389,N_3122);
or U5014 (N_5014,N_4360,N_3749);
and U5015 (N_5015,N_3112,N_4310);
or U5016 (N_5016,N_3362,N_3270);
nor U5017 (N_5017,N_3309,N_4101);
or U5018 (N_5018,N_4348,N_3476);
or U5019 (N_5019,N_3381,N_4203);
nand U5020 (N_5020,N_3027,N_3782);
and U5021 (N_5021,N_3026,N_3485);
or U5022 (N_5022,N_3414,N_3287);
xnor U5023 (N_5023,N_4277,N_3729);
and U5024 (N_5024,N_4264,N_3883);
and U5025 (N_5025,N_3717,N_3610);
or U5026 (N_5026,N_4362,N_4208);
and U5027 (N_5027,N_4355,N_3428);
nor U5028 (N_5028,N_3990,N_4453);
nand U5029 (N_5029,N_4102,N_3520);
nand U5030 (N_5030,N_3746,N_4248);
nand U5031 (N_5031,N_4222,N_3224);
or U5032 (N_5032,N_3377,N_3148);
or U5033 (N_5033,N_4331,N_3632);
or U5034 (N_5034,N_3383,N_3911);
nor U5035 (N_5035,N_3341,N_4478);
or U5036 (N_5036,N_4133,N_4188);
nor U5037 (N_5037,N_4267,N_4259);
nor U5038 (N_5038,N_3690,N_4373);
nand U5039 (N_5039,N_3029,N_4321);
or U5040 (N_5040,N_3482,N_3315);
or U5041 (N_5041,N_3938,N_3442);
and U5042 (N_5042,N_4487,N_4426);
nand U5043 (N_5043,N_3418,N_4062);
and U5044 (N_5044,N_3795,N_4003);
nor U5045 (N_5045,N_4460,N_3229);
xnor U5046 (N_5046,N_3066,N_3860);
nand U5047 (N_5047,N_3521,N_4095);
or U5048 (N_5048,N_3166,N_3901);
nand U5049 (N_5049,N_3169,N_4254);
nand U5050 (N_5050,N_3576,N_3923);
nor U5051 (N_5051,N_3075,N_3523);
nor U5052 (N_5052,N_3739,N_3265);
nand U5053 (N_5053,N_3152,N_3943);
nor U5054 (N_5054,N_3259,N_3295);
and U5055 (N_5055,N_4015,N_3434);
nand U5056 (N_5056,N_4219,N_3811);
and U5057 (N_5057,N_4244,N_3426);
or U5058 (N_5058,N_3070,N_4153);
nand U5059 (N_5059,N_3839,N_4306);
xor U5060 (N_5060,N_3059,N_3599);
xnor U5061 (N_5061,N_3820,N_4251);
and U5062 (N_5062,N_3142,N_4084);
and U5063 (N_5063,N_3951,N_3929);
and U5064 (N_5064,N_3958,N_3961);
or U5065 (N_5065,N_3904,N_4333);
and U5066 (N_5066,N_3471,N_4050);
nand U5067 (N_5067,N_3968,N_3102);
nand U5068 (N_5068,N_4382,N_4288);
or U5069 (N_5069,N_3785,N_4227);
nand U5070 (N_5070,N_3660,N_4083);
and U5071 (N_5071,N_4085,N_3028);
and U5072 (N_5072,N_3249,N_3205);
nand U5073 (N_5073,N_4146,N_3714);
nand U5074 (N_5074,N_3589,N_4137);
or U5075 (N_5075,N_4431,N_4114);
nand U5076 (N_5076,N_3889,N_3460);
nor U5077 (N_5077,N_3370,N_4000);
and U5078 (N_5078,N_4316,N_3165);
nor U5079 (N_5079,N_3529,N_3772);
and U5080 (N_5080,N_3598,N_3695);
nand U5081 (N_5081,N_3094,N_3917);
nand U5082 (N_5082,N_3604,N_4339);
or U5083 (N_5083,N_4481,N_3042);
and U5084 (N_5084,N_4446,N_3541);
nand U5085 (N_5085,N_3314,N_3840);
nand U5086 (N_5086,N_3609,N_3874);
nand U5087 (N_5087,N_4143,N_4197);
or U5088 (N_5088,N_3289,N_3877);
nor U5089 (N_5089,N_3390,N_4004);
xnor U5090 (N_5090,N_4175,N_3559);
and U5091 (N_5091,N_3073,N_4177);
and U5092 (N_5092,N_4459,N_3792);
or U5093 (N_5093,N_3267,N_4378);
and U5094 (N_5094,N_3600,N_3415);
and U5095 (N_5095,N_3606,N_3033);
and U5096 (N_5096,N_3149,N_3810);
nor U5097 (N_5097,N_4258,N_3025);
xor U5098 (N_5098,N_3173,N_4284);
or U5099 (N_5099,N_3551,N_3463);
nor U5100 (N_5100,N_3401,N_3668);
nor U5101 (N_5101,N_4123,N_4441);
and U5102 (N_5102,N_3515,N_3946);
nor U5103 (N_5103,N_4480,N_3618);
xnor U5104 (N_5104,N_3565,N_4496);
xor U5105 (N_5105,N_3662,N_3411);
nor U5106 (N_5106,N_3136,N_3087);
nor U5107 (N_5107,N_3796,N_3583);
and U5108 (N_5108,N_3009,N_3629);
and U5109 (N_5109,N_4323,N_3347);
nor U5110 (N_5110,N_3344,N_3956);
nor U5111 (N_5111,N_3947,N_3803);
or U5112 (N_5112,N_3980,N_3812);
xnor U5113 (N_5113,N_3367,N_3833);
nor U5114 (N_5114,N_4206,N_3465);
and U5115 (N_5115,N_4420,N_3736);
or U5116 (N_5116,N_3770,N_4302);
or U5117 (N_5117,N_3046,N_4367);
or U5118 (N_5118,N_3062,N_3540);
nor U5119 (N_5119,N_3719,N_3490);
nor U5120 (N_5120,N_3679,N_3013);
and U5121 (N_5121,N_3474,N_4438);
nor U5122 (N_5122,N_3342,N_3763);
nand U5123 (N_5123,N_3580,N_3685);
nand U5124 (N_5124,N_3190,N_4291);
xnor U5125 (N_5125,N_4403,N_3213);
nor U5126 (N_5126,N_3311,N_4217);
or U5127 (N_5127,N_3869,N_4327);
or U5128 (N_5128,N_3544,N_3940);
nand U5129 (N_5129,N_3140,N_3324);
and U5130 (N_5130,N_3495,N_3393);
and U5131 (N_5131,N_3768,N_3243);
nand U5132 (N_5132,N_3294,N_4399);
and U5133 (N_5133,N_3360,N_3675);
nand U5134 (N_5134,N_4294,N_3005);
xnor U5135 (N_5135,N_3394,N_4071);
and U5136 (N_5136,N_3065,N_3555);
nor U5137 (N_5137,N_3841,N_3560);
nand U5138 (N_5138,N_3120,N_3378);
or U5139 (N_5139,N_3453,N_4287);
and U5140 (N_5140,N_4158,N_4005);
or U5141 (N_5141,N_3325,N_4301);
or U5142 (N_5142,N_3650,N_3209);
nand U5143 (N_5143,N_4214,N_3925);
nor U5144 (N_5144,N_4312,N_3469);
nor U5145 (N_5145,N_3245,N_3430);
and U5146 (N_5146,N_3167,N_3546);
and U5147 (N_5147,N_3223,N_3117);
nand U5148 (N_5148,N_4147,N_3189);
or U5149 (N_5149,N_3914,N_3602);
nor U5150 (N_5150,N_4124,N_3915);
nand U5151 (N_5151,N_4028,N_3304);
nor U5152 (N_5152,N_4374,N_3843);
nand U5153 (N_5153,N_4096,N_3203);
and U5154 (N_5154,N_3621,N_3905);
nand U5155 (N_5155,N_3193,N_3969);
nand U5156 (N_5156,N_3354,N_3395);
nor U5157 (N_5157,N_4414,N_4424);
nor U5158 (N_5158,N_3131,N_4436);
or U5159 (N_5159,N_3528,N_3004);
or U5160 (N_5160,N_4273,N_3538);
or U5161 (N_5161,N_3706,N_4351);
and U5162 (N_5162,N_3007,N_3935);
nand U5163 (N_5163,N_4061,N_3483);
and U5164 (N_5164,N_4011,N_3125);
nor U5165 (N_5165,N_3828,N_3531);
or U5166 (N_5166,N_4404,N_4274);
or U5167 (N_5167,N_4135,N_4226);
nand U5168 (N_5168,N_3601,N_3250);
or U5169 (N_5169,N_4415,N_3155);
xor U5170 (N_5170,N_4249,N_4343);
nand U5171 (N_5171,N_4041,N_3588);
nand U5172 (N_5172,N_3727,N_4108);
or U5173 (N_5173,N_4194,N_4088);
or U5174 (N_5174,N_4263,N_3906);
nand U5175 (N_5175,N_3766,N_3220);
nor U5176 (N_5176,N_3835,N_4216);
and U5177 (N_5177,N_3903,N_3503);
or U5178 (N_5178,N_3204,N_4280);
or U5179 (N_5179,N_3774,N_3878);
xor U5180 (N_5180,N_3081,N_3088);
nand U5181 (N_5181,N_3386,N_3143);
xnor U5182 (N_5182,N_4491,N_3481);
nor U5183 (N_5183,N_3790,N_3241);
xnor U5184 (N_5184,N_3654,N_4396);
and U5185 (N_5185,N_3941,N_3896);
nor U5186 (N_5186,N_4247,N_3522);
or U5187 (N_5187,N_3733,N_3574);
and U5188 (N_5188,N_4375,N_4211);
nor U5189 (N_5189,N_4074,N_3753);
and U5190 (N_5190,N_4166,N_3924);
xor U5191 (N_5191,N_4416,N_4238);
or U5192 (N_5192,N_4319,N_3057);
and U5193 (N_5193,N_3787,N_4052);
nand U5194 (N_5194,N_3251,N_3132);
or U5195 (N_5195,N_3688,N_3851);
nor U5196 (N_5196,N_3922,N_4161);
and U5197 (N_5197,N_3185,N_4430);
or U5198 (N_5198,N_3247,N_4012);
nor U5199 (N_5199,N_4111,N_3064);
nor U5200 (N_5200,N_3697,N_3862);
xor U5201 (N_5201,N_3992,N_3308);
and U5202 (N_5202,N_3804,N_4495);
or U5203 (N_5203,N_4068,N_4064);
nand U5204 (N_5204,N_4444,N_4045);
nor U5205 (N_5205,N_3949,N_4458);
nand U5206 (N_5206,N_4371,N_4435);
and U5207 (N_5207,N_3942,N_4304);
nand U5208 (N_5208,N_4452,N_4213);
and U5209 (N_5209,N_3900,N_4141);
nand U5210 (N_5210,N_4450,N_3955);
nand U5211 (N_5211,N_3657,N_3891);
or U5212 (N_5212,N_3861,N_3786);
and U5213 (N_5213,N_4232,N_3525);
and U5214 (N_5214,N_3486,N_4482);
and U5215 (N_5215,N_4038,N_3137);
nand U5216 (N_5216,N_3730,N_4464);
nor U5217 (N_5217,N_4170,N_3156);
nor U5218 (N_5218,N_4497,N_4234);
xnor U5219 (N_5219,N_4484,N_4059);
nand U5220 (N_5220,N_4210,N_3099);
nand U5221 (N_5221,N_4060,N_4298);
nand U5222 (N_5222,N_3856,N_4340);
or U5223 (N_5223,N_4268,N_3374);
nand U5224 (N_5224,N_3384,N_3585);
or U5225 (N_5225,N_3388,N_4076);
and U5226 (N_5226,N_3613,N_3080);
and U5227 (N_5227,N_4035,N_3593);
or U5228 (N_5228,N_3579,N_3135);
xnor U5229 (N_5229,N_3640,N_3926);
nand U5230 (N_5230,N_4100,N_3637);
and U5231 (N_5231,N_4429,N_4297);
and U5232 (N_5232,N_3255,N_4065);
nand U5233 (N_5233,N_3077,N_3506);
nand U5234 (N_5234,N_3171,N_3196);
nor U5235 (N_5235,N_3932,N_4173);
xor U5236 (N_5236,N_3478,N_3822);
nand U5237 (N_5237,N_4184,N_3829);
xnor U5238 (N_5238,N_4155,N_4338);
and U5239 (N_5239,N_3086,N_3895);
or U5240 (N_5240,N_3713,N_3207);
and U5241 (N_5241,N_3996,N_3492);
nor U5242 (N_5242,N_3994,N_3154);
nor U5243 (N_5243,N_3513,N_4241);
nand U5244 (N_5244,N_4072,N_3920);
xor U5245 (N_5245,N_3752,N_3392);
nand U5246 (N_5246,N_3337,N_3124);
and U5247 (N_5247,N_3284,N_3814);
or U5248 (N_5248,N_4493,N_4200);
nand U5249 (N_5249,N_3078,N_4189);
nor U5250 (N_5250,N_3633,N_3597);
and U5251 (N_5251,N_3376,N_3661);
nand U5252 (N_5252,N_3759,N_3179);
or U5253 (N_5253,N_3149,N_3796);
nand U5254 (N_5254,N_3856,N_4010);
xor U5255 (N_5255,N_3546,N_4499);
nand U5256 (N_5256,N_3035,N_3623);
nand U5257 (N_5257,N_3869,N_4165);
or U5258 (N_5258,N_3606,N_3214);
and U5259 (N_5259,N_4381,N_4048);
nor U5260 (N_5260,N_3721,N_3372);
and U5261 (N_5261,N_3778,N_4100);
nor U5262 (N_5262,N_4172,N_4073);
and U5263 (N_5263,N_3234,N_3159);
and U5264 (N_5264,N_3945,N_3571);
xor U5265 (N_5265,N_4151,N_3000);
and U5266 (N_5266,N_3318,N_3978);
and U5267 (N_5267,N_3464,N_4402);
and U5268 (N_5268,N_4113,N_3521);
nor U5269 (N_5269,N_4113,N_3032);
or U5270 (N_5270,N_3748,N_3615);
and U5271 (N_5271,N_4069,N_3604);
xor U5272 (N_5272,N_3498,N_4181);
xnor U5273 (N_5273,N_4175,N_3845);
nand U5274 (N_5274,N_3850,N_3900);
and U5275 (N_5275,N_3367,N_3201);
xor U5276 (N_5276,N_4156,N_3920);
xor U5277 (N_5277,N_3193,N_3485);
nand U5278 (N_5278,N_3795,N_4356);
nand U5279 (N_5279,N_3154,N_3971);
or U5280 (N_5280,N_3825,N_3344);
nor U5281 (N_5281,N_3637,N_4281);
or U5282 (N_5282,N_3947,N_3354);
and U5283 (N_5283,N_3001,N_4399);
xor U5284 (N_5284,N_3574,N_4019);
or U5285 (N_5285,N_4073,N_4256);
nand U5286 (N_5286,N_3963,N_4458);
nand U5287 (N_5287,N_4471,N_4018);
nor U5288 (N_5288,N_3523,N_3622);
and U5289 (N_5289,N_4046,N_4477);
or U5290 (N_5290,N_3601,N_3734);
nand U5291 (N_5291,N_4260,N_3059);
nand U5292 (N_5292,N_3198,N_3099);
nor U5293 (N_5293,N_3474,N_4428);
nand U5294 (N_5294,N_3123,N_3614);
nor U5295 (N_5295,N_3094,N_3220);
nor U5296 (N_5296,N_4310,N_3797);
or U5297 (N_5297,N_3001,N_3681);
and U5298 (N_5298,N_4185,N_3305);
nor U5299 (N_5299,N_4269,N_3517);
nor U5300 (N_5300,N_4068,N_3367);
nor U5301 (N_5301,N_3742,N_4334);
or U5302 (N_5302,N_3826,N_4032);
xor U5303 (N_5303,N_3825,N_3120);
nand U5304 (N_5304,N_3352,N_4345);
nand U5305 (N_5305,N_4290,N_4298);
and U5306 (N_5306,N_4435,N_4161);
nor U5307 (N_5307,N_3478,N_3862);
or U5308 (N_5308,N_3527,N_4413);
and U5309 (N_5309,N_4470,N_3056);
xor U5310 (N_5310,N_3853,N_3200);
xor U5311 (N_5311,N_4028,N_4352);
and U5312 (N_5312,N_4245,N_3439);
xor U5313 (N_5313,N_3644,N_3612);
and U5314 (N_5314,N_3356,N_4476);
nor U5315 (N_5315,N_3254,N_3393);
nor U5316 (N_5316,N_3850,N_4401);
or U5317 (N_5317,N_3951,N_3345);
or U5318 (N_5318,N_3813,N_3684);
nand U5319 (N_5319,N_3413,N_4099);
or U5320 (N_5320,N_4137,N_4165);
or U5321 (N_5321,N_3900,N_4011);
nand U5322 (N_5322,N_4401,N_4057);
xnor U5323 (N_5323,N_3962,N_4378);
nor U5324 (N_5324,N_3012,N_3814);
nand U5325 (N_5325,N_3828,N_3048);
nor U5326 (N_5326,N_4134,N_4400);
and U5327 (N_5327,N_4264,N_3204);
nor U5328 (N_5328,N_3297,N_3712);
nor U5329 (N_5329,N_3478,N_3626);
nand U5330 (N_5330,N_3143,N_4492);
and U5331 (N_5331,N_3259,N_3319);
nand U5332 (N_5332,N_4443,N_3626);
or U5333 (N_5333,N_4353,N_4095);
nand U5334 (N_5334,N_4282,N_3492);
nor U5335 (N_5335,N_4320,N_3888);
and U5336 (N_5336,N_3095,N_3097);
and U5337 (N_5337,N_3893,N_4484);
and U5338 (N_5338,N_4136,N_3858);
or U5339 (N_5339,N_4297,N_3670);
or U5340 (N_5340,N_3445,N_3141);
and U5341 (N_5341,N_3853,N_4102);
nand U5342 (N_5342,N_4100,N_3755);
xnor U5343 (N_5343,N_4194,N_4258);
and U5344 (N_5344,N_4148,N_3421);
and U5345 (N_5345,N_3604,N_4367);
xor U5346 (N_5346,N_4370,N_4212);
or U5347 (N_5347,N_3084,N_3926);
nand U5348 (N_5348,N_4043,N_4356);
nand U5349 (N_5349,N_3793,N_3739);
or U5350 (N_5350,N_3393,N_4148);
or U5351 (N_5351,N_4239,N_3140);
nand U5352 (N_5352,N_3655,N_3023);
nand U5353 (N_5353,N_3143,N_3856);
nor U5354 (N_5354,N_3353,N_3399);
or U5355 (N_5355,N_3446,N_3363);
xnor U5356 (N_5356,N_3825,N_4419);
and U5357 (N_5357,N_4252,N_3251);
nor U5358 (N_5358,N_3832,N_4247);
and U5359 (N_5359,N_3254,N_4116);
nand U5360 (N_5360,N_3326,N_3915);
nor U5361 (N_5361,N_4420,N_3056);
nand U5362 (N_5362,N_3814,N_3130);
nor U5363 (N_5363,N_3423,N_4079);
nand U5364 (N_5364,N_3318,N_3692);
or U5365 (N_5365,N_3957,N_4148);
and U5366 (N_5366,N_3815,N_3838);
nand U5367 (N_5367,N_4182,N_4376);
or U5368 (N_5368,N_4422,N_4313);
or U5369 (N_5369,N_4471,N_4494);
xor U5370 (N_5370,N_4339,N_4417);
or U5371 (N_5371,N_3873,N_3299);
nor U5372 (N_5372,N_3693,N_4095);
nor U5373 (N_5373,N_3731,N_3978);
nand U5374 (N_5374,N_3328,N_3310);
or U5375 (N_5375,N_4459,N_4069);
or U5376 (N_5376,N_4278,N_4067);
and U5377 (N_5377,N_3012,N_3841);
nor U5378 (N_5378,N_3614,N_4351);
nand U5379 (N_5379,N_3694,N_3970);
and U5380 (N_5380,N_3952,N_3407);
nor U5381 (N_5381,N_3365,N_3055);
nand U5382 (N_5382,N_4380,N_4129);
nor U5383 (N_5383,N_4390,N_4447);
xnor U5384 (N_5384,N_3580,N_4346);
xnor U5385 (N_5385,N_4410,N_3886);
or U5386 (N_5386,N_3914,N_3191);
nor U5387 (N_5387,N_4193,N_4019);
or U5388 (N_5388,N_4195,N_3735);
nand U5389 (N_5389,N_3942,N_3949);
nand U5390 (N_5390,N_3237,N_4159);
nand U5391 (N_5391,N_4148,N_4486);
xor U5392 (N_5392,N_3283,N_3060);
and U5393 (N_5393,N_3269,N_4242);
nor U5394 (N_5394,N_3139,N_3223);
and U5395 (N_5395,N_3232,N_3341);
and U5396 (N_5396,N_3340,N_4161);
xor U5397 (N_5397,N_3965,N_4336);
and U5398 (N_5398,N_3374,N_4031);
and U5399 (N_5399,N_3779,N_3673);
or U5400 (N_5400,N_3132,N_3586);
nand U5401 (N_5401,N_3564,N_4255);
and U5402 (N_5402,N_3876,N_3952);
or U5403 (N_5403,N_4380,N_3154);
nand U5404 (N_5404,N_3009,N_3314);
and U5405 (N_5405,N_3165,N_4172);
and U5406 (N_5406,N_3973,N_3085);
nand U5407 (N_5407,N_3243,N_4135);
or U5408 (N_5408,N_3221,N_3395);
nand U5409 (N_5409,N_3984,N_3037);
nand U5410 (N_5410,N_3311,N_4146);
nor U5411 (N_5411,N_4021,N_3062);
and U5412 (N_5412,N_3485,N_3856);
xor U5413 (N_5413,N_4103,N_4347);
xnor U5414 (N_5414,N_3482,N_3059);
and U5415 (N_5415,N_3892,N_4448);
xor U5416 (N_5416,N_4061,N_3891);
and U5417 (N_5417,N_3964,N_3687);
nor U5418 (N_5418,N_4394,N_3254);
nand U5419 (N_5419,N_3823,N_3817);
nand U5420 (N_5420,N_3855,N_3658);
nor U5421 (N_5421,N_4432,N_4217);
nor U5422 (N_5422,N_3677,N_3850);
or U5423 (N_5423,N_3325,N_4267);
nand U5424 (N_5424,N_3477,N_3541);
nor U5425 (N_5425,N_4079,N_3799);
nor U5426 (N_5426,N_3646,N_3727);
xnor U5427 (N_5427,N_3895,N_4360);
and U5428 (N_5428,N_4318,N_4073);
and U5429 (N_5429,N_3343,N_4399);
xor U5430 (N_5430,N_3822,N_3334);
xnor U5431 (N_5431,N_3056,N_4171);
nand U5432 (N_5432,N_3694,N_3794);
nor U5433 (N_5433,N_4172,N_3246);
nand U5434 (N_5434,N_3260,N_4339);
or U5435 (N_5435,N_3436,N_3214);
and U5436 (N_5436,N_3057,N_4346);
and U5437 (N_5437,N_4492,N_4080);
xor U5438 (N_5438,N_3701,N_3946);
and U5439 (N_5439,N_4359,N_4188);
and U5440 (N_5440,N_3102,N_4249);
or U5441 (N_5441,N_3564,N_3636);
nand U5442 (N_5442,N_3804,N_3732);
and U5443 (N_5443,N_4403,N_3867);
or U5444 (N_5444,N_3672,N_3935);
or U5445 (N_5445,N_3806,N_3040);
nand U5446 (N_5446,N_3572,N_3557);
nand U5447 (N_5447,N_3814,N_4259);
and U5448 (N_5448,N_4495,N_3448);
xnor U5449 (N_5449,N_4291,N_3306);
nand U5450 (N_5450,N_4392,N_3592);
and U5451 (N_5451,N_4203,N_3495);
and U5452 (N_5452,N_3359,N_3990);
or U5453 (N_5453,N_3534,N_3810);
nand U5454 (N_5454,N_3231,N_3620);
or U5455 (N_5455,N_4095,N_3760);
nand U5456 (N_5456,N_3783,N_3384);
and U5457 (N_5457,N_3810,N_4414);
nor U5458 (N_5458,N_3616,N_4229);
nor U5459 (N_5459,N_3015,N_3885);
and U5460 (N_5460,N_4458,N_4355);
nor U5461 (N_5461,N_4277,N_4091);
or U5462 (N_5462,N_3289,N_3700);
or U5463 (N_5463,N_3870,N_4327);
nand U5464 (N_5464,N_3112,N_3228);
xnor U5465 (N_5465,N_4232,N_3504);
and U5466 (N_5466,N_3482,N_3966);
nand U5467 (N_5467,N_4073,N_4353);
nor U5468 (N_5468,N_3792,N_3759);
and U5469 (N_5469,N_3062,N_4304);
or U5470 (N_5470,N_4267,N_3513);
or U5471 (N_5471,N_3642,N_4215);
and U5472 (N_5472,N_4073,N_3655);
or U5473 (N_5473,N_3838,N_4415);
and U5474 (N_5474,N_4126,N_3995);
nor U5475 (N_5475,N_4443,N_3803);
or U5476 (N_5476,N_3595,N_3377);
or U5477 (N_5477,N_3862,N_4349);
or U5478 (N_5478,N_3818,N_3839);
nor U5479 (N_5479,N_4003,N_4258);
nor U5480 (N_5480,N_3416,N_3784);
or U5481 (N_5481,N_3980,N_3070);
xnor U5482 (N_5482,N_4308,N_3934);
nand U5483 (N_5483,N_3396,N_3931);
nor U5484 (N_5484,N_4483,N_3803);
nand U5485 (N_5485,N_3302,N_3618);
or U5486 (N_5486,N_3206,N_3303);
or U5487 (N_5487,N_3973,N_3229);
and U5488 (N_5488,N_3151,N_4425);
nand U5489 (N_5489,N_3273,N_3322);
nand U5490 (N_5490,N_4492,N_4240);
nand U5491 (N_5491,N_3781,N_3627);
and U5492 (N_5492,N_4185,N_3223);
nor U5493 (N_5493,N_3022,N_3315);
nor U5494 (N_5494,N_4425,N_3650);
or U5495 (N_5495,N_4354,N_3083);
nand U5496 (N_5496,N_3990,N_4216);
or U5497 (N_5497,N_4276,N_3690);
nor U5498 (N_5498,N_3348,N_3086);
nand U5499 (N_5499,N_4346,N_3696);
xor U5500 (N_5500,N_4315,N_3363);
nand U5501 (N_5501,N_4439,N_4327);
and U5502 (N_5502,N_3937,N_3260);
nor U5503 (N_5503,N_4486,N_3982);
and U5504 (N_5504,N_3370,N_3863);
nand U5505 (N_5505,N_3177,N_3817);
nor U5506 (N_5506,N_4218,N_4250);
and U5507 (N_5507,N_3757,N_4341);
nor U5508 (N_5508,N_3024,N_3357);
nor U5509 (N_5509,N_4152,N_3398);
nand U5510 (N_5510,N_3096,N_4011);
nand U5511 (N_5511,N_4466,N_3464);
xor U5512 (N_5512,N_3470,N_3791);
nand U5513 (N_5513,N_3666,N_3588);
nor U5514 (N_5514,N_3043,N_4024);
and U5515 (N_5515,N_3982,N_3522);
and U5516 (N_5516,N_3584,N_4359);
or U5517 (N_5517,N_3073,N_4457);
or U5518 (N_5518,N_3124,N_3178);
xnor U5519 (N_5519,N_4159,N_3123);
nand U5520 (N_5520,N_3690,N_3648);
or U5521 (N_5521,N_4483,N_3996);
and U5522 (N_5522,N_3654,N_4160);
and U5523 (N_5523,N_3488,N_3467);
xor U5524 (N_5524,N_3347,N_4193);
and U5525 (N_5525,N_3345,N_4265);
nand U5526 (N_5526,N_4269,N_3217);
nor U5527 (N_5527,N_4020,N_4303);
nand U5528 (N_5528,N_3702,N_4212);
and U5529 (N_5529,N_4024,N_3806);
and U5530 (N_5530,N_4112,N_4155);
nand U5531 (N_5531,N_3739,N_3935);
and U5532 (N_5532,N_3930,N_3606);
or U5533 (N_5533,N_3683,N_3229);
or U5534 (N_5534,N_4256,N_4489);
nand U5535 (N_5535,N_4041,N_3216);
or U5536 (N_5536,N_4378,N_3435);
and U5537 (N_5537,N_3327,N_3605);
nand U5538 (N_5538,N_3962,N_3396);
and U5539 (N_5539,N_3854,N_3323);
and U5540 (N_5540,N_3988,N_4085);
or U5541 (N_5541,N_4498,N_4067);
xor U5542 (N_5542,N_3835,N_3232);
nand U5543 (N_5543,N_4416,N_3681);
nand U5544 (N_5544,N_3011,N_3455);
and U5545 (N_5545,N_4277,N_3487);
xor U5546 (N_5546,N_4127,N_3841);
and U5547 (N_5547,N_3017,N_3857);
or U5548 (N_5548,N_3848,N_3515);
nor U5549 (N_5549,N_3300,N_3337);
xnor U5550 (N_5550,N_3892,N_3826);
or U5551 (N_5551,N_3684,N_3533);
or U5552 (N_5552,N_3499,N_4076);
nor U5553 (N_5553,N_3643,N_3723);
nor U5554 (N_5554,N_3880,N_4319);
xnor U5555 (N_5555,N_3717,N_3465);
nor U5556 (N_5556,N_3353,N_3146);
or U5557 (N_5557,N_4183,N_3777);
and U5558 (N_5558,N_3222,N_3026);
nand U5559 (N_5559,N_4032,N_3654);
and U5560 (N_5560,N_3089,N_3979);
or U5561 (N_5561,N_4106,N_4343);
nor U5562 (N_5562,N_3044,N_3672);
and U5563 (N_5563,N_4109,N_4212);
and U5564 (N_5564,N_3935,N_3142);
nor U5565 (N_5565,N_4042,N_4236);
nand U5566 (N_5566,N_3641,N_3999);
nand U5567 (N_5567,N_3180,N_3153);
nand U5568 (N_5568,N_4120,N_4382);
and U5569 (N_5569,N_4020,N_3820);
and U5570 (N_5570,N_4313,N_3626);
or U5571 (N_5571,N_4220,N_3957);
xor U5572 (N_5572,N_4266,N_3086);
nand U5573 (N_5573,N_3495,N_4449);
nand U5574 (N_5574,N_3598,N_3747);
and U5575 (N_5575,N_3957,N_3490);
nor U5576 (N_5576,N_3627,N_4007);
nand U5577 (N_5577,N_4239,N_3641);
or U5578 (N_5578,N_4125,N_3605);
or U5579 (N_5579,N_3582,N_3595);
or U5580 (N_5580,N_4055,N_3112);
nor U5581 (N_5581,N_3026,N_3601);
or U5582 (N_5582,N_3174,N_3666);
nand U5583 (N_5583,N_3671,N_4195);
xnor U5584 (N_5584,N_3694,N_3102);
and U5585 (N_5585,N_4160,N_3811);
nand U5586 (N_5586,N_4256,N_3923);
xnor U5587 (N_5587,N_4264,N_4162);
or U5588 (N_5588,N_3210,N_3423);
xnor U5589 (N_5589,N_4134,N_3415);
nor U5590 (N_5590,N_4225,N_3003);
nand U5591 (N_5591,N_4047,N_4234);
nand U5592 (N_5592,N_4148,N_4388);
or U5593 (N_5593,N_3857,N_3838);
nand U5594 (N_5594,N_3037,N_3504);
or U5595 (N_5595,N_4260,N_3107);
and U5596 (N_5596,N_3868,N_4417);
or U5597 (N_5597,N_4329,N_3601);
or U5598 (N_5598,N_3836,N_4190);
and U5599 (N_5599,N_4124,N_4068);
nand U5600 (N_5600,N_3630,N_3516);
nor U5601 (N_5601,N_4048,N_4153);
and U5602 (N_5602,N_3124,N_3189);
nand U5603 (N_5603,N_4125,N_4376);
and U5604 (N_5604,N_3861,N_3808);
nand U5605 (N_5605,N_4077,N_3354);
xnor U5606 (N_5606,N_4332,N_4226);
or U5607 (N_5607,N_4412,N_3109);
and U5608 (N_5608,N_4239,N_3498);
nor U5609 (N_5609,N_3172,N_4096);
nand U5610 (N_5610,N_3613,N_3505);
or U5611 (N_5611,N_4275,N_4197);
nand U5612 (N_5612,N_3837,N_4454);
or U5613 (N_5613,N_4032,N_3347);
xor U5614 (N_5614,N_3402,N_3943);
nand U5615 (N_5615,N_4196,N_4385);
nand U5616 (N_5616,N_3794,N_4377);
xor U5617 (N_5617,N_4250,N_3038);
nand U5618 (N_5618,N_4130,N_4197);
xnor U5619 (N_5619,N_3192,N_3324);
and U5620 (N_5620,N_4183,N_4012);
nand U5621 (N_5621,N_3174,N_3782);
and U5622 (N_5622,N_3592,N_3123);
nor U5623 (N_5623,N_4362,N_3066);
nand U5624 (N_5624,N_3235,N_3447);
nand U5625 (N_5625,N_4400,N_3275);
nor U5626 (N_5626,N_3442,N_3147);
nor U5627 (N_5627,N_4380,N_4080);
and U5628 (N_5628,N_3172,N_4463);
and U5629 (N_5629,N_3828,N_4138);
nand U5630 (N_5630,N_3978,N_4212);
or U5631 (N_5631,N_3789,N_4130);
or U5632 (N_5632,N_3004,N_4107);
nand U5633 (N_5633,N_3407,N_3318);
or U5634 (N_5634,N_4052,N_3171);
or U5635 (N_5635,N_3252,N_4394);
or U5636 (N_5636,N_3566,N_3944);
and U5637 (N_5637,N_4151,N_3462);
nand U5638 (N_5638,N_4284,N_3406);
xnor U5639 (N_5639,N_3785,N_4234);
and U5640 (N_5640,N_3225,N_3842);
nand U5641 (N_5641,N_3865,N_3401);
and U5642 (N_5642,N_3893,N_4041);
or U5643 (N_5643,N_3618,N_4222);
nand U5644 (N_5644,N_4203,N_3319);
or U5645 (N_5645,N_4337,N_3523);
nand U5646 (N_5646,N_4141,N_3520);
nand U5647 (N_5647,N_3975,N_3502);
nor U5648 (N_5648,N_3266,N_3644);
xor U5649 (N_5649,N_3166,N_4297);
or U5650 (N_5650,N_4172,N_3319);
nand U5651 (N_5651,N_3817,N_3432);
or U5652 (N_5652,N_3692,N_3101);
and U5653 (N_5653,N_3371,N_3907);
nand U5654 (N_5654,N_3433,N_3819);
and U5655 (N_5655,N_3557,N_4153);
nand U5656 (N_5656,N_4235,N_4194);
nor U5657 (N_5657,N_3527,N_3747);
nand U5658 (N_5658,N_4176,N_3854);
nand U5659 (N_5659,N_4212,N_3034);
and U5660 (N_5660,N_4470,N_3320);
nor U5661 (N_5661,N_3376,N_4244);
nor U5662 (N_5662,N_4441,N_3597);
and U5663 (N_5663,N_4141,N_3399);
or U5664 (N_5664,N_3705,N_3913);
nand U5665 (N_5665,N_4250,N_3933);
xnor U5666 (N_5666,N_3136,N_3757);
and U5667 (N_5667,N_3143,N_4387);
nor U5668 (N_5668,N_3683,N_3591);
and U5669 (N_5669,N_3525,N_4334);
nor U5670 (N_5670,N_4064,N_3152);
xnor U5671 (N_5671,N_3543,N_4064);
nand U5672 (N_5672,N_3763,N_4356);
nor U5673 (N_5673,N_3195,N_4152);
nor U5674 (N_5674,N_3298,N_4112);
and U5675 (N_5675,N_3827,N_4360);
and U5676 (N_5676,N_4015,N_3397);
and U5677 (N_5677,N_4397,N_3198);
nand U5678 (N_5678,N_3591,N_3107);
or U5679 (N_5679,N_4274,N_3130);
nor U5680 (N_5680,N_3679,N_3084);
or U5681 (N_5681,N_3642,N_3764);
nand U5682 (N_5682,N_3174,N_3142);
nor U5683 (N_5683,N_3184,N_4166);
nand U5684 (N_5684,N_3909,N_3170);
nor U5685 (N_5685,N_3830,N_3362);
or U5686 (N_5686,N_3480,N_3244);
nor U5687 (N_5687,N_3687,N_3919);
or U5688 (N_5688,N_3186,N_4405);
and U5689 (N_5689,N_3795,N_3640);
or U5690 (N_5690,N_4461,N_3253);
and U5691 (N_5691,N_3519,N_4456);
nor U5692 (N_5692,N_3572,N_4304);
or U5693 (N_5693,N_4289,N_4325);
nand U5694 (N_5694,N_3009,N_4107);
and U5695 (N_5695,N_3092,N_3899);
nor U5696 (N_5696,N_4433,N_3479);
nand U5697 (N_5697,N_3394,N_3684);
and U5698 (N_5698,N_4112,N_3853);
and U5699 (N_5699,N_3291,N_3272);
or U5700 (N_5700,N_3594,N_3753);
nand U5701 (N_5701,N_4119,N_3523);
or U5702 (N_5702,N_4018,N_4463);
and U5703 (N_5703,N_3587,N_4136);
or U5704 (N_5704,N_3623,N_3408);
or U5705 (N_5705,N_3865,N_3031);
and U5706 (N_5706,N_3971,N_4239);
or U5707 (N_5707,N_3193,N_3881);
or U5708 (N_5708,N_3808,N_3448);
nand U5709 (N_5709,N_4078,N_3469);
nand U5710 (N_5710,N_3114,N_4065);
nor U5711 (N_5711,N_3580,N_3621);
nand U5712 (N_5712,N_4439,N_4058);
nand U5713 (N_5713,N_3138,N_3781);
and U5714 (N_5714,N_3277,N_3092);
or U5715 (N_5715,N_4278,N_3833);
xor U5716 (N_5716,N_4429,N_3573);
nand U5717 (N_5717,N_3146,N_3950);
nor U5718 (N_5718,N_3825,N_4268);
nor U5719 (N_5719,N_4095,N_3067);
nand U5720 (N_5720,N_4164,N_3008);
and U5721 (N_5721,N_4101,N_4166);
or U5722 (N_5722,N_4376,N_3671);
and U5723 (N_5723,N_4265,N_4120);
nor U5724 (N_5724,N_3122,N_3802);
and U5725 (N_5725,N_3645,N_3010);
nand U5726 (N_5726,N_3625,N_4394);
nor U5727 (N_5727,N_3351,N_3319);
xor U5728 (N_5728,N_3788,N_3643);
nor U5729 (N_5729,N_4097,N_3888);
and U5730 (N_5730,N_3539,N_4444);
and U5731 (N_5731,N_4311,N_3757);
and U5732 (N_5732,N_3448,N_3521);
xor U5733 (N_5733,N_4419,N_3231);
or U5734 (N_5734,N_3782,N_3756);
and U5735 (N_5735,N_3108,N_3871);
nand U5736 (N_5736,N_4220,N_3591);
or U5737 (N_5737,N_3922,N_3597);
nor U5738 (N_5738,N_3295,N_3249);
nor U5739 (N_5739,N_3763,N_3137);
xor U5740 (N_5740,N_3174,N_3640);
nor U5741 (N_5741,N_3316,N_3513);
or U5742 (N_5742,N_3705,N_4303);
nand U5743 (N_5743,N_4141,N_4272);
nand U5744 (N_5744,N_4123,N_4198);
or U5745 (N_5745,N_4363,N_3175);
nor U5746 (N_5746,N_4268,N_4311);
xnor U5747 (N_5747,N_4048,N_3229);
nor U5748 (N_5748,N_4121,N_4448);
nand U5749 (N_5749,N_3898,N_3811);
or U5750 (N_5750,N_3828,N_3777);
nor U5751 (N_5751,N_4087,N_3179);
nand U5752 (N_5752,N_3626,N_3200);
xnor U5753 (N_5753,N_4194,N_4460);
nor U5754 (N_5754,N_3127,N_3032);
and U5755 (N_5755,N_3527,N_3877);
nand U5756 (N_5756,N_3141,N_4070);
nand U5757 (N_5757,N_3161,N_3046);
and U5758 (N_5758,N_3758,N_3716);
nor U5759 (N_5759,N_3893,N_3558);
or U5760 (N_5760,N_3971,N_3625);
nor U5761 (N_5761,N_4291,N_3003);
xnor U5762 (N_5762,N_3783,N_3972);
nor U5763 (N_5763,N_4124,N_3692);
and U5764 (N_5764,N_3390,N_3713);
nand U5765 (N_5765,N_3464,N_4149);
nand U5766 (N_5766,N_3673,N_3680);
or U5767 (N_5767,N_3106,N_3491);
and U5768 (N_5768,N_4132,N_3025);
or U5769 (N_5769,N_3859,N_3284);
nor U5770 (N_5770,N_3916,N_3345);
nor U5771 (N_5771,N_3825,N_4080);
nor U5772 (N_5772,N_4221,N_3466);
xor U5773 (N_5773,N_4368,N_4021);
nor U5774 (N_5774,N_3792,N_4385);
nor U5775 (N_5775,N_3857,N_3262);
or U5776 (N_5776,N_4030,N_3126);
and U5777 (N_5777,N_4496,N_3023);
and U5778 (N_5778,N_3059,N_3526);
or U5779 (N_5779,N_3801,N_3961);
and U5780 (N_5780,N_4483,N_4373);
xor U5781 (N_5781,N_3075,N_3332);
or U5782 (N_5782,N_3389,N_3325);
and U5783 (N_5783,N_3817,N_4176);
or U5784 (N_5784,N_4143,N_3273);
and U5785 (N_5785,N_4463,N_3861);
xor U5786 (N_5786,N_4211,N_3617);
xnor U5787 (N_5787,N_4335,N_3844);
and U5788 (N_5788,N_3863,N_3818);
nand U5789 (N_5789,N_4290,N_3276);
nand U5790 (N_5790,N_3071,N_3902);
nand U5791 (N_5791,N_3304,N_3906);
xnor U5792 (N_5792,N_3887,N_4089);
nand U5793 (N_5793,N_3239,N_3478);
nor U5794 (N_5794,N_3901,N_4313);
nand U5795 (N_5795,N_3469,N_4497);
nor U5796 (N_5796,N_4371,N_4223);
and U5797 (N_5797,N_4001,N_3524);
and U5798 (N_5798,N_4186,N_4151);
and U5799 (N_5799,N_3770,N_3890);
xnor U5800 (N_5800,N_3011,N_3956);
xnor U5801 (N_5801,N_3275,N_3400);
nor U5802 (N_5802,N_3314,N_3339);
and U5803 (N_5803,N_4283,N_4001);
or U5804 (N_5804,N_4409,N_4010);
and U5805 (N_5805,N_3097,N_3062);
nand U5806 (N_5806,N_3499,N_3387);
xnor U5807 (N_5807,N_3525,N_3582);
nand U5808 (N_5808,N_4338,N_3098);
and U5809 (N_5809,N_3404,N_4208);
xor U5810 (N_5810,N_4378,N_3586);
and U5811 (N_5811,N_3456,N_3268);
or U5812 (N_5812,N_3698,N_3057);
or U5813 (N_5813,N_4243,N_3058);
and U5814 (N_5814,N_3813,N_3091);
and U5815 (N_5815,N_4231,N_3770);
nand U5816 (N_5816,N_4406,N_3088);
or U5817 (N_5817,N_3744,N_3570);
and U5818 (N_5818,N_3644,N_3484);
xnor U5819 (N_5819,N_4170,N_3592);
nor U5820 (N_5820,N_3287,N_4323);
and U5821 (N_5821,N_3474,N_4479);
nand U5822 (N_5822,N_3821,N_3254);
nor U5823 (N_5823,N_3512,N_4099);
nor U5824 (N_5824,N_4310,N_3392);
and U5825 (N_5825,N_4077,N_4143);
and U5826 (N_5826,N_4412,N_4472);
and U5827 (N_5827,N_3938,N_4271);
or U5828 (N_5828,N_3742,N_3368);
and U5829 (N_5829,N_3705,N_3943);
and U5830 (N_5830,N_3021,N_4333);
and U5831 (N_5831,N_3662,N_4197);
or U5832 (N_5832,N_3947,N_3034);
xnor U5833 (N_5833,N_3038,N_3276);
nand U5834 (N_5834,N_4238,N_3167);
and U5835 (N_5835,N_3750,N_4306);
nand U5836 (N_5836,N_4376,N_4231);
and U5837 (N_5837,N_3517,N_3054);
nand U5838 (N_5838,N_4452,N_3048);
xnor U5839 (N_5839,N_3516,N_3560);
nand U5840 (N_5840,N_3226,N_3849);
nand U5841 (N_5841,N_3968,N_3337);
nor U5842 (N_5842,N_3381,N_4063);
nand U5843 (N_5843,N_3524,N_3411);
xnor U5844 (N_5844,N_4262,N_3334);
nand U5845 (N_5845,N_3746,N_3942);
nand U5846 (N_5846,N_3227,N_3365);
and U5847 (N_5847,N_4030,N_4001);
nand U5848 (N_5848,N_3774,N_3238);
and U5849 (N_5849,N_3931,N_3446);
xnor U5850 (N_5850,N_3031,N_3721);
nand U5851 (N_5851,N_4302,N_3671);
and U5852 (N_5852,N_3402,N_3932);
nor U5853 (N_5853,N_3189,N_3064);
and U5854 (N_5854,N_4052,N_3725);
and U5855 (N_5855,N_4097,N_4407);
xor U5856 (N_5856,N_4265,N_3014);
nor U5857 (N_5857,N_3382,N_3771);
or U5858 (N_5858,N_3316,N_3532);
nor U5859 (N_5859,N_4460,N_3215);
nand U5860 (N_5860,N_3067,N_4362);
nor U5861 (N_5861,N_3190,N_3523);
nand U5862 (N_5862,N_3128,N_3532);
or U5863 (N_5863,N_3071,N_3080);
nand U5864 (N_5864,N_3983,N_4438);
nand U5865 (N_5865,N_3699,N_4397);
nand U5866 (N_5866,N_4070,N_3418);
and U5867 (N_5867,N_4129,N_3751);
nand U5868 (N_5868,N_3967,N_3450);
and U5869 (N_5869,N_3739,N_4497);
and U5870 (N_5870,N_3119,N_3395);
nand U5871 (N_5871,N_4032,N_4099);
nor U5872 (N_5872,N_4486,N_3015);
nand U5873 (N_5873,N_4327,N_4017);
nand U5874 (N_5874,N_4238,N_3236);
or U5875 (N_5875,N_4173,N_3759);
nand U5876 (N_5876,N_3351,N_3452);
xor U5877 (N_5877,N_4418,N_3577);
or U5878 (N_5878,N_4485,N_3723);
and U5879 (N_5879,N_4395,N_3286);
nand U5880 (N_5880,N_3383,N_3778);
xnor U5881 (N_5881,N_4041,N_4083);
nand U5882 (N_5882,N_3361,N_4147);
nand U5883 (N_5883,N_3081,N_4326);
or U5884 (N_5884,N_3075,N_3462);
and U5885 (N_5885,N_3540,N_3230);
or U5886 (N_5886,N_3102,N_3329);
xor U5887 (N_5887,N_3376,N_3549);
nor U5888 (N_5888,N_3413,N_3610);
or U5889 (N_5889,N_3967,N_4204);
nand U5890 (N_5890,N_3714,N_4389);
nand U5891 (N_5891,N_3731,N_4458);
nand U5892 (N_5892,N_3634,N_3090);
or U5893 (N_5893,N_3517,N_3833);
nor U5894 (N_5894,N_4371,N_4464);
nor U5895 (N_5895,N_4178,N_3883);
nand U5896 (N_5896,N_3839,N_3918);
nor U5897 (N_5897,N_3213,N_4368);
xnor U5898 (N_5898,N_3056,N_3619);
nand U5899 (N_5899,N_3149,N_3457);
and U5900 (N_5900,N_4134,N_3917);
xor U5901 (N_5901,N_3927,N_4180);
xnor U5902 (N_5902,N_3849,N_4248);
nand U5903 (N_5903,N_3990,N_3317);
nor U5904 (N_5904,N_3930,N_3394);
nand U5905 (N_5905,N_3713,N_3172);
nor U5906 (N_5906,N_3930,N_3470);
nand U5907 (N_5907,N_3142,N_4451);
nor U5908 (N_5908,N_4452,N_3609);
nor U5909 (N_5909,N_3559,N_3371);
or U5910 (N_5910,N_3020,N_4165);
or U5911 (N_5911,N_3527,N_4101);
nand U5912 (N_5912,N_3845,N_3634);
or U5913 (N_5913,N_3569,N_3260);
nand U5914 (N_5914,N_3241,N_4166);
nand U5915 (N_5915,N_4295,N_3185);
nor U5916 (N_5916,N_3693,N_4313);
nand U5917 (N_5917,N_3115,N_3215);
nor U5918 (N_5918,N_3277,N_3752);
and U5919 (N_5919,N_4289,N_3462);
nor U5920 (N_5920,N_3747,N_3289);
nor U5921 (N_5921,N_3546,N_3373);
and U5922 (N_5922,N_3169,N_4370);
or U5923 (N_5923,N_4235,N_4153);
or U5924 (N_5924,N_4259,N_3713);
nor U5925 (N_5925,N_4484,N_3081);
or U5926 (N_5926,N_3728,N_3004);
nor U5927 (N_5927,N_3969,N_3834);
nor U5928 (N_5928,N_3515,N_3416);
nand U5929 (N_5929,N_3869,N_3218);
xnor U5930 (N_5930,N_3752,N_3984);
and U5931 (N_5931,N_3901,N_3333);
nor U5932 (N_5932,N_4412,N_3628);
xor U5933 (N_5933,N_3480,N_3824);
and U5934 (N_5934,N_4055,N_3854);
nand U5935 (N_5935,N_3093,N_4284);
nand U5936 (N_5936,N_4319,N_3130);
or U5937 (N_5937,N_3956,N_3580);
or U5938 (N_5938,N_3486,N_3557);
nand U5939 (N_5939,N_3394,N_3077);
xnor U5940 (N_5940,N_4235,N_3145);
nor U5941 (N_5941,N_3547,N_3146);
or U5942 (N_5942,N_3244,N_4292);
nor U5943 (N_5943,N_4313,N_4307);
nand U5944 (N_5944,N_3025,N_4348);
and U5945 (N_5945,N_4234,N_4432);
xor U5946 (N_5946,N_3035,N_3701);
or U5947 (N_5947,N_3743,N_3062);
or U5948 (N_5948,N_4304,N_3251);
nor U5949 (N_5949,N_4003,N_3606);
nand U5950 (N_5950,N_3935,N_3960);
nand U5951 (N_5951,N_3367,N_4202);
nand U5952 (N_5952,N_4206,N_4370);
or U5953 (N_5953,N_3721,N_4174);
and U5954 (N_5954,N_3836,N_3710);
xnor U5955 (N_5955,N_3752,N_4038);
or U5956 (N_5956,N_3723,N_3807);
xor U5957 (N_5957,N_3575,N_4000);
nor U5958 (N_5958,N_3339,N_3271);
and U5959 (N_5959,N_3764,N_4433);
or U5960 (N_5960,N_4433,N_4256);
xnor U5961 (N_5961,N_4300,N_3037);
or U5962 (N_5962,N_3357,N_4153);
or U5963 (N_5963,N_4491,N_3755);
nor U5964 (N_5964,N_3559,N_3654);
nand U5965 (N_5965,N_4134,N_4218);
nand U5966 (N_5966,N_4396,N_3168);
and U5967 (N_5967,N_4200,N_3175);
or U5968 (N_5968,N_3340,N_3997);
or U5969 (N_5969,N_4435,N_3406);
nor U5970 (N_5970,N_3159,N_4157);
nor U5971 (N_5971,N_3726,N_3327);
or U5972 (N_5972,N_3704,N_4295);
and U5973 (N_5973,N_4309,N_3065);
nand U5974 (N_5974,N_3103,N_3764);
and U5975 (N_5975,N_3354,N_3610);
and U5976 (N_5976,N_3609,N_3605);
and U5977 (N_5977,N_3110,N_3089);
nand U5978 (N_5978,N_3361,N_3921);
nand U5979 (N_5979,N_3802,N_3984);
and U5980 (N_5980,N_3942,N_3302);
nor U5981 (N_5981,N_3575,N_3496);
and U5982 (N_5982,N_3848,N_4399);
or U5983 (N_5983,N_3642,N_3047);
xnor U5984 (N_5984,N_3424,N_3553);
xnor U5985 (N_5985,N_3858,N_3886);
or U5986 (N_5986,N_4043,N_3818);
or U5987 (N_5987,N_3323,N_3157);
nand U5988 (N_5988,N_3858,N_3745);
or U5989 (N_5989,N_4301,N_3054);
or U5990 (N_5990,N_4247,N_4263);
and U5991 (N_5991,N_3490,N_4029);
nand U5992 (N_5992,N_4420,N_4316);
or U5993 (N_5993,N_3803,N_3523);
nand U5994 (N_5994,N_3377,N_3263);
or U5995 (N_5995,N_3986,N_3047);
and U5996 (N_5996,N_3963,N_4180);
or U5997 (N_5997,N_3623,N_3307);
and U5998 (N_5998,N_3673,N_4407);
nor U5999 (N_5999,N_4213,N_3149);
nor U6000 (N_6000,N_4924,N_5436);
nand U6001 (N_6001,N_5690,N_5636);
nor U6002 (N_6002,N_5120,N_5352);
and U6003 (N_6003,N_5357,N_5629);
or U6004 (N_6004,N_4735,N_4827);
and U6005 (N_6005,N_4821,N_5347);
nand U6006 (N_6006,N_5465,N_5018);
nand U6007 (N_6007,N_5002,N_4739);
and U6008 (N_6008,N_5066,N_4622);
and U6009 (N_6009,N_5333,N_5976);
or U6010 (N_6010,N_5116,N_5965);
nor U6011 (N_6011,N_5878,N_4585);
and U6012 (N_6012,N_5140,N_5703);
nand U6013 (N_6013,N_5183,N_4526);
nor U6014 (N_6014,N_5454,N_5627);
nand U6015 (N_6015,N_5173,N_5893);
and U6016 (N_6016,N_5185,N_4772);
or U6017 (N_6017,N_5412,N_5594);
nor U6018 (N_6018,N_4665,N_4653);
and U6019 (N_6019,N_4696,N_4999);
nand U6020 (N_6020,N_5902,N_5962);
and U6021 (N_6021,N_5798,N_5907);
nor U6022 (N_6022,N_5157,N_5283);
xor U6023 (N_6023,N_5607,N_5030);
nor U6024 (N_6024,N_4859,N_5418);
and U6025 (N_6025,N_5348,N_5325);
and U6026 (N_6026,N_5067,N_4824);
nand U6027 (N_6027,N_4656,N_5133);
and U6028 (N_6028,N_5245,N_5788);
or U6029 (N_6029,N_5573,N_5318);
or U6030 (N_6030,N_4941,N_4955);
nand U6031 (N_6031,N_4841,N_4671);
nand U6032 (N_6032,N_5240,N_5933);
nor U6033 (N_6033,N_4576,N_5851);
xor U6034 (N_6034,N_5389,N_5857);
xnor U6035 (N_6035,N_4706,N_5153);
xor U6036 (N_6036,N_5166,N_4970);
or U6037 (N_6037,N_5138,N_4719);
xnor U6038 (N_6038,N_5428,N_4601);
or U6039 (N_6039,N_4915,N_5600);
nand U6040 (N_6040,N_5281,N_5984);
or U6041 (N_6041,N_4789,N_5992);
nor U6042 (N_6042,N_5795,N_5892);
and U6043 (N_6043,N_4853,N_5786);
or U6044 (N_6044,N_5403,N_4583);
nand U6045 (N_6045,N_4663,N_5450);
nor U6046 (N_6046,N_4618,N_5043);
nand U6047 (N_6047,N_4906,N_4595);
or U6048 (N_6048,N_5154,N_5186);
xor U6049 (N_6049,N_5731,N_5365);
or U6050 (N_6050,N_4549,N_4614);
nand U6051 (N_6051,N_4638,N_5622);
or U6052 (N_6052,N_4972,N_4582);
or U6053 (N_6053,N_5343,N_4947);
nand U6054 (N_6054,N_4515,N_5397);
or U6055 (N_6055,N_5394,N_5051);
nor U6056 (N_6056,N_4973,N_5496);
nor U6057 (N_6057,N_5306,N_5423);
nand U6058 (N_6058,N_4758,N_5220);
and U6059 (N_6059,N_5430,N_5815);
xnor U6060 (N_6060,N_5947,N_5083);
and U6061 (N_6061,N_5888,N_5257);
or U6062 (N_6062,N_5075,N_5275);
xor U6063 (N_6063,N_5168,N_4654);
nand U6064 (N_6064,N_5122,N_5085);
or U6065 (N_6065,N_5855,N_5970);
and U6066 (N_6066,N_5049,N_4991);
and U6067 (N_6067,N_4545,N_4554);
or U6068 (N_6068,N_5337,N_4863);
nand U6069 (N_6069,N_4651,N_4895);
nand U6070 (N_6070,N_5334,N_4943);
or U6071 (N_6071,N_4860,N_5784);
or U6072 (N_6072,N_5382,N_5648);
nand U6073 (N_6073,N_5442,N_5940);
nand U6074 (N_6074,N_5805,N_5112);
nand U6075 (N_6075,N_5799,N_5521);
and U6076 (N_6076,N_4976,N_5022);
or U6077 (N_6077,N_5929,N_4971);
and U6078 (N_6078,N_5835,N_5781);
nor U6079 (N_6079,N_5647,N_4996);
nor U6080 (N_6080,N_5399,N_5272);
and U6081 (N_6081,N_5820,N_5277);
nor U6082 (N_6082,N_5744,N_5726);
and U6083 (N_6083,N_5409,N_5144);
or U6084 (N_6084,N_4982,N_4746);
and U6085 (N_6085,N_5385,N_4801);
nand U6086 (N_6086,N_5814,N_5960);
and U6087 (N_6087,N_4988,N_4850);
and U6088 (N_6088,N_4676,N_5639);
or U6089 (N_6089,N_4517,N_4542);
nand U6090 (N_6090,N_5871,N_4535);
nor U6091 (N_6091,N_5364,N_4926);
and U6092 (N_6092,N_4751,N_5367);
and U6093 (N_6093,N_4786,N_5128);
or U6094 (N_6094,N_4954,N_4997);
nor U6095 (N_6095,N_5735,N_4537);
nand U6096 (N_6096,N_5803,N_5955);
nand U6097 (N_6097,N_5194,N_5342);
nand U6098 (N_6098,N_4810,N_5187);
nor U6099 (N_6099,N_5581,N_4717);
or U6100 (N_6100,N_5538,N_4512);
xnor U6101 (N_6101,N_5407,N_5303);
nand U6102 (N_6102,N_5826,N_5503);
nor U6103 (N_6103,N_5410,N_4538);
and U6104 (N_6104,N_4780,N_5130);
nor U6105 (N_6105,N_4686,N_4829);
or U6106 (N_6106,N_4889,N_4781);
nor U6107 (N_6107,N_5440,N_5501);
xnor U6108 (N_6108,N_5369,N_4811);
and U6109 (N_6109,N_5967,N_5966);
nand U6110 (N_6110,N_5628,N_4502);
nand U6111 (N_6111,N_5338,N_5926);
nand U6112 (N_6112,N_5139,N_5142);
and U6113 (N_6113,N_5613,N_5523);
xor U6114 (N_6114,N_4704,N_4787);
and U6115 (N_6115,N_4655,N_5322);
and U6116 (N_6116,N_5722,N_5730);
or U6117 (N_6117,N_5096,N_4870);
nand U6118 (N_6118,N_5679,N_5042);
or U6119 (N_6119,N_5807,N_5493);
and U6120 (N_6120,N_4547,N_5565);
nor U6121 (N_6121,N_5414,N_5961);
and U6122 (N_6122,N_5813,N_5003);
and U6123 (N_6123,N_5775,N_4925);
nand U6124 (N_6124,N_4743,N_4961);
nor U6125 (N_6125,N_4729,N_4530);
and U6126 (N_6126,N_4568,N_5525);
and U6127 (N_6127,N_5356,N_5330);
nand U6128 (N_6128,N_4581,N_5585);
nor U6129 (N_6129,N_5270,N_5274);
nand U6130 (N_6130,N_4892,N_5649);
nand U6131 (N_6131,N_5780,N_5809);
nand U6132 (N_6132,N_5542,N_4580);
nand U6133 (N_6133,N_5502,N_4843);
or U6134 (N_6134,N_5045,N_5904);
nand U6135 (N_6135,N_5368,N_4837);
and U6136 (N_6136,N_4833,N_4513);
or U6137 (N_6137,N_4596,N_4744);
or U6138 (N_6138,N_5172,N_4510);
nand U6139 (N_6139,N_5297,N_5101);
or U6140 (N_6140,N_4886,N_4817);
and U6141 (N_6141,N_5611,N_5812);
and U6142 (N_6142,N_5526,N_4528);
nand U6143 (N_6143,N_5971,N_4505);
nand U6144 (N_6144,N_5919,N_5181);
or U6145 (N_6145,N_5569,N_5623);
or U6146 (N_6146,N_5259,N_5329);
and U6147 (N_6147,N_5602,N_5323);
and U6148 (N_6148,N_5125,N_4957);
nand U6149 (N_6149,N_5842,N_5863);
and U6150 (N_6150,N_5055,N_5008);
nor U6151 (N_6151,N_4808,N_5559);
or U6152 (N_6152,N_4534,N_5106);
and U6153 (N_6153,N_5054,N_5527);
xnor U6154 (N_6154,N_4936,N_5141);
or U6155 (N_6155,N_5062,N_4983);
nor U6156 (N_6156,N_5201,N_5883);
nor U6157 (N_6157,N_4600,N_5882);
and U6158 (N_6158,N_4894,N_4834);
nor U6159 (N_6159,N_5988,N_5715);
nor U6160 (N_6160,N_4763,N_5574);
and U6161 (N_6161,N_5561,N_5529);
or U6162 (N_6162,N_5664,N_5249);
or U6163 (N_6163,N_5875,N_5353);
nor U6164 (N_6164,N_5531,N_5912);
nand U6165 (N_6165,N_5519,N_5408);
nand U6166 (N_6166,N_4927,N_5522);
xnor U6167 (N_6167,N_4883,N_5858);
or U6168 (N_6168,N_4873,N_5876);
xor U6169 (N_6169,N_5152,N_4847);
or U6170 (N_6170,N_5189,N_4571);
and U6171 (N_6171,N_5472,N_5650);
nor U6172 (N_6172,N_4586,N_5089);
nand U6173 (N_6173,N_4902,N_4670);
xnor U6174 (N_6174,N_5244,N_5760);
nor U6175 (N_6175,N_5006,N_5580);
or U6176 (N_6176,N_5068,N_5630);
or U6177 (N_6177,N_4501,N_5366);
nor U6178 (N_6178,N_5891,N_5248);
or U6179 (N_6179,N_5453,N_5834);
or U6180 (N_6180,N_5918,N_4774);
nor U6181 (N_6181,N_5791,N_5593);
and U6182 (N_6182,N_4525,N_4740);
and U6183 (N_6183,N_5900,N_5642);
and U6184 (N_6184,N_4575,N_4572);
nor U6185 (N_6185,N_5738,N_5102);
and U6186 (N_6186,N_4745,N_5591);
nand U6187 (N_6187,N_5354,N_5767);
and U6188 (N_6188,N_5056,N_5041);
nand U6189 (N_6189,N_5090,N_4711);
or U6190 (N_6190,N_5945,N_5806);
nor U6191 (N_6191,N_4881,N_5737);
nor U6192 (N_6192,N_5708,N_4627);
nand U6193 (N_6193,N_4845,N_5824);
or U6194 (N_6194,N_5897,N_5914);
nand U6195 (N_6195,N_5683,N_4669);
or U6196 (N_6196,N_4564,N_5321);
or U6197 (N_6197,N_4519,N_5156);
nor U6198 (N_6198,N_5686,N_5804);
nor U6199 (N_6199,N_5175,N_4977);
and U6200 (N_6200,N_5656,N_4802);
nor U6201 (N_6201,N_5584,N_4604);
nor U6202 (N_6202,N_4675,N_4911);
nand U6203 (N_6203,N_5980,N_5073);
or U6204 (N_6204,N_4862,N_4963);
and U6205 (N_6205,N_5692,N_4923);
or U6206 (N_6206,N_5400,N_5727);
nor U6207 (N_6207,N_5047,N_4796);
nand U6208 (N_6208,N_5011,N_5115);
nand U6209 (N_6209,N_4668,N_4685);
or U6210 (N_6210,N_4979,N_5905);
nand U6211 (N_6211,N_5015,N_5605);
nand U6212 (N_6212,N_5202,N_4569);
nor U6213 (N_6213,N_4650,N_4708);
nand U6214 (N_6214,N_4967,N_4523);
and U6215 (N_6215,N_4728,N_4921);
and U6216 (N_6216,N_5570,N_5590);
or U6217 (N_6217,N_5467,N_4854);
nor U6218 (N_6218,N_5586,N_4855);
nor U6219 (N_6219,N_4590,N_5147);
nand U6220 (N_6220,N_5359,N_4705);
and U6221 (N_6221,N_5084,N_5608);
nor U6222 (N_6222,N_5361,N_5852);
nand U6223 (N_6223,N_5749,N_5494);
or U6224 (N_6224,N_5668,N_4541);
nand U6225 (N_6225,N_5770,N_5982);
xor U6226 (N_6226,N_5064,N_4664);
and U6227 (N_6227,N_5217,N_4775);
nand U6228 (N_6228,N_4964,N_4688);
nor U6229 (N_6229,N_5801,N_5719);
nand U6230 (N_6230,N_5524,N_4874);
nor U6231 (N_6231,N_4896,N_5732);
and U6232 (N_6232,N_5200,N_5118);
nor U6233 (N_6233,N_5010,N_5014);
nand U6234 (N_6234,N_5930,N_4840);
xnor U6235 (N_6235,N_5360,N_4691);
nor U6236 (N_6236,N_5178,N_4956);
nor U6237 (N_6237,N_4898,N_4805);
nand U6238 (N_6238,N_4509,N_5645);
and U6239 (N_6239,N_4531,N_4648);
nor U6240 (N_6240,N_5298,N_4624);
and U6241 (N_6241,N_5922,N_5093);
and U6242 (N_6242,N_5340,N_5293);
xnor U6243 (N_6243,N_4507,N_4905);
xor U6244 (N_6244,N_5953,N_5633);
nor U6245 (N_6245,N_4912,N_5913);
or U6246 (N_6246,N_4842,N_4642);
nor U6247 (N_6247,N_5950,N_5381);
nor U6248 (N_6248,N_4752,N_5934);
xor U6249 (N_6249,N_5983,N_5192);
nand U6250 (N_6250,N_5616,N_4969);
nand U6251 (N_6251,N_5682,N_5597);
and U6252 (N_6252,N_5477,N_4804);
or U6253 (N_6253,N_5550,N_5512);
nand U6254 (N_6254,N_5673,N_5239);
and U6255 (N_6255,N_4734,N_4560);
and U6256 (N_6256,N_5854,N_5225);
nand U6257 (N_6257,N_4563,N_5520);
nor U6258 (N_6258,N_5371,N_5489);
and U6259 (N_6259,N_5718,N_4871);
nor U6260 (N_6260,N_5571,N_4754);
nor U6261 (N_6261,N_5449,N_5458);
or U6262 (N_6262,N_4682,N_4949);
or U6263 (N_6263,N_4684,N_5743);
or U6264 (N_6264,N_5320,N_4712);
nand U6265 (N_6265,N_5537,N_5541);
xnor U6266 (N_6266,N_5660,N_5474);
or U6267 (N_6267,N_5242,N_4965);
nor U6268 (N_6268,N_5941,N_5704);
nand U6269 (N_6269,N_4672,N_4681);
nor U6270 (N_6270,N_4861,N_4904);
nand U6271 (N_6271,N_4613,N_5326);
nand U6272 (N_6272,N_5562,N_5059);
and U6273 (N_6273,N_4985,N_5507);
and U6274 (N_6274,N_5310,N_5532);
and U6275 (N_6275,N_5091,N_5880);
or U6276 (N_6276,N_5100,N_4768);
nand U6277 (N_6277,N_5994,N_5032);
nor U6278 (N_6278,N_4832,N_4720);
nor U6279 (N_6279,N_4931,N_5355);
nor U6280 (N_6280,N_5794,N_5747);
xor U6281 (N_6281,N_4918,N_4723);
nor U6282 (N_6282,N_4929,N_4646);
or U6283 (N_6283,N_5251,N_4631);
nor U6284 (N_6284,N_5688,N_4749);
nor U6285 (N_6285,N_5517,N_4968);
nand U6286 (N_6286,N_5495,N_5990);
and U6287 (N_6287,N_4984,N_4643);
xor U6288 (N_6288,N_5335,N_5536);
and U6289 (N_6289,N_4913,N_5071);
and U6290 (N_6290,N_4553,N_4959);
or U6291 (N_6291,N_5697,N_5533);
and U6292 (N_6292,N_5241,N_5237);
nand U6293 (N_6293,N_4594,N_4556);
nor U6294 (N_6294,N_5074,N_5161);
xor U6295 (N_6295,N_5973,N_5634);
nor U6296 (N_6296,N_5210,N_5752);
nor U6297 (N_6297,N_5438,N_5013);
xor U6298 (N_6298,N_5619,N_5906);
or U6299 (N_6299,N_5651,N_5425);
nand U6300 (N_6300,N_4699,N_5817);
or U6301 (N_6301,N_5105,N_5386);
nand U6302 (N_6302,N_5534,N_5946);
nor U6303 (N_6303,N_5596,N_4753);
nor U6304 (N_6304,N_4989,N_5921);
nor U6305 (N_6305,N_5687,N_4701);
nand U6306 (N_6306,N_4544,N_4514);
nand U6307 (N_6307,N_5543,N_4818);
and U6308 (N_6308,N_4522,N_5702);
or U6309 (N_6309,N_5564,N_5848);
and U6310 (N_6310,N_5927,N_5491);
nand U6311 (N_6311,N_5721,N_4756);
and U6312 (N_6312,N_5016,N_5300);
xnor U6313 (N_6313,N_5264,N_5589);
nor U6314 (N_6314,N_5741,N_4962);
nor U6315 (N_6315,N_4659,N_4605);
nand U6316 (N_6316,N_5107,N_4707);
xor U6317 (N_6317,N_5868,N_5755);
xor U6318 (N_6318,N_5195,N_4597);
nor U6319 (N_6319,N_5680,N_5592);
nor U6320 (N_6320,N_4748,N_5579);
or U6321 (N_6321,N_4782,N_4606);
or U6322 (N_6322,N_5802,N_5705);
xor U6323 (N_6323,N_5513,N_4848);
nand U6324 (N_6324,N_5317,N_5345);
or U6325 (N_6325,N_5557,N_5873);
nand U6326 (N_6326,N_4966,N_4567);
nand U6327 (N_6327,N_4950,N_5291);
or U6328 (N_6328,N_5516,N_5475);
xor U6329 (N_6329,N_5215,N_4865);
and U6330 (N_6330,N_4867,N_5974);
or U6331 (N_6331,N_4697,N_5424);
nand U6332 (N_6332,N_5218,N_5065);
nor U6333 (N_6333,N_4689,N_5968);
xnor U6334 (N_6334,N_4875,N_4718);
xnor U6335 (N_6335,N_4673,N_5724);
and U6336 (N_6336,N_4809,N_5838);
nand U6337 (N_6337,N_5545,N_5977);
nand U6338 (N_6338,N_5626,N_5208);
nand U6339 (N_6339,N_4790,N_5793);
or U6340 (N_6340,N_5243,N_5388);
nor U6341 (N_6341,N_5080,N_5265);
xor U6342 (N_6342,N_5952,N_5832);
nand U6343 (N_6343,N_4511,N_5991);
or U6344 (N_6344,N_4900,N_5553);
and U6345 (N_6345,N_4884,N_4795);
nand U6346 (N_6346,N_4932,N_5928);
or U6347 (N_6347,N_5989,N_5746);
nand U6348 (N_6348,N_5742,N_5774);
and U6349 (N_6349,N_4558,N_5836);
or U6350 (N_6350,N_5695,N_4897);
or U6351 (N_6351,N_5375,N_5641);
or U6352 (N_6352,N_4917,N_4727);
nand U6353 (N_6353,N_5999,N_5253);
nor U6354 (N_6354,N_4798,N_5479);
or U6355 (N_6355,N_5700,N_5728);
nand U6356 (N_6356,N_5769,N_5279);
xor U6357 (N_6357,N_4760,N_5844);
nor U6358 (N_6358,N_5177,N_4557);
xnor U6359 (N_6359,N_5850,N_4777);
or U6360 (N_6360,N_5869,N_4693);
and U6361 (N_6361,N_5123,N_4658);
nor U6362 (N_6362,N_4639,N_5510);
nand U6363 (N_6363,N_5483,N_5609);
nor U6364 (N_6364,N_5095,N_5540);
or U6365 (N_6365,N_4539,N_4715);
nor U6366 (N_6366,N_4724,N_5575);
or U6367 (N_6367,N_5987,N_5435);
and U6368 (N_6368,N_5829,N_4910);
xor U6369 (N_6369,N_4611,N_5745);
and U6370 (N_6370,N_5124,N_5572);
and U6371 (N_6371,N_4791,N_4617);
and U6372 (N_6372,N_5768,N_4820);
nand U6373 (N_6373,N_5459,N_4687);
nand U6374 (N_6374,N_4822,N_5577);
and U6375 (N_6375,N_5547,N_5757);
xnor U6376 (N_6376,N_5380,N_4540);
nor U6377 (N_6377,N_5576,N_4879);
nor U6378 (N_6378,N_5363,N_5797);
nor U6379 (N_6379,N_4793,N_5840);
and U6380 (N_6380,N_4641,N_4920);
nand U6381 (N_6381,N_5406,N_5886);
and U6382 (N_6382,N_5415,N_5484);
nor U6383 (N_6383,N_5916,N_4703);
nand U6384 (N_6384,N_5772,N_5614);
xnor U6385 (N_6385,N_4766,N_5909);
and U6386 (N_6386,N_5088,N_5699);
xor U6387 (N_6387,N_5170,N_4958);
xnor U6388 (N_6388,N_5870,N_5402);
and U6389 (N_6389,N_5563,N_4937);
xor U6390 (N_6390,N_5923,N_4771);
and U6391 (N_6391,N_5482,N_5127);
nand U6392 (N_6392,N_5765,N_4978);
and U6393 (N_6393,N_4593,N_5944);
and U6394 (N_6394,N_5587,N_5263);
and U6395 (N_6395,N_5694,N_4635);
and U6396 (N_6396,N_5932,N_5789);
nand U6397 (N_6397,N_5485,N_5227);
nor U6398 (N_6398,N_5885,N_5787);
and U6399 (N_6399,N_5693,N_4647);
xor U6400 (N_6400,N_4946,N_5404);
and U6401 (N_6401,N_5480,N_5956);
nand U6402 (N_6402,N_5669,N_5969);
nand U6403 (N_6403,N_4713,N_4661);
or U6404 (N_6404,N_5996,N_5504);
or U6405 (N_6405,N_5129,N_4797);
nand U6406 (N_6406,N_5098,N_4710);
nor U6407 (N_6407,N_5206,N_5332);
and U6408 (N_6408,N_5691,N_5924);
nor U6409 (N_6409,N_5295,N_5327);
nand U6410 (N_6410,N_5384,N_4858);
and U6411 (N_6411,N_4573,N_5289);
nor U6412 (N_6412,N_5164,N_5285);
or U6413 (N_6413,N_5763,N_5552);
xnor U6414 (N_6414,N_4868,N_5224);
and U6415 (N_6415,N_4799,N_5935);
nor U6416 (N_6416,N_5292,N_5535);
and U6417 (N_6417,N_5009,N_5908);
nor U6418 (N_6418,N_5723,N_5060);
nor U6419 (N_6419,N_4807,N_4527);
or U6420 (N_6420,N_4919,N_5050);
nor U6421 (N_6421,N_5603,N_4750);
xnor U6422 (N_6422,N_4998,N_5392);
nand U6423 (N_6423,N_4599,N_5448);
or U6424 (N_6424,N_5081,N_5612);
xnor U6425 (N_6425,N_5837,N_5655);
and U6426 (N_6426,N_4764,N_5346);
or U6427 (N_6427,N_5024,N_5460);
nand U6428 (N_6428,N_5136,N_5667);
or U6429 (N_6429,N_4993,N_5387);
or U6430 (N_6430,N_4776,N_5548);
xnor U6431 (N_6431,N_5443,N_5461);
or U6432 (N_6432,N_5758,N_5676);
nor U6433 (N_6433,N_5720,N_4944);
or U6434 (N_6434,N_4636,N_5750);
or U6435 (N_6435,N_5761,N_4826);
or U6436 (N_6436,N_5427,N_5733);
or U6437 (N_6437,N_5311,N_4767);
nor U6438 (N_6438,N_5920,N_4588);
xnor U6439 (N_6439,N_5997,N_5350);
and U6440 (N_6440,N_5094,N_5915);
and U6441 (N_6441,N_4662,N_5282);
nor U6442 (N_6442,N_4633,N_5092);
nand U6443 (N_6443,N_5273,N_5864);
nor U6444 (N_6444,N_5505,N_5811);
or U6445 (N_6445,N_5665,N_4788);
nor U6446 (N_6446,N_5294,N_5549);
or U6447 (N_6447,N_4695,N_5426);
nor U6448 (N_6448,N_5963,N_4922);
nor U6449 (N_6449,N_5268,N_5511);
or U6450 (N_6450,N_4851,N_4629);
nor U6451 (N_6451,N_5033,N_4813);
or U6452 (N_6452,N_5391,N_4762);
nor U6453 (N_6453,N_5146,N_5250);
or U6454 (N_6454,N_5822,N_5238);
nor U6455 (N_6455,N_5646,N_5119);
or U6456 (N_6456,N_5452,N_4570);
nand U6457 (N_6457,N_4935,N_5663);
and U6458 (N_6458,N_5213,N_5978);
and U6459 (N_6459,N_5198,N_5005);
or U6460 (N_6460,N_4856,N_5260);
nor U6461 (N_6461,N_5276,N_4846);
nor U6462 (N_6462,N_5556,N_5712);
nor U6463 (N_6463,N_5903,N_5027);
or U6464 (N_6464,N_5508,N_4616);
xor U6465 (N_6465,N_5211,N_5939);
or U6466 (N_6466,N_5618,N_5578);
or U6467 (N_6467,N_5221,N_5284);
and U6468 (N_6468,N_4852,N_4891);
nor U6469 (N_6469,N_5860,N_4869);
and U6470 (N_6470,N_5302,N_5286);
nand U6471 (N_6471,N_5530,N_5349);
nand U6472 (N_6472,N_5895,N_4566);
or U6473 (N_6473,N_4652,N_5190);
nand U6474 (N_6474,N_5143,N_4714);
nand U6475 (N_6475,N_5995,N_5445);
or U6476 (N_6476,N_4960,N_5267);
or U6477 (N_6477,N_4736,N_5214);
nor U6478 (N_6478,N_5894,N_5470);
nor U6479 (N_6479,N_5204,N_5176);
and U6480 (N_6480,N_5038,N_4814);
nor U6481 (N_6481,N_5782,N_5203);
nor U6482 (N_6482,N_5653,N_5847);
nor U6483 (N_6483,N_4546,N_5823);
nand U6484 (N_6484,N_4678,N_5979);
and U6485 (N_6485,N_5631,N_5053);
and U6486 (N_6486,N_5299,N_5643);
nand U6487 (N_6487,N_5437,N_5658);
nor U6488 (N_6488,N_4579,N_4737);
xnor U6489 (N_6489,N_5149,N_5236);
nand U6490 (N_6490,N_5019,N_5471);
and U6491 (N_6491,N_5061,N_4612);
nor U6492 (N_6492,N_5827,N_5601);
or U6493 (N_6493,N_5785,N_5684);
and U6494 (N_6494,N_5598,N_4857);
nor U6495 (N_6495,N_5207,N_5839);
nor U6496 (N_6496,N_5887,N_5810);
nand U6497 (N_6497,N_4907,N_4640);
nor U6498 (N_6498,N_5393,N_5677);
nor U6499 (N_6499,N_5476,N_5280);
nand U6500 (N_6500,N_5981,N_5487);
nor U6501 (N_6501,N_5351,N_4940);
or U6502 (N_6502,N_4503,N_5539);
nor U6503 (N_6503,N_5457,N_5943);
nor U6504 (N_6504,N_5833,N_4504);
nand U6505 (N_6505,N_5959,N_5985);
nor U6506 (N_6506,N_5439,N_5148);
nor U6507 (N_6507,N_5287,N_4533);
or U6508 (N_6508,N_4598,N_5498);
nand U6509 (N_6509,N_5163,N_4864);
nand U6510 (N_6510,N_5751,N_5948);
nand U6511 (N_6511,N_5158,N_4903);
nor U6512 (N_6512,N_5954,N_5222);
or U6513 (N_6513,N_5174,N_4939);
nor U6514 (N_6514,N_5271,N_4690);
nand U6515 (N_6515,N_5278,N_5017);
xor U6516 (N_6516,N_5862,N_4757);
xor U6517 (N_6517,N_4830,N_5023);
nand U6518 (N_6518,N_5396,N_4942);
and U6519 (N_6519,N_4784,N_4823);
nand U6520 (N_6520,N_4849,N_5754);
xor U6521 (N_6521,N_5313,N_5319);
nand U6522 (N_6522,N_5421,N_5499);
nor U6523 (N_6523,N_5429,N_5012);
nor U6524 (N_6524,N_5736,N_4644);
nand U6525 (N_6525,N_4794,N_5254);
nor U6526 (N_6526,N_4778,N_5086);
nor U6527 (N_6527,N_4574,N_4901);
xnor U6528 (N_6528,N_5020,N_5191);
nand U6529 (N_6529,N_4608,N_5219);
nor U6530 (N_6530,N_5776,N_4765);
or U6531 (N_6531,N_5000,N_5235);
and U6532 (N_6532,N_4628,N_4700);
xnor U6533 (N_6533,N_4773,N_5604);
or U6534 (N_6534,N_5740,N_5644);
and U6535 (N_6535,N_5606,N_5420);
xor U6536 (N_6536,N_5867,N_4819);
nand U6537 (N_6537,N_4785,N_5304);
nand U6538 (N_6538,N_5753,N_4559);
and U6539 (N_6539,N_5942,N_5707);
xnor U6540 (N_6540,N_4742,N_4521);
and U6541 (N_6541,N_5566,N_5104);
nand U6542 (N_6542,N_5167,N_4645);
or U6543 (N_6543,N_5696,N_5159);
or U6544 (N_6544,N_5975,N_4592);
and U6545 (N_6545,N_4938,N_5560);
or U6546 (N_6546,N_4816,N_5151);
and U6547 (N_6547,N_4591,N_5205);
or U6548 (N_6548,N_5790,N_5567);
or U6549 (N_6549,N_5040,N_5938);
nand U6550 (N_6550,N_5121,N_4888);
or U6551 (N_6551,N_5082,N_5180);
nand U6552 (N_6552,N_5621,N_5884);
and U6553 (N_6553,N_5145,N_5481);
or U6554 (N_6554,N_5662,N_5232);
and U6555 (N_6555,N_5678,N_5773);
or U6556 (N_6556,N_5230,N_4520);
nor U6557 (N_6557,N_5113,N_5659);
or U6558 (N_6558,N_5028,N_5711);
or U6559 (N_6559,N_5312,N_5717);
xnor U6560 (N_6560,N_4885,N_5052);
nand U6561 (N_6561,N_5037,N_4880);
and U6562 (N_6562,N_5544,N_4709);
xor U6563 (N_6563,N_5137,N_5898);
nand U6564 (N_6564,N_5258,N_5110);
nor U6565 (N_6565,N_5057,N_5555);
nand U6566 (N_6566,N_4621,N_5077);
xor U6567 (N_6567,N_4887,N_5890);
and U6568 (N_6568,N_4725,N_4952);
nand U6569 (N_6569,N_5097,N_5433);
or U6570 (N_6570,N_5554,N_4508);
nor U6571 (N_6571,N_5039,N_5255);
xnor U6572 (N_6572,N_5395,N_4987);
nand U6573 (N_6573,N_5308,N_4550);
and U6574 (N_6574,N_4994,N_5689);
nand U6575 (N_6575,N_4619,N_4721);
nor U6576 (N_6576,N_5949,N_5706);
or U6577 (N_6577,N_5331,N_5464);
and U6578 (N_6578,N_5374,N_4930);
and U6579 (N_6579,N_5288,N_5160);
or U6580 (N_6580,N_4666,N_5290);
or U6581 (N_6581,N_5079,N_5800);
nor U6582 (N_6582,N_5500,N_5972);
or U6583 (N_6583,N_4948,N_5131);
or U6584 (N_6584,N_5640,N_5411);
or U6585 (N_6585,N_5226,N_4634);
nand U6586 (N_6586,N_4928,N_4914);
xor U6587 (N_6587,N_4683,N_5182);
nand U6588 (N_6588,N_4909,N_5764);
or U6589 (N_6589,N_5796,N_5262);
xor U6590 (N_6590,N_4899,N_4610);
xor U6591 (N_6591,N_5951,N_5468);
nand U6592 (N_6592,N_4561,N_5212);
and U6593 (N_6593,N_4716,N_4732);
and U6594 (N_6594,N_5007,N_4838);
and U6595 (N_6595,N_4995,N_5625);
nor U6596 (N_6596,N_5911,N_5674);
and U6597 (N_6597,N_5638,N_5506);
nor U6598 (N_6598,N_4677,N_4980);
and U6599 (N_6599,N_5216,N_5048);
or U6600 (N_6600,N_4518,N_5199);
or U6601 (N_6601,N_4882,N_4529);
xnor U6602 (N_6602,N_4945,N_4698);
and U6603 (N_6603,N_4702,N_5432);
nor U6604 (N_6604,N_5766,N_5087);
and U6605 (N_6605,N_5324,N_4615);
and U6606 (N_6606,N_5756,N_5316);
or U6607 (N_6607,N_5026,N_5617);
nand U6608 (N_6608,N_5405,N_5431);
nand U6609 (N_6609,N_5383,N_5378);
nand U6610 (N_6610,N_4609,N_4674);
and U6611 (N_6611,N_5229,N_5046);
or U6612 (N_6612,N_5599,N_4625);
nand U6613 (N_6613,N_5734,N_5463);
nor U6614 (N_6614,N_4679,N_5269);
or U6615 (N_6615,N_5296,N_5469);
nand U6616 (N_6616,N_5473,N_5193);
nand U6617 (N_6617,N_5358,N_4836);
or U6618 (N_6618,N_5710,N_4524);
or U6619 (N_6619,N_5114,N_5486);
and U6620 (N_6620,N_5256,N_4500);
nand U6621 (N_6621,N_4548,N_4792);
nand U6622 (N_6622,N_5309,N_5035);
or U6623 (N_6623,N_5362,N_5725);
or U6624 (N_6624,N_5896,N_5964);
and U6625 (N_6625,N_5624,N_4831);
nor U6626 (N_6626,N_5398,N_5266);
nor U6627 (N_6627,N_5029,N_5135);
nor U6628 (N_6628,N_4532,N_4872);
nor U6629 (N_6629,N_5551,N_4908);
and U6630 (N_6630,N_4825,N_5936);
or U6631 (N_6631,N_5654,N_5004);
nor U6632 (N_6632,N_5716,N_5762);
nor U6633 (N_6633,N_4878,N_5126);
nor U6634 (N_6634,N_5681,N_5390);
and U6635 (N_6635,N_4761,N_5830);
and U6636 (N_6636,N_5488,N_5261);
and U6637 (N_6637,N_5998,N_5841);
nand U6638 (N_6638,N_5492,N_5377);
nor U6639 (N_6639,N_5117,N_5610);
nand U6640 (N_6640,N_5957,N_5635);
and U6641 (N_6641,N_5413,N_5314);
nor U6642 (N_6642,N_5441,N_5165);
nand U6643 (N_6643,N_5620,N_4516);
nand U6644 (N_6644,N_5076,N_5179);
nand U6645 (N_6645,N_4632,N_5671);
xnor U6646 (N_6646,N_4990,N_4660);
or U6647 (N_6647,N_5134,N_5456);
nor U6648 (N_6648,N_5373,N_5771);
xnor U6649 (N_6649,N_5958,N_5184);
nor U6650 (N_6650,N_5058,N_4779);
nand U6651 (N_6651,N_5209,N_4551);
nor U6652 (N_6652,N_5582,N_5595);
and U6653 (N_6653,N_4876,N_5874);
or U6654 (N_6654,N_5111,N_5370);
and U6655 (N_6655,N_5307,N_5821);
nor U6656 (N_6656,N_4806,N_4741);
xnor U6657 (N_6657,N_4726,N_5034);
nor U6658 (N_6658,N_5714,N_5070);
nand U6659 (N_6659,N_4733,N_5759);
nor U6660 (N_6660,N_4890,N_4844);
or U6661 (N_6661,N_5701,N_4620);
nor U6662 (N_6662,N_4589,N_5879);
and U6663 (N_6663,N_5344,N_5231);
and U6664 (N_6664,N_4934,N_4694);
or U6665 (N_6665,N_4747,N_5831);
xor U6666 (N_6666,N_5247,N_5881);
and U6667 (N_6667,N_4828,N_5478);
nor U6668 (N_6668,N_5818,N_5889);
nor U6669 (N_6669,N_5661,N_5986);
or U6670 (N_6670,N_5108,N_5025);
nand U6671 (N_6671,N_5583,N_5069);
and U6672 (N_6672,N_4584,N_5422);
or U6673 (N_6673,N_4578,N_5078);
or U6674 (N_6674,N_4770,N_5861);
or U6675 (N_6675,N_5588,N_5568);
or U6676 (N_6676,N_4552,N_4587);
xor U6677 (N_6677,N_5808,N_4769);
and U6678 (N_6678,N_5021,N_4543);
or U6679 (N_6679,N_5099,N_5937);
nand U6680 (N_6680,N_4893,N_5865);
nor U6681 (N_6681,N_4835,N_5828);
or U6682 (N_6682,N_4536,N_5917);
nand U6683 (N_6683,N_5223,N_5509);
nand U6684 (N_6684,N_5859,N_5171);
or U6685 (N_6685,N_5376,N_5637);
nor U6686 (N_6686,N_5899,N_4839);
nand U6687 (N_6687,N_5072,N_5196);
nor U6688 (N_6688,N_4951,N_5853);
and U6689 (N_6689,N_4630,N_5063);
nand U6690 (N_6690,N_5849,N_5709);
or U6691 (N_6691,N_5528,N_5546);
nand U6692 (N_6692,N_5109,N_4602);
nor U6693 (N_6693,N_5518,N_5856);
xnor U6694 (N_6694,N_4812,N_5328);
nand U6695 (N_6695,N_5558,N_5514);
nor U6696 (N_6696,N_4974,N_5825);
nor U6697 (N_6697,N_4603,N_5417);
and U6698 (N_6698,N_5490,N_4986);
and U6699 (N_6699,N_5031,N_5729);
and U6700 (N_6700,N_4649,N_5672);
nand U6701 (N_6701,N_4953,N_5315);
nand U6702 (N_6702,N_5845,N_5675);
and U6703 (N_6703,N_4657,N_5401);
nor U6704 (N_6704,N_5748,N_5462);
nor U6705 (N_6705,N_5816,N_5103);
nand U6706 (N_6706,N_5843,N_5372);
nor U6707 (N_6707,N_5233,N_5713);
and U6708 (N_6708,N_4623,N_5779);
nand U6709 (N_6709,N_5783,N_5925);
nor U6710 (N_6710,N_5305,N_4755);
nand U6711 (N_6711,N_4680,N_4506);
nor U6712 (N_6712,N_5234,N_4692);
nand U6713 (N_6713,N_5447,N_4800);
and U6714 (N_6714,N_4916,N_5993);
and U6715 (N_6715,N_4607,N_4738);
or U6716 (N_6716,N_5657,N_5455);
and U6717 (N_6717,N_4866,N_5044);
xor U6718 (N_6718,N_5652,N_5777);
or U6719 (N_6719,N_5670,N_4783);
or U6720 (N_6720,N_5819,N_4730);
and U6721 (N_6721,N_5778,N_5872);
or U6722 (N_6722,N_5632,N_5197);
or U6723 (N_6723,N_5901,N_4555);
nor U6724 (N_6724,N_4803,N_5379);
nor U6725 (N_6725,N_5446,N_4981);
or U6726 (N_6726,N_5336,N_5615);
or U6727 (N_6727,N_5132,N_5910);
and U6728 (N_6728,N_5252,N_5846);
nand U6729 (N_6729,N_4992,N_4565);
nor U6730 (N_6730,N_4877,N_5877);
nand U6731 (N_6731,N_4562,N_4667);
nor U6732 (N_6732,N_4975,N_5866);
nor U6733 (N_6733,N_5419,N_5150);
xor U6734 (N_6734,N_5444,N_5931);
nand U6735 (N_6735,N_5792,N_4626);
nor U6736 (N_6736,N_5434,N_5466);
nand U6737 (N_6737,N_5228,N_4759);
xnor U6738 (N_6738,N_5515,N_5739);
and U6739 (N_6739,N_4933,N_5155);
nor U6740 (N_6740,N_5188,N_5339);
xor U6741 (N_6741,N_5497,N_4722);
nand U6742 (N_6742,N_5169,N_5666);
xor U6743 (N_6743,N_4815,N_5341);
nand U6744 (N_6744,N_4577,N_5416);
nor U6745 (N_6745,N_4731,N_4637);
or U6746 (N_6746,N_5036,N_5451);
or U6747 (N_6747,N_5685,N_5001);
nor U6748 (N_6748,N_5246,N_5698);
nand U6749 (N_6749,N_5301,N_5162);
nor U6750 (N_6750,N_5644,N_5110);
or U6751 (N_6751,N_5443,N_4969);
nand U6752 (N_6752,N_4623,N_4900);
or U6753 (N_6753,N_5040,N_5816);
nand U6754 (N_6754,N_5619,N_4560);
or U6755 (N_6755,N_5584,N_4647);
or U6756 (N_6756,N_4819,N_4712);
nor U6757 (N_6757,N_5273,N_5410);
or U6758 (N_6758,N_5235,N_5878);
and U6759 (N_6759,N_5234,N_4795);
nor U6760 (N_6760,N_5547,N_5820);
nor U6761 (N_6761,N_4812,N_5453);
or U6762 (N_6762,N_4897,N_4688);
xnor U6763 (N_6763,N_4952,N_5412);
xnor U6764 (N_6764,N_5225,N_5985);
nand U6765 (N_6765,N_5633,N_5207);
nand U6766 (N_6766,N_5277,N_4879);
nand U6767 (N_6767,N_4903,N_4661);
nor U6768 (N_6768,N_5292,N_5690);
nor U6769 (N_6769,N_4834,N_4753);
or U6770 (N_6770,N_4666,N_5447);
and U6771 (N_6771,N_5145,N_4931);
and U6772 (N_6772,N_4888,N_4667);
xnor U6773 (N_6773,N_4725,N_5080);
and U6774 (N_6774,N_5119,N_4854);
nand U6775 (N_6775,N_5475,N_5777);
nor U6776 (N_6776,N_5421,N_5556);
or U6777 (N_6777,N_5479,N_4944);
xnor U6778 (N_6778,N_5613,N_5641);
nand U6779 (N_6779,N_4763,N_4583);
nand U6780 (N_6780,N_4764,N_5382);
xnor U6781 (N_6781,N_4883,N_5618);
and U6782 (N_6782,N_5405,N_5748);
and U6783 (N_6783,N_4696,N_4983);
nor U6784 (N_6784,N_5165,N_5941);
nand U6785 (N_6785,N_4675,N_5569);
nand U6786 (N_6786,N_4791,N_5114);
and U6787 (N_6787,N_5252,N_5996);
and U6788 (N_6788,N_4781,N_4807);
or U6789 (N_6789,N_4666,N_5952);
nand U6790 (N_6790,N_5698,N_5534);
xor U6791 (N_6791,N_5126,N_5332);
and U6792 (N_6792,N_5804,N_5139);
xor U6793 (N_6793,N_5123,N_4918);
and U6794 (N_6794,N_4963,N_5676);
and U6795 (N_6795,N_4525,N_5854);
xor U6796 (N_6796,N_5070,N_5317);
and U6797 (N_6797,N_5120,N_5634);
nand U6798 (N_6798,N_4633,N_5382);
nand U6799 (N_6799,N_4664,N_5075);
nand U6800 (N_6800,N_5694,N_5298);
or U6801 (N_6801,N_5026,N_4972);
or U6802 (N_6802,N_5544,N_4702);
nand U6803 (N_6803,N_4564,N_5027);
nand U6804 (N_6804,N_5256,N_5561);
xor U6805 (N_6805,N_4672,N_4867);
or U6806 (N_6806,N_4804,N_5841);
nor U6807 (N_6807,N_4543,N_5810);
or U6808 (N_6808,N_5296,N_4878);
or U6809 (N_6809,N_4893,N_4821);
or U6810 (N_6810,N_4999,N_4812);
nor U6811 (N_6811,N_4679,N_5203);
or U6812 (N_6812,N_4769,N_5420);
and U6813 (N_6813,N_4767,N_5291);
or U6814 (N_6814,N_5191,N_4933);
or U6815 (N_6815,N_4618,N_4543);
nor U6816 (N_6816,N_4754,N_5338);
xnor U6817 (N_6817,N_4785,N_4909);
nand U6818 (N_6818,N_5319,N_5293);
or U6819 (N_6819,N_4723,N_4873);
nand U6820 (N_6820,N_5348,N_5033);
or U6821 (N_6821,N_5787,N_5075);
nor U6822 (N_6822,N_5869,N_5826);
or U6823 (N_6823,N_4541,N_4690);
nor U6824 (N_6824,N_4505,N_5165);
or U6825 (N_6825,N_4744,N_5434);
nand U6826 (N_6826,N_5059,N_5004);
nand U6827 (N_6827,N_5526,N_5784);
or U6828 (N_6828,N_4921,N_5081);
or U6829 (N_6829,N_5413,N_5758);
and U6830 (N_6830,N_5123,N_5516);
nand U6831 (N_6831,N_4843,N_5173);
nand U6832 (N_6832,N_5083,N_5607);
nor U6833 (N_6833,N_5248,N_4945);
nand U6834 (N_6834,N_5330,N_4965);
nor U6835 (N_6835,N_5070,N_5087);
or U6836 (N_6836,N_5589,N_5916);
nand U6837 (N_6837,N_5401,N_4931);
or U6838 (N_6838,N_5133,N_5879);
nand U6839 (N_6839,N_4932,N_5443);
xnor U6840 (N_6840,N_5467,N_4844);
and U6841 (N_6841,N_4698,N_4701);
nor U6842 (N_6842,N_4570,N_5171);
nand U6843 (N_6843,N_5501,N_5598);
nor U6844 (N_6844,N_4863,N_5059);
or U6845 (N_6845,N_5710,N_4974);
nand U6846 (N_6846,N_5940,N_5728);
and U6847 (N_6847,N_5570,N_5350);
xnor U6848 (N_6848,N_4601,N_4778);
and U6849 (N_6849,N_5138,N_4902);
and U6850 (N_6850,N_4674,N_5312);
or U6851 (N_6851,N_4751,N_5011);
or U6852 (N_6852,N_4684,N_5027);
or U6853 (N_6853,N_5404,N_5776);
and U6854 (N_6854,N_4888,N_5690);
nor U6855 (N_6855,N_5399,N_4612);
and U6856 (N_6856,N_5064,N_4887);
xnor U6857 (N_6857,N_5709,N_5343);
and U6858 (N_6858,N_4602,N_5175);
nor U6859 (N_6859,N_5127,N_5110);
nor U6860 (N_6860,N_5060,N_5908);
and U6861 (N_6861,N_5824,N_4527);
nand U6862 (N_6862,N_4673,N_5289);
nand U6863 (N_6863,N_5628,N_4824);
xnor U6864 (N_6864,N_5972,N_5022);
nand U6865 (N_6865,N_4695,N_5775);
and U6866 (N_6866,N_4792,N_4944);
and U6867 (N_6867,N_5779,N_5954);
nand U6868 (N_6868,N_4949,N_5372);
and U6869 (N_6869,N_5044,N_4765);
and U6870 (N_6870,N_4873,N_5786);
nand U6871 (N_6871,N_4799,N_5830);
or U6872 (N_6872,N_5410,N_5863);
and U6873 (N_6873,N_5828,N_4596);
nand U6874 (N_6874,N_5501,N_5178);
nand U6875 (N_6875,N_5859,N_4719);
nand U6876 (N_6876,N_5356,N_5014);
or U6877 (N_6877,N_5631,N_5195);
and U6878 (N_6878,N_4960,N_5835);
nand U6879 (N_6879,N_4890,N_4902);
nor U6880 (N_6880,N_4672,N_5832);
nor U6881 (N_6881,N_5858,N_5663);
and U6882 (N_6882,N_5248,N_5456);
or U6883 (N_6883,N_5899,N_5381);
nor U6884 (N_6884,N_5935,N_5835);
nand U6885 (N_6885,N_4955,N_4511);
nor U6886 (N_6886,N_5049,N_4527);
or U6887 (N_6887,N_5659,N_5702);
or U6888 (N_6888,N_5660,N_5051);
xor U6889 (N_6889,N_5778,N_5963);
nor U6890 (N_6890,N_5980,N_4968);
nand U6891 (N_6891,N_4546,N_5544);
nand U6892 (N_6892,N_4769,N_5732);
nor U6893 (N_6893,N_5188,N_4570);
or U6894 (N_6894,N_4579,N_5257);
nand U6895 (N_6895,N_5992,N_4918);
or U6896 (N_6896,N_5964,N_5518);
nand U6897 (N_6897,N_5045,N_5985);
or U6898 (N_6898,N_5056,N_4997);
and U6899 (N_6899,N_5386,N_5392);
nor U6900 (N_6900,N_4899,N_4832);
nor U6901 (N_6901,N_5598,N_5861);
or U6902 (N_6902,N_4872,N_5877);
nor U6903 (N_6903,N_5825,N_5713);
and U6904 (N_6904,N_5277,N_4768);
and U6905 (N_6905,N_4697,N_5926);
nor U6906 (N_6906,N_5695,N_5383);
nor U6907 (N_6907,N_5838,N_5311);
or U6908 (N_6908,N_4930,N_4561);
nor U6909 (N_6909,N_4652,N_5531);
and U6910 (N_6910,N_4950,N_5202);
xnor U6911 (N_6911,N_5541,N_5125);
nand U6912 (N_6912,N_5930,N_5434);
and U6913 (N_6913,N_4859,N_5011);
or U6914 (N_6914,N_5645,N_5863);
and U6915 (N_6915,N_5674,N_5677);
and U6916 (N_6916,N_5846,N_4510);
nand U6917 (N_6917,N_4734,N_4631);
nand U6918 (N_6918,N_4788,N_4997);
or U6919 (N_6919,N_5682,N_4548);
nor U6920 (N_6920,N_5471,N_5589);
nand U6921 (N_6921,N_4824,N_5317);
and U6922 (N_6922,N_5138,N_4616);
or U6923 (N_6923,N_4698,N_5466);
and U6924 (N_6924,N_5490,N_5658);
nand U6925 (N_6925,N_4586,N_4734);
and U6926 (N_6926,N_4943,N_5128);
nand U6927 (N_6927,N_5647,N_4544);
nand U6928 (N_6928,N_4939,N_5227);
and U6929 (N_6929,N_5538,N_5470);
nand U6930 (N_6930,N_4960,N_5940);
or U6931 (N_6931,N_4725,N_5455);
xnor U6932 (N_6932,N_5100,N_5901);
nand U6933 (N_6933,N_5587,N_5233);
nand U6934 (N_6934,N_5738,N_5500);
xor U6935 (N_6935,N_5311,N_5360);
and U6936 (N_6936,N_5100,N_5919);
and U6937 (N_6937,N_4712,N_4500);
nor U6938 (N_6938,N_5446,N_4952);
nand U6939 (N_6939,N_5786,N_4504);
and U6940 (N_6940,N_4687,N_4752);
and U6941 (N_6941,N_5526,N_4828);
xor U6942 (N_6942,N_5503,N_5878);
nor U6943 (N_6943,N_5483,N_4620);
nand U6944 (N_6944,N_4842,N_5263);
or U6945 (N_6945,N_5086,N_4897);
or U6946 (N_6946,N_5801,N_4824);
nand U6947 (N_6947,N_5756,N_4946);
or U6948 (N_6948,N_4805,N_4963);
nor U6949 (N_6949,N_4636,N_4890);
nand U6950 (N_6950,N_5447,N_5742);
and U6951 (N_6951,N_4832,N_5442);
nand U6952 (N_6952,N_5956,N_5811);
nand U6953 (N_6953,N_4553,N_5361);
or U6954 (N_6954,N_5567,N_5428);
or U6955 (N_6955,N_5512,N_5200);
and U6956 (N_6956,N_5711,N_5603);
xor U6957 (N_6957,N_5043,N_4617);
or U6958 (N_6958,N_5769,N_5217);
xnor U6959 (N_6959,N_4963,N_5519);
or U6960 (N_6960,N_4976,N_4558);
and U6961 (N_6961,N_5942,N_5952);
xnor U6962 (N_6962,N_5439,N_4907);
nor U6963 (N_6963,N_5922,N_5726);
nor U6964 (N_6964,N_5932,N_5969);
and U6965 (N_6965,N_5514,N_5271);
nor U6966 (N_6966,N_5595,N_5867);
and U6967 (N_6967,N_5690,N_5510);
and U6968 (N_6968,N_5023,N_5409);
or U6969 (N_6969,N_5776,N_4887);
nand U6970 (N_6970,N_4508,N_5982);
nor U6971 (N_6971,N_5477,N_5843);
and U6972 (N_6972,N_4675,N_5106);
nor U6973 (N_6973,N_5092,N_5388);
or U6974 (N_6974,N_4870,N_5998);
and U6975 (N_6975,N_4838,N_5296);
and U6976 (N_6976,N_5660,N_4638);
and U6977 (N_6977,N_5932,N_4750);
or U6978 (N_6978,N_4801,N_5009);
nand U6979 (N_6979,N_4583,N_5968);
nand U6980 (N_6980,N_4503,N_4945);
or U6981 (N_6981,N_4820,N_5941);
and U6982 (N_6982,N_5293,N_4999);
xnor U6983 (N_6983,N_5214,N_5927);
nor U6984 (N_6984,N_5333,N_5619);
nor U6985 (N_6985,N_5803,N_4718);
nand U6986 (N_6986,N_4626,N_5807);
nand U6987 (N_6987,N_5778,N_5374);
nor U6988 (N_6988,N_5502,N_5190);
xor U6989 (N_6989,N_4534,N_5232);
nand U6990 (N_6990,N_5203,N_5071);
nand U6991 (N_6991,N_5214,N_5240);
and U6992 (N_6992,N_4944,N_5820);
nor U6993 (N_6993,N_5624,N_5252);
nor U6994 (N_6994,N_5016,N_5309);
or U6995 (N_6995,N_5223,N_5477);
and U6996 (N_6996,N_5927,N_5292);
nor U6997 (N_6997,N_5989,N_4625);
nor U6998 (N_6998,N_5063,N_4968);
and U6999 (N_6999,N_4689,N_5314);
and U7000 (N_7000,N_5376,N_4501);
nand U7001 (N_7001,N_4728,N_5974);
xor U7002 (N_7002,N_4946,N_5338);
nand U7003 (N_7003,N_5660,N_4660);
nand U7004 (N_7004,N_4972,N_5173);
or U7005 (N_7005,N_4726,N_5628);
and U7006 (N_7006,N_5897,N_5932);
and U7007 (N_7007,N_5402,N_4860);
xor U7008 (N_7008,N_5656,N_4945);
and U7009 (N_7009,N_4785,N_5756);
xor U7010 (N_7010,N_5010,N_5354);
or U7011 (N_7011,N_5436,N_5779);
nor U7012 (N_7012,N_5809,N_5401);
nor U7013 (N_7013,N_5833,N_5945);
nand U7014 (N_7014,N_4527,N_4708);
or U7015 (N_7015,N_5048,N_5633);
and U7016 (N_7016,N_4917,N_5706);
and U7017 (N_7017,N_5994,N_5054);
or U7018 (N_7018,N_4577,N_4976);
xnor U7019 (N_7019,N_4807,N_5055);
nand U7020 (N_7020,N_5558,N_5722);
or U7021 (N_7021,N_5709,N_5350);
and U7022 (N_7022,N_4534,N_5231);
nor U7023 (N_7023,N_5697,N_5558);
xnor U7024 (N_7024,N_4715,N_5234);
and U7025 (N_7025,N_4634,N_5862);
xnor U7026 (N_7026,N_5302,N_5096);
and U7027 (N_7027,N_4696,N_5094);
and U7028 (N_7028,N_5378,N_4886);
nand U7029 (N_7029,N_5781,N_5550);
nand U7030 (N_7030,N_5524,N_5139);
or U7031 (N_7031,N_5160,N_5544);
nor U7032 (N_7032,N_5932,N_5735);
and U7033 (N_7033,N_5603,N_5435);
nor U7034 (N_7034,N_4542,N_5269);
nand U7035 (N_7035,N_5660,N_4547);
xor U7036 (N_7036,N_4799,N_5588);
and U7037 (N_7037,N_5738,N_5437);
or U7038 (N_7038,N_4613,N_5179);
and U7039 (N_7039,N_4570,N_5975);
and U7040 (N_7040,N_4557,N_5809);
nand U7041 (N_7041,N_4688,N_4561);
nand U7042 (N_7042,N_4696,N_5981);
nor U7043 (N_7043,N_5794,N_5529);
and U7044 (N_7044,N_4721,N_5220);
nand U7045 (N_7045,N_5196,N_5267);
nand U7046 (N_7046,N_4526,N_5792);
nand U7047 (N_7047,N_5099,N_4852);
nor U7048 (N_7048,N_5427,N_5290);
nand U7049 (N_7049,N_4749,N_5164);
or U7050 (N_7050,N_4941,N_4783);
or U7051 (N_7051,N_5404,N_5376);
and U7052 (N_7052,N_5927,N_4984);
nand U7053 (N_7053,N_5009,N_5551);
nor U7054 (N_7054,N_4950,N_5308);
nor U7055 (N_7055,N_5657,N_5707);
and U7056 (N_7056,N_5105,N_5253);
and U7057 (N_7057,N_4647,N_5109);
nand U7058 (N_7058,N_5616,N_4648);
nor U7059 (N_7059,N_4953,N_4645);
or U7060 (N_7060,N_4511,N_4554);
or U7061 (N_7061,N_5274,N_4542);
and U7062 (N_7062,N_5537,N_4512);
nand U7063 (N_7063,N_5678,N_5754);
nand U7064 (N_7064,N_5031,N_5672);
nand U7065 (N_7065,N_5870,N_4572);
nand U7066 (N_7066,N_4667,N_5249);
or U7067 (N_7067,N_4663,N_4979);
xor U7068 (N_7068,N_5737,N_5082);
nor U7069 (N_7069,N_4684,N_5945);
and U7070 (N_7070,N_4859,N_5352);
and U7071 (N_7071,N_4506,N_5831);
nor U7072 (N_7072,N_5728,N_5758);
and U7073 (N_7073,N_5027,N_5659);
nand U7074 (N_7074,N_4596,N_4806);
nand U7075 (N_7075,N_4877,N_4506);
nor U7076 (N_7076,N_5129,N_5851);
xnor U7077 (N_7077,N_5809,N_5357);
xnor U7078 (N_7078,N_4714,N_5346);
nor U7079 (N_7079,N_5775,N_5801);
nor U7080 (N_7080,N_5032,N_5912);
nor U7081 (N_7081,N_5424,N_4559);
nand U7082 (N_7082,N_5355,N_4747);
xor U7083 (N_7083,N_4547,N_4840);
and U7084 (N_7084,N_4669,N_4893);
nand U7085 (N_7085,N_5855,N_4999);
or U7086 (N_7086,N_4937,N_5132);
and U7087 (N_7087,N_5556,N_4947);
xor U7088 (N_7088,N_5127,N_5029);
or U7089 (N_7089,N_4763,N_5280);
or U7090 (N_7090,N_4938,N_5793);
or U7091 (N_7091,N_5840,N_5810);
or U7092 (N_7092,N_5384,N_5523);
or U7093 (N_7093,N_5288,N_4886);
and U7094 (N_7094,N_4812,N_4862);
and U7095 (N_7095,N_5513,N_4703);
and U7096 (N_7096,N_5242,N_5010);
nor U7097 (N_7097,N_4807,N_4857);
nor U7098 (N_7098,N_5943,N_5483);
nand U7099 (N_7099,N_5747,N_4650);
or U7100 (N_7100,N_5806,N_5124);
or U7101 (N_7101,N_5056,N_5335);
nor U7102 (N_7102,N_5797,N_5769);
nor U7103 (N_7103,N_5962,N_4855);
nor U7104 (N_7104,N_5059,N_5117);
nor U7105 (N_7105,N_5212,N_5943);
xnor U7106 (N_7106,N_5637,N_5471);
or U7107 (N_7107,N_4986,N_5609);
nor U7108 (N_7108,N_5367,N_5831);
nand U7109 (N_7109,N_5100,N_5640);
nand U7110 (N_7110,N_5237,N_5084);
nand U7111 (N_7111,N_5653,N_5558);
and U7112 (N_7112,N_5917,N_5487);
or U7113 (N_7113,N_5777,N_5478);
xor U7114 (N_7114,N_5385,N_4644);
nand U7115 (N_7115,N_5135,N_4976);
xnor U7116 (N_7116,N_5963,N_5511);
and U7117 (N_7117,N_4742,N_5789);
and U7118 (N_7118,N_5468,N_5031);
xor U7119 (N_7119,N_5622,N_4550);
nor U7120 (N_7120,N_5500,N_5067);
and U7121 (N_7121,N_5446,N_4773);
or U7122 (N_7122,N_5447,N_5754);
nor U7123 (N_7123,N_5321,N_5457);
xor U7124 (N_7124,N_5045,N_4982);
nor U7125 (N_7125,N_5931,N_5393);
or U7126 (N_7126,N_4957,N_5631);
xor U7127 (N_7127,N_5278,N_5383);
and U7128 (N_7128,N_5631,N_4979);
and U7129 (N_7129,N_4550,N_4992);
and U7130 (N_7130,N_5994,N_5563);
nor U7131 (N_7131,N_5792,N_4650);
and U7132 (N_7132,N_5148,N_4799);
xnor U7133 (N_7133,N_5920,N_5648);
nand U7134 (N_7134,N_4912,N_4810);
xnor U7135 (N_7135,N_5033,N_5819);
nand U7136 (N_7136,N_5557,N_4837);
nor U7137 (N_7137,N_5130,N_5257);
nand U7138 (N_7138,N_5351,N_5343);
nand U7139 (N_7139,N_5320,N_5068);
nand U7140 (N_7140,N_5970,N_5480);
or U7141 (N_7141,N_5094,N_5306);
nand U7142 (N_7142,N_5817,N_5380);
and U7143 (N_7143,N_4677,N_4545);
nand U7144 (N_7144,N_4789,N_5294);
nand U7145 (N_7145,N_5833,N_5210);
nand U7146 (N_7146,N_5742,N_5556);
and U7147 (N_7147,N_4559,N_5686);
and U7148 (N_7148,N_5073,N_5453);
nand U7149 (N_7149,N_4550,N_4966);
nand U7150 (N_7150,N_4599,N_5879);
nand U7151 (N_7151,N_4579,N_5066);
nor U7152 (N_7152,N_5824,N_4877);
nand U7153 (N_7153,N_4730,N_4926);
nor U7154 (N_7154,N_5603,N_5832);
and U7155 (N_7155,N_4512,N_5754);
or U7156 (N_7156,N_5411,N_4809);
and U7157 (N_7157,N_4699,N_4805);
nand U7158 (N_7158,N_4668,N_5826);
or U7159 (N_7159,N_5857,N_4930);
or U7160 (N_7160,N_5039,N_5527);
nand U7161 (N_7161,N_5639,N_5585);
and U7162 (N_7162,N_5887,N_5778);
nand U7163 (N_7163,N_5988,N_5602);
and U7164 (N_7164,N_5377,N_5124);
nand U7165 (N_7165,N_5303,N_5998);
xor U7166 (N_7166,N_5177,N_5134);
and U7167 (N_7167,N_4947,N_5420);
nand U7168 (N_7168,N_5603,N_5590);
and U7169 (N_7169,N_5484,N_5476);
nand U7170 (N_7170,N_5253,N_4835);
nand U7171 (N_7171,N_5766,N_5630);
nor U7172 (N_7172,N_4722,N_5695);
nor U7173 (N_7173,N_4544,N_5318);
or U7174 (N_7174,N_5742,N_5859);
and U7175 (N_7175,N_5612,N_5844);
or U7176 (N_7176,N_4597,N_4828);
or U7177 (N_7177,N_4519,N_5451);
and U7178 (N_7178,N_5668,N_5545);
xnor U7179 (N_7179,N_4524,N_5510);
nor U7180 (N_7180,N_5925,N_5260);
and U7181 (N_7181,N_5285,N_5106);
and U7182 (N_7182,N_4736,N_4942);
nor U7183 (N_7183,N_4504,N_5967);
or U7184 (N_7184,N_5540,N_5016);
nor U7185 (N_7185,N_5800,N_5510);
xor U7186 (N_7186,N_5321,N_4987);
or U7187 (N_7187,N_4666,N_5376);
and U7188 (N_7188,N_5500,N_5710);
nor U7189 (N_7189,N_5844,N_5629);
nor U7190 (N_7190,N_4948,N_5692);
nor U7191 (N_7191,N_5278,N_5900);
nor U7192 (N_7192,N_5641,N_5954);
nor U7193 (N_7193,N_5878,N_5295);
and U7194 (N_7194,N_4872,N_5393);
or U7195 (N_7195,N_5106,N_5325);
xnor U7196 (N_7196,N_5322,N_4787);
and U7197 (N_7197,N_5396,N_4518);
or U7198 (N_7198,N_5523,N_4515);
nor U7199 (N_7199,N_4844,N_5413);
nor U7200 (N_7200,N_5913,N_5530);
and U7201 (N_7201,N_5760,N_5100);
and U7202 (N_7202,N_5696,N_5262);
xor U7203 (N_7203,N_5516,N_4710);
nor U7204 (N_7204,N_5651,N_4641);
xor U7205 (N_7205,N_4743,N_5298);
nand U7206 (N_7206,N_5187,N_5119);
xor U7207 (N_7207,N_4700,N_5085);
xor U7208 (N_7208,N_4523,N_5092);
xnor U7209 (N_7209,N_5421,N_4872);
or U7210 (N_7210,N_4964,N_5004);
nand U7211 (N_7211,N_5398,N_5019);
and U7212 (N_7212,N_5993,N_5852);
nor U7213 (N_7213,N_5301,N_5303);
or U7214 (N_7214,N_5200,N_4605);
xor U7215 (N_7215,N_5402,N_5486);
nor U7216 (N_7216,N_4724,N_5668);
nor U7217 (N_7217,N_4786,N_5051);
nor U7218 (N_7218,N_4859,N_5409);
and U7219 (N_7219,N_5500,N_5434);
or U7220 (N_7220,N_5316,N_4567);
or U7221 (N_7221,N_5820,N_5247);
nor U7222 (N_7222,N_4610,N_5756);
and U7223 (N_7223,N_5664,N_5155);
nor U7224 (N_7224,N_5505,N_5407);
xor U7225 (N_7225,N_5781,N_5725);
and U7226 (N_7226,N_4683,N_4884);
nor U7227 (N_7227,N_5854,N_4844);
or U7228 (N_7228,N_5584,N_5490);
or U7229 (N_7229,N_5816,N_4819);
nor U7230 (N_7230,N_5991,N_5437);
nor U7231 (N_7231,N_5705,N_5452);
nor U7232 (N_7232,N_5315,N_4855);
and U7233 (N_7233,N_5071,N_5230);
or U7234 (N_7234,N_5124,N_5710);
nor U7235 (N_7235,N_5157,N_4568);
xor U7236 (N_7236,N_4535,N_5630);
nor U7237 (N_7237,N_5843,N_4622);
or U7238 (N_7238,N_4715,N_4767);
or U7239 (N_7239,N_4550,N_5496);
nor U7240 (N_7240,N_5017,N_4591);
nand U7241 (N_7241,N_5558,N_5224);
nand U7242 (N_7242,N_5449,N_5411);
nand U7243 (N_7243,N_5639,N_4523);
nor U7244 (N_7244,N_5102,N_4798);
nand U7245 (N_7245,N_4757,N_5021);
nor U7246 (N_7246,N_5694,N_4793);
nor U7247 (N_7247,N_4530,N_5067);
nand U7248 (N_7248,N_5757,N_4762);
nand U7249 (N_7249,N_4571,N_4678);
nand U7250 (N_7250,N_5008,N_5787);
nand U7251 (N_7251,N_4621,N_5112);
nand U7252 (N_7252,N_5761,N_5620);
xnor U7253 (N_7253,N_4685,N_5460);
nor U7254 (N_7254,N_4533,N_4843);
nand U7255 (N_7255,N_5151,N_4789);
nor U7256 (N_7256,N_4519,N_5516);
or U7257 (N_7257,N_5396,N_4772);
nor U7258 (N_7258,N_4915,N_5284);
nor U7259 (N_7259,N_5896,N_5401);
and U7260 (N_7260,N_5488,N_5985);
nor U7261 (N_7261,N_5985,N_5109);
nor U7262 (N_7262,N_4605,N_4816);
nand U7263 (N_7263,N_5984,N_5640);
nor U7264 (N_7264,N_5250,N_5287);
or U7265 (N_7265,N_5848,N_5940);
and U7266 (N_7266,N_5738,N_5772);
nor U7267 (N_7267,N_5947,N_5131);
and U7268 (N_7268,N_5538,N_5952);
nand U7269 (N_7269,N_4902,N_5359);
nand U7270 (N_7270,N_5563,N_5280);
nor U7271 (N_7271,N_4595,N_5779);
xor U7272 (N_7272,N_5585,N_5825);
or U7273 (N_7273,N_5055,N_4777);
nand U7274 (N_7274,N_5281,N_5912);
or U7275 (N_7275,N_4720,N_4601);
nand U7276 (N_7276,N_5237,N_5225);
nor U7277 (N_7277,N_4766,N_5868);
nor U7278 (N_7278,N_5138,N_5579);
or U7279 (N_7279,N_4820,N_4719);
nand U7280 (N_7280,N_5421,N_5521);
or U7281 (N_7281,N_4911,N_5196);
nand U7282 (N_7282,N_4718,N_4978);
xor U7283 (N_7283,N_4892,N_5323);
nand U7284 (N_7284,N_5611,N_5042);
and U7285 (N_7285,N_5897,N_4811);
nor U7286 (N_7286,N_4661,N_4757);
nor U7287 (N_7287,N_5464,N_4616);
xor U7288 (N_7288,N_4688,N_5680);
or U7289 (N_7289,N_4935,N_4574);
nor U7290 (N_7290,N_5850,N_4765);
nor U7291 (N_7291,N_5596,N_4628);
nand U7292 (N_7292,N_4588,N_5340);
nand U7293 (N_7293,N_4958,N_5412);
or U7294 (N_7294,N_4784,N_5656);
nand U7295 (N_7295,N_5351,N_5390);
nand U7296 (N_7296,N_5939,N_5822);
xor U7297 (N_7297,N_5152,N_5214);
and U7298 (N_7298,N_5496,N_4542);
nand U7299 (N_7299,N_5993,N_5372);
nor U7300 (N_7300,N_4590,N_5101);
nor U7301 (N_7301,N_5504,N_5896);
xor U7302 (N_7302,N_4505,N_5436);
and U7303 (N_7303,N_5160,N_4872);
nand U7304 (N_7304,N_5856,N_4607);
nand U7305 (N_7305,N_5423,N_5212);
xnor U7306 (N_7306,N_5167,N_4993);
or U7307 (N_7307,N_5495,N_4524);
and U7308 (N_7308,N_5189,N_5522);
nor U7309 (N_7309,N_5081,N_4888);
or U7310 (N_7310,N_5527,N_5267);
nand U7311 (N_7311,N_4986,N_4774);
nor U7312 (N_7312,N_5567,N_5484);
and U7313 (N_7313,N_4942,N_5319);
nand U7314 (N_7314,N_4691,N_4952);
and U7315 (N_7315,N_5468,N_4534);
nor U7316 (N_7316,N_5076,N_5442);
nand U7317 (N_7317,N_5541,N_4710);
or U7318 (N_7318,N_5333,N_5792);
nor U7319 (N_7319,N_5442,N_4766);
nor U7320 (N_7320,N_4540,N_5794);
and U7321 (N_7321,N_4649,N_4566);
and U7322 (N_7322,N_5253,N_4819);
xnor U7323 (N_7323,N_5524,N_4601);
nor U7324 (N_7324,N_4585,N_4805);
xor U7325 (N_7325,N_5575,N_5822);
or U7326 (N_7326,N_5593,N_4533);
nor U7327 (N_7327,N_4894,N_5724);
nor U7328 (N_7328,N_5637,N_5157);
and U7329 (N_7329,N_4556,N_4504);
nand U7330 (N_7330,N_4857,N_5077);
and U7331 (N_7331,N_4756,N_5042);
nand U7332 (N_7332,N_5809,N_5943);
and U7333 (N_7333,N_4651,N_4842);
nand U7334 (N_7334,N_4992,N_4702);
nor U7335 (N_7335,N_5039,N_5873);
nand U7336 (N_7336,N_5862,N_4663);
nor U7337 (N_7337,N_5443,N_5789);
or U7338 (N_7338,N_4935,N_5273);
nor U7339 (N_7339,N_5655,N_5380);
nor U7340 (N_7340,N_4902,N_4770);
or U7341 (N_7341,N_5807,N_4709);
and U7342 (N_7342,N_5447,N_5668);
or U7343 (N_7343,N_4934,N_5864);
and U7344 (N_7344,N_4720,N_5250);
or U7345 (N_7345,N_5763,N_5827);
nor U7346 (N_7346,N_5893,N_4718);
or U7347 (N_7347,N_5653,N_4560);
nor U7348 (N_7348,N_5706,N_5207);
or U7349 (N_7349,N_5632,N_5427);
nand U7350 (N_7350,N_4590,N_5226);
and U7351 (N_7351,N_4813,N_4902);
nand U7352 (N_7352,N_5741,N_5436);
and U7353 (N_7353,N_5254,N_5461);
nand U7354 (N_7354,N_5612,N_4715);
nand U7355 (N_7355,N_5340,N_5439);
nand U7356 (N_7356,N_5588,N_5060);
nor U7357 (N_7357,N_5690,N_5986);
or U7358 (N_7358,N_5748,N_5077);
or U7359 (N_7359,N_4642,N_5665);
or U7360 (N_7360,N_5192,N_5109);
xnor U7361 (N_7361,N_5009,N_4785);
and U7362 (N_7362,N_5942,N_5775);
nor U7363 (N_7363,N_5773,N_5445);
and U7364 (N_7364,N_4717,N_5616);
and U7365 (N_7365,N_5020,N_5665);
and U7366 (N_7366,N_4517,N_5865);
nor U7367 (N_7367,N_5963,N_5019);
nor U7368 (N_7368,N_5168,N_5518);
or U7369 (N_7369,N_4521,N_4589);
or U7370 (N_7370,N_5707,N_4971);
xor U7371 (N_7371,N_5002,N_4539);
or U7372 (N_7372,N_5238,N_4509);
or U7373 (N_7373,N_5349,N_5472);
xor U7374 (N_7374,N_4875,N_4953);
and U7375 (N_7375,N_5367,N_4698);
nor U7376 (N_7376,N_5587,N_5312);
nor U7377 (N_7377,N_4631,N_5260);
and U7378 (N_7378,N_5414,N_5704);
or U7379 (N_7379,N_4894,N_5356);
xnor U7380 (N_7380,N_4909,N_5975);
and U7381 (N_7381,N_5507,N_4541);
nand U7382 (N_7382,N_4962,N_5721);
nor U7383 (N_7383,N_5385,N_5116);
xnor U7384 (N_7384,N_5312,N_4893);
nand U7385 (N_7385,N_5192,N_5854);
or U7386 (N_7386,N_5457,N_5887);
nor U7387 (N_7387,N_4951,N_4502);
and U7388 (N_7388,N_4982,N_5100);
xor U7389 (N_7389,N_5313,N_4585);
nor U7390 (N_7390,N_4795,N_4556);
nor U7391 (N_7391,N_5032,N_4803);
or U7392 (N_7392,N_4857,N_5288);
or U7393 (N_7393,N_5127,N_4752);
nand U7394 (N_7394,N_5363,N_4596);
nor U7395 (N_7395,N_5536,N_5962);
nor U7396 (N_7396,N_5646,N_5986);
nor U7397 (N_7397,N_5267,N_5009);
nor U7398 (N_7398,N_5027,N_5492);
xnor U7399 (N_7399,N_5910,N_5579);
nor U7400 (N_7400,N_5838,N_4626);
nor U7401 (N_7401,N_5009,N_4748);
nand U7402 (N_7402,N_5066,N_5413);
nor U7403 (N_7403,N_5925,N_5814);
and U7404 (N_7404,N_4634,N_5611);
or U7405 (N_7405,N_5051,N_4886);
nand U7406 (N_7406,N_4954,N_4922);
nand U7407 (N_7407,N_4739,N_4821);
or U7408 (N_7408,N_5095,N_5558);
nor U7409 (N_7409,N_4866,N_5915);
or U7410 (N_7410,N_5657,N_5218);
nand U7411 (N_7411,N_4615,N_5591);
or U7412 (N_7412,N_4618,N_4829);
nand U7413 (N_7413,N_5658,N_5566);
or U7414 (N_7414,N_4522,N_5718);
and U7415 (N_7415,N_5482,N_4968);
xor U7416 (N_7416,N_5907,N_5898);
nand U7417 (N_7417,N_5921,N_4986);
nor U7418 (N_7418,N_5101,N_5269);
nor U7419 (N_7419,N_5522,N_5188);
nand U7420 (N_7420,N_5162,N_5073);
nor U7421 (N_7421,N_5990,N_4999);
nor U7422 (N_7422,N_5713,N_5441);
nor U7423 (N_7423,N_5291,N_4530);
and U7424 (N_7424,N_4998,N_5978);
or U7425 (N_7425,N_4594,N_4660);
nand U7426 (N_7426,N_5544,N_5363);
and U7427 (N_7427,N_5632,N_4589);
xor U7428 (N_7428,N_5511,N_5675);
or U7429 (N_7429,N_4820,N_5294);
nor U7430 (N_7430,N_4714,N_5711);
nand U7431 (N_7431,N_5685,N_5560);
nand U7432 (N_7432,N_4990,N_5435);
and U7433 (N_7433,N_4744,N_4758);
nor U7434 (N_7434,N_5369,N_4667);
or U7435 (N_7435,N_5248,N_5923);
nand U7436 (N_7436,N_5530,N_5078);
nor U7437 (N_7437,N_5177,N_4519);
and U7438 (N_7438,N_5210,N_4590);
nor U7439 (N_7439,N_5054,N_5173);
xnor U7440 (N_7440,N_4576,N_5778);
nand U7441 (N_7441,N_4816,N_4507);
nand U7442 (N_7442,N_5774,N_4621);
or U7443 (N_7443,N_4884,N_5257);
nand U7444 (N_7444,N_5371,N_5711);
nand U7445 (N_7445,N_5396,N_5118);
nor U7446 (N_7446,N_5368,N_5731);
nor U7447 (N_7447,N_5606,N_5563);
xnor U7448 (N_7448,N_5149,N_4990);
or U7449 (N_7449,N_5603,N_4779);
nor U7450 (N_7450,N_5336,N_4851);
xor U7451 (N_7451,N_4548,N_4818);
and U7452 (N_7452,N_4753,N_4773);
nand U7453 (N_7453,N_4532,N_4513);
or U7454 (N_7454,N_5068,N_5218);
nor U7455 (N_7455,N_5841,N_4568);
or U7456 (N_7456,N_5380,N_4660);
nor U7457 (N_7457,N_5096,N_5161);
nand U7458 (N_7458,N_5315,N_5512);
or U7459 (N_7459,N_4859,N_5681);
or U7460 (N_7460,N_5591,N_5660);
nand U7461 (N_7461,N_5872,N_5395);
or U7462 (N_7462,N_5343,N_5645);
nor U7463 (N_7463,N_4921,N_4938);
or U7464 (N_7464,N_4524,N_5407);
or U7465 (N_7465,N_5086,N_4543);
and U7466 (N_7466,N_5435,N_5397);
nand U7467 (N_7467,N_5776,N_5480);
xor U7468 (N_7468,N_5119,N_5246);
or U7469 (N_7469,N_4864,N_5335);
or U7470 (N_7470,N_5886,N_5975);
and U7471 (N_7471,N_4743,N_5518);
or U7472 (N_7472,N_5039,N_5876);
and U7473 (N_7473,N_5959,N_5158);
or U7474 (N_7474,N_5117,N_5184);
and U7475 (N_7475,N_5993,N_5516);
nor U7476 (N_7476,N_5150,N_4579);
nand U7477 (N_7477,N_5254,N_4575);
xor U7478 (N_7478,N_5375,N_4969);
and U7479 (N_7479,N_5445,N_4846);
nand U7480 (N_7480,N_5924,N_4655);
nor U7481 (N_7481,N_5455,N_5255);
nor U7482 (N_7482,N_4704,N_5870);
or U7483 (N_7483,N_5048,N_5265);
nand U7484 (N_7484,N_5830,N_5284);
nor U7485 (N_7485,N_4906,N_4592);
or U7486 (N_7486,N_5896,N_4905);
nand U7487 (N_7487,N_5207,N_5140);
nor U7488 (N_7488,N_5732,N_4840);
or U7489 (N_7489,N_5177,N_5218);
nand U7490 (N_7490,N_5953,N_5335);
or U7491 (N_7491,N_5949,N_4523);
nor U7492 (N_7492,N_5352,N_5914);
or U7493 (N_7493,N_5492,N_4905);
nor U7494 (N_7494,N_5545,N_5160);
nand U7495 (N_7495,N_4910,N_5860);
xor U7496 (N_7496,N_4893,N_5809);
and U7497 (N_7497,N_5209,N_5165);
nand U7498 (N_7498,N_4896,N_5298);
or U7499 (N_7499,N_5172,N_4829);
nand U7500 (N_7500,N_7076,N_6563);
and U7501 (N_7501,N_6789,N_7128);
nor U7502 (N_7502,N_7004,N_6330);
nand U7503 (N_7503,N_7364,N_6309);
nor U7504 (N_7504,N_6977,N_6541);
nor U7505 (N_7505,N_6101,N_6104);
or U7506 (N_7506,N_7101,N_6471);
and U7507 (N_7507,N_6362,N_6239);
and U7508 (N_7508,N_6686,N_6581);
nand U7509 (N_7509,N_7480,N_6653);
nor U7510 (N_7510,N_6633,N_7475);
nor U7511 (N_7511,N_6407,N_6442);
or U7512 (N_7512,N_6978,N_7226);
or U7513 (N_7513,N_6358,N_6922);
and U7514 (N_7514,N_6934,N_6771);
or U7515 (N_7515,N_7313,N_7441);
nand U7516 (N_7516,N_7381,N_7366);
nand U7517 (N_7517,N_6738,N_7301);
or U7518 (N_7518,N_7114,N_6074);
or U7519 (N_7519,N_7136,N_6796);
and U7520 (N_7520,N_6122,N_6770);
xnor U7521 (N_7521,N_6228,N_6158);
or U7522 (N_7522,N_6012,N_6129);
or U7523 (N_7523,N_7311,N_7115);
nand U7524 (N_7524,N_6534,N_7474);
nand U7525 (N_7525,N_6982,N_6544);
xnor U7526 (N_7526,N_7410,N_6002);
xor U7527 (N_7527,N_7359,N_6613);
and U7528 (N_7528,N_7195,N_6916);
or U7529 (N_7529,N_6831,N_6298);
nor U7530 (N_7530,N_6269,N_6612);
and U7531 (N_7531,N_7434,N_6828);
nor U7532 (N_7532,N_7223,N_6510);
or U7533 (N_7533,N_7310,N_6657);
or U7534 (N_7534,N_7220,N_7224);
xor U7535 (N_7535,N_7215,N_6338);
nor U7536 (N_7536,N_6179,N_6683);
nor U7537 (N_7537,N_7140,N_6460);
and U7538 (N_7538,N_7249,N_7367);
and U7539 (N_7539,N_7360,N_6675);
or U7540 (N_7540,N_7113,N_6087);
nand U7541 (N_7541,N_7148,N_7125);
xor U7542 (N_7542,N_6804,N_7336);
nor U7543 (N_7543,N_7210,N_7078);
nor U7544 (N_7544,N_6660,N_6661);
nor U7545 (N_7545,N_6601,N_6229);
nor U7546 (N_7546,N_6145,N_6996);
nor U7547 (N_7547,N_6281,N_7216);
nand U7548 (N_7548,N_6291,N_7044);
nor U7549 (N_7549,N_6760,N_6640);
nand U7550 (N_7550,N_6328,N_6718);
or U7551 (N_7551,N_6435,N_7478);
nor U7552 (N_7552,N_7071,N_7376);
nor U7553 (N_7553,N_6997,N_6154);
nand U7554 (N_7554,N_6602,N_6234);
nor U7555 (N_7555,N_7244,N_6860);
nor U7556 (N_7556,N_6149,N_6008);
or U7557 (N_7557,N_7425,N_6808);
and U7558 (N_7558,N_7124,N_6036);
nor U7559 (N_7559,N_6722,N_6626);
xor U7560 (N_7560,N_6577,N_6324);
or U7561 (N_7561,N_6375,N_6483);
nor U7562 (N_7562,N_6908,N_7116);
nand U7563 (N_7563,N_6028,N_7279);
xor U7564 (N_7564,N_6265,N_7253);
and U7565 (N_7565,N_6513,N_6866);
or U7566 (N_7566,N_6021,N_6851);
nand U7567 (N_7567,N_6800,N_7119);
nor U7568 (N_7568,N_6632,N_6905);
nand U7569 (N_7569,N_6004,N_6401);
nand U7570 (N_7570,N_7447,N_6636);
and U7571 (N_7571,N_6098,N_6197);
and U7572 (N_7572,N_6352,N_6668);
or U7573 (N_7573,N_6462,N_6238);
and U7574 (N_7574,N_6505,N_7179);
and U7575 (N_7575,N_7137,N_7315);
or U7576 (N_7576,N_6748,N_7386);
or U7577 (N_7577,N_7048,N_6132);
nand U7578 (N_7578,N_6628,N_6568);
xor U7579 (N_7579,N_6425,N_6807);
and U7580 (N_7580,N_6936,N_6123);
nor U7581 (N_7581,N_6220,N_6517);
nor U7582 (N_7582,N_6015,N_6662);
nor U7583 (N_7583,N_6932,N_6904);
and U7584 (N_7584,N_7056,N_7399);
or U7585 (N_7585,N_6003,N_7324);
xor U7586 (N_7586,N_6210,N_7344);
and U7587 (N_7587,N_6912,N_6852);
nand U7588 (N_7588,N_6337,N_6560);
or U7589 (N_7589,N_7337,N_6350);
nand U7590 (N_7590,N_6455,N_6516);
nor U7591 (N_7591,N_6797,N_6452);
or U7592 (N_7592,N_7123,N_6398);
xnor U7593 (N_7593,N_6507,N_7174);
nor U7594 (N_7594,N_7126,N_7018);
and U7595 (N_7595,N_6838,N_7012);
nand U7596 (N_7596,N_6832,N_6751);
and U7597 (N_7597,N_6485,N_6684);
and U7598 (N_7598,N_6928,N_6092);
nand U7599 (N_7599,N_6524,N_6607);
nor U7600 (N_7600,N_6884,N_6713);
or U7601 (N_7601,N_7192,N_7194);
or U7602 (N_7602,N_7422,N_6217);
nor U7603 (N_7603,N_6424,N_6902);
nor U7604 (N_7604,N_6499,N_7038);
xnor U7605 (N_7605,N_6528,N_6892);
nand U7606 (N_7606,N_7015,N_6476);
or U7607 (N_7607,N_6813,N_6081);
or U7608 (N_7608,N_6288,N_6365);
nor U7609 (N_7609,N_7321,N_6681);
or U7610 (N_7610,N_7055,N_6227);
xnor U7611 (N_7611,N_6161,N_6196);
xor U7612 (N_7612,N_7118,N_6259);
nand U7613 (N_7613,N_6392,N_6169);
nor U7614 (N_7614,N_6631,N_7104);
nor U7615 (N_7615,N_6065,N_6105);
or U7616 (N_7616,N_6715,N_7189);
nand U7617 (N_7617,N_6182,N_7146);
nand U7618 (N_7618,N_6275,N_6189);
or U7619 (N_7619,N_6068,N_6351);
nor U7620 (N_7620,N_6692,N_6746);
or U7621 (N_7621,N_6047,N_7283);
and U7622 (N_7622,N_6609,N_6589);
nand U7623 (N_7623,N_6836,N_6556);
or U7624 (N_7624,N_7369,N_6233);
nor U7625 (N_7625,N_7257,N_6914);
or U7626 (N_7626,N_6150,N_6787);
nand U7627 (N_7627,N_6484,N_6585);
nor U7628 (N_7628,N_6010,N_7288);
or U7629 (N_7629,N_6744,N_6946);
and U7630 (N_7630,N_6215,N_6745);
and U7631 (N_7631,N_6390,N_6638);
nor U7632 (N_7632,N_7162,N_7089);
and U7633 (N_7633,N_7286,N_6942);
nand U7634 (N_7634,N_6898,N_6409);
nand U7635 (N_7635,N_6418,N_7485);
nor U7636 (N_7636,N_7456,N_7496);
nand U7637 (N_7637,N_6237,N_6877);
and U7638 (N_7638,N_6523,N_6880);
or U7639 (N_7639,N_6385,N_6784);
nor U7640 (N_7640,N_6303,N_6389);
xor U7641 (N_7641,N_6340,N_6393);
or U7642 (N_7642,N_7268,N_6211);
or U7643 (N_7643,N_6815,N_6985);
or U7644 (N_7644,N_7197,N_6933);
xnor U7645 (N_7645,N_6467,N_6194);
nor U7646 (N_7646,N_6768,N_7302);
nand U7647 (N_7647,N_7394,N_6976);
xnor U7648 (N_7648,N_6473,N_7212);
nand U7649 (N_7649,N_6553,N_6830);
nand U7650 (N_7650,N_7296,N_6168);
nor U7651 (N_7651,N_6926,N_6060);
nor U7652 (N_7652,N_6377,N_7380);
or U7653 (N_7653,N_6302,N_6475);
nand U7654 (N_7654,N_6776,N_6809);
nand U7655 (N_7655,N_6135,N_7297);
xnor U7656 (N_7656,N_6598,N_6103);
nand U7657 (N_7657,N_7050,N_7154);
or U7658 (N_7658,N_6336,N_7499);
nor U7659 (N_7659,N_6370,N_6138);
nor U7660 (N_7660,N_6993,N_6487);
nand U7661 (N_7661,N_6588,N_7266);
nand U7662 (N_7662,N_6468,N_6176);
and U7663 (N_7663,N_6856,N_6212);
xnor U7664 (N_7664,N_7051,N_6514);
nor U7665 (N_7665,N_6868,N_7455);
or U7666 (N_7666,N_6757,N_6248);
and U7667 (N_7667,N_6551,N_6665);
or U7668 (N_7668,N_6463,N_6980);
nor U7669 (N_7669,N_7213,N_7241);
nand U7670 (N_7670,N_7246,N_6650);
nand U7671 (N_7671,N_6753,N_7488);
and U7672 (N_7672,N_6699,N_6919);
or U7673 (N_7673,N_6506,N_7013);
nand U7674 (N_7674,N_6383,N_7027);
nor U7675 (N_7675,N_6395,N_7219);
nand U7676 (N_7676,N_6219,N_6444);
xor U7677 (N_7677,N_7003,N_6294);
or U7678 (N_7678,N_7267,N_7346);
or U7679 (N_7679,N_6059,N_6678);
nand U7680 (N_7680,N_7443,N_7368);
or U7681 (N_7681,N_6043,N_7068);
and U7682 (N_7682,N_6153,N_6165);
nor U7683 (N_7683,N_6373,N_7152);
and U7684 (N_7684,N_6243,N_7487);
and U7685 (N_7685,N_7402,N_7159);
nor U7686 (N_7686,N_7396,N_6561);
nor U7687 (N_7687,N_7338,N_7479);
and U7688 (N_7688,N_6694,N_6488);
and U7689 (N_7689,N_7393,N_6806);
nand U7690 (N_7690,N_7299,N_6357);
and U7691 (N_7691,N_6525,N_7000);
nand U7692 (N_7692,N_6141,N_6077);
nor U7693 (N_7693,N_7200,N_7132);
and U7694 (N_7694,N_6071,N_7130);
nand U7695 (N_7695,N_6136,N_6769);
nand U7696 (N_7696,N_7362,N_7149);
or U7697 (N_7697,N_6995,N_7327);
and U7698 (N_7698,N_6225,N_6817);
nand U7699 (N_7699,N_6083,N_7014);
nand U7700 (N_7700,N_6862,N_7122);
and U7701 (N_7701,N_6436,N_7463);
or U7702 (N_7702,N_6735,N_7363);
or U7703 (N_7703,N_6014,N_7188);
nand U7704 (N_7704,N_6948,N_7322);
nand U7705 (N_7705,N_6387,N_6170);
nor U7706 (N_7706,N_6438,N_6282);
or U7707 (N_7707,N_6610,N_7205);
or U7708 (N_7708,N_6825,N_7211);
and U7709 (N_7709,N_6752,N_6572);
or U7710 (N_7710,N_6501,N_6031);
nand U7711 (N_7711,N_6889,N_6479);
nand U7712 (N_7712,N_6736,N_6209);
nor U7713 (N_7713,N_6850,N_7454);
and U7714 (N_7714,N_6166,N_7082);
and U7715 (N_7715,N_7371,N_7289);
or U7716 (N_7716,N_6063,N_6845);
or U7717 (N_7717,N_6251,N_7251);
nand U7718 (N_7718,N_6214,N_7440);
and U7719 (N_7719,N_6207,N_6155);
nor U7720 (N_7720,N_6262,N_7234);
nand U7721 (N_7721,N_6224,N_6600);
nand U7722 (N_7722,N_6882,N_7351);
or U7723 (N_7723,N_7052,N_6593);
nor U7724 (N_7724,N_7398,N_6440);
and U7725 (N_7725,N_7292,N_6950);
and U7726 (N_7726,N_6443,N_6920);
or U7727 (N_7727,N_7030,N_6348);
nand U7728 (N_7728,N_6979,N_6205);
and U7729 (N_7729,N_6594,N_6543);
or U7730 (N_7730,N_6725,N_7383);
nand U7731 (N_7731,N_6241,N_7080);
or U7732 (N_7732,N_7262,N_7198);
and U7733 (N_7733,N_6026,N_6072);
nand U7734 (N_7734,N_7158,N_6273);
and U7735 (N_7735,N_6669,N_7084);
xnor U7736 (N_7736,N_6529,N_7049);
or U7737 (N_7737,N_6426,N_7291);
or U7738 (N_7738,N_6875,N_6639);
and U7739 (N_7739,N_7491,N_7106);
or U7740 (N_7740,N_7497,N_6379);
or U7741 (N_7741,N_7339,N_6819);
nor U7742 (N_7742,N_6361,N_6865);
nand U7743 (N_7743,N_7260,N_6788);
nand U7744 (N_7744,N_7156,N_7145);
xor U7745 (N_7745,N_6526,N_6296);
xor U7746 (N_7746,N_7350,N_7007);
or U7747 (N_7747,N_6971,N_6230);
or U7748 (N_7748,N_6550,N_6890);
nand U7749 (N_7749,N_6128,N_7281);
and U7750 (N_7750,N_6542,N_6203);
or U7751 (N_7751,N_6846,N_7435);
or U7752 (N_7752,N_7466,N_7202);
and U7753 (N_7753,N_6508,N_6967);
nor U7754 (N_7754,N_6690,N_6082);
nand U7755 (N_7755,N_7066,N_6419);
and U7756 (N_7756,N_7284,N_6022);
or U7757 (N_7757,N_7046,N_6777);
nand U7758 (N_7758,N_6897,N_6765);
or U7759 (N_7759,N_7025,N_6642);
nand U7760 (N_7760,N_6781,N_6558);
or U7761 (N_7761,N_6750,N_6486);
xor U7762 (N_7762,N_7388,N_6300);
or U7763 (N_7763,N_7319,N_6935);
or U7764 (N_7764,N_6963,N_7153);
xor U7765 (N_7765,N_7254,N_6187);
nor U7766 (N_7766,N_6530,N_6456);
or U7767 (N_7767,N_7385,N_6726);
and U7768 (N_7768,N_6354,N_6672);
xor U7769 (N_7769,N_7181,N_6078);
and U7770 (N_7770,N_7175,N_6886);
nand U7771 (N_7771,N_6006,N_7459);
xnor U7772 (N_7772,N_7377,N_6140);
and U7773 (N_7773,N_7273,N_7083);
nand U7774 (N_7774,N_7218,N_7473);
and U7775 (N_7775,N_6420,N_6869);
nor U7776 (N_7776,N_6625,N_6763);
nand U7777 (N_7777,N_6023,N_6941);
or U7778 (N_7778,N_6423,N_7476);
or U7779 (N_7779,N_6156,N_7438);
nor U7780 (N_7780,N_6459,N_7340);
nor U7781 (N_7781,N_7177,N_7043);
and U7782 (N_7782,N_6547,N_7418);
and U7783 (N_7783,N_6791,N_6872);
nor U7784 (N_7784,N_6493,N_6533);
and U7785 (N_7785,N_6490,N_7102);
and U7786 (N_7786,N_6091,N_7471);
nor U7787 (N_7787,N_6064,N_6498);
or U7788 (N_7788,N_6366,N_6305);
nand U7789 (N_7789,N_7467,N_7180);
nor U7790 (N_7790,N_7120,N_6536);
xor U7791 (N_7791,N_6306,N_6685);
nand U7792 (N_7792,N_7108,N_6283);
or U7793 (N_7793,N_6062,N_6364);
nor U7794 (N_7794,N_6772,N_6111);
nor U7795 (N_7795,N_6144,N_6076);
and U7796 (N_7796,N_7121,N_6937);
or U7797 (N_7797,N_6386,N_6005);
or U7798 (N_7798,N_7411,N_6312);
or U7799 (N_7799,N_6421,N_7345);
nand U7800 (N_7800,N_7464,N_6925);
and U7801 (N_7801,N_6712,N_7323);
nand U7802 (N_7802,N_7064,N_6818);
nor U7803 (N_7803,N_6604,N_6019);
nor U7804 (N_7804,N_6635,N_7240);
and U7805 (N_7805,N_6570,N_7428);
nor U7806 (N_7806,N_6268,N_7230);
nor U7807 (N_7807,N_6974,N_6097);
and U7808 (N_7808,N_6126,N_6671);
nand U7809 (N_7809,N_6794,N_7493);
or U7810 (N_7810,N_7436,N_7494);
nand U7811 (N_7811,N_7235,N_7330);
or U7812 (N_7812,N_6380,N_6399);
nand U7813 (N_7813,N_6199,N_6198);
or U7814 (N_7814,N_6325,N_6962);
or U7815 (N_7815,N_6066,N_7375);
nor U7816 (N_7816,N_6881,N_7278);
nor U7817 (N_7817,N_6775,N_7392);
xnor U7818 (N_7818,N_7199,N_7193);
or U7819 (N_7819,N_6374,N_7002);
nor U7820 (N_7820,N_6108,N_6762);
or U7821 (N_7821,N_6645,N_6367);
xor U7822 (N_7822,N_7404,N_7495);
or U7823 (N_7823,N_6052,N_7264);
nand U7824 (N_7824,N_7352,N_6322);
and U7825 (N_7825,N_7307,N_6044);
nand U7826 (N_7826,N_6109,N_7217);
xnor U7827 (N_7827,N_7075,N_6040);
or U7828 (N_7828,N_6160,N_7444);
or U7829 (N_7829,N_6427,N_6587);
nor U7830 (N_7830,N_6319,N_7209);
or U7831 (N_7831,N_6069,N_6359);
nor U7832 (N_7832,N_7333,N_6532);
nand U7833 (N_7833,N_7127,N_7184);
and U7834 (N_7834,N_6027,N_6576);
nand U7835 (N_7835,N_6855,N_6095);
nand U7836 (N_7836,N_7185,N_6901);
nand U7837 (N_7837,N_7135,N_6231);
and U7838 (N_7838,N_6519,N_7400);
nand U7839 (N_7839,N_6058,N_7225);
nor U7840 (N_7840,N_7486,N_6308);
nand U7841 (N_7841,N_6535,N_6864);
nand U7842 (N_7842,N_6793,N_6249);
nor U7843 (N_7843,N_7017,N_6255);
or U7844 (N_7844,N_6958,N_7335);
or U7845 (N_7845,N_6464,N_6049);
nand U7846 (N_7846,N_6481,N_6816);
and U7847 (N_7847,N_6676,N_6117);
and U7848 (N_7848,N_6313,N_6801);
or U7849 (N_7849,N_6988,N_6437);
xor U7850 (N_7850,N_6133,N_7356);
and U7851 (N_7851,N_6622,N_6729);
nand U7852 (N_7852,N_6964,N_7353);
or U7853 (N_7853,N_7059,N_6698);
nand U7854 (N_7854,N_7477,N_7168);
nand U7855 (N_7855,N_7354,N_6191);
or U7856 (N_7856,N_6706,N_6887);
nor U7857 (N_7857,N_6422,N_6840);
and U7858 (N_7858,N_7370,N_7206);
or U7859 (N_7859,N_6264,N_7160);
nor U7860 (N_7860,N_7274,N_6579);
xnor U7861 (N_7861,N_7415,N_6431);
nand U7862 (N_7862,N_7306,N_6280);
or U7863 (N_7863,N_6042,N_6822);
nor U7864 (N_7864,N_6990,N_6973);
or U7865 (N_7865,N_7147,N_6918);
or U7866 (N_7866,N_6039,N_6057);
or U7867 (N_7867,N_6106,N_7221);
and U7868 (N_7868,N_6883,N_6000);
xnor U7869 (N_7869,N_7290,N_6316);
nand U7870 (N_7870,N_6402,N_6837);
xor U7871 (N_7871,N_6293,N_6917);
and U7872 (N_7872,N_6414,N_6037);
and U7873 (N_7873,N_6998,N_6606);
xor U7874 (N_7874,N_6708,N_7196);
and U7875 (N_7875,N_6311,N_6157);
or U7876 (N_7876,N_6124,N_7419);
and U7877 (N_7877,N_6720,N_7134);
nor U7878 (N_7878,N_7063,N_6952);
nor U7879 (N_7879,N_7379,N_6267);
nor U7880 (N_7880,N_6343,N_6461);
xnor U7881 (N_7881,N_6216,N_6152);
nor U7882 (N_7882,N_6798,N_6276);
or U7883 (N_7883,N_6586,N_6093);
or U7884 (N_7884,N_6299,N_7142);
or U7885 (N_7885,N_7484,N_6175);
nor U7886 (N_7886,N_6256,N_7239);
nand U7887 (N_7887,N_6323,N_6183);
xnor U7888 (N_7888,N_6240,N_6749);
or U7889 (N_7889,N_6943,N_6629);
nand U7890 (N_7890,N_6200,N_6193);
or U7891 (N_7891,N_6252,N_6045);
or U7892 (N_7892,N_6709,N_7207);
nand U7893 (N_7893,N_6700,N_6289);
nor U7894 (N_7894,N_7277,N_7250);
nand U7895 (N_7895,N_7141,N_6446);
xor U7896 (N_7896,N_6342,N_7062);
nand U7897 (N_7897,N_6274,N_6945);
or U7898 (N_7898,N_6566,N_6349);
nand U7899 (N_7899,N_7332,N_7403);
or U7900 (N_7900,N_6658,N_6292);
nor U7901 (N_7901,N_6397,N_6208);
xor U7902 (N_7902,N_6792,N_7016);
xnor U7903 (N_7903,N_6391,N_6070);
nand U7904 (N_7904,N_7412,N_7107);
and U7905 (N_7905,N_6732,N_7261);
nand U7906 (N_7906,N_6120,N_6286);
or U7907 (N_7907,N_6384,N_6655);
nor U7908 (N_7908,N_7431,N_6496);
nor U7909 (N_7909,N_7155,N_7328);
nand U7910 (N_7910,N_7294,N_7416);
nor U7911 (N_7911,N_7163,N_6400);
nor U7912 (N_7912,N_7243,N_6489);
or U7913 (N_7913,N_6584,N_6253);
or U7914 (N_7914,N_7090,N_6719);
nor U7915 (N_7915,N_7058,N_6876);
nand U7916 (N_7916,N_6773,N_6782);
or U7917 (N_7917,N_6592,N_6304);
or U7918 (N_7918,N_6670,N_7252);
nand U7919 (N_7919,N_6954,N_7161);
nand U7920 (N_7920,N_6582,N_7458);
nand U7921 (N_7921,N_7426,N_7365);
xnor U7922 (N_7922,N_6016,N_6186);
or U7923 (N_7923,N_7001,N_6404);
and U7924 (N_7924,N_6465,N_6754);
nand U7925 (N_7925,N_6991,N_6067);
or U7926 (N_7926,N_6279,N_6618);
nor U7927 (N_7927,N_6314,N_6915);
xnor U7928 (N_7928,N_7405,N_6693);
and U7929 (N_7929,N_7378,N_6531);
nor U7930 (N_7930,N_6651,N_7138);
and U7931 (N_7931,N_7304,N_6272);
and U7932 (N_7932,N_6767,N_6250);
or U7933 (N_7933,N_6148,N_6223);
nand U7934 (N_7934,N_7280,N_6024);
or U7935 (N_7935,N_6583,N_7139);
or U7936 (N_7936,N_6608,N_6457);
or U7937 (N_7937,N_6664,N_7490);
and U7938 (N_7938,N_7395,N_7097);
and U7939 (N_7939,N_6679,N_6774);
nand U7940 (N_7940,N_6647,N_6521);
nand U7941 (N_7941,N_7437,N_6951);
and U7942 (N_7942,N_7110,N_6546);
nand U7943 (N_7943,N_7167,N_7100);
and U7944 (N_7944,N_7343,N_6737);
and U7945 (N_7945,N_6226,N_6730);
nor U7946 (N_7946,N_7407,N_7325);
xor U7947 (N_7947,N_6260,N_7074);
or U7948 (N_7948,N_7451,N_7079);
or U7949 (N_7949,N_6873,N_7287);
and U7950 (N_7950,N_6346,N_6620);
or U7951 (N_7951,N_6764,N_6127);
and U7952 (N_7952,N_6329,N_6758);
and U7953 (N_7953,N_6567,N_6032);
or U7954 (N_7954,N_6871,N_6910);
and U7955 (N_7955,N_7229,N_6717);
nand U7956 (N_7956,N_6739,N_7109);
and U7957 (N_7957,N_7057,N_7171);
and U7958 (N_7958,N_6245,N_7111);
xnor U7959 (N_7959,N_6167,N_6151);
nor U7960 (N_7960,N_6646,N_7040);
nor U7961 (N_7961,N_7093,N_6644);
nor U7962 (N_7962,N_6966,N_6957);
xnor U7963 (N_7963,N_6376,N_6527);
nand U7964 (N_7964,N_6595,N_6430);
or U7965 (N_7965,N_7316,N_6482);
nand U7966 (N_7966,N_6334,N_6724);
nand U7967 (N_7967,N_6703,N_7092);
nand U7968 (N_7968,N_7498,N_7008);
nand U7969 (N_7969,N_7429,N_6320);
nand U7970 (N_7970,N_6017,N_7019);
nand U7971 (N_7971,N_6164,N_6331);
nand U7972 (N_7972,N_6025,N_6537);
or U7973 (N_7973,N_6080,N_6913);
and U7974 (N_7974,N_7430,N_6803);
nand U7975 (N_7975,N_6450,N_6181);
or U7976 (N_7976,N_6474,N_7483);
nand U7977 (N_7977,N_7298,N_7245);
or U7978 (N_7978,N_6053,N_7157);
and U7979 (N_7979,N_7481,N_6623);
and U7980 (N_7980,N_6929,N_6921);
or U7981 (N_7981,N_6001,N_7423);
or U7982 (N_7982,N_6820,N_6900);
and U7983 (N_7983,N_7087,N_6073);
and U7984 (N_7984,N_6184,N_6518);
xor U7985 (N_7985,N_7237,N_6824);
and U7986 (N_7986,N_7112,N_6949);
nand U7987 (N_7987,N_6778,N_6756);
or U7988 (N_7988,N_7421,N_6137);
and U7989 (N_7989,N_7453,N_6254);
or U7990 (N_7990,N_6826,N_7236);
or U7991 (N_7991,N_6038,N_7265);
nor U7992 (N_7992,N_6562,N_7144);
xor U7993 (N_7993,N_7047,N_6335);
or U7994 (N_7994,N_6477,N_7006);
and U7995 (N_7995,N_7293,N_7427);
nor U7996 (N_7996,N_6641,N_6163);
or U7997 (N_7997,N_6497,N_6134);
nand U7998 (N_7998,N_6494,N_6372);
xor U7999 (N_7999,N_6843,N_7329);
nor U8000 (N_8000,N_7269,N_7233);
or U8001 (N_8001,N_6147,N_6020);
nor U8002 (N_8002,N_7073,N_6761);
and U8003 (N_8003,N_6054,N_7373);
or U8004 (N_8004,N_7347,N_6984);
and U8005 (N_8005,N_6033,N_7131);
or U8006 (N_8006,N_6682,N_6740);
xor U8007 (N_8007,N_6502,N_7117);
nand U8008 (N_8008,N_6310,N_6723);
or U8009 (N_8009,N_6805,N_6295);
or U8010 (N_8010,N_6649,N_6206);
or U8011 (N_8011,N_7341,N_6347);
nor U8012 (N_8012,N_6515,N_6110);
and U8013 (N_8013,N_6891,N_6088);
and U8014 (N_8014,N_6728,N_7039);
or U8015 (N_8015,N_6192,N_7420);
or U8016 (N_8016,N_7035,N_7029);
nand U8017 (N_8017,N_7314,N_6989);
and U8018 (N_8018,N_6857,N_7256);
nor U8019 (N_8019,N_6333,N_6290);
nand U8020 (N_8020,N_6125,N_7037);
xnor U8021 (N_8021,N_7096,N_6451);
nand U8022 (N_8022,N_6895,N_7406);
and U8023 (N_8023,N_6522,N_6114);
xnor U8024 (N_8024,N_7258,N_6180);
or U8025 (N_8025,N_6999,N_6204);
nor U8026 (N_8026,N_6096,N_7417);
nor U8027 (N_8027,N_7465,N_7271);
nor U8028 (N_8028,N_6086,N_7248);
nor U8029 (N_8029,N_6548,N_6834);
nor U8030 (N_8030,N_6119,N_7372);
nor U8031 (N_8031,N_6326,N_6858);
or U8032 (N_8032,N_6909,N_6178);
and U8033 (N_8033,N_7446,N_7176);
and U8034 (N_8034,N_7492,N_7320);
or U8035 (N_8035,N_6590,N_6634);
xor U8036 (N_8036,N_6842,N_7143);
nand U8037 (N_8037,N_6406,N_6257);
and U8038 (N_8038,N_7067,N_6955);
and U8039 (N_8039,N_6416,N_6603);
nor U8040 (N_8040,N_7033,N_7091);
and U8041 (N_8041,N_6055,N_6242);
xor U8042 (N_8042,N_6557,N_7358);
xnor U8043 (N_8043,N_6970,N_6571);
and U8044 (N_8044,N_6983,N_6079);
nor U8045 (N_8045,N_7263,N_6131);
xnor U8046 (N_8046,N_6986,N_6554);
and U8047 (N_8047,N_7081,N_6599);
nand U8048 (N_8048,N_6823,N_6378);
nor U8049 (N_8049,N_6394,N_6663);
nor U8050 (N_8050,N_6747,N_7285);
or U8051 (N_8051,N_6130,N_7169);
nand U8052 (N_8052,N_7445,N_7300);
and U8053 (N_8053,N_7334,N_7103);
and U8054 (N_8054,N_7374,N_7070);
and U8055 (N_8055,N_6931,N_6927);
xor U8056 (N_8056,N_6142,N_6013);
or U8057 (N_8057,N_7098,N_6261);
nor U8058 (N_8058,N_6624,N_6539);
nor U8059 (N_8059,N_6666,N_7390);
nor U8060 (N_8060,N_6332,N_7389);
or U8061 (N_8061,N_6266,N_6353);
nand U8062 (N_8062,N_6448,N_6716);
xnor U8063 (N_8063,N_6630,N_6388);
or U8064 (N_8064,N_6923,N_7452);
or U8065 (N_8065,N_7065,N_7442);
nor U8066 (N_8066,N_7413,N_6617);
nor U8067 (N_8067,N_6433,N_7187);
nor U8068 (N_8068,N_6034,N_7391);
and U8069 (N_8069,N_7086,N_6691);
xor U8070 (N_8070,N_6432,N_7305);
nand U8071 (N_8071,N_7023,N_7317);
nor U8072 (N_8072,N_6509,N_6491);
or U8073 (N_8073,N_7010,N_6345);
nand U8074 (N_8074,N_7077,N_6454);
or U8075 (N_8075,N_7222,N_6863);
or U8076 (N_8076,N_6428,N_6520);
xor U8077 (N_8077,N_6721,N_6545);
xor U8078 (N_8078,N_7178,N_6185);
xnor U8079 (N_8079,N_6939,N_6689);
nor U8080 (N_8080,N_7045,N_6270);
and U8081 (N_8081,N_6048,N_6619);
nand U8082 (N_8082,N_6263,N_6968);
nor U8083 (N_8083,N_6849,N_6994);
nor U8084 (N_8084,N_6879,N_6500);
nand U8085 (N_8085,N_6540,N_6162);
or U8086 (N_8086,N_7303,N_6969);
xor U8087 (N_8087,N_7088,N_7227);
nand U8088 (N_8088,N_7295,N_6466);
nand U8089 (N_8089,N_6177,N_6959);
and U8090 (N_8090,N_7357,N_6041);
and U8091 (N_8091,N_7449,N_6236);
nand U8092 (N_8092,N_7034,N_6470);
and U8093 (N_8093,N_7272,N_7318);
or U8094 (N_8094,N_6411,N_7469);
nor U8095 (N_8095,N_7433,N_6030);
nand U8096 (N_8096,N_6960,N_7094);
nand U8097 (N_8097,N_7165,N_6615);
and U8098 (N_8098,N_6173,N_7036);
or U8099 (N_8099,N_6235,N_7041);
nor U8100 (N_8100,N_6356,N_7247);
and U8101 (N_8101,N_6453,N_6643);
xor U8102 (N_8102,N_7439,N_7208);
xnor U8103 (N_8103,N_6621,N_6696);
nand U8104 (N_8104,N_7022,N_6287);
nand U8105 (N_8105,N_6171,N_6050);
or U8106 (N_8106,N_6405,N_6835);
and U8107 (N_8107,N_7276,N_6190);
or U8108 (N_8108,N_6085,N_6673);
or U8109 (N_8109,N_6677,N_6555);
and U8110 (N_8110,N_6702,N_6369);
xnor U8111 (N_8111,N_7401,N_6201);
nand U8112 (N_8112,N_6870,N_7164);
nor U8113 (N_8113,N_7172,N_7182);
nor U8114 (N_8114,N_7099,N_6439);
nand U8115 (N_8115,N_6195,N_6102);
nand U8116 (N_8116,N_6814,N_6659);
nor U8117 (N_8117,N_6785,N_6321);
nor U8118 (N_8118,N_7409,N_6341);
xor U8119 (N_8119,N_6888,N_6107);
xor U8120 (N_8120,N_7186,N_7270);
or U8121 (N_8121,N_6564,N_6829);
nand U8122 (N_8122,N_7031,N_6591);
xnor U8123 (N_8123,N_7183,N_7462);
and U8124 (N_8124,N_6099,N_7053);
and U8125 (N_8125,N_6853,N_6731);
nor U8126 (N_8126,N_7482,N_6218);
and U8127 (N_8127,N_6575,N_7282);
nand U8128 (N_8128,N_7312,N_6172);
or U8129 (N_8129,N_6987,N_6742);
and U8130 (N_8130,N_6848,N_7069);
and U8131 (N_8131,N_6911,N_6116);
xnor U8132 (N_8132,N_6258,N_6903);
and U8133 (N_8133,N_7414,N_6859);
nor U8134 (N_8134,N_6100,N_6188);
xnor U8135 (N_8135,N_6247,N_6445);
or U8136 (N_8136,N_7382,N_6799);
and U8137 (N_8137,N_6118,N_6811);
and U8138 (N_8138,N_7275,N_6596);
nor U8139 (N_8139,N_6574,N_6637);
and U8140 (N_8140,N_6680,N_6429);
xor U8141 (N_8141,N_6113,N_6301);
and U8142 (N_8142,N_7009,N_7085);
and U8143 (N_8143,N_6552,N_7024);
or U8144 (N_8144,N_6580,N_6790);
or U8145 (N_8145,N_6472,N_7072);
or U8146 (N_8146,N_6307,N_7461);
nor U8147 (N_8147,N_6906,N_6648);
nor U8148 (N_8148,N_6874,N_6478);
nor U8149 (N_8149,N_6495,N_7020);
or U8150 (N_8150,N_6046,N_6766);
nor U8151 (N_8151,N_6363,N_7397);
and U8152 (N_8152,N_6896,N_6755);
nand U8153 (N_8153,N_6847,N_6449);
or U8154 (N_8154,N_7190,N_6315);
xnor U8155 (N_8155,N_7472,N_6035);
xor U8156 (N_8156,N_6317,N_7151);
and U8157 (N_8157,N_6759,N_6894);
or U8158 (N_8158,N_7228,N_6714);
and U8159 (N_8159,N_6011,N_6654);
xnor U8160 (N_8160,N_6410,N_7028);
xnor U8161 (N_8161,N_6121,N_7432);
and U8162 (N_8162,N_6961,N_6833);
nor U8163 (N_8163,N_6741,N_6009);
and U8164 (N_8164,N_6981,N_7105);
and U8165 (N_8165,N_6297,N_6018);
and U8166 (N_8166,N_7448,N_6710);
nand U8167 (N_8167,N_6221,N_6812);
nand U8168 (N_8168,N_6938,N_6396);
nand U8169 (N_8169,N_7348,N_6878);
and U8170 (N_8170,N_6417,N_6907);
and U8171 (N_8171,N_6975,N_6965);
nor U8172 (N_8172,N_6232,N_7450);
xnor U8173 (N_8173,N_6707,N_6075);
nor U8174 (N_8174,N_6051,N_7384);
nor U8175 (N_8175,N_6246,N_7214);
nor U8176 (N_8176,N_6780,N_6511);
or U8177 (N_8177,N_6786,N_6344);
xor U8178 (N_8178,N_6627,N_6705);
or U8179 (N_8179,N_6089,N_7489);
nand U8180 (N_8180,N_6339,N_6318);
nand U8181 (N_8181,N_7308,N_6360);
nand U8182 (N_8182,N_6795,N_6569);
and U8183 (N_8183,N_6854,N_6434);
nand U8184 (N_8184,N_7238,N_6573);
and U8185 (N_8185,N_6867,N_6159);
nor U8186 (N_8186,N_6084,N_6953);
nor U8187 (N_8187,N_6704,N_6841);
or U8188 (N_8188,N_6139,N_6559);
nor U8189 (N_8189,N_7349,N_7095);
xnor U8190 (N_8190,N_6827,N_6408);
nand U8191 (N_8191,N_7232,N_6007);
or U8192 (N_8192,N_6174,N_7355);
nand U8193 (N_8193,N_7150,N_6578);
xnor U8194 (N_8194,N_7309,N_6278);
nand U8195 (N_8195,N_6565,N_7191);
nand U8196 (N_8196,N_7042,N_6112);
and U8197 (N_8197,N_6492,N_6652);
or U8198 (N_8198,N_6924,N_7457);
nand U8199 (N_8199,N_6549,N_7204);
and U8200 (N_8200,N_6413,N_6094);
nor U8201 (N_8201,N_6885,N_7231);
xnor U8202 (N_8202,N_6899,N_7060);
nor U8203 (N_8203,N_6893,N_6844);
nand U8204 (N_8204,N_6605,N_7061);
and U8205 (N_8205,N_6972,N_7259);
nor U8206 (N_8206,N_6674,N_6611);
and U8207 (N_8207,N_7387,N_6355);
xnor U8208 (N_8208,N_6956,N_6090);
nand U8209 (N_8209,N_6480,N_6115);
nand U8210 (N_8210,N_6271,N_6944);
nand U8211 (N_8211,N_6503,N_6368);
nor U8212 (N_8212,N_7361,N_6382);
nand U8213 (N_8213,N_6779,N_7408);
or U8214 (N_8214,N_7032,N_7201);
nand U8215 (N_8215,N_6284,N_6202);
and U8216 (N_8216,N_6469,N_6743);
xor U8217 (N_8217,N_6839,N_7424);
nand U8218 (N_8218,N_6381,N_6667);
and U8219 (N_8219,N_7026,N_6711);
nand U8220 (N_8220,N_6597,N_6447);
nor U8221 (N_8221,N_6701,N_6783);
nor U8222 (N_8222,N_6056,N_6327);
nand U8223 (N_8223,N_7470,N_7129);
and U8224 (N_8224,N_6415,N_6697);
nand U8225 (N_8225,N_7326,N_6810);
nor U8226 (N_8226,N_6930,N_6143);
or U8227 (N_8227,N_6688,N_7021);
nor U8228 (N_8228,N_7133,N_6538);
nand U8229 (N_8229,N_7011,N_6244);
or U8230 (N_8230,N_6061,N_6412);
nand U8231 (N_8231,N_7242,N_7255);
and U8232 (N_8232,N_6821,N_6512);
xor U8233 (N_8233,N_7005,N_7173);
or U8234 (N_8234,N_6947,N_6277);
xor U8235 (N_8235,N_7342,N_6616);
nand U8236 (N_8236,N_6734,N_7166);
or U8237 (N_8237,N_6733,N_6861);
and U8238 (N_8238,N_6687,N_6222);
and U8239 (N_8239,N_6403,N_6285);
xnor U8240 (N_8240,N_7054,N_6441);
xnor U8241 (N_8241,N_6458,N_6727);
or U8242 (N_8242,N_7203,N_6029);
or U8243 (N_8243,N_6371,N_6504);
xnor U8244 (N_8244,N_7331,N_7468);
nand U8245 (N_8245,N_7460,N_7170);
xnor U8246 (N_8246,N_6940,N_6802);
nand U8247 (N_8247,N_6146,N_6992);
xnor U8248 (N_8248,N_6695,N_6614);
and U8249 (N_8249,N_6213,N_6656);
and U8250 (N_8250,N_6061,N_6337);
or U8251 (N_8251,N_6618,N_6510);
and U8252 (N_8252,N_7458,N_7439);
or U8253 (N_8253,N_7306,N_7493);
or U8254 (N_8254,N_6161,N_7335);
or U8255 (N_8255,N_7328,N_6361);
and U8256 (N_8256,N_6704,N_7494);
nor U8257 (N_8257,N_7161,N_6027);
or U8258 (N_8258,N_6852,N_6709);
or U8259 (N_8259,N_7436,N_6773);
nand U8260 (N_8260,N_6855,N_6984);
or U8261 (N_8261,N_7270,N_7397);
nor U8262 (N_8262,N_6122,N_7462);
and U8263 (N_8263,N_6826,N_6338);
nor U8264 (N_8264,N_6289,N_7257);
and U8265 (N_8265,N_6814,N_7492);
and U8266 (N_8266,N_7323,N_6319);
nand U8267 (N_8267,N_6846,N_7294);
nor U8268 (N_8268,N_6522,N_6899);
nand U8269 (N_8269,N_6799,N_6164);
and U8270 (N_8270,N_7370,N_7193);
or U8271 (N_8271,N_7433,N_6610);
xnor U8272 (N_8272,N_7214,N_6676);
and U8273 (N_8273,N_6529,N_6585);
and U8274 (N_8274,N_7275,N_6655);
nor U8275 (N_8275,N_7247,N_6427);
and U8276 (N_8276,N_7193,N_7211);
nand U8277 (N_8277,N_7282,N_6121);
nand U8278 (N_8278,N_7169,N_6615);
nand U8279 (N_8279,N_7391,N_6049);
nor U8280 (N_8280,N_6165,N_6928);
xnor U8281 (N_8281,N_6767,N_6406);
nand U8282 (N_8282,N_6341,N_7011);
nand U8283 (N_8283,N_6983,N_7361);
or U8284 (N_8284,N_6967,N_6568);
or U8285 (N_8285,N_6350,N_6495);
and U8286 (N_8286,N_6526,N_6352);
nor U8287 (N_8287,N_6026,N_6832);
and U8288 (N_8288,N_6596,N_6044);
or U8289 (N_8289,N_6206,N_6587);
and U8290 (N_8290,N_6272,N_6882);
or U8291 (N_8291,N_6061,N_7067);
nor U8292 (N_8292,N_6619,N_6146);
nor U8293 (N_8293,N_7154,N_6023);
nor U8294 (N_8294,N_6057,N_7151);
and U8295 (N_8295,N_6824,N_6609);
nand U8296 (N_8296,N_6183,N_7013);
nor U8297 (N_8297,N_6534,N_6204);
xor U8298 (N_8298,N_6283,N_6757);
nand U8299 (N_8299,N_6621,N_7016);
and U8300 (N_8300,N_6441,N_6523);
or U8301 (N_8301,N_6980,N_6776);
or U8302 (N_8302,N_6783,N_6444);
and U8303 (N_8303,N_7163,N_6675);
nand U8304 (N_8304,N_6157,N_6645);
nor U8305 (N_8305,N_7138,N_7319);
and U8306 (N_8306,N_6013,N_7195);
or U8307 (N_8307,N_6046,N_6620);
or U8308 (N_8308,N_6916,N_7004);
nor U8309 (N_8309,N_7233,N_7489);
nor U8310 (N_8310,N_6180,N_7296);
xnor U8311 (N_8311,N_6592,N_6445);
and U8312 (N_8312,N_6884,N_6279);
or U8313 (N_8313,N_6511,N_6106);
nor U8314 (N_8314,N_7334,N_6117);
nand U8315 (N_8315,N_6312,N_6023);
and U8316 (N_8316,N_6270,N_6229);
or U8317 (N_8317,N_6076,N_6688);
nand U8318 (N_8318,N_6721,N_6029);
nor U8319 (N_8319,N_7383,N_6068);
nand U8320 (N_8320,N_7237,N_7058);
and U8321 (N_8321,N_6832,N_7064);
xor U8322 (N_8322,N_7056,N_7167);
nand U8323 (N_8323,N_7218,N_7396);
nor U8324 (N_8324,N_7099,N_6509);
and U8325 (N_8325,N_6272,N_6321);
and U8326 (N_8326,N_6012,N_6464);
nor U8327 (N_8327,N_7236,N_6025);
and U8328 (N_8328,N_7082,N_6907);
and U8329 (N_8329,N_6384,N_6919);
nor U8330 (N_8330,N_6548,N_6678);
nand U8331 (N_8331,N_6570,N_6381);
and U8332 (N_8332,N_6775,N_6373);
nor U8333 (N_8333,N_7136,N_6401);
nand U8334 (N_8334,N_6282,N_6296);
xnor U8335 (N_8335,N_7150,N_6491);
or U8336 (N_8336,N_6186,N_6863);
nor U8337 (N_8337,N_6377,N_6159);
and U8338 (N_8338,N_7172,N_6115);
xor U8339 (N_8339,N_6937,N_7062);
or U8340 (N_8340,N_6254,N_6919);
nor U8341 (N_8341,N_7422,N_7246);
xor U8342 (N_8342,N_6157,N_6032);
nor U8343 (N_8343,N_6810,N_7480);
or U8344 (N_8344,N_6639,N_7471);
and U8345 (N_8345,N_6464,N_6942);
nand U8346 (N_8346,N_6452,N_7065);
xnor U8347 (N_8347,N_7412,N_7097);
nor U8348 (N_8348,N_7288,N_6555);
and U8349 (N_8349,N_6443,N_6134);
nor U8350 (N_8350,N_7186,N_7334);
nor U8351 (N_8351,N_7280,N_6656);
or U8352 (N_8352,N_6391,N_7423);
nand U8353 (N_8353,N_6220,N_6381);
and U8354 (N_8354,N_6118,N_7441);
or U8355 (N_8355,N_7223,N_7350);
and U8356 (N_8356,N_7440,N_6675);
or U8357 (N_8357,N_6442,N_6888);
xor U8358 (N_8358,N_7229,N_6461);
or U8359 (N_8359,N_6461,N_7482);
and U8360 (N_8360,N_6837,N_6290);
nor U8361 (N_8361,N_6454,N_6020);
nor U8362 (N_8362,N_6625,N_6843);
and U8363 (N_8363,N_6955,N_7243);
nand U8364 (N_8364,N_7087,N_6671);
or U8365 (N_8365,N_7365,N_6342);
or U8366 (N_8366,N_6792,N_6742);
nand U8367 (N_8367,N_6998,N_7431);
xor U8368 (N_8368,N_6951,N_7134);
and U8369 (N_8369,N_7024,N_6934);
nand U8370 (N_8370,N_7014,N_7004);
and U8371 (N_8371,N_7258,N_7310);
nor U8372 (N_8372,N_7211,N_6497);
and U8373 (N_8373,N_6145,N_7293);
and U8374 (N_8374,N_6143,N_6368);
nor U8375 (N_8375,N_6138,N_7039);
or U8376 (N_8376,N_7079,N_6688);
or U8377 (N_8377,N_6272,N_7284);
or U8378 (N_8378,N_6025,N_7096);
nand U8379 (N_8379,N_6344,N_6443);
nand U8380 (N_8380,N_6319,N_6738);
nor U8381 (N_8381,N_6350,N_6866);
or U8382 (N_8382,N_6030,N_7083);
xnor U8383 (N_8383,N_6574,N_7441);
nand U8384 (N_8384,N_6664,N_6235);
and U8385 (N_8385,N_6794,N_6792);
nand U8386 (N_8386,N_6301,N_7292);
or U8387 (N_8387,N_6852,N_6310);
nor U8388 (N_8388,N_7304,N_6269);
nand U8389 (N_8389,N_6567,N_7308);
nand U8390 (N_8390,N_7233,N_7190);
nand U8391 (N_8391,N_6632,N_6895);
and U8392 (N_8392,N_7248,N_6506);
or U8393 (N_8393,N_6778,N_6677);
and U8394 (N_8394,N_7109,N_7466);
and U8395 (N_8395,N_6631,N_7427);
and U8396 (N_8396,N_6960,N_7421);
or U8397 (N_8397,N_7011,N_6848);
nor U8398 (N_8398,N_6791,N_6649);
or U8399 (N_8399,N_7395,N_6349);
or U8400 (N_8400,N_7032,N_6465);
xnor U8401 (N_8401,N_7445,N_6596);
nor U8402 (N_8402,N_6233,N_7493);
nor U8403 (N_8403,N_6201,N_6656);
or U8404 (N_8404,N_6023,N_6903);
nor U8405 (N_8405,N_7377,N_6892);
nor U8406 (N_8406,N_7282,N_7306);
nor U8407 (N_8407,N_6412,N_6133);
and U8408 (N_8408,N_7497,N_6450);
and U8409 (N_8409,N_6147,N_6896);
nand U8410 (N_8410,N_7260,N_6900);
and U8411 (N_8411,N_6156,N_6829);
and U8412 (N_8412,N_6584,N_6186);
xor U8413 (N_8413,N_7152,N_6838);
nand U8414 (N_8414,N_7188,N_6415);
nand U8415 (N_8415,N_6908,N_6607);
or U8416 (N_8416,N_6697,N_7398);
and U8417 (N_8417,N_6129,N_7314);
or U8418 (N_8418,N_6643,N_6488);
and U8419 (N_8419,N_7464,N_6728);
and U8420 (N_8420,N_7187,N_7064);
nand U8421 (N_8421,N_6531,N_6286);
nor U8422 (N_8422,N_7148,N_6164);
and U8423 (N_8423,N_6260,N_7080);
nor U8424 (N_8424,N_6223,N_6011);
or U8425 (N_8425,N_7000,N_6865);
nor U8426 (N_8426,N_7375,N_7451);
or U8427 (N_8427,N_6076,N_6171);
nand U8428 (N_8428,N_7259,N_6559);
xnor U8429 (N_8429,N_6288,N_6761);
and U8430 (N_8430,N_7404,N_6602);
nor U8431 (N_8431,N_7440,N_6728);
xnor U8432 (N_8432,N_7044,N_6794);
and U8433 (N_8433,N_6781,N_6673);
nand U8434 (N_8434,N_6418,N_6588);
nor U8435 (N_8435,N_6009,N_7267);
nand U8436 (N_8436,N_7376,N_6151);
or U8437 (N_8437,N_6057,N_7233);
nor U8438 (N_8438,N_6881,N_6615);
nor U8439 (N_8439,N_6179,N_7136);
or U8440 (N_8440,N_6353,N_7129);
nor U8441 (N_8441,N_6106,N_7195);
nand U8442 (N_8442,N_7290,N_6857);
nand U8443 (N_8443,N_7010,N_6632);
nand U8444 (N_8444,N_7311,N_6854);
xnor U8445 (N_8445,N_6197,N_7221);
and U8446 (N_8446,N_6617,N_6634);
xnor U8447 (N_8447,N_6186,N_6775);
xor U8448 (N_8448,N_6563,N_6017);
nand U8449 (N_8449,N_6141,N_7243);
or U8450 (N_8450,N_6900,N_6692);
nand U8451 (N_8451,N_7220,N_6659);
nand U8452 (N_8452,N_6496,N_6337);
and U8453 (N_8453,N_6604,N_6775);
xor U8454 (N_8454,N_7338,N_7056);
and U8455 (N_8455,N_6416,N_6033);
nand U8456 (N_8456,N_6546,N_6248);
or U8457 (N_8457,N_6884,N_6409);
nor U8458 (N_8458,N_6463,N_6255);
nand U8459 (N_8459,N_7178,N_7238);
nand U8460 (N_8460,N_6157,N_6209);
or U8461 (N_8461,N_7335,N_6207);
and U8462 (N_8462,N_6855,N_6093);
or U8463 (N_8463,N_6334,N_6378);
xnor U8464 (N_8464,N_7065,N_6083);
nor U8465 (N_8465,N_7379,N_6492);
nor U8466 (N_8466,N_7010,N_7091);
nand U8467 (N_8467,N_6019,N_6158);
and U8468 (N_8468,N_6808,N_6830);
and U8469 (N_8469,N_6283,N_6411);
or U8470 (N_8470,N_6871,N_7024);
nand U8471 (N_8471,N_7335,N_7077);
nand U8472 (N_8472,N_7182,N_7104);
xor U8473 (N_8473,N_6802,N_7436);
or U8474 (N_8474,N_6945,N_6124);
nand U8475 (N_8475,N_6604,N_6337);
or U8476 (N_8476,N_6502,N_6969);
or U8477 (N_8477,N_7179,N_6242);
or U8478 (N_8478,N_7154,N_7499);
nor U8479 (N_8479,N_7229,N_6611);
or U8480 (N_8480,N_7372,N_6361);
or U8481 (N_8481,N_7262,N_6576);
or U8482 (N_8482,N_7020,N_7143);
and U8483 (N_8483,N_6883,N_7346);
xnor U8484 (N_8484,N_6638,N_6797);
and U8485 (N_8485,N_7314,N_7091);
nand U8486 (N_8486,N_6342,N_7075);
nor U8487 (N_8487,N_6743,N_7202);
or U8488 (N_8488,N_7400,N_6771);
and U8489 (N_8489,N_6701,N_6259);
nand U8490 (N_8490,N_7462,N_6669);
or U8491 (N_8491,N_6098,N_6719);
nand U8492 (N_8492,N_6597,N_6769);
or U8493 (N_8493,N_6368,N_6249);
nor U8494 (N_8494,N_6925,N_6772);
nand U8495 (N_8495,N_6367,N_7230);
nor U8496 (N_8496,N_7219,N_7345);
nand U8497 (N_8497,N_6591,N_7212);
nand U8498 (N_8498,N_6357,N_7260);
or U8499 (N_8499,N_6322,N_6252);
nand U8500 (N_8500,N_6201,N_6106);
and U8501 (N_8501,N_6977,N_6173);
or U8502 (N_8502,N_6462,N_6366);
and U8503 (N_8503,N_6569,N_7425);
nand U8504 (N_8504,N_7391,N_6662);
xnor U8505 (N_8505,N_6363,N_7032);
or U8506 (N_8506,N_7422,N_7344);
nor U8507 (N_8507,N_7169,N_7019);
nor U8508 (N_8508,N_6988,N_7408);
nor U8509 (N_8509,N_6892,N_6517);
or U8510 (N_8510,N_6234,N_7332);
nor U8511 (N_8511,N_6563,N_6166);
xnor U8512 (N_8512,N_7422,N_6081);
xnor U8513 (N_8513,N_6472,N_6397);
nand U8514 (N_8514,N_6506,N_6498);
or U8515 (N_8515,N_6140,N_6552);
nor U8516 (N_8516,N_7095,N_6597);
or U8517 (N_8517,N_7068,N_7205);
xor U8518 (N_8518,N_7019,N_6904);
or U8519 (N_8519,N_7477,N_7040);
and U8520 (N_8520,N_6002,N_6095);
xnor U8521 (N_8521,N_6229,N_6931);
nor U8522 (N_8522,N_7461,N_6749);
nand U8523 (N_8523,N_6904,N_6155);
or U8524 (N_8524,N_6469,N_7453);
xor U8525 (N_8525,N_6225,N_7234);
and U8526 (N_8526,N_6723,N_7170);
xor U8527 (N_8527,N_6205,N_6732);
nor U8528 (N_8528,N_7456,N_6919);
and U8529 (N_8529,N_6380,N_6771);
and U8530 (N_8530,N_6459,N_7065);
and U8531 (N_8531,N_7295,N_6746);
nor U8532 (N_8532,N_6690,N_6317);
or U8533 (N_8533,N_6470,N_6784);
nor U8534 (N_8534,N_6294,N_6140);
and U8535 (N_8535,N_6960,N_7098);
and U8536 (N_8536,N_6970,N_7203);
and U8537 (N_8537,N_6200,N_6336);
or U8538 (N_8538,N_6257,N_6519);
nand U8539 (N_8539,N_6659,N_6810);
or U8540 (N_8540,N_7030,N_7466);
or U8541 (N_8541,N_7476,N_7364);
nor U8542 (N_8542,N_6110,N_6212);
and U8543 (N_8543,N_6816,N_6635);
or U8544 (N_8544,N_6692,N_6960);
xnor U8545 (N_8545,N_6953,N_6036);
or U8546 (N_8546,N_6357,N_7177);
nor U8547 (N_8547,N_6584,N_7351);
and U8548 (N_8548,N_7290,N_6246);
or U8549 (N_8549,N_6430,N_6568);
nor U8550 (N_8550,N_6522,N_6730);
and U8551 (N_8551,N_6097,N_6877);
or U8552 (N_8552,N_6330,N_6938);
and U8553 (N_8553,N_7208,N_6192);
nand U8554 (N_8554,N_6342,N_6808);
nand U8555 (N_8555,N_7289,N_6108);
or U8556 (N_8556,N_6608,N_6339);
nor U8557 (N_8557,N_7377,N_6413);
or U8558 (N_8558,N_6081,N_6830);
or U8559 (N_8559,N_7104,N_6244);
nand U8560 (N_8560,N_7057,N_7201);
nor U8561 (N_8561,N_7058,N_6264);
nor U8562 (N_8562,N_7445,N_6046);
and U8563 (N_8563,N_6076,N_6763);
and U8564 (N_8564,N_6337,N_7052);
or U8565 (N_8565,N_7264,N_6715);
nand U8566 (N_8566,N_6172,N_6883);
nand U8567 (N_8567,N_6197,N_7315);
nand U8568 (N_8568,N_6447,N_6022);
or U8569 (N_8569,N_7110,N_7493);
nand U8570 (N_8570,N_6573,N_6647);
nand U8571 (N_8571,N_6292,N_7096);
and U8572 (N_8572,N_7454,N_7336);
nor U8573 (N_8573,N_7046,N_6246);
and U8574 (N_8574,N_6296,N_6975);
or U8575 (N_8575,N_7361,N_6431);
or U8576 (N_8576,N_6802,N_6302);
nand U8577 (N_8577,N_7339,N_6923);
nand U8578 (N_8578,N_7226,N_7092);
or U8579 (N_8579,N_7249,N_6161);
or U8580 (N_8580,N_7218,N_6104);
nand U8581 (N_8581,N_7138,N_7047);
or U8582 (N_8582,N_7135,N_7228);
nor U8583 (N_8583,N_6296,N_7340);
or U8584 (N_8584,N_6227,N_6106);
nor U8585 (N_8585,N_6718,N_7243);
nand U8586 (N_8586,N_7380,N_7331);
nand U8587 (N_8587,N_6381,N_7449);
nand U8588 (N_8588,N_6850,N_7058);
or U8589 (N_8589,N_6770,N_6545);
nor U8590 (N_8590,N_6240,N_6822);
or U8591 (N_8591,N_6687,N_6390);
xor U8592 (N_8592,N_7384,N_6327);
and U8593 (N_8593,N_6950,N_6049);
xor U8594 (N_8594,N_7411,N_6718);
or U8595 (N_8595,N_6706,N_6145);
and U8596 (N_8596,N_6341,N_7117);
xnor U8597 (N_8597,N_6395,N_6136);
and U8598 (N_8598,N_6150,N_6204);
nor U8599 (N_8599,N_6457,N_7294);
nor U8600 (N_8600,N_7297,N_7031);
nand U8601 (N_8601,N_6370,N_7496);
and U8602 (N_8602,N_6866,N_6855);
and U8603 (N_8603,N_7189,N_7253);
or U8604 (N_8604,N_6982,N_7358);
or U8605 (N_8605,N_6992,N_6949);
xnor U8606 (N_8606,N_6127,N_7162);
and U8607 (N_8607,N_6452,N_6503);
nor U8608 (N_8608,N_7104,N_7296);
xor U8609 (N_8609,N_6067,N_6919);
nand U8610 (N_8610,N_6437,N_7220);
nor U8611 (N_8611,N_6452,N_7379);
and U8612 (N_8612,N_7010,N_7454);
nor U8613 (N_8613,N_6685,N_6220);
or U8614 (N_8614,N_6337,N_6208);
and U8615 (N_8615,N_7092,N_6651);
nor U8616 (N_8616,N_7315,N_6841);
and U8617 (N_8617,N_6135,N_6201);
nand U8618 (N_8618,N_7131,N_6016);
and U8619 (N_8619,N_6779,N_6349);
nor U8620 (N_8620,N_6330,N_6401);
nor U8621 (N_8621,N_6207,N_6838);
nor U8622 (N_8622,N_6189,N_6113);
nor U8623 (N_8623,N_7226,N_6564);
nor U8624 (N_8624,N_7047,N_6005);
and U8625 (N_8625,N_6910,N_6790);
xor U8626 (N_8626,N_6746,N_7460);
and U8627 (N_8627,N_6470,N_6488);
nand U8628 (N_8628,N_7196,N_6151);
or U8629 (N_8629,N_7273,N_6239);
or U8630 (N_8630,N_6354,N_6682);
nor U8631 (N_8631,N_7340,N_7409);
nor U8632 (N_8632,N_6591,N_6992);
nor U8633 (N_8633,N_6498,N_6755);
and U8634 (N_8634,N_6720,N_6639);
xnor U8635 (N_8635,N_6324,N_6728);
xor U8636 (N_8636,N_6414,N_6111);
and U8637 (N_8637,N_6737,N_6113);
nand U8638 (N_8638,N_7417,N_7341);
and U8639 (N_8639,N_7194,N_6820);
and U8640 (N_8640,N_6594,N_6652);
and U8641 (N_8641,N_7413,N_6930);
or U8642 (N_8642,N_6790,N_7166);
and U8643 (N_8643,N_7370,N_6778);
and U8644 (N_8644,N_7052,N_6987);
nand U8645 (N_8645,N_6073,N_6282);
and U8646 (N_8646,N_7342,N_6058);
and U8647 (N_8647,N_6981,N_6124);
nand U8648 (N_8648,N_7374,N_6639);
nor U8649 (N_8649,N_6201,N_6586);
xor U8650 (N_8650,N_6718,N_7386);
nor U8651 (N_8651,N_6364,N_6585);
or U8652 (N_8652,N_6721,N_7035);
xnor U8653 (N_8653,N_6638,N_6338);
nor U8654 (N_8654,N_7111,N_6426);
or U8655 (N_8655,N_6400,N_7177);
xnor U8656 (N_8656,N_6441,N_7112);
and U8657 (N_8657,N_7116,N_6825);
nor U8658 (N_8658,N_6994,N_7434);
or U8659 (N_8659,N_6169,N_6343);
nand U8660 (N_8660,N_6273,N_6563);
or U8661 (N_8661,N_6642,N_7447);
and U8662 (N_8662,N_7379,N_6412);
nand U8663 (N_8663,N_7085,N_6814);
or U8664 (N_8664,N_7310,N_6463);
nand U8665 (N_8665,N_7086,N_6938);
or U8666 (N_8666,N_6083,N_7105);
nor U8667 (N_8667,N_7443,N_6911);
and U8668 (N_8668,N_6887,N_6828);
or U8669 (N_8669,N_7376,N_7499);
or U8670 (N_8670,N_6912,N_6575);
and U8671 (N_8671,N_6318,N_6802);
nand U8672 (N_8672,N_6666,N_6021);
and U8673 (N_8673,N_6514,N_6597);
and U8674 (N_8674,N_7122,N_6556);
xnor U8675 (N_8675,N_7057,N_7132);
or U8676 (N_8676,N_6046,N_7022);
or U8677 (N_8677,N_6708,N_6250);
xor U8678 (N_8678,N_7321,N_6754);
and U8679 (N_8679,N_6697,N_7194);
nand U8680 (N_8680,N_6645,N_6042);
and U8681 (N_8681,N_6794,N_6159);
and U8682 (N_8682,N_6340,N_7433);
or U8683 (N_8683,N_6152,N_6823);
or U8684 (N_8684,N_6894,N_6153);
and U8685 (N_8685,N_7282,N_6522);
nor U8686 (N_8686,N_6827,N_7408);
nor U8687 (N_8687,N_6466,N_6776);
or U8688 (N_8688,N_6958,N_6268);
and U8689 (N_8689,N_6344,N_6798);
nand U8690 (N_8690,N_7408,N_7228);
nand U8691 (N_8691,N_6183,N_6003);
or U8692 (N_8692,N_6576,N_7022);
nor U8693 (N_8693,N_7002,N_7292);
nand U8694 (N_8694,N_7020,N_7209);
nand U8695 (N_8695,N_7283,N_7285);
nand U8696 (N_8696,N_6568,N_6800);
nor U8697 (N_8697,N_6960,N_7436);
nor U8698 (N_8698,N_6887,N_7467);
nor U8699 (N_8699,N_6142,N_6674);
nor U8700 (N_8700,N_6369,N_7185);
nand U8701 (N_8701,N_6819,N_6341);
or U8702 (N_8702,N_6158,N_6646);
or U8703 (N_8703,N_6900,N_7340);
or U8704 (N_8704,N_6661,N_6879);
nor U8705 (N_8705,N_7396,N_6959);
xor U8706 (N_8706,N_6443,N_7303);
nand U8707 (N_8707,N_6606,N_6482);
nor U8708 (N_8708,N_7153,N_6357);
nand U8709 (N_8709,N_7438,N_7035);
or U8710 (N_8710,N_7282,N_7066);
or U8711 (N_8711,N_7247,N_6683);
or U8712 (N_8712,N_7008,N_7276);
or U8713 (N_8713,N_6486,N_6147);
nor U8714 (N_8714,N_6549,N_7082);
nand U8715 (N_8715,N_6180,N_7147);
and U8716 (N_8716,N_7097,N_6818);
nand U8717 (N_8717,N_6902,N_6435);
nand U8718 (N_8718,N_6760,N_6744);
nor U8719 (N_8719,N_7455,N_6121);
and U8720 (N_8720,N_6844,N_6398);
xnor U8721 (N_8721,N_6824,N_6929);
and U8722 (N_8722,N_6916,N_6264);
nor U8723 (N_8723,N_6031,N_6086);
nand U8724 (N_8724,N_7188,N_6000);
nand U8725 (N_8725,N_7456,N_6435);
or U8726 (N_8726,N_6573,N_6655);
nor U8727 (N_8727,N_6174,N_7018);
nand U8728 (N_8728,N_6098,N_6297);
xor U8729 (N_8729,N_6616,N_6908);
nor U8730 (N_8730,N_7427,N_6604);
and U8731 (N_8731,N_6373,N_6578);
nand U8732 (N_8732,N_6021,N_6744);
xnor U8733 (N_8733,N_7353,N_7403);
and U8734 (N_8734,N_7334,N_6722);
or U8735 (N_8735,N_6035,N_6334);
nor U8736 (N_8736,N_6119,N_7045);
nand U8737 (N_8737,N_6810,N_6774);
xnor U8738 (N_8738,N_7036,N_6465);
nand U8739 (N_8739,N_7179,N_7200);
and U8740 (N_8740,N_6871,N_7321);
nand U8741 (N_8741,N_7426,N_6340);
nand U8742 (N_8742,N_7225,N_6642);
nor U8743 (N_8743,N_6293,N_7460);
xnor U8744 (N_8744,N_7378,N_6709);
and U8745 (N_8745,N_6222,N_7143);
and U8746 (N_8746,N_6895,N_6153);
nand U8747 (N_8747,N_6243,N_6191);
or U8748 (N_8748,N_6955,N_6141);
or U8749 (N_8749,N_7126,N_6009);
nand U8750 (N_8750,N_6007,N_7187);
and U8751 (N_8751,N_7071,N_7442);
or U8752 (N_8752,N_6208,N_7032);
xnor U8753 (N_8753,N_7206,N_6397);
nor U8754 (N_8754,N_7381,N_7075);
xor U8755 (N_8755,N_7160,N_6300);
xnor U8756 (N_8756,N_6650,N_6460);
or U8757 (N_8757,N_6444,N_6121);
nand U8758 (N_8758,N_7377,N_6681);
nand U8759 (N_8759,N_6185,N_6353);
nand U8760 (N_8760,N_6139,N_7037);
or U8761 (N_8761,N_6210,N_6122);
and U8762 (N_8762,N_6632,N_6313);
or U8763 (N_8763,N_6846,N_7068);
and U8764 (N_8764,N_7141,N_7056);
nand U8765 (N_8765,N_6491,N_6757);
or U8766 (N_8766,N_6341,N_6009);
nand U8767 (N_8767,N_6713,N_6541);
nand U8768 (N_8768,N_6867,N_6537);
nand U8769 (N_8769,N_6487,N_7289);
xor U8770 (N_8770,N_6744,N_6935);
nand U8771 (N_8771,N_7192,N_6446);
or U8772 (N_8772,N_7039,N_6189);
nand U8773 (N_8773,N_6779,N_6661);
or U8774 (N_8774,N_6491,N_6658);
and U8775 (N_8775,N_7017,N_6871);
and U8776 (N_8776,N_6148,N_6593);
nor U8777 (N_8777,N_7281,N_6108);
and U8778 (N_8778,N_6897,N_7473);
and U8779 (N_8779,N_6838,N_6210);
nand U8780 (N_8780,N_7377,N_7139);
and U8781 (N_8781,N_7348,N_7173);
or U8782 (N_8782,N_7109,N_7163);
or U8783 (N_8783,N_7284,N_6466);
and U8784 (N_8784,N_6394,N_6061);
nor U8785 (N_8785,N_6739,N_7381);
and U8786 (N_8786,N_6589,N_6456);
xnor U8787 (N_8787,N_6335,N_7377);
or U8788 (N_8788,N_6371,N_7277);
and U8789 (N_8789,N_6359,N_6213);
nand U8790 (N_8790,N_6309,N_6876);
nor U8791 (N_8791,N_6423,N_6292);
nand U8792 (N_8792,N_6926,N_6668);
nor U8793 (N_8793,N_6455,N_6961);
nor U8794 (N_8794,N_6705,N_6674);
xnor U8795 (N_8795,N_6445,N_6109);
or U8796 (N_8796,N_6109,N_7000);
or U8797 (N_8797,N_6602,N_6277);
nor U8798 (N_8798,N_6541,N_7116);
nor U8799 (N_8799,N_6752,N_7171);
and U8800 (N_8800,N_7094,N_6195);
nor U8801 (N_8801,N_6960,N_7111);
and U8802 (N_8802,N_7012,N_7021);
nor U8803 (N_8803,N_7448,N_6487);
nor U8804 (N_8804,N_7041,N_6531);
nor U8805 (N_8805,N_6002,N_6818);
nand U8806 (N_8806,N_6717,N_7363);
nor U8807 (N_8807,N_6992,N_6315);
nor U8808 (N_8808,N_7408,N_6992);
nor U8809 (N_8809,N_6263,N_6892);
xor U8810 (N_8810,N_6745,N_6309);
and U8811 (N_8811,N_7234,N_6858);
nand U8812 (N_8812,N_7191,N_7463);
or U8813 (N_8813,N_6973,N_6691);
or U8814 (N_8814,N_6354,N_6752);
nor U8815 (N_8815,N_6834,N_6697);
nor U8816 (N_8816,N_7080,N_7293);
or U8817 (N_8817,N_6250,N_7189);
nor U8818 (N_8818,N_7443,N_6088);
nand U8819 (N_8819,N_6666,N_6002);
and U8820 (N_8820,N_6813,N_7245);
or U8821 (N_8821,N_6523,N_6010);
and U8822 (N_8822,N_6291,N_7353);
and U8823 (N_8823,N_7408,N_7229);
nand U8824 (N_8824,N_7197,N_6406);
xnor U8825 (N_8825,N_6158,N_6041);
or U8826 (N_8826,N_7278,N_6924);
or U8827 (N_8827,N_6509,N_6612);
nand U8828 (N_8828,N_6310,N_7263);
or U8829 (N_8829,N_7213,N_6596);
or U8830 (N_8830,N_6355,N_7325);
or U8831 (N_8831,N_6699,N_6013);
and U8832 (N_8832,N_6900,N_7366);
nand U8833 (N_8833,N_6631,N_6550);
nor U8834 (N_8834,N_6840,N_6680);
nor U8835 (N_8835,N_6464,N_7404);
or U8836 (N_8836,N_6226,N_7365);
and U8837 (N_8837,N_6841,N_6468);
xor U8838 (N_8838,N_7074,N_7382);
nand U8839 (N_8839,N_6887,N_6755);
or U8840 (N_8840,N_6630,N_6029);
xnor U8841 (N_8841,N_6968,N_7248);
and U8842 (N_8842,N_6296,N_7317);
or U8843 (N_8843,N_6074,N_6494);
and U8844 (N_8844,N_7285,N_6426);
nand U8845 (N_8845,N_6939,N_6443);
nor U8846 (N_8846,N_7212,N_6744);
xor U8847 (N_8847,N_6297,N_7223);
and U8848 (N_8848,N_6051,N_6582);
or U8849 (N_8849,N_6965,N_6768);
or U8850 (N_8850,N_6511,N_6348);
xor U8851 (N_8851,N_7234,N_6864);
nand U8852 (N_8852,N_6248,N_6915);
nor U8853 (N_8853,N_6270,N_6716);
and U8854 (N_8854,N_6461,N_7151);
and U8855 (N_8855,N_7159,N_6529);
nand U8856 (N_8856,N_7358,N_6496);
or U8857 (N_8857,N_6900,N_6825);
nor U8858 (N_8858,N_6884,N_6984);
or U8859 (N_8859,N_7435,N_6177);
nor U8860 (N_8860,N_6280,N_6133);
nand U8861 (N_8861,N_6465,N_6130);
and U8862 (N_8862,N_6611,N_6402);
nand U8863 (N_8863,N_7298,N_6591);
nor U8864 (N_8864,N_7258,N_6989);
nor U8865 (N_8865,N_7447,N_6921);
nand U8866 (N_8866,N_6034,N_6483);
nand U8867 (N_8867,N_6213,N_6304);
nor U8868 (N_8868,N_6000,N_6776);
nand U8869 (N_8869,N_7417,N_7303);
nor U8870 (N_8870,N_6689,N_6345);
and U8871 (N_8871,N_6321,N_6162);
nand U8872 (N_8872,N_6578,N_7087);
nor U8873 (N_8873,N_6643,N_6762);
nand U8874 (N_8874,N_6492,N_6178);
and U8875 (N_8875,N_7245,N_7430);
and U8876 (N_8876,N_6829,N_6478);
and U8877 (N_8877,N_6495,N_6564);
and U8878 (N_8878,N_7206,N_6839);
or U8879 (N_8879,N_6037,N_7347);
nor U8880 (N_8880,N_7147,N_6808);
xnor U8881 (N_8881,N_6801,N_6007);
and U8882 (N_8882,N_6282,N_6216);
nor U8883 (N_8883,N_6963,N_6909);
nor U8884 (N_8884,N_7465,N_6732);
and U8885 (N_8885,N_7054,N_6267);
or U8886 (N_8886,N_6422,N_6830);
or U8887 (N_8887,N_6995,N_7262);
and U8888 (N_8888,N_6525,N_6011);
and U8889 (N_8889,N_6329,N_6937);
or U8890 (N_8890,N_6942,N_7078);
nand U8891 (N_8891,N_7461,N_6199);
nand U8892 (N_8892,N_6631,N_6962);
or U8893 (N_8893,N_7379,N_7028);
nand U8894 (N_8894,N_6362,N_6591);
and U8895 (N_8895,N_6503,N_7455);
nand U8896 (N_8896,N_6026,N_6189);
nand U8897 (N_8897,N_6105,N_7437);
or U8898 (N_8898,N_6164,N_6693);
nor U8899 (N_8899,N_7313,N_6084);
nor U8900 (N_8900,N_6496,N_6137);
nand U8901 (N_8901,N_7031,N_7127);
or U8902 (N_8902,N_6532,N_6608);
or U8903 (N_8903,N_7353,N_6982);
or U8904 (N_8904,N_7211,N_7034);
nor U8905 (N_8905,N_7139,N_7068);
nor U8906 (N_8906,N_6248,N_7118);
or U8907 (N_8907,N_6604,N_6450);
and U8908 (N_8908,N_6417,N_6815);
and U8909 (N_8909,N_6275,N_6492);
nor U8910 (N_8910,N_6285,N_6159);
xor U8911 (N_8911,N_7217,N_7072);
xor U8912 (N_8912,N_6678,N_6668);
xor U8913 (N_8913,N_6872,N_6194);
nor U8914 (N_8914,N_6071,N_6694);
and U8915 (N_8915,N_7432,N_7484);
nand U8916 (N_8916,N_7180,N_6480);
nor U8917 (N_8917,N_6435,N_6397);
and U8918 (N_8918,N_6928,N_6909);
or U8919 (N_8919,N_7144,N_6950);
xnor U8920 (N_8920,N_6507,N_6776);
nor U8921 (N_8921,N_7257,N_7405);
nand U8922 (N_8922,N_6186,N_6003);
nor U8923 (N_8923,N_6231,N_7391);
and U8924 (N_8924,N_7217,N_6768);
nand U8925 (N_8925,N_7062,N_6623);
xor U8926 (N_8926,N_6723,N_6546);
and U8927 (N_8927,N_7381,N_6645);
nor U8928 (N_8928,N_6589,N_6147);
or U8929 (N_8929,N_7443,N_7454);
or U8930 (N_8930,N_6908,N_7170);
nor U8931 (N_8931,N_6027,N_7278);
or U8932 (N_8932,N_6878,N_6620);
nor U8933 (N_8933,N_7346,N_6823);
or U8934 (N_8934,N_6966,N_6515);
or U8935 (N_8935,N_6709,N_6907);
nor U8936 (N_8936,N_6733,N_6312);
nor U8937 (N_8937,N_6668,N_6020);
or U8938 (N_8938,N_6108,N_6142);
and U8939 (N_8939,N_6627,N_7441);
nor U8940 (N_8940,N_7136,N_7399);
or U8941 (N_8941,N_6900,N_6787);
and U8942 (N_8942,N_6760,N_6968);
or U8943 (N_8943,N_6404,N_7135);
and U8944 (N_8944,N_6291,N_7307);
and U8945 (N_8945,N_6537,N_7075);
and U8946 (N_8946,N_6200,N_6114);
and U8947 (N_8947,N_7225,N_7250);
or U8948 (N_8948,N_7078,N_6891);
nand U8949 (N_8949,N_6027,N_6716);
and U8950 (N_8950,N_7283,N_6514);
and U8951 (N_8951,N_7060,N_6142);
and U8952 (N_8952,N_7231,N_6469);
nand U8953 (N_8953,N_6563,N_6417);
or U8954 (N_8954,N_6993,N_7238);
or U8955 (N_8955,N_6295,N_6961);
nor U8956 (N_8956,N_7465,N_7233);
nor U8957 (N_8957,N_7305,N_6298);
xnor U8958 (N_8958,N_6242,N_6918);
or U8959 (N_8959,N_6507,N_6718);
xnor U8960 (N_8960,N_6309,N_7299);
nand U8961 (N_8961,N_6387,N_6931);
or U8962 (N_8962,N_6740,N_7499);
and U8963 (N_8963,N_7047,N_6024);
nand U8964 (N_8964,N_6054,N_7124);
nor U8965 (N_8965,N_6396,N_6613);
nand U8966 (N_8966,N_7360,N_6671);
nor U8967 (N_8967,N_7493,N_6375);
nor U8968 (N_8968,N_6215,N_7239);
and U8969 (N_8969,N_6453,N_7498);
or U8970 (N_8970,N_6100,N_6204);
and U8971 (N_8971,N_6116,N_7396);
nand U8972 (N_8972,N_6202,N_6281);
nand U8973 (N_8973,N_6981,N_6510);
nand U8974 (N_8974,N_7316,N_6376);
nor U8975 (N_8975,N_6516,N_6221);
or U8976 (N_8976,N_6426,N_6626);
nand U8977 (N_8977,N_6173,N_6712);
nand U8978 (N_8978,N_6519,N_6929);
nand U8979 (N_8979,N_7349,N_7006);
nand U8980 (N_8980,N_6347,N_6525);
nor U8981 (N_8981,N_6748,N_6399);
or U8982 (N_8982,N_6038,N_6840);
xor U8983 (N_8983,N_6312,N_7462);
nor U8984 (N_8984,N_6654,N_6053);
or U8985 (N_8985,N_6827,N_7208);
and U8986 (N_8986,N_6117,N_6705);
or U8987 (N_8987,N_6869,N_6461);
nand U8988 (N_8988,N_6909,N_7332);
nor U8989 (N_8989,N_6393,N_7043);
nor U8990 (N_8990,N_6433,N_6682);
or U8991 (N_8991,N_6562,N_6195);
xor U8992 (N_8992,N_6840,N_7303);
nand U8993 (N_8993,N_6058,N_6679);
nand U8994 (N_8994,N_6609,N_6607);
nor U8995 (N_8995,N_6935,N_6031);
nand U8996 (N_8996,N_6306,N_7214);
nand U8997 (N_8997,N_6883,N_7295);
nand U8998 (N_8998,N_6351,N_6878);
and U8999 (N_8999,N_6615,N_6391);
or U9000 (N_9000,N_8816,N_7611);
and U9001 (N_9001,N_7770,N_8498);
or U9002 (N_9002,N_8933,N_7805);
or U9003 (N_9003,N_8096,N_8900);
nand U9004 (N_9004,N_7606,N_8731);
or U9005 (N_9005,N_7901,N_8046);
and U9006 (N_9006,N_8334,N_7858);
or U9007 (N_9007,N_8296,N_7904);
nor U9008 (N_9008,N_8438,N_8412);
nor U9009 (N_9009,N_7616,N_8315);
or U9010 (N_9010,N_7953,N_8607);
or U9011 (N_9011,N_7669,N_7703);
nand U9012 (N_9012,N_8828,N_7954);
nand U9013 (N_9013,N_8026,N_7879);
and U9014 (N_9014,N_8734,N_7543);
or U9015 (N_9015,N_8467,N_7614);
nor U9016 (N_9016,N_7756,N_7689);
or U9017 (N_9017,N_8157,N_7682);
and U9018 (N_9018,N_8718,N_8437);
or U9019 (N_9019,N_7965,N_7629);
nand U9020 (N_9020,N_8529,N_7857);
nor U9021 (N_9021,N_7664,N_7736);
nand U9022 (N_9022,N_8672,N_8358);
and U9023 (N_9023,N_7711,N_8683);
and U9024 (N_9024,N_8175,N_7655);
nand U9025 (N_9025,N_7557,N_8912);
nor U9026 (N_9026,N_8509,N_8924);
and U9027 (N_9027,N_8201,N_8658);
nor U9028 (N_9028,N_7727,N_8777);
or U9029 (N_9029,N_8899,N_8324);
nand U9030 (N_9030,N_8551,N_8294);
nand U9031 (N_9031,N_8176,N_8878);
nor U9032 (N_9032,N_8156,N_8927);
and U9033 (N_9033,N_8775,N_7880);
and U9034 (N_9034,N_8633,N_8081);
nand U9035 (N_9035,N_7994,N_8302);
and U9036 (N_9036,N_7725,N_8946);
or U9037 (N_9037,N_8055,N_7995);
and U9038 (N_9038,N_7673,N_8231);
nor U9039 (N_9039,N_8392,N_7983);
or U9040 (N_9040,N_8763,N_8812);
or U9041 (N_9041,N_8552,N_8217);
or U9042 (N_9042,N_8240,N_8316);
nor U9043 (N_9043,N_8182,N_8928);
or U9044 (N_9044,N_8239,N_8515);
or U9045 (N_9045,N_8979,N_8123);
nand U9046 (N_9046,N_7838,N_7530);
xnor U9047 (N_9047,N_8838,N_8139);
nor U9048 (N_9048,N_7848,N_8114);
or U9049 (N_9049,N_7704,N_8428);
nand U9050 (N_9050,N_8003,N_8132);
nor U9051 (N_9051,N_7870,N_8257);
nand U9052 (N_9052,N_7944,N_8192);
or U9053 (N_9053,N_8715,N_8908);
nor U9054 (N_9054,N_8312,N_7849);
nand U9055 (N_9055,N_8477,N_8459);
xnor U9056 (N_9056,N_8343,N_7729);
and U9057 (N_9057,N_8999,N_8195);
nor U9058 (N_9058,N_8407,N_8864);
and U9059 (N_9059,N_7815,N_8295);
nand U9060 (N_9060,N_8987,N_8199);
xnor U9061 (N_9061,N_7897,N_7713);
nor U9062 (N_9062,N_7856,N_8062);
nor U9063 (N_9063,N_8090,N_8546);
and U9064 (N_9064,N_8751,N_8948);
or U9065 (N_9065,N_8663,N_7911);
nor U9066 (N_9066,N_7651,N_8406);
and U9067 (N_9067,N_7505,N_8506);
or U9068 (N_9068,N_7973,N_8242);
and U9069 (N_9069,N_8189,N_7896);
or U9070 (N_9070,N_7720,N_8198);
and U9071 (N_9071,N_8920,N_7674);
nand U9072 (N_9072,N_8208,N_7641);
xnor U9073 (N_9073,N_8889,N_8961);
or U9074 (N_9074,N_8616,N_8004);
nand U9075 (N_9075,N_8502,N_8023);
or U9076 (N_9076,N_8747,N_8468);
nand U9077 (N_9077,N_8105,N_8807);
and U9078 (N_9078,N_8103,N_7663);
nor U9079 (N_9079,N_8101,N_8339);
nor U9080 (N_9080,N_7974,N_8771);
and U9081 (N_9081,N_7508,N_8568);
or U9082 (N_9082,N_8749,N_8142);
and U9083 (N_9083,N_8014,N_8153);
or U9084 (N_9084,N_8443,N_8656);
or U9085 (N_9085,N_7997,N_8687);
nor U9086 (N_9086,N_8094,N_8365);
and U9087 (N_9087,N_7722,N_8678);
nand U9088 (N_9088,N_7827,N_8440);
nand U9089 (N_9089,N_8093,N_7752);
nor U9090 (N_9090,N_7726,N_8901);
nor U9091 (N_9091,N_7889,N_7649);
or U9092 (N_9092,N_8832,N_8915);
and U9093 (N_9093,N_8660,N_8914);
and U9094 (N_9094,N_8880,N_7812);
nand U9095 (N_9095,N_8333,N_8635);
nand U9096 (N_9096,N_7886,N_7922);
nand U9097 (N_9097,N_8845,N_7573);
and U9098 (N_9098,N_8364,N_7613);
nor U9099 (N_9099,N_8919,N_8609);
or U9100 (N_9100,N_8562,N_8266);
xnor U9101 (N_9101,N_8359,N_7843);
nor U9102 (N_9102,N_8868,N_8320);
and U9103 (N_9103,N_7580,N_8967);
and U9104 (N_9104,N_8367,N_8408);
or U9105 (N_9105,N_7630,N_7788);
or U9106 (N_9106,N_8022,N_7619);
nor U9107 (N_9107,N_7891,N_7855);
or U9108 (N_9108,N_8808,N_8642);
and U9109 (N_9109,N_8177,N_8457);
nor U9110 (N_9110,N_7554,N_7877);
or U9111 (N_9111,N_8196,N_8416);
or U9112 (N_9112,N_8647,N_8215);
and U9113 (N_9113,N_8471,N_7626);
nand U9114 (N_9114,N_8073,N_8719);
xor U9115 (N_9115,N_8473,N_8701);
nand U9116 (N_9116,N_7688,N_8779);
and U9117 (N_9117,N_8492,N_8826);
nor U9118 (N_9118,N_7793,N_8284);
or U9119 (N_9119,N_8051,N_7768);
and U9120 (N_9120,N_8482,N_7790);
nor U9121 (N_9121,N_7942,N_8265);
and U9122 (N_9122,N_8465,N_7938);
nand U9123 (N_9123,N_7662,N_8422);
nand U9124 (N_9124,N_7832,N_8038);
nand U9125 (N_9125,N_8382,N_8882);
or U9126 (N_9126,N_8223,N_8335);
or U9127 (N_9127,N_7550,N_8847);
nand U9128 (N_9128,N_8301,N_8236);
nand U9129 (N_9129,N_8614,N_8224);
nand U9130 (N_9130,N_8227,N_8735);
nor U9131 (N_9131,N_7975,N_7825);
nor U9132 (N_9132,N_8789,N_8013);
nand U9133 (N_9133,N_8544,N_8274);
and U9134 (N_9134,N_7590,N_7724);
and U9135 (N_9135,N_8824,N_8171);
nor U9136 (N_9136,N_7615,N_7648);
xor U9137 (N_9137,N_7912,N_8653);
nand U9138 (N_9138,N_7513,N_8446);
xnor U9139 (N_9139,N_8149,N_8572);
nand U9140 (N_9140,N_8563,N_8361);
nand U9141 (N_9141,N_7928,N_8929);
or U9142 (N_9142,N_8084,N_8557);
or U9143 (N_9143,N_7739,N_8478);
xor U9144 (N_9144,N_8819,N_8263);
and U9145 (N_9145,N_7665,N_7956);
or U9146 (N_9146,N_8800,N_8330);
or U9147 (N_9147,N_8430,N_8110);
nor U9148 (N_9148,N_8728,N_7656);
nand U9149 (N_9149,N_8996,N_8982);
nor U9150 (N_9150,N_7562,N_7581);
nor U9151 (N_9151,N_8876,N_8232);
nand U9152 (N_9152,N_8148,N_8435);
and U9153 (N_9153,N_8601,N_8993);
and U9154 (N_9154,N_8526,N_7525);
nor U9155 (N_9155,N_8372,N_8949);
and U9156 (N_9156,N_8721,N_7887);
xnor U9157 (N_9157,N_7851,N_7524);
nand U9158 (N_9158,N_8292,N_8336);
and U9159 (N_9159,N_8785,N_8293);
or U9160 (N_9160,N_8268,N_8469);
nand U9161 (N_9161,N_7538,N_7868);
or U9162 (N_9162,N_8277,N_7698);
nand U9163 (N_9163,N_7966,N_7892);
xnor U9164 (N_9164,N_8858,N_7534);
nor U9165 (N_9165,N_7706,N_7523);
or U9166 (N_9166,N_8540,N_8490);
xnor U9167 (N_9167,N_7671,N_7708);
and U9168 (N_9168,N_8803,N_8956);
nand U9169 (N_9169,N_8822,N_7740);
or U9170 (N_9170,N_8748,N_8470);
nor U9171 (N_9171,N_8012,N_8424);
nor U9172 (N_9172,N_8829,N_8100);
and U9173 (N_9173,N_8381,N_7795);
nand U9174 (N_9174,N_8671,N_8860);
and U9175 (N_9175,N_7542,N_7936);
nor U9176 (N_9176,N_8611,N_8973);
xor U9177 (N_9177,N_8898,N_7946);
nand U9178 (N_9178,N_8054,N_8072);
xnor U9179 (N_9179,N_7916,N_7559);
or U9180 (N_9180,N_8584,N_7783);
nand U9181 (N_9181,N_7863,N_8684);
xnor U9182 (N_9182,N_8798,N_8442);
or U9183 (N_9183,N_8821,N_8953);
and U9184 (N_9184,N_7748,N_8995);
or U9185 (N_9185,N_8892,N_8906);
nand U9186 (N_9186,N_8200,N_7835);
nand U9187 (N_9187,N_8657,N_8629);
xnor U9188 (N_9188,N_7607,N_8709);
nand U9189 (N_9189,N_8244,N_8386);
or U9190 (N_9190,N_8089,N_8079);
xnor U9191 (N_9191,N_8885,N_7890);
xor U9192 (N_9192,N_8505,N_7931);
nand U9193 (N_9193,N_8074,N_7785);
nor U9194 (N_9194,N_8087,N_8311);
and U9195 (N_9195,N_8269,N_8379);
nor U9196 (N_9196,N_8698,N_8427);
and U9197 (N_9197,N_7751,N_8141);
and U9198 (N_9198,N_8532,N_7798);
nor U9199 (N_9199,N_7802,N_8045);
nand U9200 (N_9200,N_8686,N_7572);
xor U9201 (N_9201,N_8517,N_7810);
nand U9202 (N_9202,N_8321,N_8793);
and U9203 (N_9203,N_8212,N_8297);
or U9204 (N_9204,N_7833,N_8971);
nor U9205 (N_9205,N_8765,N_7503);
nand U9206 (N_9206,N_8666,N_8143);
nor U9207 (N_9207,N_8733,N_8969);
nor U9208 (N_9208,N_8802,N_7899);
nand U9209 (N_9209,N_8581,N_7757);
nor U9210 (N_9210,N_8165,N_8398);
or U9211 (N_9211,N_8275,N_8636);
or U9212 (N_9212,N_8724,N_8495);
nand U9213 (N_9213,N_8942,N_7707);
or U9214 (N_9214,N_8817,N_8944);
xor U9215 (N_9215,N_7509,N_8740);
xor U9216 (N_9216,N_7624,N_7691);
nor U9217 (N_9217,N_7558,N_7749);
and U9218 (N_9218,N_8456,N_7551);
and U9219 (N_9219,N_8389,N_8272);
or U9220 (N_9220,N_8039,N_8503);
nor U9221 (N_9221,N_7579,N_8550);
and U9222 (N_9222,N_7881,N_7610);
nand U9223 (N_9223,N_8426,N_8126);
nor U9224 (N_9224,N_8871,N_7950);
nor U9225 (N_9225,N_7668,N_8623);
nor U9226 (N_9226,N_8064,N_8606);
and U9227 (N_9227,N_7737,N_8936);
nand U9228 (N_9228,N_8814,N_8097);
or U9229 (N_9229,N_8910,N_8075);
nand U9230 (N_9230,N_8166,N_8308);
nor U9231 (N_9231,N_8590,N_7556);
nand U9232 (N_9232,N_8851,N_8583);
nor U9233 (N_9233,N_8145,N_8564);
and U9234 (N_9234,N_8566,N_8388);
nand U9235 (N_9235,N_8491,N_8325);
xnor U9236 (N_9236,N_8884,N_8019);
or U9237 (N_9237,N_8151,N_8638);
and U9238 (N_9238,N_8863,N_7937);
and U9239 (N_9239,N_8521,N_8360);
or U9240 (N_9240,N_8342,N_8797);
and U9241 (N_9241,N_7709,N_7955);
and U9242 (N_9242,N_8685,N_7700);
nor U9243 (N_9243,N_7638,N_8511);
nand U9244 (N_9244,N_7634,N_8837);
nand U9245 (N_9245,N_7609,N_8256);
nor U9246 (N_9246,N_8820,N_7758);
nor U9247 (N_9247,N_7791,N_7745);
nor U9248 (N_9248,N_8744,N_8366);
or U9249 (N_9249,N_8131,N_7660);
nand U9250 (N_9250,N_7893,N_7658);
or U9251 (N_9251,N_8739,N_7985);
or U9252 (N_9252,N_8181,N_7970);
and U9253 (N_9253,N_8397,N_8830);
and U9254 (N_9254,N_8643,N_7667);
nor U9255 (N_9255,N_7883,N_8780);
nor U9256 (N_9256,N_7731,N_7741);
nor U9257 (N_9257,N_8329,N_7536);
xnor U9258 (N_9258,N_8825,N_8138);
or U9259 (N_9259,N_8649,N_8447);
nand U9260 (N_9260,N_8596,N_8624);
nor U9261 (N_9261,N_8534,N_8692);
nor U9262 (N_9262,N_8547,N_8732);
nand U9263 (N_9263,N_8385,N_8931);
and U9264 (N_9264,N_8394,N_8909);
nand U9265 (N_9265,N_8271,N_8720);
nor U9266 (N_9266,N_7876,N_8781);
and U9267 (N_9267,N_7566,N_8690);
or U9268 (N_9268,N_7774,N_7586);
nand U9269 (N_9269,N_7993,N_8625);
nand U9270 (N_9270,N_8917,N_8449);
and U9271 (N_9271,N_8696,N_8567);
xor U9272 (N_9272,N_8620,N_8813);
nor U9273 (N_9273,N_7823,N_8980);
xnor U9274 (N_9274,N_8648,N_7939);
nor U9275 (N_9275,N_8483,N_7560);
and U9276 (N_9276,N_8486,N_7569);
nor U9277 (N_9277,N_7697,N_8621);
nor U9278 (N_9278,N_8879,N_8702);
nor U9279 (N_9279,N_7921,N_7981);
or U9280 (N_9280,N_8834,N_8537);
or U9281 (N_9281,N_8608,N_7753);
or U9282 (N_9282,N_8553,N_8006);
and U9283 (N_9283,N_8270,N_8527);
xnor U9284 (N_9284,N_7618,N_8957);
or U9285 (N_9285,N_7786,N_8988);
or U9286 (N_9286,N_8368,N_8627);
nand U9287 (N_9287,N_8766,N_8036);
or U9288 (N_9288,N_8031,N_7661);
nand U9289 (N_9289,N_8091,N_8178);
nand U9290 (N_9290,N_8764,N_8076);
or U9291 (N_9291,N_8060,N_8183);
nand U9292 (N_9292,N_7597,N_7695);
nor U9293 (N_9293,N_7617,N_8536);
or U9294 (N_9294,N_8887,N_7959);
and U9295 (N_9295,N_8501,N_8654);
or U9296 (N_9296,N_7602,N_8591);
or U9297 (N_9297,N_8512,N_8711);
or U9298 (N_9298,N_7522,N_7742);
or U9299 (N_9299,N_8080,N_7504);
nor U9300 (N_9300,N_8314,N_8356);
nor U9301 (N_9301,N_8147,N_8282);
nor U9302 (N_9302,N_8082,N_8938);
nand U9303 (N_9303,N_7719,N_8016);
nand U9304 (N_9304,N_8790,N_7799);
and U9305 (N_9305,N_8523,N_8574);
or U9306 (N_9306,N_8795,N_8518);
and U9307 (N_9307,N_8053,N_7867);
and U9308 (N_9308,N_7565,N_7564);
xor U9309 (N_9309,N_8264,N_7779);
and U9310 (N_9310,N_8307,N_8363);
or U9311 (N_9311,N_8890,N_8811);
nor U9312 (N_9312,N_8716,N_8921);
nor U9313 (N_9313,N_8859,N_8250);
nor U9314 (N_9314,N_8576,N_8283);
nand U9315 (N_9315,N_7642,N_8886);
nand U9316 (N_9316,N_7919,N_8083);
xnor U9317 (N_9317,N_8228,N_7782);
or U9318 (N_9318,N_8150,N_8078);
and U9319 (N_9319,N_8216,N_8436);
nor U9320 (N_9320,N_8810,N_8682);
xnor U9321 (N_9321,N_7781,N_8209);
nor U9322 (N_9322,N_7888,N_8894);
nor U9323 (N_9323,N_8262,N_8380);
nand U9324 (N_9324,N_8488,N_7920);
and U9325 (N_9325,N_7771,N_7678);
or U9326 (N_9326,N_8603,N_8659);
or U9327 (N_9327,N_8345,N_7780);
nand U9328 (N_9328,N_7644,N_8565);
and U9329 (N_9329,N_8255,N_8298);
xnor U9330 (N_9330,N_8299,N_8514);
nand U9331 (N_9331,N_8410,N_7958);
xor U9332 (N_9332,N_7807,N_8222);
and U9333 (N_9333,N_8856,N_7968);
nand U9334 (N_9334,N_8180,N_7519);
nor U9335 (N_9335,N_8778,N_8758);
nand U9336 (N_9336,N_8130,N_8044);
or U9337 (N_9337,N_7643,N_8007);
and U9338 (N_9338,N_8990,N_8855);
nand U9339 (N_9339,N_8761,N_7675);
nand U9340 (N_9340,N_7913,N_8997);
nor U9341 (N_9341,N_7754,N_8185);
and U9342 (N_9342,N_7631,N_8742);
and U9343 (N_9343,N_8129,N_8652);
or U9344 (N_9344,N_7940,N_8005);
nand U9345 (N_9345,N_8186,N_7670);
or U9346 (N_9346,N_8695,N_8754);
xor U9347 (N_9347,N_8598,N_7633);
or U9348 (N_9348,N_8383,N_8137);
and U9349 (N_9349,N_8613,N_8937);
or U9350 (N_9350,N_7702,N_8873);
nand U9351 (N_9351,N_8461,N_7862);
and U9352 (N_9352,N_8122,N_8500);
and U9353 (N_9353,N_7765,N_8531);
nor U9354 (N_9354,N_7518,N_8809);
xor U9355 (N_9355,N_8421,N_7932);
nand U9356 (N_9356,N_8767,N_8088);
or U9357 (N_9357,N_7875,N_8403);
nor U9358 (N_9358,N_8539,N_8787);
nand U9359 (N_9359,N_8786,N_7577);
and U9360 (N_9360,N_7585,N_8869);
or U9361 (N_9361,N_7517,N_8705);
or U9362 (N_9362,N_7900,N_8370);
or U9363 (N_9363,N_8011,N_8628);
or U9364 (N_9364,N_8475,N_8164);
and U9365 (N_9365,N_8230,N_7694);
nand U9366 (N_9366,N_8943,N_8225);
or U9367 (N_9367,N_7860,N_8922);
and U9368 (N_9368,N_8689,N_8445);
nand U9369 (N_9369,N_7532,N_8327);
and U9370 (N_9370,N_8400,N_8877);
or U9371 (N_9371,N_8507,N_8736);
or U9372 (N_9372,N_8881,N_8688);
nor U9373 (N_9373,N_7687,N_8840);
nand U9374 (N_9374,N_8234,N_8415);
and U9375 (N_9375,N_8211,N_7728);
xor U9376 (N_9376,N_8725,N_7787);
or U9377 (N_9377,N_8681,N_7846);
and U9378 (N_9378,N_8450,N_7679);
and U9379 (N_9379,N_7845,N_8926);
nand U9380 (N_9380,N_8480,N_8753);
nand U9381 (N_9381,N_7917,N_7604);
xnor U9382 (N_9382,N_7811,N_8612);
nand U9383 (N_9383,N_8099,N_8499);
or U9384 (N_9384,N_7962,N_8025);
nand U9385 (N_9385,N_7555,N_8896);
nand U9386 (N_9386,N_8977,N_8190);
nand U9387 (N_9387,N_8116,N_8313);
nand U9388 (N_9388,N_8947,N_8441);
xnor U9389 (N_9389,N_8173,N_7501);
or U9390 (N_9390,N_8543,N_7574);
nand U9391 (N_9391,N_7646,N_8641);
xnor U9392 (N_9392,N_7526,N_8246);
nand U9393 (N_9393,N_8463,N_8548);
nor U9394 (N_9394,N_8842,N_8554);
nand U9395 (N_9395,N_7990,N_8911);
and U9396 (N_9396,N_8951,N_8714);
nor U9397 (N_9397,N_8384,N_8113);
nor U9398 (N_9398,N_8849,N_8570);
or U9399 (N_9399,N_7537,N_7767);
nor U9400 (N_9400,N_8163,N_8419);
nand U9401 (N_9401,N_8640,N_8118);
and U9402 (N_9402,N_8516,N_8791);
or U9403 (N_9403,N_7878,N_8423);
nor U9404 (N_9404,N_8462,N_7608);
nor U9405 (N_9405,N_8144,N_8675);
and U9406 (N_9406,N_7699,N_7963);
and U9407 (N_9407,N_8644,N_7822);
nand U9408 (N_9408,N_8350,N_8960);
xnor U9409 (N_9409,N_8852,N_7831);
nor U9410 (N_9410,N_8989,N_7945);
nand U9411 (N_9411,N_8452,N_7601);
xnor U9412 (N_9412,N_8699,N_7763);
nand U9413 (N_9413,N_7563,N_8226);
and U9414 (N_9414,N_8835,N_8895);
nand U9415 (N_9415,N_7969,N_8586);
and U9416 (N_9416,N_8903,N_8804);
xnor U9417 (N_9417,N_8008,N_7659);
nand U9418 (N_9418,N_8362,N_8579);
nor U9419 (N_9419,N_8261,N_7844);
nor U9420 (N_9420,N_8288,N_7808);
and U9421 (N_9421,N_8393,N_7850);
nand U9422 (N_9422,N_8160,N_8972);
or U9423 (N_9423,N_8095,N_7588);
and U9424 (N_9424,N_8794,N_8872);
and U9425 (N_9425,N_8349,N_7949);
nor U9426 (N_9426,N_7578,N_8976);
nor U9427 (N_9427,N_7693,N_8155);
xor U9428 (N_9428,N_7636,N_7571);
or U9429 (N_9429,N_8328,N_8941);
and U9430 (N_9430,N_8245,N_7506);
nand U9431 (N_9431,N_7803,N_8770);
nor U9432 (N_9432,N_8745,N_8267);
and U9433 (N_9433,N_8970,N_8237);
or U9434 (N_9434,N_7847,N_8479);
nand U9435 (N_9435,N_7764,N_7773);
nor U9436 (N_9436,N_8276,N_8152);
nor U9437 (N_9437,N_8218,N_8755);
or U9438 (N_9438,N_7898,N_8454);
and U9439 (N_9439,N_7853,N_7800);
and U9440 (N_9440,N_7914,N_7977);
or U9441 (N_9441,N_7951,N_8853);
nand U9442 (N_9442,N_8622,N_7620);
nand U9443 (N_9443,N_7511,N_8700);
or U9444 (N_9444,N_8994,N_8319);
nor U9445 (N_9445,N_7657,N_7929);
nor U9446 (N_9446,N_8975,N_8792);
or U9447 (N_9447,N_8214,N_7701);
or U9448 (N_9448,N_8619,N_8846);
or U9449 (N_9449,N_8009,N_7941);
xor U9450 (N_9450,N_7869,N_8634);
nor U9451 (N_9451,N_8252,N_7818);
or U9452 (N_9452,N_8374,N_8027);
or U9453 (N_9453,N_8525,N_8741);
nor U9454 (N_9454,N_8844,N_8371);
nor U9455 (N_9455,N_7794,N_8578);
xor U9456 (N_9456,N_8528,N_8866);
nand U9457 (N_9457,N_7570,N_7640);
or U9458 (N_9458,N_8431,N_7821);
nand U9459 (N_9459,N_8575,N_8992);
and U9460 (N_9460,N_7734,N_8848);
nand U9461 (N_9461,N_8414,N_8061);
nor U9462 (N_9462,N_8776,N_8254);
xor U9463 (N_9463,N_8229,N_8839);
nor U9464 (N_9464,N_8533,N_8448);
nand U9465 (N_9465,N_8893,N_8453);
or U9466 (N_9466,N_7804,N_7905);
and U9467 (N_9467,N_8930,N_7516);
or U9468 (N_9468,N_7684,N_8286);
nor U9469 (N_9469,N_8135,N_7784);
and U9470 (N_9470,N_7813,N_7605);
and U9471 (N_9471,N_7769,N_8411);
nand U9472 (N_9472,N_8115,N_8273);
xor U9473 (N_9473,N_8762,N_8092);
nand U9474 (N_9474,N_7625,N_8541);
nor U9475 (N_9475,N_7594,N_8179);
and U9476 (N_9476,N_7653,N_8418);
nand U9477 (N_9477,N_7507,N_8655);
nor U9478 (N_9478,N_8413,N_7836);
nor U9479 (N_9479,N_8907,N_8605);
nand U9480 (N_9480,N_8140,N_8668);
nor U9481 (N_9481,N_7820,N_8592);
nand U9482 (N_9482,N_8773,N_7903);
or U9483 (N_9483,N_7512,N_8018);
and U9484 (N_9484,N_8168,N_8119);
nand U9485 (N_9485,N_7801,N_8604);
and U9486 (N_9486,N_8112,N_7872);
nor U9487 (N_9487,N_8207,N_8952);
nand U9488 (N_9488,N_7612,N_8184);
nor U9489 (N_9489,N_8357,N_8836);
or U9490 (N_9490,N_7839,N_8235);
or U9491 (N_9491,N_8058,N_8867);
or U9492 (N_9492,N_7621,N_7593);
xnor U9493 (N_9493,N_8950,N_8587);
nor U9494 (N_9494,N_7760,N_8494);
and U9495 (N_9495,N_8376,N_7906);
xnor U9496 (N_9496,N_8958,N_8662);
nor U9497 (N_9497,N_7743,N_8743);
and U9498 (N_9498,N_7652,N_8978);
nand U9499 (N_9499,N_8650,N_7943);
nand U9500 (N_9500,N_8504,N_8309);
nand U9501 (N_9501,N_8555,N_8354);
nor U9502 (N_9502,N_8108,N_7539);
and U9503 (N_9503,N_7841,N_8726);
nand U9504 (N_9504,N_8351,N_8353);
nor U9505 (N_9505,N_8059,N_8593);
or U9506 (N_9506,N_8905,N_8259);
and U9507 (N_9507,N_7837,N_7712);
nand U9508 (N_9508,N_8213,N_8052);
nand U9509 (N_9509,N_8481,N_8998);
and U9510 (N_9510,N_7816,N_8047);
nor U9511 (N_9511,N_8496,N_8615);
nor U9512 (N_9512,N_8974,N_8077);
nor U9513 (N_9513,N_8843,N_8722);
nand U9514 (N_9514,N_8954,N_7967);
or U9515 (N_9515,N_8805,N_8281);
nor U9516 (N_9516,N_7680,N_8940);
and U9517 (N_9517,N_8759,N_8870);
or U9518 (N_9518,N_7982,N_8127);
nor U9519 (N_9519,N_8983,N_8344);
nor U9520 (N_9520,N_8375,N_7777);
nand U9521 (N_9521,N_7744,N_7755);
nand U9522 (N_9522,N_7514,N_7567);
nand U9523 (N_9523,N_8918,N_8818);
or U9524 (N_9524,N_8932,N_7639);
nand U9525 (N_9525,N_8788,N_8444);
and U9526 (N_9526,N_7730,N_8841);
nor U9527 (N_9527,N_8015,N_7871);
xnor U9528 (N_9528,N_8310,N_7545);
xnor U9529 (N_9529,N_8670,N_8965);
or U9530 (N_9530,N_7582,N_7540);
or U9531 (N_9531,N_8519,N_8387);
and U9532 (N_9532,N_7873,N_8158);
and U9533 (N_9533,N_8964,N_7535);
nand U9534 (N_9534,N_8535,N_8174);
nand U9535 (N_9535,N_7635,N_7806);
and U9536 (N_9536,N_8631,N_8959);
nand U9537 (N_9537,N_7716,N_8318);
nand U9538 (N_9538,N_7548,N_8585);
or U9539 (N_9539,N_8752,N_8569);
or U9540 (N_9540,N_7925,N_8727);
xor U9541 (N_9541,N_8815,N_8050);
nor U9542 (N_9542,N_8056,N_8278);
and U9543 (N_9543,N_7834,N_7685);
nor U9544 (N_9544,N_8188,N_7692);
xor U9545 (N_9545,N_8597,N_8154);
or U9546 (N_9546,N_8355,N_8065);
nand U9547 (N_9547,N_8134,N_8280);
nand U9548 (N_9548,N_8035,N_7852);
nor U9549 (N_9549,N_8962,N_8939);
xnor U9550 (N_9550,N_8042,N_8104);
nand U9551 (N_9551,N_8966,N_8645);
or U9552 (N_9552,N_7986,N_8904);
nor U9553 (N_9553,N_7987,N_8107);
xor U9554 (N_9554,N_8340,N_8279);
nand U9555 (N_9555,N_7840,N_8210);
or U9556 (N_9556,N_8001,N_8024);
or U9557 (N_9557,N_8233,N_8399);
nor U9558 (N_9558,N_8674,N_8600);
and U9559 (N_9559,N_8756,N_8850);
or U9560 (N_9560,N_8677,N_8000);
nor U9561 (N_9561,N_8049,N_8560);
and U9562 (N_9562,N_8862,N_8673);
nand U9563 (N_9563,N_8322,N_7909);
nand U9564 (N_9564,N_8348,N_8723);
and U9565 (N_9565,N_8630,N_7894);
nor U9566 (N_9566,N_7759,N_8664);
and U9567 (N_9567,N_7627,N_7515);
or U9568 (N_9568,N_8432,N_8128);
and U9569 (N_9569,N_7576,N_8875);
and U9570 (N_9570,N_8854,N_8806);
or U9571 (N_9571,N_8133,N_7918);
xor U9572 (N_9572,N_8667,N_7948);
and U9573 (N_9573,N_8187,N_8203);
and U9574 (N_9574,N_7772,N_7829);
and U9575 (N_9575,N_7761,N_8404);
nor U9576 (N_9576,N_7861,N_7738);
or U9577 (N_9577,N_7589,N_7592);
or U9578 (N_9578,N_8883,N_8402);
nand U9579 (N_9579,N_8002,N_8066);
nand U9580 (N_9580,N_7984,N_8561);
xor U9581 (N_9581,N_8861,N_7676);
nand U9582 (N_9582,N_7677,N_7902);
or U9583 (N_9583,N_8258,N_8617);
xnor U9584 (N_9584,N_8704,N_8285);
and U9585 (N_9585,N_8474,N_7718);
nor U9586 (N_9586,N_8395,N_8455);
and U9587 (N_9587,N_8341,N_8484);
nand U9588 (N_9588,N_8037,N_8558);
and U9589 (N_9589,N_8439,N_8300);
or U9590 (N_9590,N_8935,N_8985);
and U9591 (N_9591,N_8925,N_7762);
and U9592 (N_9592,N_7797,N_7696);
xor U9593 (N_9593,N_7732,N_8458);
nand U9594 (N_9594,N_7884,N_8799);
nand U9595 (N_9595,N_8618,N_8085);
and U9596 (N_9596,N_7961,N_7575);
nor U9597 (N_9597,N_7778,N_7672);
nand U9598 (N_9598,N_8191,N_7972);
nor U9599 (N_9599,N_8161,N_7715);
nand U9600 (N_9600,N_7717,N_8595);
nor U9601 (N_9601,N_7952,N_7561);
or U9602 (N_9602,N_8923,N_7647);
and U9603 (N_9603,N_7705,N_8429);
nor U9604 (N_9604,N_7637,N_8542);
or U9605 (N_9605,N_8017,N_8691);
nand U9606 (N_9606,N_8493,N_8121);
nand U9607 (N_9607,N_8833,N_7792);
nand U9608 (N_9608,N_8068,N_7598);
or U9609 (N_9609,N_7842,N_8305);
xnor U9610 (N_9610,N_8865,N_8373);
nand U9611 (N_9611,N_7628,N_8651);
nand U9612 (N_9612,N_8020,N_8069);
or U9613 (N_9613,N_8010,N_8243);
or U9614 (N_9614,N_7528,N_8106);
or U9615 (N_9615,N_7544,N_8680);
nand U9616 (N_9616,N_7866,N_8710);
nand U9617 (N_9617,N_8610,N_7747);
and U9618 (N_9618,N_7735,N_7666);
and U9619 (N_9619,N_8098,N_8888);
nand U9620 (N_9620,N_8057,N_8111);
and U9621 (N_9621,N_8290,N_8289);
nand U9622 (N_9622,N_8489,N_8991);
xnor U9623 (N_9623,N_7714,N_8782);
and U9624 (N_9624,N_8485,N_8206);
and U9625 (N_9625,N_7529,N_8248);
nand U9626 (N_9626,N_8169,N_8396);
and U9627 (N_9627,N_8326,N_7595);
nand U9628 (N_9628,N_8425,N_8117);
nor U9629 (N_9629,N_8508,N_8984);
nand U9630 (N_9630,N_8639,N_8029);
and U9631 (N_9631,N_8086,N_8464);
and U9632 (N_9632,N_8679,N_8497);
or U9633 (N_9633,N_7681,N_8712);
and U9634 (N_9634,N_7531,N_7927);
nand U9635 (N_9635,N_8347,N_8304);
or U9636 (N_9636,N_7733,N_8067);
or U9637 (N_9637,N_8238,N_7541);
nor U9638 (N_9638,N_7947,N_7895);
or U9639 (N_9639,N_7996,N_7930);
xnor U9640 (N_9640,N_8417,N_8750);
and U9641 (N_9641,N_7632,N_7746);
nor U9642 (N_9642,N_8571,N_7502);
or U9643 (N_9643,N_8708,N_8205);
or U9644 (N_9644,N_8040,N_7915);
or U9645 (N_9645,N_7971,N_8472);
or U9646 (N_9646,N_8323,N_8730);
nand U9647 (N_9647,N_8594,N_8221);
and U9648 (N_9648,N_7766,N_8522);
or U9649 (N_9649,N_7553,N_7908);
or U9650 (N_9650,N_8071,N_8599);
or U9651 (N_9651,N_8030,N_8390);
or U9652 (N_9652,N_8409,N_8021);
nand U9653 (N_9653,N_7988,N_8251);
nor U9654 (N_9654,N_8033,N_8028);
or U9655 (N_9655,N_8317,N_8193);
or U9656 (N_9656,N_7552,N_8916);
nor U9657 (N_9657,N_8588,N_8434);
or U9658 (N_9658,N_7583,N_8768);
nand U9659 (N_9659,N_7510,N_8968);
and U9660 (N_9660,N_8291,N_8986);
nor U9661 (N_9661,N_8202,N_8693);
nand U9662 (N_9662,N_7710,N_7645);
and U9663 (N_9663,N_7935,N_8034);
and U9664 (N_9664,N_8204,N_7960);
or U9665 (N_9665,N_7979,N_8466);
xor U9666 (N_9666,N_8287,N_8159);
and U9667 (N_9667,N_8626,N_8783);
nand U9668 (N_9668,N_7596,N_7591);
nand U9669 (N_9669,N_8378,N_8573);
nor U9670 (N_9670,N_8247,N_7568);
nor U9671 (N_9671,N_8109,N_7584);
nand U9672 (N_9672,N_8665,N_8170);
or U9673 (N_9673,N_8241,N_7989);
nor U9674 (N_9674,N_7980,N_8757);
and U9675 (N_9675,N_7690,N_8661);
nor U9676 (N_9676,N_8580,N_8219);
or U9677 (N_9677,N_8857,N_7964);
nand U9678 (N_9678,N_7828,N_7978);
nand U9679 (N_9679,N_8513,N_8831);
xnor U9680 (N_9680,N_7520,N_7933);
nor U9681 (N_9681,N_8577,N_7874);
and U9682 (N_9682,N_8694,N_7809);
or U9683 (N_9683,N_7926,N_8697);
nand U9684 (N_9684,N_8902,N_8549);
nand U9685 (N_9685,N_7521,N_7923);
nand U9686 (N_9686,N_8784,N_8337);
or U9687 (N_9687,N_8897,N_7500);
nand U9688 (N_9688,N_8405,N_7910);
or U9689 (N_9689,N_8487,N_8136);
nor U9690 (N_9690,N_7865,N_7622);
or U9691 (N_9691,N_7824,N_8043);
nor U9692 (N_9692,N_7533,N_8070);
and U9693 (N_9693,N_8729,N_8827);
nor U9694 (N_9694,N_7599,N_8891);
or U9695 (N_9695,N_7999,N_8524);
nor U9696 (N_9696,N_7817,N_8162);
nor U9697 (N_9697,N_7527,N_8874);
or U9698 (N_9698,N_7789,N_7998);
nor U9699 (N_9699,N_8559,N_8703);
or U9700 (N_9700,N_7623,N_8124);
or U9701 (N_9701,N_8981,N_8172);
xnor U9702 (N_9702,N_8377,N_8769);
and U9703 (N_9703,N_8796,N_8737);
and U9704 (N_9704,N_8451,N_8476);
or U9705 (N_9705,N_8538,N_8401);
nor U9706 (N_9706,N_7654,N_8253);
xnor U9707 (N_9707,N_8913,N_7600);
nand U9708 (N_9708,N_7723,N_7750);
and U9709 (N_9709,N_8041,N_7814);
and U9710 (N_9710,N_8510,N_8646);
nand U9711 (N_9711,N_8197,N_8801);
nor U9712 (N_9712,N_7882,N_8707);
or U9713 (N_9713,N_8717,N_7796);
nand U9714 (N_9714,N_7826,N_8602);
nor U9715 (N_9715,N_7775,N_8303);
nor U9716 (N_9716,N_8063,N_8220);
or U9717 (N_9717,N_7683,N_7587);
nor U9718 (N_9718,N_7907,N_7976);
or U9719 (N_9719,N_8120,N_8146);
xor U9720 (N_9720,N_8706,N_8260);
or U9721 (N_9721,N_8738,N_8945);
or U9722 (N_9722,N_8331,N_7819);
xor U9723 (N_9723,N_8332,N_7549);
nand U9724 (N_9724,N_8420,N_8346);
nor U9725 (N_9725,N_7992,N_8746);
nor U9726 (N_9726,N_7864,N_7721);
and U9727 (N_9727,N_7686,N_7957);
or U9728 (N_9728,N_8460,N_8306);
or U9729 (N_9729,N_8676,N_8582);
and U9730 (N_9730,N_7854,N_8102);
nand U9731 (N_9731,N_7547,N_7830);
or U9732 (N_9732,N_8823,N_8249);
nand U9733 (N_9733,N_8032,N_8774);
nor U9734 (N_9734,N_8934,N_8433);
nand U9735 (N_9735,N_8556,N_8530);
nand U9736 (N_9736,N_7885,N_7934);
nor U9737 (N_9737,N_8963,N_7650);
nor U9738 (N_9738,N_8352,N_8955);
nand U9739 (N_9739,N_8167,N_8545);
or U9740 (N_9740,N_8125,N_7546);
nand U9741 (N_9741,N_8669,N_8637);
nor U9742 (N_9742,N_8520,N_7859);
nand U9743 (N_9743,N_8632,N_8338);
and U9744 (N_9744,N_8369,N_8048);
nor U9745 (N_9745,N_8391,N_7991);
and U9746 (N_9746,N_8772,N_8760);
and U9747 (N_9747,N_8589,N_7603);
and U9748 (N_9748,N_8194,N_7924);
or U9749 (N_9749,N_8713,N_7776);
nor U9750 (N_9750,N_7551,N_7864);
or U9751 (N_9751,N_8185,N_7708);
or U9752 (N_9752,N_8309,N_8552);
nand U9753 (N_9753,N_8380,N_8632);
nor U9754 (N_9754,N_7663,N_8273);
nor U9755 (N_9755,N_8664,N_7798);
or U9756 (N_9756,N_8540,N_8955);
and U9757 (N_9757,N_8178,N_7758);
xnor U9758 (N_9758,N_8830,N_8421);
nor U9759 (N_9759,N_7627,N_7917);
or U9760 (N_9760,N_8303,N_8757);
or U9761 (N_9761,N_8441,N_8395);
or U9762 (N_9762,N_7727,N_8450);
nand U9763 (N_9763,N_8793,N_7510);
and U9764 (N_9764,N_8960,N_7822);
nor U9765 (N_9765,N_8313,N_8588);
or U9766 (N_9766,N_8999,N_7889);
xor U9767 (N_9767,N_8332,N_7904);
nand U9768 (N_9768,N_8187,N_7810);
nor U9769 (N_9769,N_8171,N_8916);
nand U9770 (N_9770,N_7835,N_8150);
and U9771 (N_9771,N_7603,N_7766);
and U9772 (N_9772,N_8660,N_8807);
nor U9773 (N_9773,N_8595,N_7814);
nand U9774 (N_9774,N_7655,N_8349);
and U9775 (N_9775,N_8438,N_7566);
and U9776 (N_9776,N_7510,N_8930);
nor U9777 (N_9777,N_8362,N_8260);
nor U9778 (N_9778,N_8491,N_7630);
and U9779 (N_9779,N_8950,N_7672);
nor U9780 (N_9780,N_8815,N_8836);
or U9781 (N_9781,N_7985,N_8321);
and U9782 (N_9782,N_8073,N_8245);
xnor U9783 (N_9783,N_7942,N_7719);
or U9784 (N_9784,N_8912,N_8010);
and U9785 (N_9785,N_8703,N_8004);
and U9786 (N_9786,N_8749,N_8121);
nand U9787 (N_9787,N_7995,N_8783);
nand U9788 (N_9788,N_7670,N_8790);
and U9789 (N_9789,N_8900,N_8613);
nand U9790 (N_9790,N_8015,N_8067);
and U9791 (N_9791,N_8808,N_7889);
and U9792 (N_9792,N_8975,N_8213);
and U9793 (N_9793,N_7541,N_8196);
and U9794 (N_9794,N_8988,N_8063);
and U9795 (N_9795,N_8877,N_8608);
or U9796 (N_9796,N_8168,N_8447);
nand U9797 (N_9797,N_8184,N_8372);
nand U9798 (N_9798,N_8733,N_8589);
or U9799 (N_9799,N_8556,N_8699);
xnor U9800 (N_9800,N_8688,N_8175);
nor U9801 (N_9801,N_8355,N_8112);
or U9802 (N_9802,N_8273,N_8706);
and U9803 (N_9803,N_8171,N_8581);
or U9804 (N_9804,N_8316,N_7622);
nand U9805 (N_9805,N_8821,N_8948);
or U9806 (N_9806,N_7838,N_7969);
nand U9807 (N_9807,N_8355,N_8221);
nor U9808 (N_9808,N_7865,N_8851);
nor U9809 (N_9809,N_8645,N_8894);
nor U9810 (N_9810,N_7610,N_8681);
or U9811 (N_9811,N_8232,N_8840);
or U9812 (N_9812,N_8228,N_8242);
xnor U9813 (N_9813,N_8634,N_8723);
nor U9814 (N_9814,N_8760,N_8820);
nand U9815 (N_9815,N_8952,N_7503);
nand U9816 (N_9816,N_8958,N_7886);
nand U9817 (N_9817,N_7866,N_7919);
and U9818 (N_9818,N_8724,N_8955);
or U9819 (N_9819,N_8296,N_7776);
and U9820 (N_9820,N_8405,N_8273);
nand U9821 (N_9821,N_7920,N_7939);
and U9822 (N_9822,N_8685,N_8691);
nand U9823 (N_9823,N_8888,N_8772);
or U9824 (N_9824,N_7592,N_8734);
or U9825 (N_9825,N_8423,N_8323);
nand U9826 (N_9826,N_8133,N_8595);
or U9827 (N_9827,N_8446,N_8305);
nor U9828 (N_9828,N_7642,N_7528);
or U9829 (N_9829,N_8477,N_8120);
nand U9830 (N_9830,N_7788,N_8890);
xor U9831 (N_9831,N_8280,N_8224);
xnor U9832 (N_9832,N_8270,N_8919);
nand U9833 (N_9833,N_8193,N_8381);
nor U9834 (N_9834,N_8235,N_8265);
nor U9835 (N_9835,N_8754,N_8822);
nand U9836 (N_9836,N_7617,N_7547);
xnor U9837 (N_9837,N_7653,N_8710);
xnor U9838 (N_9838,N_7998,N_8737);
and U9839 (N_9839,N_8947,N_7657);
nor U9840 (N_9840,N_8029,N_8509);
nor U9841 (N_9841,N_8383,N_7709);
nand U9842 (N_9842,N_8169,N_8960);
nor U9843 (N_9843,N_8815,N_8509);
xnor U9844 (N_9844,N_7583,N_8394);
nor U9845 (N_9845,N_8995,N_8747);
nor U9846 (N_9846,N_8921,N_7934);
and U9847 (N_9847,N_8165,N_8379);
nor U9848 (N_9848,N_7855,N_7970);
nand U9849 (N_9849,N_8507,N_8331);
or U9850 (N_9850,N_7994,N_7518);
nand U9851 (N_9851,N_7605,N_7673);
nor U9852 (N_9852,N_7847,N_7512);
and U9853 (N_9853,N_8552,N_8305);
nand U9854 (N_9854,N_8675,N_7929);
nand U9855 (N_9855,N_7565,N_8834);
and U9856 (N_9856,N_8348,N_8586);
and U9857 (N_9857,N_7723,N_8338);
nor U9858 (N_9858,N_7891,N_8074);
nor U9859 (N_9859,N_8084,N_7513);
nor U9860 (N_9860,N_8293,N_7885);
nand U9861 (N_9861,N_8962,N_8082);
and U9862 (N_9862,N_7592,N_8253);
or U9863 (N_9863,N_8544,N_8576);
nor U9864 (N_9864,N_8864,N_7723);
and U9865 (N_9865,N_8509,N_8941);
nor U9866 (N_9866,N_8800,N_8993);
nor U9867 (N_9867,N_8617,N_7944);
and U9868 (N_9868,N_8069,N_8815);
nand U9869 (N_9869,N_8574,N_8741);
or U9870 (N_9870,N_7604,N_8327);
and U9871 (N_9871,N_7926,N_8557);
and U9872 (N_9872,N_7505,N_7875);
and U9873 (N_9873,N_8808,N_8470);
nand U9874 (N_9874,N_8312,N_8384);
nor U9875 (N_9875,N_8450,N_7757);
nor U9876 (N_9876,N_7960,N_8134);
or U9877 (N_9877,N_8391,N_8709);
or U9878 (N_9878,N_8525,N_8904);
nor U9879 (N_9879,N_8476,N_7718);
and U9880 (N_9880,N_8151,N_8053);
or U9881 (N_9881,N_7692,N_7902);
nand U9882 (N_9882,N_8950,N_7886);
nand U9883 (N_9883,N_8065,N_7979);
nand U9884 (N_9884,N_8418,N_7647);
nand U9885 (N_9885,N_7836,N_8918);
or U9886 (N_9886,N_8609,N_8462);
or U9887 (N_9887,N_8653,N_7770);
nor U9888 (N_9888,N_8015,N_8285);
xor U9889 (N_9889,N_8052,N_8735);
and U9890 (N_9890,N_8130,N_8157);
xnor U9891 (N_9891,N_7955,N_8661);
nand U9892 (N_9892,N_7826,N_8843);
and U9893 (N_9893,N_8091,N_8606);
and U9894 (N_9894,N_7783,N_7965);
nor U9895 (N_9895,N_8370,N_8405);
nor U9896 (N_9896,N_7803,N_7544);
nand U9897 (N_9897,N_8707,N_8652);
and U9898 (N_9898,N_8570,N_8667);
nand U9899 (N_9899,N_8407,N_8903);
nand U9900 (N_9900,N_7755,N_7917);
nand U9901 (N_9901,N_8959,N_8713);
nor U9902 (N_9902,N_8592,N_8436);
nand U9903 (N_9903,N_8611,N_8692);
xnor U9904 (N_9904,N_8917,N_7844);
xor U9905 (N_9905,N_8324,N_7685);
and U9906 (N_9906,N_8854,N_8900);
or U9907 (N_9907,N_8483,N_7848);
xnor U9908 (N_9908,N_8431,N_8528);
and U9909 (N_9909,N_8453,N_8870);
or U9910 (N_9910,N_8047,N_7981);
and U9911 (N_9911,N_8404,N_7948);
and U9912 (N_9912,N_8085,N_8585);
and U9913 (N_9913,N_7912,N_8359);
or U9914 (N_9914,N_7580,N_8199);
nor U9915 (N_9915,N_8483,N_8209);
nand U9916 (N_9916,N_8236,N_7962);
nor U9917 (N_9917,N_7651,N_7886);
nor U9918 (N_9918,N_7606,N_7969);
and U9919 (N_9919,N_7702,N_7649);
nand U9920 (N_9920,N_7785,N_8120);
or U9921 (N_9921,N_8329,N_7567);
or U9922 (N_9922,N_8992,N_8314);
nand U9923 (N_9923,N_7773,N_8745);
nand U9924 (N_9924,N_8737,N_8776);
or U9925 (N_9925,N_8378,N_7811);
nand U9926 (N_9926,N_8272,N_7779);
and U9927 (N_9927,N_8150,N_8231);
or U9928 (N_9928,N_8593,N_8052);
or U9929 (N_9929,N_7935,N_8930);
or U9930 (N_9930,N_8071,N_7576);
nand U9931 (N_9931,N_7578,N_8747);
and U9932 (N_9932,N_8985,N_7896);
or U9933 (N_9933,N_8100,N_8613);
nand U9934 (N_9934,N_8042,N_7730);
or U9935 (N_9935,N_7867,N_8393);
nand U9936 (N_9936,N_8538,N_8674);
or U9937 (N_9937,N_8640,N_7847);
nor U9938 (N_9938,N_8448,N_7868);
nand U9939 (N_9939,N_8679,N_8249);
nand U9940 (N_9940,N_8210,N_8206);
or U9941 (N_9941,N_7533,N_7982);
and U9942 (N_9942,N_8308,N_8884);
and U9943 (N_9943,N_7773,N_7944);
and U9944 (N_9944,N_7930,N_8722);
nand U9945 (N_9945,N_8219,N_7975);
nor U9946 (N_9946,N_8766,N_7545);
nand U9947 (N_9947,N_8609,N_7905);
and U9948 (N_9948,N_8064,N_8004);
nor U9949 (N_9949,N_7997,N_8533);
xnor U9950 (N_9950,N_7721,N_8098);
nor U9951 (N_9951,N_8666,N_8220);
or U9952 (N_9952,N_8813,N_8782);
and U9953 (N_9953,N_8249,N_8527);
and U9954 (N_9954,N_8786,N_8511);
nor U9955 (N_9955,N_8796,N_8396);
nor U9956 (N_9956,N_7799,N_8079);
or U9957 (N_9957,N_8351,N_7606);
and U9958 (N_9958,N_7715,N_8365);
nor U9959 (N_9959,N_7922,N_8473);
nor U9960 (N_9960,N_8989,N_8184);
nor U9961 (N_9961,N_8580,N_7645);
nor U9962 (N_9962,N_8381,N_8731);
nor U9963 (N_9963,N_8368,N_8437);
nand U9964 (N_9964,N_7720,N_7808);
nor U9965 (N_9965,N_8122,N_8067);
or U9966 (N_9966,N_8048,N_7741);
nand U9967 (N_9967,N_8738,N_7572);
xnor U9968 (N_9968,N_8900,N_7550);
and U9969 (N_9969,N_7829,N_8721);
and U9970 (N_9970,N_8439,N_8766);
nand U9971 (N_9971,N_7944,N_7852);
and U9972 (N_9972,N_8600,N_8962);
nand U9973 (N_9973,N_8562,N_8610);
or U9974 (N_9974,N_8513,N_7629);
nand U9975 (N_9975,N_7856,N_8402);
nor U9976 (N_9976,N_7916,N_8409);
nor U9977 (N_9977,N_8411,N_8616);
and U9978 (N_9978,N_8433,N_8120);
nand U9979 (N_9979,N_8570,N_8260);
xnor U9980 (N_9980,N_8333,N_8176);
nor U9981 (N_9981,N_8232,N_7849);
nor U9982 (N_9982,N_8891,N_8298);
nor U9983 (N_9983,N_8717,N_7539);
nand U9984 (N_9984,N_8020,N_8853);
nor U9985 (N_9985,N_7754,N_7731);
and U9986 (N_9986,N_7753,N_8059);
nand U9987 (N_9987,N_7620,N_8005);
nand U9988 (N_9988,N_8939,N_7590);
and U9989 (N_9989,N_7516,N_8252);
nand U9990 (N_9990,N_8346,N_8505);
nand U9991 (N_9991,N_8388,N_8932);
nor U9992 (N_9992,N_7751,N_8776);
and U9993 (N_9993,N_8321,N_8773);
nand U9994 (N_9994,N_8449,N_8172);
and U9995 (N_9995,N_7695,N_8281);
and U9996 (N_9996,N_8908,N_8746);
or U9997 (N_9997,N_8066,N_8620);
nor U9998 (N_9998,N_8234,N_8755);
nand U9999 (N_9999,N_8635,N_7956);
nor U10000 (N_10000,N_7666,N_7551);
nor U10001 (N_10001,N_8125,N_7529);
nand U10002 (N_10002,N_8174,N_7774);
or U10003 (N_10003,N_8946,N_8150);
nand U10004 (N_10004,N_7567,N_7650);
and U10005 (N_10005,N_7828,N_7690);
or U10006 (N_10006,N_7612,N_8654);
nor U10007 (N_10007,N_7546,N_8915);
nor U10008 (N_10008,N_8491,N_8219);
or U10009 (N_10009,N_8165,N_7640);
or U10010 (N_10010,N_8171,N_8379);
and U10011 (N_10011,N_8585,N_8492);
nand U10012 (N_10012,N_8880,N_8109);
or U10013 (N_10013,N_7926,N_8980);
or U10014 (N_10014,N_7634,N_8464);
or U10015 (N_10015,N_7859,N_8036);
nand U10016 (N_10016,N_8617,N_8337);
xor U10017 (N_10017,N_8370,N_7571);
and U10018 (N_10018,N_8149,N_8440);
and U10019 (N_10019,N_8201,N_8019);
or U10020 (N_10020,N_7774,N_7875);
or U10021 (N_10021,N_7738,N_8504);
nand U10022 (N_10022,N_7794,N_7741);
nor U10023 (N_10023,N_7711,N_8841);
nand U10024 (N_10024,N_7782,N_8170);
xor U10025 (N_10025,N_8140,N_7720);
nor U10026 (N_10026,N_7765,N_7809);
and U10027 (N_10027,N_7750,N_7514);
nor U10028 (N_10028,N_8705,N_8865);
or U10029 (N_10029,N_8966,N_8174);
nor U10030 (N_10030,N_8713,N_8707);
and U10031 (N_10031,N_7714,N_8332);
xor U10032 (N_10032,N_8970,N_8436);
nor U10033 (N_10033,N_8235,N_7642);
and U10034 (N_10034,N_7530,N_8467);
or U10035 (N_10035,N_8216,N_8801);
and U10036 (N_10036,N_8130,N_8398);
nor U10037 (N_10037,N_7593,N_7760);
nor U10038 (N_10038,N_7763,N_7857);
and U10039 (N_10039,N_8890,N_7981);
and U10040 (N_10040,N_8237,N_8327);
and U10041 (N_10041,N_8194,N_7699);
nor U10042 (N_10042,N_7513,N_8807);
or U10043 (N_10043,N_7741,N_8886);
nand U10044 (N_10044,N_8098,N_7689);
nor U10045 (N_10045,N_8031,N_7860);
or U10046 (N_10046,N_7588,N_7566);
nand U10047 (N_10047,N_8729,N_7685);
or U10048 (N_10048,N_7834,N_8571);
and U10049 (N_10049,N_7805,N_8064);
or U10050 (N_10050,N_8585,N_8868);
and U10051 (N_10051,N_8527,N_8310);
nand U10052 (N_10052,N_8876,N_7917);
xor U10053 (N_10053,N_7895,N_8539);
nor U10054 (N_10054,N_8367,N_8568);
or U10055 (N_10055,N_8492,N_8804);
and U10056 (N_10056,N_8225,N_8650);
nor U10057 (N_10057,N_7678,N_8954);
or U10058 (N_10058,N_8122,N_8807);
or U10059 (N_10059,N_8967,N_7722);
and U10060 (N_10060,N_7653,N_7548);
nand U10061 (N_10061,N_8746,N_8020);
nand U10062 (N_10062,N_8931,N_8840);
nor U10063 (N_10063,N_8822,N_8165);
nor U10064 (N_10064,N_8831,N_8663);
and U10065 (N_10065,N_8193,N_7981);
nand U10066 (N_10066,N_7922,N_8184);
and U10067 (N_10067,N_8880,N_8461);
nor U10068 (N_10068,N_8056,N_8062);
or U10069 (N_10069,N_8016,N_7967);
xnor U10070 (N_10070,N_8138,N_7755);
and U10071 (N_10071,N_8991,N_7716);
nand U10072 (N_10072,N_8086,N_8597);
nor U10073 (N_10073,N_8880,N_8870);
nor U10074 (N_10074,N_8476,N_8099);
nor U10075 (N_10075,N_8954,N_8100);
or U10076 (N_10076,N_7594,N_7836);
nor U10077 (N_10077,N_8281,N_8986);
or U10078 (N_10078,N_7542,N_7763);
nand U10079 (N_10079,N_8634,N_8113);
or U10080 (N_10080,N_7865,N_8405);
and U10081 (N_10081,N_8353,N_8227);
nor U10082 (N_10082,N_8088,N_8019);
nor U10083 (N_10083,N_8402,N_8088);
nor U10084 (N_10084,N_7939,N_7980);
nor U10085 (N_10085,N_8703,N_7970);
and U10086 (N_10086,N_8282,N_8285);
and U10087 (N_10087,N_8627,N_7505);
and U10088 (N_10088,N_7611,N_8072);
nand U10089 (N_10089,N_7664,N_7672);
xor U10090 (N_10090,N_7844,N_7706);
nor U10091 (N_10091,N_8464,N_7823);
and U10092 (N_10092,N_8647,N_8854);
xor U10093 (N_10093,N_7636,N_8465);
or U10094 (N_10094,N_7995,N_7555);
nor U10095 (N_10095,N_8379,N_8534);
or U10096 (N_10096,N_7524,N_8550);
nor U10097 (N_10097,N_8615,N_7950);
nor U10098 (N_10098,N_8371,N_8068);
nor U10099 (N_10099,N_8534,N_7745);
nand U10100 (N_10100,N_8996,N_7528);
or U10101 (N_10101,N_8167,N_7515);
xor U10102 (N_10102,N_7733,N_8273);
and U10103 (N_10103,N_8222,N_8326);
and U10104 (N_10104,N_8227,N_7590);
nor U10105 (N_10105,N_7552,N_8642);
xnor U10106 (N_10106,N_7863,N_8488);
nand U10107 (N_10107,N_7768,N_8375);
nand U10108 (N_10108,N_7679,N_8148);
and U10109 (N_10109,N_7676,N_7873);
nand U10110 (N_10110,N_7614,N_8227);
nand U10111 (N_10111,N_8441,N_8283);
nand U10112 (N_10112,N_8106,N_8992);
and U10113 (N_10113,N_8524,N_8754);
nor U10114 (N_10114,N_7541,N_8825);
or U10115 (N_10115,N_8620,N_8168);
or U10116 (N_10116,N_8731,N_8070);
nor U10117 (N_10117,N_7741,N_7772);
nor U10118 (N_10118,N_8978,N_7774);
nor U10119 (N_10119,N_8762,N_7871);
and U10120 (N_10120,N_7933,N_7807);
or U10121 (N_10121,N_8593,N_7829);
nor U10122 (N_10122,N_8750,N_8499);
or U10123 (N_10123,N_7967,N_8734);
and U10124 (N_10124,N_8182,N_8930);
nand U10125 (N_10125,N_8113,N_8654);
and U10126 (N_10126,N_8430,N_8819);
or U10127 (N_10127,N_8695,N_8663);
nand U10128 (N_10128,N_8555,N_8723);
and U10129 (N_10129,N_7698,N_8073);
nand U10130 (N_10130,N_7614,N_8805);
or U10131 (N_10131,N_7768,N_8070);
nand U10132 (N_10132,N_7689,N_8955);
or U10133 (N_10133,N_8354,N_8902);
or U10134 (N_10134,N_8537,N_7514);
nand U10135 (N_10135,N_8183,N_8229);
and U10136 (N_10136,N_8234,N_8059);
xnor U10137 (N_10137,N_7915,N_7900);
nand U10138 (N_10138,N_7586,N_8135);
nand U10139 (N_10139,N_8113,N_8636);
or U10140 (N_10140,N_7877,N_8044);
nand U10141 (N_10141,N_7912,N_8761);
nor U10142 (N_10142,N_8875,N_8205);
and U10143 (N_10143,N_8966,N_8347);
nand U10144 (N_10144,N_7627,N_8083);
or U10145 (N_10145,N_7746,N_8756);
and U10146 (N_10146,N_8860,N_7586);
nand U10147 (N_10147,N_8638,N_7921);
nand U10148 (N_10148,N_7662,N_8005);
nor U10149 (N_10149,N_8148,N_7941);
and U10150 (N_10150,N_7905,N_7880);
nor U10151 (N_10151,N_7623,N_8305);
or U10152 (N_10152,N_8639,N_8173);
nor U10153 (N_10153,N_8318,N_8744);
or U10154 (N_10154,N_8410,N_8025);
xnor U10155 (N_10155,N_8538,N_8817);
and U10156 (N_10156,N_8155,N_8104);
and U10157 (N_10157,N_8516,N_7893);
nand U10158 (N_10158,N_7513,N_8447);
or U10159 (N_10159,N_7682,N_8807);
xnor U10160 (N_10160,N_8984,N_7898);
nor U10161 (N_10161,N_8816,N_8993);
and U10162 (N_10162,N_7593,N_7818);
xor U10163 (N_10163,N_7951,N_7785);
nor U10164 (N_10164,N_8718,N_8291);
or U10165 (N_10165,N_7840,N_8516);
nor U10166 (N_10166,N_8909,N_8069);
nand U10167 (N_10167,N_7524,N_7974);
nand U10168 (N_10168,N_8271,N_8250);
nand U10169 (N_10169,N_8049,N_8059);
or U10170 (N_10170,N_8300,N_8284);
and U10171 (N_10171,N_8877,N_7926);
nor U10172 (N_10172,N_8964,N_8166);
or U10173 (N_10173,N_7726,N_8817);
or U10174 (N_10174,N_7711,N_8694);
or U10175 (N_10175,N_8860,N_7507);
or U10176 (N_10176,N_8279,N_8735);
and U10177 (N_10177,N_8102,N_8153);
nor U10178 (N_10178,N_7787,N_8604);
nor U10179 (N_10179,N_8897,N_8917);
and U10180 (N_10180,N_8356,N_8370);
nor U10181 (N_10181,N_8677,N_7967);
and U10182 (N_10182,N_7696,N_7659);
and U10183 (N_10183,N_8901,N_8129);
nand U10184 (N_10184,N_8591,N_8362);
and U10185 (N_10185,N_7656,N_8560);
nand U10186 (N_10186,N_7520,N_7786);
or U10187 (N_10187,N_8407,N_7996);
or U10188 (N_10188,N_7684,N_7734);
and U10189 (N_10189,N_7748,N_8234);
or U10190 (N_10190,N_7644,N_7618);
xnor U10191 (N_10191,N_8245,N_7911);
nor U10192 (N_10192,N_7650,N_8384);
or U10193 (N_10193,N_8543,N_7838);
nor U10194 (N_10194,N_7911,N_7602);
nand U10195 (N_10195,N_8428,N_8003);
nand U10196 (N_10196,N_8018,N_8734);
or U10197 (N_10197,N_7751,N_8530);
xnor U10198 (N_10198,N_8519,N_8245);
nor U10199 (N_10199,N_8910,N_7891);
nand U10200 (N_10200,N_8730,N_8844);
nand U10201 (N_10201,N_8865,N_7679);
or U10202 (N_10202,N_8426,N_7778);
or U10203 (N_10203,N_7547,N_7852);
nor U10204 (N_10204,N_8149,N_7671);
and U10205 (N_10205,N_8170,N_8928);
and U10206 (N_10206,N_8235,N_8771);
xor U10207 (N_10207,N_8392,N_7749);
nand U10208 (N_10208,N_8888,N_8145);
or U10209 (N_10209,N_8251,N_8675);
and U10210 (N_10210,N_8367,N_7740);
or U10211 (N_10211,N_8276,N_8622);
nand U10212 (N_10212,N_8141,N_8577);
nor U10213 (N_10213,N_8315,N_8977);
or U10214 (N_10214,N_7614,N_7998);
nor U10215 (N_10215,N_8677,N_8161);
nor U10216 (N_10216,N_8634,N_7635);
or U10217 (N_10217,N_8194,N_8191);
and U10218 (N_10218,N_7521,N_8733);
nor U10219 (N_10219,N_7585,N_8420);
nor U10220 (N_10220,N_8145,N_8732);
xor U10221 (N_10221,N_8096,N_8504);
nor U10222 (N_10222,N_7610,N_8412);
and U10223 (N_10223,N_7612,N_7868);
or U10224 (N_10224,N_7734,N_7618);
xor U10225 (N_10225,N_8261,N_8071);
nor U10226 (N_10226,N_8099,N_8021);
nor U10227 (N_10227,N_8722,N_8347);
or U10228 (N_10228,N_7540,N_8956);
and U10229 (N_10229,N_8801,N_8520);
nor U10230 (N_10230,N_8365,N_8637);
xor U10231 (N_10231,N_8215,N_7674);
xnor U10232 (N_10232,N_8466,N_7659);
or U10233 (N_10233,N_8335,N_8779);
nor U10234 (N_10234,N_7528,N_8016);
nor U10235 (N_10235,N_7785,N_7968);
and U10236 (N_10236,N_8283,N_7742);
nor U10237 (N_10237,N_8302,N_7645);
nand U10238 (N_10238,N_8054,N_8505);
nand U10239 (N_10239,N_7871,N_8695);
nand U10240 (N_10240,N_8118,N_8525);
nor U10241 (N_10241,N_7570,N_8288);
nand U10242 (N_10242,N_8855,N_7769);
nor U10243 (N_10243,N_8810,N_7695);
nand U10244 (N_10244,N_8469,N_8615);
and U10245 (N_10245,N_7768,N_7746);
and U10246 (N_10246,N_8691,N_8295);
and U10247 (N_10247,N_8355,N_8371);
and U10248 (N_10248,N_8162,N_8405);
and U10249 (N_10249,N_8930,N_8456);
nand U10250 (N_10250,N_7571,N_8951);
xor U10251 (N_10251,N_8037,N_7795);
nand U10252 (N_10252,N_7861,N_7823);
and U10253 (N_10253,N_8767,N_7869);
and U10254 (N_10254,N_7693,N_8121);
and U10255 (N_10255,N_8674,N_7725);
and U10256 (N_10256,N_8613,N_8904);
or U10257 (N_10257,N_8267,N_8375);
xnor U10258 (N_10258,N_7585,N_8430);
nand U10259 (N_10259,N_7671,N_8437);
xnor U10260 (N_10260,N_8057,N_7882);
xnor U10261 (N_10261,N_7940,N_8073);
nand U10262 (N_10262,N_8945,N_8914);
nand U10263 (N_10263,N_8341,N_8948);
and U10264 (N_10264,N_7644,N_7791);
nand U10265 (N_10265,N_8940,N_7777);
or U10266 (N_10266,N_8006,N_8145);
xor U10267 (N_10267,N_8841,N_8114);
or U10268 (N_10268,N_7783,N_8908);
nor U10269 (N_10269,N_8663,N_7854);
and U10270 (N_10270,N_8987,N_8327);
or U10271 (N_10271,N_8374,N_8970);
or U10272 (N_10272,N_8818,N_7638);
nor U10273 (N_10273,N_8281,N_8648);
xnor U10274 (N_10274,N_8650,N_8206);
or U10275 (N_10275,N_8729,N_8052);
and U10276 (N_10276,N_8003,N_8288);
or U10277 (N_10277,N_7660,N_7822);
xor U10278 (N_10278,N_8830,N_8118);
and U10279 (N_10279,N_7609,N_8253);
nand U10280 (N_10280,N_8937,N_8393);
and U10281 (N_10281,N_7559,N_8043);
or U10282 (N_10282,N_8373,N_8107);
nor U10283 (N_10283,N_8172,N_8865);
and U10284 (N_10284,N_8286,N_8633);
nor U10285 (N_10285,N_8460,N_8649);
nand U10286 (N_10286,N_8401,N_8805);
and U10287 (N_10287,N_8496,N_8570);
xnor U10288 (N_10288,N_8107,N_8672);
or U10289 (N_10289,N_7732,N_7794);
or U10290 (N_10290,N_8409,N_8302);
nor U10291 (N_10291,N_8675,N_8375);
or U10292 (N_10292,N_8863,N_7703);
nand U10293 (N_10293,N_7913,N_8415);
xnor U10294 (N_10294,N_8028,N_8942);
and U10295 (N_10295,N_8098,N_8724);
nor U10296 (N_10296,N_8354,N_8969);
xnor U10297 (N_10297,N_8427,N_8181);
xnor U10298 (N_10298,N_8432,N_7619);
xor U10299 (N_10299,N_8610,N_8194);
xor U10300 (N_10300,N_7640,N_7884);
or U10301 (N_10301,N_7942,N_8985);
nor U10302 (N_10302,N_8725,N_7699);
and U10303 (N_10303,N_8777,N_7583);
and U10304 (N_10304,N_7849,N_7569);
and U10305 (N_10305,N_8911,N_8525);
nand U10306 (N_10306,N_8081,N_7546);
and U10307 (N_10307,N_8012,N_7772);
nor U10308 (N_10308,N_8106,N_8423);
and U10309 (N_10309,N_8258,N_7884);
and U10310 (N_10310,N_8271,N_8960);
nand U10311 (N_10311,N_7555,N_8194);
nand U10312 (N_10312,N_8197,N_8273);
and U10313 (N_10313,N_8825,N_7557);
and U10314 (N_10314,N_7840,N_8528);
xor U10315 (N_10315,N_7737,N_7993);
or U10316 (N_10316,N_8497,N_8868);
and U10317 (N_10317,N_8015,N_7615);
nand U10318 (N_10318,N_7691,N_7663);
and U10319 (N_10319,N_8762,N_8477);
or U10320 (N_10320,N_8574,N_8243);
or U10321 (N_10321,N_7966,N_8925);
nor U10322 (N_10322,N_8354,N_8843);
or U10323 (N_10323,N_8756,N_8197);
or U10324 (N_10324,N_7595,N_7905);
nand U10325 (N_10325,N_7734,N_8931);
nor U10326 (N_10326,N_7668,N_7949);
and U10327 (N_10327,N_7775,N_8864);
nand U10328 (N_10328,N_7920,N_8669);
nor U10329 (N_10329,N_8889,N_8933);
or U10330 (N_10330,N_7664,N_8954);
nand U10331 (N_10331,N_7785,N_8406);
or U10332 (N_10332,N_7800,N_7737);
nor U10333 (N_10333,N_7887,N_8323);
or U10334 (N_10334,N_8734,N_7555);
nor U10335 (N_10335,N_8752,N_8851);
or U10336 (N_10336,N_7619,N_8323);
nor U10337 (N_10337,N_8351,N_7642);
or U10338 (N_10338,N_7821,N_8610);
nor U10339 (N_10339,N_8381,N_8444);
or U10340 (N_10340,N_8578,N_7706);
nor U10341 (N_10341,N_7923,N_8372);
nand U10342 (N_10342,N_7715,N_7582);
nor U10343 (N_10343,N_8660,N_7980);
and U10344 (N_10344,N_8001,N_8454);
or U10345 (N_10345,N_8737,N_7941);
and U10346 (N_10346,N_8959,N_8237);
xor U10347 (N_10347,N_8219,N_8232);
and U10348 (N_10348,N_8281,N_8334);
or U10349 (N_10349,N_8165,N_8405);
or U10350 (N_10350,N_8682,N_7716);
and U10351 (N_10351,N_7571,N_7888);
and U10352 (N_10352,N_7729,N_7835);
or U10353 (N_10353,N_8937,N_7974);
or U10354 (N_10354,N_8837,N_8801);
nand U10355 (N_10355,N_8102,N_7869);
and U10356 (N_10356,N_8039,N_7636);
or U10357 (N_10357,N_8384,N_8689);
or U10358 (N_10358,N_8130,N_8936);
xor U10359 (N_10359,N_7632,N_7823);
or U10360 (N_10360,N_8812,N_7510);
nand U10361 (N_10361,N_7676,N_8308);
nand U10362 (N_10362,N_8345,N_8916);
nand U10363 (N_10363,N_7891,N_8861);
nor U10364 (N_10364,N_7892,N_8191);
nor U10365 (N_10365,N_7580,N_8290);
and U10366 (N_10366,N_8966,N_8270);
and U10367 (N_10367,N_7972,N_8659);
or U10368 (N_10368,N_8180,N_8916);
xor U10369 (N_10369,N_8063,N_8166);
and U10370 (N_10370,N_8972,N_7824);
and U10371 (N_10371,N_8483,N_7654);
nand U10372 (N_10372,N_8397,N_8509);
and U10373 (N_10373,N_7937,N_8733);
nand U10374 (N_10374,N_8138,N_8994);
or U10375 (N_10375,N_8574,N_8873);
xnor U10376 (N_10376,N_7539,N_8801);
nand U10377 (N_10377,N_8291,N_8902);
and U10378 (N_10378,N_7893,N_8130);
or U10379 (N_10379,N_8214,N_8327);
and U10380 (N_10380,N_8929,N_7527);
nor U10381 (N_10381,N_8823,N_8503);
or U10382 (N_10382,N_7531,N_8701);
or U10383 (N_10383,N_8051,N_7778);
nor U10384 (N_10384,N_7857,N_8525);
or U10385 (N_10385,N_7963,N_8562);
nor U10386 (N_10386,N_8571,N_8662);
or U10387 (N_10387,N_7760,N_7879);
nor U10388 (N_10388,N_8276,N_8273);
nor U10389 (N_10389,N_7690,N_8465);
nand U10390 (N_10390,N_8539,N_8101);
nand U10391 (N_10391,N_8401,N_8870);
nand U10392 (N_10392,N_8535,N_7851);
xor U10393 (N_10393,N_8776,N_8009);
or U10394 (N_10394,N_7669,N_8133);
nor U10395 (N_10395,N_8405,N_7974);
nor U10396 (N_10396,N_8862,N_8711);
and U10397 (N_10397,N_7642,N_7547);
nand U10398 (N_10398,N_8028,N_8713);
or U10399 (N_10399,N_8634,N_8728);
nor U10400 (N_10400,N_8443,N_8176);
or U10401 (N_10401,N_8582,N_7518);
and U10402 (N_10402,N_8273,N_8870);
or U10403 (N_10403,N_8801,N_8852);
and U10404 (N_10404,N_8822,N_8802);
xor U10405 (N_10405,N_8476,N_8309);
nor U10406 (N_10406,N_7623,N_8203);
nor U10407 (N_10407,N_8017,N_7923);
nor U10408 (N_10408,N_8288,N_8923);
or U10409 (N_10409,N_8938,N_8546);
and U10410 (N_10410,N_7696,N_8494);
xor U10411 (N_10411,N_8633,N_8709);
nand U10412 (N_10412,N_7567,N_8528);
or U10413 (N_10413,N_7701,N_8173);
nand U10414 (N_10414,N_8612,N_7741);
and U10415 (N_10415,N_8496,N_7559);
and U10416 (N_10416,N_8759,N_8026);
or U10417 (N_10417,N_8371,N_8069);
and U10418 (N_10418,N_7835,N_7866);
nor U10419 (N_10419,N_7571,N_8905);
nor U10420 (N_10420,N_8606,N_7636);
or U10421 (N_10421,N_8316,N_8301);
or U10422 (N_10422,N_8478,N_8466);
xor U10423 (N_10423,N_8142,N_8302);
nand U10424 (N_10424,N_7550,N_8565);
xnor U10425 (N_10425,N_8450,N_8310);
nor U10426 (N_10426,N_8424,N_8498);
and U10427 (N_10427,N_8776,N_8984);
nand U10428 (N_10428,N_8587,N_8133);
nor U10429 (N_10429,N_8648,N_8421);
nand U10430 (N_10430,N_8072,N_8637);
and U10431 (N_10431,N_8925,N_7897);
xnor U10432 (N_10432,N_8019,N_8988);
and U10433 (N_10433,N_7642,N_8036);
or U10434 (N_10434,N_7878,N_8752);
nand U10435 (N_10435,N_7700,N_8525);
nor U10436 (N_10436,N_7992,N_8749);
or U10437 (N_10437,N_7568,N_7721);
or U10438 (N_10438,N_8495,N_7834);
nand U10439 (N_10439,N_8329,N_8489);
or U10440 (N_10440,N_8363,N_7926);
nor U10441 (N_10441,N_8499,N_8522);
nand U10442 (N_10442,N_7848,N_8534);
nor U10443 (N_10443,N_8200,N_8606);
nand U10444 (N_10444,N_8835,N_7745);
nand U10445 (N_10445,N_7812,N_8865);
or U10446 (N_10446,N_8318,N_7966);
and U10447 (N_10447,N_8762,N_8167);
and U10448 (N_10448,N_7696,N_7573);
and U10449 (N_10449,N_8723,N_7858);
nand U10450 (N_10450,N_8053,N_8038);
and U10451 (N_10451,N_7616,N_8158);
nand U10452 (N_10452,N_8820,N_7858);
nor U10453 (N_10453,N_7698,N_8253);
nor U10454 (N_10454,N_8054,N_8925);
and U10455 (N_10455,N_8500,N_8592);
nand U10456 (N_10456,N_8878,N_8063);
nand U10457 (N_10457,N_8816,N_8677);
nand U10458 (N_10458,N_8890,N_7578);
nor U10459 (N_10459,N_8349,N_7775);
nor U10460 (N_10460,N_7974,N_8591);
and U10461 (N_10461,N_7897,N_8162);
nor U10462 (N_10462,N_8473,N_7919);
or U10463 (N_10463,N_8212,N_7783);
xnor U10464 (N_10464,N_8389,N_7961);
and U10465 (N_10465,N_8364,N_7634);
nor U10466 (N_10466,N_8737,N_8307);
or U10467 (N_10467,N_8198,N_8058);
nand U10468 (N_10468,N_8418,N_7501);
nor U10469 (N_10469,N_8809,N_8960);
and U10470 (N_10470,N_7806,N_8678);
nor U10471 (N_10471,N_7798,N_8632);
and U10472 (N_10472,N_8780,N_8026);
or U10473 (N_10473,N_8536,N_8626);
nand U10474 (N_10474,N_8874,N_8112);
and U10475 (N_10475,N_8090,N_8082);
nor U10476 (N_10476,N_8248,N_8058);
nor U10477 (N_10477,N_8158,N_8413);
and U10478 (N_10478,N_8515,N_7837);
or U10479 (N_10479,N_8893,N_8660);
nand U10480 (N_10480,N_7712,N_7630);
nor U10481 (N_10481,N_8458,N_8802);
nand U10482 (N_10482,N_8278,N_8432);
or U10483 (N_10483,N_7936,N_8718);
and U10484 (N_10484,N_8577,N_8908);
xor U10485 (N_10485,N_7644,N_7637);
nor U10486 (N_10486,N_8186,N_8234);
nand U10487 (N_10487,N_7607,N_7553);
nor U10488 (N_10488,N_8374,N_7593);
xnor U10489 (N_10489,N_7649,N_8802);
or U10490 (N_10490,N_8519,N_7561);
and U10491 (N_10491,N_7676,N_8417);
and U10492 (N_10492,N_7803,N_7609);
or U10493 (N_10493,N_8042,N_7694);
nor U10494 (N_10494,N_8408,N_7957);
or U10495 (N_10495,N_8292,N_7592);
and U10496 (N_10496,N_8921,N_8147);
or U10497 (N_10497,N_7647,N_8541);
nor U10498 (N_10498,N_8311,N_8025);
or U10499 (N_10499,N_8934,N_8467);
and U10500 (N_10500,N_9468,N_10119);
nand U10501 (N_10501,N_10325,N_9601);
nor U10502 (N_10502,N_10042,N_10236);
or U10503 (N_10503,N_9883,N_9831);
xor U10504 (N_10504,N_10417,N_9543);
or U10505 (N_10505,N_9137,N_9642);
nor U10506 (N_10506,N_9788,N_9747);
or U10507 (N_10507,N_10321,N_9520);
and U10508 (N_10508,N_10403,N_9057);
and U10509 (N_10509,N_9536,N_9746);
nand U10510 (N_10510,N_9807,N_9308);
or U10511 (N_10511,N_10212,N_10137);
and U10512 (N_10512,N_9312,N_9272);
nor U10513 (N_10513,N_10012,N_10110);
or U10514 (N_10514,N_9313,N_9292);
xnor U10515 (N_10515,N_9623,N_9247);
nand U10516 (N_10516,N_9935,N_9342);
nor U10517 (N_10517,N_10335,N_9832);
nand U10518 (N_10518,N_9201,N_9123);
and U10519 (N_10519,N_10438,N_9855);
nand U10520 (N_10520,N_9439,N_9955);
xor U10521 (N_10521,N_9640,N_9989);
and U10522 (N_10522,N_9327,N_9671);
xor U10523 (N_10523,N_9084,N_9534);
xnor U10524 (N_10524,N_9514,N_9353);
nand U10525 (N_10525,N_10054,N_9230);
xor U10526 (N_10526,N_9693,N_9843);
or U10527 (N_10527,N_10105,N_9530);
nand U10528 (N_10528,N_9522,N_9714);
and U10529 (N_10529,N_10306,N_9618);
xnor U10530 (N_10530,N_9824,N_10388);
nand U10531 (N_10531,N_10223,N_9347);
and U10532 (N_10532,N_9134,N_9600);
nor U10533 (N_10533,N_9146,N_9262);
nor U10534 (N_10534,N_9849,N_10351);
nor U10535 (N_10535,N_9748,N_9836);
or U10536 (N_10536,N_9578,N_10375);
or U10537 (N_10537,N_10469,N_9075);
nor U10538 (N_10538,N_9248,N_9890);
or U10539 (N_10539,N_10220,N_9983);
nor U10540 (N_10540,N_10046,N_10314);
or U10541 (N_10541,N_10350,N_9840);
nor U10542 (N_10542,N_9772,N_9669);
xnor U10543 (N_10543,N_9677,N_9016);
xnor U10544 (N_10544,N_9310,N_9885);
or U10545 (N_10545,N_9765,N_9856);
xnor U10546 (N_10546,N_9968,N_10151);
xnor U10547 (N_10547,N_9304,N_10201);
nand U10548 (N_10548,N_10297,N_9394);
nand U10549 (N_10549,N_9863,N_10273);
nor U10550 (N_10550,N_9839,N_9834);
xor U10551 (N_10551,N_10034,N_9925);
and U10552 (N_10552,N_10455,N_9244);
or U10553 (N_10553,N_9859,N_9160);
or U10554 (N_10554,N_10198,N_9553);
nor U10555 (N_10555,N_10292,N_9675);
nor U10556 (N_10556,N_9239,N_9710);
nand U10557 (N_10557,N_9797,N_9546);
nand U10558 (N_10558,N_10287,N_10473);
nor U10559 (N_10559,N_9131,N_10424);
and U10560 (N_10560,N_9787,N_10193);
and U10561 (N_10561,N_10153,N_10421);
nand U10562 (N_10562,N_9791,N_9480);
xor U10563 (N_10563,N_9705,N_9185);
xor U10564 (N_10564,N_9919,N_10470);
or U10565 (N_10565,N_9343,N_10372);
and U10566 (N_10566,N_9178,N_9398);
or U10567 (N_10567,N_9172,N_9489);
nor U10568 (N_10568,N_10165,N_10032);
and U10569 (N_10569,N_9187,N_9626);
and U10570 (N_10570,N_10047,N_10057);
nand U10571 (N_10571,N_9574,N_10011);
nor U10572 (N_10572,N_10466,N_9805);
and U10573 (N_10573,N_9028,N_9109);
or U10574 (N_10574,N_9961,N_9275);
and U10575 (N_10575,N_9656,N_10142);
nor U10576 (N_10576,N_9736,N_10000);
nor U10577 (N_10577,N_9512,N_10363);
or U10578 (N_10578,N_9529,N_9683);
nand U10579 (N_10579,N_9778,N_9357);
nor U10580 (N_10580,N_9331,N_9022);
nor U10581 (N_10581,N_9587,N_9781);
and U10582 (N_10582,N_9375,N_10065);
nor U10583 (N_10583,N_9196,N_9257);
nand U10584 (N_10584,N_9061,N_10191);
nand U10585 (N_10585,N_9999,N_10126);
nor U10586 (N_10586,N_10208,N_9515);
or U10587 (N_10587,N_10019,N_9287);
xnor U10588 (N_10588,N_9161,N_10373);
and U10589 (N_10589,N_10060,N_10252);
nand U10590 (N_10590,N_9270,N_9742);
or U10591 (N_10591,N_10393,N_10104);
or U10592 (N_10592,N_10410,N_10213);
or U10593 (N_10593,N_10471,N_9660);
or U10594 (N_10594,N_10026,N_9804);
or U10595 (N_10595,N_10205,N_9361);
nor U10596 (N_10596,N_9090,N_10086);
or U10597 (N_10597,N_9619,N_9898);
or U10598 (N_10598,N_10443,N_9940);
or U10599 (N_10599,N_9909,N_10286);
nand U10600 (N_10600,N_9848,N_9337);
nand U10601 (N_10601,N_10474,N_9975);
or U10602 (N_10602,N_9088,N_9967);
xnor U10603 (N_10603,N_10380,N_10312);
or U10604 (N_10604,N_9702,N_9294);
nor U10605 (N_10605,N_10446,N_10094);
or U10606 (N_10606,N_9826,N_10371);
nor U10607 (N_10607,N_9535,N_10237);
nor U10608 (N_10608,N_9105,N_9737);
nand U10609 (N_10609,N_10376,N_10285);
and U10610 (N_10610,N_9221,N_9860);
and U10611 (N_10611,N_9127,N_9140);
nor U10612 (N_10612,N_10281,N_10345);
nor U10613 (N_10613,N_9756,N_10310);
or U10614 (N_10614,N_9235,N_10342);
nor U10615 (N_10615,N_10445,N_9667);
nor U10616 (N_10616,N_9401,N_10255);
nor U10617 (N_10617,N_9857,N_10313);
nor U10618 (N_10618,N_9567,N_9699);
and U10619 (N_10619,N_9540,N_9444);
nor U10620 (N_10620,N_9130,N_10066);
nor U10621 (N_10621,N_10383,N_9021);
and U10622 (N_10622,N_9243,N_10044);
nand U10623 (N_10623,N_9385,N_10181);
or U10624 (N_10624,N_10095,N_9470);
and U10625 (N_10625,N_10250,N_9823);
and U10626 (N_10626,N_10028,N_9513);
or U10627 (N_10627,N_9175,N_9670);
nand U10628 (N_10628,N_10093,N_9582);
nor U10629 (N_10629,N_9420,N_9220);
nor U10630 (N_10630,N_10251,N_9501);
and U10631 (N_10631,N_9124,N_10226);
nand U10632 (N_10632,N_10200,N_9593);
nand U10633 (N_10633,N_10341,N_9426);
or U10634 (N_10634,N_9841,N_9232);
nand U10635 (N_10635,N_9641,N_9685);
nor U10636 (N_10636,N_9065,N_9590);
nand U10637 (N_10637,N_9815,N_10112);
nand U10638 (N_10638,N_9231,N_9228);
nor U10639 (N_10639,N_9472,N_9672);
or U10640 (N_10640,N_10140,N_10268);
or U10641 (N_10641,N_10298,N_9006);
nor U10642 (N_10642,N_10280,N_9700);
nor U10643 (N_10643,N_9711,N_10358);
nand U10644 (N_10644,N_10259,N_9360);
or U10645 (N_10645,N_10348,N_9528);
nand U10646 (N_10646,N_9946,N_10378);
nand U10647 (N_10647,N_9729,N_9000);
nand U10648 (N_10648,N_9956,N_10049);
nor U10649 (N_10649,N_10009,N_10149);
nand U10650 (N_10650,N_9643,N_10027);
nor U10651 (N_10651,N_9052,N_10081);
and U10652 (N_10652,N_10077,N_10048);
nor U10653 (N_10653,N_9499,N_10486);
xor U10654 (N_10654,N_10420,N_10414);
or U10655 (N_10655,N_10072,N_9267);
xor U10656 (N_10656,N_9192,N_9876);
and U10657 (N_10657,N_9169,N_9566);
nand U10658 (N_10658,N_10202,N_9094);
nor U10659 (N_10659,N_10478,N_10395);
and U10660 (N_10660,N_9808,N_10155);
or U10661 (N_10661,N_9450,N_9419);
xor U10662 (N_10662,N_9900,N_10001);
or U10663 (N_10663,N_9068,N_9100);
nand U10664 (N_10664,N_9403,N_10228);
nor U10665 (N_10665,N_9026,N_10107);
nand U10666 (N_10666,N_10441,N_9942);
or U10667 (N_10667,N_10016,N_9421);
or U10668 (N_10668,N_9117,N_9965);
and U10669 (N_10669,N_10007,N_9769);
and U10670 (N_10670,N_9259,N_10389);
or U10671 (N_10671,N_9690,N_10248);
nand U10672 (N_10672,N_10234,N_10418);
and U10673 (N_10673,N_9960,N_9812);
xnor U10674 (N_10674,N_9929,N_9001);
and U10675 (N_10675,N_10139,N_10260);
nor U10676 (N_10676,N_9892,N_10467);
or U10677 (N_10677,N_10023,N_9085);
or U10678 (N_10678,N_9417,N_9396);
nor U10679 (N_10679,N_9933,N_9833);
nor U10680 (N_10680,N_10294,N_10387);
nor U10681 (N_10681,N_9324,N_9370);
nor U10682 (N_10682,N_9462,N_9821);
and U10683 (N_10683,N_10033,N_10305);
nor U10684 (N_10684,N_10308,N_10098);
and U10685 (N_10685,N_10422,N_9527);
nor U10686 (N_10686,N_9490,N_10452);
or U10687 (N_10687,N_10152,N_10085);
and U10688 (N_10688,N_9521,N_9377);
nand U10689 (N_10689,N_9138,N_10481);
nor U10690 (N_10690,N_10493,N_9982);
or U10691 (N_10691,N_9901,N_9121);
nor U10692 (N_10692,N_9936,N_10039);
nand U10693 (N_10693,N_9415,N_9801);
or U10694 (N_10694,N_9697,N_9557);
or U10695 (N_10695,N_9295,N_10491);
and U10696 (N_10696,N_9237,N_9612);
nor U10697 (N_10697,N_9977,N_9318);
xnor U10698 (N_10698,N_10360,N_10123);
nor U10699 (N_10699,N_9344,N_10122);
xor U10700 (N_10700,N_10425,N_9128);
nand U10701 (N_10701,N_9770,N_9195);
or U10702 (N_10702,N_9950,N_10293);
and U10703 (N_10703,N_9261,N_10357);
xor U10704 (N_10704,N_9277,N_9779);
and U10705 (N_10705,N_9283,N_9648);
or U10706 (N_10706,N_9718,N_9233);
and U10707 (N_10707,N_9477,N_9363);
or U10708 (N_10708,N_9329,N_10218);
nand U10709 (N_10709,N_9658,N_10235);
and U10710 (N_10710,N_9483,N_9142);
and U10711 (N_10711,N_9197,N_9102);
and U10712 (N_10712,N_9761,N_10430);
nand U10713 (N_10713,N_9251,N_9254);
nand U10714 (N_10714,N_9614,N_10003);
or U10715 (N_10715,N_9456,N_10326);
or U10716 (N_10716,N_10472,N_9202);
nand U10717 (N_10717,N_9630,N_10055);
xnor U10718 (N_10718,N_10008,N_10307);
xnor U10719 (N_10719,N_10192,N_10215);
and U10720 (N_10720,N_9906,N_9273);
and U10721 (N_10721,N_10329,N_10270);
or U10722 (N_10722,N_9114,N_9638);
and U10723 (N_10723,N_9015,N_9382);
xor U10724 (N_10724,N_10261,N_9923);
nor U10725 (N_10725,N_9112,N_9517);
xnor U10726 (N_10726,N_10459,N_9381);
and U10727 (N_10727,N_9298,N_9795);
nor U10728 (N_10728,N_9030,N_9176);
or U10729 (N_10729,N_9636,N_10128);
nand U10730 (N_10730,N_9887,N_10475);
and U10731 (N_10731,N_9384,N_9984);
nor U10732 (N_10732,N_9106,N_10454);
nand U10733 (N_10733,N_10015,N_9926);
or U10734 (N_10734,N_10020,N_10490);
nor U10735 (N_10735,N_9739,N_10242);
or U10736 (N_10736,N_9973,N_9720);
nor U10737 (N_10737,N_10300,N_9537);
and U10738 (N_10738,N_10427,N_9631);
and U10739 (N_10739,N_9869,N_9943);
xnor U10740 (N_10740,N_10017,N_10460);
nand U10741 (N_10741,N_9013,N_9628);
and U10742 (N_10742,N_9931,N_10245);
nor U10743 (N_10743,N_9749,N_10290);
nand U10744 (N_10744,N_10143,N_9023);
and U10745 (N_10745,N_10349,N_9511);
nor U10746 (N_10746,N_10340,N_10171);
or U10747 (N_10747,N_10332,N_10036);
or U10748 (N_10748,N_9241,N_9880);
xnor U10749 (N_10749,N_9181,N_9492);
or U10750 (N_10750,N_9358,N_9249);
and U10751 (N_10751,N_9692,N_9264);
or U10752 (N_10752,N_10492,N_9089);
xor U10753 (N_10753,N_9621,N_9240);
or U10754 (N_10754,N_9723,N_10180);
and U10755 (N_10755,N_9051,N_9830);
and U10756 (N_10756,N_9035,N_10090);
xor U10757 (N_10757,N_9014,N_10434);
nor U10758 (N_10758,N_9177,N_10322);
or U10759 (N_10759,N_9316,N_10439);
or U10760 (N_10760,N_9903,N_9713);
nand U10761 (N_10761,N_9562,N_10240);
nand U10762 (N_10762,N_9616,N_10083);
and U10763 (N_10763,N_10185,N_9584);
nor U10764 (N_10764,N_9019,N_9661);
and U10765 (N_10765,N_10070,N_9657);
or U10766 (N_10766,N_9971,N_9115);
xnor U10767 (N_10767,N_9063,N_9751);
nand U10768 (N_10768,N_9286,N_9482);
nand U10769 (N_10769,N_9730,N_9969);
and U10770 (N_10770,N_9340,N_9838);
nor U10771 (N_10771,N_9203,N_10415);
nor U10772 (N_10772,N_10056,N_9633);
and U10773 (N_10773,N_9620,N_9405);
nand U10774 (N_10774,N_10338,N_10121);
nand U10775 (N_10775,N_10224,N_10204);
xor U10776 (N_10776,N_9551,N_9605);
and U10777 (N_10777,N_10416,N_9409);
or U10778 (N_10778,N_9425,N_9596);
nor U10779 (N_10779,N_9875,N_9622);
and U10780 (N_10780,N_10227,N_9990);
nand U10781 (N_10781,N_9953,N_10161);
nand U10782 (N_10782,N_9904,N_9045);
and U10783 (N_10783,N_9759,N_9200);
or U10784 (N_10784,N_9367,N_10315);
and U10785 (N_10785,N_9122,N_9207);
or U10786 (N_10786,N_9217,N_10244);
nand U10787 (N_10787,N_9418,N_9054);
nand U10788 (N_10788,N_9315,N_9256);
nand U10789 (N_10789,N_10377,N_9864);
nand U10790 (N_10790,N_9012,N_10246);
or U10791 (N_10791,N_10409,N_10346);
nand U10792 (N_10792,N_9432,N_10262);
or U10793 (N_10793,N_9825,N_10206);
nor U10794 (N_10794,N_9414,N_10480);
or U10795 (N_10795,N_10067,N_9351);
nor U10796 (N_10796,N_10203,N_9828);
nor U10797 (N_10797,N_9884,N_9509);
nand U10798 (N_10798,N_9664,N_9074);
nor U10799 (N_10799,N_10396,N_10159);
nor U10800 (N_10800,N_10356,N_10099);
nor U10801 (N_10801,N_9569,N_9916);
nor U10802 (N_10802,N_9970,N_10238);
nor U10803 (N_10803,N_9947,N_9847);
or U10804 (N_10804,N_9629,N_9773);
or U10805 (N_10805,N_9091,N_9570);
nand U10806 (N_10806,N_10219,N_10097);
or U10807 (N_10807,N_10146,N_9033);
nor U10808 (N_10808,N_9060,N_10068);
xor U10809 (N_10809,N_9948,N_9281);
nand U10810 (N_10810,N_9905,N_9050);
and U10811 (N_10811,N_9558,N_9937);
or U10812 (N_10812,N_9625,N_10010);
nand U10813 (N_10813,N_9502,N_9149);
nor U10814 (N_10814,N_9009,N_9678);
nand U10815 (N_10815,N_10482,N_10113);
xor U10816 (N_10816,N_9250,N_9996);
or U10817 (N_10817,N_9481,N_9560);
or U10818 (N_10818,N_9182,N_9992);
nand U10819 (N_10819,N_9222,N_9252);
and U10820 (N_10820,N_10269,N_9007);
or U10821 (N_10821,N_9046,N_9959);
nand U10822 (N_10822,N_10476,N_9585);
nand U10823 (N_10823,N_10370,N_9066);
or U10824 (N_10824,N_9067,N_9446);
and U10825 (N_10825,N_9238,N_9780);
nand U10826 (N_10826,N_10074,N_9615);
and U10827 (N_10827,N_9205,N_10407);
nor U10828 (N_10828,N_10216,N_9811);
and U10829 (N_10829,N_9917,N_10164);
and U10830 (N_10830,N_9032,N_9921);
and U10831 (N_10831,N_9912,N_10144);
or U10832 (N_10832,N_10186,N_9423);
and U10833 (N_10833,N_9634,N_9236);
nor U10834 (N_10834,N_9886,N_9966);
or U10835 (N_10835,N_9728,N_10089);
nand U10836 (N_10836,N_10172,N_10317);
nor U10837 (N_10837,N_9888,N_9803);
nor U10838 (N_10838,N_10177,N_9209);
nand U10839 (N_10839,N_9784,N_9647);
nand U10840 (N_10840,N_9186,N_9938);
or U10841 (N_10841,N_10004,N_9741);
nand U10842 (N_10842,N_10384,N_9579);
nand U10843 (N_10843,N_9979,N_10276);
or U10844 (N_10844,N_9654,N_9465);
and U10845 (N_10845,N_9056,N_9300);
nor U10846 (N_10846,N_10222,N_10231);
nand U10847 (N_10847,N_9592,N_9433);
nor U10848 (N_10848,N_10062,N_10311);
and U10849 (N_10849,N_10133,N_9098);
nor U10850 (N_10850,N_9323,N_9101);
nand U10851 (N_10851,N_9599,N_10175);
and U10852 (N_10852,N_10385,N_10359);
nor U10853 (N_10853,N_9204,N_9524);
nor U10854 (N_10854,N_9424,N_10129);
nor U10855 (N_10855,N_9168,N_10025);
nor U10856 (N_10856,N_9504,N_9594);
or U10857 (N_10857,N_9734,N_9920);
and U10858 (N_10858,N_9167,N_10479);
and U10859 (N_10859,N_9216,N_9305);
or U10860 (N_10860,N_9258,N_9174);
xor U10861 (N_10861,N_9716,N_10499);
and U10862 (N_10862,N_9133,N_10189);
nor U10863 (N_10863,N_9364,N_10103);
xnor U10864 (N_10864,N_9047,N_9954);
nor U10865 (N_10865,N_10254,N_9696);
and U10866 (N_10866,N_9348,N_9406);
or U10867 (N_10867,N_10145,N_10134);
or U10868 (N_10868,N_10006,N_9473);
xnor U10869 (N_10869,N_9764,N_9279);
or U10870 (N_10870,N_10431,N_10368);
nand U10871 (N_10871,N_9952,N_10432);
nand U10872 (N_10872,N_9548,N_10013);
or U10873 (N_10873,N_9763,N_10108);
and U10874 (N_10874,N_10465,N_9388);
and U10875 (N_10875,N_9055,N_9379);
and U10876 (N_10876,N_9336,N_10188);
nand U10877 (N_10877,N_10309,N_10328);
or U10878 (N_10878,N_9188,N_9915);
nand U10879 (N_10879,N_9666,N_9872);
or U10880 (N_10880,N_9479,N_9891);
nor U10881 (N_10881,N_9507,N_9577);
xor U10882 (N_10882,N_9373,N_10265);
or U10883 (N_10883,N_9302,N_9113);
and U10884 (N_10884,N_9735,N_9345);
nor U10885 (N_10885,N_10498,N_10024);
nand U10886 (N_10886,N_9044,N_9438);
nor U10887 (N_10887,N_9039,N_9285);
nor U10888 (N_10888,N_10058,N_9156);
nor U10889 (N_10889,N_9556,N_9376);
nor U10890 (N_10890,N_9907,N_10154);
and U10891 (N_10891,N_9136,N_10263);
and U10892 (N_10892,N_10195,N_9568);
xnor U10893 (N_10893,N_10196,N_9873);
or U10894 (N_10894,N_10495,N_9341);
or U10895 (N_10895,N_9389,N_9194);
nand U10896 (N_10896,N_10247,N_10063);
or U10897 (N_10897,N_10080,N_9087);
or U10898 (N_10898,N_9107,N_9164);
xnor U10899 (N_10899,N_9410,N_9260);
nor U10900 (N_10900,N_9299,N_10158);
and U10901 (N_10901,N_9284,N_9191);
and U10902 (N_10902,N_10367,N_9062);
nand U10903 (N_10903,N_10485,N_9624);
nand U10904 (N_10904,N_9722,N_9366);
nand U10905 (N_10905,N_9994,N_9523);
nor U10906 (N_10906,N_9190,N_9311);
xor U10907 (N_10907,N_9986,N_10316);
or U10908 (N_10908,N_9707,N_10365);
nand U10909 (N_10909,N_10302,N_9682);
nand U10910 (N_10910,N_9036,N_9386);
nand U10911 (N_10911,N_9269,N_10423);
xnor U10912 (N_10912,N_9048,N_9399);
or U10913 (N_10913,N_9846,N_9372);
nor U10914 (N_10914,N_9505,N_9064);
nor U10915 (N_10915,N_9813,N_10391);
nor U10916 (N_10916,N_10253,N_9027);
xnor U10917 (N_10917,N_10497,N_9725);
nor U10918 (N_10918,N_9245,N_10069);
and U10919 (N_10919,N_9212,N_9387);
or U10920 (N_10920,N_10116,N_9096);
and U10921 (N_10921,N_10464,N_10225);
xor U10922 (N_10922,N_10320,N_10076);
nand U10923 (N_10923,N_10343,N_10102);
nor U10924 (N_10924,N_9093,N_9162);
or U10925 (N_10925,N_9715,N_9867);
or U10926 (N_10926,N_9354,N_9980);
and U10927 (N_10927,N_9290,N_10400);
or U10928 (N_10928,N_10401,N_9488);
xnor U10929 (N_10929,N_9893,N_9427);
and U10930 (N_10930,N_9645,N_9724);
nand U10931 (N_10931,N_9908,N_9229);
or U10932 (N_10932,N_9783,N_9934);
nor U10933 (N_10933,N_9053,N_10364);
or U10934 (N_10934,N_9475,N_10106);
xnor U10935 (N_10935,N_9173,N_9148);
nand U10936 (N_10936,N_10162,N_10406);
or U10937 (N_10937,N_9180,N_9208);
xor U10938 (N_10938,N_9701,N_9317);
nand U10939 (N_10939,N_9355,N_9708);
and U10940 (N_10940,N_9226,N_9144);
nand U10941 (N_10941,N_10433,N_9147);
nand U10942 (N_10942,N_10092,N_9330);
or U10943 (N_10943,N_9827,N_9108);
or U10944 (N_10944,N_9371,N_9400);
and U10945 (N_10945,N_9293,N_9964);
or U10946 (N_10946,N_10117,N_9581);
or U10947 (N_10947,N_10279,N_9829);
xnor U10948 (N_10948,N_9227,N_9911);
or U10949 (N_10949,N_9754,N_9602);
and U10950 (N_10950,N_9662,N_9003);
nor U10951 (N_10951,N_9031,N_10413);
or U10952 (N_10952,N_9842,N_10374);
and U10953 (N_10953,N_9163,N_10043);
or U10954 (N_10954,N_9798,N_9782);
xnor U10955 (N_10955,N_9151,N_10319);
nand U10956 (N_10956,N_9681,N_10484);
and U10957 (N_10957,N_10289,N_10419);
nor U10958 (N_10958,N_9991,N_10052);
or U10959 (N_10959,N_9404,N_9913);
nor U10960 (N_10960,N_9896,N_9265);
or U10961 (N_10961,N_9266,N_9453);
xnor U10962 (N_10962,N_10239,N_9246);
nand U10963 (N_10963,N_9766,N_9213);
nand U10964 (N_10964,N_9278,N_10035);
and U10965 (N_10965,N_9609,N_9183);
or U10966 (N_10966,N_10053,N_10148);
xnor U10967 (N_10967,N_9613,N_10337);
nor U10968 (N_10968,N_9727,N_9119);
nor U10969 (N_10969,N_10211,N_9339);
nor U10970 (N_10970,N_9485,N_10029);
or U10971 (N_10971,N_10487,N_9476);
nor U10972 (N_10972,N_10379,N_9271);
nand U10973 (N_10973,N_9851,N_10135);
or U10974 (N_10974,N_9171,N_9794);
nor U10975 (N_10975,N_10169,N_9120);
nor U10976 (N_10976,N_9326,N_9985);
or U10977 (N_10977,N_10002,N_9649);
and U10978 (N_10978,N_9274,N_10429);
xor U10979 (N_10979,N_9814,N_9165);
and U10980 (N_10980,N_10115,N_10241);
nand U10981 (N_10981,N_10426,N_10369);
nand U10982 (N_10982,N_10404,N_9058);
nand U10983 (N_10983,N_9038,N_10440);
and U10984 (N_10984,N_9333,N_10174);
xnor U10985 (N_10985,N_9002,N_9059);
nor U10986 (N_10986,N_9758,N_9242);
and U10987 (N_10987,N_9487,N_10453);
nand U10988 (N_10988,N_9402,N_9976);
xor U10989 (N_10989,N_10272,N_9750);
or U10990 (N_10990,N_10277,N_9478);
and U10991 (N_10991,N_10477,N_9069);
or U10992 (N_10992,N_9184,N_10127);
nor U10993 (N_10993,N_9894,N_10182);
and U10994 (N_10994,N_9853,N_9210);
or U10995 (N_10995,N_9451,N_9455);
and U10996 (N_10996,N_10283,N_10167);
and U10997 (N_10997,N_9500,N_9790);
and U10998 (N_10998,N_9611,N_9755);
nand U10999 (N_10999,N_9576,N_9591);
or U11000 (N_11000,N_9951,N_9844);
or U11001 (N_11001,N_9665,N_9319);
or U11002 (N_11002,N_10232,N_10339);
and U11003 (N_11003,N_9125,N_9436);
nor U11004 (N_11004,N_9679,N_9206);
or U11005 (N_11005,N_10021,N_9775);
nor U11006 (N_11006,N_9443,N_9070);
and U11007 (N_11007,N_9706,N_9819);
nor U11008 (N_11008,N_9255,N_10394);
xor U11009 (N_11009,N_9496,N_10207);
nand U11010 (N_11010,N_9663,N_9603);
and U11011 (N_11011,N_9467,N_9158);
or U11012 (N_11012,N_9253,N_9944);
nand U11013 (N_11013,N_9118,N_10096);
nor U11014 (N_11014,N_9154,N_9322);
or U11015 (N_11015,N_10405,N_10136);
nand U11016 (N_11016,N_10412,N_9320);
nor U11017 (N_11017,N_9332,N_9767);
nand U11018 (N_11018,N_9025,N_10458);
and U11019 (N_11019,N_9695,N_9752);
nand U11020 (N_11020,N_10296,N_9306);
nor U11021 (N_11021,N_9738,N_9494);
xor U11022 (N_11022,N_9099,N_9092);
and U11023 (N_11023,N_9545,N_9328);
or U11024 (N_11024,N_10050,N_10079);
or U11025 (N_11025,N_9471,N_9732);
nand U11026 (N_11026,N_9449,N_9411);
nand U11027 (N_11027,N_9549,N_10073);
or U11028 (N_11028,N_9506,N_9837);
or U11029 (N_11029,N_9349,N_10451);
or U11030 (N_11030,N_9368,N_10091);
or U11031 (N_11031,N_9081,N_10267);
nand U11032 (N_11032,N_10411,N_9157);
and U11033 (N_11033,N_9442,N_9538);
nor U11034 (N_11034,N_9314,N_10299);
and U11035 (N_11035,N_10295,N_9949);
nand U11036 (N_11036,N_9651,N_10038);
nor U11037 (N_11037,N_9460,N_10301);
nand U11038 (N_11038,N_9301,N_9441);
and U11039 (N_11039,N_9882,N_10399);
nor U11040 (N_11040,N_9225,N_9080);
xnor U11041 (N_11041,N_9362,N_9532);
or U11042 (N_11042,N_10304,N_9428);
or U11043 (N_11043,N_9733,N_9586);
nand U11044 (N_11044,N_9753,N_9796);
nand U11045 (N_11045,N_9785,N_9924);
or U11046 (N_11046,N_9632,N_9902);
nor U11047 (N_11047,N_10266,N_10461);
nor U11048 (N_11048,N_9604,N_10282);
xnor U11049 (N_11049,N_9910,N_9588);
nand U11050 (N_11050,N_9365,N_9957);
xor U11051 (N_11051,N_10138,N_9868);
nor U11052 (N_11052,N_9288,N_9575);
nand U11053 (N_11053,N_9486,N_10436);
xnor U11054 (N_11054,N_9135,N_10352);
and U11055 (N_11055,N_9852,N_9395);
nand U11056 (N_11056,N_10408,N_9352);
and U11057 (N_11057,N_10284,N_10022);
nor U11058 (N_11058,N_9607,N_9617);
and U11059 (N_11059,N_10187,N_10183);
or U11060 (N_11060,N_9170,N_9595);
or U11061 (N_11061,N_9214,N_9383);
xnor U11062 (N_11062,N_9004,N_9580);
nand U11063 (N_11063,N_9744,N_10330);
or U11064 (N_11064,N_10168,N_9608);
nor U11065 (N_11065,N_9498,N_10447);
nor U11066 (N_11066,N_10210,N_9082);
or U11067 (N_11067,N_10449,N_9211);
and U11068 (N_11068,N_10258,N_9571);
nor U11069 (N_11069,N_9215,N_9786);
and U11070 (N_11070,N_9457,N_9199);
and U11071 (N_11071,N_10179,N_10229);
xnor U11072 (N_11072,N_9745,N_9930);
nand U11073 (N_11073,N_9573,N_9635);
nand U11074 (N_11074,N_10291,N_10173);
and U11075 (N_11075,N_10444,N_10456);
and U11076 (N_11076,N_10157,N_9793);
nor U11077 (N_11077,N_9963,N_9198);
nand U11078 (N_11078,N_9407,N_10132);
or U11079 (N_11079,N_9110,N_9430);
nand U11080 (N_11080,N_10463,N_10264);
xnor U11081 (N_11081,N_9644,N_9011);
xnor U11082 (N_11082,N_10120,N_9380);
and U11083 (N_11083,N_10323,N_9429);
or U11084 (N_11084,N_9334,N_9495);
or U11085 (N_11085,N_10397,N_10435);
nand U11086 (N_11086,N_9743,N_9223);
and U11087 (N_11087,N_9461,N_9731);
nor U11088 (N_11088,N_10209,N_9234);
nor U11089 (N_11089,N_9932,N_9639);
nor U11090 (N_11090,N_9895,N_9854);
and U11091 (N_11091,N_9987,N_10184);
or U11092 (N_11092,N_9129,N_9889);
nand U11093 (N_11093,N_9760,N_9564);
nand U11094 (N_11094,N_9469,N_9143);
and U11095 (N_11095,N_10366,N_9768);
nor U11096 (N_11096,N_9282,N_9071);
and U11097 (N_11097,N_10124,N_9589);
or U11098 (N_11098,N_10214,N_10061);
and U11099 (N_11099,N_9655,N_9159);
nor U11100 (N_11100,N_9193,N_9870);
or U11101 (N_11101,N_9653,N_9034);
and U11102 (N_11102,N_9777,N_9694);
xnor U11103 (N_11103,N_10194,N_9981);
nand U11104 (N_11104,N_9493,N_9550);
nand U11105 (N_11105,N_10288,N_9397);
or U11106 (N_11106,N_9878,N_9774);
nor U11107 (N_11107,N_9024,N_10450);
nor U11108 (N_11108,N_9789,N_9525);
nand U11109 (N_11109,N_9392,N_9437);
or U11110 (N_11110,N_10354,N_9704);
and U11111 (N_11111,N_10088,N_9598);
nor U11112 (N_11112,N_10170,N_9497);
and U11113 (N_11113,N_9817,N_9877);
nand U11114 (N_11114,N_10327,N_9041);
or U11115 (N_11115,N_9879,N_10496);
nand U11116 (N_11116,N_9572,N_9583);
and U11117 (N_11117,N_9776,N_9927);
and U11118 (N_11118,N_9650,N_10040);
or U11119 (N_11119,N_9757,N_9544);
nand U11120 (N_11120,N_9762,N_9531);
nand U11121 (N_11121,N_10141,N_9998);
and U11122 (N_11122,N_9565,N_9652);
nand U11123 (N_11123,N_9684,N_9459);
or U11124 (N_11124,N_9547,N_9555);
nand U11125 (N_11125,N_9463,N_9721);
nor U11126 (N_11126,N_10468,N_9219);
nand U11127 (N_11127,N_9978,N_10361);
and U11128 (N_11128,N_9918,N_9218);
nor U11129 (N_11129,N_9610,N_9037);
or U11130 (N_11130,N_9268,N_9086);
xor U11131 (N_11131,N_9073,N_9291);
nor U11132 (N_11132,N_9542,N_10150);
nand U11133 (N_11133,N_9413,N_9809);
nor U11134 (N_11134,N_10230,N_10125);
nor U11135 (N_11135,N_9861,N_9850);
or U11136 (N_11136,N_9116,N_10355);
or U11137 (N_11137,N_10243,N_10278);
xnor U11138 (N_11138,N_9503,N_9029);
or U11139 (N_11139,N_9712,N_10160);
nand U11140 (N_11140,N_9431,N_9224);
and U11141 (N_11141,N_9818,N_10178);
nor U11142 (N_11142,N_10163,N_10030);
or U11143 (N_11143,N_10166,N_9356);
and U11144 (N_11144,N_9448,N_10156);
nor U11145 (N_11145,N_10084,N_9103);
or U11146 (N_11146,N_9408,N_9726);
nor U11147 (N_11147,N_10118,N_9079);
nand U11148 (N_11148,N_9637,N_10147);
and U11149 (N_11149,N_9139,N_9719);
xor U11150 (N_11150,N_9464,N_10014);
xor U11151 (N_11151,N_9689,N_10489);
and U11152 (N_11152,N_9307,N_10109);
nor U11153 (N_11153,N_9017,N_9881);
or U11154 (N_11154,N_10018,N_9454);
nand U11155 (N_11155,N_9155,N_9049);
nand U11156 (N_11156,N_9554,N_10217);
nor U11157 (N_11157,N_9416,N_9280);
and U11158 (N_11158,N_9297,N_9802);
and U11159 (N_11159,N_10041,N_9659);
or U11160 (N_11160,N_9126,N_9533);
xor U11161 (N_11161,N_10362,N_9152);
nor U11162 (N_11162,N_9958,N_9997);
nor U11163 (N_11163,N_9083,N_10333);
nor U11164 (N_11164,N_10101,N_9799);
xnor U11165 (N_11165,N_9508,N_9717);
and U11166 (N_11166,N_9179,N_9412);
or U11167 (N_11167,N_9350,N_9321);
nand U11168 (N_11168,N_10075,N_9008);
and U11169 (N_11169,N_10386,N_9519);
xor U11170 (N_11170,N_10064,N_9541);
nor U11171 (N_11171,N_9561,N_9816);
and U11172 (N_11172,N_10392,N_10344);
nand U11173 (N_11173,N_9072,N_10045);
nand U11174 (N_11174,N_10031,N_9422);
and U11175 (N_11175,N_9440,N_9132);
and U11176 (N_11176,N_10318,N_10111);
nor U11177 (N_11177,N_10488,N_9899);
nor U11178 (N_11178,N_9874,N_9686);
nand U11179 (N_11179,N_10071,N_10457);
and U11180 (N_11180,N_9325,N_10462);
or U11181 (N_11181,N_9434,N_9771);
xor U11182 (N_11182,N_9076,N_9378);
and U11183 (N_11183,N_9995,N_9822);
nand U11184 (N_11184,N_10190,N_10176);
nor U11185 (N_11185,N_9688,N_9865);
or U11186 (N_11186,N_10353,N_9552);
and U11187 (N_11187,N_10078,N_9871);
nand U11188 (N_11188,N_9962,N_9597);
nor U11189 (N_11189,N_9941,N_9674);
or U11190 (N_11190,N_9928,N_9691);
and U11191 (N_11191,N_10428,N_9668);
nand U11192 (N_11192,N_9393,N_10381);
xor U11193 (N_11193,N_9491,N_9338);
nor U11194 (N_11194,N_9646,N_10037);
and U11195 (N_11195,N_10131,N_9309);
and U11196 (N_11196,N_9993,N_10051);
nand U11197 (N_11197,N_9042,N_9810);
or U11198 (N_11198,N_9740,N_9020);
and U11199 (N_11199,N_9145,N_10382);
nor U11200 (N_11200,N_10130,N_10324);
and U11201 (N_11201,N_9559,N_9335);
or U11202 (N_11202,N_10114,N_9703);
nor U11203 (N_11203,N_9939,N_10100);
nand U11204 (N_11204,N_9018,N_9458);
nand U11205 (N_11205,N_10257,N_10437);
and U11206 (N_11206,N_9095,N_9866);
and U11207 (N_11207,N_9518,N_9835);
or U11208 (N_11208,N_10274,N_9673);
and U11209 (N_11209,N_9390,N_9296);
or U11210 (N_11210,N_10398,N_9516);
nor U11211 (N_11211,N_9539,N_9845);
nand U11212 (N_11212,N_9627,N_10087);
nor U11213 (N_11213,N_9141,N_10275);
nand U11214 (N_11214,N_9687,N_10197);
nand U11215 (N_11215,N_9303,N_9040);
nand U11216 (N_11216,N_10347,N_9445);
nor U11217 (N_11217,N_9078,N_9150);
nor U11218 (N_11218,N_9526,N_9452);
or U11219 (N_11219,N_9680,N_9474);
nor U11220 (N_11220,N_9510,N_9676);
or U11221 (N_11221,N_10390,N_9005);
and U11222 (N_11222,N_9897,N_9922);
and U11223 (N_11223,N_9945,N_10483);
and U11224 (N_11224,N_9153,N_9806);
xor U11225 (N_11225,N_9974,N_10005);
or U11226 (N_11226,N_10233,N_10442);
xor U11227 (N_11227,N_9972,N_9097);
nand U11228 (N_11228,N_10249,N_10221);
nor U11229 (N_11229,N_10303,N_9447);
nand U11230 (N_11230,N_9466,N_9988);
nor U11231 (N_11231,N_10402,N_9484);
and U11232 (N_11232,N_10331,N_10334);
nand U11233 (N_11233,N_9104,N_9914);
nand U11234 (N_11234,N_10336,N_10199);
or U11235 (N_11235,N_9189,N_10448);
nor U11236 (N_11236,N_9289,N_9435);
xor U11237 (N_11237,N_9709,N_9010);
or U11238 (N_11238,N_10494,N_10059);
nand U11239 (N_11239,N_9359,N_9606);
nand U11240 (N_11240,N_9792,N_9369);
and U11241 (N_11241,N_9862,N_9563);
xor U11242 (N_11242,N_9800,N_9698);
nor U11243 (N_11243,N_9263,N_9374);
nand U11244 (N_11244,N_10256,N_9346);
or U11245 (N_11245,N_9043,N_9858);
and U11246 (N_11246,N_9391,N_10082);
or U11247 (N_11247,N_9820,N_9166);
nand U11248 (N_11248,N_9077,N_9111);
nand U11249 (N_11249,N_10271,N_9276);
nor U11250 (N_11250,N_9740,N_10113);
or U11251 (N_11251,N_10330,N_10010);
nand U11252 (N_11252,N_9062,N_10411);
nand U11253 (N_11253,N_9476,N_10130);
nand U11254 (N_11254,N_9338,N_9221);
or U11255 (N_11255,N_10057,N_10165);
nand U11256 (N_11256,N_9143,N_9249);
or U11257 (N_11257,N_9986,N_9003);
or U11258 (N_11258,N_9444,N_9072);
nand U11259 (N_11259,N_10205,N_9113);
nand U11260 (N_11260,N_9821,N_10298);
or U11261 (N_11261,N_9840,N_9127);
and U11262 (N_11262,N_9646,N_10422);
or U11263 (N_11263,N_9078,N_9066);
nand U11264 (N_11264,N_10280,N_9735);
nand U11265 (N_11265,N_10452,N_10308);
and U11266 (N_11266,N_9660,N_9130);
and U11267 (N_11267,N_10180,N_9254);
nor U11268 (N_11268,N_9891,N_9642);
xor U11269 (N_11269,N_9913,N_9807);
nand U11270 (N_11270,N_9753,N_9350);
xnor U11271 (N_11271,N_9774,N_9847);
nor U11272 (N_11272,N_10005,N_9098);
nand U11273 (N_11273,N_9115,N_10020);
nand U11274 (N_11274,N_10098,N_10348);
and U11275 (N_11275,N_10360,N_9699);
or U11276 (N_11276,N_9759,N_9365);
or U11277 (N_11277,N_10365,N_9989);
nor U11278 (N_11278,N_10252,N_9358);
or U11279 (N_11279,N_9002,N_10210);
and U11280 (N_11280,N_10411,N_10485);
or U11281 (N_11281,N_9113,N_10079);
and U11282 (N_11282,N_10336,N_10032);
xnor U11283 (N_11283,N_9415,N_10000);
xnor U11284 (N_11284,N_10497,N_9515);
nand U11285 (N_11285,N_9883,N_10417);
or U11286 (N_11286,N_10397,N_9000);
nor U11287 (N_11287,N_9599,N_10185);
or U11288 (N_11288,N_9971,N_10111);
and U11289 (N_11289,N_9417,N_9681);
nor U11290 (N_11290,N_10092,N_9322);
or U11291 (N_11291,N_10422,N_9044);
and U11292 (N_11292,N_10140,N_9233);
or U11293 (N_11293,N_9439,N_9015);
nor U11294 (N_11294,N_9446,N_10211);
xor U11295 (N_11295,N_9709,N_10443);
nand U11296 (N_11296,N_9431,N_9433);
nand U11297 (N_11297,N_9949,N_9145);
or U11298 (N_11298,N_9078,N_9002);
or U11299 (N_11299,N_9907,N_10492);
nor U11300 (N_11300,N_10226,N_10375);
and U11301 (N_11301,N_9253,N_10459);
and U11302 (N_11302,N_10498,N_9475);
nor U11303 (N_11303,N_9442,N_9217);
nand U11304 (N_11304,N_9256,N_9287);
nand U11305 (N_11305,N_9603,N_10383);
and U11306 (N_11306,N_9653,N_9350);
nand U11307 (N_11307,N_9307,N_9070);
or U11308 (N_11308,N_9205,N_9014);
or U11309 (N_11309,N_9199,N_9782);
nand U11310 (N_11310,N_9871,N_9731);
and U11311 (N_11311,N_9749,N_9149);
nor U11312 (N_11312,N_9200,N_10182);
nand U11313 (N_11313,N_9178,N_9193);
nor U11314 (N_11314,N_9933,N_9942);
nand U11315 (N_11315,N_9833,N_9323);
nor U11316 (N_11316,N_9994,N_9751);
and U11317 (N_11317,N_10154,N_9094);
nand U11318 (N_11318,N_9441,N_9629);
nand U11319 (N_11319,N_9435,N_10347);
or U11320 (N_11320,N_9456,N_9812);
and U11321 (N_11321,N_9829,N_9806);
or U11322 (N_11322,N_9822,N_9806);
xnor U11323 (N_11323,N_9652,N_9182);
nor U11324 (N_11324,N_9385,N_9554);
nor U11325 (N_11325,N_10425,N_10016);
nor U11326 (N_11326,N_9901,N_9290);
nand U11327 (N_11327,N_10059,N_9781);
nand U11328 (N_11328,N_9889,N_9229);
and U11329 (N_11329,N_10221,N_9882);
xnor U11330 (N_11330,N_9779,N_9466);
or U11331 (N_11331,N_9177,N_9073);
xnor U11332 (N_11332,N_9591,N_9113);
and U11333 (N_11333,N_10448,N_9712);
and U11334 (N_11334,N_10345,N_9970);
nor U11335 (N_11335,N_9385,N_9574);
or U11336 (N_11336,N_10324,N_9006);
nand U11337 (N_11337,N_10395,N_10442);
nand U11338 (N_11338,N_9894,N_9443);
or U11339 (N_11339,N_9164,N_10368);
nand U11340 (N_11340,N_10492,N_9173);
nand U11341 (N_11341,N_10477,N_9480);
nand U11342 (N_11342,N_9037,N_9590);
or U11343 (N_11343,N_9870,N_9230);
xnor U11344 (N_11344,N_9898,N_9405);
xor U11345 (N_11345,N_9859,N_9385);
or U11346 (N_11346,N_10414,N_9030);
and U11347 (N_11347,N_9030,N_9837);
nand U11348 (N_11348,N_10109,N_10021);
and U11349 (N_11349,N_10178,N_9026);
nor U11350 (N_11350,N_9129,N_9926);
xnor U11351 (N_11351,N_10254,N_9088);
or U11352 (N_11352,N_10267,N_9415);
and U11353 (N_11353,N_9950,N_10366);
nand U11354 (N_11354,N_9963,N_9699);
xnor U11355 (N_11355,N_9159,N_9107);
and U11356 (N_11356,N_9602,N_10244);
nand U11357 (N_11357,N_9047,N_9555);
or U11358 (N_11358,N_10239,N_10188);
and U11359 (N_11359,N_9885,N_10020);
or U11360 (N_11360,N_10130,N_9420);
xor U11361 (N_11361,N_9873,N_9518);
or U11362 (N_11362,N_9998,N_9679);
and U11363 (N_11363,N_10341,N_9929);
and U11364 (N_11364,N_9038,N_9863);
or U11365 (N_11365,N_10438,N_10204);
nand U11366 (N_11366,N_9548,N_9219);
nor U11367 (N_11367,N_10131,N_10192);
nor U11368 (N_11368,N_9916,N_9622);
and U11369 (N_11369,N_9603,N_9455);
nand U11370 (N_11370,N_10345,N_9559);
xnor U11371 (N_11371,N_10068,N_10169);
nor U11372 (N_11372,N_9422,N_10095);
or U11373 (N_11373,N_9422,N_9711);
and U11374 (N_11374,N_9016,N_9660);
or U11375 (N_11375,N_9631,N_10169);
and U11376 (N_11376,N_9005,N_10099);
and U11377 (N_11377,N_10198,N_9972);
xor U11378 (N_11378,N_10361,N_9982);
and U11379 (N_11379,N_9305,N_10431);
and U11380 (N_11380,N_9722,N_10174);
nor U11381 (N_11381,N_10197,N_9457);
and U11382 (N_11382,N_10035,N_9502);
and U11383 (N_11383,N_9151,N_9507);
and U11384 (N_11384,N_9557,N_9635);
and U11385 (N_11385,N_9028,N_9313);
and U11386 (N_11386,N_9565,N_10214);
nand U11387 (N_11387,N_9958,N_9208);
and U11388 (N_11388,N_9729,N_10265);
nor U11389 (N_11389,N_9742,N_9469);
xor U11390 (N_11390,N_10489,N_9507);
or U11391 (N_11391,N_9416,N_9502);
or U11392 (N_11392,N_10403,N_9849);
or U11393 (N_11393,N_10454,N_9280);
nor U11394 (N_11394,N_9273,N_9592);
or U11395 (N_11395,N_10153,N_10275);
and U11396 (N_11396,N_10038,N_10293);
and U11397 (N_11397,N_10006,N_9684);
and U11398 (N_11398,N_9753,N_9930);
or U11399 (N_11399,N_9546,N_9133);
or U11400 (N_11400,N_9754,N_9984);
nor U11401 (N_11401,N_9097,N_9978);
nand U11402 (N_11402,N_10108,N_9382);
nand U11403 (N_11403,N_9635,N_10480);
or U11404 (N_11404,N_9546,N_9668);
or U11405 (N_11405,N_9919,N_10317);
and U11406 (N_11406,N_10288,N_10307);
nand U11407 (N_11407,N_9675,N_9924);
and U11408 (N_11408,N_9463,N_9974);
and U11409 (N_11409,N_10163,N_10239);
or U11410 (N_11410,N_9715,N_9180);
xnor U11411 (N_11411,N_9166,N_9767);
and U11412 (N_11412,N_9052,N_9354);
or U11413 (N_11413,N_10414,N_9560);
nor U11414 (N_11414,N_10023,N_9368);
nand U11415 (N_11415,N_9076,N_10383);
nand U11416 (N_11416,N_10262,N_9909);
or U11417 (N_11417,N_9352,N_10033);
nor U11418 (N_11418,N_9615,N_10204);
nand U11419 (N_11419,N_9515,N_10390);
xor U11420 (N_11420,N_9446,N_9719);
nor U11421 (N_11421,N_9614,N_9932);
or U11422 (N_11422,N_10447,N_9633);
nand U11423 (N_11423,N_9967,N_9933);
xor U11424 (N_11424,N_10055,N_9308);
or U11425 (N_11425,N_9726,N_9310);
or U11426 (N_11426,N_10202,N_9025);
nand U11427 (N_11427,N_9751,N_9641);
and U11428 (N_11428,N_9732,N_9131);
and U11429 (N_11429,N_9173,N_9042);
nand U11430 (N_11430,N_10134,N_10236);
xnor U11431 (N_11431,N_9470,N_9742);
or U11432 (N_11432,N_9539,N_9384);
nor U11433 (N_11433,N_9774,N_9337);
or U11434 (N_11434,N_9082,N_9376);
nor U11435 (N_11435,N_9731,N_9446);
nand U11436 (N_11436,N_10055,N_9634);
and U11437 (N_11437,N_10375,N_9310);
xnor U11438 (N_11438,N_9800,N_9500);
or U11439 (N_11439,N_9212,N_9082);
or U11440 (N_11440,N_9857,N_10158);
or U11441 (N_11441,N_9037,N_9313);
nor U11442 (N_11442,N_9856,N_9624);
xnor U11443 (N_11443,N_10474,N_9230);
and U11444 (N_11444,N_10134,N_9091);
and U11445 (N_11445,N_9409,N_10469);
or U11446 (N_11446,N_9097,N_9676);
nor U11447 (N_11447,N_10251,N_9506);
nand U11448 (N_11448,N_9814,N_9269);
or U11449 (N_11449,N_9341,N_9786);
nand U11450 (N_11450,N_10138,N_9858);
nor U11451 (N_11451,N_10317,N_9589);
nor U11452 (N_11452,N_10243,N_9415);
nor U11453 (N_11453,N_10457,N_9459);
xor U11454 (N_11454,N_9617,N_9866);
or U11455 (N_11455,N_10007,N_9689);
nor U11456 (N_11456,N_9801,N_9988);
nor U11457 (N_11457,N_9714,N_9171);
xnor U11458 (N_11458,N_10448,N_9208);
or U11459 (N_11459,N_9107,N_9408);
or U11460 (N_11460,N_9798,N_9671);
xnor U11461 (N_11461,N_9016,N_10356);
or U11462 (N_11462,N_10470,N_10298);
nand U11463 (N_11463,N_9256,N_9810);
or U11464 (N_11464,N_9452,N_10155);
nor U11465 (N_11465,N_9261,N_9212);
nand U11466 (N_11466,N_9415,N_9772);
xnor U11467 (N_11467,N_9417,N_9628);
nand U11468 (N_11468,N_9847,N_9745);
or U11469 (N_11469,N_9330,N_9228);
and U11470 (N_11470,N_9391,N_9326);
and U11471 (N_11471,N_9215,N_9974);
nand U11472 (N_11472,N_9102,N_9317);
and U11473 (N_11473,N_9518,N_9235);
xnor U11474 (N_11474,N_10458,N_9754);
and U11475 (N_11475,N_9225,N_9056);
nand U11476 (N_11476,N_10442,N_9393);
nand U11477 (N_11477,N_9733,N_9318);
and U11478 (N_11478,N_10384,N_9892);
or U11479 (N_11479,N_9377,N_9940);
and U11480 (N_11480,N_9587,N_9064);
nand U11481 (N_11481,N_9785,N_9546);
or U11482 (N_11482,N_9524,N_10137);
nor U11483 (N_11483,N_10194,N_9565);
or U11484 (N_11484,N_9973,N_9065);
nor U11485 (N_11485,N_9943,N_10327);
and U11486 (N_11486,N_9259,N_9522);
nand U11487 (N_11487,N_9979,N_9758);
nand U11488 (N_11488,N_10146,N_10480);
or U11489 (N_11489,N_9843,N_9425);
nor U11490 (N_11490,N_9580,N_9919);
or U11491 (N_11491,N_9127,N_9443);
nor U11492 (N_11492,N_9041,N_9635);
and U11493 (N_11493,N_9280,N_9182);
and U11494 (N_11494,N_10422,N_9227);
or U11495 (N_11495,N_10475,N_9533);
nand U11496 (N_11496,N_10102,N_9190);
and U11497 (N_11497,N_10136,N_10209);
or U11498 (N_11498,N_9636,N_9028);
xor U11499 (N_11499,N_9693,N_9185);
or U11500 (N_11500,N_9784,N_10173);
nor U11501 (N_11501,N_9303,N_10099);
and U11502 (N_11502,N_10464,N_10473);
or U11503 (N_11503,N_10108,N_9798);
nand U11504 (N_11504,N_9006,N_9328);
or U11505 (N_11505,N_10251,N_9465);
and U11506 (N_11506,N_10244,N_9964);
xnor U11507 (N_11507,N_9946,N_9403);
nand U11508 (N_11508,N_9129,N_9731);
nor U11509 (N_11509,N_9269,N_10362);
or U11510 (N_11510,N_9041,N_9528);
and U11511 (N_11511,N_10213,N_10185);
and U11512 (N_11512,N_9689,N_9919);
nand U11513 (N_11513,N_9023,N_10017);
xnor U11514 (N_11514,N_10334,N_10088);
or U11515 (N_11515,N_10147,N_9552);
and U11516 (N_11516,N_9821,N_9857);
xnor U11517 (N_11517,N_9618,N_9542);
or U11518 (N_11518,N_9822,N_10126);
nand U11519 (N_11519,N_9039,N_9542);
nor U11520 (N_11520,N_9944,N_9177);
nand U11521 (N_11521,N_10252,N_9898);
nor U11522 (N_11522,N_9683,N_10420);
nor U11523 (N_11523,N_9299,N_10053);
nand U11524 (N_11524,N_10036,N_10071);
nand U11525 (N_11525,N_9262,N_9078);
and U11526 (N_11526,N_10200,N_9548);
or U11527 (N_11527,N_9788,N_9096);
nand U11528 (N_11528,N_9745,N_9886);
and U11529 (N_11529,N_9801,N_10422);
nor U11530 (N_11530,N_9831,N_9952);
or U11531 (N_11531,N_10061,N_9698);
nand U11532 (N_11532,N_9561,N_9342);
nand U11533 (N_11533,N_10255,N_10070);
nand U11534 (N_11534,N_9233,N_10416);
or U11535 (N_11535,N_9490,N_9569);
nand U11536 (N_11536,N_9343,N_10055);
nor U11537 (N_11537,N_10096,N_10083);
nor U11538 (N_11538,N_9834,N_9530);
or U11539 (N_11539,N_9409,N_9788);
or U11540 (N_11540,N_10155,N_10289);
nor U11541 (N_11541,N_10180,N_9744);
and U11542 (N_11542,N_9366,N_9781);
or U11543 (N_11543,N_9670,N_9933);
nor U11544 (N_11544,N_9151,N_10411);
and U11545 (N_11545,N_9732,N_10317);
xor U11546 (N_11546,N_10385,N_9892);
nor U11547 (N_11547,N_9211,N_9436);
nor U11548 (N_11548,N_10244,N_9586);
xnor U11549 (N_11549,N_9665,N_10426);
nand U11550 (N_11550,N_9225,N_9492);
nor U11551 (N_11551,N_10319,N_9745);
or U11552 (N_11552,N_10352,N_10483);
and U11553 (N_11553,N_9784,N_10208);
and U11554 (N_11554,N_9360,N_9303);
or U11555 (N_11555,N_10467,N_10247);
or U11556 (N_11556,N_9615,N_10397);
and U11557 (N_11557,N_9559,N_9983);
nor U11558 (N_11558,N_9968,N_9217);
and U11559 (N_11559,N_9693,N_10399);
nand U11560 (N_11560,N_9459,N_10464);
nand U11561 (N_11561,N_9488,N_10243);
and U11562 (N_11562,N_9972,N_9935);
or U11563 (N_11563,N_9751,N_10098);
or U11564 (N_11564,N_9110,N_9715);
and U11565 (N_11565,N_9384,N_10296);
and U11566 (N_11566,N_10485,N_9887);
nor U11567 (N_11567,N_10200,N_9630);
nor U11568 (N_11568,N_9774,N_9114);
and U11569 (N_11569,N_10130,N_9203);
nand U11570 (N_11570,N_9016,N_9213);
xor U11571 (N_11571,N_9093,N_9289);
and U11572 (N_11572,N_9306,N_9895);
and U11573 (N_11573,N_10343,N_9929);
xor U11574 (N_11574,N_10436,N_10020);
and U11575 (N_11575,N_9825,N_9051);
or U11576 (N_11576,N_9832,N_10154);
or U11577 (N_11577,N_9291,N_10243);
nor U11578 (N_11578,N_9365,N_9927);
or U11579 (N_11579,N_10407,N_10073);
nand U11580 (N_11580,N_9594,N_9492);
nor U11581 (N_11581,N_10296,N_10259);
nand U11582 (N_11582,N_10424,N_10090);
xnor U11583 (N_11583,N_9211,N_9763);
or U11584 (N_11584,N_9924,N_9014);
nor U11585 (N_11585,N_9191,N_10006);
nor U11586 (N_11586,N_9801,N_9634);
or U11587 (N_11587,N_9021,N_9650);
and U11588 (N_11588,N_9868,N_9452);
nor U11589 (N_11589,N_10381,N_9373);
nor U11590 (N_11590,N_9549,N_9686);
nand U11591 (N_11591,N_10375,N_9124);
or U11592 (N_11592,N_9934,N_10337);
or U11593 (N_11593,N_9744,N_9046);
or U11594 (N_11594,N_9964,N_9351);
nand U11595 (N_11595,N_9871,N_10022);
nor U11596 (N_11596,N_9701,N_9623);
nand U11597 (N_11597,N_10014,N_10384);
nor U11598 (N_11598,N_9698,N_10100);
and U11599 (N_11599,N_9623,N_10426);
and U11600 (N_11600,N_9442,N_9091);
or U11601 (N_11601,N_9047,N_10223);
or U11602 (N_11602,N_9317,N_9463);
nor U11603 (N_11603,N_10292,N_10020);
and U11604 (N_11604,N_10470,N_10323);
and U11605 (N_11605,N_9284,N_10471);
or U11606 (N_11606,N_9608,N_9963);
or U11607 (N_11607,N_10209,N_9560);
and U11608 (N_11608,N_9612,N_10195);
or U11609 (N_11609,N_9519,N_9981);
nand U11610 (N_11610,N_9614,N_10332);
or U11611 (N_11611,N_9394,N_9313);
or U11612 (N_11612,N_9119,N_9691);
and U11613 (N_11613,N_9775,N_9846);
and U11614 (N_11614,N_9231,N_9912);
nor U11615 (N_11615,N_10123,N_9656);
and U11616 (N_11616,N_10199,N_9878);
and U11617 (N_11617,N_9759,N_9672);
or U11618 (N_11618,N_9737,N_9778);
nand U11619 (N_11619,N_10024,N_9129);
or U11620 (N_11620,N_9982,N_9851);
and U11621 (N_11621,N_9451,N_9879);
nand U11622 (N_11622,N_10462,N_9414);
or U11623 (N_11623,N_10435,N_9818);
xor U11624 (N_11624,N_9035,N_10424);
or U11625 (N_11625,N_10207,N_9841);
nand U11626 (N_11626,N_9433,N_9799);
and U11627 (N_11627,N_10383,N_9364);
nor U11628 (N_11628,N_9840,N_9045);
or U11629 (N_11629,N_10187,N_9794);
and U11630 (N_11630,N_9293,N_10211);
or U11631 (N_11631,N_9373,N_10376);
nand U11632 (N_11632,N_10046,N_10358);
nand U11633 (N_11633,N_9862,N_9974);
or U11634 (N_11634,N_10126,N_10349);
nand U11635 (N_11635,N_10344,N_10173);
xnor U11636 (N_11636,N_9586,N_9273);
nand U11637 (N_11637,N_9735,N_10216);
xnor U11638 (N_11638,N_9852,N_9442);
and U11639 (N_11639,N_9736,N_9348);
or U11640 (N_11640,N_10270,N_9215);
or U11641 (N_11641,N_9915,N_10353);
xor U11642 (N_11642,N_10138,N_9204);
nor U11643 (N_11643,N_10395,N_9717);
xor U11644 (N_11644,N_9748,N_9258);
and U11645 (N_11645,N_10437,N_10405);
nand U11646 (N_11646,N_10357,N_10487);
nor U11647 (N_11647,N_9710,N_9478);
or U11648 (N_11648,N_9460,N_9188);
or U11649 (N_11649,N_10348,N_9271);
and U11650 (N_11650,N_9086,N_9311);
and U11651 (N_11651,N_9506,N_9379);
and U11652 (N_11652,N_9630,N_9381);
nand U11653 (N_11653,N_9480,N_9481);
nor U11654 (N_11654,N_9997,N_10278);
nand U11655 (N_11655,N_10225,N_10351);
xor U11656 (N_11656,N_9462,N_9636);
and U11657 (N_11657,N_9933,N_9342);
or U11658 (N_11658,N_9768,N_10199);
and U11659 (N_11659,N_9404,N_9835);
or U11660 (N_11660,N_10499,N_9454);
nor U11661 (N_11661,N_9432,N_10033);
or U11662 (N_11662,N_10025,N_9447);
or U11663 (N_11663,N_10253,N_9439);
and U11664 (N_11664,N_10238,N_10223);
and U11665 (N_11665,N_9924,N_9930);
nand U11666 (N_11666,N_10132,N_9237);
nor U11667 (N_11667,N_9699,N_9572);
or U11668 (N_11668,N_10420,N_9499);
xnor U11669 (N_11669,N_9837,N_10221);
or U11670 (N_11670,N_9782,N_10410);
xor U11671 (N_11671,N_9439,N_9748);
nand U11672 (N_11672,N_9672,N_9838);
or U11673 (N_11673,N_9619,N_9412);
nand U11674 (N_11674,N_9276,N_10445);
nand U11675 (N_11675,N_9896,N_9063);
nand U11676 (N_11676,N_9567,N_9343);
and U11677 (N_11677,N_9211,N_9957);
nor U11678 (N_11678,N_9725,N_9874);
and U11679 (N_11679,N_9080,N_9424);
nand U11680 (N_11680,N_9878,N_9397);
or U11681 (N_11681,N_9356,N_10454);
and U11682 (N_11682,N_9451,N_9422);
or U11683 (N_11683,N_10133,N_9582);
or U11684 (N_11684,N_9520,N_9693);
and U11685 (N_11685,N_9247,N_9917);
or U11686 (N_11686,N_10268,N_10280);
nand U11687 (N_11687,N_9858,N_9031);
or U11688 (N_11688,N_10122,N_9492);
nor U11689 (N_11689,N_9182,N_9452);
and U11690 (N_11690,N_9126,N_9263);
nand U11691 (N_11691,N_9504,N_10185);
and U11692 (N_11692,N_9115,N_9211);
or U11693 (N_11693,N_10262,N_10232);
nor U11694 (N_11694,N_9254,N_9532);
and U11695 (N_11695,N_10203,N_9595);
or U11696 (N_11696,N_9250,N_10419);
and U11697 (N_11697,N_9508,N_9874);
xnor U11698 (N_11698,N_9074,N_9494);
or U11699 (N_11699,N_10115,N_9911);
and U11700 (N_11700,N_9933,N_9353);
or U11701 (N_11701,N_9785,N_9821);
nor U11702 (N_11702,N_9223,N_9227);
and U11703 (N_11703,N_10369,N_10496);
nand U11704 (N_11704,N_10475,N_10431);
nand U11705 (N_11705,N_9227,N_9889);
nor U11706 (N_11706,N_9925,N_10232);
or U11707 (N_11707,N_9415,N_9523);
nand U11708 (N_11708,N_9785,N_9425);
nor U11709 (N_11709,N_9603,N_9080);
and U11710 (N_11710,N_9481,N_10114);
nand U11711 (N_11711,N_9756,N_10498);
nor U11712 (N_11712,N_9320,N_9081);
nor U11713 (N_11713,N_9080,N_9568);
and U11714 (N_11714,N_9864,N_9352);
nand U11715 (N_11715,N_9576,N_10061);
nor U11716 (N_11716,N_9288,N_9354);
nand U11717 (N_11717,N_9768,N_9287);
or U11718 (N_11718,N_9550,N_9879);
or U11719 (N_11719,N_9170,N_10377);
nor U11720 (N_11720,N_9076,N_10471);
nor U11721 (N_11721,N_9256,N_9282);
nor U11722 (N_11722,N_10470,N_9967);
nor U11723 (N_11723,N_9567,N_9023);
or U11724 (N_11724,N_9330,N_10011);
nand U11725 (N_11725,N_9831,N_9601);
nor U11726 (N_11726,N_9974,N_10174);
nand U11727 (N_11727,N_10005,N_10461);
nor U11728 (N_11728,N_9985,N_9695);
xor U11729 (N_11729,N_9825,N_10040);
xnor U11730 (N_11730,N_10108,N_10391);
nor U11731 (N_11731,N_9989,N_9539);
nand U11732 (N_11732,N_9015,N_9396);
or U11733 (N_11733,N_9849,N_9551);
and U11734 (N_11734,N_10400,N_9043);
nor U11735 (N_11735,N_10471,N_10402);
or U11736 (N_11736,N_9509,N_10170);
or U11737 (N_11737,N_9101,N_9723);
nand U11738 (N_11738,N_9362,N_10095);
or U11739 (N_11739,N_10352,N_10193);
nand U11740 (N_11740,N_9471,N_9806);
and U11741 (N_11741,N_9502,N_9316);
xnor U11742 (N_11742,N_10322,N_9124);
and U11743 (N_11743,N_10133,N_9375);
and U11744 (N_11744,N_10189,N_10311);
xor U11745 (N_11745,N_9008,N_9773);
nor U11746 (N_11746,N_9764,N_9019);
nor U11747 (N_11747,N_9174,N_10125);
nand U11748 (N_11748,N_9958,N_9922);
and U11749 (N_11749,N_9759,N_9197);
nor U11750 (N_11750,N_10096,N_9906);
or U11751 (N_11751,N_10448,N_9917);
or U11752 (N_11752,N_10188,N_9627);
and U11753 (N_11753,N_9637,N_10208);
nand U11754 (N_11754,N_9414,N_9672);
nand U11755 (N_11755,N_10346,N_9513);
xnor U11756 (N_11756,N_9293,N_9925);
nand U11757 (N_11757,N_10119,N_9613);
nor U11758 (N_11758,N_9701,N_9409);
nor U11759 (N_11759,N_9614,N_10325);
nand U11760 (N_11760,N_9639,N_10375);
nand U11761 (N_11761,N_10423,N_10474);
and U11762 (N_11762,N_10057,N_9218);
nor U11763 (N_11763,N_9977,N_9213);
xnor U11764 (N_11764,N_10386,N_10473);
nor U11765 (N_11765,N_10278,N_10439);
or U11766 (N_11766,N_9933,N_10144);
nand U11767 (N_11767,N_10381,N_9209);
nor U11768 (N_11768,N_10420,N_10316);
or U11769 (N_11769,N_9864,N_9306);
and U11770 (N_11770,N_9874,N_10187);
and U11771 (N_11771,N_9429,N_9522);
or U11772 (N_11772,N_9227,N_9534);
or U11773 (N_11773,N_10067,N_9579);
or U11774 (N_11774,N_10139,N_9370);
xnor U11775 (N_11775,N_9117,N_10393);
and U11776 (N_11776,N_10257,N_9766);
xor U11777 (N_11777,N_10234,N_10236);
nand U11778 (N_11778,N_9363,N_10330);
nand U11779 (N_11779,N_10168,N_10367);
xor U11780 (N_11780,N_10052,N_9819);
nor U11781 (N_11781,N_9471,N_9153);
and U11782 (N_11782,N_10223,N_10336);
or U11783 (N_11783,N_9206,N_9604);
nor U11784 (N_11784,N_9599,N_9840);
and U11785 (N_11785,N_9871,N_9113);
nor U11786 (N_11786,N_10219,N_9098);
xor U11787 (N_11787,N_9542,N_9569);
and U11788 (N_11788,N_9095,N_9847);
nor U11789 (N_11789,N_9405,N_9307);
and U11790 (N_11790,N_9822,N_9655);
and U11791 (N_11791,N_9343,N_9980);
nand U11792 (N_11792,N_9741,N_9776);
and U11793 (N_11793,N_9300,N_10074);
nor U11794 (N_11794,N_10370,N_9001);
and U11795 (N_11795,N_9170,N_9888);
or U11796 (N_11796,N_9842,N_9028);
nor U11797 (N_11797,N_9268,N_9750);
and U11798 (N_11798,N_10023,N_9628);
nor U11799 (N_11799,N_10296,N_9596);
nor U11800 (N_11800,N_9215,N_10009);
or U11801 (N_11801,N_10360,N_9866);
or U11802 (N_11802,N_10289,N_10365);
nand U11803 (N_11803,N_10294,N_9379);
and U11804 (N_11804,N_10022,N_10386);
nor U11805 (N_11805,N_10403,N_9424);
and U11806 (N_11806,N_9176,N_9475);
and U11807 (N_11807,N_9575,N_9846);
nor U11808 (N_11808,N_10381,N_9363);
xnor U11809 (N_11809,N_10259,N_10148);
or U11810 (N_11810,N_9724,N_9424);
or U11811 (N_11811,N_9233,N_10049);
nor U11812 (N_11812,N_9257,N_10116);
nand U11813 (N_11813,N_9403,N_9947);
xor U11814 (N_11814,N_10119,N_10086);
nor U11815 (N_11815,N_9664,N_9963);
nand U11816 (N_11816,N_10174,N_10383);
and U11817 (N_11817,N_9918,N_9386);
or U11818 (N_11818,N_10005,N_9015);
and U11819 (N_11819,N_10107,N_9538);
nor U11820 (N_11820,N_10360,N_9202);
and U11821 (N_11821,N_9513,N_9609);
nand U11822 (N_11822,N_9841,N_10063);
or U11823 (N_11823,N_9167,N_10394);
nor U11824 (N_11824,N_9414,N_9221);
xnor U11825 (N_11825,N_9499,N_10352);
nor U11826 (N_11826,N_9877,N_9004);
nand U11827 (N_11827,N_10230,N_9551);
nand U11828 (N_11828,N_9777,N_9041);
nand U11829 (N_11829,N_9546,N_9249);
and U11830 (N_11830,N_9729,N_9049);
nand U11831 (N_11831,N_9011,N_9762);
or U11832 (N_11832,N_10134,N_10480);
nand U11833 (N_11833,N_9046,N_9136);
nand U11834 (N_11834,N_10225,N_10281);
and U11835 (N_11835,N_9783,N_9209);
and U11836 (N_11836,N_10095,N_9223);
and U11837 (N_11837,N_10464,N_9319);
nor U11838 (N_11838,N_9072,N_9240);
or U11839 (N_11839,N_10450,N_9829);
nand U11840 (N_11840,N_9527,N_9512);
or U11841 (N_11841,N_9310,N_10264);
or U11842 (N_11842,N_9833,N_9505);
nor U11843 (N_11843,N_9705,N_9239);
nor U11844 (N_11844,N_9147,N_9886);
nand U11845 (N_11845,N_9335,N_9657);
nor U11846 (N_11846,N_9124,N_9850);
or U11847 (N_11847,N_9721,N_9492);
nand U11848 (N_11848,N_9159,N_9702);
and U11849 (N_11849,N_10344,N_9743);
and U11850 (N_11850,N_10246,N_9540);
and U11851 (N_11851,N_10358,N_9703);
or U11852 (N_11852,N_9519,N_9997);
or U11853 (N_11853,N_10077,N_9077);
nor U11854 (N_11854,N_10160,N_10333);
nand U11855 (N_11855,N_9714,N_9122);
nor U11856 (N_11856,N_10257,N_10206);
or U11857 (N_11857,N_9079,N_9338);
xor U11858 (N_11858,N_10384,N_9626);
nor U11859 (N_11859,N_9733,N_9828);
or U11860 (N_11860,N_9211,N_9920);
nor U11861 (N_11861,N_9677,N_9181);
nand U11862 (N_11862,N_10436,N_9960);
nor U11863 (N_11863,N_9397,N_9381);
nor U11864 (N_11864,N_9597,N_9030);
nand U11865 (N_11865,N_9441,N_10189);
and U11866 (N_11866,N_9617,N_9482);
or U11867 (N_11867,N_9115,N_10044);
nand U11868 (N_11868,N_10164,N_9157);
nor U11869 (N_11869,N_10076,N_10094);
nand U11870 (N_11870,N_10232,N_10100);
and U11871 (N_11871,N_9387,N_9287);
nor U11872 (N_11872,N_9241,N_10354);
and U11873 (N_11873,N_10381,N_9804);
nor U11874 (N_11874,N_9688,N_9610);
xor U11875 (N_11875,N_9600,N_9411);
nand U11876 (N_11876,N_10125,N_9897);
and U11877 (N_11877,N_10462,N_9905);
xnor U11878 (N_11878,N_9388,N_9995);
or U11879 (N_11879,N_10345,N_10033);
or U11880 (N_11880,N_10012,N_9546);
nand U11881 (N_11881,N_9065,N_9670);
nand U11882 (N_11882,N_9678,N_9510);
xnor U11883 (N_11883,N_10143,N_9663);
nand U11884 (N_11884,N_9227,N_9287);
nand U11885 (N_11885,N_10480,N_10496);
nor U11886 (N_11886,N_10393,N_9855);
nand U11887 (N_11887,N_10143,N_9632);
nand U11888 (N_11888,N_9193,N_9349);
nor U11889 (N_11889,N_9228,N_9289);
or U11890 (N_11890,N_9566,N_9076);
nor U11891 (N_11891,N_9003,N_10475);
or U11892 (N_11892,N_9332,N_9708);
nor U11893 (N_11893,N_10338,N_9128);
and U11894 (N_11894,N_9414,N_9524);
nand U11895 (N_11895,N_9301,N_9780);
or U11896 (N_11896,N_9548,N_9063);
nand U11897 (N_11897,N_9488,N_9343);
nor U11898 (N_11898,N_9244,N_10040);
nor U11899 (N_11899,N_9577,N_9995);
nor U11900 (N_11900,N_9690,N_9160);
nor U11901 (N_11901,N_10258,N_10121);
nor U11902 (N_11902,N_10428,N_9119);
and U11903 (N_11903,N_10313,N_9127);
nor U11904 (N_11904,N_9272,N_9703);
nand U11905 (N_11905,N_10175,N_10014);
and U11906 (N_11906,N_9202,N_10043);
nor U11907 (N_11907,N_9332,N_9590);
and U11908 (N_11908,N_9604,N_9849);
nor U11909 (N_11909,N_9456,N_9155);
or U11910 (N_11910,N_9934,N_10054);
and U11911 (N_11911,N_9501,N_10156);
nor U11912 (N_11912,N_10352,N_10300);
and U11913 (N_11913,N_10199,N_9182);
or U11914 (N_11914,N_9087,N_10461);
and U11915 (N_11915,N_9056,N_10245);
nor U11916 (N_11916,N_9820,N_10414);
nor U11917 (N_11917,N_10377,N_10288);
and U11918 (N_11918,N_10242,N_10006);
nand U11919 (N_11919,N_9991,N_9759);
or U11920 (N_11920,N_9985,N_9768);
nor U11921 (N_11921,N_10425,N_10315);
and U11922 (N_11922,N_10344,N_10045);
or U11923 (N_11923,N_9813,N_9251);
or U11924 (N_11924,N_9518,N_10368);
or U11925 (N_11925,N_9347,N_10224);
and U11926 (N_11926,N_9658,N_9435);
nor U11927 (N_11927,N_9799,N_10261);
nand U11928 (N_11928,N_10257,N_10259);
and U11929 (N_11929,N_10050,N_9851);
nand U11930 (N_11930,N_9974,N_9658);
or U11931 (N_11931,N_10300,N_10355);
nor U11932 (N_11932,N_9294,N_10135);
nor U11933 (N_11933,N_10331,N_9759);
or U11934 (N_11934,N_9119,N_9784);
or U11935 (N_11935,N_10120,N_10005);
and U11936 (N_11936,N_10080,N_9868);
and U11937 (N_11937,N_9119,N_9449);
xor U11938 (N_11938,N_9427,N_10342);
and U11939 (N_11939,N_10302,N_10097);
nand U11940 (N_11940,N_9733,N_10181);
nor U11941 (N_11941,N_9286,N_10145);
nor U11942 (N_11942,N_10255,N_9469);
or U11943 (N_11943,N_10046,N_9828);
or U11944 (N_11944,N_9143,N_10139);
nor U11945 (N_11945,N_9010,N_9746);
nor U11946 (N_11946,N_9021,N_10192);
or U11947 (N_11947,N_10247,N_9844);
nand U11948 (N_11948,N_10246,N_10368);
nand U11949 (N_11949,N_9942,N_9289);
or U11950 (N_11950,N_10192,N_9627);
nand U11951 (N_11951,N_9828,N_9980);
or U11952 (N_11952,N_9609,N_9422);
nor U11953 (N_11953,N_10406,N_9289);
nand U11954 (N_11954,N_9613,N_9934);
nand U11955 (N_11955,N_9628,N_9533);
nor U11956 (N_11956,N_10422,N_9103);
or U11957 (N_11957,N_9684,N_9855);
xnor U11958 (N_11958,N_10011,N_9520);
nor U11959 (N_11959,N_10091,N_9390);
nand U11960 (N_11960,N_10438,N_9045);
nor U11961 (N_11961,N_10168,N_9030);
or U11962 (N_11962,N_9258,N_9854);
nand U11963 (N_11963,N_10482,N_9316);
xor U11964 (N_11964,N_10311,N_10191);
and U11965 (N_11965,N_10102,N_9966);
nor U11966 (N_11966,N_10057,N_9080);
nand U11967 (N_11967,N_9507,N_9422);
and U11968 (N_11968,N_10183,N_10023);
and U11969 (N_11969,N_9993,N_9742);
xor U11970 (N_11970,N_9743,N_9358);
nor U11971 (N_11971,N_10147,N_9964);
and U11972 (N_11972,N_10134,N_9814);
nand U11973 (N_11973,N_9902,N_9658);
and U11974 (N_11974,N_9828,N_9494);
or U11975 (N_11975,N_9599,N_9646);
or U11976 (N_11976,N_10011,N_9657);
and U11977 (N_11977,N_9160,N_9494);
nand U11978 (N_11978,N_10052,N_9670);
or U11979 (N_11979,N_9769,N_10036);
and U11980 (N_11980,N_9822,N_10051);
nor U11981 (N_11981,N_10052,N_9203);
xor U11982 (N_11982,N_9413,N_9522);
nand U11983 (N_11983,N_10442,N_9656);
and U11984 (N_11984,N_9699,N_9977);
xnor U11985 (N_11985,N_9825,N_9557);
nand U11986 (N_11986,N_9063,N_9001);
or U11987 (N_11987,N_9961,N_10040);
or U11988 (N_11988,N_9599,N_9119);
nor U11989 (N_11989,N_9255,N_9142);
nand U11990 (N_11990,N_9000,N_10073);
nand U11991 (N_11991,N_10125,N_9606);
nand U11992 (N_11992,N_9518,N_10334);
nand U11993 (N_11993,N_9756,N_9695);
nor U11994 (N_11994,N_9928,N_9997);
xor U11995 (N_11995,N_10112,N_9221);
nand U11996 (N_11996,N_10465,N_9015);
nor U11997 (N_11997,N_10285,N_9916);
nor U11998 (N_11998,N_9606,N_9337);
and U11999 (N_11999,N_10489,N_9682);
nor U12000 (N_12000,N_11954,N_11280);
nand U12001 (N_12001,N_11398,N_11900);
or U12002 (N_12002,N_11069,N_11381);
nor U12003 (N_12003,N_11419,N_11046);
nor U12004 (N_12004,N_10706,N_10764);
nor U12005 (N_12005,N_11603,N_10709);
nor U12006 (N_12006,N_10525,N_11783);
or U12007 (N_12007,N_11786,N_11943);
nor U12008 (N_12008,N_10843,N_10530);
nand U12009 (N_12009,N_11146,N_11974);
nor U12010 (N_12010,N_10559,N_11357);
and U12011 (N_12011,N_11145,N_11843);
xor U12012 (N_12012,N_11952,N_10840);
nor U12013 (N_12013,N_10575,N_11576);
nand U12014 (N_12014,N_10894,N_11653);
and U12015 (N_12015,N_11578,N_11527);
nand U12016 (N_12016,N_11554,N_10993);
nand U12017 (N_12017,N_11832,N_10650);
or U12018 (N_12018,N_10985,N_11841);
and U12019 (N_12019,N_10952,N_11712);
nand U12020 (N_12020,N_11018,N_11403);
nand U12021 (N_12021,N_11243,N_10513);
nor U12022 (N_12022,N_11656,N_10554);
nand U12023 (N_12023,N_10589,N_11983);
and U12024 (N_12024,N_11686,N_11186);
nand U12025 (N_12025,N_11861,N_11256);
nor U12026 (N_12026,N_10850,N_11925);
xor U12027 (N_12027,N_10870,N_10614);
and U12028 (N_12028,N_11168,N_11026);
xor U12029 (N_12029,N_10681,N_11246);
and U12030 (N_12030,N_11912,N_11676);
nand U12031 (N_12031,N_11274,N_10904);
nor U12032 (N_12032,N_10700,N_10760);
and U12033 (N_12033,N_10991,N_11063);
nand U12034 (N_12034,N_11379,N_11140);
nand U12035 (N_12035,N_11557,N_11804);
nor U12036 (N_12036,N_11725,N_10787);
or U12037 (N_12037,N_10823,N_11327);
or U12038 (N_12038,N_11188,N_11698);
nand U12039 (N_12039,N_11992,N_11484);
nor U12040 (N_12040,N_11780,N_10624);
xor U12041 (N_12041,N_11593,N_11628);
and U12042 (N_12042,N_11364,N_10770);
or U12043 (N_12043,N_11680,N_10601);
and U12044 (N_12044,N_11109,N_11015);
or U12045 (N_12045,N_11907,N_11956);
or U12046 (N_12046,N_10917,N_10617);
nand U12047 (N_12047,N_11930,N_10890);
xor U12048 (N_12048,N_10779,N_11763);
nand U12049 (N_12049,N_11309,N_11059);
xnor U12050 (N_12050,N_10645,N_11029);
and U12051 (N_12051,N_11028,N_11201);
nor U12052 (N_12052,N_11815,N_11363);
and U12053 (N_12053,N_10853,N_11771);
and U12054 (N_12054,N_10822,N_11344);
nand U12055 (N_12055,N_11794,N_11627);
nand U12056 (N_12056,N_11629,N_11996);
nor U12057 (N_12057,N_10631,N_10519);
or U12058 (N_12058,N_10983,N_10921);
nand U12059 (N_12059,N_11784,N_10864);
or U12060 (N_12060,N_11916,N_10500);
and U12061 (N_12061,N_11333,N_11547);
nor U12062 (N_12062,N_11453,N_10916);
nand U12063 (N_12063,N_11761,N_10830);
nor U12064 (N_12064,N_11049,N_11623);
and U12065 (N_12065,N_11689,N_11612);
nor U12066 (N_12066,N_10641,N_11194);
or U12067 (N_12067,N_11287,N_11448);
nor U12068 (N_12068,N_10563,N_11733);
nand U12069 (N_12069,N_11849,N_11569);
nor U12070 (N_12070,N_10911,N_10810);
or U12071 (N_12071,N_11110,N_10762);
and U12072 (N_12072,N_11641,N_11831);
nor U12073 (N_12073,N_11105,N_11335);
and U12074 (N_12074,N_11347,N_11673);
xnor U12075 (N_12075,N_11820,N_10714);
xnor U12076 (N_12076,N_11971,N_11944);
or U12077 (N_12077,N_10794,N_11747);
and U12078 (N_12078,N_11542,N_10998);
nor U12079 (N_12079,N_11568,N_11217);
and U12080 (N_12080,N_11423,N_11240);
nand U12081 (N_12081,N_11856,N_11577);
or U12082 (N_12082,N_11894,N_11991);
nand U12083 (N_12083,N_11164,N_11989);
or U12084 (N_12084,N_10701,N_10982);
or U12085 (N_12085,N_11865,N_10776);
nand U12086 (N_12086,N_11898,N_10652);
nand U12087 (N_12087,N_10551,N_11955);
and U12088 (N_12088,N_11125,N_11416);
or U12089 (N_12089,N_11456,N_10646);
nor U12090 (N_12090,N_11135,N_10935);
nor U12091 (N_12091,N_11812,N_11058);
nand U12092 (N_12092,N_11715,N_11077);
nor U12093 (N_12093,N_10540,N_10777);
and U12094 (N_12094,N_11138,N_11850);
and U12095 (N_12095,N_11765,N_11891);
or U12096 (N_12096,N_11480,N_11390);
nand U12097 (N_12097,N_11404,N_11187);
and U12098 (N_12098,N_10541,N_10665);
nor U12099 (N_12099,N_11495,N_11253);
nand U12100 (N_12100,N_11963,N_10817);
xnor U12101 (N_12101,N_11184,N_11793);
nor U12102 (N_12102,N_10842,N_11303);
nand U12103 (N_12103,N_11061,N_11905);
or U12104 (N_12104,N_11910,N_11677);
nand U12105 (N_12105,N_11332,N_11739);
nand U12106 (N_12106,N_11814,N_11090);
nor U12107 (N_12107,N_11491,N_11566);
xor U12108 (N_12108,N_11479,N_11076);
or U12109 (N_12109,N_11564,N_11565);
nor U12110 (N_12110,N_11293,N_11417);
nand U12111 (N_12111,N_10898,N_11034);
or U12112 (N_12112,N_11042,N_10891);
and U12113 (N_12113,N_11133,N_11399);
or U12114 (N_12114,N_11579,N_11618);
or U12115 (N_12115,N_11543,N_10736);
nor U12116 (N_12116,N_10604,N_11769);
nor U12117 (N_12117,N_11016,N_10675);
or U12118 (N_12118,N_11790,N_11070);
or U12119 (N_12119,N_10611,N_11518);
xor U12120 (N_12120,N_11397,N_11643);
nand U12121 (N_12121,N_11463,N_10855);
and U12122 (N_12122,N_10832,N_10887);
and U12123 (N_12123,N_11734,N_10806);
nor U12124 (N_12124,N_11613,N_11402);
and U12125 (N_12125,N_11007,N_11878);
nor U12126 (N_12126,N_11489,N_10883);
nand U12127 (N_12127,N_11252,N_10637);
or U12128 (N_12128,N_10958,N_10612);
nand U12129 (N_12129,N_11047,N_11539);
and U12130 (N_12130,N_11350,N_11057);
and U12131 (N_12131,N_11189,N_10673);
xor U12132 (N_12132,N_11004,N_10862);
nand U12133 (N_12133,N_11202,N_10735);
and U12134 (N_12134,N_11156,N_11107);
and U12135 (N_12135,N_11270,N_11866);
nand U12136 (N_12136,N_11927,N_11592);
nor U12137 (N_12137,N_11979,N_11153);
and U12138 (N_12138,N_11774,N_11251);
nand U12139 (N_12139,N_11699,N_11314);
nor U12140 (N_12140,N_10821,N_11354);
and U12141 (N_12141,N_10802,N_11696);
nor U12142 (N_12142,N_11097,N_11174);
nor U12143 (N_12143,N_11638,N_10992);
or U12144 (N_12144,N_11228,N_11072);
or U12145 (N_12145,N_11237,N_11436);
xor U12146 (N_12146,N_11120,N_11710);
nor U12147 (N_12147,N_11501,N_11407);
xnor U12148 (N_12148,N_11241,N_11606);
and U12149 (N_12149,N_11544,N_11719);
or U12150 (N_12150,N_10741,N_11289);
and U12151 (N_12151,N_11386,N_11585);
nand U12152 (N_12152,N_11721,N_11867);
nor U12153 (N_12153,N_11266,N_11204);
nand U12154 (N_12154,N_11869,N_10786);
or U12155 (N_12155,N_11258,N_10763);
and U12156 (N_12156,N_10867,N_10682);
nand U12157 (N_12157,N_11520,N_10980);
nor U12158 (N_12158,N_10871,N_11119);
nand U12159 (N_12159,N_11352,N_11834);
nor U12160 (N_12160,N_11385,N_10963);
nor U12161 (N_12161,N_11646,N_11493);
nor U12162 (N_12162,N_11446,N_11773);
and U12163 (N_12163,N_11651,N_11548);
nor U12164 (N_12164,N_10987,N_10945);
and U12165 (N_12165,N_11079,N_11755);
and U12166 (N_12166,N_11805,N_11321);
or U12167 (N_12167,N_11249,N_11497);
or U12168 (N_12168,N_11358,N_11770);
nand U12169 (N_12169,N_11908,N_11737);
or U12170 (N_12170,N_11950,N_11506);
xnor U12171 (N_12171,N_10978,N_11600);
and U12172 (N_12172,N_11626,N_10922);
nor U12173 (N_12173,N_11191,N_11876);
nor U12174 (N_12174,N_11563,N_11467);
xnor U12175 (N_12175,N_11648,N_11959);
nand U12176 (N_12176,N_10726,N_10825);
nor U12177 (N_12177,N_10708,N_10946);
and U12178 (N_12178,N_10590,N_11857);
nor U12179 (N_12179,N_11278,N_11683);
nor U12180 (N_12180,N_10717,N_10649);
and U12181 (N_12181,N_11296,N_11978);
and U12182 (N_12182,N_11504,N_10640);
and U12183 (N_12183,N_10954,N_11408);
and U12184 (N_12184,N_11155,N_10550);
nand U12185 (N_12185,N_10561,N_11516);
nor U12186 (N_12186,N_11045,N_11384);
nor U12187 (N_12187,N_10731,N_11764);
or U12188 (N_12188,N_10973,N_11162);
nand U12189 (N_12189,N_11895,N_11224);
nor U12190 (N_12190,N_10555,N_10635);
and U12191 (N_12191,N_11687,N_11019);
and U12192 (N_12192,N_11366,N_11942);
or U12193 (N_12193,N_11893,N_10704);
and U12194 (N_12194,N_10512,N_11036);
nor U12195 (N_12195,N_11681,N_10934);
nor U12196 (N_12196,N_10974,N_11782);
nand U12197 (N_12197,N_11115,N_11055);
nand U12198 (N_12198,N_10620,N_11250);
nor U12199 (N_12199,N_11132,N_11797);
and U12200 (N_12200,N_11661,N_11836);
or U12201 (N_12201,N_11081,N_11432);
or U12202 (N_12202,N_11746,N_11065);
nor U12203 (N_12203,N_11195,N_11167);
and U12204 (N_12204,N_11203,N_10885);
or U12205 (N_12205,N_11339,N_11473);
or U12206 (N_12206,N_11904,N_11617);
nor U12207 (N_12207,N_10615,N_11371);
or U12208 (N_12208,N_10995,N_11172);
and U12209 (N_12209,N_11556,N_10899);
nor U12210 (N_12210,N_11255,N_10877);
nor U12211 (N_12211,N_11645,N_10568);
xnor U12212 (N_12212,N_10651,N_11788);
xnor U12213 (N_12213,N_11796,N_10844);
xor U12214 (N_12214,N_10677,N_10566);
nor U12215 (N_12215,N_10805,N_11177);
nor U12216 (N_12216,N_11795,N_10795);
nor U12217 (N_12217,N_11888,N_11791);
and U12218 (N_12218,N_10502,N_10836);
and U12219 (N_12219,N_10654,N_11136);
or U12220 (N_12220,N_11035,N_11359);
and U12221 (N_12221,N_10831,N_10629);
nor U12222 (N_12222,N_10558,N_11117);
and U12223 (N_12223,N_10564,N_11343);
or U12224 (N_12224,N_11915,N_11089);
or U12225 (N_12225,N_10577,N_11968);
xor U12226 (N_12226,N_11225,N_10979);
nor U12227 (N_12227,N_10543,N_10546);
nor U12228 (N_12228,N_10626,N_10851);
or U12229 (N_12229,N_11748,N_11349);
nand U12230 (N_12230,N_10503,N_10607);
nor U12231 (N_12231,N_11477,N_11936);
nor U12232 (N_12232,N_10661,N_11524);
nand U12233 (N_12233,N_11123,N_11662);
nor U12234 (N_12234,N_11458,N_10854);
nand U12235 (N_12235,N_10723,N_11918);
nor U12236 (N_12236,N_10955,N_11348);
or U12237 (N_12237,N_11512,N_10940);
or U12238 (N_12238,N_11031,N_11011);
or U12239 (N_12239,N_11259,N_10548);
and U12240 (N_12240,N_10660,N_11260);
and U12241 (N_12241,N_11199,N_11754);
nand U12242 (N_12242,N_11395,N_11426);
and U12243 (N_12243,N_11190,N_10508);
or U12244 (N_12244,N_11005,N_10884);
and U12245 (N_12245,N_11457,N_10518);
nand U12246 (N_12246,N_11941,N_11766);
nand U12247 (N_12247,N_11383,N_10610);
or U12248 (N_12248,N_10553,N_11778);
or U12249 (N_12249,N_11736,N_10729);
and U12250 (N_12250,N_11387,N_11127);
and U12251 (N_12251,N_11415,N_10863);
nand U12252 (N_12252,N_10734,N_10964);
nand U12253 (N_12253,N_11649,N_11267);
or U12254 (N_12254,N_11037,N_11660);
nand U12255 (N_12255,N_11032,N_11789);
nor U12256 (N_12256,N_11609,N_11232);
and U12257 (N_12257,N_11206,N_11242);
and U12258 (N_12258,N_11095,N_11562);
xnor U12259 (N_12259,N_11647,N_11500);
nor U12260 (N_12260,N_11182,N_10861);
nor U12261 (N_12261,N_11560,N_10919);
nand U12262 (N_12262,N_10695,N_11903);
nor U12263 (N_12263,N_10730,N_11223);
and U12264 (N_12264,N_11707,N_11892);
nor U12265 (N_12265,N_11210,N_11147);
or U12266 (N_12266,N_11422,N_11842);
or U12267 (N_12267,N_10638,N_11434);
or U12268 (N_12268,N_11541,N_10597);
nand U12269 (N_12269,N_11482,N_11312);
nand U12270 (N_12270,N_11839,N_11702);
nand U12271 (N_12271,N_10686,N_11367);
and U12272 (N_12272,N_11664,N_11311);
and U12273 (N_12273,N_10606,N_11048);
and U12274 (N_12274,N_11284,N_11179);
nand U12275 (N_12275,N_10849,N_11551);
and U12276 (N_12276,N_11205,N_10902);
nor U12277 (N_12277,N_10986,N_11040);
and U12278 (N_12278,N_11990,N_11604);
and U12279 (N_12279,N_10534,N_10981);
xor U12280 (N_12280,N_11802,N_11411);
nand U12281 (N_12281,N_10759,N_10509);
nor U12282 (N_12282,N_11175,N_11444);
and U12283 (N_12283,N_11985,N_11414);
or U12284 (N_12284,N_11083,N_10752);
and U12285 (N_12285,N_10712,N_10959);
nand U12286 (N_12286,N_11957,N_11939);
and U12287 (N_12287,N_10784,N_11762);
nand U12288 (N_12288,N_11540,N_11010);
and U12289 (N_12289,N_10878,N_10608);
and U12290 (N_12290,N_11014,N_10718);
nand U12291 (N_12291,N_11071,N_10803);
or U12292 (N_12292,N_11599,N_11508);
nand U12293 (N_12293,N_11487,N_10965);
or U12294 (N_12294,N_11803,N_11858);
or U12295 (N_12295,N_11811,N_11126);
xnor U12296 (N_12296,N_11180,N_11062);
or U12297 (N_12297,N_11502,N_11781);
xnor U12298 (N_12298,N_11166,N_11142);
or U12299 (N_12299,N_11741,N_11101);
nand U12300 (N_12300,N_10727,N_11345);
nand U12301 (N_12301,N_10761,N_11525);
and U12302 (N_12302,N_11932,N_10679);
nand U12303 (N_12303,N_11396,N_10594);
nand U12304 (N_12304,N_11817,N_11148);
xor U12305 (N_12305,N_10670,N_10848);
xor U12306 (N_12306,N_10684,N_10804);
or U12307 (N_12307,N_11521,N_10600);
and U12308 (N_12308,N_10990,N_10807);
xnor U12309 (N_12309,N_11854,N_11039);
nor U12310 (N_12310,N_10865,N_11052);
or U12311 (N_12311,N_11538,N_11496);
or U12312 (N_12312,N_11519,N_10815);
nand U12313 (N_12313,N_11587,N_11533);
and U12314 (N_12314,N_11933,N_11685);
nand U12315 (N_12315,N_11675,N_10538);
nor U12316 (N_12316,N_11144,N_10957);
nand U12317 (N_12317,N_11598,N_11478);
nor U12318 (N_12318,N_11033,N_11075);
nand U12319 (N_12319,N_11041,N_10627);
nor U12320 (N_12320,N_11437,N_10536);
nor U12321 (N_12321,N_11368,N_11558);
and U12322 (N_12322,N_11691,N_11318);
nand U12323 (N_12323,N_11486,N_10725);
and U12324 (N_12324,N_10542,N_11792);
or U12325 (N_12325,N_11238,N_11948);
nor U12326 (N_12326,N_10720,N_11433);
or U12327 (N_12327,N_11580,N_10621);
and U12328 (N_12328,N_11356,N_11678);
nor U12329 (N_12329,N_11470,N_10814);
nand U12330 (N_12330,N_11295,N_10873);
nand U12331 (N_12331,N_11726,N_11813);
nand U12332 (N_12332,N_11134,N_10926);
and U12333 (N_12333,N_11342,N_10977);
nor U12334 (N_12334,N_11614,N_11254);
and U12335 (N_12335,N_11964,N_10740);
nor U12336 (N_12336,N_11799,N_11161);
nand U12337 (N_12337,N_11716,N_10783);
nand U12338 (N_12338,N_11216,N_10869);
and U12339 (N_12339,N_11392,N_11980);
and U12340 (N_12340,N_11636,N_10808);
xnor U12341 (N_12341,N_10676,N_11022);
xor U12342 (N_12342,N_11735,N_11233);
nand U12343 (N_12343,N_11818,N_10703);
nand U12344 (N_12344,N_11275,N_11310);
or U12345 (N_12345,N_11550,N_11994);
or U12346 (N_12346,N_11438,N_11515);
nand U12347 (N_12347,N_11810,N_11337);
nand U12348 (N_12348,N_10947,N_11672);
xnor U12349 (N_12349,N_10892,N_10586);
nor U12350 (N_12350,N_11002,N_11116);
or U12351 (N_12351,N_11322,N_10596);
nor U12352 (N_12352,N_11909,N_11882);
or U12353 (N_12353,N_11986,N_11196);
nand U12354 (N_12354,N_10966,N_11087);
nor U12355 (N_12355,N_10790,N_11693);
nand U12356 (N_12356,N_11530,N_10571);
or U12357 (N_12357,N_11277,N_11692);
nand U12358 (N_12358,N_11244,N_11630);
xor U12359 (N_12359,N_10782,N_10644);
and U12360 (N_12360,N_11522,N_10860);
xor U12361 (N_12361,N_11001,N_10758);
nand U12362 (N_12362,N_11601,N_11043);
and U12363 (N_12363,N_11605,N_10839);
and U12364 (N_12364,N_11257,N_11513);
nor U12365 (N_12365,N_11624,N_11472);
and U12366 (N_12366,N_10886,N_11999);
and U12367 (N_12367,N_10915,N_11376);
or U12368 (N_12368,N_11634,N_11452);
or U12369 (N_12369,N_11911,N_11425);
nor U12370 (N_12370,N_10948,N_10587);
nor U12371 (N_12371,N_11124,N_11331);
or U12372 (N_12372,N_11724,N_11768);
and U12373 (N_12373,N_11118,N_10507);
nor U12374 (N_12374,N_10569,N_11084);
or U12375 (N_12375,N_11879,N_11325);
xnor U12376 (N_12376,N_11129,N_10636);
or U12377 (N_12377,N_11192,N_10667);
and U12378 (N_12378,N_11787,N_11141);
nor U12379 (N_12379,N_10771,N_10552);
or U12380 (N_12380,N_11406,N_10699);
and U12381 (N_12381,N_11459,N_11870);
nand U12382 (N_12382,N_11485,N_10933);
nor U12383 (N_12383,N_11705,N_10602);
nand U12384 (N_12384,N_11104,N_11292);
xor U12385 (N_12385,N_11455,N_10920);
and U12386 (N_12386,N_11610,N_11775);
and U12387 (N_12387,N_10715,N_11073);
and U12388 (N_12388,N_11102,N_10925);
and U12389 (N_12389,N_11722,N_11785);
nor U12390 (N_12390,N_11960,N_10719);
nor U12391 (N_12391,N_11583,N_11272);
and U12392 (N_12392,N_11380,N_11465);
nor U12393 (N_12393,N_11976,N_11663);
nand U12394 (N_12394,N_11706,N_11896);
and U12395 (N_12395,N_11163,N_11170);
nor U12396 (N_12396,N_10798,N_11669);
or U12397 (N_12397,N_11476,N_11723);
nand U12398 (N_12398,N_11341,N_11239);
xor U12399 (N_12399,N_11466,N_10657);
nor U12400 (N_12400,N_11469,N_11248);
or U12401 (N_12401,N_10801,N_10625);
or U12402 (N_12402,N_11670,N_11505);
xor U12403 (N_12403,N_11640,N_11091);
and U12404 (N_12404,N_10511,N_10756);
nor U12405 (N_12405,N_10506,N_10895);
or U12406 (N_12406,N_11409,N_11833);
nand U12407 (N_12407,N_11958,N_11632);
nand U12408 (N_12408,N_11509,N_10789);
and U12409 (N_12409,N_10927,N_11528);
nand U12410 (N_12410,N_11222,N_11114);
nand U12411 (N_12411,N_10609,N_10984);
xnor U12412 (N_12412,N_10747,N_11567);
nor U12413 (N_12413,N_11286,N_11961);
nand U12414 (N_12414,N_11300,N_11382);
nor U12415 (N_12415,N_11086,N_11622);
and U12416 (N_12416,N_10595,N_11682);
nor U12417 (N_12417,N_10592,N_11099);
nand U12418 (N_12418,N_11092,N_11510);
and U12419 (N_12419,N_11428,N_10888);
nand U12420 (N_12420,N_11602,N_11729);
or U12421 (N_12421,N_10733,N_11657);
and U12422 (N_12422,N_10616,N_11226);
or U12423 (N_12423,N_11694,N_11873);
nor U12424 (N_12424,N_11862,N_11088);
or U12425 (N_12425,N_10793,N_11334);
nor U12426 (N_12426,N_11424,N_11633);
nor U12427 (N_12427,N_11919,N_11975);
and U12428 (N_12428,N_11574,N_11265);
or U12429 (N_12429,N_10580,N_11420);
or U12430 (N_12430,N_11926,N_11157);
or U12431 (N_12431,N_11362,N_11208);
or U12432 (N_12432,N_11100,N_10938);
and U12433 (N_12433,N_10994,N_11695);
and U12434 (N_12434,N_10653,N_11658);
or U12435 (N_12435,N_11094,N_11283);
and U12436 (N_12436,N_11713,N_11835);
or U12437 (N_12437,N_11688,N_11826);
nand U12438 (N_12438,N_11877,N_10574);
and U12439 (N_12439,N_10539,N_11809);
xnor U12440 (N_12440,N_11207,N_10527);
and U12441 (N_12441,N_11532,N_11679);
nand U12442 (N_12442,N_11340,N_11394);
or U12443 (N_12443,N_10944,N_11461);
or U12444 (N_12444,N_11171,N_10531);
nand U12445 (N_12445,N_10576,N_10953);
or U12446 (N_12446,N_11375,N_10929);
and U12447 (N_12447,N_11130,N_11159);
or U12448 (N_12448,N_11374,N_10827);
nor U12449 (N_12449,N_11315,N_11655);
nor U12450 (N_12450,N_11897,N_11523);
nand U12451 (N_12451,N_10785,N_11066);
xnor U12452 (N_12452,N_10713,N_10685);
or U12453 (N_12453,N_11236,N_10603);
xnor U12454 (N_12454,N_10749,N_11131);
and U12455 (N_12455,N_10724,N_10581);
nand U12456 (N_12456,N_11276,N_10750);
nand U12457 (N_12457,N_11981,N_11330);
xnor U12458 (N_12458,N_10562,N_11591);
or U12459 (N_12459,N_10769,N_10874);
or U12460 (N_12460,N_11749,N_10544);
and U12461 (N_12461,N_11137,N_10868);
or U12462 (N_12462,N_11855,N_11701);
xor U12463 (N_12463,N_10989,N_11213);
nor U12464 (N_12464,N_11586,N_11742);
xnor U12465 (N_12465,N_10755,N_11853);
xor U12466 (N_12466,N_11665,N_11984);
or U12467 (N_12467,N_10751,N_11846);
or U12468 (N_12468,N_10767,N_11973);
or U12469 (N_12469,N_11013,N_11752);
nand U12470 (N_12470,N_11700,N_11625);
xor U12471 (N_12471,N_11393,N_11173);
and U12472 (N_12472,N_10634,N_10598);
xor U12473 (N_12473,N_10950,N_10722);
and U12474 (N_12474,N_11447,N_10668);
nand U12475 (N_12475,N_10694,N_11418);
nand U12476 (N_12476,N_11413,N_10570);
or U12477 (N_12477,N_11776,N_11498);
xor U12478 (N_12478,N_10693,N_11934);
nand U12479 (N_12479,N_11490,N_11871);
nand U12480 (N_12480,N_11012,N_10672);
nor U12481 (N_12481,N_11160,N_11008);
and U12482 (N_12482,N_11758,N_10866);
nand U12483 (N_12483,N_11139,N_11261);
or U12484 (N_12484,N_11728,N_11299);
xnor U12485 (N_12485,N_11745,N_11652);
nand U12486 (N_12486,N_10765,N_11922);
and U12487 (N_12487,N_11667,N_10689);
xor U12488 (N_12488,N_11970,N_10516);
or U12489 (N_12489,N_11531,N_11056);
and U12490 (N_12490,N_10690,N_10572);
nor U12491 (N_12491,N_11306,N_11020);
and U12492 (N_12492,N_10876,N_10753);
xnor U12493 (N_12493,N_10528,N_10924);
or U12494 (N_12494,N_11078,N_10584);
nand U12495 (N_12495,N_11581,N_10772);
nand U12496 (N_12496,N_10930,N_10941);
xnor U12497 (N_12497,N_11806,N_11552);
nor U12498 (N_12498,N_10556,N_11355);
nor U12499 (N_12499,N_11914,N_11442);
nand U12500 (N_12500,N_11684,N_11499);
xnor U12501 (N_12501,N_11285,N_10857);
and U12502 (N_12502,N_11517,N_11727);
nor U12503 (N_12503,N_11112,N_11945);
nor U12504 (N_12504,N_11328,N_11731);
nand U12505 (N_12505,N_11017,N_11370);
nand U12506 (N_12506,N_11962,N_11229);
nand U12507 (N_12507,N_10968,N_10943);
or U12508 (N_12508,N_11928,N_11825);
and U12509 (N_12509,N_11740,N_11098);
nand U12510 (N_12510,N_10970,N_11313);
and U12511 (N_12511,N_10656,N_11571);
nor U12512 (N_12512,N_11845,N_10716);
nor U12513 (N_12513,N_11150,N_11732);
nor U12514 (N_12514,N_11711,N_10856);
and U12515 (N_12515,N_11209,N_11537);
or U12516 (N_12516,N_11573,N_11108);
and U12517 (N_12517,N_10613,N_10619);
or U12518 (N_12518,N_11772,N_10529);
and U12519 (N_12519,N_10744,N_11534);
xnor U12520 (N_12520,N_10923,N_10847);
xor U12521 (N_12521,N_11263,N_11924);
or U12522 (N_12522,N_10960,N_10882);
and U12523 (N_12523,N_10545,N_10505);
nor U12524 (N_12524,N_11471,N_10812);
or U12525 (N_12525,N_11848,N_11351);
nand U12526 (N_12526,N_11429,N_10858);
and U12527 (N_12527,N_11621,N_11360);
nand U12528 (N_12528,N_11931,N_11317);
nand U12529 (N_12529,N_11902,N_11273);
and U12530 (N_12530,N_10872,N_11822);
xnor U12531 (N_12531,N_11546,N_11654);
nor U12532 (N_12532,N_11307,N_10648);
nor U12533 (N_12533,N_11947,N_11864);
and U12534 (N_12534,N_11492,N_10939);
or U12535 (N_12535,N_10547,N_10845);
nor U12536 (N_12536,N_10766,N_11800);
nand U12537 (N_12537,N_10510,N_11181);
and U12538 (N_12538,N_11050,N_10800);
nor U12539 (N_12539,N_10622,N_11993);
nand U12540 (N_12540,N_11113,N_11324);
and U12541 (N_12541,N_10692,N_10639);
and U12542 (N_12542,N_10520,N_10897);
nor U12543 (N_12543,N_10514,N_11807);
or U12544 (N_12544,N_11575,N_11128);
nand U12545 (N_12545,N_11619,N_10824);
nor U12546 (N_12546,N_10523,N_11860);
and U12547 (N_12547,N_11709,N_10738);
xor U12548 (N_12548,N_11443,N_10573);
nor U12549 (N_12549,N_11671,N_11951);
and U12550 (N_12550,N_11435,N_11064);
nor U12551 (N_12551,N_11096,N_11427);
nor U12552 (N_12552,N_10737,N_11863);
nor U12553 (N_12553,N_11995,N_11178);
nand U12554 (N_12554,N_11545,N_11218);
nand U12555 (N_12555,N_11106,N_11221);
and U12556 (N_12556,N_11291,N_11756);
and U12557 (N_12557,N_11074,N_11757);
or U12558 (N_12558,N_11234,N_11451);
nand U12559 (N_12559,N_10671,N_11885);
xor U12560 (N_12560,N_11391,N_11561);
nor U12561 (N_12561,N_10702,N_10819);
or U12562 (N_12562,N_11597,N_11365);
xor U12563 (N_12563,N_10837,N_11247);
nor U12564 (N_12564,N_11219,N_11044);
nor U12565 (N_12565,N_11589,N_10746);
and U12566 (N_12566,N_10663,N_10859);
nor U12567 (N_12567,N_10811,N_11481);
nand U12568 (N_12568,N_11053,N_10710);
nor U12569 (N_12569,N_10743,N_11085);
or U12570 (N_12570,N_11720,N_10618);
or U12571 (N_12571,N_11751,N_10937);
nand U12572 (N_12572,N_11889,N_10852);
nor U12573 (N_12573,N_11165,N_10826);
and U12574 (N_12574,N_11559,N_10829);
nor U12575 (N_12575,N_11666,N_11103);
nand U12576 (N_12576,N_10630,N_11838);
nor U12577 (N_12577,N_11886,N_11021);
xor U12578 (N_12578,N_10961,N_11494);
nor U12579 (N_12579,N_11935,N_11967);
or U12580 (N_12580,N_11212,N_10909);
or U12581 (N_12581,N_11025,N_11753);
nand U12582 (N_12582,N_11801,N_11197);
nand U12583 (N_12583,N_11966,N_10903);
nor U12584 (N_12584,N_11744,N_11290);
nand U12585 (N_12585,N_11149,N_10768);
nor U12586 (N_12586,N_11988,N_10788);
nor U12587 (N_12587,N_11308,N_10818);
nor U12588 (N_12588,N_10928,N_11193);
or U12589 (N_12589,N_11302,N_10688);
or U12590 (N_12590,N_11441,N_11859);
nand U12591 (N_12591,N_10905,N_10900);
or U12592 (N_12592,N_11439,N_11828);
nand U12593 (N_12593,N_11875,N_10780);
and U12594 (N_12594,N_10579,N_11767);
or U12595 (N_12595,N_11006,N_11389);
or U12596 (N_12596,N_10698,N_10599);
nand U12597 (N_12597,N_11268,N_11183);
or U12598 (N_12598,N_10951,N_11323);
xnor U12599 (N_12599,N_11827,N_10585);
or U12600 (N_12600,N_10889,N_11326);
nor U12601 (N_12601,N_11030,N_10666);
or U12602 (N_12602,N_11449,N_11608);
nand U12603 (N_12603,N_10683,N_11635);
nand U12604 (N_12604,N_10623,N_11288);
or U12605 (N_12605,N_11111,N_11690);
or U12606 (N_12606,N_11294,N_10647);
and U12607 (N_12607,N_10778,N_10834);
and U12608 (N_12608,N_11514,N_11987);
nand U12609 (N_12609,N_11464,N_11868);
nand U12610 (N_12610,N_11151,N_11169);
and U12611 (N_12611,N_11998,N_10949);
and U12612 (N_12612,N_11642,N_10820);
nor U12613 (N_12613,N_11401,N_11929);
nor U12614 (N_12614,N_11421,N_10691);
or U12615 (N_12615,N_10680,N_10655);
and U12616 (N_12616,N_10797,N_11068);
nor U12617 (N_12617,N_11369,N_11852);
nor U12618 (N_12618,N_11121,N_11594);
and U12619 (N_12619,N_11588,N_11697);
nand U12620 (N_12620,N_11844,N_11483);
nor U12621 (N_12621,N_11823,N_10971);
or U12622 (N_12622,N_11227,N_11759);
nand U12623 (N_12623,N_10526,N_11946);
or U12624 (N_12624,N_11000,N_11329);
nor U12625 (N_12625,N_10732,N_11582);
and U12626 (N_12626,N_11024,N_11440);
and U12627 (N_12627,N_11346,N_10754);
nor U12628 (N_12628,N_11320,N_11220);
nor U12629 (N_12629,N_11198,N_11874);
and U12630 (N_12630,N_11570,N_11297);
and U12631 (N_12631,N_10896,N_10658);
xor U12632 (N_12632,N_10549,N_11837);
nor U12633 (N_12633,N_11884,N_10532);
or U12634 (N_12634,N_11185,N_11282);
nand U12635 (N_12635,N_11659,N_11887);
xor U12636 (N_12636,N_11830,N_11264);
or U12637 (N_12637,N_10567,N_10605);
nor U12638 (N_12638,N_10956,N_10583);
nor U12639 (N_12639,N_11430,N_11215);
nor U12640 (N_12640,N_10932,N_10662);
or U12641 (N_12641,N_11122,N_11840);
xnor U12642 (N_12642,N_11997,N_10914);
nand U12643 (N_12643,N_10969,N_11639);
nand U12644 (N_12644,N_11338,N_11881);
nand U12645 (N_12645,N_11880,N_11474);
nor U12646 (N_12646,N_10999,N_11901);
and U12647 (N_12647,N_11304,N_11230);
nand U12648 (N_12648,N_10535,N_10910);
and U12649 (N_12649,N_11503,N_11631);
nand U12650 (N_12650,N_10643,N_11316);
nor U12651 (N_12651,N_11982,N_11431);
nand U12652 (N_12652,N_11615,N_11301);
and U12653 (N_12653,N_11674,N_11899);
xnor U12654 (N_12654,N_11023,N_11507);
nand U12655 (N_12655,N_11906,N_11271);
or U12656 (N_12656,N_11231,N_11152);
or U12657 (N_12657,N_11262,N_11760);
and U12658 (N_12658,N_10813,N_10664);
and U12659 (N_12659,N_11027,N_11938);
nor U12660 (N_12660,N_10988,N_11003);
and U12661 (N_12661,N_10809,N_11607);
nand U12662 (N_12662,N_10775,N_10838);
and U12663 (N_12663,N_10841,N_10976);
or U12664 (N_12664,N_11535,N_10816);
and U12665 (N_12665,N_11595,N_11200);
nor U12666 (N_12666,N_11596,N_10628);
nor U12667 (N_12667,N_10557,N_11009);
xor U12668 (N_12668,N_10591,N_10517);
and U12669 (N_12669,N_10588,N_11410);
xor U12670 (N_12670,N_11269,N_11620);
or U12671 (N_12671,N_10997,N_11611);
nor U12672 (N_12672,N_11388,N_11245);
nand U12673 (N_12673,N_11176,N_10942);
xnor U12674 (N_12674,N_11779,N_10582);
nand U12675 (N_12675,N_10757,N_11743);
nand U12676 (N_12676,N_11377,N_10687);
or U12677 (N_12677,N_10522,N_10875);
and U12678 (N_12678,N_11038,N_10674);
or U12679 (N_12679,N_11644,N_11450);
or U12680 (N_12680,N_10881,N_11353);
nand U12681 (N_12681,N_10697,N_11305);
xor U12682 (N_12682,N_11279,N_10537);
and U12683 (N_12683,N_10774,N_11953);
and U12684 (N_12684,N_11703,N_11584);
or U12685 (N_12685,N_11214,N_10901);
nor U12686 (N_12686,N_10745,N_10633);
and U12687 (N_12687,N_10833,N_10962);
nor U12688 (N_12688,N_11920,N_11154);
nor U12689 (N_12689,N_11714,N_10796);
nor U12690 (N_12690,N_10893,N_11526);
and U12691 (N_12691,N_10835,N_10828);
or U12692 (N_12692,N_11378,N_11718);
or U12693 (N_12693,N_10879,N_11921);
or U12694 (N_12694,N_11821,N_10678);
nand U12695 (N_12695,N_10906,N_11460);
or U12696 (N_12696,N_11158,N_10880);
and U12697 (N_12697,N_11738,N_11475);
nor U12698 (N_12698,N_11816,N_10907);
nor U12699 (N_12699,N_10972,N_10504);
or U12700 (N_12700,N_11400,N_11298);
xnor U12701 (N_12701,N_11412,N_11445);
or U12702 (N_12702,N_11373,N_11143);
or U12703 (N_12703,N_10781,N_10967);
nand U12704 (N_12704,N_10515,N_11051);
nand U12705 (N_12705,N_10521,N_10728);
or U12706 (N_12706,N_11851,N_11965);
and U12707 (N_12707,N_10593,N_11668);
and U12708 (N_12708,N_10975,N_11372);
nand U12709 (N_12709,N_11977,N_11529);
or U12710 (N_12710,N_10931,N_10996);
nor U12711 (N_12711,N_10711,N_11717);
nand U12712 (N_12712,N_11940,N_11872);
xnor U12713 (N_12713,N_11553,N_11824);
nor U12714 (N_12714,N_10791,N_11468);
or U12715 (N_12715,N_11913,N_10632);
xor U12716 (N_12716,N_11777,N_11650);
nand U12717 (N_12717,N_11704,N_11847);
or U12718 (N_12718,N_11462,N_11555);
nand U12719 (N_12719,N_10913,N_10918);
and U12720 (N_12720,N_10799,N_11949);
nor U12721 (N_12721,N_10578,N_11082);
xor U12722 (N_12722,N_11890,N_11361);
and U12723 (N_12723,N_11211,N_11572);
nor U12724 (N_12724,N_10707,N_10908);
nor U12725 (N_12725,N_10846,N_11488);
xor U12726 (N_12726,N_10773,N_11883);
nor U12727 (N_12727,N_11235,N_11336);
or U12728 (N_12728,N_11281,N_11549);
nor U12729 (N_12729,N_11808,N_11054);
nand U12730 (N_12730,N_11937,N_11829);
and U12731 (N_12731,N_11454,N_11590);
or U12732 (N_12732,N_11730,N_10696);
or U12733 (N_12733,N_11060,N_11637);
nand U12734 (N_12734,N_11080,N_11708);
nand U12735 (N_12735,N_11319,N_10642);
xor U12736 (N_12736,N_10659,N_11511);
or U12737 (N_12737,N_10669,N_11616);
xor U12738 (N_12738,N_11972,N_10565);
nor U12739 (N_12739,N_10912,N_10705);
and U12740 (N_12740,N_10742,N_11798);
xnor U12741 (N_12741,N_11819,N_10739);
and U12742 (N_12742,N_11093,N_11917);
nor U12743 (N_12743,N_11750,N_10501);
nor U12744 (N_12744,N_10792,N_11067);
or U12745 (N_12745,N_11923,N_11536);
nor U12746 (N_12746,N_10936,N_10524);
nor U12747 (N_12747,N_10748,N_10560);
and U12748 (N_12748,N_11969,N_10721);
xnor U12749 (N_12749,N_11405,N_10533);
nor U12750 (N_12750,N_10928,N_11060);
xnor U12751 (N_12751,N_10749,N_11088);
or U12752 (N_12752,N_11339,N_11009);
and U12753 (N_12753,N_11344,N_11764);
nor U12754 (N_12754,N_10727,N_11207);
nand U12755 (N_12755,N_10570,N_10663);
and U12756 (N_12756,N_10992,N_11433);
nor U12757 (N_12757,N_10642,N_11037);
or U12758 (N_12758,N_10564,N_11337);
xor U12759 (N_12759,N_11655,N_11652);
nand U12760 (N_12760,N_10905,N_11652);
and U12761 (N_12761,N_11716,N_11950);
nand U12762 (N_12762,N_11834,N_11848);
nor U12763 (N_12763,N_11202,N_11199);
xor U12764 (N_12764,N_10602,N_11731);
and U12765 (N_12765,N_10662,N_10673);
nor U12766 (N_12766,N_11616,N_10582);
nand U12767 (N_12767,N_11195,N_11446);
and U12768 (N_12768,N_11787,N_10822);
and U12769 (N_12769,N_11160,N_11530);
nand U12770 (N_12770,N_11959,N_11732);
and U12771 (N_12771,N_11332,N_11450);
nor U12772 (N_12772,N_10896,N_11118);
nand U12773 (N_12773,N_11929,N_10509);
or U12774 (N_12774,N_11780,N_11753);
nor U12775 (N_12775,N_11452,N_11815);
nand U12776 (N_12776,N_11816,N_11944);
xnor U12777 (N_12777,N_11231,N_10596);
or U12778 (N_12778,N_11038,N_11471);
nor U12779 (N_12779,N_11001,N_11913);
nor U12780 (N_12780,N_11162,N_11294);
nor U12781 (N_12781,N_10685,N_11536);
and U12782 (N_12782,N_10510,N_11157);
and U12783 (N_12783,N_11176,N_10817);
nor U12784 (N_12784,N_11494,N_11070);
nor U12785 (N_12785,N_11882,N_10673);
or U12786 (N_12786,N_10773,N_11539);
or U12787 (N_12787,N_11556,N_11942);
xnor U12788 (N_12788,N_10721,N_10905);
and U12789 (N_12789,N_11784,N_11692);
and U12790 (N_12790,N_11195,N_10794);
xor U12791 (N_12791,N_10843,N_10526);
nand U12792 (N_12792,N_10798,N_10567);
nor U12793 (N_12793,N_10939,N_10508);
or U12794 (N_12794,N_11329,N_11588);
or U12795 (N_12795,N_11074,N_10551);
xnor U12796 (N_12796,N_11972,N_11475);
or U12797 (N_12797,N_11964,N_10669);
nand U12798 (N_12798,N_11322,N_11918);
nand U12799 (N_12799,N_11382,N_10602);
nor U12800 (N_12800,N_11996,N_10931);
or U12801 (N_12801,N_10631,N_11954);
nor U12802 (N_12802,N_11326,N_11197);
nand U12803 (N_12803,N_11218,N_11021);
and U12804 (N_12804,N_11271,N_11446);
or U12805 (N_12805,N_10548,N_10571);
and U12806 (N_12806,N_11224,N_10695);
nand U12807 (N_12807,N_11347,N_10736);
or U12808 (N_12808,N_11271,N_10582);
and U12809 (N_12809,N_10600,N_11590);
or U12810 (N_12810,N_10889,N_11246);
nand U12811 (N_12811,N_11553,N_10739);
and U12812 (N_12812,N_11247,N_11740);
nor U12813 (N_12813,N_10845,N_11206);
and U12814 (N_12814,N_10877,N_11490);
or U12815 (N_12815,N_11330,N_11224);
and U12816 (N_12816,N_11094,N_11492);
or U12817 (N_12817,N_10792,N_11375);
nand U12818 (N_12818,N_11131,N_11629);
xor U12819 (N_12819,N_10736,N_11795);
or U12820 (N_12820,N_11413,N_11938);
and U12821 (N_12821,N_11722,N_10502);
nor U12822 (N_12822,N_11741,N_11133);
nor U12823 (N_12823,N_11010,N_10709);
nand U12824 (N_12824,N_11547,N_10670);
or U12825 (N_12825,N_10860,N_11549);
or U12826 (N_12826,N_11892,N_11407);
and U12827 (N_12827,N_11945,N_11466);
or U12828 (N_12828,N_11363,N_10948);
nor U12829 (N_12829,N_11549,N_10962);
nor U12830 (N_12830,N_10718,N_11163);
nand U12831 (N_12831,N_10784,N_10544);
and U12832 (N_12832,N_11151,N_11060);
nand U12833 (N_12833,N_10967,N_11107);
or U12834 (N_12834,N_10655,N_10930);
nor U12835 (N_12835,N_10558,N_11194);
and U12836 (N_12836,N_11861,N_11863);
xor U12837 (N_12837,N_10969,N_10572);
nor U12838 (N_12838,N_11311,N_10896);
nor U12839 (N_12839,N_11096,N_11002);
or U12840 (N_12840,N_11322,N_11964);
nor U12841 (N_12841,N_11881,N_10740);
and U12842 (N_12842,N_10541,N_11970);
xor U12843 (N_12843,N_11233,N_11318);
and U12844 (N_12844,N_10836,N_11313);
or U12845 (N_12845,N_11669,N_11280);
or U12846 (N_12846,N_11509,N_10924);
nor U12847 (N_12847,N_11415,N_10530);
nand U12848 (N_12848,N_10957,N_10696);
nand U12849 (N_12849,N_11930,N_11889);
nand U12850 (N_12850,N_10816,N_11779);
or U12851 (N_12851,N_10762,N_11619);
nor U12852 (N_12852,N_11619,N_10607);
or U12853 (N_12853,N_10969,N_11971);
or U12854 (N_12854,N_10631,N_11432);
and U12855 (N_12855,N_11509,N_10999);
and U12856 (N_12856,N_11458,N_11686);
or U12857 (N_12857,N_10577,N_11776);
and U12858 (N_12858,N_11264,N_10939);
xor U12859 (N_12859,N_11622,N_10517);
xnor U12860 (N_12860,N_10996,N_11456);
nand U12861 (N_12861,N_10771,N_11854);
nand U12862 (N_12862,N_10706,N_11094);
and U12863 (N_12863,N_11288,N_11133);
nor U12864 (N_12864,N_10949,N_11810);
nand U12865 (N_12865,N_11225,N_11035);
or U12866 (N_12866,N_10796,N_10580);
nor U12867 (N_12867,N_11501,N_11360);
xnor U12868 (N_12868,N_11289,N_11667);
nand U12869 (N_12869,N_11284,N_11802);
nor U12870 (N_12870,N_10842,N_10751);
and U12871 (N_12871,N_11964,N_10635);
or U12872 (N_12872,N_11017,N_11719);
nand U12873 (N_12873,N_11484,N_11275);
xor U12874 (N_12874,N_10601,N_11391);
or U12875 (N_12875,N_10886,N_11753);
or U12876 (N_12876,N_11439,N_11474);
nor U12877 (N_12877,N_10790,N_11268);
nand U12878 (N_12878,N_11631,N_11167);
nand U12879 (N_12879,N_10919,N_11966);
and U12880 (N_12880,N_11885,N_11999);
nand U12881 (N_12881,N_11759,N_11659);
xor U12882 (N_12882,N_11284,N_10698);
and U12883 (N_12883,N_10565,N_10916);
nand U12884 (N_12884,N_10762,N_10579);
nand U12885 (N_12885,N_11125,N_11495);
and U12886 (N_12886,N_10647,N_11210);
or U12887 (N_12887,N_10527,N_11168);
nor U12888 (N_12888,N_11659,N_11840);
nand U12889 (N_12889,N_11649,N_10762);
nor U12890 (N_12890,N_11285,N_11293);
and U12891 (N_12891,N_11542,N_11612);
or U12892 (N_12892,N_10645,N_10956);
or U12893 (N_12893,N_11986,N_10619);
nand U12894 (N_12894,N_11804,N_11312);
or U12895 (N_12895,N_11257,N_11588);
xor U12896 (N_12896,N_11906,N_11523);
and U12897 (N_12897,N_11903,N_11352);
and U12898 (N_12898,N_10873,N_11067);
xnor U12899 (N_12899,N_11925,N_11592);
or U12900 (N_12900,N_11077,N_11520);
and U12901 (N_12901,N_10694,N_11840);
and U12902 (N_12902,N_10771,N_10754);
nor U12903 (N_12903,N_11992,N_11755);
nor U12904 (N_12904,N_10934,N_10599);
or U12905 (N_12905,N_11049,N_11019);
and U12906 (N_12906,N_10718,N_10788);
and U12907 (N_12907,N_10765,N_10518);
and U12908 (N_12908,N_11584,N_11477);
nor U12909 (N_12909,N_11141,N_11750);
xnor U12910 (N_12910,N_11745,N_10547);
or U12911 (N_12911,N_11765,N_11432);
and U12912 (N_12912,N_11498,N_11681);
or U12913 (N_12913,N_11077,N_11158);
xnor U12914 (N_12914,N_10937,N_11946);
nand U12915 (N_12915,N_11554,N_11004);
or U12916 (N_12916,N_11722,N_11799);
nor U12917 (N_12917,N_11375,N_11898);
nor U12918 (N_12918,N_11865,N_11776);
nand U12919 (N_12919,N_10591,N_11241);
and U12920 (N_12920,N_10620,N_11863);
nand U12921 (N_12921,N_11403,N_11499);
or U12922 (N_12922,N_10754,N_10930);
nand U12923 (N_12923,N_11971,N_11793);
or U12924 (N_12924,N_11184,N_11975);
or U12925 (N_12925,N_10620,N_10945);
xnor U12926 (N_12926,N_11895,N_10915);
or U12927 (N_12927,N_11461,N_11931);
xor U12928 (N_12928,N_10649,N_11192);
nor U12929 (N_12929,N_11327,N_10649);
nor U12930 (N_12930,N_11325,N_11883);
or U12931 (N_12931,N_10814,N_11314);
or U12932 (N_12932,N_10733,N_11472);
nand U12933 (N_12933,N_11476,N_10815);
and U12934 (N_12934,N_11651,N_11038);
or U12935 (N_12935,N_11255,N_11850);
nand U12936 (N_12936,N_11658,N_11286);
or U12937 (N_12937,N_11783,N_10769);
nand U12938 (N_12938,N_11243,N_11750);
and U12939 (N_12939,N_10600,N_11458);
nand U12940 (N_12940,N_11351,N_11615);
nand U12941 (N_12941,N_11876,N_10734);
nor U12942 (N_12942,N_11530,N_11776);
nor U12943 (N_12943,N_11939,N_10580);
or U12944 (N_12944,N_11886,N_11166);
nor U12945 (N_12945,N_11914,N_10663);
nand U12946 (N_12946,N_11882,N_11832);
nand U12947 (N_12947,N_10711,N_10549);
nand U12948 (N_12948,N_11993,N_11360);
and U12949 (N_12949,N_11237,N_10528);
nor U12950 (N_12950,N_11197,N_10709);
and U12951 (N_12951,N_11772,N_10726);
nand U12952 (N_12952,N_10933,N_11615);
nor U12953 (N_12953,N_10694,N_10925);
nand U12954 (N_12954,N_10655,N_10886);
and U12955 (N_12955,N_11779,N_11407);
and U12956 (N_12956,N_11687,N_11442);
nor U12957 (N_12957,N_11402,N_11978);
or U12958 (N_12958,N_10622,N_10906);
or U12959 (N_12959,N_10683,N_11974);
or U12960 (N_12960,N_11260,N_11448);
nor U12961 (N_12961,N_11904,N_10622);
nor U12962 (N_12962,N_11579,N_11843);
or U12963 (N_12963,N_11742,N_11080);
nor U12964 (N_12964,N_11286,N_11076);
or U12965 (N_12965,N_11569,N_10989);
nand U12966 (N_12966,N_11234,N_11704);
nand U12967 (N_12967,N_10652,N_11008);
or U12968 (N_12968,N_11686,N_10509);
nand U12969 (N_12969,N_10792,N_11048);
nand U12970 (N_12970,N_11081,N_11428);
xnor U12971 (N_12971,N_11827,N_11180);
nor U12972 (N_12972,N_11707,N_11710);
and U12973 (N_12973,N_11585,N_10776);
xnor U12974 (N_12974,N_10551,N_10749);
or U12975 (N_12975,N_11798,N_11278);
or U12976 (N_12976,N_11619,N_10944);
nor U12977 (N_12977,N_10729,N_11857);
or U12978 (N_12978,N_11965,N_10966);
nand U12979 (N_12979,N_11830,N_10815);
nand U12980 (N_12980,N_11004,N_11709);
and U12981 (N_12981,N_10753,N_10538);
nor U12982 (N_12982,N_11369,N_11602);
or U12983 (N_12983,N_11049,N_10756);
or U12984 (N_12984,N_10750,N_11215);
or U12985 (N_12985,N_11390,N_11594);
nand U12986 (N_12986,N_10633,N_11747);
nand U12987 (N_12987,N_11413,N_10885);
and U12988 (N_12988,N_11627,N_11014);
nand U12989 (N_12989,N_11931,N_10835);
and U12990 (N_12990,N_10989,N_11877);
or U12991 (N_12991,N_10753,N_10794);
and U12992 (N_12992,N_11448,N_11283);
and U12993 (N_12993,N_11336,N_10889);
or U12994 (N_12994,N_11804,N_11243);
or U12995 (N_12995,N_11863,N_11616);
nor U12996 (N_12996,N_11223,N_11106);
nand U12997 (N_12997,N_11984,N_10519);
nand U12998 (N_12998,N_11521,N_11708);
nor U12999 (N_12999,N_11002,N_11439);
and U13000 (N_13000,N_10884,N_11703);
nor U13001 (N_13001,N_11469,N_11730);
or U13002 (N_13002,N_11017,N_10570);
or U13003 (N_13003,N_11527,N_11417);
nor U13004 (N_13004,N_10831,N_10504);
nor U13005 (N_13005,N_11409,N_11125);
or U13006 (N_13006,N_11519,N_11995);
nand U13007 (N_13007,N_10821,N_11926);
nor U13008 (N_13008,N_10954,N_11997);
and U13009 (N_13009,N_11801,N_10736);
nor U13010 (N_13010,N_11253,N_11082);
and U13011 (N_13011,N_11092,N_11519);
and U13012 (N_13012,N_10676,N_11964);
and U13013 (N_13013,N_10555,N_11920);
or U13014 (N_13014,N_11303,N_10912);
nand U13015 (N_13015,N_11952,N_11793);
and U13016 (N_13016,N_11377,N_11668);
nand U13017 (N_13017,N_11307,N_11937);
and U13018 (N_13018,N_10864,N_11904);
xor U13019 (N_13019,N_11051,N_11211);
and U13020 (N_13020,N_11216,N_11000);
and U13021 (N_13021,N_11635,N_10659);
or U13022 (N_13022,N_10588,N_10695);
or U13023 (N_13023,N_11006,N_11851);
and U13024 (N_13024,N_10877,N_11914);
and U13025 (N_13025,N_10632,N_11194);
nand U13026 (N_13026,N_10730,N_11640);
nand U13027 (N_13027,N_11378,N_11391);
nand U13028 (N_13028,N_11623,N_10820);
or U13029 (N_13029,N_11076,N_11982);
nand U13030 (N_13030,N_11794,N_11418);
or U13031 (N_13031,N_10752,N_11008);
xor U13032 (N_13032,N_11658,N_10681);
nand U13033 (N_13033,N_10722,N_11721);
nand U13034 (N_13034,N_10761,N_10991);
and U13035 (N_13035,N_11156,N_10655);
nor U13036 (N_13036,N_11292,N_10733);
or U13037 (N_13037,N_11300,N_11964);
nor U13038 (N_13038,N_10797,N_10833);
nor U13039 (N_13039,N_11077,N_11591);
or U13040 (N_13040,N_11180,N_11684);
nor U13041 (N_13041,N_11888,N_11334);
nor U13042 (N_13042,N_11407,N_11346);
or U13043 (N_13043,N_11761,N_11471);
nor U13044 (N_13044,N_10519,N_11300);
nor U13045 (N_13045,N_11200,N_11655);
or U13046 (N_13046,N_10735,N_11991);
nand U13047 (N_13047,N_11455,N_10780);
nor U13048 (N_13048,N_11170,N_10756);
or U13049 (N_13049,N_11969,N_10915);
nand U13050 (N_13050,N_11558,N_10698);
and U13051 (N_13051,N_10618,N_11920);
nand U13052 (N_13052,N_10546,N_10941);
or U13053 (N_13053,N_10559,N_11445);
and U13054 (N_13054,N_11365,N_10669);
nor U13055 (N_13055,N_11244,N_11153);
or U13056 (N_13056,N_11999,N_11129);
nand U13057 (N_13057,N_10988,N_11261);
xnor U13058 (N_13058,N_10899,N_11204);
nor U13059 (N_13059,N_11541,N_11031);
or U13060 (N_13060,N_10917,N_11994);
and U13061 (N_13061,N_11268,N_11404);
nand U13062 (N_13062,N_10919,N_11096);
and U13063 (N_13063,N_10728,N_11741);
nand U13064 (N_13064,N_10952,N_10707);
nand U13065 (N_13065,N_11284,N_11422);
or U13066 (N_13066,N_11406,N_11864);
and U13067 (N_13067,N_11972,N_10904);
nor U13068 (N_13068,N_11146,N_11689);
or U13069 (N_13069,N_10541,N_11418);
and U13070 (N_13070,N_10517,N_11424);
nand U13071 (N_13071,N_10981,N_10984);
nand U13072 (N_13072,N_11824,N_11859);
nand U13073 (N_13073,N_11887,N_11336);
and U13074 (N_13074,N_10852,N_11637);
nand U13075 (N_13075,N_11656,N_10882);
or U13076 (N_13076,N_11830,N_11439);
and U13077 (N_13077,N_11160,N_11187);
nand U13078 (N_13078,N_11018,N_10876);
or U13079 (N_13079,N_11114,N_11567);
xor U13080 (N_13080,N_11763,N_11610);
nor U13081 (N_13081,N_11914,N_10854);
xnor U13082 (N_13082,N_11705,N_11544);
nand U13083 (N_13083,N_11492,N_10796);
nand U13084 (N_13084,N_11550,N_11249);
xor U13085 (N_13085,N_11683,N_10867);
or U13086 (N_13086,N_11400,N_11119);
and U13087 (N_13087,N_10594,N_11089);
and U13088 (N_13088,N_11965,N_11431);
xor U13089 (N_13089,N_11934,N_10773);
nand U13090 (N_13090,N_11900,N_11530);
or U13091 (N_13091,N_10631,N_11068);
and U13092 (N_13092,N_11633,N_11135);
nand U13093 (N_13093,N_11566,N_11814);
nand U13094 (N_13094,N_11348,N_11198);
nor U13095 (N_13095,N_11125,N_10713);
nand U13096 (N_13096,N_11956,N_11431);
nand U13097 (N_13097,N_11956,N_10670);
nor U13098 (N_13098,N_10826,N_11324);
and U13099 (N_13099,N_11644,N_11815);
nor U13100 (N_13100,N_10978,N_11534);
nor U13101 (N_13101,N_11185,N_11348);
or U13102 (N_13102,N_10669,N_10531);
or U13103 (N_13103,N_11423,N_10590);
and U13104 (N_13104,N_10688,N_11155);
and U13105 (N_13105,N_11333,N_11687);
nand U13106 (N_13106,N_10517,N_11872);
and U13107 (N_13107,N_10558,N_11946);
or U13108 (N_13108,N_11741,N_10692);
nor U13109 (N_13109,N_11987,N_11580);
nand U13110 (N_13110,N_11436,N_11161);
or U13111 (N_13111,N_10792,N_10978);
nand U13112 (N_13112,N_10871,N_10974);
or U13113 (N_13113,N_11146,N_11991);
nand U13114 (N_13114,N_11388,N_11369);
and U13115 (N_13115,N_11930,N_10856);
and U13116 (N_13116,N_10883,N_10928);
and U13117 (N_13117,N_11570,N_10572);
nand U13118 (N_13118,N_10621,N_11714);
or U13119 (N_13119,N_11131,N_11307);
nor U13120 (N_13120,N_10552,N_10519);
and U13121 (N_13121,N_11774,N_11044);
or U13122 (N_13122,N_10580,N_11785);
nor U13123 (N_13123,N_11872,N_11647);
or U13124 (N_13124,N_11302,N_11771);
nor U13125 (N_13125,N_11079,N_11686);
or U13126 (N_13126,N_10981,N_11570);
or U13127 (N_13127,N_11192,N_10707);
or U13128 (N_13128,N_11368,N_11121);
or U13129 (N_13129,N_11432,N_11103);
xor U13130 (N_13130,N_10944,N_11832);
and U13131 (N_13131,N_10698,N_11323);
or U13132 (N_13132,N_11896,N_11833);
and U13133 (N_13133,N_11822,N_11427);
or U13134 (N_13134,N_10720,N_10776);
nor U13135 (N_13135,N_10763,N_11326);
or U13136 (N_13136,N_10975,N_10960);
or U13137 (N_13137,N_11721,N_11877);
nor U13138 (N_13138,N_11620,N_10875);
nand U13139 (N_13139,N_11943,N_11351);
and U13140 (N_13140,N_11953,N_11132);
or U13141 (N_13141,N_11171,N_10692);
nand U13142 (N_13142,N_11932,N_10864);
nand U13143 (N_13143,N_11371,N_11342);
and U13144 (N_13144,N_10767,N_10757);
or U13145 (N_13145,N_11773,N_11801);
and U13146 (N_13146,N_11939,N_11905);
nand U13147 (N_13147,N_10900,N_10518);
nand U13148 (N_13148,N_11070,N_11898);
nor U13149 (N_13149,N_10878,N_10739);
xor U13150 (N_13150,N_10671,N_11871);
and U13151 (N_13151,N_10717,N_11815);
nand U13152 (N_13152,N_10596,N_11779);
and U13153 (N_13153,N_11740,N_11946);
and U13154 (N_13154,N_11383,N_11430);
nand U13155 (N_13155,N_11032,N_11993);
nand U13156 (N_13156,N_11059,N_10767);
or U13157 (N_13157,N_10918,N_11718);
nor U13158 (N_13158,N_11492,N_11460);
or U13159 (N_13159,N_10643,N_11569);
xnor U13160 (N_13160,N_11753,N_11350);
nor U13161 (N_13161,N_11964,N_11121);
or U13162 (N_13162,N_11231,N_11642);
and U13163 (N_13163,N_11760,N_11685);
nor U13164 (N_13164,N_10961,N_10643);
nand U13165 (N_13165,N_10980,N_11242);
or U13166 (N_13166,N_10926,N_10849);
nand U13167 (N_13167,N_11771,N_10724);
or U13168 (N_13168,N_11584,N_11133);
nand U13169 (N_13169,N_11300,N_10722);
nand U13170 (N_13170,N_11028,N_10737);
nand U13171 (N_13171,N_11068,N_10774);
nor U13172 (N_13172,N_11964,N_11974);
and U13173 (N_13173,N_11844,N_10891);
and U13174 (N_13174,N_11737,N_11388);
nor U13175 (N_13175,N_11856,N_10710);
nand U13176 (N_13176,N_11612,N_10544);
and U13177 (N_13177,N_11557,N_10674);
or U13178 (N_13178,N_11297,N_10538);
nor U13179 (N_13179,N_11751,N_11646);
nor U13180 (N_13180,N_11523,N_11122);
nor U13181 (N_13181,N_11072,N_11989);
and U13182 (N_13182,N_11993,N_11544);
nor U13183 (N_13183,N_11842,N_11506);
nor U13184 (N_13184,N_10834,N_11523);
and U13185 (N_13185,N_10678,N_10847);
nor U13186 (N_13186,N_11895,N_11228);
xor U13187 (N_13187,N_11444,N_11422);
nand U13188 (N_13188,N_10730,N_11496);
xor U13189 (N_13189,N_11879,N_11740);
nand U13190 (N_13190,N_10981,N_11532);
or U13191 (N_13191,N_11393,N_10663);
and U13192 (N_13192,N_10689,N_11657);
xor U13193 (N_13193,N_10528,N_11368);
nand U13194 (N_13194,N_11444,N_11418);
xor U13195 (N_13195,N_11271,N_10848);
nand U13196 (N_13196,N_10923,N_11448);
nand U13197 (N_13197,N_11044,N_11353);
or U13198 (N_13198,N_11630,N_11311);
and U13199 (N_13199,N_11785,N_11900);
nor U13200 (N_13200,N_11473,N_11640);
nor U13201 (N_13201,N_11584,N_11656);
and U13202 (N_13202,N_10816,N_11638);
nand U13203 (N_13203,N_11198,N_10909);
or U13204 (N_13204,N_11781,N_10615);
xnor U13205 (N_13205,N_11475,N_11425);
nand U13206 (N_13206,N_11751,N_10691);
nand U13207 (N_13207,N_11804,N_11817);
nor U13208 (N_13208,N_11784,N_11080);
xor U13209 (N_13209,N_11802,N_10702);
nor U13210 (N_13210,N_11517,N_10900);
nand U13211 (N_13211,N_10744,N_11548);
nor U13212 (N_13212,N_10707,N_10859);
nand U13213 (N_13213,N_11214,N_10821);
xnor U13214 (N_13214,N_11429,N_10793);
nor U13215 (N_13215,N_10880,N_11252);
or U13216 (N_13216,N_10962,N_11601);
nand U13217 (N_13217,N_11645,N_11043);
nand U13218 (N_13218,N_11236,N_10787);
nand U13219 (N_13219,N_10840,N_11692);
and U13220 (N_13220,N_10943,N_10671);
xor U13221 (N_13221,N_11365,N_11844);
nand U13222 (N_13222,N_10941,N_11610);
and U13223 (N_13223,N_11489,N_11456);
xor U13224 (N_13224,N_10751,N_10966);
nand U13225 (N_13225,N_11764,N_11574);
nand U13226 (N_13226,N_10689,N_10567);
xor U13227 (N_13227,N_10505,N_10783);
nor U13228 (N_13228,N_11307,N_10951);
and U13229 (N_13229,N_11939,N_11705);
or U13230 (N_13230,N_11382,N_10639);
or U13231 (N_13231,N_10866,N_10925);
and U13232 (N_13232,N_11710,N_11121);
and U13233 (N_13233,N_10917,N_11645);
and U13234 (N_13234,N_10779,N_11649);
nand U13235 (N_13235,N_10588,N_10610);
nand U13236 (N_13236,N_10701,N_11715);
and U13237 (N_13237,N_11997,N_11046);
or U13238 (N_13238,N_11160,N_10687);
nor U13239 (N_13239,N_11606,N_10709);
or U13240 (N_13240,N_10894,N_11409);
and U13241 (N_13241,N_11437,N_11738);
or U13242 (N_13242,N_10643,N_11835);
and U13243 (N_13243,N_10511,N_11016);
and U13244 (N_13244,N_11122,N_10601);
nor U13245 (N_13245,N_10682,N_11604);
and U13246 (N_13246,N_11569,N_11880);
xnor U13247 (N_13247,N_11053,N_10553);
nor U13248 (N_13248,N_11212,N_11116);
and U13249 (N_13249,N_11262,N_11962);
or U13250 (N_13250,N_11830,N_10782);
or U13251 (N_13251,N_11541,N_11760);
xor U13252 (N_13252,N_11087,N_11333);
or U13253 (N_13253,N_11424,N_10567);
xor U13254 (N_13254,N_10812,N_10630);
or U13255 (N_13255,N_10876,N_11335);
and U13256 (N_13256,N_11132,N_11473);
or U13257 (N_13257,N_11608,N_11733);
nand U13258 (N_13258,N_11396,N_11907);
nand U13259 (N_13259,N_10928,N_11609);
nand U13260 (N_13260,N_11046,N_10527);
xor U13261 (N_13261,N_11332,N_11356);
nand U13262 (N_13262,N_11646,N_10840);
and U13263 (N_13263,N_10797,N_11934);
nand U13264 (N_13264,N_11232,N_11485);
nand U13265 (N_13265,N_11069,N_10713);
or U13266 (N_13266,N_10720,N_10781);
nor U13267 (N_13267,N_11550,N_11555);
nor U13268 (N_13268,N_10708,N_10653);
nor U13269 (N_13269,N_10652,N_10974);
or U13270 (N_13270,N_11552,N_10992);
and U13271 (N_13271,N_11771,N_11469);
and U13272 (N_13272,N_11580,N_11171);
nor U13273 (N_13273,N_11254,N_11049);
or U13274 (N_13274,N_11893,N_11866);
nor U13275 (N_13275,N_10559,N_11160);
nand U13276 (N_13276,N_10668,N_10785);
nor U13277 (N_13277,N_11936,N_10561);
xor U13278 (N_13278,N_11771,N_10635);
nand U13279 (N_13279,N_10786,N_11566);
or U13280 (N_13280,N_11768,N_11437);
or U13281 (N_13281,N_10737,N_11673);
nand U13282 (N_13282,N_10615,N_10596);
or U13283 (N_13283,N_11799,N_10636);
and U13284 (N_13284,N_11658,N_10541);
and U13285 (N_13285,N_10933,N_10947);
or U13286 (N_13286,N_10933,N_11155);
and U13287 (N_13287,N_11303,N_11225);
nor U13288 (N_13288,N_11448,N_11288);
nand U13289 (N_13289,N_11825,N_11157);
or U13290 (N_13290,N_10799,N_11525);
or U13291 (N_13291,N_11071,N_11710);
and U13292 (N_13292,N_11341,N_10784);
and U13293 (N_13293,N_11393,N_10725);
nand U13294 (N_13294,N_11961,N_11931);
xnor U13295 (N_13295,N_11799,N_10692);
nor U13296 (N_13296,N_10660,N_11994);
and U13297 (N_13297,N_11432,N_11943);
nor U13298 (N_13298,N_11598,N_11405);
nor U13299 (N_13299,N_11897,N_11098);
nor U13300 (N_13300,N_11592,N_10875);
and U13301 (N_13301,N_10843,N_11534);
and U13302 (N_13302,N_11192,N_11952);
or U13303 (N_13303,N_11982,N_10824);
and U13304 (N_13304,N_10746,N_10867);
and U13305 (N_13305,N_11607,N_11268);
nand U13306 (N_13306,N_10592,N_11190);
nor U13307 (N_13307,N_11885,N_10780);
or U13308 (N_13308,N_10583,N_11940);
and U13309 (N_13309,N_11307,N_11414);
nand U13310 (N_13310,N_11751,N_11231);
nor U13311 (N_13311,N_11932,N_11427);
nor U13312 (N_13312,N_11518,N_11063);
or U13313 (N_13313,N_11528,N_11489);
and U13314 (N_13314,N_10868,N_11488);
nand U13315 (N_13315,N_11936,N_11260);
xnor U13316 (N_13316,N_10624,N_11367);
xnor U13317 (N_13317,N_11732,N_10819);
nand U13318 (N_13318,N_10921,N_10974);
and U13319 (N_13319,N_11564,N_11716);
xor U13320 (N_13320,N_11327,N_11628);
nor U13321 (N_13321,N_11943,N_11673);
and U13322 (N_13322,N_11188,N_10892);
nor U13323 (N_13323,N_10861,N_11439);
or U13324 (N_13324,N_10799,N_10570);
nand U13325 (N_13325,N_11437,N_11002);
or U13326 (N_13326,N_10684,N_11564);
and U13327 (N_13327,N_11114,N_10801);
nand U13328 (N_13328,N_11476,N_11308);
or U13329 (N_13329,N_11325,N_11724);
nand U13330 (N_13330,N_11457,N_10710);
nand U13331 (N_13331,N_10873,N_10942);
nor U13332 (N_13332,N_11772,N_11719);
and U13333 (N_13333,N_11690,N_11986);
or U13334 (N_13334,N_11240,N_10669);
nor U13335 (N_13335,N_11541,N_11030);
nand U13336 (N_13336,N_11240,N_11431);
and U13337 (N_13337,N_11694,N_11916);
nor U13338 (N_13338,N_10794,N_11518);
and U13339 (N_13339,N_11425,N_11825);
or U13340 (N_13340,N_10655,N_10864);
and U13341 (N_13341,N_11401,N_11466);
and U13342 (N_13342,N_11884,N_10626);
nor U13343 (N_13343,N_10926,N_11306);
or U13344 (N_13344,N_11820,N_10834);
nand U13345 (N_13345,N_10909,N_11736);
nor U13346 (N_13346,N_11844,N_11623);
or U13347 (N_13347,N_10528,N_11866);
nor U13348 (N_13348,N_11263,N_11640);
and U13349 (N_13349,N_11608,N_11095);
nand U13350 (N_13350,N_11300,N_11850);
or U13351 (N_13351,N_11606,N_11750);
or U13352 (N_13352,N_11353,N_10754);
and U13353 (N_13353,N_11736,N_11734);
nor U13354 (N_13354,N_10524,N_10949);
nor U13355 (N_13355,N_10869,N_11766);
xnor U13356 (N_13356,N_11575,N_11748);
nand U13357 (N_13357,N_10906,N_11228);
nor U13358 (N_13358,N_11694,N_10572);
nand U13359 (N_13359,N_10554,N_10790);
nor U13360 (N_13360,N_10536,N_11967);
or U13361 (N_13361,N_11040,N_11842);
or U13362 (N_13362,N_11075,N_11575);
nand U13363 (N_13363,N_10584,N_11360);
nor U13364 (N_13364,N_11483,N_11811);
and U13365 (N_13365,N_10888,N_10901);
nand U13366 (N_13366,N_10567,N_11275);
nand U13367 (N_13367,N_10627,N_10813);
and U13368 (N_13368,N_10543,N_11216);
nand U13369 (N_13369,N_11199,N_10815);
nor U13370 (N_13370,N_10709,N_11330);
xor U13371 (N_13371,N_11214,N_11765);
or U13372 (N_13372,N_11760,N_10961);
and U13373 (N_13373,N_11487,N_10899);
or U13374 (N_13374,N_11398,N_11620);
nand U13375 (N_13375,N_11809,N_11666);
nand U13376 (N_13376,N_11332,N_11509);
nor U13377 (N_13377,N_10898,N_11614);
nand U13378 (N_13378,N_10622,N_11094);
nor U13379 (N_13379,N_10822,N_11438);
xnor U13380 (N_13380,N_11454,N_11046);
and U13381 (N_13381,N_10786,N_11907);
nor U13382 (N_13382,N_10925,N_10965);
nor U13383 (N_13383,N_11482,N_11863);
or U13384 (N_13384,N_10627,N_11756);
and U13385 (N_13385,N_11882,N_11358);
or U13386 (N_13386,N_11653,N_11522);
nor U13387 (N_13387,N_10668,N_11960);
nand U13388 (N_13388,N_10725,N_10528);
xnor U13389 (N_13389,N_11920,N_11987);
and U13390 (N_13390,N_10514,N_11442);
nand U13391 (N_13391,N_11197,N_11852);
or U13392 (N_13392,N_11526,N_11862);
and U13393 (N_13393,N_11017,N_11871);
and U13394 (N_13394,N_11321,N_11422);
nand U13395 (N_13395,N_11369,N_11153);
nand U13396 (N_13396,N_11166,N_11320);
xor U13397 (N_13397,N_11525,N_11826);
xnor U13398 (N_13398,N_10940,N_10947);
or U13399 (N_13399,N_11504,N_11913);
or U13400 (N_13400,N_11634,N_11441);
nand U13401 (N_13401,N_11221,N_11725);
or U13402 (N_13402,N_11728,N_10949);
or U13403 (N_13403,N_11237,N_10986);
or U13404 (N_13404,N_11038,N_11906);
xor U13405 (N_13405,N_11941,N_10601);
or U13406 (N_13406,N_11606,N_11911);
and U13407 (N_13407,N_11545,N_10558);
or U13408 (N_13408,N_10746,N_10646);
or U13409 (N_13409,N_11708,N_11774);
nor U13410 (N_13410,N_10885,N_11219);
nor U13411 (N_13411,N_11212,N_11651);
or U13412 (N_13412,N_10824,N_11900);
nand U13413 (N_13413,N_11500,N_11628);
or U13414 (N_13414,N_11605,N_10782);
and U13415 (N_13415,N_11050,N_11196);
or U13416 (N_13416,N_11711,N_11487);
or U13417 (N_13417,N_11290,N_10566);
and U13418 (N_13418,N_11404,N_11585);
nand U13419 (N_13419,N_11310,N_11922);
or U13420 (N_13420,N_10508,N_11421);
and U13421 (N_13421,N_11379,N_11552);
nor U13422 (N_13422,N_11309,N_10918);
nand U13423 (N_13423,N_10850,N_10758);
and U13424 (N_13424,N_10913,N_10969);
and U13425 (N_13425,N_11128,N_11915);
or U13426 (N_13426,N_11294,N_10700);
nor U13427 (N_13427,N_11919,N_11750);
or U13428 (N_13428,N_11234,N_11059);
and U13429 (N_13429,N_10619,N_11727);
nand U13430 (N_13430,N_10513,N_11758);
and U13431 (N_13431,N_11850,N_10617);
or U13432 (N_13432,N_11554,N_11492);
nor U13433 (N_13433,N_11163,N_10667);
or U13434 (N_13434,N_10689,N_10820);
and U13435 (N_13435,N_11615,N_11734);
nor U13436 (N_13436,N_11122,N_11412);
nand U13437 (N_13437,N_10717,N_11861);
nand U13438 (N_13438,N_11056,N_11364);
nand U13439 (N_13439,N_10580,N_11788);
nand U13440 (N_13440,N_10879,N_11235);
or U13441 (N_13441,N_11366,N_11502);
nand U13442 (N_13442,N_10880,N_11631);
or U13443 (N_13443,N_11526,N_10655);
nand U13444 (N_13444,N_11193,N_10917);
or U13445 (N_13445,N_11463,N_11758);
or U13446 (N_13446,N_11313,N_11020);
nor U13447 (N_13447,N_10517,N_10782);
nor U13448 (N_13448,N_11572,N_11108);
nand U13449 (N_13449,N_11854,N_11057);
nor U13450 (N_13450,N_10797,N_11093);
or U13451 (N_13451,N_11116,N_11463);
nor U13452 (N_13452,N_10513,N_10618);
nand U13453 (N_13453,N_10647,N_11391);
nor U13454 (N_13454,N_10854,N_10702);
nand U13455 (N_13455,N_10669,N_11856);
or U13456 (N_13456,N_11403,N_11601);
or U13457 (N_13457,N_10579,N_11404);
nand U13458 (N_13458,N_11919,N_10684);
or U13459 (N_13459,N_11894,N_11266);
or U13460 (N_13460,N_11493,N_10692);
and U13461 (N_13461,N_11440,N_11837);
nand U13462 (N_13462,N_10783,N_11466);
xnor U13463 (N_13463,N_10845,N_10961);
nor U13464 (N_13464,N_11064,N_11067);
nor U13465 (N_13465,N_10644,N_10968);
nor U13466 (N_13466,N_11038,N_11971);
or U13467 (N_13467,N_11957,N_11784);
and U13468 (N_13468,N_11668,N_11773);
xor U13469 (N_13469,N_11737,N_11789);
nand U13470 (N_13470,N_10603,N_10979);
nand U13471 (N_13471,N_10610,N_11513);
nand U13472 (N_13472,N_11007,N_10720);
nand U13473 (N_13473,N_10796,N_11852);
nand U13474 (N_13474,N_11879,N_10985);
xor U13475 (N_13475,N_11624,N_10850);
and U13476 (N_13476,N_10808,N_11863);
or U13477 (N_13477,N_10803,N_10832);
nand U13478 (N_13478,N_11183,N_10852);
and U13479 (N_13479,N_11899,N_11619);
or U13480 (N_13480,N_10769,N_11429);
nand U13481 (N_13481,N_11673,N_11134);
or U13482 (N_13482,N_11171,N_11403);
or U13483 (N_13483,N_11947,N_10801);
nand U13484 (N_13484,N_10970,N_10974);
nor U13485 (N_13485,N_10641,N_10837);
nor U13486 (N_13486,N_11524,N_10702);
nor U13487 (N_13487,N_10700,N_11309);
xor U13488 (N_13488,N_11696,N_11610);
nor U13489 (N_13489,N_11177,N_11876);
and U13490 (N_13490,N_11366,N_10640);
nor U13491 (N_13491,N_11281,N_10813);
and U13492 (N_13492,N_11151,N_11173);
nor U13493 (N_13493,N_11183,N_11173);
or U13494 (N_13494,N_10960,N_10859);
nand U13495 (N_13495,N_11609,N_11799);
and U13496 (N_13496,N_11158,N_11841);
nor U13497 (N_13497,N_10824,N_10507);
and U13498 (N_13498,N_10932,N_10558);
xor U13499 (N_13499,N_11181,N_10668);
nor U13500 (N_13500,N_12929,N_13335);
nand U13501 (N_13501,N_12428,N_12959);
and U13502 (N_13502,N_12990,N_12489);
and U13503 (N_13503,N_12019,N_12739);
and U13504 (N_13504,N_12340,N_12993);
nor U13505 (N_13505,N_12385,N_13445);
and U13506 (N_13506,N_13333,N_13074);
or U13507 (N_13507,N_13196,N_13255);
nand U13508 (N_13508,N_12017,N_12774);
xnor U13509 (N_13509,N_12136,N_12087);
nand U13510 (N_13510,N_12764,N_12514);
nand U13511 (N_13511,N_13221,N_13262);
and U13512 (N_13512,N_13397,N_12826);
xor U13513 (N_13513,N_12072,N_13085);
or U13514 (N_13514,N_12734,N_12889);
nor U13515 (N_13515,N_13101,N_12838);
nand U13516 (N_13516,N_12283,N_12098);
xnor U13517 (N_13517,N_12078,N_13207);
nand U13518 (N_13518,N_13378,N_12462);
nor U13519 (N_13519,N_13171,N_13423);
nand U13520 (N_13520,N_12309,N_12789);
or U13521 (N_13521,N_12873,N_13156);
or U13522 (N_13522,N_12580,N_13016);
nor U13523 (N_13523,N_12595,N_12563);
and U13524 (N_13524,N_13341,N_12408);
or U13525 (N_13525,N_13012,N_13048);
xnor U13526 (N_13526,N_13417,N_12175);
and U13527 (N_13527,N_12241,N_12676);
and U13528 (N_13528,N_13244,N_12191);
and U13529 (N_13529,N_12083,N_12479);
or U13530 (N_13530,N_12026,N_12837);
nand U13531 (N_13531,N_12028,N_12797);
nor U13532 (N_13532,N_12937,N_12830);
nand U13533 (N_13533,N_12074,N_12402);
or U13534 (N_13534,N_12944,N_12605);
nand U13535 (N_13535,N_12742,N_13425);
and U13536 (N_13536,N_12575,N_12424);
nand U13537 (N_13537,N_13038,N_13226);
xor U13538 (N_13538,N_13322,N_13260);
and U13539 (N_13539,N_12427,N_12973);
nand U13540 (N_13540,N_12438,N_12051);
nor U13541 (N_13541,N_13302,N_12561);
nor U13542 (N_13542,N_12986,N_12354);
or U13543 (N_13543,N_12529,N_13309);
or U13544 (N_13544,N_12378,N_12669);
or U13545 (N_13545,N_13407,N_13312);
and U13546 (N_13546,N_12075,N_12685);
nor U13547 (N_13547,N_12750,N_12222);
nand U13548 (N_13548,N_13352,N_12598);
or U13549 (N_13549,N_12339,N_12876);
xor U13550 (N_13550,N_12433,N_12673);
nand U13551 (N_13551,N_12347,N_12371);
or U13552 (N_13552,N_12934,N_12457);
nand U13553 (N_13553,N_13144,N_13223);
or U13554 (N_13554,N_12955,N_12294);
nand U13555 (N_13555,N_12795,N_12059);
nor U13556 (N_13556,N_12054,N_12333);
nand U13557 (N_13557,N_13245,N_12148);
nor U13558 (N_13558,N_12454,N_12705);
or U13559 (N_13559,N_12202,N_12270);
nor U13560 (N_13560,N_12541,N_12288);
nand U13561 (N_13561,N_12056,N_13443);
or U13562 (N_13562,N_13096,N_12829);
nand U13563 (N_13563,N_13225,N_12055);
nand U13564 (N_13564,N_12966,N_12280);
nor U13565 (N_13565,N_12787,N_12981);
and U13566 (N_13566,N_12160,N_13284);
nand U13567 (N_13567,N_12694,N_12636);
nand U13568 (N_13568,N_12022,N_12802);
nor U13569 (N_13569,N_12994,N_13020);
or U13570 (N_13570,N_13203,N_12825);
and U13571 (N_13571,N_12084,N_12620);
or U13572 (N_13572,N_13356,N_13165);
or U13573 (N_13573,N_12883,N_13186);
and U13574 (N_13574,N_13305,N_12670);
nand U13575 (N_13575,N_12409,N_12388);
or U13576 (N_13576,N_12783,N_13167);
nor U13577 (N_13577,N_13436,N_13174);
nor U13578 (N_13578,N_13337,N_13396);
or U13579 (N_13579,N_12477,N_12183);
or U13580 (N_13580,N_12090,N_12284);
nor U13581 (N_13581,N_12046,N_12648);
or U13582 (N_13582,N_12027,N_13192);
and U13583 (N_13583,N_13442,N_12184);
nor U13584 (N_13584,N_13115,N_13209);
or U13585 (N_13585,N_13460,N_12237);
xnor U13586 (N_13586,N_13044,N_13040);
nor U13587 (N_13587,N_13150,N_12667);
or U13588 (N_13588,N_13433,N_13461);
nor U13589 (N_13589,N_13109,N_12156);
nor U13590 (N_13590,N_13348,N_12935);
nor U13591 (N_13591,N_12060,N_12145);
and U13592 (N_13592,N_12239,N_12258);
and U13593 (N_13593,N_12912,N_12749);
or U13594 (N_13594,N_12193,N_12520);
xnor U13595 (N_13595,N_13147,N_13298);
or U13596 (N_13596,N_12804,N_12296);
nand U13597 (N_13597,N_13440,N_12708);
and U13598 (N_13598,N_12821,N_13354);
nor U13599 (N_13599,N_12456,N_12586);
or U13600 (N_13600,N_12967,N_12257);
nor U13601 (N_13601,N_12686,N_12133);
nor U13602 (N_13602,N_12816,N_12422);
xnor U13603 (N_13603,N_12681,N_13353);
or U13604 (N_13604,N_12310,N_12482);
xor U13605 (N_13605,N_13202,N_12475);
nand U13606 (N_13606,N_13463,N_13416);
nor U13607 (N_13607,N_12800,N_12140);
nor U13608 (N_13608,N_12387,N_12707);
and U13609 (N_13609,N_12961,N_13492);
nand U13610 (N_13610,N_12608,N_13068);
nor U13611 (N_13611,N_12604,N_12397);
nand U13612 (N_13612,N_13448,N_12762);
and U13613 (N_13613,N_12557,N_12246);
nand U13614 (N_13614,N_12903,N_12556);
and U13615 (N_13615,N_12615,N_12177);
and U13616 (N_13616,N_12171,N_12814);
nor U13617 (N_13617,N_12358,N_12068);
or U13618 (N_13618,N_12813,N_12585);
and U13619 (N_13619,N_12793,N_12871);
nor U13620 (N_13620,N_13329,N_12139);
and U13621 (N_13621,N_12914,N_13213);
and U13622 (N_13622,N_13400,N_12303);
nand U13623 (N_13623,N_12911,N_12208);
nor U13624 (N_13624,N_12850,N_12500);
nand U13625 (N_13625,N_12539,N_13208);
nand U13626 (N_13626,N_12227,N_12516);
or U13627 (N_13627,N_12909,N_12497);
or U13628 (N_13628,N_12719,N_12809);
nor U13629 (N_13629,N_12581,N_13043);
or U13630 (N_13630,N_12647,N_13283);
xor U13631 (N_13631,N_13137,N_12213);
and U13632 (N_13632,N_12041,N_12508);
and U13633 (N_13633,N_12063,N_12755);
xnor U13634 (N_13634,N_12013,N_13266);
and U13635 (N_13635,N_13424,N_12253);
nand U13636 (N_13636,N_12852,N_12958);
or U13637 (N_13637,N_13494,N_13128);
nor U13638 (N_13638,N_12592,N_13268);
or U13639 (N_13639,N_13285,N_12070);
or U13640 (N_13640,N_12554,N_13472);
nand U13641 (N_13641,N_13406,N_13429);
nand U13642 (N_13642,N_13111,N_12372);
nand U13643 (N_13643,N_12437,N_12077);
nor U13644 (N_13644,N_13270,N_13452);
nor U13645 (N_13645,N_13130,N_12664);
or U13646 (N_13646,N_12741,N_12815);
or U13647 (N_13647,N_12025,N_13325);
nor U13648 (N_13648,N_12000,N_13166);
and U13649 (N_13649,N_13185,N_12528);
and U13650 (N_13650,N_13087,N_12638);
nand U13651 (N_13651,N_13491,N_12015);
or U13652 (N_13652,N_12609,N_12969);
xor U13653 (N_13653,N_13287,N_12375);
or U13654 (N_13654,N_13292,N_12550);
nand U13655 (N_13655,N_12064,N_13453);
or U13656 (N_13656,N_13133,N_12234);
or U13657 (N_13657,N_12709,N_12281);
or U13658 (N_13658,N_13269,N_13434);
or U13659 (N_13659,N_12440,N_13071);
and U13660 (N_13660,N_13141,N_12735);
nor U13661 (N_13661,N_12349,N_12405);
or U13662 (N_13662,N_13035,N_12185);
nand U13663 (N_13663,N_13172,N_12357);
or U13664 (N_13664,N_13490,N_13454);
and U13665 (N_13665,N_13427,N_13100);
and U13666 (N_13666,N_13409,N_13250);
xor U13667 (N_13667,N_12124,N_13475);
xor U13668 (N_13668,N_13449,N_13138);
and U13669 (N_13669,N_12492,N_12506);
or U13670 (N_13670,N_12522,N_12841);
nor U13671 (N_13671,N_13211,N_13008);
nor U13672 (N_13672,N_12590,N_13456);
nand U13673 (N_13673,N_12212,N_12461);
and U13674 (N_13674,N_12110,N_12355);
nand U13675 (N_13675,N_12524,N_12119);
nand U13676 (N_13676,N_12326,N_12768);
nor U13677 (N_13677,N_12302,N_12766);
and U13678 (N_13678,N_13464,N_12146);
nand U13679 (N_13679,N_12555,N_13224);
and U13680 (N_13680,N_12618,N_12147);
xnor U13681 (N_13681,N_13243,N_12373);
or U13682 (N_13682,N_13194,N_12786);
nor U13683 (N_13683,N_13170,N_12248);
nand U13684 (N_13684,N_12763,N_12938);
nand U13685 (N_13685,N_13098,N_12316);
nor U13686 (N_13686,N_12920,N_13009);
nor U13687 (N_13687,N_12361,N_12509);
nand U13688 (N_13688,N_12626,N_12352);
xnor U13689 (N_13689,N_13181,N_12268);
nand U13690 (N_13690,N_13272,N_13437);
nor U13691 (N_13691,N_12877,N_12058);
nor U13692 (N_13692,N_12105,N_12836);
nor U13693 (N_13693,N_12919,N_12259);
or U13694 (N_13694,N_12754,N_12570);
nor U13695 (N_13695,N_12215,N_12292);
nand U13696 (N_13696,N_13049,N_12818);
or U13697 (N_13697,N_13187,N_12382);
or U13698 (N_13698,N_12484,N_12229);
nand U13699 (N_13699,N_12896,N_12471);
or U13700 (N_13700,N_12782,N_12964);
nor U13701 (N_13701,N_12926,N_13139);
nor U13702 (N_13702,N_12891,N_12502);
or U13703 (N_13703,N_12526,N_13183);
nand U13704 (N_13704,N_12225,N_13360);
or U13705 (N_13705,N_12957,N_13466);
or U13706 (N_13706,N_13076,N_12855);
nand U13707 (N_13707,N_13383,N_13499);
xnor U13708 (N_13708,N_12666,N_13246);
xnor U13709 (N_13709,N_12389,N_12398);
nor U13710 (N_13710,N_12602,N_12984);
or U13711 (N_13711,N_12157,N_12857);
nor U13712 (N_13712,N_12899,N_12182);
nor U13713 (N_13713,N_12845,N_12571);
xnor U13714 (N_13714,N_12455,N_13294);
and U13715 (N_13715,N_13120,N_13343);
and U13716 (N_13716,N_13457,N_13247);
or U13717 (N_13717,N_13495,N_13164);
and U13718 (N_13718,N_12654,N_13386);
nand U13719 (N_13719,N_13034,N_12188);
and U13720 (N_13720,N_12429,N_13350);
or U13721 (N_13721,N_12662,N_12576);
xnor U13722 (N_13722,N_13162,N_12180);
or U13723 (N_13723,N_13249,N_12419);
nand U13724 (N_13724,N_12971,N_12822);
nor U13725 (N_13725,N_13093,N_13146);
or U13726 (N_13726,N_12819,N_12628);
and U13727 (N_13727,N_13042,N_13197);
nand U13728 (N_13728,N_12067,N_12487);
nand U13729 (N_13729,N_12478,N_12946);
or U13730 (N_13730,N_13389,N_13136);
and U13731 (N_13731,N_13411,N_13430);
or U13732 (N_13732,N_12210,N_12312);
nor U13733 (N_13733,N_13124,N_12173);
nand U13734 (N_13734,N_12179,N_12949);
nand U13735 (N_13735,N_13338,N_13019);
or U13736 (N_13736,N_12368,N_12345);
nand U13737 (N_13737,N_13073,N_12097);
and U13738 (N_13738,N_13403,N_13267);
nand U13739 (N_13739,N_13308,N_12359);
and U13740 (N_13740,N_12942,N_13301);
nand U13741 (N_13741,N_12341,N_12360);
nand U13742 (N_13742,N_13024,N_13095);
nand U13743 (N_13743,N_13496,N_12843);
and U13744 (N_13744,N_12204,N_13345);
nand U13745 (N_13745,N_12040,N_13013);
or U13746 (N_13746,N_12412,N_13288);
or U13747 (N_13747,N_12186,N_12413);
and U13748 (N_13748,N_12030,N_12863);
or U13749 (N_13749,N_13078,N_13401);
nand U13750 (N_13750,N_13127,N_12441);
nor U13751 (N_13751,N_13241,N_13478);
or U13752 (N_13752,N_12245,N_12727);
xor U13753 (N_13753,N_12176,N_13069);
or U13754 (N_13754,N_12925,N_13077);
nor U13755 (N_13755,N_12144,N_12167);
nor U13756 (N_13756,N_12610,N_12677);
nor U13757 (N_13757,N_13376,N_12260);
nand U13758 (N_13758,N_12726,N_12537);
and U13759 (N_13759,N_12223,N_12024);
or U13760 (N_13760,N_12542,N_12315);
or U13761 (N_13761,N_12458,N_13113);
nand U13762 (N_13762,N_12982,N_12323);
or U13763 (N_13763,N_12614,N_13210);
nor U13764 (N_13764,N_12760,N_13498);
nand U13765 (N_13765,N_13182,N_12747);
xnor U13766 (N_13766,N_12624,N_13015);
and U13767 (N_13767,N_12699,N_12111);
or U13768 (N_13768,N_12893,N_12640);
nor U13769 (N_13769,N_13045,N_12189);
nor U13770 (N_13770,N_12279,N_12639);
or U13771 (N_13771,N_13118,N_13299);
or U13772 (N_13772,N_12864,N_13307);
nand U13773 (N_13773,N_13296,N_12470);
nand U13774 (N_13774,N_12701,N_13029);
xor U13775 (N_13775,N_13289,N_12807);
and U13776 (N_13776,N_12534,N_12518);
nand U13777 (N_13777,N_13334,N_13198);
nor U13778 (N_13778,N_12770,N_13094);
nor U13779 (N_13779,N_12858,N_13479);
nand U13780 (N_13780,N_12660,N_12803);
nand U13781 (N_13781,N_12558,N_12692);
and U13782 (N_13782,N_13254,N_13017);
xnor U13783 (N_13783,N_12383,N_12684);
and U13784 (N_13784,N_13158,N_12289);
or U13785 (N_13785,N_12379,N_12621);
and U13786 (N_13786,N_13143,N_12794);
or U13787 (N_13787,N_12351,N_13263);
nor U13788 (N_13788,N_13340,N_12295);
or U13789 (N_13789,N_12715,N_12560);
or U13790 (N_13790,N_12645,N_12898);
nand U13791 (N_13791,N_13151,N_13199);
nand U13792 (N_13792,N_12443,N_12103);
and U13793 (N_13793,N_13253,N_13107);
nor U13794 (N_13794,N_12150,N_12082);
and U13795 (N_13795,N_12474,N_13030);
nor U13796 (N_13796,N_12014,N_12356);
xnor U13797 (N_13797,N_13276,N_12431);
and U13798 (N_13798,N_12153,N_12512);
or U13799 (N_13799,N_13233,N_12329);
and U13800 (N_13800,N_12525,N_12037);
or U13801 (N_13801,N_12406,N_13374);
nor U13802 (N_13802,N_12653,N_12988);
or U13803 (N_13803,N_12744,N_12214);
nand U13804 (N_13804,N_12828,N_12767);
nand U13805 (N_13805,N_13324,N_12266);
and U13806 (N_13806,N_12276,N_12697);
nor U13807 (N_13807,N_12038,N_13470);
and U13808 (N_13808,N_12820,N_12086);
and U13809 (N_13809,N_12285,N_13175);
and U13810 (N_13810,N_13311,N_12343);
nand U13811 (N_13811,N_12833,N_12317);
nand U13812 (N_13812,N_12721,N_12886);
or U13813 (N_13813,N_13300,N_13372);
and U13814 (N_13814,N_12076,N_13195);
nor U13815 (N_13815,N_12094,N_12112);
and U13816 (N_13816,N_13359,N_13149);
nor U13817 (N_13817,N_12880,N_12890);
or U13818 (N_13818,N_12466,N_12495);
or U13819 (N_13819,N_12272,N_12313);
and U13820 (N_13820,N_12009,N_13026);
and U13821 (N_13821,N_12254,N_12761);
nor U13822 (N_13822,N_12467,N_13435);
and U13823 (N_13823,N_12932,N_13327);
or U13824 (N_13824,N_13082,N_13191);
or U13825 (N_13825,N_12567,N_12305);
nor U13826 (N_13826,N_13483,N_12631);
nor U13827 (N_13827,N_13316,N_12835);
xor U13828 (N_13828,N_12120,N_12562);
nor U13829 (N_13829,N_12123,N_12531);
nor U13830 (N_13830,N_12100,N_13297);
xnor U13831 (N_13831,N_12021,N_12998);
nand U13832 (N_13832,N_13381,N_12551);
and U13833 (N_13833,N_12847,N_13471);
or U13834 (N_13834,N_12092,N_12436);
nand U13835 (N_13835,N_13368,N_13375);
xnor U13836 (N_13836,N_12217,N_12970);
or U13837 (N_13837,N_12972,N_12665);
or U13838 (N_13838,N_12733,N_13215);
or U13839 (N_13839,N_12849,N_13361);
nor U13840 (N_13840,N_12299,N_12334);
nor U13841 (N_13841,N_13025,N_13488);
nand U13842 (N_13842,N_12403,N_12776);
or U13843 (N_13843,N_12933,N_12447);
or U13844 (N_13844,N_12104,N_12872);
and U13845 (N_13845,N_12348,N_12163);
or U13846 (N_13846,N_13135,N_12494);
nor U13847 (N_13847,N_12805,N_12897);
nand U13848 (N_13848,N_12706,N_12549);
and U13849 (N_13849,N_12772,N_13291);
or U13850 (N_13850,N_12095,N_12485);
and U13851 (N_13851,N_12751,N_12195);
nor U13852 (N_13852,N_13455,N_13132);
nor U13853 (N_13853,N_13286,N_13477);
and U13854 (N_13854,N_13336,N_12012);
nor U13855 (N_13855,N_12577,N_12391);
xnor U13856 (N_13856,N_13066,N_12113);
xor U13857 (N_13857,N_12724,N_12251);
nand U13858 (N_13858,N_13328,N_13265);
nor U13859 (N_13859,N_12381,N_13205);
or U13860 (N_13860,N_12158,N_12996);
nand U13861 (N_13861,N_12756,N_12769);
nor U13862 (N_13862,N_12736,N_12565);
nor U13863 (N_13863,N_12507,N_12612);
nand U13864 (N_13864,N_12364,N_12318);
and U13865 (N_13865,N_13154,N_12510);
nand U13866 (N_13866,N_13256,N_12960);
or U13867 (N_13867,N_12196,N_13160);
and U13868 (N_13868,N_12350,N_12481);
nor U13869 (N_13869,N_12106,N_12216);
xor U13870 (N_13870,N_12892,N_13168);
nand U13871 (N_13871,N_13273,N_12298);
nand U13872 (N_13872,N_13102,N_12201);
nand U13873 (N_13873,N_12366,N_12005);
and U13874 (N_13874,N_12704,N_12301);
nor U13875 (N_13875,N_13419,N_13331);
or U13876 (N_13876,N_12152,N_12211);
and U13877 (N_13877,N_12533,N_12472);
and U13878 (N_13878,N_13121,N_12989);
or U13879 (N_13879,N_12796,N_13306);
nand U13880 (N_13880,N_13067,N_12226);
nand U13881 (N_13881,N_12047,N_13036);
and U13882 (N_13882,N_12799,N_12320);
nand U13883 (N_13883,N_12032,N_13362);
nand U13884 (N_13884,N_12080,N_12194);
or U13885 (N_13885,N_12716,N_13380);
nand U13886 (N_13886,N_12941,N_13486);
nor U13887 (N_13887,N_12035,N_12328);
and U13888 (N_13888,N_13476,N_12342);
and U13889 (N_13889,N_12808,N_13371);
xor U13890 (N_13890,N_13410,N_13326);
or U13891 (N_13891,N_12728,N_12093);
nor U13892 (N_13892,N_12962,N_12931);
nand U13893 (N_13893,N_13467,N_12780);
nor U13894 (N_13894,N_13161,N_12633);
or U13895 (N_13895,N_13450,N_12231);
nand U13896 (N_13896,N_12865,N_13114);
nor U13897 (N_13897,N_13365,N_12033);
nand U13898 (N_13898,N_12170,N_12250);
or U13899 (N_13899,N_13317,N_12307);
or U13900 (N_13900,N_12731,N_12940);
nand U13901 (N_13901,N_12757,N_12582);
or U13902 (N_13902,N_12505,N_13408);
nand U13903 (N_13903,N_12922,N_12066);
nand U13904 (N_13904,N_13028,N_12114);
and U13905 (N_13905,N_13023,N_12134);
xor U13906 (N_13906,N_12752,N_12668);
nand U13907 (N_13907,N_13364,N_13257);
nand U13908 (N_13908,N_12753,N_12846);
or U13909 (N_13909,N_13458,N_13055);
nor U13910 (N_13910,N_13119,N_12882);
or U13911 (N_13911,N_13480,N_12221);
and U13912 (N_13912,N_12209,N_13485);
and U13913 (N_13913,N_12943,N_13145);
nor U13914 (N_13914,N_12930,N_12162);
nand U13915 (N_13915,N_12597,N_12995);
and U13916 (N_13916,N_13056,N_12240);
xnor U13917 (N_13917,N_12695,N_13431);
nand U13918 (N_13918,N_12135,N_12978);
or U13919 (N_13919,N_12236,N_12997);
and U13920 (N_13920,N_12801,N_13219);
xnor U13921 (N_13921,N_12884,N_12448);
or U13922 (N_13922,N_12523,N_12513);
nor U13923 (N_13923,N_12778,N_12252);
xor U13924 (N_13924,N_12566,N_13259);
nor U13925 (N_13925,N_13384,N_12218);
nor U13926 (N_13926,N_12601,N_12324);
nand U13927 (N_13927,N_13193,N_12274);
nand U13928 (N_13928,N_12939,N_12517);
or U13929 (N_13929,N_12564,N_12255);
xnor U13930 (N_13930,N_13062,N_13080);
nor U13931 (N_13931,N_12854,N_12203);
and U13932 (N_13932,N_12434,N_12738);
nand U13933 (N_13933,N_12418,N_12860);
nand U13934 (N_13934,N_12853,N_12362);
or U13935 (N_13935,N_13293,N_13451);
or U13936 (N_13936,N_12411,N_12444);
or U13937 (N_13937,N_12369,N_12057);
nor U13938 (N_13938,N_12219,N_12344);
nor U13939 (N_13939,N_12975,N_12016);
nor U13940 (N_13940,N_12449,N_12875);
or U13941 (N_13941,N_12616,N_12792);
nand U13942 (N_13942,N_13321,N_13057);
or U13943 (N_13943,N_12979,N_12593);
nand U13944 (N_13944,N_12401,N_12546);
nor U13945 (N_13945,N_13465,N_12242);
and U13946 (N_13946,N_12839,N_13358);
nor U13947 (N_13947,N_13280,N_12483);
or U13948 (N_13948,N_12445,N_12174);
and U13949 (N_13949,N_12325,N_12088);
or U13950 (N_13950,N_13385,N_13125);
or U13951 (N_13951,N_13278,N_12954);
or U13952 (N_13952,N_12126,N_12758);
and U13953 (N_13953,N_12712,N_12798);
nor U13954 (N_13954,N_12453,N_12337);
or U13955 (N_13955,N_12023,N_12936);
nand U13956 (N_13956,N_12420,N_13279);
or U13957 (N_13957,N_13319,N_12096);
and U13958 (N_13958,N_13104,N_12062);
nand U13959 (N_13959,N_12894,N_12553);
or U13960 (N_13960,N_12907,N_12137);
nand U13961 (N_13961,N_12029,N_12691);
and U13962 (N_13962,N_12034,N_12273);
and U13963 (N_13963,N_12407,N_12637);
or U13964 (N_13964,N_13126,N_13313);
nand U13965 (N_13965,N_13060,N_12071);
and U13966 (N_13966,N_12777,N_13002);
nor U13967 (N_13967,N_12233,N_12459);
xnor U13968 (N_13968,N_12569,N_13347);
and U13969 (N_13969,N_12790,N_12568);
nand U13970 (N_13970,N_13075,N_12806);
or U13971 (N_13971,N_12746,N_12031);
or U13972 (N_13972,N_12504,N_12149);
xor U13973 (N_13973,N_13474,N_13152);
nor U13974 (N_13974,N_13447,N_12322);
nand U13975 (N_13975,N_12414,N_12039);
and U13976 (N_13976,N_12991,N_12644);
nor U13977 (N_13977,N_13370,N_13373);
or U13978 (N_13978,N_13123,N_12651);
or U13979 (N_13979,N_13081,N_12390);
nor U13980 (N_13980,N_13050,N_12924);
nor U13981 (N_13981,N_12151,N_13180);
nor U13982 (N_13982,N_13421,N_13088);
nand U13983 (N_13983,N_13462,N_12338);
nor U13984 (N_13984,N_12468,N_12916);
nand U13985 (N_13985,N_12655,N_13155);
and U13986 (N_13986,N_12910,N_13404);
and U13987 (N_13987,N_12396,N_13179);
nand U13988 (N_13988,N_12658,N_12611);
xnor U13989 (N_13989,N_13058,N_13320);
and U13990 (N_13990,N_12974,N_12885);
or U13991 (N_13991,N_13281,N_13234);
nand U13992 (N_13992,N_13242,N_13415);
or U13993 (N_13993,N_12044,N_13201);
xor U13994 (N_13994,N_12951,N_13148);
and U13995 (N_13995,N_12109,N_12154);
nor U13996 (N_13996,N_12464,N_13190);
and U13997 (N_13997,N_12824,N_13304);
and U13998 (N_13998,N_12143,N_12125);
nor U13999 (N_13999,N_13391,N_12649);
nand U14000 (N_14000,N_12713,N_13059);
nand U14001 (N_14001,N_12107,N_12331);
or U14002 (N_14002,N_13252,N_12859);
nor U14003 (N_14003,N_13099,N_13212);
and U14004 (N_14004,N_12410,N_13332);
and U14005 (N_14005,N_12129,N_12450);
nand U14006 (N_14006,N_13173,N_12061);
or U14007 (N_14007,N_12574,N_12486);
and U14008 (N_14008,N_12048,N_12834);
nand U14009 (N_14009,N_13007,N_12392);
xor U14010 (N_14010,N_12547,N_12386);
nand U14011 (N_14011,N_13037,N_12050);
or U14012 (N_14012,N_12395,N_12130);
xor U14013 (N_14013,N_13047,N_12629);
and U14014 (N_14014,N_12052,N_13072);
and U14015 (N_14015,N_13006,N_12915);
xnor U14016 (N_14016,N_13222,N_13387);
and U14017 (N_14017,N_13200,N_13097);
nor U14018 (N_14018,N_12085,N_12627);
or U14019 (N_14019,N_13163,N_12900);
nand U14020 (N_14020,N_12927,N_12244);
nand U14021 (N_14021,N_12263,N_12588);
and U14022 (N_14022,N_12155,N_12099);
nor U14023 (N_14023,N_12043,N_13277);
nor U14024 (N_14024,N_12945,N_12635);
and U14025 (N_14025,N_12172,N_12142);
and U14026 (N_14026,N_13303,N_13232);
nand U14027 (N_14027,N_12874,N_12878);
nor U14028 (N_14028,N_12536,N_12122);
xor U14029 (N_14029,N_12327,N_12277);
or U14030 (N_14030,N_12164,N_13178);
and U14031 (N_14031,N_13402,N_12131);
nor U14032 (N_14032,N_12073,N_12404);
nand U14033 (N_14033,N_12901,N_12527);
nor U14034 (N_14034,N_13070,N_12121);
nand U14035 (N_14035,N_12652,N_13344);
nand U14036 (N_14036,N_13004,N_12178);
or U14037 (N_14037,N_13129,N_13351);
nor U14038 (N_14038,N_12473,N_12451);
or U14039 (N_14039,N_12346,N_12690);
and U14040 (N_14040,N_12007,N_13240);
nand U14041 (N_14041,N_12700,N_12895);
or U14042 (N_14042,N_13206,N_12249);
xor U14043 (N_14043,N_12535,N_12425);
and U14044 (N_14044,N_13388,N_13134);
and U14045 (N_14045,N_13122,N_12165);
nand U14046 (N_14046,N_13227,N_12321);
nor U14047 (N_14047,N_13177,N_13230);
or U14048 (N_14048,N_12623,N_12696);
or U14049 (N_14049,N_12374,N_12603);
or U14050 (N_14050,N_12049,N_13063);
nand U14051 (N_14051,N_12332,N_12247);
nor U14052 (N_14052,N_12319,N_12663);
nand U14053 (N_14053,N_12659,N_12267);
nand U14054 (N_14054,N_13339,N_12490);
xnor U14055 (N_14055,N_13001,N_12788);
and U14056 (N_14056,N_12856,N_12725);
and U14057 (N_14057,N_12619,N_13248);
and U14058 (N_14058,N_12235,N_12169);
and U14059 (N_14059,N_12573,N_12906);
nand U14060 (N_14060,N_13412,N_12674);
nor U14061 (N_14061,N_12544,N_13418);
nand U14062 (N_14062,N_12519,N_12844);
and U14063 (N_14063,N_12717,N_12282);
and U14064 (N_14064,N_12224,N_13011);
nand U14065 (N_14065,N_12465,N_12679);
nand U14066 (N_14066,N_12187,N_13346);
and U14067 (N_14067,N_13112,N_13000);
nor U14068 (N_14068,N_13239,N_12559);
nand U14069 (N_14069,N_12496,N_12773);
nor U14070 (N_14070,N_12748,N_13110);
nor U14071 (N_14071,N_12521,N_12928);
nor U14072 (N_14072,N_12290,N_12232);
xnor U14073 (N_14073,N_12887,N_12308);
nor U14074 (N_14074,N_12421,N_12908);
nand U14075 (N_14075,N_12269,N_12643);
or U14076 (N_14076,N_13382,N_12197);
or U14077 (N_14077,N_13189,N_12950);
nand U14078 (N_14078,N_13444,N_13493);
and U14079 (N_14079,N_12740,N_13349);
xnor U14080 (N_14080,N_13214,N_12415);
or U14081 (N_14081,N_12622,N_12399);
or U14082 (N_14082,N_12384,N_13229);
and U14083 (N_14083,N_13083,N_12881);
nor U14084 (N_14084,N_12842,N_12702);
nand U14085 (N_14085,N_13315,N_13395);
or U14086 (N_14086,N_12287,N_12488);
or U14087 (N_14087,N_12400,N_13184);
nand U14088 (N_14088,N_13422,N_12300);
nand U14089 (N_14089,N_12599,N_12530);
xnor U14090 (N_14090,N_13218,N_12613);
or U14091 (N_14091,N_12956,N_12493);
or U14092 (N_14092,N_12036,N_13032);
and U14093 (N_14093,N_13188,N_12671);
nand U14094 (N_14094,N_13484,N_12192);
nand U14095 (N_14095,N_12646,N_12661);
nand U14096 (N_14096,N_13489,N_12784);
nor U14097 (N_14097,N_12293,N_12118);
nor U14098 (N_14098,N_13231,N_12718);
nand U14099 (N_14099,N_13216,N_12190);
nand U14100 (N_14100,N_12460,N_12584);
nor U14101 (N_14101,N_13392,N_13399);
nor U14102 (N_14102,N_12683,N_13090);
and U14103 (N_14103,N_13027,N_12335);
nor U14104 (N_14104,N_12869,N_12963);
nor U14105 (N_14105,N_12917,N_12480);
and U14106 (N_14106,N_13367,N_12168);
nand U14107 (N_14107,N_12128,N_12866);
xor U14108 (N_14108,N_12442,N_13169);
and U14109 (N_14109,N_12579,N_12003);
nor U14110 (N_14110,N_12423,N_12840);
nand U14111 (N_14111,N_12377,N_13405);
or U14112 (N_14112,N_12430,N_13393);
nor U14113 (N_14113,N_13459,N_12548);
or U14114 (N_14114,N_12132,N_12089);
nand U14115 (N_14115,N_12722,N_12688);
nor U14116 (N_14116,N_12261,N_12115);
nand U14117 (N_14117,N_12256,N_13275);
or U14118 (N_14118,N_13379,N_13238);
or U14119 (N_14119,N_12775,N_12968);
and U14120 (N_14120,N_13441,N_12687);
or U14121 (N_14121,N_13022,N_12004);
or U14122 (N_14122,N_13159,N_13236);
or U14123 (N_14123,N_13005,N_13432);
nor U14124 (N_14124,N_12265,N_12511);
and U14125 (N_14125,N_12977,N_13426);
or U14126 (N_14126,N_12116,N_12714);
or U14127 (N_14127,N_13394,N_13377);
nor U14128 (N_14128,N_12617,N_12286);
or U14129 (N_14129,N_13366,N_13258);
or U14130 (N_14130,N_13217,N_13108);
or U14131 (N_14131,N_12730,N_12330);
or U14132 (N_14132,N_12435,N_12069);
nor U14133 (N_14133,N_12020,N_12607);
xor U14134 (N_14134,N_13204,N_12867);
and U14135 (N_14135,N_12630,N_13117);
nand U14136 (N_14136,N_12091,N_13251);
nor U14137 (N_14137,N_12503,N_12642);
and U14138 (N_14138,N_13264,N_13271);
nor U14139 (N_14139,N_12540,N_12002);
and U14140 (N_14140,N_12306,N_13235);
or U14141 (N_14141,N_13355,N_12304);
and U14142 (N_14142,N_13086,N_13310);
or U14143 (N_14143,N_12376,N_12992);
or U14144 (N_14144,N_12297,N_12823);
or U14145 (N_14145,N_12948,N_12275);
or U14146 (N_14146,N_12811,N_13323);
nor U14147 (N_14147,N_12220,N_12965);
and U14148 (N_14148,N_13021,N_13220);
or U14149 (N_14149,N_13469,N_13084);
nand U14150 (N_14150,N_13330,N_13342);
and U14151 (N_14151,N_12181,N_13438);
and U14152 (N_14152,N_13092,N_12710);
nand U14153 (N_14153,N_12827,N_12732);
or U14154 (N_14154,N_12680,N_12678);
and U14155 (N_14155,N_12606,N_12625);
or U14156 (N_14156,N_12001,N_12765);
nor U14157 (N_14157,N_12947,N_12426);
or U14158 (N_14158,N_12779,N_12672);
and U14159 (N_14159,N_12238,N_13140);
xnor U14160 (N_14160,N_13282,N_12501);
nor U14161 (N_14161,N_12812,N_12952);
and U14162 (N_14162,N_12264,N_12532);
nor U14163 (N_14163,N_12499,N_13468);
nand U14164 (N_14164,N_12861,N_12737);
nor U14165 (N_14165,N_13079,N_12656);
nor U14166 (N_14166,N_12831,N_12980);
nand U14167 (N_14167,N_12987,N_12745);
or U14168 (N_14168,N_12353,N_13103);
and U14169 (N_14169,N_12311,N_13106);
and U14170 (N_14170,N_13295,N_12953);
nand U14171 (N_14171,N_13054,N_13116);
nand U14172 (N_14172,N_12291,N_12689);
nor U14173 (N_14173,N_13039,N_13065);
or U14174 (N_14174,N_12600,N_12729);
nand U14175 (N_14175,N_12228,N_12166);
xnor U14176 (N_14176,N_12278,N_12634);
nand U14177 (N_14177,N_12081,N_13237);
nand U14178 (N_14178,N_12650,N_12583);
nand U14179 (N_14179,N_12079,N_13010);
and U14180 (N_14180,N_12921,N_12198);
nand U14181 (N_14181,N_12791,N_12785);
or U14182 (N_14182,N_12703,N_12446);
nor U14183 (N_14183,N_12552,N_13089);
nor U14184 (N_14184,N_13153,N_13290);
xor U14185 (N_14185,N_12578,N_12810);
or U14186 (N_14186,N_12008,N_12879);
nor U14187 (N_14187,N_12983,N_12589);
xnor U14188 (N_14188,N_13031,N_12498);
nand U14189 (N_14189,N_12596,N_12675);
nor U14190 (N_14190,N_12271,N_12045);
or U14191 (N_14191,N_12452,N_12011);
and U14192 (N_14192,N_12380,N_13041);
and U14193 (N_14193,N_12018,N_13033);
or U14194 (N_14194,N_13369,N_12851);
or U14195 (N_14195,N_12416,N_12759);
xor U14196 (N_14196,N_12587,N_13318);
nor U14197 (N_14197,N_12417,N_12367);
and U14198 (N_14198,N_13481,N_12682);
or U14199 (N_14199,N_12632,N_13420);
xor U14200 (N_14200,N_13064,N_13439);
nor U14201 (N_14201,N_12053,N_13390);
and U14202 (N_14202,N_12711,N_12127);
or U14203 (N_14203,N_12870,N_12010);
nor U14204 (N_14204,N_12976,N_12363);
and U14205 (N_14205,N_12545,N_12904);
and U14206 (N_14206,N_12262,N_12572);
nor U14207 (N_14207,N_12199,N_12006);
nor U14208 (N_14208,N_12230,N_12723);
nand U14209 (N_14209,N_13091,N_12161);
nor U14210 (N_14210,N_12515,N_12594);
nor U14211 (N_14211,N_12463,N_13228);
nand U14212 (N_14212,N_12817,N_13053);
and U14213 (N_14213,N_12207,N_12476);
nor U14214 (N_14214,N_13497,N_12985);
nor U14215 (N_14215,N_12913,N_12918);
and U14216 (N_14216,N_13473,N_12469);
nor U14217 (N_14217,N_12432,N_12862);
xnor U14218 (N_14218,N_13261,N_12108);
nor U14219 (N_14219,N_12693,N_12117);
and U14220 (N_14220,N_12159,N_13157);
or U14221 (N_14221,N_13487,N_12491);
nand U14222 (N_14222,N_12141,N_13061);
nand U14223 (N_14223,N_12042,N_12138);
nor U14224 (N_14224,N_12370,N_13046);
nand U14225 (N_14225,N_13176,N_12641);
and U14226 (N_14226,N_12243,N_13428);
xor U14227 (N_14227,N_12771,N_13357);
or U14228 (N_14228,N_13414,N_13398);
or U14229 (N_14229,N_12543,N_12888);
nand U14230 (N_14230,N_12205,N_12439);
nor U14231 (N_14231,N_13274,N_12905);
nand U14232 (N_14232,N_13051,N_13363);
nor U14233 (N_14233,N_12102,N_13314);
xnor U14234 (N_14234,N_12538,N_13003);
or U14235 (N_14235,N_12832,N_13413);
or U14236 (N_14236,N_13446,N_13018);
and U14237 (N_14237,N_12999,N_13131);
nor U14238 (N_14238,N_12868,N_12848);
and U14239 (N_14239,N_13105,N_13142);
nor U14240 (N_14240,N_12065,N_12720);
and U14241 (N_14241,N_12206,N_12591);
xnor U14242 (N_14242,N_13014,N_12923);
or U14243 (N_14243,N_12101,N_12743);
and U14244 (N_14244,N_12698,N_13482);
nor U14245 (N_14245,N_12365,N_12393);
and U14246 (N_14246,N_12902,N_12314);
or U14247 (N_14247,N_12200,N_13052);
and U14248 (N_14248,N_12781,N_12336);
nand U14249 (N_14249,N_12394,N_12657);
and U14250 (N_14250,N_12274,N_13449);
nor U14251 (N_14251,N_12576,N_13104);
or U14252 (N_14252,N_12275,N_12995);
xor U14253 (N_14253,N_12921,N_12356);
xnor U14254 (N_14254,N_13054,N_13327);
nor U14255 (N_14255,N_12939,N_12312);
or U14256 (N_14256,N_12232,N_13135);
xnor U14257 (N_14257,N_12171,N_13004);
nand U14258 (N_14258,N_12686,N_12597);
nand U14259 (N_14259,N_13178,N_13086);
nor U14260 (N_14260,N_13267,N_13146);
nor U14261 (N_14261,N_12193,N_12873);
or U14262 (N_14262,N_12239,N_12291);
or U14263 (N_14263,N_13017,N_12136);
xnor U14264 (N_14264,N_12198,N_12344);
nor U14265 (N_14265,N_12155,N_12279);
and U14266 (N_14266,N_12460,N_13133);
xnor U14267 (N_14267,N_13457,N_13113);
xnor U14268 (N_14268,N_12700,N_12819);
and U14269 (N_14269,N_12569,N_13222);
or U14270 (N_14270,N_12382,N_13414);
nand U14271 (N_14271,N_12874,N_12407);
nand U14272 (N_14272,N_13098,N_12124);
nand U14273 (N_14273,N_13474,N_12157);
and U14274 (N_14274,N_12305,N_12186);
nand U14275 (N_14275,N_13128,N_12953);
and U14276 (N_14276,N_12399,N_12076);
or U14277 (N_14277,N_13338,N_12095);
nand U14278 (N_14278,N_12895,N_13037);
or U14279 (N_14279,N_12827,N_12259);
and U14280 (N_14280,N_12780,N_13136);
and U14281 (N_14281,N_13496,N_12705);
and U14282 (N_14282,N_13139,N_12431);
or U14283 (N_14283,N_12758,N_12669);
xor U14284 (N_14284,N_12896,N_12381);
or U14285 (N_14285,N_12320,N_13216);
nor U14286 (N_14286,N_12365,N_13042);
nand U14287 (N_14287,N_12667,N_12731);
or U14288 (N_14288,N_12157,N_12984);
and U14289 (N_14289,N_13358,N_12216);
nor U14290 (N_14290,N_13486,N_13321);
and U14291 (N_14291,N_12476,N_12270);
and U14292 (N_14292,N_12052,N_12210);
nand U14293 (N_14293,N_12408,N_12565);
nand U14294 (N_14294,N_13200,N_12103);
and U14295 (N_14295,N_13471,N_13210);
nor U14296 (N_14296,N_12219,N_12204);
or U14297 (N_14297,N_12830,N_12960);
nand U14298 (N_14298,N_12850,N_12231);
and U14299 (N_14299,N_12790,N_12314);
or U14300 (N_14300,N_13170,N_12559);
nor U14301 (N_14301,N_12909,N_12920);
xnor U14302 (N_14302,N_12578,N_12580);
or U14303 (N_14303,N_12831,N_12948);
nand U14304 (N_14304,N_13043,N_12197);
nand U14305 (N_14305,N_12460,N_12476);
xnor U14306 (N_14306,N_12475,N_12418);
and U14307 (N_14307,N_12332,N_13082);
xor U14308 (N_14308,N_13025,N_12750);
nor U14309 (N_14309,N_12257,N_12788);
nand U14310 (N_14310,N_12752,N_12489);
and U14311 (N_14311,N_13377,N_12458);
nor U14312 (N_14312,N_13173,N_13264);
and U14313 (N_14313,N_12185,N_12152);
or U14314 (N_14314,N_12059,N_12697);
or U14315 (N_14315,N_12254,N_12033);
xnor U14316 (N_14316,N_12410,N_12166);
xnor U14317 (N_14317,N_12735,N_13123);
nor U14318 (N_14318,N_12818,N_13008);
or U14319 (N_14319,N_12842,N_13099);
nor U14320 (N_14320,N_13325,N_12102);
and U14321 (N_14321,N_13047,N_12364);
xnor U14322 (N_14322,N_12859,N_12014);
and U14323 (N_14323,N_12730,N_12549);
nand U14324 (N_14324,N_13307,N_13397);
and U14325 (N_14325,N_12589,N_12509);
or U14326 (N_14326,N_12013,N_12214);
or U14327 (N_14327,N_13399,N_13286);
or U14328 (N_14328,N_13198,N_13131);
or U14329 (N_14329,N_13252,N_12417);
nand U14330 (N_14330,N_12144,N_12114);
and U14331 (N_14331,N_13256,N_13062);
nor U14332 (N_14332,N_13089,N_13420);
or U14333 (N_14333,N_12201,N_12587);
or U14334 (N_14334,N_13292,N_13341);
xnor U14335 (N_14335,N_12841,N_12014);
xnor U14336 (N_14336,N_12505,N_12687);
nor U14337 (N_14337,N_12706,N_13168);
nand U14338 (N_14338,N_13354,N_12806);
or U14339 (N_14339,N_13342,N_12469);
nand U14340 (N_14340,N_12388,N_12973);
nand U14341 (N_14341,N_13104,N_12906);
and U14342 (N_14342,N_12254,N_12385);
and U14343 (N_14343,N_12281,N_12886);
nand U14344 (N_14344,N_13358,N_13021);
and U14345 (N_14345,N_12380,N_12226);
nor U14346 (N_14346,N_12015,N_12857);
and U14347 (N_14347,N_12527,N_13255);
nand U14348 (N_14348,N_12697,N_13227);
nand U14349 (N_14349,N_12066,N_12026);
or U14350 (N_14350,N_13065,N_13189);
nor U14351 (N_14351,N_13320,N_13011);
and U14352 (N_14352,N_12868,N_13035);
and U14353 (N_14353,N_12624,N_12827);
nand U14354 (N_14354,N_12778,N_12333);
or U14355 (N_14355,N_12824,N_12942);
nor U14356 (N_14356,N_12712,N_13431);
and U14357 (N_14357,N_13451,N_12089);
or U14358 (N_14358,N_12681,N_12382);
nand U14359 (N_14359,N_12147,N_12200);
xnor U14360 (N_14360,N_12937,N_12172);
nor U14361 (N_14361,N_12881,N_13326);
or U14362 (N_14362,N_12646,N_13183);
nand U14363 (N_14363,N_12626,N_12345);
xnor U14364 (N_14364,N_12844,N_12773);
nor U14365 (N_14365,N_12364,N_12834);
and U14366 (N_14366,N_13046,N_12748);
nand U14367 (N_14367,N_12041,N_12308);
nand U14368 (N_14368,N_13205,N_13035);
nor U14369 (N_14369,N_12468,N_13361);
xnor U14370 (N_14370,N_12448,N_12941);
xor U14371 (N_14371,N_12597,N_12539);
nor U14372 (N_14372,N_12018,N_12445);
nand U14373 (N_14373,N_12319,N_12966);
or U14374 (N_14374,N_12487,N_12486);
and U14375 (N_14375,N_13406,N_12009);
nor U14376 (N_14376,N_12560,N_13022);
nor U14377 (N_14377,N_12074,N_12051);
and U14378 (N_14378,N_13465,N_13089);
nand U14379 (N_14379,N_12983,N_13202);
xnor U14380 (N_14380,N_12538,N_13275);
nand U14381 (N_14381,N_12344,N_12610);
xor U14382 (N_14382,N_12885,N_13372);
nor U14383 (N_14383,N_13112,N_12843);
and U14384 (N_14384,N_13332,N_13212);
nand U14385 (N_14385,N_12213,N_12541);
nor U14386 (N_14386,N_12699,N_12518);
nand U14387 (N_14387,N_13180,N_13127);
or U14388 (N_14388,N_12732,N_12722);
or U14389 (N_14389,N_12287,N_13218);
and U14390 (N_14390,N_12681,N_12103);
or U14391 (N_14391,N_13147,N_12358);
xnor U14392 (N_14392,N_12254,N_13452);
and U14393 (N_14393,N_13261,N_12024);
nand U14394 (N_14394,N_12824,N_12397);
and U14395 (N_14395,N_12329,N_13109);
xor U14396 (N_14396,N_13413,N_12567);
and U14397 (N_14397,N_13035,N_13475);
or U14398 (N_14398,N_12205,N_12309);
or U14399 (N_14399,N_12871,N_12638);
nor U14400 (N_14400,N_13331,N_13053);
xnor U14401 (N_14401,N_12920,N_13313);
xor U14402 (N_14402,N_13119,N_12426);
nand U14403 (N_14403,N_12662,N_12628);
or U14404 (N_14404,N_12017,N_12057);
nor U14405 (N_14405,N_12929,N_13445);
or U14406 (N_14406,N_12502,N_12699);
nor U14407 (N_14407,N_13028,N_12614);
nor U14408 (N_14408,N_13327,N_13122);
nand U14409 (N_14409,N_12933,N_13363);
xor U14410 (N_14410,N_12512,N_12822);
nor U14411 (N_14411,N_12445,N_12278);
nand U14412 (N_14412,N_12963,N_12187);
and U14413 (N_14413,N_12719,N_12839);
and U14414 (N_14414,N_13373,N_12053);
nand U14415 (N_14415,N_13108,N_13402);
and U14416 (N_14416,N_12814,N_13144);
xnor U14417 (N_14417,N_12905,N_12260);
or U14418 (N_14418,N_12663,N_12666);
nand U14419 (N_14419,N_12431,N_12065);
and U14420 (N_14420,N_12551,N_12525);
xnor U14421 (N_14421,N_12034,N_12928);
nor U14422 (N_14422,N_13105,N_12932);
nor U14423 (N_14423,N_13244,N_12049);
or U14424 (N_14424,N_12151,N_12072);
nor U14425 (N_14425,N_12566,N_13007);
or U14426 (N_14426,N_12075,N_12146);
xnor U14427 (N_14427,N_12916,N_12269);
xor U14428 (N_14428,N_12197,N_12691);
nor U14429 (N_14429,N_13250,N_13084);
xor U14430 (N_14430,N_13166,N_12038);
nand U14431 (N_14431,N_12669,N_12292);
nand U14432 (N_14432,N_13371,N_12579);
or U14433 (N_14433,N_12483,N_13071);
nand U14434 (N_14434,N_12682,N_12772);
xnor U14435 (N_14435,N_12078,N_13452);
or U14436 (N_14436,N_12588,N_12954);
or U14437 (N_14437,N_12175,N_12928);
nor U14438 (N_14438,N_12585,N_12506);
or U14439 (N_14439,N_12707,N_12756);
xnor U14440 (N_14440,N_13291,N_12940);
nor U14441 (N_14441,N_12965,N_13408);
or U14442 (N_14442,N_12116,N_12566);
nor U14443 (N_14443,N_13429,N_12411);
nor U14444 (N_14444,N_12405,N_12440);
nand U14445 (N_14445,N_12586,N_12345);
or U14446 (N_14446,N_12213,N_13288);
and U14447 (N_14447,N_12019,N_12318);
xnor U14448 (N_14448,N_12791,N_12215);
and U14449 (N_14449,N_12349,N_12820);
nor U14450 (N_14450,N_12580,N_12648);
nand U14451 (N_14451,N_12786,N_12225);
nand U14452 (N_14452,N_13015,N_13399);
nand U14453 (N_14453,N_13491,N_12838);
nor U14454 (N_14454,N_13469,N_12961);
or U14455 (N_14455,N_13499,N_12840);
xnor U14456 (N_14456,N_12861,N_12296);
nor U14457 (N_14457,N_12487,N_13033);
or U14458 (N_14458,N_13483,N_12988);
nor U14459 (N_14459,N_12574,N_12592);
and U14460 (N_14460,N_13022,N_13229);
xnor U14461 (N_14461,N_12283,N_12132);
nor U14462 (N_14462,N_13481,N_13144);
and U14463 (N_14463,N_12225,N_12667);
and U14464 (N_14464,N_13108,N_12120);
or U14465 (N_14465,N_12309,N_13116);
or U14466 (N_14466,N_13372,N_12472);
and U14467 (N_14467,N_12461,N_12990);
nor U14468 (N_14468,N_12690,N_12508);
nand U14469 (N_14469,N_12931,N_12279);
nor U14470 (N_14470,N_12229,N_12039);
xnor U14471 (N_14471,N_13228,N_12832);
or U14472 (N_14472,N_12982,N_13436);
or U14473 (N_14473,N_13071,N_13360);
nor U14474 (N_14474,N_13481,N_12713);
nand U14475 (N_14475,N_12121,N_12063);
or U14476 (N_14476,N_12949,N_12201);
and U14477 (N_14477,N_13221,N_12585);
or U14478 (N_14478,N_12222,N_13235);
nor U14479 (N_14479,N_12985,N_12833);
or U14480 (N_14480,N_13176,N_12773);
and U14481 (N_14481,N_13168,N_12296);
and U14482 (N_14482,N_13309,N_12470);
xnor U14483 (N_14483,N_12703,N_12803);
nor U14484 (N_14484,N_12026,N_13363);
and U14485 (N_14485,N_12667,N_12205);
nand U14486 (N_14486,N_12506,N_13045);
nand U14487 (N_14487,N_12862,N_12508);
nor U14488 (N_14488,N_12071,N_12474);
nor U14489 (N_14489,N_13405,N_13440);
or U14490 (N_14490,N_13341,N_13326);
and U14491 (N_14491,N_12649,N_12234);
or U14492 (N_14492,N_13284,N_12230);
nand U14493 (N_14493,N_12104,N_12874);
nor U14494 (N_14494,N_12748,N_12346);
or U14495 (N_14495,N_13046,N_13021);
xnor U14496 (N_14496,N_13032,N_12081);
or U14497 (N_14497,N_13011,N_13048);
nor U14498 (N_14498,N_12438,N_12982);
and U14499 (N_14499,N_13158,N_13073);
nor U14500 (N_14500,N_12433,N_12993);
and U14501 (N_14501,N_12709,N_12704);
nand U14502 (N_14502,N_13338,N_12901);
nor U14503 (N_14503,N_12679,N_12693);
nand U14504 (N_14504,N_12398,N_12732);
or U14505 (N_14505,N_12039,N_12526);
or U14506 (N_14506,N_12384,N_12870);
and U14507 (N_14507,N_13483,N_12648);
xor U14508 (N_14508,N_12003,N_13340);
nor U14509 (N_14509,N_12154,N_12164);
xor U14510 (N_14510,N_13216,N_13466);
xnor U14511 (N_14511,N_12872,N_12637);
nand U14512 (N_14512,N_12971,N_12815);
and U14513 (N_14513,N_12306,N_13122);
nor U14514 (N_14514,N_12972,N_12724);
and U14515 (N_14515,N_13134,N_12562);
nor U14516 (N_14516,N_13181,N_12049);
nor U14517 (N_14517,N_12503,N_12779);
and U14518 (N_14518,N_12977,N_13138);
or U14519 (N_14519,N_13164,N_12618);
or U14520 (N_14520,N_12204,N_13136);
nand U14521 (N_14521,N_13270,N_13334);
xnor U14522 (N_14522,N_12773,N_12251);
xor U14523 (N_14523,N_12622,N_12100);
or U14524 (N_14524,N_12733,N_12872);
nor U14525 (N_14525,N_13466,N_12857);
and U14526 (N_14526,N_13172,N_12506);
xor U14527 (N_14527,N_12853,N_12196);
and U14528 (N_14528,N_12787,N_13287);
or U14529 (N_14529,N_12322,N_12162);
or U14530 (N_14530,N_13270,N_12934);
or U14531 (N_14531,N_12984,N_12803);
and U14532 (N_14532,N_12700,N_13035);
xnor U14533 (N_14533,N_12876,N_12996);
nor U14534 (N_14534,N_12889,N_12150);
nor U14535 (N_14535,N_13433,N_12016);
nor U14536 (N_14536,N_13134,N_13370);
nand U14537 (N_14537,N_12935,N_12757);
or U14538 (N_14538,N_13189,N_13299);
or U14539 (N_14539,N_12116,N_12775);
or U14540 (N_14540,N_12521,N_12246);
nand U14541 (N_14541,N_12234,N_12162);
or U14542 (N_14542,N_13263,N_13459);
or U14543 (N_14543,N_13383,N_13094);
and U14544 (N_14544,N_12484,N_12940);
nand U14545 (N_14545,N_12515,N_13227);
nor U14546 (N_14546,N_12037,N_13313);
or U14547 (N_14547,N_12835,N_13090);
nand U14548 (N_14548,N_12292,N_12590);
or U14549 (N_14549,N_12555,N_12983);
xor U14550 (N_14550,N_12796,N_12015);
or U14551 (N_14551,N_13076,N_12490);
nand U14552 (N_14552,N_13244,N_13257);
or U14553 (N_14553,N_13292,N_12428);
xnor U14554 (N_14554,N_13187,N_12603);
nand U14555 (N_14555,N_12207,N_13320);
xor U14556 (N_14556,N_13478,N_13389);
nor U14557 (N_14557,N_12327,N_13115);
nor U14558 (N_14558,N_12487,N_12719);
nor U14559 (N_14559,N_12140,N_12297);
nor U14560 (N_14560,N_12885,N_13352);
nor U14561 (N_14561,N_13380,N_13137);
nor U14562 (N_14562,N_12043,N_12717);
nor U14563 (N_14563,N_13096,N_12465);
nor U14564 (N_14564,N_12980,N_12565);
nand U14565 (N_14565,N_12732,N_12841);
and U14566 (N_14566,N_12830,N_12744);
nor U14567 (N_14567,N_13277,N_13107);
or U14568 (N_14568,N_13074,N_12118);
nand U14569 (N_14569,N_12062,N_12899);
xor U14570 (N_14570,N_13287,N_13041);
or U14571 (N_14571,N_12775,N_12742);
or U14572 (N_14572,N_12378,N_12135);
nor U14573 (N_14573,N_13117,N_12385);
and U14574 (N_14574,N_12410,N_13419);
or U14575 (N_14575,N_12839,N_12577);
nand U14576 (N_14576,N_13479,N_13354);
or U14577 (N_14577,N_12704,N_13315);
or U14578 (N_14578,N_13126,N_12552);
and U14579 (N_14579,N_12132,N_12431);
or U14580 (N_14580,N_12218,N_12031);
or U14581 (N_14581,N_12607,N_12862);
or U14582 (N_14582,N_12716,N_13485);
nor U14583 (N_14583,N_12581,N_12916);
nand U14584 (N_14584,N_12134,N_12198);
and U14585 (N_14585,N_12834,N_13268);
xor U14586 (N_14586,N_12828,N_12592);
xor U14587 (N_14587,N_13353,N_13343);
nor U14588 (N_14588,N_13318,N_12791);
and U14589 (N_14589,N_12691,N_12162);
xnor U14590 (N_14590,N_12807,N_13378);
nor U14591 (N_14591,N_12719,N_12580);
and U14592 (N_14592,N_13120,N_13119);
xor U14593 (N_14593,N_12487,N_12634);
nor U14594 (N_14594,N_12021,N_12346);
nand U14595 (N_14595,N_12878,N_12090);
nor U14596 (N_14596,N_12814,N_13062);
or U14597 (N_14597,N_13394,N_13186);
and U14598 (N_14598,N_12762,N_12446);
xnor U14599 (N_14599,N_12074,N_12851);
or U14600 (N_14600,N_12373,N_12601);
or U14601 (N_14601,N_12166,N_12960);
xor U14602 (N_14602,N_12615,N_12091);
xnor U14603 (N_14603,N_12260,N_12421);
and U14604 (N_14604,N_13063,N_13461);
or U14605 (N_14605,N_13459,N_13017);
and U14606 (N_14606,N_12256,N_13005);
nand U14607 (N_14607,N_13275,N_13063);
nand U14608 (N_14608,N_12705,N_13180);
or U14609 (N_14609,N_12419,N_13183);
or U14610 (N_14610,N_12226,N_12275);
xor U14611 (N_14611,N_12934,N_13011);
and U14612 (N_14612,N_13273,N_12307);
xor U14613 (N_14613,N_13164,N_12716);
nand U14614 (N_14614,N_12112,N_12943);
nor U14615 (N_14615,N_12635,N_12996);
nand U14616 (N_14616,N_12421,N_12766);
nand U14617 (N_14617,N_13300,N_12564);
nor U14618 (N_14618,N_12073,N_12785);
or U14619 (N_14619,N_13173,N_12985);
or U14620 (N_14620,N_12732,N_12813);
or U14621 (N_14621,N_12147,N_13071);
and U14622 (N_14622,N_12761,N_12637);
and U14623 (N_14623,N_12538,N_12412);
or U14624 (N_14624,N_13098,N_12990);
xnor U14625 (N_14625,N_13270,N_12173);
and U14626 (N_14626,N_12404,N_12688);
and U14627 (N_14627,N_12261,N_12981);
xor U14628 (N_14628,N_12102,N_12745);
nand U14629 (N_14629,N_13006,N_12711);
and U14630 (N_14630,N_12325,N_12674);
nand U14631 (N_14631,N_12944,N_13442);
or U14632 (N_14632,N_12546,N_12302);
or U14633 (N_14633,N_12949,N_13216);
nor U14634 (N_14634,N_13475,N_12722);
xnor U14635 (N_14635,N_12622,N_12849);
and U14636 (N_14636,N_12070,N_13097);
nand U14637 (N_14637,N_12799,N_12978);
xor U14638 (N_14638,N_13370,N_12327);
nor U14639 (N_14639,N_13338,N_12808);
nand U14640 (N_14640,N_12274,N_12879);
nor U14641 (N_14641,N_13465,N_13069);
nor U14642 (N_14642,N_13302,N_13136);
nor U14643 (N_14643,N_13073,N_12234);
or U14644 (N_14644,N_12697,N_12286);
nand U14645 (N_14645,N_12879,N_12044);
nand U14646 (N_14646,N_13270,N_12511);
xor U14647 (N_14647,N_12745,N_12049);
nand U14648 (N_14648,N_13011,N_12864);
nor U14649 (N_14649,N_13408,N_13390);
or U14650 (N_14650,N_13342,N_12183);
nand U14651 (N_14651,N_13226,N_12198);
xnor U14652 (N_14652,N_12195,N_13016);
nand U14653 (N_14653,N_12189,N_12432);
xor U14654 (N_14654,N_12991,N_13485);
nand U14655 (N_14655,N_12984,N_12417);
nor U14656 (N_14656,N_13381,N_13109);
and U14657 (N_14657,N_13340,N_12473);
xnor U14658 (N_14658,N_12585,N_12787);
and U14659 (N_14659,N_12415,N_12700);
and U14660 (N_14660,N_12985,N_12288);
nand U14661 (N_14661,N_13233,N_12336);
nand U14662 (N_14662,N_12920,N_13094);
or U14663 (N_14663,N_12424,N_12909);
nor U14664 (N_14664,N_13243,N_12150);
xor U14665 (N_14665,N_12299,N_12198);
nand U14666 (N_14666,N_12875,N_12058);
nand U14667 (N_14667,N_12858,N_13169);
xor U14668 (N_14668,N_13098,N_13296);
nand U14669 (N_14669,N_13082,N_13259);
nor U14670 (N_14670,N_13459,N_12806);
and U14671 (N_14671,N_12832,N_12181);
nand U14672 (N_14672,N_12097,N_13042);
or U14673 (N_14673,N_12282,N_12183);
nor U14674 (N_14674,N_12078,N_13447);
nor U14675 (N_14675,N_12167,N_12841);
xor U14676 (N_14676,N_13034,N_12827);
nor U14677 (N_14677,N_13094,N_12403);
nor U14678 (N_14678,N_13332,N_12342);
nor U14679 (N_14679,N_13497,N_13364);
xnor U14680 (N_14680,N_13413,N_13373);
nand U14681 (N_14681,N_12640,N_12783);
nor U14682 (N_14682,N_13095,N_12803);
nor U14683 (N_14683,N_13182,N_13160);
or U14684 (N_14684,N_12808,N_12297);
and U14685 (N_14685,N_13476,N_12776);
and U14686 (N_14686,N_12113,N_12743);
and U14687 (N_14687,N_12412,N_13294);
xnor U14688 (N_14688,N_12952,N_13185);
nand U14689 (N_14689,N_12677,N_12313);
nand U14690 (N_14690,N_12128,N_13092);
or U14691 (N_14691,N_12092,N_12208);
nor U14692 (N_14692,N_13116,N_12635);
and U14693 (N_14693,N_13061,N_12262);
and U14694 (N_14694,N_12902,N_12285);
nor U14695 (N_14695,N_13417,N_12623);
nor U14696 (N_14696,N_12564,N_13202);
and U14697 (N_14697,N_12341,N_12206);
nand U14698 (N_14698,N_12073,N_12880);
nand U14699 (N_14699,N_13439,N_13385);
nor U14700 (N_14700,N_12406,N_13497);
nand U14701 (N_14701,N_13019,N_12267);
nand U14702 (N_14702,N_12685,N_12170);
nor U14703 (N_14703,N_12749,N_12800);
and U14704 (N_14704,N_13459,N_12783);
or U14705 (N_14705,N_12509,N_12387);
or U14706 (N_14706,N_12742,N_12113);
or U14707 (N_14707,N_12028,N_12734);
xor U14708 (N_14708,N_12665,N_13188);
and U14709 (N_14709,N_13179,N_12857);
nor U14710 (N_14710,N_12156,N_13348);
or U14711 (N_14711,N_12195,N_13102);
or U14712 (N_14712,N_12354,N_12446);
nand U14713 (N_14713,N_12289,N_12110);
or U14714 (N_14714,N_12811,N_12966);
nand U14715 (N_14715,N_12529,N_12025);
nand U14716 (N_14716,N_12811,N_12027);
or U14717 (N_14717,N_13416,N_13316);
nor U14718 (N_14718,N_13189,N_12293);
nand U14719 (N_14719,N_12691,N_12279);
nor U14720 (N_14720,N_12829,N_12399);
or U14721 (N_14721,N_13104,N_12374);
nor U14722 (N_14722,N_12617,N_12032);
and U14723 (N_14723,N_13361,N_13333);
or U14724 (N_14724,N_13151,N_12275);
xor U14725 (N_14725,N_12629,N_12126);
and U14726 (N_14726,N_12967,N_12263);
and U14727 (N_14727,N_12477,N_12441);
nand U14728 (N_14728,N_13122,N_13439);
nand U14729 (N_14729,N_12440,N_12433);
and U14730 (N_14730,N_12331,N_12736);
nand U14731 (N_14731,N_12129,N_13217);
nand U14732 (N_14732,N_12286,N_12501);
nand U14733 (N_14733,N_13019,N_13066);
or U14734 (N_14734,N_12734,N_12962);
nor U14735 (N_14735,N_12526,N_12227);
xnor U14736 (N_14736,N_13192,N_12223);
xor U14737 (N_14737,N_12489,N_13447);
nor U14738 (N_14738,N_12049,N_12286);
nor U14739 (N_14739,N_13199,N_12628);
or U14740 (N_14740,N_13383,N_13060);
nor U14741 (N_14741,N_12803,N_12439);
and U14742 (N_14742,N_12338,N_12656);
or U14743 (N_14743,N_12944,N_12662);
nand U14744 (N_14744,N_12391,N_12839);
nor U14745 (N_14745,N_13435,N_12348);
and U14746 (N_14746,N_13026,N_12284);
and U14747 (N_14747,N_13407,N_12937);
xnor U14748 (N_14748,N_12782,N_12800);
nor U14749 (N_14749,N_13018,N_13226);
nand U14750 (N_14750,N_13129,N_13030);
or U14751 (N_14751,N_13048,N_12777);
nor U14752 (N_14752,N_13487,N_12367);
and U14753 (N_14753,N_13451,N_12075);
nor U14754 (N_14754,N_12416,N_13158);
nor U14755 (N_14755,N_12221,N_12428);
or U14756 (N_14756,N_12480,N_13212);
or U14757 (N_14757,N_12953,N_13099);
or U14758 (N_14758,N_12533,N_12339);
nand U14759 (N_14759,N_12396,N_12180);
and U14760 (N_14760,N_13108,N_12465);
nor U14761 (N_14761,N_12042,N_12073);
and U14762 (N_14762,N_12079,N_13105);
nand U14763 (N_14763,N_12796,N_12266);
nand U14764 (N_14764,N_12142,N_12408);
and U14765 (N_14765,N_13161,N_12235);
or U14766 (N_14766,N_12707,N_12751);
nor U14767 (N_14767,N_12452,N_12590);
nand U14768 (N_14768,N_13112,N_12947);
nor U14769 (N_14769,N_13212,N_12616);
nor U14770 (N_14770,N_13116,N_12408);
and U14771 (N_14771,N_12879,N_12510);
or U14772 (N_14772,N_12476,N_12553);
xor U14773 (N_14773,N_12280,N_12487);
or U14774 (N_14774,N_12823,N_12656);
or U14775 (N_14775,N_13135,N_12408);
and U14776 (N_14776,N_12683,N_12772);
nand U14777 (N_14777,N_13373,N_12378);
nor U14778 (N_14778,N_12951,N_12006);
or U14779 (N_14779,N_12488,N_13420);
xnor U14780 (N_14780,N_12169,N_12642);
xnor U14781 (N_14781,N_12974,N_13498);
and U14782 (N_14782,N_13142,N_12405);
nand U14783 (N_14783,N_12146,N_13132);
nor U14784 (N_14784,N_13042,N_12246);
xnor U14785 (N_14785,N_12008,N_12575);
nor U14786 (N_14786,N_12736,N_12499);
and U14787 (N_14787,N_12784,N_12092);
and U14788 (N_14788,N_12910,N_12740);
or U14789 (N_14789,N_12026,N_12321);
or U14790 (N_14790,N_12980,N_13102);
or U14791 (N_14791,N_12127,N_13076);
xor U14792 (N_14792,N_12648,N_12941);
or U14793 (N_14793,N_12166,N_12959);
nor U14794 (N_14794,N_12788,N_13401);
nor U14795 (N_14795,N_13352,N_13190);
nand U14796 (N_14796,N_12779,N_12684);
and U14797 (N_14797,N_12152,N_13121);
nor U14798 (N_14798,N_12386,N_13118);
xor U14799 (N_14799,N_12053,N_12174);
nand U14800 (N_14800,N_12823,N_12706);
xor U14801 (N_14801,N_13032,N_12344);
nor U14802 (N_14802,N_12254,N_12122);
nand U14803 (N_14803,N_12658,N_12078);
and U14804 (N_14804,N_13091,N_12515);
nand U14805 (N_14805,N_13003,N_12778);
nand U14806 (N_14806,N_12160,N_13141);
and U14807 (N_14807,N_12993,N_13027);
and U14808 (N_14808,N_12305,N_12817);
or U14809 (N_14809,N_12096,N_13303);
and U14810 (N_14810,N_12749,N_13127);
nand U14811 (N_14811,N_12928,N_12515);
nor U14812 (N_14812,N_12506,N_12775);
nor U14813 (N_14813,N_13471,N_13421);
nand U14814 (N_14814,N_12813,N_12310);
and U14815 (N_14815,N_12110,N_13301);
or U14816 (N_14816,N_13472,N_12305);
xnor U14817 (N_14817,N_12635,N_13387);
nor U14818 (N_14818,N_12141,N_12706);
and U14819 (N_14819,N_13130,N_13276);
nand U14820 (N_14820,N_12650,N_12993);
xor U14821 (N_14821,N_13475,N_12744);
nor U14822 (N_14822,N_12961,N_12599);
or U14823 (N_14823,N_12062,N_12289);
nand U14824 (N_14824,N_12306,N_12116);
xor U14825 (N_14825,N_12261,N_12091);
nand U14826 (N_14826,N_12839,N_13096);
nand U14827 (N_14827,N_13484,N_12461);
or U14828 (N_14828,N_13273,N_12744);
nor U14829 (N_14829,N_12658,N_13467);
and U14830 (N_14830,N_13257,N_12752);
xnor U14831 (N_14831,N_13307,N_12496);
and U14832 (N_14832,N_13374,N_12065);
nand U14833 (N_14833,N_13481,N_12220);
nor U14834 (N_14834,N_12190,N_13210);
and U14835 (N_14835,N_12456,N_13369);
nor U14836 (N_14836,N_12727,N_13282);
and U14837 (N_14837,N_13160,N_12706);
nor U14838 (N_14838,N_13460,N_13325);
or U14839 (N_14839,N_13476,N_12445);
or U14840 (N_14840,N_12739,N_12684);
and U14841 (N_14841,N_12818,N_13038);
or U14842 (N_14842,N_12984,N_13054);
nor U14843 (N_14843,N_12887,N_12827);
nand U14844 (N_14844,N_12418,N_12245);
xor U14845 (N_14845,N_12274,N_12887);
and U14846 (N_14846,N_13231,N_13023);
nor U14847 (N_14847,N_12725,N_13138);
nor U14848 (N_14848,N_12604,N_12037);
nand U14849 (N_14849,N_13437,N_13077);
nor U14850 (N_14850,N_12398,N_12126);
and U14851 (N_14851,N_13054,N_12864);
or U14852 (N_14852,N_12623,N_12437);
nand U14853 (N_14853,N_13426,N_12692);
and U14854 (N_14854,N_12633,N_12090);
and U14855 (N_14855,N_12700,N_12708);
nor U14856 (N_14856,N_12826,N_13449);
nor U14857 (N_14857,N_12011,N_13382);
or U14858 (N_14858,N_12980,N_12015);
and U14859 (N_14859,N_12387,N_12237);
nor U14860 (N_14860,N_13106,N_12869);
xnor U14861 (N_14861,N_12838,N_13330);
nor U14862 (N_14862,N_12174,N_13371);
xnor U14863 (N_14863,N_13091,N_12987);
nor U14864 (N_14864,N_12123,N_13425);
and U14865 (N_14865,N_13387,N_12111);
nand U14866 (N_14866,N_13207,N_13401);
nand U14867 (N_14867,N_13163,N_12289);
nand U14868 (N_14868,N_12020,N_12429);
and U14869 (N_14869,N_12473,N_13278);
nor U14870 (N_14870,N_12055,N_12429);
nand U14871 (N_14871,N_12130,N_12954);
or U14872 (N_14872,N_12115,N_13317);
nor U14873 (N_14873,N_12013,N_12755);
xnor U14874 (N_14874,N_13419,N_12162);
or U14875 (N_14875,N_12342,N_13107);
or U14876 (N_14876,N_12489,N_12166);
nand U14877 (N_14877,N_13342,N_12427);
and U14878 (N_14878,N_13264,N_13370);
or U14879 (N_14879,N_12934,N_12643);
and U14880 (N_14880,N_13186,N_13137);
nand U14881 (N_14881,N_12015,N_13161);
and U14882 (N_14882,N_12830,N_12403);
or U14883 (N_14883,N_13248,N_12304);
and U14884 (N_14884,N_13261,N_12156);
and U14885 (N_14885,N_12758,N_12078);
nand U14886 (N_14886,N_12033,N_13083);
nor U14887 (N_14887,N_12724,N_12948);
nor U14888 (N_14888,N_12976,N_13063);
nand U14889 (N_14889,N_12522,N_12541);
nor U14890 (N_14890,N_12109,N_12718);
nor U14891 (N_14891,N_13125,N_12668);
nor U14892 (N_14892,N_12004,N_13439);
xnor U14893 (N_14893,N_12966,N_12856);
xor U14894 (N_14894,N_13420,N_13110);
nand U14895 (N_14895,N_12827,N_13023);
xor U14896 (N_14896,N_13236,N_12703);
nor U14897 (N_14897,N_12548,N_12720);
nand U14898 (N_14898,N_12692,N_12767);
nand U14899 (N_14899,N_12214,N_12601);
or U14900 (N_14900,N_12977,N_12112);
nand U14901 (N_14901,N_12561,N_12246);
nand U14902 (N_14902,N_13492,N_12113);
nand U14903 (N_14903,N_12913,N_12430);
and U14904 (N_14904,N_13147,N_12417);
and U14905 (N_14905,N_12508,N_12719);
nor U14906 (N_14906,N_13457,N_13313);
and U14907 (N_14907,N_12837,N_12264);
and U14908 (N_14908,N_12675,N_12022);
nand U14909 (N_14909,N_12664,N_12584);
nor U14910 (N_14910,N_12229,N_12253);
nor U14911 (N_14911,N_12842,N_12009);
and U14912 (N_14912,N_12924,N_12559);
and U14913 (N_14913,N_13456,N_13123);
nand U14914 (N_14914,N_12847,N_12232);
and U14915 (N_14915,N_12573,N_13327);
and U14916 (N_14916,N_13123,N_12390);
nand U14917 (N_14917,N_12233,N_13480);
nand U14918 (N_14918,N_13349,N_13436);
nor U14919 (N_14919,N_12142,N_13110);
nand U14920 (N_14920,N_12919,N_13471);
or U14921 (N_14921,N_12301,N_12977);
nor U14922 (N_14922,N_13476,N_13242);
and U14923 (N_14923,N_13306,N_12118);
xor U14924 (N_14924,N_12612,N_13326);
nand U14925 (N_14925,N_12744,N_13361);
and U14926 (N_14926,N_13402,N_12627);
nor U14927 (N_14927,N_12928,N_13041);
and U14928 (N_14928,N_12530,N_12711);
xnor U14929 (N_14929,N_13240,N_12352);
or U14930 (N_14930,N_12539,N_12096);
and U14931 (N_14931,N_12181,N_12908);
and U14932 (N_14932,N_12322,N_12895);
and U14933 (N_14933,N_12576,N_12440);
nand U14934 (N_14934,N_13434,N_13275);
nor U14935 (N_14935,N_12512,N_13066);
nand U14936 (N_14936,N_13279,N_12082);
nand U14937 (N_14937,N_12985,N_12170);
and U14938 (N_14938,N_12797,N_12235);
nor U14939 (N_14939,N_12056,N_12985);
or U14940 (N_14940,N_12842,N_12830);
nand U14941 (N_14941,N_12157,N_12877);
xnor U14942 (N_14942,N_12332,N_12452);
or U14943 (N_14943,N_12419,N_12758);
nand U14944 (N_14944,N_13110,N_13003);
nand U14945 (N_14945,N_13207,N_12361);
nor U14946 (N_14946,N_12176,N_12452);
nor U14947 (N_14947,N_13138,N_13467);
and U14948 (N_14948,N_13480,N_13151);
and U14949 (N_14949,N_12452,N_12955);
and U14950 (N_14950,N_13305,N_12610);
nor U14951 (N_14951,N_12393,N_12751);
or U14952 (N_14952,N_13197,N_13336);
nand U14953 (N_14953,N_12382,N_12994);
or U14954 (N_14954,N_13308,N_12464);
nor U14955 (N_14955,N_12911,N_12864);
or U14956 (N_14956,N_12854,N_12719);
nand U14957 (N_14957,N_12697,N_12717);
nor U14958 (N_14958,N_13152,N_12155);
nor U14959 (N_14959,N_12838,N_13380);
or U14960 (N_14960,N_12817,N_13139);
or U14961 (N_14961,N_13027,N_12100);
or U14962 (N_14962,N_13183,N_12847);
xor U14963 (N_14963,N_13085,N_12892);
nand U14964 (N_14964,N_13371,N_13158);
and U14965 (N_14965,N_12598,N_12061);
and U14966 (N_14966,N_12412,N_12577);
nor U14967 (N_14967,N_13496,N_12164);
and U14968 (N_14968,N_12488,N_12540);
or U14969 (N_14969,N_12842,N_12805);
xor U14970 (N_14970,N_12691,N_12001);
nand U14971 (N_14971,N_13195,N_12164);
nand U14972 (N_14972,N_12589,N_12457);
and U14973 (N_14973,N_12228,N_12983);
or U14974 (N_14974,N_12875,N_12606);
or U14975 (N_14975,N_13498,N_12317);
or U14976 (N_14976,N_12140,N_12021);
or U14977 (N_14977,N_12609,N_12727);
nand U14978 (N_14978,N_13072,N_12438);
nand U14979 (N_14979,N_12208,N_13433);
xnor U14980 (N_14980,N_12452,N_13483);
nand U14981 (N_14981,N_12229,N_12338);
and U14982 (N_14982,N_12387,N_12326);
or U14983 (N_14983,N_12179,N_12134);
nand U14984 (N_14984,N_12013,N_12112);
nor U14985 (N_14985,N_12795,N_12376);
xor U14986 (N_14986,N_12787,N_13293);
or U14987 (N_14987,N_13049,N_13005);
nor U14988 (N_14988,N_12351,N_13147);
and U14989 (N_14989,N_13304,N_12937);
or U14990 (N_14990,N_12698,N_12580);
nand U14991 (N_14991,N_12184,N_12489);
and U14992 (N_14992,N_12691,N_12844);
and U14993 (N_14993,N_12223,N_13496);
nor U14994 (N_14994,N_12116,N_12524);
nand U14995 (N_14995,N_12151,N_12481);
nand U14996 (N_14996,N_12268,N_12231);
or U14997 (N_14997,N_13379,N_12957);
nor U14998 (N_14998,N_12171,N_13317);
nor U14999 (N_14999,N_12360,N_12940);
or UO_0 (O_0,N_14743,N_14253);
or UO_1 (O_1,N_14319,N_14492);
and UO_2 (O_2,N_14036,N_13841);
nand UO_3 (O_3,N_13737,N_14884);
or UO_4 (O_4,N_14927,N_14370);
nor UO_5 (O_5,N_14602,N_13630);
or UO_6 (O_6,N_14216,N_13536);
nor UO_7 (O_7,N_14828,N_14397);
and UO_8 (O_8,N_14413,N_13704);
nand UO_9 (O_9,N_14192,N_14145);
nor UO_10 (O_10,N_14543,N_14475);
and UO_11 (O_11,N_14798,N_14570);
nor UO_12 (O_12,N_14060,N_14598);
nor UO_13 (O_13,N_14968,N_13669);
nor UO_14 (O_14,N_14883,N_13905);
nand UO_15 (O_15,N_14215,N_13789);
nand UO_16 (O_16,N_14423,N_14173);
nor UO_17 (O_17,N_14635,N_13592);
xnor UO_18 (O_18,N_14749,N_13582);
or UO_19 (O_19,N_13634,N_14843);
xor UO_20 (O_20,N_14810,N_14086);
nor UO_21 (O_21,N_14594,N_14252);
nor UO_22 (O_22,N_14693,N_13939);
nand UO_23 (O_23,N_14524,N_14110);
xor UO_24 (O_24,N_14988,N_13940);
or UO_25 (O_25,N_14646,N_14129);
nand UO_26 (O_26,N_14160,N_13728);
and UO_27 (O_27,N_14963,N_14276);
and UO_28 (O_28,N_13963,N_14074);
nor UO_29 (O_29,N_14244,N_14981);
nor UO_30 (O_30,N_14915,N_14035);
or UO_31 (O_31,N_14738,N_14403);
nand UO_32 (O_32,N_14499,N_14596);
nand UO_33 (O_33,N_13810,N_13616);
nor UO_34 (O_34,N_13894,N_13666);
and UO_35 (O_35,N_14661,N_13547);
nand UO_36 (O_36,N_13542,N_14518);
nor UO_37 (O_37,N_14766,N_14158);
nor UO_38 (O_38,N_13613,N_14357);
nor UO_39 (O_39,N_14925,N_14010);
nor UO_40 (O_40,N_14666,N_14529);
nand UO_41 (O_41,N_14474,N_14973);
nand UO_42 (O_42,N_14838,N_13842);
nor UO_43 (O_43,N_14502,N_13752);
nor UO_44 (O_44,N_14029,N_14681);
xnor UO_45 (O_45,N_14366,N_13720);
nand UO_46 (O_46,N_14942,N_14669);
or UO_47 (O_47,N_13927,N_13748);
xor UO_48 (O_48,N_13667,N_14262);
nor UO_49 (O_49,N_14378,N_14909);
and UO_50 (O_50,N_13836,N_14923);
and UO_51 (O_51,N_14194,N_13987);
or UO_52 (O_52,N_13791,N_13936);
nand UO_53 (O_53,N_14470,N_14002);
and UO_54 (O_54,N_14339,N_14419);
and UO_55 (O_55,N_14450,N_14875);
or UO_56 (O_56,N_14852,N_14658);
and UO_57 (O_57,N_14612,N_14157);
and UO_58 (O_58,N_13850,N_14428);
nand UO_59 (O_59,N_14579,N_14146);
or UO_60 (O_60,N_14355,N_14633);
or UO_61 (O_61,N_14618,N_13769);
nor UO_62 (O_62,N_14053,N_14954);
and UO_63 (O_63,N_14928,N_14685);
xor UO_64 (O_64,N_14437,N_14171);
or UO_65 (O_65,N_13935,N_14608);
or UO_66 (O_66,N_13937,N_14085);
or UO_67 (O_67,N_13952,N_14358);
nand UO_68 (O_68,N_14407,N_14985);
nand UO_69 (O_69,N_14730,N_13636);
and UO_70 (O_70,N_14193,N_14603);
nor UO_71 (O_71,N_14087,N_14426);
or UO_72 (O_72,N_13717,N_14815);
and UO_73 (O_73,N_13610,N_14090);
nor UO_74 (O_74,N_14684,N_14716);
nor UO_75 (O_75,N_14264,N_14638);
and UO_76 (O_76,N_14991,N_14007);
xnor UO_77 (O_77,N_14369,N_14978);
nor UO_78 (O_78,N_13982,N_13639);
nor UO_79 (O_79,N_13568,N_14567);
or UO_80 (O_80,N_14694,N_13853);
nor UO_81 (O_81,N_14208,N_14333);
and UO_82 (O_82,N_14563,N_14170);
xnor UO_83 (O_83,N_13744,N_13594);
nand UO_84 (O_84,N_13687,N_14288);
nand UO_85 (O_85,N_13924,N_13825);
xnor UO_86 (O_86,N_14381,N_14095);
or UO_87 (O_87,N_13673,N_14780);
or UO_88 (O_88,N_14817,N_14962);
or UO_89 (O_89,N_13807,N_13620);
and UO_90 (O_90,N_14682,N_13545);
or UO_91 (O_91,N_14523,N_13538);
xor UO_92 (O_92,N_14575,N_13915);
nor UO_93 (O_93,N_13816,N_13938);
nand UO_94 (O_94,N_14398,N_14860);
nand UO_95 (O_95,N_14167,N_14237);
and UO_96 (O_96,N_14917,N_13897);
or UO_97 (O_97,N_14334,N_13797);
nand UO_98 (O_98,N_14561,N_14512);
or UO_99 (O_99,N_14178,N_14112);
nor UO_100 (O_100,N_13925,N_13901);
nand UO_101 (O_101,N_14105,N_13862);
nand UO_102 (O_102,N_13556,N_13962);
nor UO_103 (O_103,N_14533,N_14506);
nand UO_104 (O_104,N_13864,N_14177);
and UO_105 (O_105,N_14839,N_14517);
and UO_106 (O_106,N_14840,N_14154);
or UO_107 (O_107,N_13882,N_13688);
nor UO_108 (O_108,N_14924,N_14332);
nand UO_109 (O_109,N_14793,N_13680);
nor UO_110 (O_110,N_14020,N_14102);
or UO_111 (O_111,N_13674,N_14240);
nand UO_112 (O_112,N_14084,N_14256);
nand UO_113 (O_113,N_13731,N_14993);
and UO_114 (O_114,N_14510,N_13931);
nor UO_115 (O_115,N_13656,N_14511);
or UO_116 (O_116,N_13892,N_13786);
nand UO_117 (O_117,N_14757,N_13524);
xnor UO_118 (O_118,N_14695,N_14786);
or UO_119 (O_119,N_14905,N_14195);
nor UO_120 (O_120,N_14149,N_13900);
nand UO_121 (O_121,N_14094,N_14077);
or UO_122 (O_122,N_14486,N_14325);
and UO_123 (O_123,N_14034,N_14813);
or UO_124 (O_124,N_14373,N_14099);
nand UO_125 (O_125,N_14812,N_14785);
nand UO_126 (O_126,N_13829,N_13911);
or UO_127 (O_127,N_14179,N_14649);
nor UO_128 (O_128,N_14043,N_13887);
nor UO_129 (O_129,N_14477,N_14736);
or UO_130 (O_130,N_14420,N_14297);
or UO_131 (O_131,N_14372,N_14304);
nor UO_132 (O_132,N_14803,N_14476);
nor UO_133 (O_133,N_13819,N_13746);
xor UO_134 (O_134,N_14630,N_13934);
nor UO_135 (O_135,N_13511,N_14634);
or UO_136 (O_136,N_14345,N_14600);
nand UO_137 (O_137,N_14848,N_14075);
or UO_138 (O_138,N_13595,N_13893);
nand UO_139 (O_139,N_14854,N_14360);
or UO_140 (O_140,N_14070,N_14218);
nor UO_141 (O_141,N_14768,N_14837);
or UO_142 (O_142,N_13615,N_14834);
xnor UO_143 (O_143,N_14759,N_13770);
or UO_144 (O_144,N_14957,N_13824);
nor UO_145 (O_145,N_14702,N_14067);
nor UO_146 (O_146,N_13908,N_13540);
or UO_147 (O_147,N_14796,N_13500);
or UO_148 (O_148,N_14125,N_14583);
or UO_149 (O_149,N_13781,N_13798);
xnor UO_150 (O_150,N_13638,N_13677);
or UO_151 (O_151,N_14096,N_14558);
nor UO_152 (O_152,N_13655,N_14960);
nand UO_153 (O_153,N_14281,N_14341);
nand UO_154 (O_154,N_13648,N_14498);
and UO_155 (O_155,N_13566,N_14525);
and UO_156 (O_156,N_14604,N_14677);
or UO_157 (O_157,N_13771,N_14710);
or UO_158 (O_158,N_13516,N_13909);
or UO_159 (O_159,N_14151,N_14436);
or UO_160 (O_160,N_14201,N_14150);
or UO_161 (O_161,N_14374,N_13676);
nand UO_162 (O_162,N_13628,N_13999);
and UO_163 (O_163,N_14557,N_14967);
or UO_164 (O_164,N_14528,N_14180);
xnor UO_165 (O_165,N_14331,N_14664);
nor UO_166 (O_166,N_13986,N_14997);
nor UO_167 (O_167,N_14811,N_14037);
or UO_168 (O_168,N_14431,N_14920);
nor UO_169 (O_169,N_13572,N_14266);
nand UO_170 (O_170,N_13753,N_14877);
or UO_171 (O_171,N_13805,N_14592);
or UO_172 (O_172,N_14109,N_14422);
nor UO_173 (O_173,N_14033,N_14655);
nor UO_174 (O_174,N_14235,N_13766);
or UO_175 (O_175,N_14019,N_14560);
or UO_176 (O_176,N_13881,N_14122);
nand UO_177 (O_177,N_14337,N_14054);
xor UO_178 (O_178,N_14340,N_14490);
nor UO_179 (O_179,N_14894,N_14184);
nor UO_180 (O_180,N_14027,N_14701);
nand UO_181 (O_181,N_14064,N_14338);
nand UO_182 (O_182,N_13692,N_14041);
or UO_183 (O_183,N_14471,N_14031);
nor UO_184 (O_184,N_13736,N_13856);
nand UO_185 (O_185,N_14222,N_14039);
nand UO_186 (O_186,N_13652,N_14800);
and UO_187 (O_187,N_14169,N_13644);
nand UO_188 (O_188,N_13812,N_13741);
or UO_189 (O_189,N_13851,N_14462);
nand UO_190 (O_190,N_14527,N_14092);
and UO_191 (O_191,N_14126,N_13989);
xor UO_192 (O_192,N_14580,N_14389);
and UO_193 (O_193,N_14872,N_14765);
nand UO_194 (O_194,N_14497,N_14998);
nor UO_195 (O_195,N_13838,N_14469);
nor UO_196 (O_196,N_13848,N_14404);
or UO_197 (O_197,N_13942,N_14994);
nor UO_198 (O_198,N_13537,N_14636);
nor UO_199 (O_199,N_14190,N_14457);
and UO_200 (O_200,N_14779,N_14613);
xnor UO_201 (O_201,N_14881,N_14001);
xnor UO_202 (O_202,N_14822,N_13928);
nor UO_203 (O_203,N_14934,N_13521);
nand UO_204 (O_204,N_14657,N_13612);
or UO_205 (O_205,N_13947,N_13926);
or UO_206 (O_206,N_14624,N_14896);
and UO_207 (O_207,N_14255,N_14764);
nand UO_208 (O_208,N_13775,N_13581);
nand UO_209 (O_209,N_14484,N_14667);
nor UO_210 (O_210,N_14703,N_14069);
and UO_211 (O_211,N_14025,N_14520);
and UO_212 (O_212,N_14248,N_14162);
and UO_213 (O_213,N_14376,N_13782);
and UO_214 (O_214,N_14047,N_14893);
nand UO_215 (O_215,N_14732,N_13750);
nor UO_216 (O_216,N_14343,N_13519);
or UO_217 (O_217,N_14841,N_14865);
and UO_218 (O_218,N_13955,N_13632);
or UO_219 (O_219,N_14665,N_13994);
nor UO_220 (O_220,N_14752,N_14969);
nand UO_221 (O_221,N_13977,N_13877);
or UO_222 (O_222,N_13678,N_14734);
nor UO_223 (O_223,N_14936,N_14287);
nor UO_224 (O_224,N_14293,N_14754);
nand UO_225 (O_225,N_14607,N_14032);
nor UO_226 (O_226,N_14356,N_14818);
xor UO_227 (O_227,N_14017,N_14088);
or UO_228 (O_228,N_14731,N_14209);
nand UO_229 (O_229,N_14675,N_14229);
nor UO_230 (O_230,N_14117,N_13948);
nand UO_231 (O_231,N_13964,N_14294);
and UO_232 (O_232,N_14223,N_13988);
and UO_233 (O_233,N_14383,N_14737);
and UO_234 (O_234,N_14004,N_14713);
nor UO_235 (O_235,N_13954,N_14652);
xnor UO_236 (O_236,N_13563,N_13528);
nor UO_237 (O_237,N_13759,N_13831);
xnor UO_238 (O_238,N_13609,N_14559);
nand UO_239 (O_239,N_13861,N_14771);
nor UO_240 (O_240,N_14071,N_14846);
and UO_241 (O_241,N_14267,N_14683);
or UO_242 (O_242,N_14787,N_14776);
nor UO_243 (O_243,N_14619,N_14246);
and UO_244 (O_244,N_14116,N_14821);
and UO_245 (O_245,N_13596,N_14021);
nor UO_246 (O_246,N_13530,N_14965);
or UO_247 (O_247,N_14433,N_14516);
nor UO_248 (O_248,N_14553,N_14999);
nand UO_249 (O_249,N_14983,N_14313);
nand UO_250 (O_250,N_13505,N_14719);
and UO_251 (O_251,N_14265,N_14717);
and UO_252 (O_252,N_13689,N_13716);
or UO_253 (O_253,N_13967,N_14012);
and UO_254 (O_254,N_14705,N_14707);
and UO_255 (O_255,N_14590,N_14830);
and UO_256 (O_256,N_14274,N_14136);
nor UO_257 (O_257,N_14172,N_14671);
and UO_258 (O_258,N_14485,N_13837);
nand UO_259 (O_259,N_14254,N_13774);
and UO_260 (O_260,N_14862,N_14213);
and UO_261 (O_261,N_14142,N_13956);
nor UO_262 (O_262,N_14714,N_14748);
nand UO_263 (O_263,N_14003,N_14250);
and UO_264 (O_264,N_14692,N_13932);
or UO_265 (O_265,N_13907,N_13990);
nand UO_266 (O_266,N_14361,N_14300);
nand UO_267 (O_267,N_14836,N_14878);
nor UO_268 (O_268,N_14447,N_14522);
xor UO_269 (O_269,N_14891,N_14750);
nor UO_270 (O_270,N_14364,N_14014);
nor UO_271 (O_271,N_14678,N_14825);
nor UO_272 (O_272,N_14296,N_13790);
and UO_273 (O_273,N_14013,N_13873);
or UO_274 (O_274,N_14211,N_14940);
xor UO_275 (O_275,N_14260,N_13527);
or UO_276 (O_276,N_14066,N_13529);
or UO_277 (O_277,N_14165,N_14480);
nand UO_278 (O_278,N_13916,N_13830);
nor UO_279 (O_279,N_14611,N_13522);
and UO_280 (O_280,N_13557,N_14008);
xor UO_281 (O_281,N_14536,N_14442);
or UO_282 (O_282,N_14299,N_13501);
xor UO_283 (O_283,N_14586,N_13761);
xnor UO_284 (O_284,N_13583,N_14239);
or UO_285 (O_285,N_14249,N_14902);
nand UO_286 (O_286,N_14532,N_14055);
nor UO_287 (O_287,N_14483,N_14310);
and UO_288 (O_288,N_14697,N_13577);
nor UO_289 (O_289,N_14774,N_13625);
nand UO_290 (O_290,N_14496,N_14541);
nor UO_291 (O_291,N_14463,N_13561);
and UO_292 (O_292,N_14315,N_14143);
nor UO_293 (O_293,N_14482,N_14236);
xnor UO_294 (O_294,N_13679,N_13675);
xnor UO_295 (O_295,N_14911,N_14514);
nor UO_296 (O_296,N_13863,N_14704);
nand UO_297 (O_297,N_14460,N_13642);
nor UO_298 (O_298,N_14804,N_14508);
or UO_299 (O_299,N_13784,N_14856);
nor UO_300 (O_300,N_14577,N_14556);
or UO_301 (O_301,N_13534,N_13649);
and UO_302 (O_302,N_14879,N_13709);
or UO_303 (O_303,N_14913,N_14466);
or UO_304 (O_304,N_13629,N_14949);
nor UO_305 (O_305,N_13777,N_14279);
nand UO_306 (O_306,N_14809,N_14059);
or UO_307 (O_307,N_13957,N_14176);
nand UO_308 (O_308,N_13525,N_13698);
or UO_309 (O_309,N_14115,N_13661);
and UO_310 (O_310,N_14984,N_14912);
nand UO_311 (O_311,N_14467,N_13941);
nand UO_312 (O_312,N_13755,N_13682);
and UO_313 (O_313,N_14724,N_14353);
or UO_314 (O_314,N_14971,N_14790);
or UO_315 (O_315,N_14980,N_14270);
nor UO_316 (O_316,N_14904,N_13912);
or UO_317 (O_317,N_14329,N_14762);
nand UO_318 (O_318,N_13754,N_13772);
or UO_319 (O_319,N_14827,N_14342);
or UO_320 (O_320,N_13532,N_13898);
nor UO_321 (O_321,N_13619,N_14368);
or UO_322 (O_322,N_14302,N_14441);
and UO_323 (O_323,N_13855,N_13502);
or UO_324 (O_324,N_14111,N_13788);
or UO_325 (O_325,N_14844,N_13724);
nor UO_326 (O_326,N_14632,N_13890);
or UO_327 (O_327,N_14500,N_14011);
nand UO_328 (O_328,N_13965,N_14722);
nor UO_329 (O_329,N_13906,N_14349);
and UO_330 (O_330,N_14406,N_14974);
or UO_331 (O_331,N_14595,N_14947);
or UO_332 (O_332,N_13813,N_14674);
or UO_333 (O_333,N_13512,N_14727);
and UO_334 (O_334,N_14979,N_14439);
nor UO_335 (O_335,N_14599,N_14620);
nor UO_336 (O_336,N_14068,N_14400);
nand UO_337 (O_337,N_14409,N_13725);
or UO_338 (O_338,N_13827,N_14321);
xnor UO_339 (O_339,N_14849,N_14166);
nand UO_340 (O_340,N_14855,N_14182);
and UO_341 (O_341,N_14198,N_14335);
nor UO_342 (O_342,N_13579,N_13588);
or UO_343 (O_343,N_13562,N_14245);
or UO_344 (O_344,N_13718,N_14568);
and UO_345 (O_345,N_14910,N_13602);
nand UO_346 (O_346,N_13668,N_13576);
or UO_347 (O_347,N_13654,N_13598);
and UO_348 (O_348,N_14259,N_14197);
and UO_349 (O_349,N_14181,N_14725);
nor UO_350 (O_350,N_14408,N_14119);
or UO_351 (O_351,N_14455,N_14729);
nand UO_352 (O_352,N_14628,N_14783);
and UO_353 (O_353,N_14347,N_14900);
nor UO_354 (O_354,N_14972,N_14537);
and UO_355 (O_355,N_13622,N_13555);
nand UO_356 (O_356,N_13930,N_14895);
or UO_357 (O_357,N_14042,N_13840);
and UO_358 (O_358,N_14833,N_13803);
nand UO_359 (O_359,N_13995,N_14359);
and UO_360 (O_360,N_14481,N_14050);
nand UO_361 (O_361,N_14380,N_13876);
and UO_362 (O_362,N_14977,N_13705);
and UO_363 (O_363,N_14100,N_14513);
xnor UO_364 (O_364,N_14073,N_14943);
nor UO_365 (O_365,N_14344,N_13695);
nand UO_366 (O_366,N_13559,N_14091);
and UO_367 (O_367,N_14203,N_13880);
nand UO_368 (O_368,N_13657,N_14775);
and UO_369 (O_369,N_13822,N_13889);
and UO_370 (O_370,N_14187,N_14141);
xnor UO_371 (O_371,N_14614,N_14770);
and UO_372 (O_372,N_13708,N_13730);
nor UO_373 (O_373,N_14626,N_13870);
or UO_374 (O_374,N_14572,N_14515);
nor UO_375 (O_375,N_14371,N_13809);
and UO_376 (O_376,N_13697,N_14609);
or UO_377 (O_377,N_13618,N_13821);
nand UO_378 (O_378,N_14418,N_14653);
and UO_379 (O_379,N_14202,N_14610);
nand UO_380 (O_380,N_13608,N_14721);
and UO_381 (O_381,N_14384,N_14637);
nand UO_382 (O_382,N_14348,N_14217);
xnor UO_383 (O_383,N_14956,N_14044);
or UO_384 (O_384,N_13611,N_13681);
or UO_385 (O_385,N_14185,N_13972);
and UO_386 (O_386,N_13979,N_13518);
nand UO_387 (O_387,N_14625,N_14552);
and UO_388 (O_388,N_13763,N_14080);
nor UO_389 (O_389,N_13739,N_14221);
or UO_390 (O_390,N_14819,N_14323);
xor UO_391 (O_391,N_14672,N_13553);
nor UO_392 (O_392,N_13533,N_14670);
nor UO_393 (O_393,N_14935,N_14464);
xor UO_394 (O_394,N_14995,N_14200);
xor UO_395 (O_395,N_13891,N_14401);
or UO_396 (O_396,N_14107,N_14689);
nor UO_397 (O_397,N_13721,N_13921);
or UO_398 (O_398,N_14326,N_14565);
nand UO_399 (O_399,N_13552,N_13968);
nand UO_400 (O_400,N_13858,N_14842);
and UO_401 (O_401,N_13513,N_14263);
nor UO_402 (O_402,N_13883,N_13606);
nand UO_403 (O_403,N_14324,N_13817);
xnor UO_404 (O_404,N_14451,N_14573);
and UO_405 (O_405,N_13773,N_14745);
xnor UO_406 (O_406,N_14161,N_13814);
and UO_407 (O_407,N_13740,N_13765);
nand UO_408 (O_408,N_14715,N_14493);
nor UO_409 (O_409,N_14089,N_14679);
nor UO_410 (O_410,N_14542,N_13846);
or UO_411 (O_411,N_14708,N_14395);
or UO_412 (O_412,N_13685,N_13756);
xor UO_413 (O_413,N_14897,N_13868);
nand UO_414 (O_414,N_14030,N_14718);
and UO_415 (O_415,N_14412,N_13729);
nand UO_416 (O_416,N_13779,N_14065);
and UO_417 (O_417,N_13768,N_14414);
and UO_418 (O_418,N_13835,N_14735);
nor UO_419 (O_419,N_14581,N_13726);
and UO_420 (O_420,N_13623,N_13564);
nand UO_421 (O_421,N_14571,N_13903);
or UO_422 (O_422,N_14238,N_13605);
xor UO_423 (O_423,N_14622,N_14549);
nor UO_424 (O_424,N_14391,N_14898);
nand UO_425 (O_425,N_14261,N_14589);
nand UO_426 (O_426,N_14396,N_14489);
and UO_427 (O_427,N_14440,N_14000);
nor UO_428 (O_428,N_14309,N_14530);
and UO_429 (O_429,N_14772,N_13742);
or UO_430 (O_430,N_14164,N_14393);
or UO_431 (O_431,N_14623,N_14465);
nand UO_432 (O_432,N_14352,N_14857);
nor UO_433 (O_433,N_14886,N_13785);
or UO_434 (O_434,N_14468,N_13515);
or UO_435 (O_435,N_14535,N_14282);
nand UO_436 (O_436,N_14307,N_14285);
xor UO_437 (O_437,N_14124,N_14488);
or UO_438 (O_438,N_14914,N_14504);
and UO_439 (O_439,N_14424,N_14421);
or UO_440 (O_440,N_13514,N_13795);
nand UO_441 (O_441,N_13637,N_14868);
and UO_442 (O_442,N_14191,N_14578);
nand UO_443 (O_443,N_13585,N_14308);
nor UO_444 (O_444,N_14687,N_14186);
nor UO_445 (O_445,N_14519,N_13607);
nand UO_446 (O_446,N_13587,N_13526);
or UO_447 (O_447,N_13749,N_14045);
and UO_448 (O_448,N_13590,N_14562);
or UO_449 (O_449,N_13546,N_14316);
and UO_450 (O_450,N_13767,N_13811);
nor UO_451 (O_451,N_13645,N_13624);
or UO_452 (O_452,N_13933,N_14133);
nor UO_453 (O_453,N_14816,N_13971);
and UO_454 (O_454,N_14631,N_14063);
nand UO_455 (O_455,N_14763,N_13860);
and UO_456 (O_456,N_13715,N_13984);
nor UO_457 (O_457,N_14507,N_13973);
xnor UO_458 (O_458,N_13544,N_13917);
nor UO_459 (O_459,N_14952,N_14847);
or UO_460 (O_460,N_14101,N_14314);
nand UO_461 (O_461,N_14009,N_14312);
or UO_462 (O_462,N_13961,N_14438);
nand UO_463 (O_463,N_14251,N_14906);
or UO_464 (O_464,N_13627,N_13554);
nor UO_465 (O_465,N_14076,N_13690);
xnor UO_466 (O_466,N_13719,N_14931);
and UO_467 (O_467,N_14038,N_13888);
or UO_468 (O_468,N_13974,N_14005);
nor UO_469 (O_469,N_14806,N_13626);
nand UO_470 (O_470,N_13806,N_14148);
nand UO_471 (O_471,N_14751,N_14922);
nand UO_472 (O_472,N_13735,N_14322);
and UO_473 (O_473,N_14907,N_13653);
or UO_474 (O_474,N_14061,N_14430);
or UO_475 (O_475,N_14680,N_14574);
xnor UO_476 (O_476,N_13843,N_13700);
and UO_477 (O_477,N_14362,N_14645);
or UO_478 (O_478,N_13738,N_13745);
or UO_479 (O_479,N_13567,N_14899);
nand UO_480 (O_480,N_14443,N_14698);
nor UO_481 (O_481,N_14823,N_14876);
nand UO_482 (O_482,N_14388,N_14642);
or UO_483 (O_483,N_13712,N_14435);
xnor UO_484 (O_484,N_14206,N_14018);
or UO_485 (O_485,N_14788,N_14807);
or UO_486 (O_486,N_14083,N_13539);
nand UO_487 (O_487,N_14880,N_14606);
or UO_488 (O_488,N_14584,N_14416);
nor UO_489 (O_489,N_13920,N_13832);
or UO_490 (O_490,N_14593,N_13647);
xor UO_491 (O_491,N_14104,N_14627);
nand UO_492 (O_492,N_14473,N_14137);
nor UO_493 (O_493,N_13981,N_13734);
and UO_494 (O_494,N_14159,N_13603);
nor UO_495 (O_495,N_14709,N_13878);
or UO_496 (O_496,N_14955,N_13584);
xnor UO_497 (O_497,N_14831,N_14275);
and UO_498 (O_498,N_14644,N_13660);
nand UO_499 (O_499,N_14970,N_14495);
and UO_500 (O_500,N_14597,N_14174);
and UO_501 (O_501,N_14448,N_14616);
and UO_502 (O_502,N_14434,N_14712);
and UO_503 (O_503,N_14121,N_14445);
nand UO_504 (O_504,N_14746,N_14103);
nor UO_505 (O_505,N_13573,N_13834);
nand UO_506 (O_506,N_14046,N_14188);
xor UO_507 (O_507,N_14621,N_14048);
nand UO_508 (O_508,N_14277,N_13943);
nor UO_509 (O_509,N_13578,N_13820);
or UO_510 (O_510,N_13796,N_14640);
nor UO_511 (O_511,N_14647,N_14247);
or UO_512 (O_512,N_14651,N_14062);
and UO_513 (O_513,N_13663,N_14346);
nand UO_514 (O_514,N_14363,N_14118);
nand UO_515 (O_515,N_13686,N_13949);
nor UO_516 (O_516,N_13683,N_14491);
and UO_517 (O_517,N_14199,N_13845);
or UO_518 (O_518,N_13565,N_14417);
xor UO_519 (O_519,N_14298,N_14888);
nor UO_520 (O_520,N_14330,N_13839);
or UO_521 (O_521,N_14521,N_13733);
xor UO_522 (O_522,N_14153,N_14548);
nor UO_523 (O_523,N_14686,N_14662);
nand UO_524 (O_524,N_14951,N_14659);
nand UO_525 (O_525,N_14959,N_14699);
nand UO_526 (O_526,N_13574,N_14526);
nor UO_527 (O_527,N_14918,N_14688);
nor UO_528 (O_528,N_14144,N_13651);
nand UO_529 (O_529,N_13991,N_13643);
and UO_530 (O_530,N_13872,N_13560);
or UO_531 (O_531,N_13758,N_14132);
and UO_532 (O_532,N_13713,N_14961);
and UO_533 (O_533,N_14458,N_14394);
xnor UO_534 (O_534,N_13662,N_14615);
and UO_535 (O_535,N_14456,N_13659);
nand UO_536 (O_536,N_13503,N_14919);
or UO_537 (O_537,N_13523,N_14538);
nand UO_538 (O_538,N_14720,N_14802);
or UO_539 (O_539,N_14273,N_14354);
and UO_540 (O_540,N_13601,N_14639);
xnor UO_541 (O_541,N_14990,N_14901);
or UO_542 (O_542,N_14629,N_14114);
and UO_543 (O_543,N_14859,N_14289);
nor UO_544 (O_544,N_14207,N_13849);
or UO_545 (O_545,N_14320,N_13996);
and UO_546 (O_546,N_14937,N_14336);
nor UO_547 (O_547,N_13672,N_14082);
nand UO_548 (O_548,N_13569,N_13641);
nand UO_549 (O_549,N_13580,N_14799);
nor UO_550 (O_550,N_14654,N_13507);
and UO_551 (O_551,N_14797,N_14452);
nand UO_552 (O_552,N_14643,N_13818);
and UO_553 (O_553,N_13950,N_14269);
and UO_554 (O_554,N_14220,N_13711);
nor UO_555 (O_555,N_14175,N_14227);
nor UO_556 (O_556,N_14382,N_13723);
nand UO_557 (O_557,N_14286,N_14231);
or UO_558 (O_558,N_14327,N_14415);
nand UO_559 (O_559,N_13671,N_14829);
nor UO_560 (O_560,N_14777,N_14134);
and UO_561 (O_561,N_13904,N_14108);
or UO_562 (O_562,N_13549,N_14271);
and UO_563 (O_563,N_13844,N_13946);
and UO_564 (O_564,N_13953,N_14411);
nor UO_565 (O_565,N_13976,N_13913);
xor UO_566 (O_566,N_14547,N_13910);
nor UO_567 (O_567,N_13640,N_14232);
or UO_568 (O_568,N_13600,N_14858);
nand UO_569 (O_569,N_14311,N_14453);
nand UO_570 (O_570,N_14773,N_14284);
nand UO_571 (O_571,N_14845,N_14147);
nand UO_572 (O_572,N_13614,N_14234);
nand UO_573 (O_573,N_14328,N_14258);
or UO_574 (O_574,N_13593,N_14617);
nand UO_575 (O_575,N_14233,N_14432);
or UO_576 (O_576,N_14152,N_14976);
xor UO_577 (O_577,N_14049,N_14975);
and UO_578 (O_578,N_14026,N_14820);
or UO_579 (O_579,N_14539,N_14230);
and UO_580 (O_580,N_14711,N_14982);
or UO_581 (O_581,N_14405,N_14784);
xor UO_582 (O_582,N_14472,N_14367);
and UO_583 (O_583,N_13757,N_14941);
nor UO_584 (O_584,N_13859,N_13776);
and UO_585 (O_585,N_13804,N_13780);
nand UO_586 (O_586,N_13783,N_13799);
nor UO_587 (O_587,N_14449,N_13959);
or UO_588 (O_588,N_14546,N_14509);
nor UO_589 (O_589,N_14290,N_14588);
or UO_590 (O_590,N_13992,N_14392);
nand UO_591 (O_591,N_14106,N_14278);
or UO_592 (O_592,N_13535,N_13801);
and UO_593 (O_593,N_14700,N_14544);
and UO_594 (O_594,N_13980,N_14022);
nor UO_595 (O_595,N_14454,N_14826);
nor UO_596 (O_596,N_14241,N_13531);
and UO_597 (O_597,N_14554,N_14814);
nand UO_598 (O_598,N_14015,N_14168);
xor UO_599 (O_599,N_14863,N_13558);
nor UO_600 (O_600,N_14016,N_13778);
and UO_601 (O_601,N_13550,N_14668);
and UO_602 (O_602,N_14257,N_14953);
or UO_603 (O_603,N_14196,N_13571);
xnor UO_604 (O_604,N_13966,N_14385);
or UO_605 (O_605,N_14587,N_14582);
and UO_606 (O_606,N_14805,N_13886);
or UO_607 (O_607,N_13826,N_14564);
nor UO_608 (O_608,N_14690,N_14051);
xor UO_609 (O_609,N_14966,N_13510);
nor UO_610 (O_610,N_14964,N_14696);
or UO_611 (O_611,N_14706,N_14058);
nor UO_612 (O_612,N_14726,N_14243);
or UO_613 (O_613,N_14079,N_14305);
and UO_614 (O_614,N_13694,N_13751);
and UO_615 (O_615,N_13978,N_14861);
nand UO_616 (O_616,N_14140,N_14410);
or UO_617 (O_617,N_14028,N_14291);
nor UO_618 (O_618,N_13604,N_14691);
nand UO_619 (O_619,N_13702,N_14156);
nand UO_620 (O_620,N_14351,N_14479);
or UO_621 (O_621,N_14996,N_14739);
nand UO_622 (O_622,N_13591,N_14873);
nand UO_623 (O_623,N_14605,N_14950);
nor UO_624 (O_624,N_14272,N_14425);
nand UO_625 (O_625,N_14429,N_14531);
and UO_626 (O_626,N_14487,N_14808);
or UO_627 (O_627,N_13857,N_13833);
or UO_628 (O_628,N_14130,N_13866);
xnor UO_629 (O_629,N_14212,N_14929);
and UO_630 (O_630,N_14318,N_14569);
and UO_631 (O_631,N_14576,N_13958);
or UO_632 (O_632,N_14306,N_14205);
nor UO_633 (O_633,N_13658,N_14283);
nor UO_634 (O_634,N_13589,N_13710);
nand UO_635 (O_635,N_13732,N_14551);
and UO_636 (O_636,N_14242,N_14078);
and UO_637 (O_637,N_13633,N_14926);
or UO_638 (O_638,N_14444,N_14778);
and UO_639 (O_639,N_14123,N_13635);
nand UO_640 (O_640,N_13869,N_14386);
or UO_641 (O_641,N_13884,N_13951);
and UO_642 (O_642,N_14601,N_14214);
or UO_643 (O_643,N_14540,N_14958);
or UO_644 (O_644,N_13997,N_14280);
and UO_645 (O_645,N_14399,N_14791);
or UO_646 (O_646,N_14545,N_14723);
nor UO_647 (O_647,N_13597,N_14885);
nor UO_648 (O_648,N_14461,N_14228);
nand UO_649 (O_649,N_13983,N_14832);
or UO_650 (O_650,N_13919,N_14870);
nor UO_651 (O_651,N_14225,N_14853);
and UO_652 (O_652,N_13506,N_14650);
nor UO_653 (O_653,N_13985,N_14938);
or UO_654 (O_654,N_14301,N_14882);
nor UO_655 (O_655,N_14585,N_14377);
nand UO_656 (O_656,N_14056,N_14566);
nand UO_657 (O_657,N_13517,N_13854);
xor UO_658 (O_658,N_13714,N_14733);
nand UO_659 (O_659,N_14534,N_14742);
nand UO_660 (O_660,N_14945,N_13548);
or UO_661 (O_661,N_13617,N_13684);
nor UO_662 (O_662,N_14932,N_14501);
xor UO_663 (O_663,N_14908,N_13802);
nor UO_664 (O_664,N_14986,N_14120);
nand UO_665 (O_665,N_13969,N_13879);
nand UO_666 (O_666,N_14226,N_13852);
nor UO_667 (O_667,N_14989,N_14040);
and UO_668 (O_668,N_13691,N_14761);
nor UO_669 (O_669,N_14903,N_13787);
and UO_670 (O_670,N_14795,N_13520);
nand UO_671 (O_671,N_14210,N_13701);
nand UO_672 (O_672,N_14155,N_13760);
and UO_673 (O_673,N_14756,N_14939);
nor UO_674 (O_674,N_13764,N_14478);
nand UO_675 (O_675,N_14139,N_14946);
nand UO_676 (O_676,N_13508,N_13847);
nor UO_677 (O_677,N_14375,N_14933);
nor UO_678 (O_678,N_13960,N_14740);
nor UO_679 (O_679,N_14728,N_13914);
nand UO_680 (O_680,N_14127,N_13944);
xnor UO_681 (O_681,N_14747,N_13896);
nor UO_682 (O_682,N_13792,N_13631);
nor UO_683 (O_683,N_14128,N_14741);
and UO_684 (O_684,N_14874,N_14641);
and UO_685 (O_685,N_14890,N_14505);
nor UO_686 (O_686,N_14676,N_13707);
nor UO_687 (O_687,N_13885,N_14268);
and UO_688 (O_688,N_13929,N_13646);
and UO_689 (O_689,N_13998,N_13621);
or UO_690 (O_690,N_13693,N_13918);
and UO_691 (O_691,N_14866,N_14921);
or UO_692 (O_692,N_14303,N_14390);
xor UO_693 (O_693,N_14887,N_13543);
nor UO_694 (O_694,N_13703,N_13970);
xor UO_695 (O_695,N_13823,N_14098);
or UO_696 (O_696,N_13509,N_14782);
nor UO_697 (O_697,N_14867,N_13575);
xnor UO_698 (O_698,N_14503,N_14992);
xor UO_699 (O_699,N_14801,N_14944);
or UO_700 (O_700,N_13828,N_13762);
nand UO_701 (O_701,N_14930,N_13945);
and UO_702 (O_702,N_13541,N_14758);
nand UO_703 (O_703,N_14591,N_14023);
nand UO_704 (O_704,N_14081,N_13993);
nand UO_705 (O_705,N_14224,N_14781);
nand UO_706 (O_706,N_14648,N_14365);
or UO_707 (O_707,N_13800,N_14317);
nand UO_708 (O_708,N_13722,N_13551);
nor UO_709 (O_709,N_14948,N_13696);
nor UO_710 (O_710,N_14072,N_13895);
and UO_711 (O_711,N_14189,N_13570);
and UO_712 (O_712,N_14052,N_14057);
or UO_713 (O_713,N_13871,N_13670);
xnor UO_714 (O_714,N_14871,N_13865);
and UO_715 (O_715,N_14744,N_14656);
or UO_716 (O_716,N_14135,N_13650);
nor UO_717 (O_717,N_13665,N_14755);
and UO_718 (O_718,N_14889,N_14769);
nand UO_719 (O_719,N_14673,N_13699);
and UO_720 (O_720,N_13794,N_14204);
and UO_721 (O_721,N_13975,N_14850);
and UO_722 (O_722,N_14789,N_14295);
or UO_723 (O_723,N_13923,N_13808);
or UO_724 (O_724,N_14792,N_14113);
nor UO_725 (O_725,N_13586,N_13743);
nor UO_726 (O_726,N_14138,N_13664);
nor UO_727 (O_727,N_14379,N_14093);
and UO_728 (O_728,N_14459,N_14916);
nor UO_729 (O_729,N_14864,N_14183);
or UO_730 (O_730,N_14892,N_14555);
or UO_731 (O_731,N_14402,N_14753);
nand UO_732 (O_732,N_14550,N_14292);
nor UO_733 (O_733,N_14794,N_13867);
nor UO_734 (O_734,N_14350,N_13875);
nand UO_735 (O_735,N_14163,N_14760);
and UO_736 (O_736,N_13874,N_14835);
nor UO_737 (O_737,N_14987,N_14660);
nor UO_738 (O_738,N_13706,N_14663);
or UO_739 (O_739,N_14494,N_13899);
nor UO_740 (O_740,N_13727,N_14427);
nand UO_741 (O_741,N_14006,N_14767);
nor UO_742 (O_742,N_14446,N_14387);
nand UO_743 (O_743,N_13747,N_14869);
nand UO_744 (O_744,N_13793,N_13815);
xnor UO_745 (O_745,N_14851,N_14024);
nand UO_746 (O_746,N_13599,N_14824);
xnor UO_747 (O_747,N_13504,N_14097);
xnor UO_748 (O_748,N_13902,N_14219);
and UO_749 (O_749,N_13922,N_14131);
xnor UO_750 (O_750,N_14036,N_14083);
or UO_751 (O_751,N_14888,N_14186);
or UO_752 (O_752,N_14387,N_14412);
nor UO_753 (O_753,N_14079,N_14942);
nand UO_754 (O_754,N_13637,N_13681);
and UO_755 (O_755,N_14160,N_14179);
or UO_756 (O_756,N_13625,N_14817);
and UO_757 (O_757,N_14241,N_14208);
nand UO_758 (O_758,N_14986,N_14367);
and UO_759 (O_759,N_14236,N_14109);
xnor UO_760 (O_760,N_14480,N_14595);
nand UO_761 (O_761,N_14737,N_13525);
nor UO_762 (O_762,N_14813,N_14314);
and UO_763 (O_763,N_14607,N_13784);
nand UO_764 (O_764,N_13538,N_13996);
xor UO_765 (O_765,N_14709,N_14008);
and UO_766 (O_766,N_14315,N_13896);
and UO_767 (O_767,N_13949,N_14913);
and UO_768 (O_768,N_14059,N_13515);
nor UO_769 (O_769,N_14407,N_13503);
nand UO_770 (O_770,N_13921,N_14311);
nor UO_771 (O_771,N_14109,N_13648);
nor UO_772 (O_772,N_14818,N_13850);
nor UO_773 (O_773,N_13583,N_14749);
nand UO_774 (O_774,N_14219,N_13541);
nand UO_775 (O_775,N_13790,N_14254);
xor UO_776 (O_776,N_14153,N_14925);
or UO_777 (O_777,N_14957,N_13994);
or UO_778 (O_778,N_14963,N_13905);
or UO_779 (O_779,N_14182,N_14857);
or UO_780 (O_780,N_14337,N_13891);
xnor UO_781 (O_781,N_14817,N_14009);
nor UO_782 (O_782,N_13672,N_13818);
xor UO_783 (O_783,N_13666,N_13534);
nand UO_784 (O_784,N_14736,N_13713);
and UO_785 (O_785,N_13720,N_13690);
and UO_786 (O_786,N_13984,N_13737);
and UO_787 (O_787,N_14508,N_13924);
nor UO_788 (O_788,N_14983,N_13626);
and UO_789 (O_789,N_14852,N_14501);
xor UO_790 (O_790,N_13790,N_14947);
and UO_791 (O_791,N_14815,N_14704);
or UO_792 (O_792,N_14883,N_13727);
and UO_793 (O_793,N_14830,N_13670);
xnor UO_794 (O_794,N_14523,N_13614);
nand UO_795 (O_795,N_14746,N_14813);
nand UO_796 (O_796,N_13694,N_13980);
or UO_797 (O_797,N_14052,N_13556);
xnor UO_798 (O_798,N_14695,N_14816);
xor UO_799 (O_799,N_14248,N_14067);
and UO_800 (O_800,N_13692,N_13818);
or UO_801 (O_801,N_14842,N_13622);
nand UO_802 (O_802,N_14117,N_13899);
or UO_803 (O_803,N_14931,N_14446);
nand UO_804 (O_804,N_14470,N_14812);
or UO_805 (O_805,N_13826,N_14461);
or UO_806 (O_806,N_14641,N_13838);
and UO_807 (O_807,N_14005,N_13583);
or UO_808 (O_808,N_14644,N_14568);
nand UO_809 (O_809,N_14659,N_13957);
xor UO_810 (O_810,N_14598,N_13865);
nand UO_811 (O_811,N_14125,N_14640);
xnor UO_812 (O_812,N_13899,N_14570);
and UO_813 (O_813,N_13904,N_13536);
or UO_814 (O_814,N_14316,N_14283);
and UO_815 (O_815,N_13653,N_13561);
or UO_816 (O_816,N_13650,N_14884);
nand UO_817 (O_817,N_13914,N_13765);
or UO_818 (O_818,N_14368,N_13876);
nand UO_819 (O_819,N_13508,N_14180);
and UO_820 (O_820,N_14594,N_14060);
and UO_821 (O_821,N_14637,N_14344);
nor UO_822 (O_822,N_14222,N_14416);
and UO_823 (O_823,N_14011,N_14995);
and UO_824 (O_824,N_13903,N_14219);
or UO_825 (O_825,N_14612,N_13932);
nor UO_826 (O_826,N_13991,N_14306);
nand UO_827 (O_827,N_14557,N_14099);
and UO_828 (O_828,N_14010,N_14158);
and UO_829 (O_829,N_13600,N_13750);
nor UO_830 (O_830,N_14211,N_13696);
nor UO_831 (O_831,N_14269,N_13971);
nor UO_832 (O_832,N_13601,N_14643);
nand UO_833 (O_833,N_13913,N_14900);
nor UO_834 (O_834,N_13833,N_13863);
nor UO_835 (O_835,N_14324,N_14208);
or UO_836 (O_836,N_14504,N_14289);
and UO_837 (O_837,N_14218,N_13631);
or UO_838 (O_838,N_13635,N_14525);
and UO_839 (O_839,N_14394,N_14876);
nor UO_840 (O_840,N_13926,N_14532);
nor UO_841 (O_841,N_14377,N_14436);
and UO_842 (O_842,N_14453,N_14528);
nor UO_843 (O_843,N_14350,N_14653);
and UO_844 (O_844,N_13559,N_14449);
nor UO_845 (O_845,N_14765,N_14745);
xor UO_846 (O_846,N_14644,N_14704);
or UO_847 (O_847,N_13848,N_13632);
nand UO_848 (O_848,N_14646,N_14114);
nor UO_849 (O_849,N_14543,N_14224);
or UO_850 (O_850,N_14487,N_14278);
and UO_851 (O_851,N_14719,N_14093);
or UO_852 (O_852,N_14400,N_14388);
xor UO_853 (O_853,N_14687,N_14415);
nor UO_854 (O_854,N_13637,N_13922);
or UO_855 (O_855,N_14185,N_14036);
or UO_856 (O_856,N_14620,N_13829);
nand UO_857 (O_857,N_13942,N_14101);
nor UO_858 (O_858,N_14445,N_14855);
or UO_859 (O_859,N_14088,N_13683);
nor UO_860 (O_860,N_14744,N_14988);
nor UO_861 (O_861,N_13599,N_13999);
nor UO_862 (O_862,N_14653,N_13515);
or UO_863 (O_863,N_14906,N_14217);
and UO_864 (O_864,N_14619,N_14748);
nor UO_865 (O_865,N_14695,N_14392);
xnor UO_866 (O_866,N_14638,N_14791);
nand UO_867 (O_867,N_14259,N_14852);
and UO_868 (O_868,N_13751,N_13779);
or UO_869 (O_869,N_14340,N_13579);
and UO_870 (O_870,N_13938,N_13592);
or UO_871 (O_871,N_13531,N_14824);
nor UO_872 (O_872,N_13697,N_14888);
nor UO_873 (O_873,N_13573,N_14787);
nor UO_874 (O_874,N_13536,N_13629);
or UO_875 (O_875,N_14152,N_14944);
or UO_876 (O_876,N_14211,N_14656);
or UO_877 (O_877,N_14652,N_14255);
or UO_878 (O_878,N_14607,N_14662);
and UO_879 (O_879,N_14893,N_13749);
and UO_880 (O_880,N_13951,N_14447);
nand UO_881 (O_881,N_13556,N_14913);
or UO_882 (O_882,N_14059,N_14923);
and UO_883 (O_883,N_13715,N_14923);
and UO_884 (O_884,N_14978,N_13774);
xor UO_885 (O_885,N_14651,N_14627);
and UO_886 (O_886,N_14999,N_13700);
or UO_887 (O_887,N_14751,N_14100);
xor UO_888 (O_888,N_14824,N_13905);
or UO_889 (O_889,N_14054,N_13962);
nor UO_890 (O_890,N_14727,N_14135);
xnor UO_891 (O_891,N_13659,N_14473);
and UO_892 (O_892,N_14026,N_14675);
or UO_893 (O_893,N_13861,N_13873);
nor UO_894 (O_894,N_14129,N_14788);
or UO_895 (O_895,N_14149,N_13531);
nand UO_896 (O_896,N_13726,N_14870);
nor UO_897 (O_897,N_14426,N_14675);
and UO_898 (O_898,N_14117,N_13582);
or UO_899 (O_899,N_14170,N_13565);
or UO_900 (O_900,N_14123,N_14979);
xnor UO_901 (O_901,N_13866,N_13970);
and UO_902 (O_902,N_14313,N_13936);
nand UO_903 (O_903,N_14550,N_14178);
or UO_904 (O_904,N_14937,N_13557);
or UO_905 (O_905,N_14780,N_14420);
nand UO_906 (O_906,N_14327,N_13628);
nor UO_907 (O_907,N_14490,N_14179);
nand UO_908 (O_908,N_13521,N_14099);
nand UO_909 (O_909,N_13841,N_13752);
nand UO_910 (O_910,N_14418,N_14037);
nor UO_911 (O_911,N_13504,N_13726);
or UO_912 (O_912,N_13538,N_14076);
xor UO_913 (O_913,N_14382,N_13588);
nor UO_914 (O_914,N_13917,N_14712);
or UO_915 (O_915,N_14592,N_14824);
or UO_916 (O_916,N_14082,N_14631);
nand UO_917 (O_917,N_13620,N_14685);
nor UO_918 (O_918,N_14880,N_14638);
or UO_919 (O_919,N_13752,N_14045);
or UO_920 (O_920,N_13641,N_14585);
and UO_921 (O_921,N_13942,N_13837);
nor UO_922 (O_922,N_13520,N_13947);
or UO_923 (O_923,N_14815,N_14386);
and UO_924 (O_924,N_13784,N_13565);
nand UO_925 (O_925,N_14715,N_14225);
xor UO_926 (O_926,N_13906,N_13790);
and UO_927 (O_927,N_13570,N_13896);
nand UO_928 (O_928,N_13977,N_14509);
nor UO_929 (O_929,N_13540,N_14430);
xor UO_930 (O_930,N_14793,N_13899);
or UO_931 (O_931,N_13597,N_13985);
nand UO_932 (O_932,N_14856,N_14134);
or UO_933 (O_933,N_14756,N_14807);
nor UO_934 (O_934,N_14727,N_14703);
and UO_935 (O_935,N_13959,N_14690);
nor UO_936 (O_936,N_14855,N_14266);
nand UO_937 (O_937,N_14223,N_13530);
nand UO_938 (O_938,N_13806,N_14210);
or UO_939 (O_939,N_14143,N_14664);
or UO_940 (O_940,N_14938,N_14727);
nand UO_941 (O_941,N_14133,N_14423);
nand UO_942 (O_942,N_13586,N_14095);
nand UO_943 (O_943,N_14954,N_13745);
or UO_944 (O_944,N_14418,N_13835);
and UO_945 (O_945,N_14049,N_13702);
nor UO_946 (O_946,N_14556,N_14544);
nand UO_947 (O_947,N_14564,N_14727);
or UO_948 (O_948,N_14122,N_14123);
or UO_949 (O_949,N_13983,N_14820);
nor UO_950 (O_950,N_13731,N_14163);
or UO_951 (O_951,N_13808,N_14274);
and UO_952 (O_952,N_13777,N_14125);
xnor UO_953 (O_953,N_14547,N_14600);
and UO_954 (O_954,N_13510,N_14575);
nand UO_955 (O_955,N_14438,N_14459);
and UO_956 (O_956,N_14966,N_14891);
nand UO_957 (O_957,N_14939,N_13795);
xor UO_958 (O_958,N_14506,N_13808);
and UO_959 (O_959,N_14581,N_13958);
xor UO_960 (O_960,N_14395,N_14251);
nand UO_961 (O_961,N_14207,N_13594);
nor UO_962 (O_962,N_14505,N_14785);
or UO_963 (O_963,N_14520,N_14765);
and UO_964 (O_964,N_14173,N_14589);
nor UO_965 (O_965,N_14771,N_14826);
and UO_966 (O_966,N_14267,N_14973);
nor UO_967 (O_967,N_14058,N_13607);
nand UO_968 (O_968,N_14401,N_14125);
nor UO_969 (O_969,N_14511,N_14925);
xor UO_970 (O_970,N_14948,N_14488);
nand UO_971 (O_971,N_14065,N_13729);
nand UO_972 (O_972,N_13852,N_14874);
or UO_973 (O_973,N_14765,N_14822);
nor UO_974 (O_974,N_14517,N_13979);
or UO_975 (O_975,N_14455,N_14676);
nand UO_976 (O_976,N_14819,N_13558);
and UO_977 (O_977,N_14388,N_14751);
xor UO_978 (O_978,N_14718,N_14815);
and UO_979 (O_979,N_14180,N_14748);
and UO_980 (O_980,N_13563,N_13864);
and UO_981 (O_981,N_14379,N_14951);
nor UO_982 (O_982,N_14093,N_14035);
or UO_983 (O_983,N_14523,N_13588);
nand UO_984 (O_984,N_14935,N_14143);
nand UO_985 (O_985,N_14011,N_13729);
or UO_986 (O_986,N_14283,N_14057);
and UO_987 (O_987,N_14409,N_14167);
nor UO_988 (O_988,N_14556,N_14671);
nor UO_989 (O_989,N_14781,N_14308);
nor UO_990 (O_990,N_13683,N_13544);
nand UO_991 (O_991,N_13730,N_14823);
nand UO_992 (O_992,N_14462,N_13821);
nand UO_993 (O_993,N_14960,N_13781);
nand UO_994 (O_994,N_14286,N_14782);
nor UO_995 (O_995,N_14161,N_14639);
nand UO_996 (O_996,N_14118,N_13582);
xor UO_997 (O_997,N_13529,N_14079);
or UO_998 (O_998,N_14530,N_14457);
nand UO_999 (O_999,N_13754,N_14891);
nor UO_1000 (O_1000,N_14270,N_14541);
xor UO_1001 (O_1001,N_13535,N_13984);
nor UO_1002 (O_1002,N_13574,N_14020);
nor UO_1003 (O_1003,N_14185,N_14861);
nor UO_1004 (O_1004,N_14095,N_14300);
nor UO_1005 (O_1005,N_14306,N_14391);
nand UO_1006 (O_1006,N_14532,N_13836);
and UO_1007 (O_1007,N_13735,N_14921);
nor UO_1008 (O_1008,N_14498,N_14389);
and UO_1009 (O_1009,N_14293,N_14290);
and UO_1010 (O_1010,N_14413,N_14972);
or UO_1011 (O_1011,N_14315,N_14939);
xor UO_1012 (O_1012,N_14493,N_13801);
or UO_1013 (O_1013,N_14984,N_14360);
nand UO_1014 (O_1014,N_14397,N_14812);
nand UO_1015 (O_1015,N_14971,N_13770);
or UO_1016 (O_1016,N_14819,N_14452);
and UO_1017 (O_1017,N_13682,N_13904);
nand UO_1018 (O_1018,N_14862,N_14135);
nand UO_1019 (O_1019,N_13653,N_13987);
or UO_1020 (O_1020,N_14326,N_14576);
or UO_1021 (O_1021,N_13575,N_14399);
or UO_1022 (O_1022,N_13713,N_13948);
and UO_1023 (O_1023,N_14489,N_13627);
nor UO_1024 (O_1024,N_13805,N_14919);
nor UO_1025 (O_1025,N_13831,N_14620);
nand UO_1026 (O_1026,N_14546,N_14276);
or UO_1027 (O_1027,N_14998,N_14898);
nand UO_1028 (O_1028,N_14134,N_14848);
and UO_1029 (O_1029,N_14216,N_14552);
or UO_1030 (O_1030,N_13610,N_14282);
nand UO_1031 (O_1031,N_13549,N_14034);
nor UO_1032 (O_1032,N_14730,N_14985);
and UO_1033 (O_1033,N_14680,N_13628);
nor UO_1034 (O_1034,N_14134,N_13511);
and UO_1035 (O_1035,N_13641,N_14481);
and UO_1036 (O_1036,N_14637,N_13780);
and UO_1037 (O_1037,N_14879,N_14883);
xor UO_1038 (O_1038,N_14009,N_13984);
and UO_1039 (O_1039,N_14754,N_14331);
nand UO_1040 (O_1040,N_13964,N_14549);
nor UO_1041 (O_1041,N_14285,N_14171);
nand UO_1042 (O_1042,N_14053,N_14152);
nand UO_1043 (O_1043,N_14466,N_14351);
nor UO_1044 (O_1044,N_13849,N_13985);
nor UO_1045 (O_1045,N_14802,N_14029);
nand UO_1046 (O_1046,N_14660,N_14818);
nand UO_1047 (O_1047,N_13661,N_14659);
or UO_1048 (O_1048,N_14954,N_13947);
nor UO_1049 (O_1049,N_14896,N_14521);
nand UO_1050 (O_1050,N_13690,N_13511);
and UO_1051 (O_1051,N_13643,N_14572);
nor UO_1052 (O_1052,N_14117,N_14300);
nor UO_1053 (O_1053,N_14959,N_13763);
nor UO_1054 (O_1054,N_14044,N_14550);
nor UO_1055 (O_1055,N_14182,N_14129);
or UO_1056 (O_1056,N_13743,N_13572);
nor UO_1057 (O_1057,N_13748,N_13506);
nor UO_1058 (O_1058,N_14871,N_14014);
and UO_1059 (O_1059,N_14786,N_14156);
or UO_1060 (O_1060,N_14714,N_14619);
nand UO_1061 (O_1061,N_13560,N_14224);
nand UO_1062 (O_1062,N_14047,N_13635);
nand UO_1063 (O_1063,N_14505,N_13770);
xnor UO_1064 (O_1064,N_14292,N_13741);
nand UO_1065 (O_1065,N_14731,N_13997);
and UO_1066 (O_1066,N_14254,N_14186);
or UO_1067 (O_1067,N_14741,N_14400);
and UO_1068 (O_1068,N_14196,N_13720);
and UO_1069 (O_1069,N_14175,N_13857);
xnor UO_1070 (O_1070,N_14454,N_13701);
nand UO_1071 (O_1071,N_14625,N_14285);
nor UO_1072 (O_1072,N_14734,N_14932);
and UO_1073 (O_1073,N_13529,N_13900);
and UO_1074 (O_1074,N_13957,N_14290);
xor UO_1075 (O_1075,N_13508,N_14713);
nor UO_1076 (O_1076,N_13734,N_14029);
or UO_1077 (O_1077,N_13879,N_14834);
nor UO_1078 (O_1078,N_13990,N_13626);
xnor UO_1079 (O_1079,N_14782,N_13953);
nor UO_1080 (O_1080,N_14658,N_14502);
nand UO_1081 (O_1081,N_14101,N_14002);
nand UO_1082 (O_1082,N_13798,N_14533);
xor UO_1083 (O_1083,N_14939,N_14410);
or UO_1084 (O_1084,N_13648,N_14787);
and UO_1085 (O_1085,N_13635,N_13582);
nand UO_1086 (O_1086,N_13530,N_13558);
or UO_1087 (O_1087,N_14387,N_14576);
xnor UO_1088 (O_1088,N_13878,N_13785);
and UO_1089 (O_1089,N_14748,N_14277);
nor UO_1090 (O_1090,N_14946,N_14813);
nor UO_1091 (O_1091,N_14220,N_13790);
or UO_1092 (O_1092,N_14144,N_14147);
nand UO_1093 (O_1093,N_14671,N_14654);
and UO_1094 (O_1094,N_14815,N_14844);
nand UO_1095 (O_1095,N_14054,N_13691);
nor UO_1096 (O_1096,N_14637,N_14964);
or UO_1097 (O_1097,N_14850,N_13553);
nor UO_1098 (O_1098,N_13703,N_14604);
and UO_1099 (O_1099,N_13689,N_14796);
nor UO_1100 (O_1100,N_14973,N_14758);
or UO_1101 (O_1101,N_14511,N_14291);
nor UO_1102 (O_1102,N_14915,N_14083);
nand UO_1103 (O_1103,N_13990,N_14365);
or UO_1104 (O_1104,N_14523,N_14957);
nand UO_1105 (O_1105,N_13684,N_14463);
nand UO_1106 (O_1106,N_13661,N_13749);
nand UO_1107 (O_1107,N_14758,N_14823);
or UO_1108 (O_1108,N_13853,N_14154);
or UO_1109 (O_1109,N_14566,N_13606);
or UO_1110 (O_1110,N_14183,N_13887);
nor UO_1111 (O_1111,N_13688,N_14018);
or UO_1112 (O_1112,N_14037,N_14009);
or UO_1113 (O_1113,N_13640,N_14330);
nor UO_1114 (O_1114,N_14315,N_13873);
nor UO_1115 (O_1115,N_14081,N_14307);
or UO_1116 (O_1116,N_13660,N_13789);
xor UO_1117 (O_1117,N_14781,N_14169);
xor UO_1118 (O_1118,N_13564,N_14038);
xor UO_1119 (O_1119,N_14168,N_14060);
nor UO_1120 (O_1120,N_13904,N_14908);
nand UO_1121 (O_1121,N_13684,N_14389);
or UO_1122 (O_1122,N_14634,N_13563);
nand UO_1123 (O_1123,N_14454,N_14061);
and UO_1124 (O_1124,N_14537,N_13956);
nor UO_1125 (O_1125,N_14249,N_13929);
xor UO_1126 (O_1126,N_13745,N_14739);
nor UO_1127 (O_1127,N_14397,N_14764);
nand UO_1128 (O_1128,N_14598,N_14038);
nor UO_1129 (O_1129,N_14531,N_13502);
nand UO_1130 (O_1130,N_14893,N_13694);
and UO_1131 (O_1131,N_14917,N_14733);
nand UO_1132 (O_1132,N_13967,N_14199);
nor UO_1133 (O_1133,N_14473,N_13724);
nand UO_1134 (O_1134,N_14006,N_14819);
nor UO_1135 (O_1135,N_13879,N_14605);
and UO_1136 (O_1136,N_13713,N_14551);
nand UO_1137 (O_1137,N_14770,N_14531);
nor UO_1138 (O_1138,N_13524,N_13674);
nand UO_1139 (O_1139,N_13916,N_14907);
nand UO_1140 (O_1140,N_14219,N_13866);
nor UO_1141 (O_1141,N_13518,N_14774);
xnor UO_1142 (O_1142,N_14156,N_13835);
nor UO_1143 (O_1143,N_14978,N_14960);
nor UO_1144 (O_1144,N_14998,N_14294);
nor UO_1145 (O_1145,N_13601,N_13604);
nor UO_1146 (O_1146,N_14609,N_14593);
or UO_1147 (O_1147,N_14755,N_14048);
or UO_1148 (O_1148,N_14897,N_13803);
nor UO_1149 (O_1149,N_13512,N_14632);
or UO_1150 (O_1150,N_13811,N_14881);
and UO_1151 (O_1151,N_14140,N_14674);
xnor UO_1152 (O_1152,N_13684,N_13891);
nand UO_1153 (O_1153,N_13950,N_13573);
and UO_1154 (O_1154,N_14413,N_14612);
or UO_1155 (O_1155,N_13771,N_14970);
and UO_1156 (O_1156,N_14204,N_14495);
nor UO_1157 (O_1157,N_13690,N_14436);
or UO_1158 (O_1158,N_13960,N_14492);
or UO_1159 (O_1159,N_13794,N_14968);
or UO_1160 (O_1160,N_14509,N_14094);
nor UO_1161 (O_1161,N_14647,N_14354);
nor UO_1162 (O_1162,N_14294,N_14863);
and UO_1163 (O_1163,N_13928,N_14694);
nor UO_1164 (O_1164,N_14716,N_14797);
and UO_1165 (O_1165,N_14743,N_14470);
and UO_1166 (O_1166,N_14494,N_13656);
or UO_1167 (O_1167,N_14605,N_14893);
nor UO_1168 (O_1168,N_14726,N_14715);
nor UO_1169 (O_1169,N_13555,N_14843);
nand UO_1170 (O_1170,N_13795,N_14557);
or UO_1171 (O_1171,N_14234,N_14365);
nand UO_1172 (O_1172,N_14127,N_14692);
nor UO_1173 (O_1173,N_13781,N_14391);
nor UO_1174 (O_1174,N_14923,N_14032);
nand UO_1175 (O_1175,N_13869,N_13806);
nor UO_1176 (O_1176,N_14405,N_14729);
xor UO_1177 (O_1177,N_14929,N_14462);
nor UO_1178 (O_1178,N_13554,N_14646);
nor UO_1179 (O_1179,N_13514,N_14685);
and UO_1180 (O_1180,N_13556,N_14512);
nand UO_1181 (O_1181,N_14501,N_14972);
or UO_1182 (O_1182,N_13708,N_13954);
or UO_1183 (O_1183,N_14577,N_14377);
or UO_1184 (O_1184,N_14264,N_14712);
and UO_1185 (O_1185,N_14714,N_14537);
or UO_1186 (O_1186,N_14619,N_14435);
nand UO_1187 (O_1187,N_13654,N_14758);
xnor UO_1188 (O_1188,N_13944,N_13705);
or UO_1189 (O_1189,N_14336,N_13629);
and UO_1190 (O_1190,N_14606,N_13756);
or UO_1191 (O_1191,N_14175,N_13664);
xor UO_1192 (O_1192,N_14469,N_14046);
nor UO_1193 (O_1193,N_14658,N_13807);
nor UO_1194 (O_1194,N_13889,N_14023);
nor UO_1195 (O_1195,N_13704,N_13834);
or UO_1196 (O_1196,N_14174,N_14946);
nor UO_1197 (O_1197,N_14496,N_14023);
or UO_1198 (O_1198,N_14189,N_14769);
or UO_1199 (O_1199,N_13724,N_14130);
or UO_1200 (O_1200,N_14328,N_13866);
and UO_1201 (O_1201,N_14072,N_14448);
and UO_1202 (O_1202,N_14640,N_14894);
nand UO_1203 (O_1203,N_13953,N_13957);
nor UO_1204 (O_1204,N_13772,N_14132);
nand UO_1205 (O_1205,N_13998,N_13592);
or UO_1206 (O_1206,N_14120,N_14918);
nor UO_1207 (O_1207,N_14166,N_13875);
and UO_1208 (O_1208,N_13622,N_14561);
nor UO_1209 (O_1209,N_13815,N_14396);
nor UO_1210 (O_1210,N_13575,N_14584);
and UO_1211 (O_1211,N_14031,N_14289);
and UO_1212 (O_1212,N_14472,N_14282);
xnor UO_1213 (O_1213,N_14616,N_14644);
and UO_1214 (O_1214,N_14551,N_13871);
nor UO_1215 (O_1215,N_14378,N_14668);
xor UO_1216 (O_1216,N_14591,N_14833);
or UO_1217 (O_1217,N_14140,N_14943);
xnor UO_1218 (O_1218,N_13531,N_14551);
and UO_1219 (O_1219,N_13679,N_14120);
nand UO_1220 (O_1220,N_14455,N_14498);
or UO_1221 (O_1221,N_13539,N_14615);
or UO_1222 (O_1222,N_14431,N_14024);
xnor UO_1223 (O_1223,N_14498,N_14560);
nor UO_1224 (O_1224,N_13969,N_14784);
nor UO_1225 (O_1225,N_14334,N_14568);
nand UO_1226 (O_1226,N_14829,N_14833);
or UO_1227 (O_1227,N_14357,N_13867);
or UO_1228 (O_1228,N_14565,N_14193);
nor UO_1229 (O_1229,N_13721,N_14519);
xor UO_1230 (O_1230,N_14367,N_14286);
nand UO_1231 (O_1231,N_13593,N_13540);
nor UO_1232 (O_1232,N_13818,N_14185);
and UO_1233 (O_1233,N_14457,N_13614);
nand UO_1234 (O_1234,N_14811,N_13692);
nand UO_1235 (O_1235,N_14764,N_14041);
nor UO_1236 (O_1236,N_13757,N_13915);
and UO_1237 (O_1237,N_14411,N_14370);
and UO_1238 (O_1238,N_14677,N_14286);
or UO_1239 (O_1239,N_14757,N_14184);
nand UO_1240 (O_1240,N_13606,N_14075);
nand UO_1241 (O_1241,N_14505,N_14014);
nor UO_1242 (O_1242,N_14467,N_13805);
or UO_1243 (O_1243,N_13708,N_14940);
or UO_1244 (O_1244,N_13560,N_13834);
and UO_1245 (O_1245,N_13705,N_14169);
or UO_1246 (O_1246,N_13912,N_13747);
nor UO_1247 (O_1247,N_14377,N_13709);
and UO_1248 (O_1248,N_13744,N_14733);
nor UO_1249 (O_1249,N_14781,N_14423);
and UO_1250 (O_1250,N_13952,N_14582);
nor UO_1251 (O_1251,N_13927,N_13704);
or UO_1252 (O_1252,N_14674,N_13574);
xor UO_1253 (O_1253,N_14570,N_14809);
and UO_1254 (O_1254,N_14001,N_14350);
nand UO_1255 (O_1255,N_14431,N_14530);
nor UO_1256 (O_1256,N_14074,N_13892);
xor UO_1257 (O_1257,N_13706,N_14863);
and UO_1258 (O_1258,N_14058,N_14258);
and UO_1259 (O_1259,N_14721,N_14883);
and UO_1260 (O_1260,N_14421,N_14852);
xnor UO_1261 (O_1261,N_13820,N_14516);
and UO_1262 (O_1262,N_13680,N_14504);
nand UO_1263 (O_1263,N_13509,N_13787);
nor UO_1264 (O_1264,N_14907,N_13887);
and UO_1265 (O_1265,N_13989,N_14700);
nor UO_1266 (O_1266,N_13690,N_13897);
or UO_1267 (O_1267,N_14987,N_14031);
nor UO_1268 (O_1268,N_14329,N_13941);
or UO_1269 (O_1269,N_14506,N_14512);
and UO_1270 (O_1270,N_14909,N_14526);
xnor UO_1271 (O_1271,N_14249,N_14001);
xor UO_1272 (O_1272,N_14967,N_14811);
nand UO_1273 (O_1273,N_13716,N_14972);
and UO_1274 (O_1274,N_14199,N_14502);
nand UO_1275 (O_1275,N_13908,N_13574);
nor UO_1276 (O_1276,N_14425,N_13967);
or UO_1277 (O_1277,N_14989,N_14851);
and UO_1278 (O_1278,N_14982,N_14092);
or UO_1279 (O_1279,N_14458,N_14280);
nand UO_1280 (O_1280,N_13615,N_14174);
nor UO_1281 (O_1281,N_14776,N_14691);
or UO_1282 (O_1282,N_13538,N_14864);
or UO_1283 (O_1283,N_14435,N_13600);
or UO_1284 (O_1284,N_14803,N_14620);
nor UO_1285 (O_1285,N_14526,N_13515);
and UO_1286 (O_1286,N_14063,N_14058);
nand UO_1287 (O_1287,N_13689,N_14557);
nand UO_1288 (O_1288,N_13754,N_14161);
nor UO_1289 (O_1289,N_14722,N_13541);
xnor UO_1290 (O_1290,N_14886,N_14380);
and UO_1291 (O_1291,N_14614,N_14753);
or UO_1292 (O_1292,N_14596,N_14001);
and UO_1293 (O_1293,N_14834,N_13658);
and UO_1294 (O_1294,N_13993,N_13834);
nor UO_1295 (O_1295,N_13730,N_14223);
nor UO_1296 (O_1296,N_13803,N_14042);
nand UO_1297 (O_1297,N_14562,N_14928);
or UO_1298 (O_1298,N_14965,N_14946);
nand UO_1299 (O_1299,N_14706,N_14288);
and UO_1300 (O_1300,N_13873,N_14022);
or UO_1301 (O_1301,N_14661,N_14903);
nand UO_1302 (O_1302,N_13533,N_14152);
nor UO_1303 (O_1303,N_14318,N_14842);
and UO_1304 (O_1304,N_14297,N_14447);
xor UO_1305 (O_1305,N_14522,N_14265);
or UO_1306 (O_1306,N_14909,N_14895);
and UO_1307 (O_1307,N_13513,N_14191);
xor UO_1308 (O_1308,N_13999,N_14351);
or UO_1309 (O_1309,N_14185,N_13672);
or UO_1310 (O_1310,N_13584,N_13657);
and UO_1311 (O_1311,N_13712,N_14561);
or UO_1312 (O_1312,N_14581,N_13520);
xnor UO_1313 (O_1313,N_14171,N_13937);
xor UO_1314 (O_1314,N_14698,N_14254);
or UO_1315 (O_1315,N_14345,N_13610);
and UO_1316 (O_1316,N_14259,N_13761);
xor UO_1317 (O_1317,N_13520,N_14938);
nand UO_1318 (O_1318,N_13815,N_13674);
nor UO_1319 (O_1319,N_13673,N_14814);
nand UO_1320 (O_1320,N_14506,N_14747);
xor UO_1321 (O_1321,N_13660,N_14013);
and UO_1322 (O_1322,N_14546,N_14191);
and UO_1323 (O_1323,N_14477,N_14839);
or UO_1324 (O_1324,N_14545,N_14205);
xor UO_1325 (O_1325,N_13773,N_14471);
or UO_1326 (O_1326,N_14413,N_13922);
or UO_1327 (O_1327,N_14414,N_14761);
or UO_1328 (O_1328,N_13859,N_13866);
nor UO_1329 (O_1329,N_14397,N_14850);
and UO_1330 (O_1330,N_13513,N_13821);
nor UO_1331 (O_1331,N_14699,N_14183);
or UO_1332 (O_1332,N_13875,N_14909);
xnor UO_1333 (O_1333,N_13666,N_14836);
nor UO_1334 (O_1334,N_14396,N_14613);
and UO_1335 (O_1335,N_14394,N_14371);
or UO_1336 (O_1336,N_14752,N_13805);
and UO_1337 (O_1337,N_13562,N_14922);
or UO_1338 (O_1338,N_14842,N_14306);
and UO_1339 (O_1339,N_14981,N_14545);
nor UO_1340 (O_1340,N_14569,N_14146);
nand UO_1341 (O_1341,N_14724,N_14903);
and UO_1342 (O_1342,N_14816,N_13590);
and UO_1343 (O_1343,N_13538,N_14747);
nor UO_1344 (O_1344,N_14665,N_14728);
nand UO_1345 (O_1345,N_13638,N_13595);
and UO_1346 (O_1346,N_13997,N_14936);
or UO_1347 (O_1347,N_14164,N_13742);
nor UO_1348 (O_1348,N_14601,N_14809);
nand UO_1349 (O_1349,N_13677,N_13734);
nor UO_1350 (O_1350,N_14152,N_14894);
nor UO_1351 (O_1351,N_13994,N_14667);
nor UO_1352 (O_1352,N_14012,N_13993);
xnor UO_1353 (O_1353,N_14462,N_14291);
nand UO_1354 (O_1354,N_14332,N_14474);
or UO_1355 (O_1355,N_14285,N_14067);
and UO_1356 (O_1356,N_14262,N_13749);
and UO_1357 (O_1357,N_14977,N_13638);
and UO_1358 (O_1358,N_13789,N_13788);
xnor UO_1359 (O_1359,N_14309,N_14871);
and UO_1360 (O_1360,N_13623,N_14515);
nand UO_1361 (O_1361,N_13628,N_13757);
nor UO_1362 (O_1362,N_13661,N_14150);
nand UO_1363 (O_1363,N_14699,N_14444);
and UO_1364 (O_1364,N_13763,N_14955);
nor UO_1365 (O_1365,N_13874,N_13958);
nand UO_1366 (O_1366,N_14448,N_14141);
and UO_1367 (O_1367,N_13801,N_13566);
or UO_1368 (O_1368,N_14562,N_13606);
xor UO_1369 (O_1369,N_13930,N_13824);
nand UO_1370 (O_1370,N_13960,N_14803);
nand UO_1371 (O_1371,N_14938,N_13573);
nor UO_1372 (O_1372,N_13902,N_14050);
nand UO_1373 (O_1373,N_13946,N_14275);
or UO_1374 (O_1374,N_14415,N_14607);
nor UO_1375 (O_1375,N_13971,N_14280);
nand UO_1376 (O_1376,N_14814,N_14256);
or UO_1377 (O_1377,N_13879,N_14019);
nand UO_1378 (O_1378,N_14544,N_14623);
nor UO_1379 (O_1379,N_14992,N_13944);
or UO_1380 (O_1380,N_14580,N_14173);
and UO_1381 (O_1381,N_13967,N_14879);
nor UO_1382 (O_1382,N_14679,N_14249);
or UO_1383 (O_1383,N_13550,N_14080);
or UO_1384 (O_1384,N_13893,N_14129);
and UO_1385 (O_1385,N_13632,N_13688);
xor UO_1386 (O_1386,N_13583,N_14747);
or UO_1387 (O_1387,N_13554,N_13509);
or UO_1388 (O_1388,N_14066,N_14812);
or UO_1389 (O_1389,N_13621,N_14705);
nand UO_1390 (O_1390,N_14405,N_14148);
and UO_1391 (O_1391,N_13835,N_14745);
nand UO_1392 (O_1392,N_14668,N_14287);
or UO_1393 (O_1393,N_13645,N_13633);
xnor UO_1394 (O_1394,N_13869,N_13611);
xnor UO_1395 (O_1395,N_13947,N_14714);
nand UO_1396 (O_1396,N_13548,N_14477);
nand UO_1397 (O_1397,N_14199,N_13947);
nor UO_1398 (O_1398,N_14059,N_14724);
nand UO_1399 (O_1399,N_14353,N_14182);
nand UO_1400 (O_1400,N_14289,N_14782);
nor UO_1401 (O_1401,N_14352,N_13929);
nor UO_1402 (O_1402,N_14558,N_14840);
nor UO_1403 (O_1403,N_14043,N_13909);
nand UO_1404 (O_1404,N_13562,N_14692);
nor UO_1405 (O_1405,N_14440,N_14527);
and UO_1406 (O_1406,N_14035,N_14954);
nand UO_1407 (O_1407,N_14250,N_14690);
or UO_1408 (O_1408,N_14700,N_14227);
nand UO_1409 (O_1409,N_13512,N_14619);
nor UO_1410 (O_1410,N_14570,N_14094);
nor UO_1411 (O_1411,N_14803,N_13952);
or UO_1412 (O_1412,N_14424,N_13730);
xor UO_1413 (O_1413,N_14439,N_14614);
nand UO_1414 (O_1414,N_14096,N_14053);
nand UO_1415 (O_1415,N_13644,N_13950);
nor UO_1416 (O_1416,N_14989,N_14306);
nor UO_1417 (O_1417,N_14090,N_13933);
xnor UO_1418 (O_1418,N_14709,N_14330);
nor UO_1419 (O_1419,N_13926,N_14926);
or UO_1420 (O_1420,N_14997,N_14269);
xnor UO_1421 (O_1421,N_13731,N_13696);
nor UO_1422 (O_1422,N_14613,N_13625);
nor UO_1423 (O_1423,N_13980,N_14167);
nand UO_1424 (O_1424,N_14165,N_14556);
nor UO_1425 (O_1425,N_13781,N_14594);
nor UO_1426 (O_1426,N_14460,N_14170);
nor UO_1427 (O_1427,N_13813,N_14504);
or UO_1428 (O_1428,N_14031,N_13988);
and UO_1429 (O_1429,N_13941,N_13748);
xnor UO_1430 (O_1430,N_13808,N_14987);
nor UO_1431 (O_1431,N_13632,N_14605);
nor UO_1432 (O_1432,N_13549,N_13502);
nor UO_1433 (O_1433,N_14815,N_14404);
and UO_1434 (O_1434,N_13710,N_14920);
nor UO_1435 (O_1435,N_14950,N_13777);
or UO_1436 (O_1436,N_14438,N_14519);
nor UO_1437 (O_1437,N_14026,N_14456);
nand UO_1438 (O_1438,N_13742,N_14969);
nand UO_1439 (O_1439,N_14263,N_14699);
xnor UO_1440 (O_1440,N_14370,N_14621);
xnor UO_1441 (O_1441,N_14539,N_14204);
nor UO_1442 (O_1442,N_13555,N_14425);
nor UO_1443 (O_1443,N_14431,N_14638);
or UO_1444 (O_1444,N_14049,N_14157);
nand UO_1445 (O_1445,N_14996,N_14744);
nand UO_1446 (O_1446,N_14165,N_14695);
or UO_1447 (O_1447,N_13944,N_13990);
nand UO_1448 (O_1448,N_14498,N_13917);
nor UO_1449 (O_1449,N_13850,N_13755);
xnor UO_1450 (O_1450,N_14270,N_14909);
nor UO_1451 (O_1451,N_13514,N_14971);
nor UO_1452 (O_1452,N_13903,N_14265);
or UO_1453 (O_1453,N_14520,N_14870);
or UO_1454 (O_1454,N_14795,N_14332);
nor UO_1455 (O_1455,N_13919,N_13849);
or UO_1456 (O_1456,N_14687,N_14272);
nand UO_1457 (O_1457,N_13581,N_14547);
nand UO_1458 (O_1458,N_14455,N_13956);
nand UO_1459 (O_1459,N_14745,N_14076);
xnor UO_1460 (O_1460,N_14753,N_14263);
or UO_1461 (O_1461,N_14776,N_14035);
and UO_1462 (O_1462,N_14436,N_13736);
and UO_1463 (O_1463,N_14220,N_14087);
nand UO_1464 (O_1464,N_13554,N_13533);
and UO_1465 (O_1465,N_14340,N_14164);
or UO_1466 (O_1466,N_14489,N_14529);
nor UO_1467 (O_1467,N_13639,N_14157);
nand UO_1468 (O_1468,N_14315,N_14694);
nor UO_1469 (O_1469,N_14302,N_13509);
nor UO_1470 (O_1470,N_14668,N_14537);
or UO_1471 (O_1471,N_14062,N_14825);
xnor UO_1472 (O_1472,N_14187,N_13828);
nor UO_1473 (O_1473,N_13987,N_14462);
nand UO_1474 (O_1474,N_14410,N_13810);
nor UO_1475 (O_1475,N_14237,N_14029);
nand UO_1476 (O_1476,N_14943,N_14345);
nor UO_1477 (O_1477,N_13851,N_14064);
and UO_1478 (O_1478,N_13961,N_14076);
and UO_1479 (O_1479,N_14637,N_14316);
or UO_1480 (O_1480,N_14182,N_14617);
and UO_1481 (O_1481,N_14052,N_14887);
xor UO_1482 (O_1482,N_14295,N_14496);
or UO_1483 (O_1483,N_14278,N_14021);
nor UO_1484 (O_1484,N_14974,N_14729);
and UO_1485 (O_1485,N_14027,N_13882);
nand UO_1486 (O_1486,N_13625,N_13700);
and UO_1487 (O_1487,N_13595,N_14154);
nand UO_1488 (O_1488,N_13913,N_13557);
and UO_1489 (O_1489,N_14776,N_13658);
or UO_1490 (O_1490,N_14503,N_14904);
and UO_1491 (O_1491,N_14336,N_14049);
nand UO_1492 (O_1492,N_13686,N_14559);
xor UO_1493 (O_1493,N_13573,N_14496);
and UO_1494 (O_1494,N_14741,N_13895);
and UO_1495 (O_1495,N_13999,N_14454);
and UO_1496 (O_1496,N_14090,N_13628);
and UO_1497 (O_1497,N_14044,N_14775);
nor UO_1498 (O_1498,N_14659,N_14700);
and UO_1499 (O_1499,N_14727,N_14754);
nand UO_1500 (O_1500,N_14568,N_14388);
or UO_1501 (O_1501,N_13710,N_14799);
nor UO_1502 (O_1502,N_13889,N_14458);
nor UO_1503 (O_1503,N_14468,N_14196);
nand UO_1504 (O_1504,N_14034,N_14658);
or UO_1505 (O_1505,N_14417,N_14444);
nor UO_1506 (O_1506,N_14502,N_14774);
and UO_1507 (O_1507,N_13531,N_14340);
nand UO_1508 (O_1508,N_14367,N_14881);
nor UO_1509 (O_1509,N_14031,N_14559);
nand UO_1510 (O_1510,N_13967,N_14680);
or UO_1511 (O_1511,N_14721,N_13534);
nand UO_1512 (O_1512,N_14520,N_13957);
or UO_1513 (O_1513,N_14829,N_13732);
or UO_1514 (O_1514,N_14485,N_14952);
or UO_1515 (O_1515,N_14046,N_13820);
and UO_1516 (O_1516,N_14437,N_14052);
and UO_1517 (O_1517,N_14708,N_14868);
nor UO_1518 (O_1518,N_14155,N_14813);
nand UO_1519 (O_1519,N_13962,N_13827);
nand UO_1520 (O_1520,N_13505,N_14838);
nor UO_1521 (O_1521,N_13780,N_13687);
and UO_1522 (O_1522,N_14680,N_14196);
nand UO_1523 (O_1523,N_14501,N_13839);
or UO_1524 (O_1524,N_14740,N_14002);
and UO_1525 (O_1525,N_13921,N_14711);
nand UO_1526 (O_1526,N_14239,N_14117);
or UO_1527 (O_1527,N_14790,N_13772);
nor UO_1528 (O_1528,N_13603,N_14119);
and UO_1529 (O_1529,N_14981,N_13555);
nand UO_1530 (O_1530,N_14074,N_13794);
nand UO_1531 (O_1531,N_13925,N_13802);
or UO_1532 (O_1532,N_13782,N_14383);
or UO_1533 (O_1533,N_14456,N_14773);
and UO_1534 (O_1534,N_14291,N_13768);
nor UO_1535 (O_1535,N_13664,N_14613);
or UO_1536 (O_1536,N_14464,N_13920);
nand UO_1537 (O_1537,N_14483,N_14006);
or UO_1538 (O_1538,N_14208,N_14309);
or UO_1539 (O_1539,N_14625,N_14052);
nand UO_1540 (O_1540,N_14531,N_14293);
or UO_1541 (O_1541,N_14629,N_14435);
or UO_1542 (O_1542,N_14992,N_13876);
nor UO_1543 (O_1543,N_13807,N_14513);
and UO_1544 (O_1544,N_14893,N_14142);
or UO_1545 (O_1545,N_14315,N_13613);
and UO_1546 (O_1546,N_14151,N_14400);
and UO_1547 (O_1547,N_14652,N_13882);
nor UO_1548 (O_1548,N_13993,N_14730);
nand UO_1549 (O_1549,N_14226,N_14259);
nand UO_1550 (O_1550,N_13952,N_14163);
and UO_1551 (O_1551,N_14382,N_13580);
or UO_1552 (O_1552,N_14557,N_13627);
or UO_1553 (O_1553,N_14470,N_14241);
nand UO_1554 (O_1554,N_13520,N_13584);
nand UO_1555 (O_1555,N_13746,N_14768);
and UO_1556 (O_1556,N_14907,N_14856);
xnor UO_1557 (O_1557,N_13681,N_13675);
or UO_1558 (O_1558,N_14625,N_14554);
and UO_1559 (O_1559,N_14711,N_14673);
or UO_1560 (O_1560,N_14326,N_13773);
xnor UO_1561 (O_1561,N_13570,N_13916);
nand UO_1562 (O_1562,N_13658,N_14078);
and UO_1563 (O_1563,N_13678,N_13937);
nor UO_1564 (O_1564,N_14040,N_14330);
nor UO_1565 (O_1565,N_14753,N_14081);
nand UO_1566 (O_1566,N_14489,N_13570);
or UO_1567 (O_1567,N_13911,N_14980);
and UO_1568 (O_1568,N_14909,N_13812);
nand UO_1569 (O_1569,N_13574,N_14226);
and UO_1570 (O_1570,N_14946,N_14237);
nor UO_1571 (O_1571,N_14439,N_13872);
and UO_1572 (O_1572,N_14782,N_13960);
or UO_1573 (O_1573,N_14618,N_14342);
nand UO_1574 (O_1574,N_13955,N_14981);
xnor UO_1575 (O_1575,N_14707,N_14622);
nor UO_1576 (O_1576,N_14847,N_13735);
or UO_1577 (O_1577,N_14493,N_14884);
or UO_1578 (O_1578,N_13596,N_14742);
nand UO_1579 (O_1579,N_14135,N_13505);
and UO_1580 (O_1580,N_14571,N_13557);
nand UO_1581 (O_1581,N_14183,N_13639);
or UO_1582 (O_1582,N_13580,N_13586);
xor UO_1583 (O_1583,N_14407,N_14334);
and UO_1584 (O_1584,N_13678,N_13622);
and UO_1585 (O_1585,N_13768,N_14826);
nand UO_1586 (O_1586,N_14623,N_13734);
nor UO_1587 (O_1587,N_14471,N_13567);
xnor UO_1588 (O_1588,N_14339,N_14540);
nor UO_1589 (O_1589,N_13592,N_13596);
and UO_1590 (O_1590,N_14139,N_13873);
nand UO_1591 (O_1591,N_14881,N_13724);
xor UO_1592 (O_1592,N_14263,N_13791);
or UO_1593 (O_1593,N_13961,N_14886);
or UO_1594 (O_1594,N_13784,N_13849);
and UO_1595 (O_1595,N_14175,N_13542);
and UO_1596 (O_1596,N_14370,N_13791);
or UO_1597 (O_1597,N_14221,N_14172);
nor UO_1598 (O_1598,N_14528,N_13784);
or UO_1599 (O_1599,N_14283,N_13989);
nor UO_1600 (O_1600,N_14124,N_13901);
and UO_1601 (O_1601,N_14537,N_14625);
or UO_1602 (O_1602,N_14186,N_14321);
nor UO_1603 (O_1603,N_14547,N_14981);
nor UO_1604 (O_1604,N_13581,N_13896);
and UO_1605 (O_1605,N_13783,N_14587);
or UO_1606 (O_1606,N_14328,N_13802);
nor UO_1607 (O_1607,N_14376,N_14127);
nand UO_1608 (O_1608,N_14108,N_14002);
or UO_1609 (O_1609,N_13958,N_13847);
nand UO_1610 (O_1610,N_14174,N_14929);
nor UO_1611 (O_1611,N_14840,N_13780);
and UO_1612 (O_1612,N_14549,N_14898);
or UO_1613 (O_1613,N_13763,N_14356);
nor UO_1614 (O_1614,N_14147,N_14460);
nand UO_1615 (O_1615,N_14939,N_14365);
nor UO_1616 (O_1616,N_13613,N_14657);
nor UO_1617 (O_1617,N_13524,N_14101);
and UO_1618 (O_1618,N_14782,N_14202);
or UO_1619 (O_1619,N_13937,N_13765);
nor UO_1620 (O_1620,N_14419,N_13596);
or UO_1621 (O_1621,N_14501,N_14497);
or UO_1622 (O_1622,N_14720,N_14847);
and UO_1623 (O_1623,N_13582,N_13806);
nor UO_1624 (O_1624,N_13631,N_14316);
nand UO_1625 (O_1625,N_13501,N_14360);
nand UO_1626 (O_1626,N_13812,N_13767);
or UO_1627 (O_1627,N_14554,N_14735);
or UO_1628 (O_1628,N_13582,N_14393);
xnor UO_1629 (O_1629,N_13830,N_14094);
nor UO_1630 (O_1630,N_13705,N_13602);
and UO_1631 (O_1631,N_14974,N_14829);
or UO_1632 (O_1632,N_14202,N_13809);
and UO_1633 (O_1633,N_13747,N_13698);
or UO_1634 (O_1634,N_13515,N_13890);
and UO_1635 (O_1635,N_14515,N_14676);
nand UO_1636 (O_1636,N_14334,N_13872);
or UO_1637 (O_1637,N_14585,N_13624);
or UO_1638 (O_1638,N_14972,N_13934);
xor UO_1639 (O_1639,N_14970,N_14851);
and UO_1640 (O_1640,N_13830,N_13722);
nor UO_1641 (O_1641,N_13528,N_14259);
and UO_1642 (O_1642,N_14583,N_14782);
xor UO_1643 (O_1643,N_14255,N_13678);
xnor UO_1644 (O_1644,N_14472,N_13981);
nor UO_1645 (O_1645,N_14488,N_14589);
nand UO_1646 (O_1646,N_14524,N_14345);
nor UO_1647 (O_1647,N_13704,N_14778);
and UO_1648 (O_1648,N_13829,N_14351);
nand UO_1649 (O_1649,N_14174,N_14515);
nor UO_1650 (O_1650,N_14507,N_14011);
or UO_1651 (O_1651,N_14501,N_14797);
nor UO_1652 (O_1652,N_14221,N_14512);
nand UO_1653 (O_1653,N_14687,N_13675);
and UO_1654 (O_1654,N_14528,N_14955);
xnor UO_1655 (O_1655,N_13518,N_13554);
nand UO_1656 (O_1656,N_14823,N_14695);
or UO_1657 (O_1657,N_14449,N_14248);
and UO_1658 (O_1658,N_14630,N_14890);
nor UO_1659 (O_1659,N_13746,N_14983);
nor UO_1660 (O_1660,N_14637,N_14498);
nor UO_1661 (O_1661,N_14988,N_13931);
or UO_1662 (O_1662,N_14998,N_14854);
or UO_1663 (O_1663,N_14358,N_14567);
nand UO_1664 (O_1664,N_14787,N_13968);
nor UO_1665 (O_1665,N_13572,N_14455);
and UO_1666 (O_1666,N_14182,N_14649);
and UO_1667 (O_1667,N_14632,N_14916);
nor UO_1668 (O_1668,N_14194,N_14373);
and UO_1669 (O_1669,N_13949,N_13591);
nand UO_1670 (O_1670,N_13666,N_14820);
nor UO_1671 (O_1671,N_14924,N_14388);
or UO_1672 (O_1672,N_14806,N_14426);
nor UO_1673 (O_1673,N_14980,N_13788);
and UO_1674 (O_1674,N_13824,N_13803);
and UO_1675 (O_1675,N_14195,N_13831);
or UO_1676 (O_1676,N_13865,N_13606);
and UO_1677 (O_1677,N_14961,N_14020);
nor UO_1678 (O_1678,N_14881,N_14423);
nor UO_1679 (O_1679,N_13758,N_13524);
nor UO_1680 (O_1680,N_13891,N_14838);
nor UO_1681 (O_1681,N_13929,N_13976);
or UO_1682 (O_1682,N_14905,N_14588);
nor UO_1683 (O_1683,N_13971,N_13792);
or UO_1684 (O_1684,N_14159,N_14689);
nand UO_1685 (O_1685,N_14039,N_14121);
nor UO_1686 (O_1686,N_13743,N_14299);
nor UO_1687 (O_1687,N_13688,N_14652);
or UO_1688 (O_1688,N_14922,N_14505);
nand UO_1689 (O_1689,N_14245,N_13911);
or UO_1690 (O_1690,N_13950,N_13584);
xor UO_1691 (O_1691,N_14924,N_14483);
nand UO_1692 (O_1692,N_14040,N_14129);
and UO_1693 (O_1693,N_13859,N_13799);
or UO_1694 (O_1694,N_14115,N_14188);
xnor UO_1695 (O_1695,N_14766,N_13891);
nor UO_1696 (O_1696,N_14906,N_13632);
or UO_1697 (O_1697,N_13577,N_13518);
and UO_1698 (O_1698,N_13737,N_13734);
and UO_1699 (O_1699,N_14099,N_13965);
and UO_1700 (O_1700,N_14002,N_14912);
nand UO_1701 (O_1701,N_14968,N_13601);
xnor UO_1702 (O_1702,N_13527,N_14759);
and UO_1703 (O_1703,N_14332,N_14255);
nand UO_1704 (O_1704,N_14114,N_14264);
nor UO_1705 (O_1705,N_14188,N_14433);
nor UO_1706 (O_1706,N_13535,N_14308);
xnor UO_1707 (O_1707,N_14003,N_14292);
or UO_1708 (O_1708,N_13636,N_14752);
nor UO_1709 (O_1709,N_14308,N_14934);
and UO_1710 (O_1710,N_14771,N_14457);
and UO_1711 (O_1711,N_14713,N_14177);
or UO_1712 (O_1712,N_14244,N_14718);
and UO_1713 (O_1713,N_13738,N_13575);
and UO_1714 (O_1714,N_14185,N_13811);
nand UO_1715 (O_1715,N_13939,N_14537);
xor UO_1716 (O_1716,N_14579,N_13817);
nand UO_1717 (O_1717,N_14453,N_13963);
and UO_1718 (O_1718,N_14738,N_13634);
nand UO_1719 (O_1719,N_14788,N_14389);
or UO_1720 (O_1720,N_14550,N_13967);
nor UO_1721 (O_1721,N_14092,N_14968);
nor UO_1722 (O_1722,N_14493,N_13507);
or UO_1723 (O_1723,N_13849,N_14035);
or UO_1724 (O_1724,N_14251,N_13506);
and UO_1725 (O_1725,N_13838,N_14032);
nand UO_1726 (O_1726,N_14134,N_13675);
nor UO_1727 (O_1727,N_14184,N_14952);
or UO_1728 (O_1728,N_13682,N_13764);
nor UO_1729 (O_1729,N_14175,N_13726);
and UO_1730 (O_1730,N_14750,N_13820);
xor UO_1731 (O_1731,N_13573,N_13627);
or UO_1732 (O_1732,N_14246,N_14442);
and UO_1733 (O_1733,N_13714,N_14574);
or UO_1734 (O_1734,N_14600,N_14543);
and UO_1735 (O_1735,N_13605,N_14151);
or UO_1736 (O_1736,N_14272,N_14208);
or UO_1737 (O_1737,N_14200,N_14145);
or UO_1738 (O_1738,N_14750,N_14459);
or UO_1739 (O_1739,N_14521,N_13794);
xnor UO_1740 (O_1740,N_14519,N_14026);
or UO_1741 (O_1741,N_14432,N_13858);
nand UO_1742 (O_1742,N_13747,N_13610);
nor UO_1743 (O_1743,N_14820,N_14786);
xnor UO_1744 (O_1744,N_14692,N_14519);
or UO_1745 (O_1745,N_14196,N_13612);
xor UO_1746 (O_1746,N_13629,N_14243);
and UO_1747 (O_1747,N_14446,N_13838);
and UO_1748 (O_1748,N_14244,N_14516);
and UO_1749 (O_1749,N_13642,N_14020);
xor UO_1750 (O_1750,N_14979,N_13836);
xor UO_1751 (O_1751,N_13869,N_14890);
nor UO_1752 (O_1752,N_14544,N_13954);
nand UO_1753 (O_1753,N_14266,N_13808);
and UO_1754 (O_1754,N_14369,N_13603);
nor UO_1755 (O_1755,N_13645,N_13635);
or UO_1756 (O_1756,N_13815,N_14983);
nor UO_1757 (O_1757,N_14663,N_14559);
and UO_1758 (O_1758,N_13827,N_14166);
or UO_1759 (O_1759,N_14487,N_13889);
xnor UO_1760 (O_1760,N_14153,N_14633);
nor UO_1761 (O_1761,N_14380,N_14074);
nor UO_1762 (O_1762,N_13632,N_14941);
or UO_1763 (O_1763,N_13804,N_14515);
or UO_1764 (O_1764,N_14848,N_13571);
and UO_1765 (O_1765,N_14832,N_13500);
or UO_1766 (O_1766,N_14284,N_14276);
or UO_1767 (O_1767,N_14397,N_14087);
and UO_1768 (O_1768,N_14341,N_14365);
nor UO_1769 (O_1769,N_14509,N_13922);
or UO_1770 (O_1770,N_14542,N_14062);
or UO_1771 (O_1771,N_14236,N_14212);
nand UO_1772 (O_1772,N_14794,N_13547);
nand UO_1773 (O_1773,N_13866,N_13691);
nand UO_1774 (O_1774,N_13909,N_14265);
or UO_1775 (O_1775,N_13764,N_14350);
nand UO_1776 (O_1776,N_14477,N_14488);
or UO_1777 (O_1777,N_14069,N_14635);
nor UO_1778 (O_1778,N_14925,N_14237);
nand UO_1779 (O_1779,N_13858,N_14282);
and UO_1780 (O_1780,N_14627,N_13608);
nor UO_1781 (O_1781,N_14171,N_14442);
xnor UO_1782 (O_1782,N_13960,N_14092);
nor UO_1783 (O_1783,N_14885,N_14607);
nor UO_1784 (O_1784,N_14203,N_14426);
nand UO_1785 (O_1785,N_14686,N_13997);
xor UO_1786 (O_1786,N_14862,N_14905);
nor UO_1787 (O_1787,N_14378,N_14962);
and UO_1788 (O_1788,N_13810,N_14165);
nand UO_1789 (O_1789,N_14903,N_14488);
and UO_1790 (O_1790,N_13781,N_13977);
or UO_1791 (O_1791,N_14014,N_14651);
xnor UO_1792 (O_1792,N_13856,N_14710);
xnor UO_1793 (O_1793,N_14955,N_14490);
nand UO_1794 (O_1794,N_14508,N_13830);
nor UO_1795 (O_1795,N_13848,N_14722);
and UO_1796 (O_1796,N_13607,N_14074);
nor UO_1797 (O_1797,N_14048,N_13833);
xnor UO_1798 (O_1798,N_13791,N_14871);
nand UO_1799 (O_1799,N_14051,N_13587);
nor UO_1800 (O_1800,N_14134,N_14831);
nand UO_1801 (O_1801,N_14470,N_13739);
and UO_1802 (O_1802,N_14231,N_13644);
nor UO_1803 (O_1803,N_14111,N_14636);
and UO_1804 (O_1804,N_14173,N_13545);
nor UO_1805 (O_1805,N_13557,N_14935);
or UO_1806 (O_1806,N_13917,N_14675);
nand UO_1807 (O_1807,N_14414,N_14043);
nand UO_1808 (O_1808,N_13876,N_14339);
nand UO_1809 (O_1809,N_14724,N_13662);
nor UO_1810 (O_1810,N_13988,N_13860);
xor UO_1811 (O_1811,N_14877,N_13850);
and UO_1812 (O_1812,N_13521,N_14980);
or UO_1813 (O_1813,N_14244,N_14440);
nand UO_1814 (O_1814,N_14741,N_13927);
nor UO_1815 (O_1815,N_14422,N_13972);
nor UO_1816 (O_1816,N_14377,N_13900);
or UO_1817 (O_1817,N_13623,N_14352);
nor UO_1818 (O_1818,N_13921,N_13648);
or UO_1819 (O_1819,N_14094,N_14585);
nor UO_1820 (O_1820,N_14257,N_14082);
nand UO_1821 (O_1821,N_13794,N_13591);
nor UO_1822 (O_1822,N_14456,N_14230);
nand UO_1823 (O_1823,N_14807,N_14876);
and UO_1824 (O_1824,N_14480,N_14547);
nand UO_1825 (O_1825,N_13950,N_13685);
nand UO_1826 (O_1826,N_13825,N_14539);
and UO_1827 (O_1827,N_14302,N_14905);
or UO_1828 (O_1828,N_13640,N_14970);
nor UO_1829 (O_1829,N_14913,N_13801);
and UO_1830 (O_1830,N_14417,N_14581);
and UO_1831 (O_1831,N_14336,N_13588);
or UO_1832 (O_1832,N_14983,N_14758);
or UO_1833 (O_1833,N_14984,N_13736);
and UO_1834 (O_1834,N_14610,N_13819);
nor UO_1835 (O_1835,N_13606,N_14545);
and UO_1836 (O_1836,N_13593,N_14744);
or UO_1837 (O_1837,N_14007,N_13510);
and UO_1838 (O_1838,N_14940,N_14286);
or UO_1839 (O_1839,N_14305,N_14526);
nand UO_1840 (O_1840,N_14816,N_14394);
nor UO_1841 (O_1841,N_14861,N_14537);
and UO_1842 (O_1842,N_13633,N_14291);
nor UO_1843 (O_1843,N_14814,N_13761);
nand UO_1844 (O_1844,N_14545,N_13644);
nor UO_1845 (O_1845,N_14452,N_14292);
xnor UO_1846 (O_1846,N_13784,N_13789);
or UO_1847 (O_1847,N_13602,N_14631);
nor UO_1848 (O_1848,N_14333,N_14227);
or UO_1849 (O_1849,N_14736,N_14894);
and UO_1850 (O_1850,N_14349,N_14621);
nand UO_1851 (O_1851,N_14135,N_14490);
or UO_1852 (O_1852,N_14091,N_14504);
and UO_1853 (O_1853,N_14608,N_14835);
and UO_1854 (O_1854,N_13506,N_13763);
nor UO_1855 (O_1855,N_13854,N_14163);
and UO_1856 (O_1856,N_13671,N_13789);
nor UO_1857 (O_1857,N_13704,N_14036);
nand UO_1858 (O_1858,N_14686,N_13954);
xor UO_1859 (O_1859,N_14907,N_13500);
and UO_1860 (O_1860,N_13818,N_14534);
nand UO_1861 (O_1861,N_13529,N_14382);
xnor UO_1862 (O_1862,N_14368,N_13630);
nor UO_1863 (O_1863,N_13636,N_14686);
nand UO_1864 (O_1864,N_14272,N_14713);
nor UO_1865 (O_1865,N_13572,N_14695);
and UO_1866 (O_1866,N_14323,N_14553);
or UO_1867 (O_1867,N_14704,N_14488);
or UO_1868 (O_1868,N_14913,N_14380);
xor UO_1869 (O_1869,N_14982,N_14960);
nor UO_1870 (O_1870,N_14625,N_13580);
nand UO_1871 (O_1871,N_14241,N_13605);
or UO_1872 (O_1872,N_14081,N_14641);
nor UO_1873 (O_1873,N_13665,N_14918);
or UO_1874 (O_1874,N_13842,N_13799);
nor UO_1875 (O_1875,N_14536,N_14319);
and UO_1876 (O_1876,N_13834,N_13593);
nor UO_1877 (O_1877,N_14631,N_14681);
nand UO_1878 (O_1878,N_14063,N_14230);
and UO_1879 (O_1879,N_14880,N_13811);
xor UO_1880 (O_1880,N_14966,N_14538);
and UO_1881 (O_1881,N_14856,N_13580);
and UO_1882 (O_1882,N_14735,N_14692);
nor UO_1883 (O_1883,N_14497,N_13777);
and UO_1884 (O_1884,N_14091,N_14098);
and UO_1885 (O_1885,N_13936,N_13861);
nand UO_1886 (O_1886,N_14818,N_14881);
nand UO_1887 (O_1887,N_14415,N_13570);
xor UO_1888 (O_1888,N_14204,N_14287);
nand UO_1889 (O_1889,N_14367,N_14032);
nand UO_1890 (O_1890,N_14353,N_13507);
nand UO_1891 (O_1891,N_13522,N_14008);
or UO_1892 (O_1892,N_14706,N_14709);
nor UO_1893 (O_1893,N_14098,N_14956);
xnor UO_1894 (O_1894,N_14002,N_14336);
nand UO_1895 (O_1895,N_14031,N_14609);
nand UO_1896 (O_1896,N_14710,N_14761);
nor UO_1897 (O_1897,N_14376,N_14733);
nand UO_1898 (O_1898,N_13682,N_13727);
and UO_1899 (O_1899,N_14979,N_13586);
nor UO_1900 (O_1900,N_14861,N_13857);
and UO_1901 (O_1901,N_14899,N_14080);
and UO_1902 (O_1902,N_14619,N_14053);
or UO_1903 (O_1903,N_14151,N_14687);
nand UO_1904 (O_1904,N_14637,N_14755);
nor UO_1905 (O_1905,N_14922,N_14767);
xnor UO_1906 (O_1906,N_13840,N_14117);
nand UO_1907 (O_1907,N_13813,N_14089);
or UO_1908 (O_1908,N_13543,N_14684);
nor UO_1909 (O_1909,N_13841,N_14260);
xor UO_1910 (O_1910,N_13750,N_14440);
or UO_1911 (O_1911,N_14648,N_14502);
and UO_1912 (O_1912,N_13881,N_14711);
nand UO_1913 (O_1913,N_13573,N_13906);
or UO_1914 (O_1914,N_14506,N_14248);
or UO_1915 (O_1915,N_14037,N_13929);
nor UO_1916 (O_1916,N_14184,N_14149);
nand UO_1917 (O_1917,N_14170,N_13990);
or UO_1918 (O_1918,N_14348,N_14212);
and UO_1919 (O_1919,N_14313,N_14474);
nor UO_1920 (O_1920,N_13669,N_14392);
and UO_1921 (O_1921,N_13524,N_13698);
nand UO_1922 (O_1922,N_14775,N_13680);
nor UO_1923 (O_1923,N_14397,N_13683);
and UO_1924 (O_1924,N_14349,N_13931);
nand UO_1925 (O_1925,N_13939,N_14847);
or UO_1926 (O_1926,N_13816,N_13873);
and UO_1927 (O_1927,N_14925,N_13946);
or UO_1928 (O_1928,N_13971,N_13998);
and UO_1929 (O_1929,N_14060,N_14500);
and UO_1930 (O_1930,N_13533,N_14687);
nand UO_1931 (O_1931,N_14093,N_13803);
or UO_1932 (O_1932,N_14553,N_14646);
xor UO_1933 (O_1933,N_14425,N_14072);
nor UO_1934 (O_1934,N_14552,N_14768);
or UO_1935 (O_1935,N_14037,N_13638);
and UO_1936 (O_1936,N_14438,N_14374);
or UO_1937 (O_1937,N_13897,N_13864);
or UO_1938 (O_1938,N_14688,N_14996);
and UO_1939 (O_1939,N_13652,N_13519);
nor UO_1940 (O_1940,N_13760,N_14056);
or UO_1941 (O_1941,N_13963,N_13537);
and UO_1942 (O_1942,N_13598,N_14119);
nand UO_1943 (O_1943,N_13507,N_14345);
xor UO_1944 (O_1944,N_13713,N_13677);
and UO_1945 (O_1945,N_14303,N_14326);
or UO_1946 (O_1946,N_14652,N_13998);
and UO_1947 (O_1947,N_13984,N_14713);
nand UO_1948 (O_1948,N_14951,N_14133);
and UO_1949 (O_1949,N_14419,N_13665);
nor UO_1950 (O_1950,N_14184,N_14648);
nor UO_1951 (O_1951,N_14484,N_14956);
nor UO_1952 (O_1952,N_14756,N_14918);
nor UO_1953 (O_1953,N_14723,N_13815);
xor UO_1954 (O_1954,N_14506,N_13841);
nor UO_1955 (O_1955,N_14988,N_13941);
nor UO_1956 (O_1956,N_14613,N_14778);
and UO_1957 (O_1957,N_13795,N_13624);
or UO_1958 (O_1958,N_14293,N_13564);
nand UO_1959 (O_1959,N_13902,N_14806);
nor UO_1960 (O_1960,N_14191,N_14673);
nand UO_1961 (O_1961,N_13628,N_14541);
nor UO_1962 (O_1962,N_13868,N_14684);
or UO_1963 (O_1963,N_14926,N_14209);
or UO_1964 (O_1964,N_14922,N_14724);
and UO_1965 (O_1965,N_13970,N_14788);
nor UO_1966 (O_1966,N_14170,N_14779);
or UO_1967 (O_1967,N_14296,N_14059);
and UO_1968 (O_1968,N_14694,N_14715);
nor UO_1969 (O_1969,N_13736,N_13751);
and UO_1970 (O_1970,N_14230,N_14752);
nand UO_1971 (O_1971,N_14297,N_14032);
or UO_1972 (O_1972,N_14660,N_14023);
xnor UO_1973 (O_1973,N_14714,N_14104);
or UO_1974 (O_1974,N_14794,N_14031);
nand UO_1975 (O_1975,N_14292,N_14744);
nor UO_1976 (O_1976,N_14230,N_14729);
nand UO_1977 (O_1977,N_13891,N_14651);
nor UO_1978 (O_1978,N_13551,N_14321);
nand UO_1979 (O_1979,N_14130,N_14910);
xnor UO_1980 (O_1980,N_13671,N_14162);
xor UO_1981 (O_1981,N_14092,N_13779);
or UO_1982 (O_1982,N_13778,N_13894);
and UO_1983 (O_1983,N_13547,N_13604);
and UO_1984 (O_1984,N_14718,N_14997);
nor UO_1985 (O_1985,N_14388,N_13543);
nor UO_1986 (O_1986,N_13922,N_13997);
or UO_1987 (O_1987,N_14687,N_14363);
and UO_1988 (O_1988,N_14522,N_14536);
xnor UO_1989 (O_1989,N_14391,N_14156);
or UO_1990 (O_1990,N_14208,N_14118);
and UO_1991 (O_1991,N_14682,N_14495);
nand UO_1992 (O_1992,N_13921,N_14950);
or UO_1993 (O_1993,N_14973,N_14983);
nor UO_1994 (O_1994,N_14323,N_14688);
nor UO_1995 (O_1995,N_13750,N_13735);
nor UO_1996 (O_1996,N_13632,N_14445);
or UO_1997 (O_1997,N_14353,N_13748);
nor UO_1998 (O_1998,N_14278,N_14605);
xnor UO_1999 (O_1999,N_13577,N_14895);
endmodule