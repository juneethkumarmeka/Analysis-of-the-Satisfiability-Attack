module basic_500_3000_500_30_levels_1xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
xnor U0 (N_0,In_497,In_172);
or U1 (N_1,In_122,In_403);
nand U2 (N_2,In_218,In_224);
nand U3 (N_3,In_204,In_390);
or U4 (N_4,In_202,In_6);
nor U5 (N_5,In_217,In_427);
and U6 (N_6,In_467,In_103);
and U7 (N_7,In_285,In_39);
nand U8 (N_8,In_64,In_233);
nor U9 (N_9,In_384,In_445);
xnor U10 (N_10,In_489,In_215);
or U11 (N_11,In_387,In_100);
or U12 (N_12,In_66,In_148);
nand U13 (N_13,In_373,In_362);
and U14 (N_14,In_134,In_53);
nand U15 (N_15,In_251,In_196);
nor U16 (N_16,In_276,In_197);
or U17 (N_17,In_42,In_379);
or U18 (N_18,In_443,In_207);
nand U19 (N_19,In_406,In_5);
and U20 (N_20,In_397,In_43);
nand U21 (N_21,In_128,In_350);
nand U22 (N_22,In_83,In_189);
nand U23 (N_23,In_319,In_392);
or U24 (N_24,In_293,In_372);
and U25 (N_25,In_322,In_308);
or U26 (N_26,In_382,In_284);
xor U27 (N_27,In_367,In_349);
or U28 (N_28,In_470,In_454);
nand U29 (N_29,In_368,In_112);
and U30 (N_30,In_416,In_330);
or U31 (N_31,In_482,In_296);
nor U32 (N_32,In_429,In_360);
nand U33 (N_33,In_81,In_272);
nand U34 (N_34,In_184,In_463);
nor U35 (N_35,In_117,In_311);
and U36 (N_36,In_388,In_194);
nand U37 (N_37,In_331,In_94);
nor U38 (N_38,In_212,In_213);
nor U39 (N_39,In_97,In_313);
or U40 (N_40,In_341,In_306);
nand U41 (N_41,In_491,In_274);
nor U42 (N_42,In_474,In_118);
nand U43 (N_43,In_23,In_89);
and U44 (N_44,In_459,In_40);
nor U45 (N_45,In_453,In_366);
or U46 (N_46,In_420,In_49);
nor U47 (N_47,In_243,In_358);
nand U48 (N_48,In_369,In_398);
or U49 (N_49,In_492,In_314);
nand U50 (N_50,In_464,In_124);
xor U51 (N_51,In_364,In_60);
nand U52 (N_52,In_37,In_150);
nor U53 (N_53,In_411,In_149);
or U54 (N_54,In_252,In_32);
or U55 (N_55,In_413,In_180);
nor U56 (N_56,In_170,In_26);
and U57 (N_57,In_163,In_181);
nor U58 (N_58,In_267,In_242);
nand U59 (N_59,In_232,In_316);
and U60 (N_60,In_383,In_50);
nand U61 (N_61,In_237,In_323);
nand U62 (N_62,In_195,In_381);
nand U63 (N_63,In_262,In_98);
nor U64 (N_64,In_404,In_386);
nor U65 (N_65,In_269,In_486);
nor U66 (N_66,In_412,In_80);
and U67 (N_67,In_498,In_407);
nand U68 (N_68,In_438,In_255);
nand U69 (N_69,In_123,In_258);
and U70 (N_70,In_54,In_2);
or U71 (N_71,In_176,In_461);
and U72 (N_72,In_199,In_10);
nand U73 (N_73,In_77,In_290);
or U74 (N_74,In_281,In_286);
and U75 (N_75,In_72,In_88);
or U76 (N_76,In_265,In_275);
or U77 (N_77,In_444,In_496);
and U78 (N_78,In_327,In_151);
or U79 (N_79,In_385,In_222);
xor U80 (N_80,In_315,In_347);
or U81 (N_81,In_428,In_377);
nor U82 (N_82,In_16,In_478);
and U83 (N_83,In_462,In_402);
or U84 (N_84,In_260,In_188);
nor U85 (N_85,In_9,In_154);
nor U86 (N_86,In_447,In_41);
and U87 (N_87,In_241,In_7);
nor U88 (N_88,In_423,In_465);
nand U89 (N_89,In_56,In_108);
and U90 (N_90,In_356,In_495);
and U91 (N_91,In_200,In_264);
or U92 (N_92,In_19,In_378);
and U93 (N_93,In_147,In_333);
and U94 (N_94,In_138,In_169);
and U95 (N_95,In_14,In_451);
or U96 (N_96,In_110,In_153);
or U97 (N_97,In_99,In_334);
or U98 (N_98,In_144,In_115);
or U99 (N_99,In_328,In_129);
nor U100 (N_100,In_305,N_89);
nand U101 (N_101,N_56,N_5);
and U102 (N_102,In_67,N_54);
xor U103 (N_103,In_292,N_90);
nor U104 (N_104,N_83,In_484);
nand U105 (N_105,In_320,In_307);
and U106 (N_106,In_399,In_488);
nand U107 (N_107,N_66,In_278);
nor U108 (N_108,N_43,In_294);
and U109 (N_109,N_23,In_125);
nor U110 (N_110,In_405,In_175);
nand U111 (N_111,In_493,N_59);
or U112 (N_112,In_321,In_186);
or U113 (N_113,In_279,N_42);
nor U114 (N_114,In_90,In_121);
nor U115 (N_115,In_177,In_193);
nand U116 (N_116,In_92,In_352);
nor U117 (N_117,In_139,In_211);
or U118 (N_118,In_337,In_299);
nor U119 (N_119,In_220,In_174);
nor U120 (N_120,In_155,In_244);
nor U121 (N_121,In_228,In_18);
nor U122 (N_122,In_430,In_436);
nor U123 (N_123,N_44,In_143);
and U124 (N_124,In_410,In_164);
nand U125 (N_125,In_400,In_257);
nor U126 (N_126,In_415,In_389);
and U127 (N_127,N_37,In_348);
and U128 (N_128,N_45,N_1);
nor U129 (N_129,In_158,In_119);
nor U130 (N_130,N_96,N_87);
or U131 (N_131,In_70,In_216);
or U132 (N_132,In_318,In_11);
or U133 (N_133,In_62,In_107);
and U134 (N_134,In_229,In_152);
and U135 (N_135,In_309,N_32);
nor U136 (N_136,N_40,In_471);
and U137 (N_137,In_345,In_393);
and U138 (N_138,In_485,In_408);
nor U139 (N_139,In_69,In_391);
nand U140 (N_140,In_190,In_450);
nor U141 (N_141,In_376,In_51);
or U142 (N_142,In_396,N_2);
nor U143 (N_143,In_487,In_490);
or U144 (N_144,In_231,In_234);
nor U145 (N_145,In_442,In_236);
and U146 (N_146,In_424,In_256);
nand U147 (N_147,N_27,In_456);
nand U148 (N_148,In_375,In_36);
and U149 (N_149,N_71,In_288);
nor U150 (N_150,In_426,N_3);
and U151 (N_151,In_95,In_418);
nor U152 (N_152,In_93,In_291);
and U153 (N_153,In_17,In_57);
and U154 (N_154,In_221,In_380);
nor U155 (N_155,In_86,N_78);
nand U156 (N_156,N_74,In_351);
xor U157 (N_157,N_52,In_120);
nor U158 (N_158,In_126,N_92);
nor U159 (N_159,N_70,In_38);
and U160 (N_160,In_287,N_29);
nor U161 (N_161,In_13,In_261);
and U162 (N_162,N_81,In_45);
nand U163 (N_163,In_340,N_72);
nor U164 (N_164,In_46,In_431);
nor U165 (N_165,In_61,N_30);
nor U166 (N_166,N_34,In_414);
and U167 (N_167,N_65,In_326);
nor U168 (N_168,N_20,In_85);
and U169 (N_169,In_223,In_310);
nand U170 (N_170,In_27,In_344);
and U171 (N_171,In_355,In_179);
or U172 (N_172,In_329,In_171);
nand U173 (N_173,In_109,N_85);
nor U174 (N_174,In_157,N_97);
and U175 (N_175,In_185,N_94);
nor U176 (N_176,In_370,N_95);
nor U177 (N_177,In_15,In_133);
nor U178 (N_178,In_448,In_214);
nand U179 (N_179,In_289,In_302);
nand U180 (N_180,N_6,In_167);
nor U181 (N_181,N_62,In_401);
nor U182 (N_182,In_254,N_76);
nor U183 (N_183,In_198,N_58);
nor U184 (N_184,In_253,In_104);
or U185 (N_185,In_28,In_187);
or U186 (N_186,In_455,In_499);
nand U187 (N_187,N_80,In_357);
nand U188 (N_188,In_248,In_162);
nand U189 (N_189,N_8,In_82);
nor U190 (N_190,In_468,In_91);
and U191 (N_191,N_33,In_342);
and U192 (N_192,N_21,In_483);
or U193 (N_193,N_75,N_28);
and U194 (N_194,In_20,N_12);
and U195 (N_195,In_249,In_280);
nand U196 (N_196,In_63,In_74);
nand U197 (N_197,In_59,In_441);
nor U198 (N_198,In_75,N_82);
or U199 (N_199,In_114,In_475);
or U200 (N_200,N_11,N_39);
and U201 (N_201,N_143,N_145);
nor U202 (N_202,In_282,N_13);
nor U203 (N_203,N_114,In_12);
or U204 (N_204,N_171,In_127);
or U205 (N_205,N_184,N_146);
or U206 (N_206,N_131,In_208);
and U207 (N_207,In_266,N_50);
and U208 (N_208,In_419,In_141);
nor U209 (N_209,In_363,In_226);
or U210 (N_210,In_161,N_77);
nor U211 (N_211,N_183,N_161);
xor U212 (N_212,N_10,In_359);
or U213 (N_213,N_129,In_371);
nor U214 (N_214,N_4,N_195);
or U215 (N_215,In_25,In_469);
nand U216 (N_216,N_35,In_191);
nor U217 (N_217,In_245,In_55);
nor U218 (N_218,In_235,N_111);
or U219 (N_219,N_125,N_180);
or U220 (N_220,In_480,N_137);
nand U221 (N_221,In_271,In_168);
nand U222 (N_222,N_176,In_84);
nor U223 (N_223,In_324,N_153);
or U224 (N_224,N_22,In_277);
or U225 (N_225,In_106,In_201);
or U226 (N_226,N_196,In_140);
nand U227 (N_227,In_142,N_79);
and U228 (N_228,N_110,In_417);
or U229 (N_229,N_69,N_194);
nor U230 (N_230,N_119,In_78);
nor U231 (N_231,In_303,In_325);
nor U232 (N_232,In_76,In_65);
nand U233 (N_233,N_19,In_210);
or U234 (N_234,In_166,N_0);
and U235 (N_235,N_166,N_168);
nand U236 (N_236,N_14,In_192);
nor U237 (N_237,In_209,N_36);
nor U238 (N_238,In_111,N_106);
nor U239 (N_239,In_52,N_107);
nor U240 (N_240,N_93,N_126);
nand U241 (N_241,In_297,In_68);
or U242 (N_242,N_118,In_48);
or U243 (N_243,N_18,N_141);
or U244 (N_244,In_434,N_158);
nand U245 (N_245,N_91,In_440);
or U246 (N_246,N_60,N_55);
nand U247 (N_247,In_268,In_263);
nor U248 (N_248,N_154,N_136);
nand U249 (N_249,N_177,N_86);
nand U250 (N_250,In_227,N_172);
nand U251 (N_251,N_144,In_466);
or U252 (N_252,In_101,In_304);
nand U253 (N_253,N_187,In_270);
nand U254 (N_254,In_259,N_115);
and U255 (N_255,N_26,In_132);
and U256 (N_256,In_301,N_38);
and U257 (N_257,In_460,N_127);
nand U258 (N_258,N_165,N_122);
or U259 (N_259,In_79,In_3);
nand U260 (N_260,In_145,In_395);
nor U261 (N_261,N_169,In_452);
nor U262 (N_262,N_84,N_191);
and U263 (N_263,N_189,In_247);
nor U264 (N_264,In_35,In_203);
and U265 (N_265,In_102,N_63);
nor U266 (N_266,N_150,N_121);
nand U267 (N_267,In_335,In_178);
and U268 (N_268,N_160,N_120);
and U269 (N_269,In_361,In_239);
or U270 (N_270,N_103,In_47);
nor U271 (N_271,N_102,In_422);
and U272 (N_272,In_439,In_8);
nor U273 (N_273,N_178,N_98);
and U274 (N_274,N_192,In_312);
nor U275 (N_275,N_113,In_116);
and U276 (N_276,In_71,N_148);
nand U277 (N_277,N_101,N_181);
nand U278 (N_278,N_135,N_112);
or U279 (N_279,In_130,In_332);
or U280 (N_280,In_33,N_57);
nor U281 (N_281,N_9,N_104);
nor U282 (N_282,N_167,N_124);
nand U283 (N_283,In_137,N_173);
xor U284 (N_284,N_51,In_425);
nor U285 (N_285,N_157,In_230);
nor U286 (N_286,In_353,N_188);
or U287 (N_287,N_53,In_338);
and U288 (N_288,In_457,In_31);
nand U289 (N_289,In_476,N_49);
or U290 (N_290,In_205,In_24);
and U291 (N_291,In_160,N_25);
or U292 (N_292,In_96,N_164);
nand U293 (N_293,N_128,In_173);
nor U294 (N_294,In_58,N_68);
nor U295 (N_295,In_30,In_29);
and U296 (N_296,In_135,In_346);
and U297 (N_297,In_22,In_433);
nor U298 (N_298,N_17,In_354);
and U299 (N_299,N_24,N_133);
and U300 (N_300,N_233,N_47);
nand U301 (N_301,N_247,N_215);
nor U302 (N_302,N_155,N_263);
nand U303 (N_303,N_240,N_99);
and U304 (N_304,N_206,In_156);
and U305 (N_305,N_253,N_209);
nor U306 (N_306,N_152,N_238);
nand U307 (N_307,In_21,N_174);
nand U308 (N_308,N_219,N_139);
and U309 (N_309,In_183,In_300);
and U310 (N_310,N_197,N_130);
and U311 (N_311,N_230,N_271);
and U312 (N_312,N_286,In_225);
and U313 (N_313,In_159,N_272);
or U314 (N_314,N_276,N_258);
nor U315 (N_315,N_248,N_190);
and U316 (N_316,N_222,In_34);
and U317 (N_317,N_198,N_204);
nor U318 (N_318,In_273,N_123);
or U319 (N_319,N_229,N_260);
or U320 (N_320,N_218,In_219);
and U321 (N_321,N_252,N_67);
or U322 (N_322,N_16,N_296);
nand U323 (N_323,In_146,N_277);
nand U324 (N_324,N_15,N_298);
nand U325 (N_325,N_227,N_175);
and U326 (N_326,N_64,N_285);
nand U327 (N_327,In_458,N_142);
nand U328 (N_328,N_283,N_294);
or U329 (N_329,N_239,In_1);
or U330 (N_330,N_138,N_156);
nand U331 (N_331,N_273,In_283);
nand U332 (N_332,N_278,N_216);
nor U333 (N_333,In_44,N_246);
and U334 (N_334,In_105,N_41);
nand U335 (N_335,N_291,N_262);
and U336 (N_336,N_226,N_88);
or U337 (N_337,N_147,In_449);
nor U338 (N_338,In_298,N_162);
nand U339 (N_339,N_185,N_236);
nor U340 (N_340,N_245,N_225);
nand U341 (N_341,N_282,In_437);
and U342 (N_342,N_241,In_165);
nor U343 (N_343,In_336,N_186);
nand U344 (N_344,N_31,In_409);
or U345 (N_345,N_280,N_274);
nand U346 (N_346,N_289,N_250);
and U347 (N_347,N_269,N_116);
and U348 (N_348,In_339,N_109);
nor U349 (N_349,In_472,In_479);
and U350 (N_350,N_46,N_200);
or U351 (N_351,In_0,N_231);
and U352 (N_352,N_179,N_265);
nor U353 (N_353,In_317,N_151);
and U354 (N_354,N_117,In_295);
nand U355 (N_355,N_105,N_48);
nor U356 (N_356,N_140,N_7);
and U357 (N_357,N_201,In_113);
nor U358 (N_358,N_224,N_259);
nor U359 (N_359,In_394,N_255);
nand U360 (N_360,N_212,N_182);
nand U361 (N_361,N_228,N_221);
nand U362 (N_362,N_264,N_293);
nor U363 (N_363,N_208,In_481);
nor U364 (N_364,N_73,N_261);
nor U365 (N_365,N_213,In_250);
or U366 (N_366,N_256,N_243);
nor U367 (N_367,In_494,In_435);
nor U368 (N_368,N_132,N_203);
nor U369 (N_369,N_290,N_223);
nor U370 (N_370,In_421,N_287);
or U371 (N_371,N_237,N_249);
nand U372 (N_372,N_61,N_266);
and U373 (N_373,N_149,N_108);
nor U374 (N_374,N_275,In_131);
nand U375 (N_375,N_299,N_210);
and U376 (N_376,N_217,In_365);
xor U377 (N_377,In_182,In_432);
nand U378 (N_378,N_292,N_235);
and U379 (N_379,N_254,In_246);
nand U380 (N_380,N_220,N_214);
nand U381 (N_381,In_343,N_297);
and U382 (N_382,N_207,N_257);
nor U383 (N_383,N_281,N_193);
nand U384 (N_384,In_240,In_238);
nor U385 (N_385,N_163,N_199);
and U386 (N_386,In_477,In_473);
or U387 (N_387,N_205,In_73);
and U388 (N_388,In_446,N_134);
nand U389 (N_389,N_100,N_211);
nor U390 (N_390,In_206,N_270);
nand U391 (N_391,N_244,N_295);
nand U392 (N_392,N_159,N_288);
nor U393 (N_393,N_279,N_268);
nor U394 (N_394,N_284,In_87);
or U395 (N_395,N_234,In_136);
nor U396 (N_396,N_232,In_374);
and U397 (N_397,In_4,N_202);
or U398 (N_398,N_242,N_267);
nand U399 (N_399,N_251,N_170);
nand U400 (N_400,N_317,N_304);
or U401 (N_401,N_325,N_301);
xnor U402 (N_402,N_378,N_315);
nor U403 (N_403,N_361,N_374);
nand U404 (N_404,N_362,N_327);
and U405 (N_405,N_329,N_397);
nand U406 (N_406,N_328,N_371);
nor U407 (N_407,N_308,N_330);
nand U408 (N_408,N_326,N_372);
nand U409 (N_409,N_360,N_346);
nand U410 (N_410,N_386,N_373);
nor U411 (N_411,N_332,N_354);
nand U412 (N_412,N_313,N_356);
or U413 (N_413,N_394,N_390);
and U414 (N_414,N_365,N_349);
nor U415 (N_415,N_369,N_359);
or U416 (N_416,N_380,N_366);
nor U417 (N_417,N_344,N_385);
or U418 (N_418,N_311,N_364);
nor U419 (N_419,N_336,N_342);
nor U420 (N_420,N_314,N_333);
or U421 (N_421,N_352,N_368);
and U422 (N_422,N_399,N_307);
and U423 (N_423,N_320,N_334);
nand U424 (N_424,N_388,N_358);
nand U425 (N_425,N_363,N_377);
and U426 (N_426,N_351,N_389);
nand U427 (N_427,N_347,N_319);
and U428 (N_428,N_393,N_387);
nor U429 (N_429,N_331,N_338);
and U430 (N_430,N_343,N_306);
and U431 (N_431,N_341,N_337);
and U432 (N_432,N_357,N_335);
nor U433 (N_433,N_391,N_379);
and U434 (N_434,N_316,N_350);
and U435 (N_435,N_345,N_395);
nor U436 (N_436,N_370,N_384);
nor U437 (N_437,N_367,N_322);
and U438 (N_438,N_398,N_318);
or U439 (N_439,N_312,N_339);
nor U440 (N_440,N_355,N_305);
nor U441 (N_441,N_309,N_323);
and U442 (N_442,N_324,N_348);
nand U443 (N_443,N_310,N_382);
nand U444 (N_444,N_302,N_321);
nand U445 (N_445,N_303,N_376);
nor U446 (N_446,N_340,N_392);
and U447 (N_447,N_383,N_353);
nor U448 (N_448,N_300,N_381);
nand U449 (N_449,N_396,N_375);
or U450 (N_450,N_367,N_399);
nor U451 (N_451,N_388,N_397);
or U452 (N_452,N_359,N_313);
and U453 (N_453,N_317,N_330);
nor U454 (N_454,N_339,N_349);
nor U455 (N_455,N_330,N_352);
nand U456 (N_456,N_355,N_343);
nor U457 (N_457,N_370,N_342);
and U458 (N_458,N_345,N_322);
or U459 (N_459,N_372,N_373);
and U460 (N_460,N_330,N_375);
or U461 (N_461,N_360,N_370);
nand U462 (N_462,N_326,N_373);
nand U463 (N_463,N_342,N_390);
or U464 (N_464,N_323,N_392);
nand U465 (N_465,N_342,N_379);
nor U466 (N_466,N_353,N_334);
nor U467 (N_467,N_360,N_341);
or U468 (N_468,N_395,N_350);
nor U469 (N_469,N_367,N_328);
or U470 (N_470,N_326,N_304);
nor U471 (N_471,N_354,N_341);
and U472 (N_472,N_329,N_352);
or U473 (N_473,N_383,N_330);
nor U474 (N_474,N_331,N_337);
nor U475 (N_475,N_334,N_387);
and U476 (N_476,N_308,N_385);
and U477 (N_477,N_387,N_349);
or U478 (N_478,N_377,N_386);
nand U479 (N_479,N_342,N_307);
and U480 (N_480,N_312,N_357);
or U481 (N_481,N_355,N_399);
or U482 (N_482,N_366,N_354);
nand U483 (N_483,N_361,N_336);
nand U484 (N_484,N_332,N_310);
nand U485 (N_485,N_371,N_351);
and U486 (N_486,N_378,N_326);
nand U487 (N_487,N_389,N_312);
nor U488 (N_488,N_392,N_369);
and U489 (N_489,N_385,N_313);
nand U490 (N_490,N_315,N_355);
and U491 (N_491,N_398,N_345);
or U492 (N_492,N_341,N_336);
nor U493 (N_493,N_343,N_380);
nand U494 (N_494,N_369,N_363);
or U495 (N_495,N_390,N_335);
nor U496 (N_496,N_359,N_336);
or U497 (N_497,N_327,N_320);
or U498 (N_498,N_344,N_318);
xnor U499 (N_499,N_372,N_307);
nand U500 (N_500,N_408,N_403);
or U501 (N_501,N_495,N_481);
nor U502 (N_502,N_478,N_492);
or U503 (N_503,N_494,N_440);
or U504 (N_504,N_467,N_426);
and U505 (N_505,N_487,N_486);
nand U506 (N_506,N_433,N_416);
nor U507 (N_507,N_483,N_401);
nand U508 (N_508,N_465,N_437);
xnor U509 (N_509,N_493,N_459);
nand U510 (N_510,N_452,N_475);
or U511 (N_511,N_407,N_446);
nand U512 (N_512,N_461,N_442);
nor U513 (N_513,N_449,N_458);
nand U514 (N_514,N_431,N_485);
or U515 (N_515,N_472,N_466);
nor U516 (N_516,N_457,N_439);
and U517 (N_517,N_456,N_482);
nor U518 (N_518,N_435,N_468);
nand U519 (N_519,N_438,N_470);
nand U520 (N_520,N_424,N_417);
nand U521 (N_521,N_432,N_491);
nor U522 (N_522,N_436,N_474);
nor U523 (N_523,N_496,N_414);
or U524 (N_524,N_413,N_455);
and U525 (N_525,N_447,N_430);
xor U526 (N_526,N_400,N_471);
or U527 (N_527,N_405,N_476);
and U528 (N_528,N_410,N_484);
nand U529 (N_529,N_477,N_404);
nor U530 (N_530,N_463,N_409);
and U531 (N_531,N_488,N_497);
or U532 (N_532,N_479,N_443);
nor U533 (N_533,N_445,N_454);
and U534 (N_534,N_460,N_499);
and U535 (N_535,N_427,N_490);
or U536 (N_536,N_489,N_453);
or U537 (N_537,N_448,N_441);
or U538 (N_538,N_421,N_469);
nand U539 (N_539,N_411,N_418);
nor U540 (N_540,N_464,N_402);
and U541 (N_541,N_498,N_428);
and U542 (N_542,N_444,N_420);
or U543 (N_543,N_412,N_473);
or U544 (N_544,N_462,N_429);
nand U545 (N_545,N_422,N_423);
and U546 (N_546,N_406,N_419);
and U547 (N_547,N_434,N_450);
or U548 (N_548,N_425,N_415);
or U549 (N_549,N_451,N_480);
or U550 (N_550,N_442,N_463);
nand U551 (N_551,N_484,N_451);
and U552 (N_552,N_421,N_433);
and U553 (N_553,N_426,N_493);
or U554 (N_554,N_473,N_435);
nand U555 (N_555,N_450,N_480);
or U556 (N_556,N_436,N_411);
and U557 (N_557,N_438,N_461);
nand U558 (N_558,N_414,N_468);
or U559 (N_559,N_403,N_470);
nor U560 (N_560,N_430,N_495);
and U561 (N_561,N_426,N_471);
nor U562 (N_562,N_433,N_408);
nor U563 (N_563,N_456,N_459);
nand U564 (N_564,N_408,N_479);
and U565 (N_565,N_409,N_422);
or U566 (N_566,N_452,N_427);
and U567 (N_567,N_420,N_469);
and U568 (N_568,N_469,N_413);
and U569 (N_569,N_489,N_408);
and U570 (N_570,N_409,N_486);
or U571 (N_571,N_415,N_437);
or U572 (N_572,N_404,N_467);
or U573 (N_573,N_425,N_444);
or U574 (N_574,N_469,N_468);
and U575 (N_575,N_400,N_461);
and U576 (N_576,N_470,N_463);
or U577 (N_577,N_465,N_460);
nor U578 (N_578,N_433,N_431);
and U579 (N_579,N_422,N_492);
and U580 (N_580,N_477,N_466);
and U581 (N_581,N_454,N_429);
nand U582 (N_582,N_413,N_433);
nor U583 (N_583,N_443,N_466);
or U584 (N_584,N_430,N_467);
and U585 (N_585,N_469,N_416);
nor U586 (N_586,N_490,N_436);
or U587 (N_587,N_405,N_495);
and U588 (N_588,N_488,N_469);
or U589 (N_589,N_492,N_406);
nor U590 (N_590,N_439,N_480);
nor U591 (N_591,N_498,N_492);
or U592 (N_592,N_451,N_472);
nor U593 (N_593,N_449,N_457);
or U594 (N_594,N_472,N_433);
nor U595 (N_595,N_463,N_483);
or U596 (N_596,N_467,N_496);
and U597 (N_597,N_431,N_444);
nand U598 (N_598,N_487,N_497);
nand U599 (N_599,N_450,N_464);
xor U600 (N_600,N_534,N_511);
and U601 (N_601,N_547,N_559);
nor U602 (N_602,N_525,N_538);
nor U603 (N_603,N_500,N_518);
or U604 (N_604,N_508,N_517);
nor U605 (N_605,N_543,N_564);
nor U606 (N_606,N_573,N_545);
and U607 (N_607,N_521,N_548);
and U608 (N_608,N_533,N_565);
or U609 (N_609,N_544,N_503);
nand U610 (N_610,N_551,N_584);
nor U611 (N_611,N_550,N_501);
and U612 (N_612,N_574,N_599);
and U613 (N_613,N_571,N_592);
nand U614 (N_614,N_590,N_583);
and U615 (N_615,N_562,N_556);
or U616 (N_616,N_549,N_568);
nand U617 (N_617,N_595,N_581);
nand U618 (N_618,N_585,N_578);
nor U619 (N_619,N_579,N_529);
nand U620 (N_620,N_558,N_519);
or U621 (N_621,N_554,N_510);
nand U622 (N_622,N_566,N_502);
or U623 (N_623,N_507,N_506);
xnor U624 (N_624,N_539,N_561);
or U625 (N_625,N_509,N_535);
nor U626 (N_626,N_580,N_582);
nand U627 (N_627,N_555,N_567);
nand U628 (N_628,N_589,N_531);
and U629 (N_629,N_575,N_536);
nor U630 (N_630,N_546,N_557);
and U631 (N_631,N_537,N_593);
or U632 (N_632,N_597,N_570);
nor U633 (N_633,N_594,N_504);
nor U634 (N_634,N_588,N_523);
and U635 (N_635,N_520,N_587);
xnor U636 (N_636,N_577,N_553);
and U637 (N_637,N_591,N_522);
nor U638 (N_638,N_552,N_560);
nand U639 (N_639,N_524,N_514);
and U640 (N_640,N_576,N_512);
nor U641 (N_641,N_527,N_528);
nand U642 (N_642,N_598,N_513);
nand U643 (N_643,N_586,N_596);
and U644 (N_644,N_540,N_572);
nand U645 (N_645,N_569,N_541);
nand U646 (N_646,N_516,N_530);
nand U647 (N_647,N_505,N_563);
nand U648 (N_648,N_542,N_515);
and U649 (N_649,N_532,N_526);
or U650 (N_650,N_575,N_542);
nor U651 (N_651,N_564,N_573);
or U652 (N_652,N_534,N_531);
and U653 (N_653,N_569,N_581);
or U654 (N_654,N_535,N_575);
nor U655 (N_655,N_553,N_580);
or U656 (N_656,N_533,N_536);
nand U657 (N_657,N_571,N_563);
or U658 (N_658,N_518,N_582);
or U659 (N_659,N_591,N_560);
nor U660 (N_660,N_534,N_524);
or U661 (N_661,N_590,N_504);
or U662 (N_662,N_515,N_571);
nand U663 (N_663,N_589,N_503);
or U664 (N_664,N_590,N_514);
and U665 (N_665,N_514,N_547);
and U666 (N_666,N_504,N_580);
nor U667 (N_667,N_569,N_561);
nor U668 (N_668,N_577,N_588);
or U669 (N_669,N_553,N_599);
nand U670 (N_670,N_581,N_562);
or U671 (N_671,N_533,N_531);
nand U672 (N_672,N_505,N_506);
nand U673 (N_673,N_509,N_505);
nor U674 (N_674,N_568,N_546);
and U675 (N_675,N_507,N_582);
and U676 (N_676,N_581,N_505);
nor U677 (N_677,N_537,N_581);
nand U678 (N_678,N_521,N_525);
nand U679 (N_679,N_566,N_532);
and U680 (N_680,N_577,N_540);
nor U681 (N_681,N_549,N_592);
or U682 (N_682,N_573,N_599);
nor U683 (N_683,N_503,N_559);
or U684 (N_684,N_567,N_592);
nand U685 (N_685,N_550,N_547);
and U686 (N_686,N_591,N_558);
nor U687 (N_687,N_593,N_511);
nand U688 (N_688,N_553,N_552);
nand U689 (N_689,N_588,N_585);
and U690 (N_690,N_500,N_554);
nor U691 (N_691,N_562,N_598);
and U692 (N_692,N_557,N_587);
and U693 (N_693,N_529,N_585);
and U694 (N_694,N_534,N_552);
or U695 (N_695,N_537,N_517);
or U696 (N_696,N_590,N_541);
or U697 (N_697,N_563,N_529);
or U698 (N_698,N_576,N_586);
and U699 (N_699,N_511,N_553);
or U700 (N_700,N_690,N_603);
nor U701 (N_701,N_614,N_661);
nor U702 (N_702,N_618,N_652);
nand U703 (N_703,N_638,N_653);
nor U704 (N_704,N_612,N_684);
nand U705 (N_705,N_639,N_688);
and U706 (N_706,N_629,N_608);
nor U707 (N_707,N_600,N_602);
or U708 (N_708,N_672,N_685);
nor U709 (N_709,N_683,N_637);
nand U710 (N_710,N_601,N_644);
and U711 (N_711,N_636,N_664);
or U712 (N_712,N_607,N_660);
nor U713 (N_713,N_673,N_650);
or U714 (N_714,N_674,N_658);
nand U715 (N_715,N_669,N_633);
nand U716 (N_716,N_611,N_694);
and U717 (N_717,N_682,N_663);
or U718 (N_718,N_656,N_628);
or U719 (N_719,N_651,N_692);
or U720 (N_720,N_666,N_689);
nand U721 (N_721,N_686,N_691);
nand U722 (N_722,N_693,N_615);
nor U723 (N_723,N_624,N_631);
nand U724 (N_724,N_632,N_675);
or U725 (N_725,N_617,N_670);
nand U726 (N_726,N_665,N_662);
or U727 (N_727,N_613,N_619);
nand U728 (N_728,N_627,N_643);
or U729 (N_729,N_626,N_655);
or U730 (N_730,N_604,N_678);
and U731 (N_731,N_654,N_695);
or U732 (N_732,N_630,N_687);
nand U733 (N_733,N_649,N_610);
nor U734 (N_734,N_648,N_641);
and U735 (N_735,N_640,N_699);
and U736 (N_736,N_698,N_659);
nor U737 (N_737,N_635,N_667);
nor U738 (N_738,N_634,N_622);
nand U739 (N_739,N_621,N_681);
nand U740 (N_740,N_680,N_645);
and U741 (N_741,N_646,N_679);
or U742 (N_742,N_676,N_671);
nor U743 (N_743,N_677,N_668);
nand U744 (N_744,N_606,N_609);
and U745 (N_745,N_620,N_657);
or U746 (N_746,N_616,N_696);
or U747 (N_747,N_697,N_605);
and U748 (N_748,N_642,N_625);
and U749 (N_749,N_623,N_647);
nand U750 (N_750,N_683,N_645);
or U751 (N_751,N_678,N_695);
or U752 (N_752,N_645,N_622);
or U753 (N_753,N_663,N_638);
nor U754 (N_754,N_668,N_615);
nand U755 (N_755,N_651,N_632);
nand U756 (N_756,N_653,N_650);
or U757 (N_757,N_667,N_607);
and U758 (N_758,N_696,N_657);
nand U759 (N_759,N_647,N_678);
and U760 (N_760,N_603,N_637);
or U761 (N_761,N_682,N_611);
nand U762 (N_762,N_696,N_611);
or U763 (N_763,N_637,N_672);
or U764 (N_764,N_666,N_693);
or U765 (N_765,N_649,N_600);
or U766 (N_766,N_631,N_678);
or U767 (N_767,N_675,N_671);
nor U768 (N_768,N_626,N_642);
or U769 (N_769,N_610,N_696);
and U770 (N_770,N_611,N_628);
or U771 (N_771,N_627,N_645);
or U772 (N_772,N_615,N_621);
and U773 (N_773,N_608,N_621);
nand U774 (N_774,N_602,N_642);
or U775 (N_775,N_626,N_615);
and U776 (N_776,N_682,N_612);
or U777 (N_777,N_680,N_647);
nand U778 (N_778,N_671,N_623);
nand U779 (N_779,N_618,N_658);
nor U780 (N_780,N_630,N_624);
nand U781 (N_781,N_640,N_677);
and U782 (N_782,N_624,N_638);
or U783 (N_783,N_614,N_617);
nand U784 (N_784,N_681,N_647);
nand U785 (N_785,N_601,N_685);
or U786 (N_786,N_673,N_674);
or U787 (N_787,N_602,N_663);
or U788 (N_788,N_621,N_695);
nand U789 (N_789,N_688,N_652);
or U790 (N_790,N_694,N_646);
and U791 (N_791,N_637,N_642);
nand U792 (N_792,N_662,N_663);
and U793 (N_793,N_622,N_690);
nand U794 (N_794,N_640,N_654);
nand U795 (N_795,N_655,N_666);
nand U796 (N_796,N_638,N_699);
nand U797 (N_797,N_611,N_641);
nor U798 (N_798,N_613,N_611);
and U799 (N_799,N_613,N_680);
nand U800 (N_800,N_713,N_744);
or U801 (N_801,N_743,N_781);
nor U802 (N_802,N_785,N_711);
nor U803 (N_803,N_731,N_786);
and U804 (N_804,N_765,N_764);
nand U805 (N_805,N_715,N_756);
nand U806 (N_806,N_772,N_746);
or U807 (N_807,N_799,N_708);
or U808 (N_808,N_794,N_728);
nor U809 (N_809,N_701,N_748);
and U810 (N_810,N_791,N_778);
nand U811 (N_811,N_766,N_740);
nor U812 (N_812,N_747,N_742);
nand U813 (N_813,N_755,N_792);
and U814 (N_814,N_779,N_733);
or U815 (N_815,N_768,N_771);
or U816 (N_816,N_723,N_754);
nand U817 (N_817,N_762,N_725);
nor U818 (N_818,N_714,N_737);
and U819 (N_819,N_710,N_790);
xnor U820 (N_820,N_752,N_727);
and U821 (N_821,N_775,N_787);
nand U822 (N_822,N_735,N_780);
nor U823 (N_823,N_770,N_793);
nor U824 (N_824,N_763,N_773);
nand U825 (N_825,N_767,N_798);
and U826 (N_826,N_745,N_783);
nand U827 (N_827,N_797,N_730);
nand U828 (N_828,N_720,N_703);
or U829 (N_829,N_719,N_758);
and U830 (N_830,N_789,N_784);
nand U831 (N_831,N_760,N_736);
nor U832 (N_832,N_729,N_712);
nor U833 (N_833,N_724,N_738);
and U834 (N_834,N_796,N_706);
nand U835 (N_835,N_717,N_761);
nand U836 (N_836,N_716,N_704);
and U837 (N_837,N_732,N_709);
xnor U838 (N_838,N_757,N_705);
and U839 (N_839,N_700,N_774);
and U840 (N_840,N_750,N_726);
nand U841 (N_841,N_734,N_722);
nor U842 (N_842,N_739,N_759);
nor U843 (N_843,N_776,N_753);
and U844 (N_844,N_769,N_718);
nor U845 (N_845,N_782,N_741);
and U846 (N_846,N_702,N_707);
nor U847 (N_847,N_749,N_788);
or U848 (N_848,N_751,N_777);
nand U849 (N_849,N_795,N_721);
and U850 (N_850,N_705,N_720);
nand U851 (N_851,N_755,N_791);
or U852 (N_852,N_710,N_747);
and U853 (N_853,N_747,N_790);
or U854 (N_854,N_732,N_707);
or U855 (N_855,N_756,N_700);
nand U856 (N_856,N_720,N_799);
nor U857 (N_857,N_789,N_739);
and U858 (N_858,N_704,N_780);
or U859 (N_859,N_781,N_766);
and U860 (N_860,N_775,N_770);
or U861 (N_861,N_758,N_746);
nor U862 (N_862,N_771,N_701);
nand U863 (N_863,N_710,N_717);
nand U864 (N_864,N_744,N_770);
nand U865 (N_865,N_739,N_715);
nor U866 (N_866,N_780,N_747);
nand U867 (N_867,N_741,N_778);
xnor U868 (N_868,N_711,N_784);
and U869 (N_869,N_786,N_775);
nor U870 (N_870,N_786,N_794);
nand U871 (N_871,N_733,N_747);
and U872 (N_872,N_731,N_744);
nand U873 (N_873,N_753,N_766);
nor U874 (N_874,N_731,N_771);
nor U875 (N_875,N_714,N_758);
or U876 (N_876,N_778,N_752);
or U877 (N_877,N_760,N_770);
nand U878 (N_878,N_724,N_778);
or U879 (N_879,N_708,N_780);
and U880 (N_880,N_711,N_780);
or U881 (N_881,N_708,N_750);
or U882 (N_882,N_708,N_716);
or U883 (N_883,N_708,N_768);
xnor U884 (N_884,N_702,N_733);
nand U885 (N_885,N_706,N_714);
or U886 (N_886,N_782,N_744);
or U887 (N_887,N_774,N_743);
and U888 (N_888,N_740,N_785);
nand U889 (N_889,N_751,N_778);
and U890 (N_890,N_733,N_713);
and U891 (N_891,N_707,N_776);
or U892 (N_892,N_716,N_748);
or U893 (N_893,N_756,N_767);
nor U894 (N_894,N_776,N_748);
nor U895 (N_895,N_765,N_726);
or U896 (N_896,N_750,N_778);
nor U897 (N_897,N_700,N_759);
nand U898 (N_898,N_730,N_760);
and U899 (N_899,N_716,N_706);
nand U900 (N_900,N_846,N_847);
nor U901 (N_901,N_876,N_875);
nor U902 (N_902,N_838,N_853);
nand U903 (N_903,N_892,N_890);
xor U904 (N_904,N_808,N_850);
or U905 (N_905,N_865,N_822);
nand U906 (N_906,N_842,N_845);
or U907 (N_907,N_898,N_863);
nor U908 (N_908,N_818,N_823);
nor U909 (N_909,N_819,N_878);
nor U910 (N_910,N_827,N_805);
nor U911 (N_911,N_862,N_891);
nand U912 (N_912,N_854,N_896);
or U913 (N_913,N_835,N_800);
nor U914 (N_914,N_857,N_836);
or U915 (N_915,N_826,N_828);
nand U916 (N_916,N_874,N_871);
and U917 (N_917,N_877,N_848);
nor U918 (N_918,N_825,N_870);
nor U919 (N_919,N_851,N_859);
or U920 (N_920,N_893,N_899);
nor U921 (N_921,N_801,N_897);
or U922 (N_922,N_821,N_858);
and U923 (N_923,N_839,N_864);
or U924 (N_924,N_849,N_873);
nand U925 (N_925,N_802,N_806);
nand U926 (N_926,N_811,N_813);
nand U927 (N_927,N_880,N_814);
or U928 (N_928,N_883,N_832);
and U929 (N_929,N_841,N_879);
or U930 (N_930,N_887,N_895);
and U931 (N_931,N_815,N_834);
nor U932 (N_932,N_816,N_833);
and U933 (N_933,N_809,N_881);
nand U934 (N_934,N_888,N_885);
nand U935 (N_935,N_810,N_812);
nand U936 (N_936,N_852,N_894);
nand U937 (N_937,N_829,N_886);
nor U938 (N_938,N_817,N_807);
nor U939 (N_939,N_837,N_824);
nor U940 (N_940,N_844,N_860);
nand U941 (N_941,N_843,N_830);
or U942 (N_942,N_861,N_882);
nand U943 (N_943,N_804,N_866);
nor U944 (N_944,N_856,N_831);
and U945 (N_945,N_820,N_803);
or U946 (N_946,N_855,N_872);
and U947 (N_947,N_884,N_840);
or U948 (N_948,N_889,N_869);
nor U949 (N_949,N_867,N_868);
and U950 (N_950,N_864,N_844);
and U951 (N_951,N_810,N_831);
and U952 (N_952,N_888,N_811);
nand U953 (N_953,N_890,N_820);
nor U954 (N_954,N_858,N_896);
and U955 (N_955,N_888,N_837);
and U956 (N_956,N_853,N_890);
nand U957 (N_957,N_886,N_866);
nor U958 (N_958,N_844,N_808);
or U959 (N_959,N_892,N_836);
or U960 (N_960,N_808,N_893);
or U961 (N_961,N_805,N_812);
or U962 (N_962,N_846,N_858);
nand U963 (N_963,N_897,N_866);
nor U964 (N_964,N_857,N_816);
or U965 (N_965,N_855,N_843);
or U966 (N_966,N_844,N_858);
or U967 (N_967,N_853,N_825);
and U968 (N_968,N_821,N_827);
and U969 (N_969,N_812,N_883);
or U970 (N_970,N_898,N_871);
and U971 (N_971,N_877,N_888);
or U972 (N_972,N_832,N_871);
nor U973 (N_973,N_898,N_864);
or U974 (N_974,N_838,N_895);
nor U975 (N_975,N_881,N_825);
nand U976 (N_976,N_855,N_853);
or U977 (N_977,N_861,N_840);
and U978 (N_978,N_800,N_880);
or U979 (N_979,N_849,N_833);
and U980 (N_980,N_842,N_802);
nor U981 (N_981,N_887,N_860);
nor U982 (N_982,N_885,N_839);
nor U983 (N_983,N_859,N_867);
and U984 (N_984,N_813,N_870);
or U985 (N_985,N_824,N_899);
and U986 (N_986,N_885,N_865);
nor U987 (N_987,N_805,N_859);
and U988 (N_988,N_833,N_802);
or U989 (N_989,N_817,N_863);
nor U990 (N_990,N_828,N_865);
and U991 (N_991,N_843,N_860);
or U992 (N_992,N_878,N_858);
and U993 (N_993,N_850,N_869);
nand U994 (N_994,N_831,N_837);
and U995 (N_995,N_875,N_851);
or U996 (N_996,N_844,N_805);
nor U997 (N_997,N_812,N_890);
nand U998 (N_998,N_823,N_882);
nor U999 (N_999,N_899,N_815);
and U1000 (N_1000,N_964,N_933);
and U1001 (N_1001,N_940,N_922);
nand U1002 (N_1002,N_920,N_907);
or U1003 (N_1003,N_945,N_925);
and U1004 (N_1004,N_921,N_990);
or U1005 (N_1005,N_927,N_986);
or U1006 (N_1006,N_948,N_995);
nand U1007 (N_1007,N_961,N_987);
nor U1008 (N_1008,N_970,N_943);
or U1009 (N_1009,N_957,N_979);
nor U1010 (N_1010,N_909,N_962);
nor U1011 (N_1011,N_997,N_911);
and U1012 (N_1012,N_978,N_981);
nor U1013 (N_1013,N_919,N_930);
and U1014 (N_1014,N_912,N_992);
nand U1015 (N_1015,N_934,N_982);
or U1016 (N_1016,N_972,N_980);
nor U1017 (N_1017,N_908,N_941);
and U1018 (N_1018,N_917,N_946);
or U1019 (N_1019,N_984,N_913);
or U1020 (N_1020,N_983,N_942);
and U1021 (N_1021,N_910,N_936);
nand U1022 (N_1022,N_974,N_903);
or U1023 (N_1023,N_956,N_967);
and U1024 (N_1024,N_991,N_939);
nor U1025 (N_1025,N_955,N_985);
and U1026 (N_1026,N_904,N_900);
and U1027 (N_1027,N_944,N_965);
and U1028 (N_1028,N_906,N_938);
and U1029 (N_1029,N_994,N_916);
or U1030 (N_1030,N_969,N_928);
and U1031 (N_1031,N_973,N_953);
nand U1032 (N_1032,N_947,N_960);
nand U1033 (N_1033,N_989,N_966);
or U1034 (N_1034,N_915,N_918);
nand U1035 (N_1035,N_999,N_954);
nand U1036 (N_1036,N_923,N_950);
nand U1037 (N_1037,N_924,N_993);
nand U1038 (N_1038,N_926,N_977);
nor U1039 (N_1039,N_935,N_996);
or U1040 (N_1040,N_988,N_937);
nor U1041 (N_1041,N_901,N_976);
nor U1042 (N_1042,N_963,N_931);
and U1043 (N_1043,N_902,N_959);
xor U1044 (N_1044,N_951,N_975);
or U1045 (N_1045,N_914,N_998);
nand U1046 (N_1046,N_929,N_932);
nand U1047 (N_1047,N_905,N_971);
nand U1048 (N_1048,N_958,N_949);
or U1049 (N_1049,N_952,N_968);
nor U1050 (N_1050,N_987,N_988);
or U1051 (N_1051,N_955,N_960);
and U1052 (N_1052,N_993,N_994);
nor U1053 (N_1053,N_975,N_968);
nor U1054 (N_1054,N_987,N_981);
or U1055 (N_1055,N_943,N_936);
nor U1056 (N_1056,N_955,N_939);
or U1057 (N_1057,N_912,N_928);
and U1058 (N_1058,N_971,N_968);
and U1059 (N_1059,N_927,N_999);
and U1060 (N_1060,N_994,N_962);
or U1061 (N_1061,N_936,N_920);
nand U1062 (N_1062,N_918,N_901);
nand U1063 (N_1063,N_927,N_966);
nor U1064 (N_1064,N_994,N_995);
nor U1065 (N_1065,N_928,N_966);
and U1066 (N_1066,N_905,N_939);
nand U1067 (N_1067,N_928,N_901);
or U1068 (N_1068,N_981,N_944);
or U1069 (N_1069,N_943,N_920);
nor U1070 (N_1070,N_920,N_978);
or U1071 (N_1071,N_942,N_998);
or U1072 (N_1072,N_967,N_930);
nand U1073 (N_1073,N_969,N_986);
and U1074 (N_1074,N_959,N_912);
nor U1075 (N_1075,N_937,N_962);
or U1076 (N_1076,N_968,N_923);
and U1077 (N_1077,N_932,N_970);
or U1078 (N_1078,N_939,N_961);
nand U1079 (N_1079,N_951,N_915);
nor U1080 (N_1080,N_997,N_968);
and U1081 (N_1081,N_926,N_998);
nand U1082 (N_1082,N_925,N_956);
nand U1083 (N_1083,N_971,N_993);
nand U1084 (N_1084,N_907,N_957);
and U1085 (N_1085,N_968,N_957);
or U1086 (N_1086,N_935,N_918);
and U1087 (N_1087,N_937,N_972);
or U1088 (N_1088,N_983,N_967);
or U1089 (N_1089,N_900,N_996);
xor U1090 (N_1090,N_984,N_949);
nand U1091 (N_1091,N_925,N_957);
nand U1092 (N_1092,N_956,N_999);
or U1093 (N_1093,N_934,N_907);
nand U1094 (N_1094,N_929,N_942);
and U1095 (N_1095,N_991,N_915);
nor U1096 (N_1096,N_977,N_924);
nand U1097 (N_1097,N_995,N_956);
nand U1098 (N_1098,N_943,N_937);
or U1099 (N_1099,N_900,N_942);
and U1100 (N_1100,N_1050,N_1056);
nand U1101 (N_1101,N_1081,N_1070);
nand U1102 (N_1102,N_1064,N_1082);
nand U1103 (N_1103,N_1089,N_1057);
nor U1104 (N_1104,N_1099,N_1069);
and U1105 (N_1105,N_1075,N_1043);
nor U1106 (N_1106,N_1080,N_1087);
nand U1107 (N_1107,N_1053,N_1006);
nor U1108 (N_1108,N_1013,N_1071);
xor U1109 (N_1109,N_1038,N_1059);
nand U1110 (N_1110,N_1046,N_1091);
or U1111 (N_1111,N_1031,N_1044);
or U1112 (N_1112,N_1065,N_1036);
and U1113 (N_1113,N_1033,N_1041);
nand U1114 (N_1114,N_1094,N_1051);
and U1115 (N_1115,N_1020,N_1042);
and U1116 (N_1116,N_1019,N_1001);
nand U1117 (N_1117,N_1025,N_1048);
or U1118 (N_1118,N_1035,N_1030);
or U1119 (N_1119,N_1098,N_1017);
or U1120 (N_1120,N_1068,N_1077);
nand U1121 (N_1121,N_1067,N_1018);
and U1122 (N_1122,N_1037,N_1097);
nand U1123 (N_1123,N_1008,N_1093);
and U1124 (N_1124,N_1049,N_1074);
nor U1125 (N_1125,N_1000,N_1088);
and U1126 (N_1126,N_1021,N_1055);
and U1127 (N_1127,N_1095,N_1007);
and U1128 (N_1128,N_1052,N_1078);
nor U1129 (N_1129,N_1029,N_1066);
nand U1130 (N_1130,N_1015,N_1039);
nor U1131 (N_1131,N_1028,N_1060);
nor U1132 (N_1132,N_1062,N_1061);
and U1133 (N_1133,N_1003,N_1040);
and U1134 (N_1134,N_1090,N_1002);
or U1135 (N_1135,N_1026,N_1073);
or U1136 (N_1136,N_1004,N_1076);
and U1137 (N_1137,N_1010,N_1032);
nand U1138 (N_1138,N_1054,N_1009);
nand U1139 (N_1139,N_1083,N_1027);
nor U1140 (N_1140,N_1024,N_1023);
or U1141 (N_1141,N_1034,N_1016);
or U1142 (N_1142,N_1072,N_1047);
nor U1143 (N_1143,N_1063,N_1086);
or U1144 (N_1144,N_1005,N_1045);
nand U1145 (N_1145,N_1058,N_1084);
and U1146 (N_1146,N_1085,N_1092);
or U1147 (N_1147,N_1096,N_1022);
nor U1148 (N_1148,N_1014,N_1079);
and U1149 (N_1149,N_1012,N_1011);
xor U1150 (N_1150,N_1090,N_1049);
and U1151 (N_1151,N_1046,N_1066);
and U1152 (N_1152,N_1052,N_1047);
xor U1153 (N_1153,N_1099,N_1048);
nor U1154 (N_1154,N_1028,N_1039);
and U1155 (N_1155,N_1051,N_1016);
and U1156 (N_1156,N_1074,N_1075);
nand U1157 (N_1157,N_1054,N_1058);
nor U1158 (N_1158,N_1095,N_1009);
nand U1159 (N_1159,N_1050,N_1055);
nor U1160 (N_1160,N_1016,N_1071);
and U1161 (N_1161,N_1052,N_1009);
nor U1162 (N_1162,N_1021,N_1059);
or U1163 (N_1163,N_1098,N_1039);
nor U1164 (N_1164,N_1036,N_1018);
nand U1165 (N_1165,N_1021,N_1056);
nor U1166 (N_1166,N_1024,N_1066);
and U1167 (N_1167,N_1088,N_1078);
nor U1168 (N_1168,N_1096,N_1042);
and U1169 (N_1169,N_1053,N_1096);
nand U1170 (N_1170,N_1030,N_1069);
nor U1171 (N_1171,N_1075,N_1042);
nor U1172 (N_1172,N_1083,N_1047);
or U1173 (N_1173,N_1008,N_1058);
nand U1174 (N_1174,N_1054,N_1063);
and U1175 (N_1175,N_1037,N_1073);
or U1176 (N_1176,N_1078,N_1063);
and U1177 (N_1177,N_1062,N_1053);
or U1178 (N_1178,N_1097,N_1003);
and U1179 (N_1179,N_1099,N_1020);
or U1180 (N_1180,N_1091,N_1031);
nor U1181 (N_1181,N_1009,N_1094);
or U1182 (N_1182,N_1008,N_1088);
or U1183 (N_1183,N_1015,N_1021);
or U1184 (N_1184,N_1074,N_1085);
and U1185 (N_1185,N_1012,N_1057);
and U1186 (N_1186,N_1027,N_1030);
or U1187 (N_1187,N_1024,N_1011);
nand U1188 (N_1188,N_1049,N_1054);
nand U1189 (N_1189,N_1047,N_1015);
nor U1190 (N_1190,N_1083,N_1017);
nand U1191 (N_1191,N_1071,N_1063);
and U1192 (N_1192,N_1003,N_1096);
nand U1193 (N_1193,N_1013,N_1015);
nor U1194 (N_1194,N_1055,N_1052);
or U1195 (N_1195,N_1016,N_1014);
or U1196 (N_1196,N_1016,N_1038);
xor U1197 (N_1197,N_1090,N_1054);
nor U1198 (N_1198,N_1017,N_1088);
nor U1199 (N_1199,N_1050,N_1047);
or U1200 (N_1200,N_1101,N_1170);
or U1201 (N_1201,N_1109,N_1189);
nand U1202 (N_1202,N_1156,N_1140);
and U1203 (N_1203,N_1118,N_1183);
and U1204 (N_1204,N_1143,N_1163);
nor U1205 (N_1205,N_1146,N_1136);
or U1206 (N_1206,N_1138,N_1115);
nor U1207 (N_1207,N_1158,N_1117);
nand U1208 (N_1208,N_1161,N_1112);
or U1209 (N_1209,N_1131,N_1165);
and U1210 (N_1210,N_1107,N_1178);
xor U1211 (N_1211,N_1121,N_1110);
nand U1212 (N_1212,N_1195,N_1173);
or U1213 (N_1213,N_1194,N_1145);
nor U1214 (N_1214,N_1114,N_1184);
and U1215 (N_1215,N_1197,N_1155);
nor U1216 (N_1216,N_1172,N_1191);
and U1217 (N_1217,N_1151,N_1174);
nor U1218 (N_1218,N_1108,N_1160);
nand U1219 (N_1219,N_1167,N_1182);
nor U1220 (N_1220,N_1148,N_1180);
or U1221 (N_1221,N_1106,N_1120);
nand U1222 (N_1222,N_1141,N_1162);
and U1223 (N_1223,N_1171,N_1147);
and U1224 (N_1224,N_1123,N_1135);
nand U1225 (N_1225,N_1185,N_1164);
and U1226 (N_1226,N_1100,N_1133);
or U1227 (N_1227,N_1157,N_1179);
and U1228 (N_1228,N_1168,N_1103);
nand U1229 (N_1229,N_1127,N_1129);
and U1230 (N_1230,N_1154,N_1113);
nand U1231 (N_1231,N_1105,N_1130);
and U1232 (N_1232,N_1102,N_1111);
or U1233 (N_1233,N_1159,N_1186);
nor U1234 (N_1234,N_1193,N_1119);
or U1235 (N_1235,N_1139,N_1198);
or U1236 (N_1236,N_1192,N_1152);
nand U1237 (N_1237,N_1190,N_1134);
or U1238 (N_1238,N_1128,N_1132);
nand U1239 (N_1239,N_1153,N_1175);
nand U1240 (N_1240,N_1125,N_1187);
nand U1241 (N_1241,N_1181,N_1124);
or U1242 (N_1242,N_1176,N_1169);
nor U1243 (N_1243,N_1116,N_1144);
xor U1244 (N_1244,N_1150,N_1122);
or U1245 (N_1245,N_1126,N_1177);
nor U1246 (N_1246,N_1188,N_1104);
nand U1247 (N_1247,N_1166,N_1149);
nand U1248 (N_1248,N_1142,N_1196);
or U1249 (N_1249,N_1199,N_1137);
and U1250 (N_1250,N_1122,N_1147);
nor U1251 (N_1251,N_1134,N_1109);
nand U1252 (N_1252,N_1164,N_1110);
and U1253 (N_1253,N_1122,N_1180);
or U1254 (N_1254,N_1114,N_1145);
nand U1255 (N_1255,N_1115,N_1155);
nor U1256 (N_1256,N_1165,N_1170);
or U1257 (N_1257,N_1187,N_1184);
and U1258 (N_1258,N_1142,N_1152);
nor U1259 (N_1259,N_1192,N_1125);
and U1260 (N_1260,N_1116,N_1115);
nand U1261 (N_1261,N_1144,N_1102);
or U1262 (N_1262,N_1107,N_1132);
and U1263 (N_1263,N_1178,N_1139);
or U1264 (N_1264,N_1191,N_1105);
and U1265 (N_1265,N_1189,N_1127);
and U1266 (N_1266,N_1143,N_1169);
and U1267 (N_1267,N_1116,N_1176);
nand U1268 (N_1268,N_1125,N_1120);
and U1269 (N_1269,N_1185,N_1116);
or U1270 (N_1270,N_1118,N_1134);
nand U1271 (N_1271,N_1174,N_1187);
nand U1272 (N_1272,N_1130,N_1152);
and U1273 (N_1273,N_1146,N_1188);
and U1274 (N_1274,N_1112,N_1138);
and U1275 (N_1275,N_1152,N_1119);
or U1276 (N_1276,N_1121,N_1107);
nand U1277 (N_1277,N_1102,N_1168);
nand U1278 (N_1278,N_1101,N_1145);
nor U1279 (N_1279,N_1157,N_1106);
or U1280 (N_1280,N_1132,N_1112);
nand U1281 (N_1281,N_1194,N_1118);
and U1282 (N_1282,N_1137,N_1173);
nor U1283 (N_1283,N_1153,N_1108);
or U1284 (N_1284,N_1120,N_1109);
nand U1285 (N_1285,N_1143,N_1147);
and U1286 (N_1286,N_1174,N_1147);
nor U1287 (N_1287,N_1118,N_1190);
nand U1288 (N_1288,N_1190,N_1174);
nor U1289 (N_1289,N_1118,N_1126);
and U1290 (N_1290,N_1112,N_1133);
and U1291 (N_1291,N_1152,N_1151);
or U1292 (N_1292,N_1106,N_1143);
or U1293 (N_1293,N_1157,N_1100);
nand U1294 (N_1294,N_1146,N_1175);
and U1295 (N_1295,N_1181,N_1110);
nand U1296 (N_1296,N_1118,N_1164);
nand U1297 (N_1297,N_1141,N_1176);
nand U1298 (N_1298,N_1132,N_1106);
nand U1299 (N_1299,N_1157,N_1153);
nor U1300 (N_1300,N_1218,N_1298);
nand U1301 (N_1301,N_1205,N_1271);
nand U1302 (N_1302,N_1238,N_1249);
nand U1303 (N_1303,N_1243,N_1242);
nor U1304 (N_1304,N_1288,N_1280);
and U1305 (N_1305,N_1237,N_1241);
nor U1306 (N_1306,N_1297,N_1270);
or U1307 (N_1307,N_1296,N_1290);
nor U1308 (N_1308,N_1299,N_1292);
nand U1309 (N_1309,N_1262,N_1287);
nand U1310 (N_1310,N_1286,N_1226);
nand U1311 (N_1311,N_1223,N_1201);
nor U1312 (N_1312,N_1265,N_1215);
or U1313 (N_1313,N_1213,N_1211);
nor U1314 (N_1314,N_1278,N_1203);
and U1315 (N_1315,N_1207,N_1214);
or U1316 (N_1316,N_1251,N_1247);
or U1317 (N_1317,N_1274,N_1260);
or U1318 (N_1318,N_1222,N_1257);
nor U1319 (N_1319,N_1235,N_1254);
nor U1320 (N_1320,N_1295,N_1277);
or U1321 (N_1321,N_1261,N_1210);
nor U1322 (N_1322,N_1227,N_1220);
or U1323 (N_1323,N_1225,N_1273);
and U1324 (N_1324,N_1276,N_1266);
and U1325 (N_1325,N_1200,N_1232);
or U1326 (N_1326,N_1275,N_1264);
or U1327 (N_1327,N_1252,N_1212);
nor U1328 (N_1328,N_1234,N_1268);
nand U1329 (N_1329,N_1245,N_1248);
nand U1330 (N_1330,N_1263,N_1289);
nor U1331 (N_1331,N_1244,N_1267);
xnor U1332 (N_1332,N_1239,N_1217);
or U1333 (N_1333,N_1202,N_1229);
or U1334 (N_1334,N_1255,N_1284);
nor U1335 (N_1335,N_1253,N_1291);
nand U1336 (N_1336,N_1269,N_1258);
nor U1337 (N_1337,N_1206,N_1208);
or U1338 (N_1338,N_1231,N_1230);
and U1339 (N_1339,N_1221,N_1283);
nand U1340 (N_1340,N_1236,N_1204);
nand U1341 (N_1341,N_1281,N_1279);
or U1342 (N_1342,N_1240,N_1282);
and U1343 (N_1343,N_1209,N_1246);
nor U1344 (N_1344,N_1293,N_1228);
nor U1345 (N_1345,N_1219,N_1256);
and U1346 (N_1346,N_1259,N_1224);
or U1347 (N_1347,N_1272,N_1294);
nand U1348 (N_1348,N_1285,N_1216);
nand U1349 (N_1349,N_1250,N_1233);
nor U1350 (N_1350,N_1219,N_1287);
and U1351 (N_1351,N_1205,N_1228);
nor U1352 (N_1352,N_1290,N_1234);
and U1353 (N_1353,N_1268,N_1202);
nor U1354 (N_1354,N_1210,N_1277);
and U1355 (N_1355,N_1233,N_1226);
nand U1356 (N_1356,N_1294,N_1278);
nand U1357 (N_1357,N_1263,N_1285);
or U1358 (N_1358,N_1298,N_1209);
and U1359 (N_1359,N_1285,N_1269);
nand U1360 (N_1360,N_1226,N_1210);
and U1361 (N_1361,N_1291,N_1234);
nor U1362 (N_1362,N_1232,N_1239);
nand U1363 (N_1363,N_1233,N_1231);
nand U1364 (N_1364,N_1221,N_1226);
and U1365 (N_1365,N_1296,N_1211);
nor U1366 (N_1366,N_1209,N_1263);
nand U1367 (N_1367,N_1243,N_1233);
nand U1368 (N_1368,N_1230,N_1280);
nand U1369 (N_1369,N_1255,N_1259);
nand U1370 (N_1370,N_1270,N_1203);
nor U1371 (N_1371,N_1240,N_1271);
nor U1372 (N_1372,N_1280,N_1258);
or U1373 (N_1373,N_1299,N_1288);
nand U1374 (N_1374,N_1288,N_1215);
nand U1375 (N_1375,N_1291,N_1217);
or U1376 (N_1376,N_1223,N_1262);
or U1377 (N_1377,N_1243,N_1216);
or U1378 (N_1378,N_1214,N_1216);
nand U1379 (N_1379,N_1260,N_1289);
nor U1380 (N_1380,N_1281,N_1248);
and U1381 (N_1381,N_1287,N_1208);
nand U1382 (N_1382,N_1277,N_1261);
or U1383 (N_1383,N_1228,N_1200);
nor U1384 (N_1384,N_1257,N_1273);
and U1385 (N_1385,N_1297,N_1282);
nand U1386 (N_1386,N_1287,N_1227);
or U1387 (N_1387,N_1268,N_1235);
nand U1388 (N_1388,N_1217,N_1247);
or U1389 (N_1389,N_1274,N_1229);
or U1390 (N_1390,N_1202,N_1233);
nor U1391 (N_1391,N_1210,N_1282);
nor U1392 (N_1392,N_1297,N_1265);
nor U1393 (N_1393,N_1293,N_1268);
and U1394 (N_1394,N_1281,N_1267);
nand U1395 (N_1395,N_1264,N_1287);
and U1396 (N_1396,N_1226,N_1252);
and U1397 (N_1397,N_1290,N_1248);
nand U1398 (N_1398,N_1227,N_1266);
xnor U1399 (N_1399,N_1215,N_1282);
nand U1400 (N_1400,N_1326,N_1379);
or U1401 (N_1401,N_1397,N_1360);
and U1402 (N_1402,N_1388,N_1398);
or U1403 (N_1403,N_1315,N_1363);
nor U1404 (N_1404,N_1334,N_1332);
nor U1405 (N_1405,N_1335,N_1338);
nand U1406 (N_1406,N_1304,N_1387);
and U1407 (N_1407,N_1324,N_1323);
and U1408 (N_1408,N_1359,N_1349);
nand U1409 (N_1409,N_1367,N_1317);
nor U1410 (N_1410,N_1394,N_1305);
or U1411 (N_1411,N_1364,N_1318);
nor U1412 (N_1412,N_1376,N_1306);
nand U1413 (N_1413,N_1389,N_1331);
or U1414 (N_1414,N_1330,N_1395);
nor U1415 (N_1415,N_1328,N_1352);
xor U1416 (N_1416,N_1355,N_1390);
nor U1417 (N_1417,N_1372,N_1357);
and U1418 (N_1418,N_1384,N_1346);
nand U1419 (N_1419,N_1343,N_1378);
nand U1420 (N_1420,N_1377,N_1307);
and U1421 (N_1421,N_1391,N_1356);
or U1422 (N_1422,N_1386,N_1353);
and U1423 (N_1423,N_1309,N_1314);
nor U1424 (N_1424,N_1344,N_1383);
or U1425 (N_1425,N_1366,N_1361);
and U1426 (N_1426,N_1347,N_1396);
nor U1427 (N_1427,N_1350,N_1340);
or U1428 (N_1428,N_1333,N_1371);
nand U1429 (N_1429,N_1319,N_1316);
nand U1430 (N_1430,N_1308,N_1385);
or U1431 (N_1431,N_1365,N_1312);
nand U1432 (N_1432,N_1322,N_1339);
and U1433 (N_1433,N_1354,N_1392);
and U1434 (N_1434,N_1348,N_1381);
nor U1435 (N_1435,N_1301,N_1300);
and U1436 (N_1436,N_1337,N_1310);
nor U1437 (N_1437,N_1351,N_1373);
nor U1438 (N_1438,N_1303,N_1342);
or U1439 (N_1439,N_1327,N_1325);
nand U1440 (N_1440,N_1362,N_1341);
and U1441 (N_1441,N_1345,N_1329);
nand U1442 (N_1442,N_1358,N_1370);
and U1443 (N_1443,N_1393,N_1320);
nand U1444 (N_1444,N_1321,N_1369);
and U1445 (N_1445,N_1302,N_1311);
nor U1446 (N_1446,N_1313,N_1375);
nand U1447 (N_1447,N_1336,N_1399);
nand U1448 (N_1448,N_1374,N_1368);
and U1449 (N_1449,N_1380,N_1382);
or U1450 (N_1450,N_1366,N_1387);
and U1451 (N_1451,N_1343,N_1360);
or U1452 (N_1452,N_1388,N_1354);
nor U1453 (N_1453,N_1379,N_1312);
nor U1454 (N_1454,N_1360,N_1310);
xnor U1455 (N_1455,N_1313,N_1343);
or U1456 (N_1456,N_1307,N_1345);
or U1457 (N_1457,N_1381,N_1309);
nand U1458 (N_1458,N_1375,N_1372);
or U1459 (N_1459,N_1313,N_1356);
nand U1460 (N_1460,N_1335,N_1361);
nor U1461 (N_1461,N_1329,N_1321);
and U1462 (N_1462,N_1363,N_1374);
or U1463 (N_1463,N_1325,N_1364);
nor U1464 (N_1464,N_1333,N_1338);
and U1465 (N_1465,N_1320,N_1369);
and U1466 (N_1466,N_1396,N_1365);
nor U1467 (N_1467,N_1379,N_1305);
or U1468 (N_1468,N_1322,N_1337);
or U1469 (N_1469,N_1311,N_1301);
nand U1470 (N_1470,N_1366,N_1362);
nor U1471 (N_1471,N_1316,N_1389);
and U1472 (N_1472,N_1388,N_1393);
or U1473 (N_1473,N_1382,N_1397);
and U1474 (N_1474,N_1326,N_1348);
or U1475 (N_1475,N_1324,N_1359);
or U1476 (N_1476,N_1314,N_1305);
nor U1477 (N_1477,N_1362,N_1391);
nand U1478 (N_1478,N_1359,N_1325);
nand U1479 (N_1479,N_1360,N_1333);
and U1480 (N_1480,N_1389,N_1312);
and U1481 (N_1481,N_1354,N_1398);
or U1482 (N_1482,N_1360,N_1331);
and U1483 (N_1483,N_1346,N_1324);
nor U1484 (N_1484,N_1363,N_1344);
nand U1485 (N_1485,N_1379,N_1331);
or U1486 (N_1486,N_1372,N_1376);
xor U1487 (N_1487,N_1325,N_1382);
nand U1488 (N_1488,N_1381,N_1390);
or U1489 (N_1489,N_1326,N_1355);
and U1490 (N_1490,N_1386,N_1330);
nand U1491 (N_1491,N_1330,N_1358);
nor U1492 (N_1492,N_1361,N_1326);
or U1493 (N_1493,N_1334,N_1392);
and U1494 (N_1494,N_1346,N_1345);
or U1495 (N_1495,N_1332,N_1307);
nand U1496 (N_1496,N_1371,N_1319);
and U1497 (N_1497,N_1333,N_1399);
nand U1498 (N_1498,N_1392,N_1349);
or U1499 (N_1499,N_1398,N_1306);
xor U1500 (N_1500,N_1452,N_1464);
nor U1501 (N_1501,N_1419,N_1402);
and U1502 (N_1502,N_1417,N_1436);
and U1503 (N_1503,N_1423,N_1477);
nor U1504 (N_1504,N_1492,N_1429);
and U1505 (N_1505,N_1406,N_1445);
and U1506 (N_1506,N_1460,N_1446);
nor U1507 (N_1507,N_1471,N_1458);
nand U1508 (N_1508,N_1414,N_1483);
and U1509 (N_1509,N_1495,N_1470);
or U1510 (N_1510,N_1403,N_1461);
and U1511 (N_1511,N_1456,N_1491);
or U1512 (N_1512,N_1444,N_1468);
nand U1513 (N_1513,N_1498,N_1463);
xor U1514 (N_1514,N_1410,N_1476);
or U1515 (N_1515,N_1481,N_1497);
and U1516 (N_1516,N_1494,N_1449);
and U1517 (N_1517,N_1408,N_1424);
and U1518 (N_1518,N_1486,N_1453);
and U1519 (N_1519,N_1465,N_1443);
and U1520 (N_1520,N_1457,N_1489);
or U1521 (N_1521,N_1480,N_1433);
nand U1522 (N_1522,N_1499,N_1473);
nand U1523 (N_1523,N_1451,N_1430);
nand U1524 (N_1524,N_1478,N_1425);
nor U1525 (N_1525,N_1441,N_1455);
xor U1526 (N_1526,N_1438,N_1411);
and U1527 (N_1527,N_1487,N_1422);
and U1528 (N_1528,N_1407,N_1413);
nand U1529 (N_1529,N_1431,N_1467);
and U1530 (N_1530,N_1482,N_1472);
nor U1531 (N_1531,N_1421,N_1475);
or U1532 (N_1532,N_1400,N_1412);
nor U1533 (N_1533,N_1493,N_1488);
nand U1534 (N_1534,N_1466,N_1479);
nor U1535 (N_1535,N_1434,N_1415);
or U1536 (N_1536,N_1416,N_1426);
and U1537 (N_1537,N_1469,N_1428);
and U1538 (N_1538,N_1420,N_1462);
nor U1539 (N_1539,N_1484,N_1437);
nor U1540 (N_1540,N_1450,N_1459);
nand U1541 (N_1541,N_1405,N_1439);
nand U1542 (N_1542,N_1409,N_1442);
or U1543 (N_1543,N_1418,N_1447);
or U1544 (N_1544,N_1474,N_1485);
and U1545 (N_1545,N_1404,N_1496);
nand U1546 (N_1546,N_1432,N_1490);
nor U1547 (N_1547,N_1448,N_1435);
and U1548 (N_1548,N_1427,N_1454);
nand U1549 (N_1549,N_1401,N_1440);
nand U1550 (N_1550,N_1463,N_1452);
nor U1551 (N_1551,N_1492,N_1493);
nor U1552 (N_1552,N_1472,N_1414);
nor U1553 (N_1553,N_1449,N_1466);
nor U1554 (N_1554,N_1425,N_1467);
and U1555 (N_1555,N_1405,N_1444);
nand U1556 (N_1556,N_1432,N_1478);
nor U1557 (N_1557,N_1483,N_1403);
nor U1558 (N_1558,N_1467,N_1448);
nand U1559 (N_1559,N_1442,N_1475);
nor U1560 (N_1560,N_1462,N_1429);
and U1561 (N_1561,N_1459,N_1426);
nor U1562 (N_1562,N_1480,N_1483);
nor U1563 (N_1563,N_1472,N_1473);
or U1564 (N_1564,N_1401,N_1459);
nor U1565 (N_1565,N_1418,N_1485);
or U1566 (N_1566,N_1462,N_1491);
nand U1567 (N_1567,N_1445,N_1405);
nand U1568 (N_1568,N_1487,N_1477);
nor U1569 (N_1569,N_1401,N_1411);
nor U1570 (N_1570,N_1466,N_1475);
and U1571 (N_1571,N_1438,N_1429);
and U1572 (N_1572,N_1446,N_1472);
or U1573 (N_1573,N_1437,N_1428);
nor U1574 (N_1574,N_1499,N_1431);
and U1575 (N_1575,N_1497,N_1462);
nor U1576 (N_1576,N_1449,N_1435);
or U1577 (N_1577,N_1459,N_1491);
and U1578 (N_1578,N_1473,N_1479);
nor U1579 (N_1579,N_1430,N_1429);
and U1580 (N_1580,N_1423,N_1436);
nand U1581 (N_1581,N_1482,N_1443);
and U1582 (N_1582,N_1415,N_1436);
nand U1583 (N_1583,N_1457,N_1428);
nand U1584 (N_1584,N_1497,N_1465);
or U1585 (N_1585,N_1469,N_1445);
nor U1586 (N_1586,N_1444,N_1461);
and U1587 (N_1587,N_1444,N_1472);
nor U1588 (N_1588,N_1430,N_1415);
nor U1589 (N_1589,N_1401,N_1438);
or U1590 (N_1590,N_1435,N_1428);
or U1591 (N_1591,N_1430,N_1499);
nor U1592 (N_1592,N_1400,N_1486);
and U1593 (N_1593,N_1485,N_1489);
nor U1594 (N_1594,N_1477,N_1413);
nor U1595 (N_1595,N_1499,N_1493);
nor U1596 (N_1596,N_1473,N_1454);
and U1597 (N_1597,N_1416,N_1412);
nand U1598 (N_1598,N_1435,N_1476);
nor U1599 (N_1599,N_1459,N_1482);
and U1600 (N_1600,N_1541,N_1554);
nand U1601 (N_1601,N_1537,N_1590);
or U1602 (N_1602,N_1565,N_1539);
nand U1603 (N_1603,N_1517,N_1566);
nand U1604 (N_1604,N_1582,N_1550);
and U1605 (N_1605,N_1536,N_1542);
and U1606 (N_1606,N_1576,N_1543);
or U1607 (N_1607,N_1595,N_1592);
nor U1608 (N_1608,N_1528,N_1545);
nor U1609 (N_1609,N_1533,N_1578);
and U1610 (N_1610,N_1527,N_1549);
nor U1611 (N_1611,N_1519,N_1573);
and U1612 (N_1612,N_1567,N_1521);
and U1613 (N_1613,N_1511,N_1574);
nor U1614 (N_1614,N_1526,N_1596);
nor U1615 (N_1615,N_1583,N_1507);
and U1616 (N_1616,N_1505,N_1531);
nand U1617 (N_1617,N_1564,N_1580);
and U1618 (N_1618,N_1508,N_1561);
and U1619 (N_1619,N_1548,N_1559);
or U1620 (N_1620,N_1597,N_1598);
and U1621 (N_1621,N_1544,N_1589);
nand U1622 (N_1622,N_1570,N_1593);
or U1623 (N_1623,N_1503,N_1551);
nor U1624 (N_1624,N_1553,N_1556);
nand U1625 (N_1625,N_1557,N_1538);
nor U1626 (N_1626,N_1586,N_1555);
nor U1627 (N_1627,N_1585,N_1530);
and U1628 (N_1628,N_1535,N_1568);
and U1629 (N_1629,N_1599,N_1501);
and U1630 (N_1630,N_1504,N_1514);
nor U1631 (N_1631,N_1525,N_1534);
nand U1632 (N_1632,N_1510,N_1513);
or U1633 (N_1633,N_1571,N_1575);
nand U1634 (N_1634,N_1588,N_1552);
or U1635 (N_1635,N_1584,N_1509);
or U1636 (N_1636,N_1562,N_1594);
or U1637 (N_1637,N_1579,N_1506);
and U1638 (N_1638,N_1569,N_1547);
nor U1639 (N_1639,N_1577,N_1523);
nand U1640 (N_1640,N_1512,N_1558);
xor U1641 (N_1641,N_1591,N_1500);
and U1642 (N_1642,N_1560,N_1520);
nor U1643 (N_1643,N_1529,N_1540);
or U1644 (N_1644,N_1516,N_1563);
and U1645 (N_1645,N_1532,N_1502);
nor U1646 (N_1646,N_1572,N_1518);
nand U1647 (N_1647,N_1524,N_1522);
nand U1648 (N_1648,N_1546,N_1515);
or U1649 (N_1649,N_1587,N_1581);
and U1650 (N_1650,N_1552,N_1510);
and U1651 (N_1651,N_1511,N_1582);
and U1652 (N_1652,N_1501,N_1552);
nor U1653 (N_1653,N_1547,N_1571);
or U1654 (N_1654,N_1570,N_1571);
or U1655 (N_1655,N_1585,N_1529);
or U1656 (N_1656,N_1538,N_1533);
or U1657 (N_1657,N_1564,N_1535);
or U1658 (N_1658,N_1593,N_1576);
or U1659 (N_1659,N_1592,N_1593);
nand U1660 (N_1660,N_1586,N_1578);
nand U1661 (N_1661,N_1567,N_1518);
nand U1662 (N_1662,N_1582,N_1563);
nor U1663 (N_1663,N_1538,N_1572);
nor U1664 (N_1664,N_1558,N_1565);
or U1665 (N_1665,N_1537,N_1572);
and U1666 (N_1666,N_1525,N_1569);
or U1667 (N_1667,N_1588,N_1526);
or U1668 (N_1668,N_1591,N_1551);
or U1669 (N_1669,N_1554,N_1543);
nor U1670 (N_1670,N_1500,N_1565);
nor U1671 (N_1671,N_1549,N_1560);
nor U1672 (N_1672,N_1541,N_1528);
and U1673 (N_1673,N_1561,N_1575);
nor U1674 (N_1674,N_1511,N_1591);
or U1675 (N_1675,N_1597,N_1534);
nand U1676 (N_1676,N_1508,N_1596);
nor U1677 (N_1677,N_1518,N_1587);
or U1678 (N_1678,N_1500,N_1588);
nand U1679 (N_1679,N_1570,N_1582);
and U1680 (N_1680,N_1566,N_1584);
nor U1681 (N_1681,N_1542,N_1510);
nor U1682 (N_1682,N_1540,N_1523);
nand U1683 (N_1683,N_1540,N_1513);
nand U1684 (N_1684,N_1579,N_1574);
and U1685 (N_1685,N_1572,N_1540);
nor U1686 (N_1686,N_1540,N_1552);
and U1687 (N_1687,N_1583,N_1513);
nand U1688 (N_1688,N_1555,N_1563);
nor U1689 (N_1689,N_1514,N_1541);
or U1690 (N_1690,N_1525,N_1522);
nor U1691 (N_1691,N_1561,N_1584);
and U1692 (N_1692,N_1588,N_1555);
and U1693 (N_1693,N_1560,N_1559);
or U1694 (N_1694,N_1576,N_1567);
nand U1695 (N_1695,N_1530,N_1538);
or U1696 (N_1696,N_1544,N_1586);
nand U1697 (N_1697,N_1576,N_1573);
nor U1698 (N_1698,N_1580,N_1543);
and U1699 (N_1699,N_1538,N_1587);
and U1700 (N_1700,N_1687,N_1603);
or U1701 (N_1701,N_1620,N_1608);
and U1702 (N_1702,N_1607,N_1669);
nor U1703 (N_1703,N_1695,N_1623);
and U1704 (N_1704,N_1678,N_1641);
and U1705 (N_1705,N_1664,N_1629);
or U1706 (N_1706,N_1665,N_1652);
or U1707 (N_1707,N_1612,N_1691);
or U1708 (N_1708,N_1628,N_1675);
and U1709 (N_1709,N_1610,N_1674);
and U1710 (N_1710,N_1686,N_1626);
or U1711 (N_1711,N_1654,N_1621);
and U1712 (N_1712,N_1643,N_1637);
or U1713 (N_1713,N_1625,N_1653);
nor U1714 (N_1714,N_1684,N_1648);
nand U1715 (N_1715,N_1646,N_1659);
nand U1716 (N_1716,N_1639,N_1614);
nand U1717 (N_1717,N_1672,N_1658);
nand U1718 (N_1718,N_1615,N_1655);
and U1719 (N_1719,N_1613,N_1680);
and U1720 (N_1720,N_1677,N_1651);
nand U1721 (N_1721,N_1668,N_1688);
and U1722 (N_1722,N_1698,N_1609);
and U1723 (N_1723,N_1671,N_1667);
or U1724 (N_1724,N_1640,N_1605);
nand U1725 (N_1725,N_1673,N_1624);
or U1726 (N_1726,N_1638,N_1611);
nor U1727 (N_1727,N_1622,N_1645);
nor U1728 (N_1728,N_1616,N_1685);
nor U1729 (N_1729,N_1602,N_1617);
or U1730 (N_1730,N_1660,N_1632);
or U1731 (N_1731,N_1636,N_1689);
and U1732 (N_1732,N_1618,N_1662);
nor U1733 (N_1733,N_1690,N_1681);
nand U1734 (N_1734,N_1642,N_1649);
and U1735 (N_1735,N_1627,N_1661);
or U1736 (N_1736,N_1699,N_1683);
or U1737 (N_1737,N_1657,N_1631);
nand U1738 (N_1738,N_1663,N_1604);
or U1739 (N_1739,N_1666,N_1682);
and U1740 (N_1740,N_1676,N_1633);
nand U1741 (N_1741,N_1693,N_1644);
and U1742 (N_1742,N_1670,N_1606);
nor U1743 (N_1743,N_1650,N_1679);
and U1744 (N_1744,N_1697,N_1634);
and U1745 (N_1745,N_1635,N_1692);
and U1746 (N_1746,N_1656,N_1630);
or U1747 (N_1747,N_1600,N_1696);
nand U1748 (N_1748,N_1647,N_1619);
nor U1749 (N_1749,N_1601,N_1694);
nor U1750 (N_1750,N_1616,N_1617);
and U1751 (N_1751,N_1683,N_1678);
nor U1752 (N_1752,N_1665,N_1677);
nand U1753 (N_1753,N_1658,N_1623);
and U1754 (N_1754,N_1682,N_1684);
or U1755 (N_1755,N_1682,N_1618);
nor U1756 (N_1756,N_1680,N_1655);
or U1757 (N_1757,N_1683,N_1607);
or U1758 (N_1758,N_1658,N_1699);
nand U1759 (N_1759,N_1697,N_1635);
nor U1760 (N_1760,N_1692,N_1647);
or U1761 (N_1761,N_1610,N_1600);
xnor U1762 (N_1762,N_1667,N_1657);
nand U1763 (N_1763,N_1653,N_1692);
or U1764 (N_1764,N_1615,N_1694);
nand U1765 (N_1765,N_1660,N_1669);
or U1766 (N_1766,N_1666,N_1686);
nor U1767 (N_1767,N_1648,N_1680);
nor U1768 (N_1768,N_1607,N_1608);
nor U1769 (N_1769,N_1653,N_1684);
and U1770 (N_1770,N_1633,N_1638);
nor U1771 (N_1771,N_1629,N_1625);
nand U1772 (N_1772,N_1661,N_1637);
or U1773 (N_1773,N_1698,N_1606);
and U1774 (N_1774,N_1651,N_1673);
and U1775 (N_1775,N_1641,N_1645);
and U1776 (N_1776,N_1644,N_1623);
and U1777 (N_1777,N_1666,N_1659);
nor U1778 (N_1778,N_1640,N_1660);
and U1779 (N_1779,N_1676,N_1667);
xnor U1780 (N_1780,N_1634,N_1684);
nand U1781 (N_1781,N_1655,N_1634);
and U1782 (N_1782,N_1629,N_1658);
and U1783 (N_1783,N_1637,N_1669);
nand U1784 (N_1784,N_1651,N_1668);
nor U1785 (N_1785,N_1691,N_1633);
nor U1786 (N_1786,N_1670,N_1688);
and U1787 (N_1787,N_1699,N_1647);
and U1788 (N_1788,N_1621,N_1677);
or U1789 (N_1789,N_1612,N_1629);
nand U1790 (N_1790,N_1633,N_1668);
nand U1791 (N_1791,N_1690,N_1607);
nor U1792 (N_1792,N_1694,N_1661);
or U1793 (N_1793,N_1642,N_1680);
nand U1794 (N_1794,N_1642,N_1670);
or U1795 (N_1795,N_1676,N_1650);
nor U1796 (N_1796,N_1636,N_1653);
or U1797 (N_1797,N_1606,N_1680);
nand U1798 (N_1798,N_1647,N_1673);
or U1799 (N_1799,N_1674,N_1697);
nor U1800 (N_1800,N_1725,N_1799);
or U1801 (N_1801,N_1778,N_1740);
and U1802 (N_1802,N_1772,N_1730);
or U1803 (N_1803,N_1733,N_1751);
nand U1804 (N_1804,N_1704,N_1794);
and U1805 (N_1805,N_1705,N_1708);
nor U1806 (N_1806,N_1786,N_1746);
nand U1807 (N_1807,N_1793,N_1780);
nand U1808 (N_1808,N_1701,N_1707);
nor U1809 (N_1809,N_1756,N_1729);
or U1810 (N_1810,N_1703,N_1763);
and U1811 (N_1811,N_1713,N_1728);
nand U1812 (N_1812,N_1770,N_1727);
or U1813 (N_1813,N_1735,N_1732);
or U1814 (N_1814,N_1744,N_1773);
or U1815 (N_1815,N_1795,N_1742);
and U1816 (N_1816,N_1789,N_1741);
nand U1817 (N_1817,N_1785,N_1757);
and U1818 (N_1818,N_1711,N_1783);
and U1819 (N_1819,N_1720,N_1726);
or U1820 (N_1820,N_1712,N_1747);
or U1821 (N_1821,N_1760,N_1767);
nand U1822 (N_1822,N_1798,N_1700);
nor U1823 (N_1823,N_1796,N_1759);
nand U1824 (N_1824,N_1771,N_1758);
nand U1825 (N_1825,N_1775,N_1749);
nand U1826 (N_1826,N_1748,N_1736);
nand U1827 (N_1827,N_1710,N_1754);
nor U1828 (N_1828,N_1716,N_1734);
nor U1829 (N_1829,N_1739,N_1709);
nand U1830 (N_1830,N_1722,N_1765);
and U1831 (N_1831,N_1718,N_1762);
or U1832 (N_1832,N_1787,N_1715);
or U1833 (N_1833,N_1750,N_1768);
and U1834 (N_1834,N_1792,N_1790);
or U1835 (N_1835,N_1714,N_1788);
and U1836 (N_1836,N_1743,N_1784);
nand U1837 (N_1837,N_1702,N_1781);
nor U1838 (N_1838,N_1717,N_1761);
nor U1839 (N_1839,N_1755,N_1721);
nand U1840 (N_1840,N_1753,N_1777);
nor U1841 (N_1841,N_1791,N_1766);
nand U1842 (N_1842,N_1724,N_1752);
or U1843 (N_1843,N_1706,N_1776);
nand U1844 (N_1844,N_1731,N_1774);
nor U1845 (N_1845,N_1723,N_1745);
or U1846 (N_1846,N_1719,N_1769);
or U1847 (N_1847,N_1764,N_1737);
nor U1848 (N_1848,N_1779,N_1782);
nand U1849 (N_1849,N_1738,N_1797);
or U1850 (N_1850,N_1781,N_1761);
nand U1851 (N_1851,N_1769,N_1799);
and U1852 (N_1852,N_1761,N_1723);
or U1853 (N_1853,N_1786,N_1771);
nand U1854 (N_1854,N_1745,N_1773);
nor U1855 (N_1855,N_1703,N_1700);
xor U1856 (N_1856,N_1733,N_1784);
or U1857 (N_1857,N_1782,N_1737);
and U1858 (N_1858,N_1736,N_1753);
nor U1859 (N_1859,N_1773,N_1777);
nand U1860 (N_1860,N_1714,N_1728);
and U1861 (N_1861,N_1713,N_1704);
and U1862 (N_1862,N_1715,N_1781);
nand U1863 (N_1863,N_1798,N_1746);
nor U1864 (N_1864,N_1771,N_1773);
nor U1865 (N_1865,N_1720,N_1777);
xor U1866 (N_1866,N_1729,N_1797);
nor U1867 (N_1867,N_1710,N_1703);
and U1868 (N_1868,N_1771,N_1792);
and U1869 (N_1869,N_1781,N_1756);
or U1870 (N_1870,N_1705,N_1784);
nor U1871 (N_1871,N_1763,N_1752);
nand U1872 (N_1872,N_1784,N_1701);
and U1873 (N_1873,N_1778,N_1718);
or U1874 (N_1874,N_1783,N_1706);
nor U1875 (N_1875,N_1745,N_1786);
or U1876 (N_1876,N_1799,N_1781);
xor U1877 (N_1877,N_1763,N_1789);
nor U1878 (N_1878,N_1751,N_1718);
and U1879 (N_1879,N_1796,N_1782);
or U1880 (N_1880,N_1760,N_1708);
nand U1881 (N_1881,N_1735,N_1704);
nand U1882 (N_1882,N_1742,N_1728);
nand U1883 (N_1883,N_1761,N_1703);
nor U1884 (N_1884,N_1730,N_1702);
and U1885 (N_1885,N_1754,N_1748);
nor U1886 (N_1886,N_1786,N_1710);
nand U1887 (N_1887,N_1758,N_1766);
nand U1888 (N_1888,N_1792,N_1732);
nor U1889 (N_1889,N_1790,N_1779);
and U1890 (N_1890,N_1707,N_1745);
nand U1891 (N_1891,N_1781,N_1748);
and U1892 (N_1892,N_1769,N_1789);
or U1893 (N_1893,N_1797,N_1712);
or U1894 (N_1894,N_1735,N_1777);
nor U1895 (N_1895,N_1795,N_1774);
or U1896 (N_1896,N_1790,N_1708);
nand U1897 (N_1897,N_1729,N_1763);
and U1898 (N_1898,N_1725,N_1765);
nand U1899 (N_1899,N_1750,N_1767);
and U1900 (N_1900,N_1876,N_1880);
and U1901 (N_1901,N_1825,N_1870);
nand U1902 (N_1902,N_1815,N_1821);
nand U1903 (N_1903,N_1841,N_1893);
and U1904 (N_1904,N_1805,N_1831);
nand U1905 (N_1905,N_1863,N_1859);
or U1906 (N_1906,N_1864,N_1819);
and U1907 (N_1907,N_1830,N_1809);
nand U1908 (N_1908,N_1873,N_1872);
or U1909 (N_1909,N_1894,N_1834);
and U1910 (N_1910,N_1806,N_1802);
nand U1911 (N_1911,N_1898,N_1858);
nand U1912 (N_1912,N_1823,N_1807);
nor U1913 (N_1913,N_1824,N_1854);
nor U1914 (N_1914,N_1849,N_1818);
nand U1915 (N_1915,N_1888,N_1857);
nand U1916 (N_1916,N_1867,N_1833);
or U1917 (N_1917,N_1839,N_1878);
nand U1918 (N_1918,N_1843,N_1853);
xor U1919 (N_1919,N_1856,N_1822);
or U1920 (N_1920,N_1847,N_1861);
and U1921 (N_1921,N_1842,N_1848);
nand U1922 (N_1922,N_1879,N_1899);
nor U1923 (N_1923,N_1845,N_1886);
or U1924 (N_1924,N_1816,N_1866);
nor U1925 (N_1925,N_1891,N_1826);
nor U1926 (N_1926,N_1812,N_1874);
or U1927 (N_1927,N_1828,N_1883);
nor U1928 (N_1928,N_1875,N_1832);
nand U1929 (N_1929,N_1810,N_1836);
nand U1930 (N_1930,N_1868,N_1887);
xnor U1931 (N_1931,N_1895,N_1877);
or U1932 (N_1932,N_1814,N_1840);
and U1933 (N_1933,N_1800,N_1889);
or U1934 (N_1934,N_1844,N_1801);
and U1935 (N_1935,N_1852,N_1871);
nand U1936 (N_1936,N_1808,N_1855);
nand U1937 (N_1937,N_1862,N_1850);
nor U1938 (N_1938,N_1851,N_1890);
nor U1939 (N_1939,N_1838,N_1835);
or U1940 (N_1940,N_1881,N_1817);
or U1941 (N_1941,N_1820,N_1896);
nor U1942 (N_1942,N_1897,N_1882);
and U1943 (N_1943,N_1865,N_1827);
nor U1944 (N_1944,N_1813,N_1804);
and U1945 (N_1945,N_1811,N_1885);
nand U1946 (N_1946,N_1837,N_1829);
and U1947 (N_1947,N_1846,N_1803);
nor U1948 (N_1948,N_1884,N_1860);
and U1949 (N_1949,N_1892,N_1869);
nor U1950 (N_1950,N_1879,N_1855);
and U1951 (N_1951,N_1809,N_1850);
and U1952 (N_1952,N_1871,N_1813);
and U1953 (N_1953,N_1826,N_1854);
nand U1954 (N_1954,N_1870,N_1887);
nor U1955 (N_1955,N_1856,N_1843);
nand U1956 (N_1956,N_1869,N_1854);
or U1957 (N_1957,N_1851,N_1879);
or U1958 (N_1958,N_1844,N_1824);
or U1959 (N_1959,N_1803,N_1867);
and U1960 (N_1960,N_1895,N_1800);
or U1961 (N_1961,N_1826,N_1804);
and U1962 (N_1962,N_1885,N_1891);
or U1963 (N_1963,N_1879,N_1807);
nand U1964 (N_1964,N_1831,N_1852);
nand U1965 (N_1965,N_1874,N_1816);
and U1966 (N_1966,N_1836,N_1805);
nand U1967 (N_1967,N_1819,N_1841);
and U1968 (N_1968,N_1830,N_1870);
nor U1969 (N_1969,N_1832,N_1889);
nand U1970 (N_1970,N_1849,N_1868);
nand U1971 (N_1971,N_1894,N_1800);
and U1972 (N_1972,N_1855,N_1824);
or U1973 (N_1973,N_1848,N_1874);
or U1974 (N_1974,N_1849,N_1844);
nor U1975 (N_1975,N_1899,N_1819);
or U1976 (N_1976,N_1802,N_1805);
nand U1977 (N_1977,N_1859,N_1846);
and U1978 (N_1978,N_1840,N_1856);
nand U1979 (N_1979,N_1887,N_1897);
or U1980 (N_1980,N_1828,N_1841);
nand U1981 (N_1981,N_1886,N_1879);
nand U1982 (N_1982,N_1825,N_1816);
nand U1983 (N_1983,N_1898,N_1846);
and U1984 (N_1984,N_1888,N_1881);
or U1985 (N_1985,N_1839,N_1884);
and U1986 (N_1986,N_1853,N_1875);
and U1987 (N_1987,N_1898,N_1897);
or U1988 (N_1988,N_1898,N_1879);
and U1989 (N_1989,N_1827,N_1806);
and U1990 (N_1990,N_1840,N_1891);
or U1991 (N_1991,N_1820,N_1859);
nand U1992 (N_1992,N_1898,N_1893);
and U1993 (N_1993,N_1841,N_1818);
nand U1994 (N_1994,N_1810,N_1847);
nand U1995 (N_1995,N_1857,N_1877);
nand U1996 (N_1996,N_1822,N_1877);
and U1997 (N_1997,N_1899,N_1810);
and U1998 (N_1998,N_1826,N_1869);
and U1999 (N_1999,N_1820,N_1854);
nand U2000 (N_2000,N_1912,N_1913);
or U2001 (N_2001,N_1981,N_1973);
and U2002 (N_2002,N_1933,N_1970);
nor U2003 (N_2003,N_1958,N_1949);
nor U2004 (N_2004,N_1979,N_1965);
or U2005 (N_2005,N_1935,N_1961);
nand U2006 (N_2006,N_1975,N_1922);
nor U2007 (N_2007,N_1944,N_1989);
nor U2008 (N_2008,N_1992,N_1903);
nand U2009 (N_2009,N_1996,N_1959);
nor U2010 (N_2010,N_1955,N_1960);
and U2011 (N_2011,N_1914,N_1938);
nand U2012 (N_2012,N_1969,N_1948);
or U2013 (N_2013,N_1939,N_1937);
or U2014 (N_2014,N_1962,N_1985);
nand U2015 (N_2015,N_1916,N_1910);
nor U2016 (N_2016,N_1905,N_1921);
or U2017 (N_2017,N_1982,N_1964);
nor U2018 (N_2018,N_1940,N_1942);
and U2019 (N_2019,N_1993,N_1909);
nand U2020 (N_2020,N_1930,N_1947);
or U2021 (N_2021,N_1978,N_1915);
nor U2022 (N_2022,N_1929,N_1932);
nor U2023 (N_2023,N_1974,N_1972);
or U2024 (N_2024,N_1934,N_1963);
or U2025 (N_2025,N_1984,N_1980);
and U2026 (N_2026,N_1906,N_1917);
and U2027 (N_2027,N_1951,N_1950);
or U2028 (N_2028,N_1995,N_1904);
and U2029 (N_2029,N_1987,N_1956);
or U2030 (N_2030,N_1911,N_1908);
nand U2031 (N_2031,N_1900,N_1943);
and U2032 (N_2032,N_1928,N_1953);
nand U2033 (N_2033,N_1983,N_1977);
and U2034 (N_2034,N_1924,N_1954);
nand U2035 (N_2035,N_1901,N_1946);
nor U2036 (N_2036,N_1976,N_1991);
nand U2037 (N_2037,N_1999,N_1988);
or U2038 (N_2038,N_1941,N_1936);
nor U2039 (N_2039,N_1907,N_1902);
nor U2040 (N_2040,N_1967,N_1931);
or U2041 (N_2041,N_1986,N_1920);
nand U2042 (N_2042,N_1968,N_1966);
nand U2043 (N_2043,N_1952,N_1925);
nand U2044 (N_2044,N_1997,N_1971);
or U2045 (N_2045,N_1919,N_1957);
nor U2046 (N_2046,N_1927,N_1918);
nor U2047 (N_2047,N_1994,N_1990);
or U2048 (N_2048,N_1998,N_1945);
or U2049 (N_2049,N_1923,N_1926);
nand U2050 (N_2050,N_1960,N_1928);
or U2051 (N_2051,N_1940,N_1929);
nor U2052 (N_2052,N_1947,N_1942);
nand U2053 (N_2053,N_1997,N_1916);
and U2054 (N_2054,N_1994,N_1991);
nand U2055 (N_2055,N_1958,N_1953);
nand U2056 (N_2056,N_1990,N_1918);
nand U2057 (N_2057,N_1968,N_1919);
or U2058 (N_2058,N_1949,N_1925);
nor U2059 (N_2059,N_1989,N_1953);
nand U2060 (N_2060,N_1985,N_1957);
nand U2061 (N_2061,N_1936,N_1969);
nor U2062 (N_2062,N_1930,N_1926);
nand U2063 (N_2063,N_1989,N_1938);
or U2064 (N_2064,N_1963,N_1973);
and U2065 (N_2065,N_1928,N_1921);
nor U2066 (N_2066,N_1920,N_1933);
or U2067 (N_2067,N_1950,N_1967);
or U2068 (N_2068,N_1970,N_1924);
or U2069 (N_2069,N_1962,N_1945);
or U2070 (N_2070,N_1925,N_1960);
nand U2071 (N_2071,N_1924,N_1965);
and U2072 (N_2072,N_1929,N_1972);
nand U2073 (N_2073,N_1969,N_1981);
nand U2074 (N_2074,N_1950,N_1997);
or U2075 (N_2075,N_1924,N_1972);
and U2076 (N_2076,N_1961,N_1937);
or U2077 (N_2077,N_1989,N_1946);
or U2078 (N_2078,N_1951,N_1945);
nor U2079 (N_2079,N_1905,N_1955);
nand U2080 (N_2080,N_1956,N_1989);
nand U2081 (N_2081,N_1996,N_1925);
or U2082 (N_2082,N_1918,N_1940);
or U2083 (N_2083,N_1931,N_1957);
nand U2084 (N_2084,N_1936,N_1904);
nand U2085 (N_2085,N_1903,N_1955);
and U2086 (N_2086,N_1953,N_1941);
nor U2087 (N_2087,N_1903,N_1913);
or U2088 (N_2088,N_1945,N_1982);
nor U2089 (N_2089,N_1930,N_1932);
nor U2090 (N_2090,N_1931,N_1908);
nor U2091 (N_2091,N_1991,N_1963);
or U2092 (N_2092,N_1933,N_1967);
or U2093 (N_2093,N_1924,N_1919);
nand U2094 (N_2094,N_1971,N_1958);
and U2095 (N_2095,N_1917,N_1963);
nor U2096 (N_2096,N_1900,N_1985);
and U2097 (N_2097,N_1993,N_1912);
or U2098 (N_2098,N_1995,N_1933);
and U2099 (N_2099,N_1999,N_1930);
nand U2100 (N_2100,N_2089,N_2095);
or U2101 (N_2101,N_2075,N_2011);
or U2102 (N_2102,N_2077,N_2078);
nor U2103 (N_2103,N_2072,N_2039);
and U2104 (N_2104,N_2027,N_2037);
or U2105 (N_2105,N_2038,N_2002);
nand U2106 (N_2106,N_2015,N_2003);
nand U2107 (N_2107,N_2099,N_2036);
nand U2108 (N_2108,N_2093,N_2045);
nor U2109 (N_2109,N_2049,N_2005);
nand U2110 (N_2110,N_2087,N_2001);
nand U2111 (N_2111,N_2030,N_2061);
nand U2112 (N_2112,N_2041,N_2048);
or U2113 (N_2113,N_2079,N_2014);
nor U2114 (N_2114,N_2084,N_2024);
or U2115 (N_2115,N_2050,N_2017);
or U2116 (N_2116,N_2035,N_2032);
and U2117 (N_2117,N_2028,N_2047);
or U2118 (N_2118,N_2069,N_2068);
nand U2119 (N_2119,N_2085,N_2090);
and U2120 (N_2120,N_2009,N_2031);
nor U2121 (N_2121,N_2096,N_2056);
and U2122 (N_2122,N_2006,N_2062);
nor U2123 (N_2123,N_2033,N_2071);
nand U2124 (N_2124,N_2020,N_2074);
or U2125 (N_2125,N_2019,N_2063);
and U2126 (N_2126,N_2064,N_2081);
nor U2127 (N_2127,N_2043,N_2023);
nand U2128 (N_2128,N_2066,N_2052);
nand U2129 (N_2129,N_2029,N_2004);
or U2130 (N_2130,N_2057,N_2091);
or U2131 (N_2131,N_2007,N_2067);
nand U2132 (N_2132,N_2016,N_2051);
and U2133 (N_2133,N_2018,N_2055);
nor U2134 (N_2134,N_2026,N_2021);
nand U2135 (N_2135,N_2012,N_2080);
nor U2136 (N_2136,N_2076,N_2073);
nor U2137 (N_2137,N_2059,N_2098);
nor U2138 (N_2138,N_2058,N_2082);
nor U2139 (N_2139,N_2046,N_2065);
nand U2140 (N_2140,N_2097,N_2088);
nand U2141 (N_2141,N_2010,N_2086);
nor U2142 (N_2142,N_2042,N_2060);
or U2143 (N_2143,N_2070,N_2040);
nand U2144 (N_2144,N_2054,N_2094);
or U2145 (N_2145,N_2044,N_2013);
or U2146 (N_2146,N_2022,N_2000);
or U2147 (N_2147,N_2008,N_2034);
nand U2148 (N_2148,N_2053,N_2083);
nor U2149 (N_2149,N_2092,N_2025);
and U2150 (N_2150,N_2049,N_2010);
nor U2151 (N_2151,N_2065,N_2086);
and U2152 (N_2152,N_2000,N_2050);
and U2153 (N_2153,N_2022,N_2035);
nor U2154 (N_2154,N_2021,N_2082);
and U2155 (N_2155,N_2032,N_2008);
or U2156 (N_2156,N_2033,N_2031);
or U2157 (N_2157,N_2040,N_2071);
nand U2158 (N_2158,N_2073,N_2080);
or U2159 (N_2159,N_2051,N_2031);
and U2160 (N_2160,N_2095,N_2070);
or U2161 (N_2161,N_2010,N_2027);
and U2162 (N_2162,N_2035,N_2052);
nand U2163 (N_2163,N_2097,N_2004);
nor U2164 (N_2164,N_2038,N_2039);
nand U2165 (N_2165,N_2097,N_2030);
or U2166 (N_2166,N_2099,N_2009);
or U2167 (N_2167,N_2065,N_2067);
nand U2168 (N_2168,N_2013,N_2070);
nand U2169 (N_2169,N_2026,N_2017);
or U2170 (N_2170,N_2042,N_2097);
nor U2171 (N_2171,N_2047,N_2097);
xnor U2172 (N_2172,N_2036,N_2018);
nor U2173 (N_2173,N_2031,N_2021);
and U2174 (N_2174,N_2027,N_2013);
xnor U2175 (N_2175,N_2079,N_2097);
nand U2176 (N_2176,N_2005,N_2045);
nand U2177 (N_2177,N_2021,N_2058);
and U2178 (N_2178,N_2072,N_2057);
or U2179 (N_2179,N_2051,N_2022);
nor U2180 (N_2180,N_2048,N_2023);
and U2181 (N_2181,N_2072,N_2007);
and U2182 (N_2182,N_2083,N_2021);
nor U2183 (N_2183,N_2004,N_2037);
or U2184 (N_2184,N_2082,N_2077);
nand U2185 (N_2185,N_2020,N_2062);
nor U2186 (N_2186,N_2027,N_2057);
nand U2187 (N_2187,N_2084,N_2052);
nand U2188 (N_2188,N_2006,N_2001);
xor U2189 (N_2189,N_2076,N_2018);
nand U2190 (N_2190,N_2083,N_2060);
nor U2191 (N_2191,N_2054,N_2012);
or U2192 (N_2192,N_2048,N_2042);
nand U2193 (N_2193,N_2068,N_2080);
nand U2194 (N_2194,N_2043,N_2002);
nand U2195 (N_2195,N_2078,N_2015);
and U2196 (N_2196,N_2008,N_2035);
nor U2197 (N_2197,N_2089,N_2007);
nand U2198 (N_2198,N_2020,N_2071);
nand U2199 (N_2199,N_2025,N_2070);
nor U2200 (N_2200,N_2142,N_2135);
nand U2201 (N_2201,N_2121,N_2187);
and U2202 (N_2202,N_2183,N_2157);
nor U2203 (N_2203,N_2151,N_2160);
nand U2204 (N_2204,N_2193,N_2106);
or U2205 (N_2205,N_2171,N_2158);
nor U2206 (N_2206,N_2130,N_2108);
or U2207 (N_2207,N_2148,N_2143);
nand U2208 (N_2208,N_2116,N_2194);
nand U2209 (N_2209,N_2112,N_2118);
nand U2210 (N_2210,N_2185,N_2196);
or U2211 (N_2211,N_2154,N_2111);
and U2212 (N_2212,N_2107,N_2129);
nor U2213 (N_2213,N_2180,N_2133);
and U2214 (N_2214,N_2140,N_2139);
nand U2215 (N_2215,N_2166,N_2147);
or U2216 (N_2216,N_2136,N_2198);
nor U2217 (N_2217,N_2181,N_2150);
or U2218 (N_2218,N_2131,N_2105);
or U2219 (N_2219,N_2192,N_2120);
and U2220 (N_2220,N_2167,N_2109);
nand U2221 (N_2221,N_2146,N_2123);
nor U2222 (N_2222,N_2101,N_2156);
or U2223 (N_2223,N_2162,N_2134);
nor U2224 (N_2224,N_2110,N_2102);
and U2225 (N_2225,N_2168,N_2104);
or U2226 (N_2226,N_2179,N_2159);
nor U2227 (N_2227,N_2172,N_2141);
nand U2228 (N_2228,N_2182,N_2144);
nor U2229 (N_2229,N_2176,N_2175);
and U2230 (N_2230,N_2170,N_2197);
and U2231 (N_2231,N_2184,N_2100);
or U2232 (N_2232,N_2155,N_2149);
nor U2233 (N_2233,N_2164,N_2145);
and U2234 (N_2234,N_2169,N_2103);
and U2235 (N_2235,N_2152,N_2137);
nand U2236 (N_2236,N_2174,N_2161);
and U2237 (N_2237,N_2119,N_2128);
or U2238 (N_2238,N_2165,N_2199);
and U2239 (N_2239,N_2124,N_2178);
nor U2240 (N_2240,N_2125,N_2191);
or U2241 (N_2241,N_2195,N_2138);
nand U2242 (N_2242,N_2127,N_2117);
nor U2243 (N_2243,N_2177,N_2114);
and U2244 (N_2244,N_2115,N_2126);
nand U2245 (N_2245,N_2188,N_2163);
and U2246 (N_2246,N_2190,N_2153);
or U2247 (N_2247,N_2122,N_2173);
or U2248 (N_2248,N_2113,N_2189);
and U2249 (N_2249,N_2186,N_2132);
nand U2250 (N_2250,N_2189,N_2194);
or U2251 (N_2251,N_2195,N_2116);
or U2252 (N_2252,N_2129,N_2119);
and U2253 (N_2253,N_2169,N_2111);
nand U2254 (N_2254,N_2118,N_2117);
nor U2255 (N_2255,N_2142,N_2106);
or U2256 (N_2256,N_2155,N_2144);
and U2257 (N_2257,N_2113,N_2148);
nand U2258 (N_2258,N_2178,N_2159);
or U2259 (N_2259,N_2196,N_2152);
nor U2260 (N_2260,N_2130,N_2188);
nand U2261 (N_2261,N_2181,N_2109);
nor U2262 (N_2262,N_2144,N_2166);
and U2263 (N_2263,N_2144,N_2124);
or U2264 (N_2264,N_2144,N_2112);
or U2265 (N_2265,N_2139,N_2132);
nor U2266 (N_2266,N_2174,N_2149);
xor U2267 (N_2267,N_2160,N_2169);
or U2268 (N_2268,N_2101,N_2152);
nand U2269 (N_2269,N_2169,N_2142);
and U2270 (N_2270,N_2103,N_2129);
and U2271 (N_2271,N_2116,N_2146);
or U2272 (N_2272,N_2145,N_2140);
nand U2273 (N_2273,N_2170,N_2135);
nand U2274 (N_2274,N_2187,N_2102);
nor U2275 (N_2275,N_2143,N_2171);
nor U2276 (N_2276,N_2125,N_2188);
nor U2277 (N_2277,N_2134,N_2126);
nor U2278 (N_2278,N_2170,N_2186);
xor U2279 (N_2279,N_2185,N_2107);
nor U2280 (N_2280,N_2167,N_2153);
nand U2281 (N_2281,N_2166,N_2181);
and U2282 (N_2282,N_2103,N_2136);
nor U2283 (N_2283,N_2125,N_2158);
or U2284 (N_2284,N_2163,N_2113);
and U2285 (N_2285,N_2130,N_2117);
or U2286 (N_2286,N_2152,N_2120);
or U2287 (N_2287,N_2157,N_2140);
or U2288 (N_2288,N_2164,N_2197);
or U2289 (N_2289,N_2182,N_2140);
nor U2290 (N_2290,N_2182,N_2108);
and U2291 (N_2291,N_2133,N_2193);
nand U2292 (N_2292,N_2120,N_2137);
or U2293 (N_2293,N_2126,N_2160);
nor U2294 (N_2294,N_2135,N_2159);
or U2295 (N_2295,N_2121,N_2167);
and U2296 (N_2296,N_2126,N_2117);
and U2297 (N_2297,N_2143,N_2157);
nand U2298 (N_2298,N_2175,N_2114);
nor U2299 (N_2299,N_2114,N_2129);
and U2300 (N_2300,N_2244,N_2269);
and U2301 (N_2301,N_2267,N_2282);
nor U2302 (N_2302,N_2294,N_2210);
nand U2303 (N_2303,N_2258,N_2281);
nand U2304 (N_2304,N_2299,N_2276);
or U2305 (N_2305,N_2209,N_2235);
nand U2306 (N_2306,N_2289,N_2242);
or U2307 (N_2307,N_2255,N_2236);
or U2308 (N_2308,N_2284,N_2241);
or U2309 (N_2309,N_2222,N_2271);
or U2310 (N_2310,N_2296,N_2273);
and U2311 (N_2311,N_2200,N_2232);
and U2312 (N_2312,N_2220,N_2215);
nor U2313 (N_2313,N_2249,N_2272);
nor U2314 (N_2314,N_2230,N_2251);
nor U2315 (N_2315,N_2203,N_2216);
or U2316 (N_2316,N_2231,N_2226);
and U2317 (N_2317,N_2297,N_2298);
or U2318 (N_2318,N_2205,N_2268);
and U2319 (N_2319,N_2275,N_2264);
nor U2320 (N_2320,N_2261,N_2290);
nand U2321 (N_2321,N_2262,N_2233);
nand U2322 (N_2322,N_2259,N_2224);
xor U2323 (N_2323,N_2201,N_2213);
nand U2324 (N_2324,N_2240,N_2263);
nor U2325 (N_2325,N_2219,N_2239);
and U2326 (N_2326,N_2274,N_2291);
nor U2327 (N_2327,N_2221,N_2204);
nor U2328 (N_2328,N_2245,N_2250);
and U2329 (N_2329,N_2247,N_2237);
nand U2330 (N_2330,N_2229,N_2243);
nand U2331 (N_2331,N_2248,N_2218);
nand U2332 (N_2332,N_2293,N_2256);
nor U2333 (N_2333,N_2227,N_2206);
nor U2334 (N_2334,N_2277,N_2246);
and U2335 (N_2335,N_2228,N_2202);
nand U2336 (N_2336,N_2280,N_2217);
or U2337 (N_2337,N_2214,N_2211);
or U2338 (N_2338,N_2254,N_2212);
nor U2339 (N_2339,N_2225,N_2270);
or U2340 (N_2340,N_2283,N_2208);
nor U2341 (N_2341,N_2286,N_2279);
or U2342 (N_2342,N_2295,N_2285);
xor U2343 (N_2343,N_2266,N_2288);
and U2344 (N_2344,N_2253,N_2223);
nor U2345 (N_2345,N_2238,N_2234);
nand U2346 (N_2346,N_2252,N_2257);
or U2347 (N_2347,N_2292,N_2207);
and U2348 (N_2348,N_2260,N_2278);
or U2349 (N_2349,N_2265,N_2287);
nor U2350 (N_2350,N_2285,N_2220);
nand U2351 (N_2351,N_2296,N_2272);
or U2352 (N_2352,N_2271,N_2294);
nand U2353 (N_2353,N_2226,N_2203);
nor U2354 (N_2354,N_2284,N_2262);
nor U2355 (N_2355,N_2298,N_2218);
nand U2356 (N_2356,N_2276,N_2282);
nand U2357 (N_2357,N_2288,N_2226);
or U2358 (N_2358,N_2268,N_2261);
and U2359 (N_2359,N_2224,N_2253);
nand U2360 (N_2360,N_2262,N_2226);
and U2361 (N_2361,N_2299,N_2234);
or U2362 (N_2362,N_2242,N_2257);
and U2363 (N_2363,N_2259,N_2215);
or U2364 (N_2364,N_2273,N_2244);
or U2365 (N_2365,N_2249,N_2297);
nand U2366 (N_2366,N_2260,N_2277);
or U2367 (N_2367,N_2278,N_2291);
nor U2368 (N_2368,N_2225,N_2265);
nor U2369 (N_2369,N_2223,N_2281);
and U2370 (N_2370,N_2275,N_2207);
xnor U2371 (N_2371,N_2277,N_2256);
or U2372 (N_2372,N_2215,N_2248);
nor U2373 (N_2373,N_2292,N_2261);
nor U2374 (N_2374,N_2202,N_2266);
nand U2375 (N_2375,N_2203,N_2278);
or U2376 (N_2376,N_2293,N_2203);
nand U2377 (N_2377,N_2270,N_2212);
or U2378 (N_2378,N_2279,N_2237);
nor U2379 (N_2379,N_2295,N_2292);
and U2380 (N_2380,N_2291,N_2236);
nor U2381 (N_2381,N_2261,N_2219);
or U2382 (N_2382,N_2239,N_2211);
nand U2383 (N_2383,N_2241,N_2256);
and U2384 (N_2384,N_2289,N_2266);
or U2385 (N_2385,N_2223,N_2225);
nand U2386 (N_2386,N_2234,N_2269);
and U2387 (N_2387,N_2212,N_2275);
nor U2388 (N_2388,N_2272,N_2282);
nor U2389 (N_2389,N_2220,N_2298);
nor U2390 (N_2390,N_2206,N_2222);
nor U2391 (N_2391,N_2231,N_2283);
nand U2392 (N_2392,N_2293,N_2211);
nand U2393 (N_2393,N_2281,N_2218);
nor U2394 (N_2394,N_2212,N_2260);
nor U2395 (N_2395,N_2299,N_2288);
nand U2396 (N_2396,N_2234,N_2207);
or U2397 (N_2397,N_2254,N_2247);
and U2398 (N_2398,N_2293,N_2228);
and U2399 (N_2399,N_2274,N_2263);
and U2400 (N_2400,N_2340,N_2366);
or U2401 (N_2401,N_2333,N_2354);
or U2402 (N_2402,N_2351,N_2385);
nand U2403 (N_2403,N_2367,N_2383);
or U2404 (N_2404,N_2310,N_2378);
nor U2405 (N_2405,N_2386,N_2313);
or U2406 (N_2406,N_2392,N_2326);
and U2407 (N_2407,N_2315,N_2369);
or U2408 (N_2408,N_2309,N_2343);
nand U2409 (N_2409,N_2382,N_2338);
or U2410 (N_2410,N_2308,N_2368);
nand U2411 (N_2411,N_2334,N_2352);
nor U2412 (N_2412,N_2396,N_2399);
nor U2413 (N_2413,N_2302,N_2388);
or U2414 (N_2414,N_2374,N_2344);
nand U2415 (N_2415,N_2335,N_2319);
or U2416 (N_2416,N_2305,N_2362);
nand U2417 (N_2417,N_2356,N_2395);
nor U2418 (N_2418,N_2306,N_2324);
and U2419 (N_2419,N_2379,N_2397);
nand U2420 (N_2420,N_2336,N_2325);
or U2421 (N_2421,N_2364,N_2301);
and U2422 (N_2422,N_2393,N_2317);
or U2423 (N_2423,N_2394,N_2375);
or U2424 (N_2424,N_2365,N_2331);
nand U2425 (N_2425,N_2384,N_2332);
and U2426 (N_2426,N_2387,N_2304);
nor U2427 (N_2427,N_2389,N_2316);
and U2428 (N_2428,N_2330,N_2360);
and U2429 (N_2429,N_2347,N_2311);
nor U2430 (N_2430,N_2350,N_2361);
nor U2431 (N_2431,N_2381,N_2358);
nor U2432 (N_2432,N_2300,N_2323);
or U2433 (N_2433,N_2398,N_2376);
nand U2434 (N_2434,N_2312,N_2345);
nor U2435 (N_2435,N_2327,N_2363);
or U2436 (N_2436,N_2346,N_2348);
and U2437 (N_2437,N_2341,N_2359);
and U2438 (N_2438,N_2320,N_2353);
nand U2439 (N_2439,N_2321,N_2371);
or U2440 (N_2440,N_2337,N_2370);
nand U2441 (N_2441,N_2390,N_2372);
or U2442 (N_2442,N_2377,N_2303);
nor U2443 (N_2443,N_2328,N_2329);
nand U2444 (N_2444,N_2307,N_2349);
nor U2445 (N_2445,N_2318,N_2355);
and U2446 (N_2446,N_2342,N_2380);
and U2447 (N_2447,N_2391,N_2322);
nand U2448 (N_2448,N_2339,N_2373);
and U2449 (N_2449,N_2314,N_2357);
and U2450 (N_2450,N_2386,N_2341);
nor U2451 (N_2451,N_2324,N_2366);
and U2452 (N_2452,N_2306,N_2344);
or U2453 (N_2453,N_2334,N_2344);
or U2454 (N_2454,N_2398,N_2323);
nor U2455 (N_2455,N_2384,N_2325);
and U2456 (N_2456,N_2375,N_2390);
or U2457 (N_2457,N_2399,N_2367);
or U2458 (N_2458,N_2359,N_2337);
nand U2459 (N_2459,N_2340,N_2391);
and U2460 (N_2460,N_2386,N_2362);
nor U2461 (N_2461,N_2396,N_2356);
or U2462 (N_2462,N_2398,N_2371);
nand U2463 (N_2463,N_2350,N_2397);
and U2464 (N_2464,N_2316,N_2371);
nor U2465 (N_2465,N_2319,N_2301);
nand U2466 (N_2466,N_2318,N_2319);
nor U2467 (N_2467,N_2363,N_2317);
nor U2468 (N_2468,N_2327,N_2389);
nor U2469 (N_2469,N_2397,N_2384);
or U2470 (N_2470,N_2395,N_2375);
and U2471 (N_2471,N_2341,N_2350);
nor U2472 (N_2472,N_2307,N_2352);
and U2473 (N_2473,N_2348,N_2306);
nand U2474 (N_2474,N_2391,N_2373);
or U2475 (N_2475,N_2373,N_2388);
or U2476 (N_2476,N_2309,N_2316);
and U2477 (N_2477,N_2331,N_2324);
or U2478 (N_2478,N_2332,N_2343);
and U2479 (N_2479,N_2300,N_2394);
or U2480 (N_2480,N_2312,N_2335);
or U2481 (N_2481,N_2365,N_2374);
nor U2482 (N_2482,N_2303,N_2388);
or U2483 (N_2483,N_2336,N_2385);
or U2484 (N_2484,N_2344,N_2373);
nand U2485 (N_2485,N_2306,N_2304);
or U2486 (N_2486,N_2341,N_2307);
or U2487 (N_2487,N_2367,N_2364);
and U2488 (N_2488,N_2385,N_2365);
nand U2489 (N_2489,N_2387,N_2362);
nand U2490 (N_2490,N_2338,N_2342);
nand U2491 (N_2491,N_2381,N_2359);
and U2492 (N_2492,N_2344,N_2330);
and U2493 (N_2493,N_2328,N_2354);
or U2494 (N_2494,N_2301,N_2322);
and U2495 (N_2495,N_2355,N_2346);
nor U2496 (N_2496,N_2309,N_2398);
and U2497 (N_2497,N_2356,N_2368);
or U2498 (N_2498,N_2399,N_2316);
nor U2499 (N_2499,N_2346,N_2352);
nor U2500 (N_2500,N_2465,N_2416);
or U2501 (N_2501,N_2456,N_2414);
or U2502 (N_2502,N_2499,N_2448);
and U2503 (N_2503,N_2410,N_2462);
nor U2504 (N_2504,N_2452,N_2463);
nand U2505 (N_2505,N_2444,N_2408);
nor U2506 (N_2506,N_2402,N_2477);
nand U2507 (N_2507,N_2445,N_2485);
nor U2508 (N_2508,N_2418,N_2484);
nor U2509 (N_2509,N_2466,N_2459);
nor U2510 (N_2510,N_2468,N_2470);
nand U2511 (N_2511,N_2483,N_2467);
nor U2512 (N_2512,N_2413,N_2469);
or U2513 (N_2513,N_2497,N_2415);
nand U2514 (N_2514,N_2482,N_2424);
or U2515 (N_2515,N_2491,N_2403);
nand U2516 (N_2516,N_2431,N_2401);
or U2517 (N_2517,N_2437,N_2450);
or U2518 (N_2518,N_2407,N_2458);
nand U2519 (N_2519,N_2446,N_2461);
nor U2520 (N_2520,N_2464,N_2423);
and U2521 (N_2521,N_2476,N_2447);
nor U2522 (N_2522,N_2471,N_2427);
and U2523 (N_2523,N_2473,N_2480);
nor U2524 (N_2524,N_2409,N_2400);
nor U2525 (N_2525,N_2493,N_2496);
or U2526 (N_2526,N_2451,N_2425);
or U2527 (N_2527,N_2495,N_2411);
nand U2528 (N_2528,N_2428,N_2435);
nand U2529 (N_2529,N_2490,N_2406);
or U2530 (N_2530,N_2436,N_2419);
nor U2531 (N_2531,N_2440,N_2439);
or U2532 (N_2532,N_2486,N_2426);
nor U2533 (N_2533,N_2441,N_2453);
nor U2534 (N_2534,N_2434,N_2474);
nor U2535 (N_2535,N_2432,N_2405);
nand U2536 (N_2536,N_2433,N_2457);
and U2537 (N_2537,N_2443,N_2460);
and U2538 (N_2538,N_2472,N_2429);
and U2539 (N_2539,N_2489,N_2487);
xnor U2540 (N_2540,N_2420,N_2455);
and U2541 (N_2541,N_2488,N_2442);
nand U2542 (N_2542,N_2449,N_2417);
nor U2543 (N_2543,N_2412,N_2479);
nand U2544 (N_2544,N_2421,N_2481);
nand U2545 (N_2545,N_2438,N_2498);
and U2546 (N_2546,N_2475,N_2494);
or U2547 (N_2547,N_2422,N_2492);
or U2548 (N_2548,N_2404,N_2430);
or U2549 (N_2549,N_2478,N_2454);
or U2550 (N_2550,N_2437,N_2447);
nand U2551 (N_2551,N_2461,N_2480);
nand U2552 (N_2552,N_2432,N_2436);
nand U2553 (N_2553,N_2487,N_2467);
nand U2554 (N_2554,N_2482,N_2473);
and U2555 (N_2555,N_2400,N_2481);
or U2556 (N_2556,N_2495,N_2474);
or U2557 (N_2557,N_2457,N_2436);
or U2558 (N_2558,N_2471,N_2470);
nor U2559 (N_2559,N_2406,N_2460);
nor U2560 (N_2560,N_2498,N_2404);
and U2561 (N_2561,N_2462,N_2426);
nand U2562 (N_2562,N_2436,N_2495);
nor U2563 (N_2563,N_2474,N_2427);
nand U2564 (N_2564,N_2446,N_2498);
or U2565 (N_2565,N_2433,N_2417);
nor U2566 (N_2566,N_2470,N_2436);
nor U2567 (N_2567,N_2480,N_2476);
or U2568 (N_2568,N_2451,N_2455);
nand U2569 (N_2569,N_2431,N_2410);
nor U2570 (N_2570,N_2483,N_2439);
nand U2571 (N_2571,N_2401,N_2452);
nor U2572 (N_2572,N_2420,N_2470);
nand U2573 (N_2573,N_2474,N_2490);
or U2574 (N_2574,N_2445,N_2479);
nand U2575 (N_2575,N_2457,N_2427);
or U2576 (N_2576,N_2462,N_2446);
or U2577 (N_2577,N_2498,N_2492);
nor U2578 (N_2578,N_2458,N_2432);
nor U2579 (N_2579,N_2405,N_2498);
and U2580 (N_2580,N_2494,N_2484);
nor U2581 (N_2581,N_2497,N_2477);
and U2582 (N_2582,N_2496,N_2478);
nand U2583 (N_2583,N_2485,N_2424);
nor U2584 (N_2584,N_2465,N_2436);
or U2585 (N_2585,N_2420,N_2432);
or U2586 (N_2586,N_2416,N_2413);
nand U2587 (N_2587,N_2476,N_2471);
or U2588 (N_2588,N_2441,N_2482);
or U2589 (N_2589,N_2415,N_2458);
or U2590 (N_2590,N_2426,N_2450);
and U2591 (N_2591,N_2440,N_2441);
nand U2592 (N_2592,N_2469,N_2466);
or U2593 (N_2593,N_2452,N_2432);
and U2594 (N_2594,N_2439,N_2468);
nand U2595 (N_2595,N_2412,N_2483);
and U2596 (N_2596,N_2409,N_2478);
nor U2597 (N_2597,N_2411,N_2410);
or U2598 (N_2598,N_2436,N_2401);
nor U2599 (N_2599,N_2443,N_2433);
nor U2600 (N_2600,N_2560,N_2505);
nor U2601 (N_2601,N_2563,N_2525);
nor U2602 (N_2602,N_2577,N_2557);
and U2603 (N_2603,N_2504,N_2559);
nor U2604 (N_2604,N_2520,N_2541);
nand U2605 (N_2605,N_2568,N_2518);
and U2606 (N_2606,N_2558,N_2521);
and U2607 (N_2607,N_2537,N_2546);
nor U2608 (N_2608,N_2527,N_2580);
nand U2609 (N_2609,N_2582,N_2579);
and U2610 (N_2610,N_2512,N_2530);
and U2611 (N_2611,N_2511,N_2567);
and U2612 (N_2612,N_2586,N_2561);
or U2613 (N_2613,N_2592,N_2535);
or U2614 (N_2614,N_2587,N_2581);
or U2615 (N_2615,N_2570,N_2532);
nand U2616 (N_2616,N_2508,N_2556);
and U2617 (N_2617,N_2545,N_2540);
and U2618 (N_2618,N_2538,N_2588);
and U2619 (N_2619,N_2510,N_2536);
and U2620 (N_2620,N_2596,N_2595);
or U2621 (N_2621,N_2503,N_2509);
nor U2622 (N_2622,N_2542,N_2516);
nor U2623 (N_2623,N_2539,N_2552);
and U2624 (N_2624,N_2524,N_2598);
or U2625 (N_2625,N_2578,N_2576);
and U2626 (N_2626,N_2548,N_2594);
and U2627 (N_2627,N_2555,N_2543);
nor U2628 (N_2628,N_2564,N_2529);
nor U2629 (N_2629,N_2574,N_2544);
or U2630 (N_2630,N_2553,N_2571);
or U2631 (N_2631,N_2501,N_2533);
and U2632 (N_2632,N_2519,N_2569);
nand U2633 (N_2633,N_2507,N_2515);
nand U2634 (N_2634,N_2506,N_2528);
nor U2635 (N_2635,N_2583,N_2589);
nor U2636 (N_2636,N_2551,N_2585);
or U2637 (N_2637,N_2591,N_2573);
or U2638 (N_2638,N_2526,N_2547);
nand U2639 (N_2639,N_2502,N_2572);
and U2640 (N_2640,N_2575,N_2593);
or U2641 (N_2641,N_2565,N_2534);
nor U2642 (N_2642,N_2566,N_2549);
nor U2643 (N_2643,N_2597,N_2517);
or U2644 (N_2644,N_2531,N_2550);
nand U2645 (N_2645,N_2514,N_2590);
nor U2646 (N_2646,N_2584,N_2562);
and U2647 (N_2647,N_2554,N_2522);
and U2648 (N_2648,N_2523,N_2500);
and U2649 (N_2649,N_2513,N_2599);
and U2650 (N_2650,N_2517,N_2504);
and U2651 (N_2651,N_2554,N_2531);
and U2652 (N_2652,N_2588,N_2502);
or U2653 (N_2653,N_2579,N_2543);
and U2654 (N_2654,N_2537,N_2540);
nor U2655 (N_2655,N_2508,N_2531);
and U2656 (N_2656,N_2587,N_2568);
nor U2657 (N_2657,N_2502,N_2503);
nand U2658 (N_2658,N_2514,N_2549);
nand U2659 (N_2659,N_2504,N_2507);
and U2660 (N_2660,N_2549,N_2570);
nand U2661 (N_2661,N_2504,N_2573);
nand U2662 (N_2662,N_2575,N_2523);
or U2663 (N_2663,N_2557,N_2502);
or U2664 (N_2664,N_2582,N_2585);
xor U2665 (N_2665,N_2598,N_2534);
or U2666 (N_2666,N_2592,N_2512);
nor U2667 (N_2667,N_2558,N_2589);
nand U2668 (N_2668,N_2587,N_2598);
or U2669 (N_2669,N_2579,N_2529);
or U2670 (N_2670,N_2544,N_2512);
or U2671 (N_2671,N_2538,N_2587);
and U2672 (N_2672,N_2548,N_2543);
or U2673 (N_2673,N_2594,N_2593);
and U2674 (N_2674,N_2568,N_2572);
and U2675 (N_2675,N_2590,N_2500);
and U2676 (N_2676,N_2520,N_2599);
nand U2677 (N_2677,N_2508,N_2583);
or U2678 (N_2678,N_2580,N_2556);
and U2679 (N_2679,N_2587,N_2565);
or U2680 (N_2680,N_2551,N_2514);
nand U2681 (N_2681,N_2573,N_2520);
or U2682 (N_2682,N_2556,N_2528);
or U2683 (N_2683,N_2510,N_2521);
nor U2684 (N_2684,N_2556,N_2542);
and U2685 (N_2685,N_2549,N_2569);
and U2686 (N_2686,N_2534,N_2593);
nand U2687 (N_2687,N_2524,N_2516);
or U2688 (N_2688,N_2523,N_2535);
and U2689 (N_2689,N_2527,N_2564);
and U2690 (N_2690,N_2538,N_2547);
or U2691 (N_2691,N_2591,N_2595);
nor U2692 (N_2692,N_2574,N_2535);
and U2693 (N_2693,N_2571,N_2527);
or U2694 (N_2694,N_2529,N_2533);
nand U2695 (N_2695,N_2537,N_2586);
and U2696 (N_2696,N_2553,N_2595);
or U2697 (N_2697,N_2534,N_2535);
and U2698 (N_2698,N_2575,N_2528);
or U2699 (N_2699,N_2555,N_2558);
nor U2700 (N_2700,N_2688,N_2616);
nand U2701 (N_2701,N_2680,N_2667);
and U2702 (N_2702,N_2681,N_2622);
nor U2703 (N_2703,N_2699,N_2634);
and U2704 (N_2704,N_2695,N_2637);
nor U2705 (N_2705,N_2678,N_2615);
nand U2706 (N_2706,N_2654,N_2609);
nor U2707 (N_2707,N_2651,N_2692);
nand U2708 (N_2708,N_2647,N_2606);
and U2709 (N_2709,N_2664,N_2646);
nand U2710 (N_2710,N_2638,N_2642);
and U2711 (N_2711,N_2644,N_2632);
nor U2712 (N_2712,N_2666,N_2633);
nor U2713 (N_2713,N_2618,N_2683);
or U2714 (N_2714,N_2628,N_2682);
xor U2715 (N_2715,N_2623,N_2619);
nor U2716 (N_2716,N_2687,N_2611);
or U2717 (N_2717,N_2657,N_2698);
nor U2718 (N_2718,N_2652,N_2641);
or U2719 (N_2719,N_2694,N_2677);
and U2720 (N_2720,N_2639,N_2603);
nor U2721 (N_2721,N_2613,N_2625);
nor U2722 (N_2722,N_2608,N_2691);
and U2723 (N_2723,N_2627,N_2671);
and U2724 (N_2724,N_2659,N_2614);
and U2725 (N_2725,N_2672,N_2624);
nor U2726 (N_2726,N_2635,N_2668);
or U2727 (N_2727,N_2653,N_2662);
nor U2728 (N_2728,N_2600,N_2670);
nor U2729 (N_2729,N_2697,N_2661);
or U2730 (N_2730,N_2656,N_2620);
nand U2731 (N_2731,N_2676,N_2686);
and U2732 (N_2732,N_2650,N_2658);
and U2733 (N_2733,N_2640,N_2601);
nor U2734 (N_2734,N_2612,N_2617);
nor U2735 (N_2735,N_2690,N_2684);
and U2736 (N_2736,N_2636,N_2631);
and U2737 (N_2737,N_2605,N_2679);
and U2738 (N_2738,N_2648,N_2693);
or U2739 (N_2739,N_2645,N_2660);
nand U2740 (N_2740,N_2602,N_2607);
nand U2741 (N_2741,N_2669,N_2649);
nor U2742 (N_2742,N_2604,N_2689);
or U2743 (N_2743,N_2643,N_2610);
and U2744 (N_2744,N_2696,N_2674);
nor U2745 (N_2745,N_2630,N_2663);
nand U2746 (N_2746,N_2675,N_2626);
or U2747 (N_2747,N_2621,N_2685);
or U2748 (N_2748,N_2665,N_2629);
or U2749 (N_2749,N_2655,N_2673);
nand U2750 (N_2750,N_2652,N_2664);
nor U2751 (N_2751,N_2675,N_2670);
nor U2752 (N_2752,N_2618,N_2612);
and U2753 (N_2753,N_2638,N_2647);
nand U2754 (N_2754,N_2687,N_2683);
and U2755 (N_2755,N_2600,N_2655);
nand U2756 (N_2756,N_2615,N_2676);
nor U2757 (N_2757,N_2627,N_2620);
nor U2758 (N_2758,N_2618,N_2619);
or U2759 (N_2759,N_2683,N_2688);
and U2760 (N_2760,N_2696,N_2678);
nor U2761 (N_2761,N_2619,N_2621);
nor U2762 (N_2762,N_2649,N_2681);
and U2763 (N_2763,N_2679,N_2665);
nand U2764 (N_2764,N_2655,N_2670);
nand U2765 (N_2765,N_2680,N_2607);
and U2766 (N_2766,N_2625,N_2657);
or U2767 (N_2767,N_2696,N_2683);
nand U2768 (N_2768,N_2656,N_2604);
nor U2769 (N_2769,N_2647,N_2660);
xnor U2770 (N_2770,N_2677,N_2621);
or U2771 (N_2771,N_2665,N_2623);
and U2772 (N_2772,N_2657,N_2624);
nand U2773 (N_2773,N_2657,N_2601);
or U2774 (N_2774,N_2682,N_2672);
nand U2775 (N_2775,N_2639,N_2604);
nand U2776 (N_2776,N_2613,N_2608);
nand U2777 (N_2777,N_2648,N_2681);
and U2778 (N_2778,N_2624,N_2688);
nand U2779 (N_2779,N_2696,N_2658);
nand U2780 (N_2780,N_2602,N_2690);
nor U2781 (N_2781,N_2699,N_2668);
nand U2782 (N_2782,N_2676,N_2632);
and U2783 (N_2783,N_2689,N_2600);
and U2784 (N_2784,N_2693,N_2667);
and U2785 (N_2785,N_2618,N_2691);
or U2786 (N_2786,N_2610,N_2693);
and U2787 (N_2787,N_2670,N_2666);
nor U2788 (N_2788,N_2640,N_2696);
and U2789 (N_2789,N_2673,N_2635);
nor U2790 (N_2790,N_2630,N_2684);
and U2791 (N_2791,N_2669,N_2608);
nand U2792 (N_2792,N_2695,N_2616);
or U2793 (N_2793,N_2656,N_2671);
nand U2794 (N_2794,N_2637,N_2648);
or U2795 (N_2795,N_2657,N_2639);
or U2796 (N_2796,N_2623,N_2680);
and U2797 (N_2797,N_2613,N_2689);
nand U2798 (N_2798,N_2643,N_2648);
or U2799 (N_2799,N_2650,N_2607);
xnor U2800 (N_2800,N_2711,N_2784);
or U2801 (N_2801,N_2767,N_2771);
nor U2802 (N_2802,N_2710,N_2743);
nand U2803 (N_2803,N_2795,N_2746);
nor U2804 (N_2804,N_2752,N_2718);
or U2805 (N_2805,N_2742,N_2732);
nor U2806 (N_2806,N_2741,N_2724);
nand U2807 (N_2807,N_2797,N_2766);
nand U2808 (N_2808,N_2799,N_2788);
or U2809 (N_2809,N_2768,N_2753);
or U2810 (N_2810,N_2761,N_2764);
nand U2811 (N_2811,N_2745,N_2770);
or U2812 (N_2812,N_2721,N_2713);
nor U2813 (N_2813,N_2791,N_2777);
nand U2814 (N_2814,N_2786,N_2730);
or U2815 (N_2815,N_2704,N_2733);
nand U2816 (N_2816,N_2790,N_2760);
or U2817 (N_2817,N_2763,N_2736);
nor U2818 (N_2818,N_2726,N_2787);
nand U2819 (N_2819,N_2757,N_2793);
nor U2820 (N_2820,N_2782,N_2723);
nor U2821 (N_2821,N_2756,N_2754);
nor U2822 (N_2822,N_2775,N_2708);
and U2823 (N_2823,N_2717,N_2744);
nor U2824 (N_2824,N_2776,N_2709);
nor U2825 (N_2825,N_2722,N_2762);
nor U2826 (N_2826,N_2728,N_2735);
nor U2827 (N_2827,N_2703,N_2794);
and U2828 (N_2828,N_2706,N_2739);
or U2829 (N_2829,N_2751,N_2749);
and U2830 (N_2830,N_2778,N_2734);
nor U2831 (N_2831,N_2748,N_2781);
and U2832 (N_2832,N_2712,N_2707);
or U2833 (N_2833,N_2701,N_2737);
or U2834 (N_2834,N_2714,N_2783);
and U2835 (N_2835,N_2758,N_2772);
or U2836 (N_2836,N_2720,N_2747);
or U2837 (N_2837,N_2769,N_2755);
nand U2838 (N_2838,N_2798,N_2773);
or U2839 (N_2839,N_2789,N_2725);
nor U2840 (N_2840,N_2779,N_2740);
nand U2841 (N_2841,N_2738,N_2729);
and U2842 (N_2842,N_2792,N_2719);
and U2843 (N_2843,N_2796,N_2759);
xor U2844 (N_2844,N_2702,N_2765);
nor U2845 (N_2845,N_2715,N_2785);
nand U2846 (N_2846,N_2774,N_2700);
or U2847 (N_2847,N_2731,N_2716);
or U2848 (N_2848,N_2750,N_2780);
nor U2849 (N_2849,N_2705,N_2727);
nor U2850 (N_2850,N_2776,N_2753);
or U2851 (N_2851,N_2781,N_2741);
and U2852 (N_2852,N_2795,N_2782);
nand U2853 (N_2853,N_2724,N_2720);
or U2854 (N_2854,N_2755,N_2763);
or U2855 (N_2855,N_2769,N_2762);
nand U2856 (N_2856,N_2776,N_2710);
or U2857 (N_2857,N_2770,N_2706);
and U2858 (N_2858,N_2746,N_2770);
and U2859 (N_2859,N_2746,N_2707);
nand U2860 (N_2860,N_2799,N_2777);
and U2861 (N_2861,N_2703,N_2772);
nand U2862 (N_2862,N_2756,N_2778);
or U2863 (N_2863,N_2727,N_2797);
nor U2864 (N_2864,N_2764,N_2737);
and U2865 (N_2865,N_2730,N_2740);
nand U2866 (N_2866,N_2762,N_2743);
or U2867 (N_2867,N_2798,N_2700);
or U2868 (N_2868,N_2772,N_2736);
and U2869 (N_2869,N_2789,N_2717);
and U2870 (N_2870,N_2717,N_2768);
or U2871 (N_2871,N_2720,N_2759);
and U2872 (N_2872,N_2706,N_2788);
nor U2873 (N_2873,N_2767,N_2774);
and U2874 (N_2874,N_2797,N_2702);
or U2875 (N_2875,N_2712,N_2756);
or U2876 (N_2876,N_2751,N_2778);
nand U2877 (N_2877,N_2779,N_2712);
and U2878 (N_2878,N_2752,N_2744);
nand U2879 (N_2879,N_2784,N_2714);
or U2880 (N_2880,N_2736,N_2735);
and U2881 (N_2881,N_2751,N_2784);
nor U2882 (N_2882,N_2751,N_2738);
or U2883 (N_2883,N_2741,N_2719);
and U2884 (N_2884,N_2737,N_2745);
nor U2885 (N_2885,N_2789,N_2720);
or U2886 (N_2886,N_2768,N_2719);
nand U2887 (N_2887,N_2794,N_2765);
nand U2888 (N_2888,N_2729,N_2750);
nand U2889 (N_2889,N_2757,N_2784);
or U2890 (N_2890,N_2733,N_2709);
and U2891 (N_2891,N_2794,N_2715);
nor U2892 (N_2892,N_2706,N_2745);
or U2893 (N_2893,N_2787,N_2719);
nor U2894 (N_2894,N_2720,N_2757);
nor U2895 (N_2895,N_2781,N_2707);
or U2896 (N_2896,N_2721,N_2738);
or U2897 (N_2897,N_2767,N_2766);
or U2898 (N_2898,N_2762,N_2775);
nor U2899 (N_2899,N_2764,N_2735);
nor U2900 (N_2900,N_2823,N_2819);
nor U2901 (N_2901,N_2808,N_2852);
or U2902 (N_2902,N_2899,N_2886);
nand U2903 (N_2903,N_2843,N_2801);
xor U2904 (N_2904,N_2854,N_2841);
nor U2905 (N_2905,N_2811,N_2879);
nand U2906 (N_2906,N_2813,N_2844);
nor U2907 (N_2907,N_2867,N_2814);
or U2908 (N_2908,N_2817,N_2875);
and U2909 (N_2909,N_2805,N_2898);
and U2910 (N_2910,N_2831,N_2868);
nor U2911 (N_2911,N_2860,N_2839);
nand U2912 (N_2912,N_2851,N_2812);
or U2913 (N_2913,N_2848,N_2894);
and U2914 (N_2914,N_2885,N_2849);
and U2915 (N_2915,N_2847,N_2846);
and U2916 (N_2916,N_2857,N_2872);
nor U2917 (N_2917,N_2830,N_2891);
nand U2918 (N_2918,N_2896,N_2858);
nand U2919 (N_2919,N_2815,N_2822);
nor U2920 (N_2920,N_2828,N_2816);
and U2921 (N_2921,N_2832,N_2825);
nor U2922 (N_2922,N_2859,N_2835);
nand U2923 (N_2923,N_2855,N_2892);
nor U2924 (N_2924,N_2804,N_2840);
or U2925 (N_2925,N_2873,N_2881);
nor U2926 (N_2926,N_2888,N_2877);
nor U2927 (N_2927,N_2826,N_2837);
nand U2928 (N_2928,N_2820,N_2806);
nor U2929 (N_2929,N_2836,N_2818);
and U2930 (N_2930,N_2807,N_2809);
nand U2931 (N_2931,N_2866,N_2865);
nor U2932 (N_2932,N_2887,N_2802);
and U2933 (N_2933,N_2827,N_2871);
and U2934 (N_2934,N_2833,N_2876);
nand U2935 (N_2935,N_2853,N_2856);
and U2936 (N_2936,N_2862,N_2884);
and U2937 (N_2937,N_2897,N_2845);
nand U2938 (N_2938,N_2803,N_2878);
and U2939 (N_2939,N_2863,N_2800);
nand U2940 (N_2940,N_2861,N_2834);
or U2941 (N_2941,N_2880,N_2883);
and U2942 (N_2942,N_2889,N_2895);
or U2943 (N_2943,N_2890,N_2874);
or U2944 (N_2944,N_2821,N_2893);
or U2945 (N_2945,N_2829,N_2824);
nand U2946 (N_2946,N_2882,N_2869);
or U2947 (N_2947,N_2810,N_2864);
or U2948 (N_2948,N_2870,N_2850);
or U2949 (N_2949,N_2842,N_2838);
nand U2950 (N_2950,N_2858,N_2845);
or U2951 (N_2951,N_2870,N_2815);
nand U2952 (N_2952,N_2877,N_2804);
or U2953 (N_2953,N_2813,N_2835);
nand U2954 (N_2954,N_2817,N_2854);
or U2955 (N_2955,N_2838,N_2889);
nor U2956 (N_2956,N_2812,N_2813);
nor U2957 (N_2957,N_2878,N_2827);
nand U2958 (N_2958,N_2824,N_2835);
or U2959 (N_2959,N_2854,N_2803);
or U2960 (N_2960,N_2864,N_2894);
or U2961 (N_2961,N_2814,N_2886);
or U2962 (N_2962,N_2873,N_2842);
nand U2963 (N_2963,N_2875,N_2893);
and U2964 (N_2964,N_2842,N_2857);
and U2965 (N_2965,N_2838,N_2802);
or U2966 (N_2966,N_2870,N_2832);
or U2967 (N_2967,N_2803,N_2852);
and U2968 (N_2968,N_2870,N_2855);
nand U2969 (N_2969,N_2838,N_2836);
and U2970 (N_2970,N_2814,N_2816);
nor U2971 (N_2971,N_2843,N_2813);
or U2972 (N_2972,N_2839,N_2849);
nand U2973 (N_2973,N_2813,N_2802);
or U2974 (N_2974,N_2886,N_2850);
nor U2975 (N_2975,N_2810,N_2876);
nor U2976 (N_2976,N_2888,N_2821);
nor U2977 (N_2977,N_2809,N_2861);
nor U2978 (N_2978,N_2899,N_2832);
or U2979 (N_2979,N_2830,N_2888);
nand U2980 (N_2980,N_2824,N_2805);
nand U2981 (N_2981,N_2806,N_2897);
nand U2982 (N_2982,N_2837,N_2809);
nand U2983 (N_2983,N_2842,N_2831);
nand U2984 (N_2984,N_2842,N_2847);
nor U2985 (N_2985,N_2868,N_2890);
nand U2986 (N_2986,N_2894,N_2889);
xor U2987 (N_2987,N_2879,N_2857);
or U2988 (N_2988,N_2858,N_2883);
nor U2989 (N_2989,N_2886,N_2870);
or U2990 (N_2990,N_2887,N_2867);
and U2991 (N_2991,N_2849,N_2832);
and U2992 (N_2992,N_2822,N_2878);
and U2993 (N_2993,N_2882,N_2821);
nor U2994 (N_2994,N_2887,N_2886);
nor U2995 (N_2995,N_2871,N_2895);
nand U2996 (N_2996,N_2814,N_2807);
and U2997 (N_2997,N_2844,N_2865);
or U2998 (N_2998,N_2851,N_2806);
nor U2999 (N_2999,N_2848,N_2880);
nand UO_0 (O_0,N_2976,N_2982);
and UO_1 (O_1,N_2935,N_2991);
nand UO_2 (O_2,N_2940,N_2998);
and UO_3 (O_3,N_2937,N_2930);
and UO_4 (O_4,N_2928,N_2994);
and UO_5 (O_5,N_2965,N_2975);
nor UO_6 (O_6,N_2933,N_2980);
or UO_7 (O_7,N_2921,N_2995);
and UO_8 (O_8,N_2952,N_2919);
nor UO_9 (O_9,N_2944,N_2984);
nor UO_10 (O_10,N_2979,N_2923);
or UO_11 (O_11,N_2904,N_2951);
and UO_12 (O_12,N_2929,N_2943);
nand UO_13 (O_13,N_2986,N_2996);
or UO_14 (O_14,N_2932,N_2992);
and UO_15 (O_15,N_2917,N_2926);
and UO_16 (O_16,N_2910,N_2956);
nand UO_17 (O_17,N_2977,N_2934);
or UO_18 (O_18,N_2974,N_2993);
nor UO_19 (O_19,N_2927,N_2957);
nand UO_20 (O_20,N_2967,N_2969);
and UO_21 (O_21,N_2949,N_2912);
and UO_22 (O_22,N_2968,N_2970);
nor UO_23 (O_23,N_2966,N_2931);
and UO_24 (O_24,N_2922,N_2990);
nor UO_25 (O_25,N_2972,N_2913);
nor UO_26 (O_26,N_2964,N_2911);
nor UO_27 (O_27,N_2983,N_2908);
nand UO_28 (O_28,N_2909,N_2918);
nor UO_29 (O_29,N_2942,N_2958);
or UO_30 (O_30,N_2978,N_2989);
nand UO_31 (O_31,N_2916,N_2948);
nand UO_32 (O_32,N_2981,N_2987);
nand UO_33 (O_33,N_2999,N_2955);
and UO_34 (O_34,N_2902,N_2941);
nand UO_35 (O_35,N_2920,N_2959);
and UO_36 (O_36,N_2945,N_2961);
nand UO_37 (O_37,N_2936,N_2963);
or UO_38 (O_38,N_2938,N_2960);
or UO_39 (O_39,N_2962,N_2973);
nand UO_40 (O_40,N_2950,N_2947);
nand UO_41 (O_41,N_2985,N_2924);
nand UO_42 (O_42,N_2971,N_2954);
or UO_43 (O_43,N_2925,N_2903);
or UO_44 (O_44,N_2907,N_2900);
or UO_45 (O_45,N_2915,N_2905);
nor UO_46 (O_46,N_2997,N_2906);
xnor UO_47 (O_47,N_2953,N_2914);
nor UO_48 (O_48,N_2939,N_2901);
and UO_49 (O_49,N_2988,N_2946);
and UO_50 (O_50,N_2969,N_2945);
nand UO_51 (O_51,N_2915,N_2920);
nor UO_52 (O_52,N_2918,N_2917);
nand UO_53 (O_53,N_2959,N_2995);
or UO_54 (O_54,N_2905,N_2998);
or UO_55 (O_55,N_2914,N_2900);
nor UO_56 (O_56,N_2962,N_2991);
nand UO_57 (O_57,N_2964,N_2959);
and UO_58 (O_58,N_2993,N_2970);
or UO_59 (O_59,N_2919,N_2926);
nand UO_60 (O_60,N_2921,N_2900);
and UO_61 (O_61,N_2986,N_2926);
and UO_62 (O_62,N_2906,N_2943);
and UO_63 (O_63,N_2949,N_2960);
nand UO_64 (O_64,N_2971,N_2925);
nand UO_65 (O_65,N_2961,N_2928);
nand UO_66 (O_66,N_2978,N_2928);
or UO_67 (O_67,N_2913,N_2939);
or UO_68 (O_68,N_2976,N_2960);
nand UO_69 (O_69,N_2978,N_2940);
and UO_70 (O_70,N_2938,N_2904);
nor UO_71 (O_71,N_2953,N_2960);
nand UO_72 (O_72,N_2970,N_2964);
or UO_73 (O_73,N_2901,N_2927);
nor UO_74 (O_74,N_2957,N_2963);
nor UO_75 (O_75,N_2944,N_2970);
or UO_76 (O_76,N_2947,N_2931);
nand UO_77 (O_77,N_2911,N_2914);
nand UO_78 (O_78,N_2932,N_2980);
nor UO_79 (O_79,N_2987,N_2995);
or UO_80 (O_80,N_2958,N_2968);
nor UO_81 (O_81,N_2993,N_2954);
nand UO_82 (O_82,N_2971,N_2998);
nand UO_83 (O_83,N_2904,N_2971);
and UO_84 (O_84,N_2920,N_2947);
and UO_85 (O_85,N_2951,N_2958);
nor UO_86 (O_86,N_2902,N_2937);
and UO_87 (O_87,N_2904,N_2979);
or UO_88 (O_88,N_2901,N_2912);
and UO_89 (O_89,N_2911,N_2934);
or UO_90 (O_90,N_2954,N_2962);
nand UO_91 (O_91,N_2989,N_2993);
and UO_92 (O_92,N_2950,N_2968);
or UO_93 (O_93,N_2992,N_2952);
nand UO_94 (O_94,N_2941,N_2994);
or UO_95 (O_95,N_2948,N_2961);
and UO_96 (O_96,N_2997,N_2916);
nor UO_97 (O_97,N_2983,N_2917);
nor UO_98 (O_98,N_2930,N_2996);
and UO_99 (O_99,N_2994,N_2985);
nor UO_100 (O_100,N_2927,N_2947);
or UO_101 (O_101,N_2946,N_2932);
nor UO_102 (O_102,N_2920,N_2929);
nor UO_103 (O_103,N_2969,N_2977);
and UO_104 (O_104,N_2901,N_2916);
nor UO_105 (O_105,N_2960,N_2947);
and UO_106 (O_106,N_2943,N_2997);
nand UO_107 (O_107,N_2986,N_2992);
nor UO_108 (O_108,N_2943,N_2996);
or UO_109 (O_109,N_2985,N_2920);
nand UO_110 (O_110,N_2985,N_2921);
nor UO_111 (O_111,N_2973,N_2967);
nor UO_112 (O_112,N_2990,N_2908);
nand UO_113 (O_113,N_2943,N_2968);
or UO_114 (O_114,N_2946,N_2900);
nor UO_115 (O_115,N_2933,N_2994);
and UO_116 (O_116,N_2948,N_2909);
nor UO_117 (O_117,N_2924,N_2979);
or UO_118 (O_118,N_2943,N_2960);
or UO_119 (O_119,N_2987,N_2982);
nor UO_120 (O_120,N_2919,N_2936);
and UO_121 (O_121,N_2997,N_2904);
and UO_122 (O_122,N_2987,N_2907);
or UO_123 (O_123,N_2993,N_2957);
nand UO_124 (O_124,N_2993,N_2960);
or UO_125 (O_125,N_2910,N_2962);
nor UO_126 (O_126,N_2990,N_2967);
nor UO_127 (O_127,N_2982,N_2933);
nor UO_128 (O_128,N_2980,N_2911);
nor UO_129 (O_129,N_2976,N_2928);
and UO_130 (O_130,N_2932,N_2907);
nand UO_131 (O_131,N_2971,N_2959);
and UO_132 (O_132,N_2962,N_2950);
or UO_133 (O_133,N_2903,N_2965);
or UO_134 (O_134,N_2937,N_2983);
nor UO_135 (O_135,N_2981,N_2948);
and UO_136 (O_136,N_2956,N_2961);
nor UO_137 (O_137,N_2963,N_2951);
and UO_138 (O_138,N_2967,N_2997);
nand UO_139 (O_139,N_2960,N_2978);
or UO_140 (O_140,N_2950,N_2940);
nand UO_141 (O_141,N_2958,N_2926);
and UO_142 (O_142,N_2952,N_2960);
nor UO_143 (O_143,N_2903,N_2904);
or UO_144 (O_144,N_2936,N_2934);
nor UO_145 (O_145,N_2920,N_2930);
nor UO_146 (O_146,N_2926,N_2916);
nor UO_147 (O_147,N_2923,N_2947);
nand UO_148 (O_148,N_2925,N_2987);
nor UO_149 (O_149,N_2953,N_2994);
or UO_150 (O_150,N_2927,N_2961);
and UO_151 (O_151,N_2919,N_2956);
nor UO_152 (O_152,N_2912,N_2996);
and UO_153 (O_153,N_2972,N_2977);
nor UO_154 (O_154,N_2992,N_2985);
and UO_155 (O_155,N_2941,N_2990);
nand UO_156 (O_156,N_2912,N_2988);
nor UO_157 (O_157,N_2928,N_2970);
nand UO_158 (O_158,N_2991,N_2989);
nor UO_159 (O_159,N_2929,N_2942);
or UO_160 (O_160,N_2934,N_2923);
nor UO_161 (O_161,N_2938,N_2931);
nor UO_162 (O_162,N_2990,N_2913);
nand UO_163 (O_163,N_2981,N_2947);
nand UO_164 (O_164,N_2957,N_2999);
and UO_165 (O_165,N_2931,N_2905);
and UO_166 (O_166,N_2911,N_2935);
and UO_167 (O_167,N_2971,N_2926);
and UO_168 (O_168,N_2961,N_2915);
or UO_169 (O_169,N_2901,N_2953);
or UO_170 (O_170,N_2972,N_2955);
or UO_171 (O_171,N_2969,N_2983);
or UO_172 (O_172,N_2920,N_2934);
and UO_173 (O_173,N_2999,N_2960);
nand UO_174 (O_174,N_2963,N_2938);
nor UO_175 (O_175,N_2984,N_2929);
nand UO_176 (O_176,N_2991,N_2995);
nand UO_177 (O_177,N_2990,N_2954);
or UO_178 (O_178,N_2908,N_2968);
or UO_179 (O_179,N_2936,N_2903);
nor UO_180 (O_180,N_2933,N_2935);
or UO_181 (O_181,N_2937,N_2904);
nand UO_182 (O_182,N_2957,N_2995);
nand UO_183 (O_183,N_2953,N_2985);
nor UO_184 (O_184,N_2977,N_2942);
nand UO_185 (O_185,N_2938,N_2997);
nor UO_186 (O_186,N_2983,N_2957);
nand UO_187 (O_187,N_2949,N_2931);
nor UO_188 (O_188,N_2949,N_2966);
and UO_189 (O_189,N_2986,N_2955);
nand UO_190 (O_190,N_2948,N_2932);
and UO_191 (O_191,N_2995,N_2961);
and UO_192 (O_192,N_2983,N_2928);
or UO_193 (O_193,N_2916,N_2905);
nor UO_194 (O_194,N_2992,N_2910);
xnor UO_195 (O_195,N_2992,N_2905);
and UO_196 (O_196,N_2965,N_2962);
nor UO_197 (O_197,N_2986,N_2942);
or UO_198 (O_198,N_2940,N_2992);
or UO_199 (O_199,N_2944,N_2950);
nand UO_200 (O_200,N_2951,N_2910);
or UO_201 (O_201,N_2933,N_2975);
nor UO_202 (O_202,N_2990,N_2976);
and UO_203 (O_203,N_2992,N_2924);
or UO_204 (O_204,N_2952,N_2976);
or UO_205 (O_205,N_2940,N_2980);
nand UO_206 (O_206,N_2995,N_2907);
or UO_207 (O_207,N_2943,N_2901);
nand UO_208 (O_208,N_2911,N_2960);
or UO_209 (O_209,N_2900,N_2999);
nand UO_210 (O_210,N_2976,N_2984);
nor UO_211 (O_211,N_2988,N_2900);
and UO_212 (O_212,N_2925,N_2964);
and UO_213 (O_213,N_2905,N_2945);
and UO_214 (O_214,N_2942,N_2978);
or UO_215 (O_215,N_2905,N_2980);
nor UO_216 (O_216,N_2945,N_2916);
and UO_217 (O_217,N_2901,N_2976);
and UO_218 (O_218,N_2929,N_2905);
or UO_219 (O_219,N_2912,N_2905);
nand UO_220 (O_220,N_2919,N_2950);
nor UO_221 (O_221,N_2932,N_2926);
or UO_222 (O_222,N_2998,N_2976);
and UO_223 (O_223,N_2957,N_2998);
and UO_224 (O_224,N_2939,N_2903);
or UO_225 (O_225,N_2940,N_2960);
nor UO_226 (O_226,N_2915,N_2974);
nor UO_227 (O_227,N_2932,N_2916);
or UO_228 (O_228,N_2942,N_2946);
nor UO_229 (O_229,N_2980,N_2951);
and UO_230 (O_230,N_2968,N_2917);
nor UO_231 (O_231,N_2937,N_2961);
and UO_232 (O_232,N_2942,N_2911);
nand UO_233 (O_233,N_2942,N_2943);
nand UO_234 (O_234,N_2961,N_2959);
nor UO_235 (O_235,N_2977,N_2981);
or UO_236 (O_236,N_2927,N_2952);
or UO_237 (O_237,N_2933,N_2940);
nor UO_238 (O_238,N_2900,N_2934);
or UO_239 (O_239,N_2913,N_2960);
nand UO_240 (O_240,N_2983,N_2900);
nand UO_241 (O_241,N_2979,N_2921);
nand UO_242 (O_242,N_2979,N_2903);
nor UO_243 (O_243,N_2958,N_2988);
nand UO_244 (O_244,N_2993,N_2945);
nor UO_245 (O_245,N_2952,N_2990);
nand UO_246 (O_246,N_2993,N_2990);
and UO_247 (O_247,N_2958,N_2965);
and UO_248 (O_248,N_2990,N_2973);
nor UO_249 (O_249,N_2915,N_2962);
and UO_250 (O_250,N_2934,N_2983);
nor UO_251 (O_251,N_2999,N_2958);
nand UO_252 (O_252,N_2957,N_2971);
nor UO_253 (O_253,N_2952,N_2931);
and UO_254 (O_254,N_2912,N_2948);
nand UO_255 (O_255,N_2970,N_2975);
nor UO_256 (O_256,N_2934,N_2992);
and UO_257 (O_257,N_2945,N_2951);
nor UO_258 (O_258,N_2948,N_2920);
nand UO_259 (O_259,N_2912,N_2953);
nor UO_260 (O_260,N_2939,N_2902);
and UO_261 (O_261,N_2902,N_2907);
or UO_262 (O_262,N_2946,N_2985);
nor UO_263 (O_263,N_2989,N_2956);
or UO_264 (O_264,N_2935,N_2936);
or UO_265 (O_265,N_2980,N_2957);
xor UO_266 (O_266,N_2929,N_2983);
nand UO_267 (O_267,N_2967,N_2951);
nor UO_268 (O_268,N_2990,N_2935);
nand UO_269 (O_269,N_2996,N_2967);
nor UO_270 (O_270,N_2948,N_2983);
or UO_271 (O_271,N_2900,N_2918);
and UO_272 (O_272,N_2995,N_2930);
nand UO_273 (O_273,N_2953,N_2974);
and UO_274 (O_274,N_2996,N_2940);
nand UO_275 (O_275,N_2971,N_2931);
and UO_276 (O_276,N_2982,N_2902);
nand UO_277 (O_277,N_2912,N_2977);
nand UO_278 (O_278,N_2977,N_2901);
nand UO_279 (O_279,N_2986,N_2934);
nand UO_280 (O_280,N_2961,N_2987);
nor UO_281 (O_281,N_2921,N_2922);
nand UO_282 (O_282,N_2913,N_2952);
or UO_283 (O_283,N_2974,N_2920);
and UO_284 (O_284,N_2977,N_2954);
nand UO_285 (O_285,N_2964,N_2937);
and UO_286 (O_286,N_2917,N_2958);
and UO_287 (O_287,N_2983,N_2903);
and UO_288 (O_288,N_2974,N_2999);
nand UO_289 (O_289,N_2940,N_2993);
nand UO_290 (O_290,N_2955,N_2950);
nand UO_291 (O_291,N_2940,N_2962);
and UO_292 (O_292,N_2930,N_2933);
nor UO_293 (O_293,N_2964,N_2995);
nor UO_294 (O_294,N_2966,N_2919);
or UO_295 (O_295,N_2917,N_2969);
and UO_296 (O_296,N_2996,N_2944);
or UO_297 (O_297,N_2953,N_2973);
nor UO_298 (O_298,N_2905,N_2968);
nand UO_299 (O_299,N_2991,N_2934);
nor UO_300 (O_300,N_2905,N_2943);
xnor UO_301 (O_301,N_2974,N_2964);
or UO_302 (O_302,N_2937,N_2996);
or UO_303 (O_303,N_2991,N_2986);
xnor UO_304 (O_304,N_2991,N_2911);
nand UO_305 (O_305,N_2945,N_2956);
nor UO_306 (O_306,N_2920,N_2913);
nor UO_307 (O_307,N_2986,N_2975);
nand UO_308 (O_308,N_2941,N_2908);
nor UO_309 (O_309,N_2975,N_2994);
and UO_310 (O_310,N_2980,N_2945);
and UO_311 (O_311,N_2945,N_2950);
nor UO_312 (O_312,N_2941,N_2951);
and UO_313 (O_313,N_2932,N_2953);
or UO_314 (O_314,N_2942,N_2976);
or UO_315 (O_315,N_2937,N_2906);
nand UO_316 (O_316,N_2914,N_2927);
nand UO_317 (O_317,N_2928,N_2927);
or UO_318 (O_318,N_2927,N_2954);
nor UO_319 (O_319,N_2989,N_2985);
and UO_320 (O_320,N_2959,N_2922);
nand UO_321 (O_321,N_2900,N_2920);
and UO_322 (O_322,N_2937,N_2967);
nand UO_323 (O_323,N_2993,N_2914);
nand UO_324 (O_324,N_2988,N_2940);
and UO_325 (O_325,N_2948,N_2915);
nor UO_326 (O_326,N_2935,N_2971);
and UO_327 (O_327,N_2930,N_2991);
or UO_328 (O_328,N_2954,N_2929);
or UO_329 (O_329,N_2944,N_2913);
or UO_330 (O_330,N_2998,N_2987);
nor UO_331 (O_331,N_2949,N_2906);
and UO_332 (O_332,N_2908,N_2918);
and UO_333 (O_333,N_2976,N_2915);
or UO_334 (O_334,N_2927,N_2953);
nand UO_335 (O_335,N_2912,N_2973);
nand UO_336 (O_336,N_2911,N_2969);
nand UO_337 (O_337,N_2999,N_2971);
or UO_338 (O_338,N_2902,N_2969);
nor UO_339 (O_339,N_2904,N_2932);
nand UO_340 (O_340,N_2957,N_2988);
and UO_341 (O_341,N_2945,N_2949);
or UO_342 (O_342,N_2949,N_2957);
nand UO_343 (O_343,N_2998,N_2963);
nand UO_344 (O_344,N_2973,N_2976);
and UO_345 (O_345,N_2960,N_2970);
nor UO_346 (O_346,N_2964,N_2931);
nand UO_347 (O_347,N_2974,N_2930);
and UO_348 (O_348,N_2909,N_2992);
and UO_349 (O_349,N_2920,N_2991);
nand UO_350 (O_350,N_2962,N_2944);
and UO_351 (O_351,N_2932,N_2962);
or UO_352 (O_352,N_2931,N_2944);
nor UO_353 (O_353,N_2983,N_2980);
nor UO_354 (O_354,N_2925,N_2917);
and UO_355 (O_355,N_2902,N_2956);
and UO_356 (O_356,N_2942,N_2933);
and UO_357 (O_357,N_2923,N_2903);
nand UO_358 (O_358,N_2910,N_2968);
nand UO_359 (O_359,N_2950,N_2986);
nor UO_360 (O_360,N_2952,N_2985);
or UO_361 (O_361,N_2942,N_2950);
nand UO_362 (O_362,N_2981,N_2915);
and UO_363 (O_363,N_2951,N_2984);
or UO_364 (O_364,N_2950,N_2952);
nand UO_365 (O_365,N_2918,N_2948);
nand UO_366 (O_366,N_2952,N_2935);
nand UO_367 (O_367,N_2984,N_2953);
nor UO_368 (O_368,N_2945,N_2907);
nand UO_369 (O_369,N_2969,N_2929);
and UO_370 (O_370,N_2963,N_2986);
nor UO_371 (O_371,N_2963,N_2910);
and UO_372 (O_372,N_2967,N_2957);
and UO_373 (O_373,N_2937,N_2965);
nand UO_374 (O_374,N_2900,N_2923);
and UO_375 (O_375,N_2974,N_2976);
and UO_376 (O_376,N_2956,N_2959);
and UO_377 (O_377,N_2918,N_2928);
nor UO_378 (O_378,N_2982,N_2923);
and UO_379 (O_379,N_2939,N_2979);
and UO_380 (O_380,N_2936,N_2975);
and UO_381 (O_381,N_2923,N_2942);
nand UO_382 (O_382,N_2985,N_2974);
or UO_383 (O_383,N_2962,N_2952);
and UO_384 (O_384,N_2902,N_2936);
or UO_385 (O_385,N_2978,N_2985);
and UO_386 (O_386,N_2914,N_2980);
or UO_387 (O_387,N_2978,N_2951);
nor UO_388 (O_388,N_2906,N_2941);
or UO_389 (O_389,N_2945,N_2979);
or UO_390 (O_390,N_2953,N_2997);
or UO_391 (O_391,N_2986,N_2965);
nor UO_392 (O_392,N_2906,N_2935);
nand UO_393 (O_393,N_2951,N_2985);
and UO_394 (O_394,N_2966,N_2967);
and UO_395 (O_395,N_2931,N_2999);
and UO_396 (O_396,N_2925,N_2940);
or UO_397 (O_397,N_2974,N_2907);
or UO_398 (O_398,N_2951,N_2999);
and UO_399 (O_399,N_2953,N_2937);
nand UO_400 (O_400,N_2933,N_2923);
nand UO_401 (O_401,N_2951,N_2994);
and UO_402 (O_402,N_2955,N_2918);
nand UO_403 (O_403,N_2982,N_2962);
nor UO_404 (O_404,N_2921,N_2983);
or UO_405 (O_405,N_2981,N_2906);
and UO_406 (O_406,N_2905,N_2959);
nand UO_407 (O_407,N_2939,N_2994);
nor UO_408 (O_408,N_2973,N_2911);
nor UO_409 (O_409,N_2972,N_2938);
or UO_410 (O_410,N_2920,N_2966);
or UO_411 (O_411,N_2969,N_2901);
and UO_412 (O_412,N_2925,N_2976);
and UO_413 (O_413,N_2976,N_2969);
or UO_414 (O_414,N_2964,N_2957);
nor UO_415 (O_415,N_2994,N_2960);
nand UO_416 (O_416,N_2934,N_2966);
or UO_417 (O_417,N_2900,N_2964);
nor UO_418 (O_418,N_2929,N_2903);
or UO_419 (O_419,N_2934,N_2940);
nand UO_420 (O_420,N_2942,N_2999);
and UO_421 (O_421,N_2938,N_2982);
nand UO_422 (O_422,N_2971,N_2914);
or UO_423 (O_423,N_2941,N_2922);
and UO_424 (O_424,N_2940,N_2913);
and UO_425 (O_425,N_2912,N_2930);
nor UO_426 (O_426,N_2916,N_2910);
and UO_427 (O_427,N_2961,N_2985);
nor UO_428 (O_428,N_2975,N_2914);
nand UO_429 (O_429,N_2971,N_2975);
nor UO_430 (O_430,N_2910,N_2918);
or UO_431 (O_431,N_2961,N_2935);
and UO_432 (O_432,N_2914,N_2942);
or UO_433 (O_433,N_2907,N_2930);
nand UO_434 (O_434,N_2900,N_2912);
or UO_435 (O_435,N_2982,N_2916);
or UO_436 (O_436,N_2961,N_2940);
nor UO_437 (O_437,N_2967,N_2986);
or UO_438 (O_438,N_2984,N_2959);
or UO_439 (O_439,N_2961,N_2962);
or UO_440 (O_440,N_2910,N_2945);
and UO_441 (O_441,N_2910,N_2975);
or UO_442 (O_442,N_2970,N_2910);
and UO_443 (O_443,N_2998,N_2947);
nor UO_444 (O_444,N_2923,N_2984);
nor UO_445 (O_445,N_2947,N_2912);
nor UO_446 (O_446,N_2913,N_2993);
or UO_447 (O_447,N_2946,N_2998);
and UO_448 (O_448,N_2951,N_2914);
and UO_449 (O_449,N_2920,N_2912);
nand UO_450 (O_450,N_2996,N_2911);
and UO_451 (O_451,N_2929,N_2930);
nor UO_452 (O_452,N_2974,N_2923);
or UO_453 (O_453,N_2958,N_2994);
or UO_454 (O_454,N_2911,N_2903);
xnor UO_455 (O_455,N_2933,N_2959);
nor UO_456 (O_456,N_2968,N_2990);
and UO_457 (O_457,N_2914,N_2921);
and UO_458 (O_458,N_2953,N_2962);
or UO_459 (O_459,N_2977,N_2925);
and UO_460 (O_460,N_2925,N_2954);
nand UO_461 (O_461,N_2912,N_2935);
or UO_462 (O_462,N_2977,N_2915);
and UO_463 (O_463,N_2940,N_2903);
nor UO_464 (O_464,N_2988,N_2956);
nor UO_465 (O_465,N_2977,N_2979);
nor UO_466 (O_466,N_2986,N_2995);
or UO_467 (O_467,N_2994,N_2914);
and UO_468 (O_468,N_2905,N_2933);
nor UO_469 (O_469,N_2931,N_2910);
and UO_470 (O_470,N_2962,N_2964);
or UO_471 (O_471,N_2941,N_2974);
or UO_472 (O_472,N_2993,N_2984);
and UO_473 (O_473,N_2956,N_2951);
and UO_474 (O_474,N_2926,N_2937);
nor UO_475 (O_475,N_2928,N_2952);
or UO_476 (O_476,N_2988,N_2970);
nor UO_477 (O_477,N_2908,N_2960);
and UO_478 (O_478,N_2987,N_2912);
or UO_479 (O_479,N_2917,N_2985);
or UO_480 (O_480,N_2968,N_2922);
nand UO_481 (O_481,N_2960,N_2945);
xnor UO_482 (O_482,N_2932,N_2965);
nor UO_483 (O_483,N_2950,N_2997);
or UO_484 (O_484,N_2974,N_2924);
or UO_485 (O_485,N_2956,N_2979);
nand UO_486 (O_486,N_2908,N_2931);
nor UO_487 (O_487,N_2950,N_2993);
or UO_488 (O_488,N_2950,N_2973);
or UO_489 (O_489,N_2939,N_2971);
and UO_490 (O_490,N_2962,N_2976);
nor UO_491 (O_491,N_2924,N_2914);
and UO_492 (O_492,N_2987,N_2970);
and UO_493 (O_493,N_2989,N_2938);
nor UO_494 (O_494,N_2961,N_2922);
nor UO_495 (O_495,N_2929,N_2968);
or UO_496 (O_496,N_2992,N_2970);
nor UO_497 (O_497,N_2908,N_2923);
nor UO_498 (O_498,N_2937,N_2963);
nand UO_499 (O_499,N_2937,N_2988);
endmodule