module basic_500_3000_500_3_levels_2xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_432,In_438);
nand U1 (N_1,In_41,In_365);
and U2 (N_2,In_418,In_214);
nand U3 (N_3,In_242,In_472);
or U4 (N_4,In_189,In_123);
and U5 (N_5,In_139,In_187);
or U6 (N_6,In_445,In_192);
and U7 (N_7,In_251,In_414);
nand U8 (N_8,In_106,In_57);
nand U9 (N_9,In_459,In_272);
and U10 (N_10,In_19,In_16);
or U11 (N_11,In_460,In_370);
nor U12 (N_12,In_380,In_399);
nor U13 (N_13,In_177,In_393);
or U14 (N_14,In_68,In_3);
nor U15 (N_15,In_250,In_437);
and U16 (N_16,In_9,In_496);
or U17 (N_17,In_311,In_264);
nor U18 (N_18,In_194,In_295);
and U19 (N_19,In_85,In_452);
nor U20 (N_20,In_153,In_353);
nor U21 (N_21,In_54,In_266);
nand U22 (N_22,In_36,In_231);
nand U23 (N_23,In_390,In_230);
or U24 (N_24,In_450,In_479);
or U25 (N_25,In_457,In_157);
or U26 (N_26,In_417,In_337);
or U27 (N_27,In_206,In_207);
and U28 (N_28,In_60,In_104);
and U29 (N_29,In_446,In_17);
nor U30 (N_30,In_132,In_70);
and U31 (N_31,In_391,In_292);
or U32 (N_32,In_345,In_50);
or U33 (N_33,In_78,In_39);
nand U34 (N_34,In_430,In_208);
and U35 (N_35,In_290,In_252);
nor U36 (N_36,In_4,In_127);
nor U37 (N_37,In_216,In_357);
and U38 (N_38,In_492,In_461);
or U39 (N_39,In_115,In_449);
or U40 (N_40,In_455,In_51);
nor U41 (N_41,In_424,In_49);
nor U42 (N_42,In_142,In_310);
and U43 (N_43,In_37,In_79);
or U44 (N_44,In_482,In_147);
nor U45 (N_45,In_302,In_98);
and U46 (N_46,In_0,In_340);
nor U47 (N_47,In_6,In_95);
nor U48 (N_48,In_465,In_176);
nor U49 (N_49,In_211,In_31);
or U50 (N_50,In_469,In_151);
nor U51 (N_51,In_277,In_169);
or U52 (N_52,In_373,In_369);
nor U53 (N_53,In_110,In_154);
nor U54 (N_54,In_382,In_166);
nand U55 (N_55,In_145,In_471);
nand U56 (N_56,In_81,In_174);
and U57 (N_57,In_210,In_124);
nor U58 (N_58,In_350,In_267);
nor U59 (N_59,In_234,In_218);
and U60 (N_60,In_140,In_35);
and U61 (N_61,In_69,In_25);
or U62 (N_62,In_338,In_90);
nor U63 (N_63,In_368,In_144);
nor U64 (N_64,In_263,In_243);
or U65 (N_65,In_120,In_395);
nand U66 (N_66,In_160,In_275);
nor U67 (N_67,In_329,In_15);
and U68 (N_68,In_423,In_257);
nand U69 (N_69,In_179,In_434);
and U70 (N_70,In_109,In_296);
nor U71 (N_71,In_255,In_273);
nand U72 (N_72,In_289,In_133);
or U73 (N_73,In_499,In_442);
nand U74 (N_74,In_235,In_413);
nor U75 (N_75,In_326,In_149);
nor U76 (N_76,In_222,In_258);
or U77 (N_77,In_347,In_197);
nor U78 (N_78,In_372,In_488);
nor U79 (N_79,In_462,In_485);
or U80 (N_80,In_265,In_431);
or U81 (N_81,In_301,In_116);
or U82 (N_82,In_335,In_362);
nand U83 (N_83,In_34,In_419);
xor U84 (N_84,In_356,In_383);
xnor U85 (N_85,In_220,In_375);
and U86 (N_86,In_240,In_40);
and U87 (N_87,In_91,In_236);
xnor U88 (N_88,In_405,In_199);
and U89 (N_89,In_312,In_108);
nand U90 (N_90,In_415,In_360);
and U91 (N_91,In_467,In_388);
or U92 (N_92,In_435,In_287);
nand U93 (N_93,In_72,In_241);
nor U94 (N_94,In_441,In_103);
nand U95 (N_95,In_336,In_215);
and U96 (N_96,In_165,In_361);
nand U97 (N_97,In_346,In_381);
nor U98 (N_98,In_233,In_268);
and U99 (N_99,In_408,In_409);
nor U100 (N_100,In_180,In_286);
nor U101 (N_101,In_254,In_88);
or U102 (N_102,In_294,In_89);
and U103 (N_103,In_293,In_348);
xor U104 (N_104,In_217,In_493);
or U105 (N_105,In_476,In_466);
nand U106 (N_106,In_196,In_280);
and U107 (N_107,In_107,In_66);
nor U108 (N_108,In_32,In_161);
nor U109 (N_109,In_158,In_453);
and U110 (N_110,In_315,In_478);
and U111 (N_111,In_397,In_253);
nor U112 (N_112,In_14,In_475);
and U113 (N_113,In_297,In_491);
nor U114 (N_114,In_170,In_93);
nand U115 (N_115,In_497,In_394);
and U116 (N_116,In_304,In_195);
nand U117 (N_117,In_178,In_205);
nor U118 (N_118,In_63,In_83);
nand U119 (N_119,In_26,In_44);
and U120 (N_120,In_184,In_392);
and U121 (N_121,In_237,In_30);
and U122 (N_122,In_136,In_288);
nand U123 (N_123,In_327,In_223);
xor U124 (N_124,In_378,In_135);
or U125 (N_125,In_244,In_247);
nand U126 (N_126,In_339,In_420);
and U127 (N_127,In_271,In_10);
and U128 (N_128,In_168,In_232);
or U129 (N_129,In_379,In_73);
nand U130 (N_130,In_384,In_96);
or U131 (N_131,In_358,In_62);
nor U132 (N_132,In_105,In_111);
nor U133 (N_133,In_422,In_480);
and U134 (N_134,In_219,In_52);
and U135 (N_135,In_427,In_55);
or U136 (N_136,In_410,In_470);
nand U137 (N_137,In_428,In_298);
or U138 (N_138,In_433,In_64);
or U139 (N_139,In_134,In_143);
xnor U140 (N_140,In_84,In_305);
nor U141 (N_141,In_8,In_316);
or U142 (N_142,In_76,In_342);
nor U143 (N_143,In_61,In_333);
or U144 (N_144,In_186,In_439);
or U145 (N_145,In_130,In_119);
and U146 (N_146,In_11,In_185);
nor U147 (N_147,In_53,In_406);
or U148 (N_148,In_43,In_213);
and U149 (N_149,In_22,In_454);
nor U150 (N_150,In_314,In_175);
nand U151 (N_151,In_285,In_278);
nor U152 (N_152,In_238,In_137);
nor U153 (N_153,In_308,In_65);
or U154 (N_154,In_448,In_239);
nand U155 (N_155,In_246,In_164);
nor U156 (N_156,In_1,In_171);
nand U157 (N_157,In_440,In_100);
or U158 (N_158,In_183,In_416);
and U159 (N_159,In_447,In_141);
or U160 (N_160,In_13,In_193);
nor U161 (N_161,In_283,In_221);
nand U162 (N_162,In_112,In_389);
or U163 (N_163,In_99,In_48);
nand U164 (N_164,In_92,In_421);
or U165 (N_165,In_398,In_458);
nor U166 (N_166,In_276,In_21);
nand U167 (N_167,In_269,In_411);
or U168 (N_168,In_279,In_260);
and U169 (N_169,In_114,In_354);
nor U170 (N_170,In_319,In_374);
or U171 (N_171,In_204,In_248);
nand U172 (N_172,In_259,In_443);
nand U173 (N_173,In_121,In_18);
xnor U174 (N_174,In_7,In_284);
nor U175 (N_175,In_494,In_261);
nor U176 (N_176,In_322,In_2);
and U177 (N_177,In_256,In_341);
or U178 (N_178,In_29,In_75);
and U179 (N_179,In_463,In_125);
and U180 (N_180,In_385,In_101);
xnor U181 (N_181,In_359,In_128);
nor U182 (N_182,In_274,In_307);
and U183 (N_183,In_377,In_456);
and U184 (N_184,In_23,In_182);
or U185 (N_185,In_403,In_489);
and U186 (N_186,In_152,In_159);
or U187 (N_187,In_483,In_364);
or U188 (N_188,In_225,In_226);
and U189 (N_189,In_396,In_270);
nand U190 (N_190,In_228,In_402);
nor U191 (N_191,In_343,In_118);
or U192 (N_192,In_464,In_202);
or U193 (N_193,In_27,In_400);
xnor U194 (N_194,In_407,In_404);
nand U195 (N_195,In_481,In_80);
nor U196 (N_196,In_321,In_209);
xnor U197 (N_197,In_371,In_74);
or U198 (N_198,In_97,In_386);
nor U199 (N_199,In_201,In_150);
nand U200 (N_200,In_58,In_498);
nand U201 (N_201,In_363,In_20);
nor U202 (N_202,In_33,In_46);
nor U203 (N_203,In_330,In_12);
nand U204 (N_204,In_200,In_425);
or U205 (N_205,In_87,In_146);
nor U206 (N_206,In_191,In_24);
and U207 (N_207,In_426,In_331);
and U208 (N_208,In_325,In_212);
nand U209 (N_209,In_300,In_67);
nor U210 (N_210,In_28,In_42);
nor U211 (N_211,In_156,In_203);
and U212 (N_212,In_282,In_291);
or U213 (N_213,In_167,In_306);
nor U214 (N_214,In_181,In_249);
or U215 (N_215,In_5,In_474);
nor U216 (N_216,In_173,In_412);
or U217 (N_217,In_303,In_495);
nand U218 (N_218,In_131,In_281);
nor U219 (N_219,In_401,In_487);
or U220 (N_220,In_436,In_320);
and U221 (N_221,In_313,In_56);
or U222 (N_222,In_148,In_86);
nor U223 (N_223,In_172,In_486);
nand U224 (N_224,In_82,In_245);
nand U225 (N_225,In_328,In_318);
nor U226 (N_226,In_198,In_323);
nand U227 (N_227,In_117,In_162);
nor U228 (N_228,In_45,In_224);
nor U229 (N_229,In_444,In_71);
and U230 (N_230,In_477,In_484);
nor U231 (N_231,In_332,In_102);
nor U232 (N_232,In_351,In_344);
nand U233 (N_233,In_367,In_129);
and U234 (N_234,In_334,In_155);
nand U235 (N_235,In_77,In_190);
or U236 (N_236,In_317,In_376);
xnor U237 (N_237,In_138,In_490);
nand U238 (N_238,In_355,In_38);
and U239 (N_239,In_429,In_366);
and U240 (N_240,In_262,In_188);
nor U241 (N_241,In_451,In_473);
nor U242 (N_242,In_59,In_126);
nand U243 (N_243,In_163,In_94);
or U244 (N_244,In_349,In_229);
or U245 (N_245,In_352,In_227);
nor U246 (N_246,In_113,In_122);
nor U247 (N_247,In_324,In_468);
or U248 (N_248,In_47,In_309);
and U249 (N_249,In_299,In_387);
and U250 (N_250,In_316,In_251);
or U251 (N_251,In_264,In_278);
nor U252 (N_252,In_272,In_16);
and U253 (N_253,In_202,In_494);
or U254 (N_254,In_167,In_260);
nor U255 (N_255,In_179,In_453);
and U256 (N_256,In_444,In_207);
nand U257 (N_257,In_130,In_84);
nand U258 (N_258,In_492,In_459);
nor U259 (N_259,In_490,In_13);
nand U260 (N_260,In_449,In_88);
nor U261 (N_261,In_73,In_478);
nor U262 (N_262,In_90,In_7);
nand U263 (N_263,In_150,In_277);
nand U264 (N_264,In_193,In_399);
and U265 (N_265,In_222,In_163);
or U266 (N_266,In_345,In_188);
nor U267 (N_267,In_351,In_154);
and U268 (N_268,In_216,In_450);
nand U269 (N_269,In_111,In_214);
nor U270 (N_270,In_1,In_299);
nor U271 (N_271,In_169,In_167);
or U272 (N_272,In_145,In_334);
or U273 (N_273,In_178,In_284);
nand U274 (N_274,In_466,In_391);
and U275 (N_275,In_333,In_202);
nand U276 (N_276,In_224,In_385);
nor U277 (N_277,In_50,In_28);
or U278 (N_278,In_458,In_293);
nand U279 (N_279,In_179,In_423);
or U280 (N_280,In_315,In_131);
nor U281 (N_281,In_25,In_283);
nand U282 (N_282,In_381,In_80);
and U283 (N_283,In_12,In_243);
nor U284 (N_284,In_240,In_187);
or U285 (N_285,In_214,In_305);
nand U286 (N_286,In_390,In_383);
nor U287 (N_287,In_146,In_454);
or U288 (N_288,In_423,In_145);
nor U289 (N_289,In_175,In_199);
nand U290 (N_290,In_173,In_275);
or U291 (N_291,In_60,In_436);
nand U292 (N_292,In_347,In_68);
nor U293 (N_293,In_236,In_128);
or U294 (N_294,In_432,In_140);
and U295 (N_295,In_35,In_397);
xor U296 (N_296,In_200,In_362);
nor U297 (N_297,In_319,In_268);
or U298 (N_298,In_471,In_253);
or U299 (N_299,In_268,In_30);
nand U300 (N_300,In_81,In_376);
or U301 (N_301,In_381,In_15);
and U302 (N_302,In_213,In_330);
nor U303 (N_303,In_305,In_385);
nand U304 (N_304,In_229,In_243);
and U305 (N_305,In_47,In_152);
or U306 (N_306,In_72,In_77);
nor U307 (N_307,In_69,In_236);
or U308 (N_308,In_288,In_372);
xnor U309 (N_309,In_164,In_251);
nand U310 (N_310,In_297,In_134);
or U311 (N_311,In_496,In_170);
nor U312 (N_312,In_34,In_458);
and U313 (N_313,In_426,In_403);
and U314 (N_314,In_408,In_223);
and U315 (N_315,In_172,In_168);
nor U316 (N_316,In_281,In_363);
and U317 (N_317,In_289,In_256);
or U318 (N_318,In_231,In_195);
and U319 (N_319,In_285,In_259);
and U320 (N_320,In_127,In_259);
nand U321 (N_321,In_200,In_33);
or U322 (N_322,In_434,In_158);
and U323 (N_323,In_282,In_312);
or U324 (N_324,In_356,In_282);
nor U325 (N_325,In_248,In_56);
nor U326 (N_326,In_445,In_146);
and U327 (N_327,In_320,In_350);
nand U328 (N_328,In_278,In_381);
nand U329 (N_329,In_223,In_65);
and U330 (N_330,In_114,In_397);
and U331 (N_331,In_2,In_85);
nor U332 (N_332,In_390,In_120);
xor U333 (N_333,In_139,In_13);
or U334 (N_334,In_37,In_162);
and U335 (N_335,In_245,In_415);
or U336 (N_336,In_27,In_132);
nor U337 (N_337,In_358,In_322);
xnor U338 (N_338,In_148,In_480);
nor U339 (N_339,In_338,In_181);
nor U340 (N_340,In_177,In_408);
nand U341 (N_341,In_273,In_225);
nor U342 (N_342,In_268,In_67);
and U343 (N_343,In_143,In_346);
nand U344 (N_344,In_243,In_234);
xor U345 (N_345,In_486,In_289);
and U346 (N_346,In_431,In_281);
or U347 (N_347,In_409,In_376);
and U348 (N_348,In_87,In_194);
nand U349 (N_349,In_397,In_294);
nor U350 (N_350,In_330,In_361);
or U351 (N_351,In_317,In_316);
nor U352 (N_352,In_21,In_361);
nand U353 (N_353,In_308,In_443);
xor U354 (N_354,In_125,In_461);
xor U355 (N_355,In_471,In_261);
nand U356 (N_356,In_266,In_376);
nand U357 (N_357,In_396,In_288);
and U358 (N_358,In_410,In_194);
or U359 (N_359,In_232,In_227);
and U360 (N_360,In_377,In_184);
nor U361 (N_361,In_257,In_331);
or U362 (N_362,In_494,In_169);
or U363 (N_363,In_479,In_274);
or U364 (N_364,In_494,In_465);
nor U365 (N_365,In_221,In_378);
nand U366 (N_366,In_47,In_371);
or U367 (N_367,In_129,In_120);
nor U368 (N_368,In_473,In_106);
and U369 (N_369,In_62,In_438);
and U370 (N_370,In_358,In_495);
nand U371 (N_371,In_241,In_283);
nand U372 (N_372,In_440,In_173);
nor U373 (N_373,In_251,In_105);
or U374 (N_374,In_480,In_372);
nor U375 (N_375,In_44,In_72);
nor U376 (N_376,In_424,In_356);
nand U377 (N_377,In_271,In_311);
nand U378 (N_378,In_284,In_444);
or U379 (N_379,In_456,In_141);
nand U380 (N_380,In_377,In_320);
and U381 (N_381,In_387,In_241);
and U382 (N_382,In_224,In_91);
nor U383 (N_383,In_282,In_244);
and U384 (N_384,In_489,In_419);
nand U385 (N_385,In_64,In_89);
and U386 (N_386,In_365,In_305);
or U387 (N_387,In_119,In_78);
nand U388 (N_388,In_364,In_262);
and U389 (N_389,In_462,In_228);
and U390 (N_390,In_214,In_11);
nand U391 (N_391,In_28,In_432);
nand U392 (N_392,In_425,In_272);
nor U393 (N_393,In_495,In_91);
nand U394 (N_394,In_203,In_341);
and U395 (N_395,In_370,In_83);
xnor U396 (N_396,In_446,In_49);
nand U397 (N_397,In_76,In_144);
or U398 (N_398,In_286,In_343);
nand U399 (N_399,In_405,In_168);
nand U400 (N_400,In_210,In_85);
nor U401 (N_401,In_425,In_185);
nand U402 (N_402,In_99,In_385);
or U403 (N_403,In_95,In_241);
and U404 (N_404,In_375,In_219);
and U405 (N_405,In_262,In_333);
and U406 (N_406,In_36,In_427);
or U407 (N_407,In_348,In_127);
nor U408 (N_408,In_366,In_113);
nand U409 (N_409,In_490,In_128);
or U410 (N_410,In_14,In_7);
nor U411 (N_411,In_94,In_209);
or U412 (N_412,In_312,In_21);
xor U413 (N_413,In_477,In_152);
nand U414 (N_414,In_405,In_155);
or U415 (N_415,In_179,In_216);
and U416 (N_416,In_443,In_314);
and U417 (N_417,In_433,In_240);
nor U418 (N_418,In_49,In_62);
or U419 (N_419,In_219,In_175);
or U420 (N_420,In_60,In_451);
and U421 (N_421,In_373,In_395);
or U422 (N_422,In_107,In_294);
or U423 (N_423,In_295,In_296);
nand U424 (N_424,In_193,In_112);
nand U425 (N_425,In_453,In_477);
or U426 (N_426,In_369,In_324);
nor U427 (N_427,In_307,In_19);
and U428 (N_428,In_220,In_402);
and U429 (N_429,In_460,In_8);
or U430 (N_430,In_406,In_122);
nor U431 (N_431,In_399,In_382);
nand U432 (N_432,In_39,In_182);
and U433 (N_433,In_97,In_438);
and U434 (N_434,In_443,In_214);
nor U435 (N_435,In_230,In_2);
nand U436 (N_436,In_129,In_306);
or U437 (N_437,In_276,In_19);
and U438 (N_438,In_208,In_56);
nor U439 (N_439,In_449,In_445);
and U440 (N_440,In_349,In_494);
xor U441 (N_441,In_263,In_122);
nor U442 (N_442,In_158,In_391);
or U443 (N_443,In_197,In_28);
and U444 (N_444,In_345,In_71);
nor U445 (N_445,In_79,In_231);
and U446 (N_446,In_358,In_184);
nor U447 (N_447,In_85,In_248);
and U448 (N_448,In_198,In_159);
nand U449 (N_449,In_254,In_499);
nand U450 (N_450,In_200,In_171);
and U451 (N_451,In_484,In_206);
nand U452 (N_452,In_14,In_227);
nand U453 (N_453,In_396,In_255);
and U454 (N_454,In_437,In_239);
nand U455 (N_455,In_96,In_294);
xnor U456 (N_456,In_301,In_401);
or U457 (N_457,In_244,In_236);
nor U458 (N_458,In_389,In_404);
or U459 (N_459,In_240,In_194);
nand U460 (N_460,In_80,In_256);
nor U461 (N_461,In_79,In_24);
nand U462 (N_462,In_220,In_321);
nor U463 (N_463,In_44,In_301);
nand U464 (N_464,In_102,In_392);
nor U465 (N_465,In_210,In_477);
and U466 (N_466,In_307,In_222);
nor U467 (N_467,In_77,In_497);
nor U468 (N_468,In_16,In_108);
nor U469 (N_469,In_451,In_496);
and U470 (N_470,In_277,In_485);
nand U471 (N_471,In_357,In_187);
nor U472 (N_472,In_123,In_21);
nand U473 (N_473,In_484,In_81);
or U474 (N_474,In_358,In_262);
nand U475 (N_475,In_391,In_26);
nand U476 (N_476,In_126,In_20);
and U477 (N_477,In_99,In_175);
and U478 (N_478,In_103,In_329);
and U479 (N_479,In_265,In_449);
and U480 (N_480,In_434,In_42);
or U481 (N_481,In_87,In_16);
nor U482 (N_482,In_40,In_50);
nor U483 (N_483,In_482,In_67);
or U484 (N_484,In_109,In_374);
nand U485 (N_485,In_301,In_54);
nor U486 (N_486,In_414,In_188);
nand U487 (N_487,In_248,In_452);
nor U488 (N_488,In_244,In_418);
nand U489 (N_489,In_290,In_93);
or U490 (N_490,In_91,In_362);
nand U491 (N_491,In_297,In_91);
nand U492 (N_492,In_252,In_440);
nand U493 (N_493,In_480,In_16);
or U494 (N_494,In_14,In_48);
or U495 (N_495,In_262,In_23);
or U496 (N_496,In_171,In_27);
nand U497 (N_497,In_302,In_119);
or U498 (N_498,In_391,In_123);
or U499 (N_499,In_357,In_470);
or U500 (N_500,In_100,In_318);
nor U501 (N_501,In_487,In_50);
or U502 (N_502,In_359,In_22);
nand U503 (N_503,In_313,In_495);
xor U504 (N_504,In_34,In_486);
nor U505 (N_505,In_187,In_138);
or U506 (N_506,In_21,In_60);
nor U507 (N_507,In_94,In_64);
nor U508 (N_508,In_92,In_475);
or U509 (N_509,In_414,In_374);
and U510 (N_510,In_32,In_497);
nand U511 (N_511,In_417,In_106);
and U512 (N_512,In_199,In_115);
or U513 (N_513,In_397,In_132);
or U514 (N_514,In_319,In_353);
nor U515 (N_515,In_281,In_261);
and U516 (N_516,In_141,In_290);
or U517 (N_517,In_224,In_336);
nand U518 (N_518,In_99,In_29);
nor U519 (N_519,In_38,In_88);
nand U520 (N_520,In_293,In_254);
nand U521 (N_521,In_283,In_273);
and U522 (N_522,In_190,In_54);
nor U523 (N_523,In_259,In_453);
nor U524 (N_524,In_17,In_474);
nand U525 (N_525,In_49,In_276);
nand U526 (N_526,In_334,In_395);
nand U527 (N_527,In_433,In_378);
and U528 (N_528,In_225,In_90);
nand U529 (N_529,In_463,In_409);
or U530 (N_530,In_307,In_167);
nand U531 (N_531,In_326,In_143);
or U532 (N_532,In_252,In_267);
nor U533 (N_533,In_490,In_127);
nor U534 (N_534,In_199,In_141);
nor U535 (N_535,In_466,In_70);
or U536 (N_536,In_261,In_56);
or U537 (N_537,In_27,In_298);
xnor U538 (N_538,In_314,In_33);
or U539 (N_539,In_252,In_282);
nor U540 (N_540,In_307,In_83);
or U541 (N_541,In_335,In_152);
nand U542 (N_542,In_178,In_415);
nand U543 (N_543,In_85,In_405);
and U544 (N_544,In_332,In_471);
nor U545 (N_545,In_411,In_494);
nand U546 (N_546,In_247,In_56);
nor U547 (N_547,In_193,In_392);
or U548 (N_548,In_378,In_356);
nand U549 (N_549,In_104,In_333);
nor U550 (N_550,In_232,In_253);
and U551 (N_551,In_379,In_350);
nor U552 (N_552,In_413,In_391);
and U553 (N_553,In_128,In_225);
nand U554 (N_554,In_344,In_159);
nor U555 (N_555,In_131,In_356);
nand U556 (N_556,In_316,In_159);
nor U557 (N_557,In_47,In_122);
nand U558 (N_558,In_87,In_406);
or U559 (N_559,In_328,In_166);
nor U560 (N_560,In_145,In_476);
nand U561 (N_561,In_129,In_485);
or U562 (N_562,In_393,In_90);
nor U563 (N_563,In_162,In_98);
nand U564 (N_564,In_322,In_119);
nand U565 (N_565,In_317,In_408);
and U566 (N_566,In_315,In_278);
and U567 (N_567,In_435,In_358);
nand U568 (N_568,In_433,In_110);
and U569 (N_569,In_303,In_322);
or U570 (N_570,In_185,In_141);
nor U571 (N_571,In_32,In_448);
nor U572 (N_572,In_72,In_284);
or U573 (N_573,In_257,In_448);
nor U574 (N_574,In_429,In_497);
nor U575 (N_575,In_300,In_240);
or U576 (N_576,In_59,In_318);
and U577 (N_577,In_31,In_229);
nor U578 (N_578,In_441,In_350);
nor U579 (N_579,In_291,In_134);
nor U580 (N_580,In_78,In_201);
or U581 (N_581,In_68,In_486);
nor U582 (N_582,In_365,In_235);
or U583 (N_583,In_362,In_482);
nor U584 (N_584,In_474,In_483);
nor U585 (N_585,In_424,In_170);
nor U586 (N_586,In_485,In_272);
nand U587 (N_587,In_455,In_230);
or U588 (N_588,In_195,In_447);
or U589 (N_589,In_80,In_442);
nor U590 (N_590,In_356,In_69);
nand U591 (N_591,In_229,In_225);
or U592 (N_592,In_484,In_195);
nor U593 (N_593,In_342,In_230);
nor U594 (N_594,In_323,In_468);
and U595 (N_595,In_27,In_333);
and U596 (N_596,In_84,In_423);
nand U597 (N_597,In_196,In_99);
or U598 (N_598,In_351,In_392);
nor U599 (N_599,In_58,In_67);
or U600 (N_600,In_80,In_54);
nor U601 (N_601,In_276,In_450);
nand U602 (N_602,In_84,In_253);
nor U603 (N_603,In_486,In_214);
nand U604 (N_604,In_27,In_477);
and U605 (N_605,In_227,In_5);
nand U606 (N_606,In_253,In_7);
or U607 (N_607,In_71,In_332);
nand U608 (N_608,In_482,In_279);
nor U609 (N_609,In_28,In_54);
or U610 (N_610,In_65,In_304);
nor U611 (N_611,In_76,In_307);
or U612 (N_612,In_423,In_455);
and U613 (N_613,In_383,In_161);
and U614 (N_614,In_292,In_329);
or U615 (N_615,In_138,In_336);
or U616 (N_616,In_250,In_20);
nand U617 (N_617,In_32,In_109);
or U618 (N_618,In_148,In_486);
or U619 (N_619,In_290,In_287);
nand U620 (N_620,In_445,In_480);
nand U621 (N_621,In_357,In_481);
nand U622 (N_622,In_200,In_90);
nand U623 (N_623,In_311,In_284);
or U624 (N_624,In_423,In_85);
or U625 (N_625,In_298,In_24);
nand U626 (N_626,In_149,In_385);
nor U627 (N_627,In_418,In_20);
or U628 (N_628,In_242,In_18);
xor U629 (N_629,In_497,In_125);
or U630 (N_630,In_464,In_204);
nor U631 (N_631,In_436,In_255);
nand U632 (N_632,In_120,In_293);
and U633 (N_633,In_65,In_395);
nand U634 (N_634,In_69,In_321);
nor U635 (N_635,In_247,In_79);
nor U636 (N_636,In_464,In_212);
xnor U637 (N_637,In_111,In_209);
and U638 (N_638,In_64,In_476);
nor U639 (N_639,In_175,In_88);
nand U640 (N_640,In_420,In_442);
nor U641 (N_641,In_434,In_233);
nor U642 (N_642,In_418,In_14);
or U643 (N_643,In_195,In_308);
and U644 (N_644,In_231,In_158);
and U645 (N_645,In_142,In_442);
nor U646 (N_646,In_408,In_27);
and U647 (N_647,In_344,In_95);
and U648 (N_648,In_205,In_69);
or U649 (N_649,In_348,In_414);
and U650 (N_650,In_362,In_128);
and U651 (N_651,In_453,In_363);
and U652 (N_652,In_212,In_347);
or U653 (N_653,In_121,In_328);
and U654 (N_654,In_140,In_224);
and U655 (N_655,In_151,In_201);
nand U656 (N_656,In_485,In_203);
nor U657 (N_657,In_324,In_20);
nor U658 (N_658,In_90,In_31);
nand U659 (N_659,In_493,In_85);
nor U660 (N_660,In_316,In_286);
nor U661 (N_661,In_35,In_52);
xnor U662 (N_662,In_225,In_411);
xor U663 (N_663,In_390,In_331);
nand U664 (N_664,In_48,In_282);
or U665 (N_665,In_493,In_441);
nor U666 (N_666,In_368,In_349);
and U667 (N_667,In_398,In_15);
nand U668 (N_668,In_407,In_147);
nand U669 (N_669,In_369,In_366);
and U670 (N_670,In_234,In_188);
or U671 (N_671,In_444,In_497);
or U672 (N_672,In_1,In_434);
and U673 (N_673,In_295,In_418);
and U674 (N_674,In_123,In_475);
and U675 (N_675,In_185,In_100);
nor U676 (N_676,In_420,In_460);
and U677 (N_677,In_134,In_160);
nand U678 (N_678,In_34,In_386);
and U679 (N_679,In_433,In_390);
nand U680 (N_680,In_211,In_397);
nor U681 (N_681,In_19,In_113);
or U682 (N_682,In_371,In_298);
nor U683 (N_683,In_136,In_459);
nor U684 (N_684,In_451,In_340);
nor U685 (N_685,In_289,In_6);
nor U686 (N_686,In_47,In_494);
nand U687 (N_687,In_254,In_185);
and U688 (N_688,In_192,In_100);
nand U689 (N_689,In_145,In_417);
xnor U690 (N_690,In_209,In_87);
nand U691 (N_691,In_451,In_336);
and U692 (N_692,In_189,In_385);
nor U693 (N_693,In_218,In_118);
and U694 (N_694,In_336,In_452);
nand U695 (N_695,In_323,In_199);
nand U696 (N_696,In_224,In_392);
and U697 (N_697,In_215,In_45);
nand U698 (N_698,In_240,In_403);
or U699 (N_699,In_369,In_207);
nand U700 (N_700,In_135,In_353);
and U701 (N_701,In_345,In_142);
and U702 (N_702,In_486,In_496);
and U703 (N_703,In_168,In_307);
nand U704 (N_704,In_461,In_262);
or U705 (N_705,In_108,In_0);
and U706 (N_706,In_115,In_84);
or U707 (N_707,In_24,In_384);
nor U708 (N_708,In_268,In_181);
nand U709 (N_709,In_277,In_305);
nor U710 (N_710,In_370,In_223);
or U711 (N_711,In_445,In_28);
or U712 (N_712,In_263,In_415);
and U713 (N_713,In_477,In_267);
and U714 (N_714,In_158,In_16);
nand U715 (N_715,In_210,In_499);
or U716 (N_716,In_252,In_498);
nand U717 (N_717,In_286,In_125);
nor U718 (N_718,In_273,In_256);
and U719 (N_719,In_366,In_285);
xnor U720 (N_720,In_291,In_447);
and U721 (N_721,In_285,In_205);
nand U722 (N_722,In_313,In_477);
nand U723 (N_723,In_456,In_363);
or U724 (N_724,In_245,In_26);
and U725 (N_725,In_341,In_60);
nand U726 (N_726,In_368,In_156);
and U727 (N_727,In_423,In_493);
nor U728 (N_728,In_88,In_339);
nor U729 (N_729,In_497,In_11);
or U730 (N_730,In_362,In_386);
nor U731 (N_731,In_316,In_413);
or U732 (N_732,In_335,In_166);
or U733 (N_733,In_23,In_114);
nand U734 (N_734,In_5,In_222);
nor U735 (N_735,In_365,In_58);
nor U736 (N_736,In_358,In_101);
and U737 (N_737,In_68,In_16);
or U738 (N_738,In_91,In_51);
and U739 (N_739,In_49,In_392);
nand U740 (N_740,In_226,In_372);
and U741 (N_741,In_156,In_344);
nand U742 (N_742,In_409,In_153);
nand U743 (N_743,In_448,In_177);
nand U744 (N_744,In_176,In_483);
nand U745 (N_745,In_310,In_269);
nand U746 (N_746,In_471,In_405);
and U747 (N_747,In_458,In_40);
nor U748 (N_748,In_35,In_33);
nor U749 (N_749,In_216,In_156);
nand U750 (N_750,In_434,In_480);
or U751 (N_751,In_180,In_236);
or U752 (N_752,In_406,In_486);
nor U753 (N_753,In_63,In_27);
or U754 (N_754,In_311,In_329);
nor U755 (N_755,In_65,In_366);
or U756 (N_756,In_476,In_69);
nand U757 (N_757,In_294,In_226);
nor U758 (N_758,In_142,In_17);
and U759 (N_759,In_91,In_49);
and U760 (N_760,In_164,In_475);
nand U761 (N_761,In_174,In_69);
or U762 (N_762,In_326,In_415);
nor U763 (N_763,In_284,In_411);
nor U764 (N_764,In_333,In_354);
nor U765 (N_765,In_104,In_178);
and U766 (N_766,In_476,In_61);
or U767 (N_767,In_275,In_394);
nand U768 (N_768,In_442,In_186);
nor U769 (N_769,In_45,In_390);
nand U770 (N_770,In_7,In_134);
and U771 (N_771,In_62,In_432);
and U772 (N_772,In_364,In_245);
and U773 (N_773,In_181,In_202);
nor U774 (N_774,In_299,In_156);
nor U775 (N_775,In_497,In_24);
or U776 (N_776,In_353,In_7);
nor U777 (N_777,In_341,In_180);
or U778 (N_778,In_423,In_262);
nand U779 (N_779,In_377,In_251);
or U780 (N_780,In_456,In_21);
nor U781 (N_781,In_104,In_259);
nor U782 (N_782,In_407,In_316);
and U783 (N_783,In_150,In_272);
nor U784 (N_784,In_332,In_177);
nand U785 (N_785,In_308,In_354);
and U786 (N_786,In_283,In_312);
xor U787 (N_787,In_64,In_179);
nand U788 (N_788,In_434,In_222);
and U789 (N_789,In_484,In_412);
or U790 (N_790,In_452,In_294);
nand U791 (N_791,In_120,In_434);
or U792 (N_792,In_355,In_82);
or U793 (N_793,In_131,In_115);
or U794 (N_794,In_397,In_28);
nor U795 (N_795,In_123,In_416);
or U796 (N_796,In_347,In_460);
xnor U797 (N_797,In_461,In_494);
nand U798 (N_798,In_315,In_45);
and U799 (N_799,In_132,In_206);
and U800 (N_800,In_154,In_451);
or U801 (N_801,In_229,In_232);
or U802 (N_802,In_492,In_85);
or U803 (N_803,In_27,In_62);
nand U804 (N_804,In_307,In_297);
nor U805 (N_805,In_49,In_335);
nand U806 (N_806,In_402,In_13);
nor U807 (N_807,In_145,In_303);
nand U808 (N_808,In_19,In_152);
and U809 (N_809,In_143,In_464);
and U810 (N_810,In_334,In_433);
or U811 (N_811,In_336,In_49);
or U812 (N_812,In_484,In_60);
and U813 (N_813,In_325,In_24);
nor U814 (N_814,In_248,In_201);
nand U815 (N_815,In_150,In_461);
nand U816 (N_816,In_448,In_169);
and U817 (N_817,In_207,In_368);
nand U818 (N_818,In_180,In_287);
nor U819 (N_819,In_316,In_90);
nor U820 (N_820,In_214,In_166);
and U821 (N_821,In_36,In_73);
and U822 (N_822,In_20,In_291);
or U823 (N_823,In_19,In_281);
xnor U824 (N_824,In_98,In_400);
nand U825 (N_825,In_244,In_35);
or U826 (N_826,In_282,In_190);
or U827 (N_827,In_86,In_74);
and U828 (N_828,In_4,In_314);
or U829 (N_829,In_21,In_173);
xor U830 (N_830,In_107,In_237);
nand U831 (N_831,In_342,In_316);
nor U832 (N_832,In_271,In_482);
or U833 (N_833,In_295,In_291);
nand U834 (N_834,In_72,In_43);
or U835 (N_835,In_351,In_329);
or U836 (N_836,In_27,In_265);
and U837 (N_837,In_395,In_67);
nand U838 (N_838,In_134,In_217);
and U839 (N_839,In_364,In_210);
nand U840 (N_840,In_399,In_307);
nand U841 (N_841,In_4,In_424);
nand U842 (N_842,In_317,In_382);
and U843 (N_843,In_391,In_183);
or U844 (N_844,In_2,In_480);
nor U845 (N_845,In_487,In_464);
and U846 (N_846,In_108,In_444);
nand U847 (N_847,In_469,In_240);
nand U848 (N_848,In_364,In_440);
and U849 (N_849,In_290,In_60);
and U850 (N_850,In_384,In_332);
or U851 (N_851,In_142,In_490);
nand U852 (N_852,In_197,In_392);
nand U853 (N_853,In_240,In_4);
nand U854 (N_854,In_201,In_174);
or U855 (N_855,In_202,In_200);
nor U856 (N_856,In_441,In_252);
or U857 (N_857,In_137,In_485);
or U858 (N_858,In_127,In_124);
nor U859 (N_859,In_371,In_53);
xnor U860 (N_860,In_221,In_403);
xor U861 (N_861,In_304,In_288);
nand U862 (N_862,In_61,In_339);
nand U863 (N_863,In_266,In_336);
and U864 (N_864,In_137,In_117);
xor U865 (N_865,In_182,In_362);
or U866 (N_866,In_442,In_280);
and U867 (N_867,In_289,In_17);
and U868 (N_868,In_197,In_337);
and U869 (N_869,In_292,In_148);
and U870 (N_870,In_241,In_29);
nand U871 (N_871,In_211,In_68);
and U872 (N_872,In_79,In_62);
nand U873 (N_873,In_355,In_9);
nor U874 (N_874,In_434,In_460);
and U875 (N_875,In_388,In_51);
or U876 (N_876,In_383,In_190);
nor U877 (N_877,In_283,In_465);
or U878 (N_878,In_106,In_327);
xnor U879 (N_879,In_282,In_102);
or U880 (N_880,In_293,In_305);
or U881 (N_881,In_390,In_480);
xnor U882 (N_882,In_327,In_42);
and U883 (N_883,In_227,In_491);
or U884 (N_884,In_114,In_96);
and U885 (N_885,In_306,In_208);
nor U886 (N_886,In_129,In_138);
nand U887 (N_887,In_372,In_240);
or U888 (N_888,In_353,In_305);
and U889 (N_889,In_102,In_162);
nor U890 (N_890,In_449,In_462);
or U891 (N_891,In_349,In_52);
and U892 (N_892,In_438,In_275);
nand U893 (N_893,In_285,In_313);
and U894 (N_894,In_131,In_302);
nor U895 (N_895,In_157,In_461);
or U896 (N_896,In_417,In_406);
and U897 (N_897,In_417,In_161);
nand U898 (N_898,In_284,In_362);
and U899 (N_899,In_227,In_351);
nand U900 (N_900,In_347,In_477);
nor U901 (N_901,In_79,In_344);
nor U902 (N_902,In_330,In_338);
and U903 (N_903,In_64,In_222);
nand U904 (N_904,In_284,In_115);
nor U905 (N_905,In_242,In_231);
or U906 (N_906,In_224,In_221);
nand U907 (N_907,In_39,In_488);
nand U908 (N_908,In_48,In_167);
nor U909 (N_909,In_119,In_38);
and U910 (N_910,In_71,In_124);
nand U911 (N_911,In_301,In_435);
nor U912 (N_912,In_5,In_373);
and U913 (N_913,In_438,In_436);
nor U914 (N_914,In_112,In_36);
and U915 (N_915,In_117,In_216);
and U916 (N_916,In_326,In_202);
or U917 (N_917,In_137,In_71);
and U918 (N_918,In_118,In_93);
and U919 (N_919,In_326,In_330);
nand U920 (N_920,In_57,In_343);
nor U921 (N_921,In_159,In_277);
nor U922 (N_922,In_239,In_410);
nand U923 (N_923,In_398,In_320);
or U924 (N_924,In_213,In_472);
nand U925 (N_925,In_440,In_315);
or U926 (N_926,In_233,In_461);
nor U927 (N_927,In_181,In_259);
nand U928 (N_928,In_217,In_499);
and U929 (N_929,In_268,In_362);
nor U930 (N_930,In_101,In_263);
nor U931 (N_931,In_123,In_472);
nor U932 (N_932,In_487,In_283);
nand U933 (N_933,In_92,In_461);
or U934 (N_934,In_335,In_135);
and U935 (N_935,In_471,In_429);
nor U936 (N_936,In_208,In_158);
and U937 (N_937,In_5,In_381);
or U938 (N_938,In_327,In_384);
nand U939 (N_939,In_434,In_196);
or U940 (N_940,In_461,In_329);
and U941 (N_941,In_483,In_473);
nand U942 (N_942,In_402,In_481);
nor U943 (N_943,In_142,In_267);
and U944 (N_944,In_492,In_491);
nand U945 (N_945,In_202,In_474);
or U946 (N_946,In_55,In_421);
nor U947 (N_947,In_419,In_238);
nand U948 (N_948,In_100,In_95);
or U949 (N_949,In_278,In_493);
nand U950 (N_950,In_31,In_475);
or U951 (N_951,In_168,In_355);
or U952 (N_952,In_466,In_356);
nand U953 (N_953,In_54,In_460);
and U954 (N_954,In_221,In_293);
and U955 (N_955,In_272,In_301);
nor U956 (N_956,In_61,In_64);
nor U957 (N_957,In_442,In_349);
nor U958 (N_958,In_484,In_73);
nor U959 (N_959,In_388,In_272);
nand U960 (N_960,In_174,In_349);
nand U961 (N_961,In_448,In_443);
nand U962 (N_962,In_296,In_357);
or U963 (N_963,In_96,In_155);
nor U964 (N_964,In_379,In_293);
nor U965 (N_965,In_158,In_413);
nand U966 (N_966,In_48,In_215);
and U967 (N_967,In_378,In_58);
nand U968 (N_968,In_408,In_11);
nor U969 (N_969,In_94,In_152);
and U970 (N_970,In_104,In_332);
or U971 (N_971,In_317,In_86);
nor U972 (N_972,In_118,In_385);
or U973 (N_973,In_177,In_63);
or U974 (N_974,In_477,In_206);
nor U975 (N_975,In_449,In_441);
or U976 (N_976,In_310,In_258);
or U977 (N_977,In_262,In_493);
nor U978 (N_978,In_465,In_71);
nor U979 (N_979,In_434,In_368);
or U980 (N_980,In_130,In_476);
and U981 (N_981,In_72,In_374);
nor U982 (N_982,In_267,In_182);
xor U983 (N_983,In_372,In_117);
nor U984 (N_984,In_75,In_272);
nor U985 (N_985,In_188,In_121);
nor U986 (N_986,In_197,In_499);
and U987 (N_987,In_97,In_67);
or U988 (N_988,In_303,In_319);
or U989 (N_989,In_82,In_227);
xor U990 (N_990,In_496,In_339);
and U991 (N_991,In_450,In_21);
nand U992 (N_992,In_164,In_54);
or U993 (N_993,In_32,In_42);
nand U994 (N_994,In_491,In_145);
nor U995 (N_995,In_322,In_380);
nor U996 (N_996,In_279,In_197);
nand U997 (N_997,In_45,In_325);
or U998 (N_998,In_73,In_350);
nand U999 (N_999,In_483,In_281);
or U1000 (N_1000,N_380,N_456);
nor U1001 (N_1001,N_269,N_83);
xnor U1002 (N_1002,N_849,N_404);
nand U1003 (N_1003,N_288,N_9);
nand U1004 (N_1004,N_785,N_876);
nor U1005 (N_1005,N_656,N_295);
nor U1006 (N_1006,N_208,N_893);
nand U1007 (N_1007,N_706,N_709);
nor U1008 (N_1008,N_987,N_58);
or U1009 (N_1009,N_17,N_582);
nand U1010 (N_1010,N_971,N_408);
nand U1011 (N_1011,N_702,N_133);
nor U1012 (N_1012,N_439,N_6);
nor U1013 (N_1013,N_914,N_34);
or U1014 (N_1014,N_326,N_529);
nand U1015 (N_1015,N_222,N_743);
nand U1016 (N_1016,N_826,N_153);
xor U1017 (N_1017,N_511,N_619);
nor U1018 (N_1018,N_409,N_719);
and U1019 (N_1019,N_866,N_349);
xor U1020 (N_1020,N_367,N_148);
nor U1021 (N_1021,N_694,N_990);
or U1022 (N_1022,N_431,N_125);
nand U1023 (N_1023,N_338,N_909);
and U1024 (N_1024,N_804,N_200);
and U1025 (N_1025,N_924,N_545);
nand U1026 (N_1026,N_438,N_926);
and U1027 (N_1027,N_220,N_811);
or U1028 (N_1028,N_616,N_848);
and U1029 (N_1029,N_972,N_746);
or U1030 (N_1030,N_318,N_834);
and U1031 (N_1031,N_855,N_308);
and U1032 (N_1032,N_37,N_24);
or U1033 (N_1033,N_809,N_937);
nand U1034 (N_1034,N_859,N_920);
or U1035 (N_1035,N_142,N_68);
nand U1036 (N_1036,N_624,N_444);
and U1037 (N_1037,N_400,N_391);
or U1038 (N_1038,N_896,N_490);
or U1039 (N_1039,N_108,N_340);
and U1040 (N_1040,N_417,N_503);
nor U1041 (N_1041,N_366,N_573);
and U1042 (N_1042,N_377,N_451);
nor U1043 (N_1043,N_690,N_369);
nor U1044 (N_1044,N_865,N_662);
nand U1045 (N_1045,N_742,N_492);
and U1046 (N_1046,N_356,N_164);
nand U1047 (N_1047,N_21,N_201);
nor U1048 (N_1048,N_922,N_415);
or U1049 (N_1049,N_891,N_176);
xnor U1050 (N_1050,N_633,N_317);
nand U1051 (N_1051,N_885,N_405);
nand U1052 (N_1052,N_685,N_111);
nor U1053 (N_1053,N_594,N_911);
nand U1054 (N_1054,N_463,N_549);
nor U1055 (N_1055,N_723,N_512);
and U1056 (N_1056,N_651,N_628);
or U1057 (N_1057,N_652,N_337);
nor U1058 (N_1058,N_581,N_315);
or U1059 (N_1059,N_999,N_192);
nand U1060 (N_1060,N_850,N_245);
or U1061 (N_1061,N_583,N_740);
and U1062 (N_1062,N_818,N_484);
nor U1063 (N_1063,N_908,N_830);
and U1064 (N_1064,N_683,N_657);
and U1065 (N_1065,N_151,N_851);
nand U1066 (N_1066,N_258,N_72);
nor U1067 (N_1067,N_278,N_747);
nor U1068 (N_1068,N_152,N_535);
or U1069 (N_1069,N_137,N_761);
or U1070 (N_1070,N_135,N_732);
nor U1071 (N_1071,N_96,N_344);
nand U1072 (N_1072,N_156,N_140);
nand U1073 (N_1073,N_973,N_109);
nand U1074 (N_1074,N_399,N_584);
or U1075 (N_1075,N_61,N_564);
nor U1076 (N_1076,N_212,N_940);
nand U1077 (N_1077,N_286,N_620);
or U1078 (N_1078,N_262,N_472);
and U1079 (N_1079,N_780,N_729);
nor U1080 (N_1080,N_884,N_668);
nor U1081 (N_1081,N_725,N_560);
and U1082 (N_1082,N_892,N_976);
and U1083 (N_1083,N_321,N_167);
nand U1084 (N_1084,N_27,N_632);
nand U1085 (N_1085,N_32,N_146);
and U1086 (N_1086,N_749,N_733);
nor U1087 (N_1087,N_226,N_939);
or U1088 (N_1088,N_697,N_888);
or U1089 (N_1089,N_460,N_99);
or U1090 (N_1090,N_559,N_397);
nor U1091 (N_1091,N_4,N_664);
and U1092 (N_1092,N_555,N_424);
and U1093 (N_1093,N_756,N_57);
and U1094 (N_1094,N_227,N_778);
and U1095 (N_1095,N_952,N_777);
nand U1096 (N_1096,N_87,N_485);
or U1097 (N_1097,N_810,N_275);
or U1098 (N_1098,N_602,N_630);
or U1099 (N_1099,N_607,N_667);
or U1100 (N_1100,N_883,N_907);
or U1101 (N_1101,N_808,N_249);
nor U1102 (N_1102,N_389,N_767);
nand U1103 (N_1103,N_363,N_770);
nor U1104 (N_1104,N_499,N_7);
nand U1105 (N_1105,N_540,N_605);
and U1106 (N_1106,N_844,N_537);
nand U1107 (N_1107,N_304,N_643);
nor U1108 (N_1108,N_414,N_606);
nor U1109 (N_1109,N_950,N_282);
and U1110 (N_1110,N_766,N_877);
xor U1111 (N_1111,N_614,N_642);
nor U1112 (N_1112,N_508,N_447);
and U1113 (N_1113,N_793,N_755);
or U1114 (N_1114,N_833,N_789);
and U1115 (N_1115,N_974,N_724);
nand U1116 (N_1116,N_62,N_285);
nor U1117 (N_1117,N_897,N_303);
nand U1118 (N_1118,N_294,N_134);
or U1119 (N_1119,N_180,N_441);
nor U1120 (N_1120,N_239,N_776);
nor U1121 (N_1121,N_145,N_116);
or U1122 (N_1122,N_591,N_122);
and U1123 (N_1123,N_775,N_375);
and U1124 (N_1124,N_647,N_434);
or U1125 (N_1125,N_173,N_211);
or U1126 (N_1126,N_556,N_121);
nand U1127 (N_1127,N_95,N_73);
nor U1128 (N_1128,N_54,N_675);
or U1129 (N_1129,N_915,N_354);
nand U1130 (N_1130,N_119,N_550);
nand U1131 (N_1131,N_539,N_791);
nor U1132 (N_1132,N_829,N_899);
nor U1133 (N_1133,N_118,N_534);
or U1134 (N_1134,N_592,N_188);
or U1135 (N_1135,N_622,N_131);
or U1136 (N_1136,N_458,N_579);
or U1137 (N_1137,N_33,N_170);
and U1138 (N_1138,N_847,N_954);
nand U1139 (N_1139,N_113,N_66);
and U1140 (N_1140,N_852,N_75);
and U1141 (N_1141,N_289,N_857);
nor U1142 (N_1142,N_823,N_696);
or U1143 (N_1143,N_816,N_70);
or U1144 (N_1144,N_727,N_936);
nor U1145 (N_1145,N_40,N_346);
xnor U1146 (N_1146,N_631,N_671);
and U1147 (N_1147,N_371,N_799);
nor U1148 (N_1148,N_645,N_445);
xor U1149 (N_1149,N_487,N_948);
nand U1150 (N_1150,N_600,N_543);
and U1151 (N_1151,N_526,N_691);
or U1152 (N_1152,N_272,N_491);
nor U1153 (N_1153,N_0,N_739);
and U1154 (N_1154,N_762,N_433);
nor U1155 (N_1155,N_677,N_428);
or U1156 (N_1156,N_895,N_280);
and U1157 (N_1157,N_566,N_726);
nand U1158 (N_1158,N_525,N_168);
and U1159 (N_1159,N_544,N_821);
or U1160 (N_1160,N_856,N_882);
and U1161 (N_1161,N_874,N_700);
nor U1162 (N_1162,N_184,N_571);
nand U1163 (N_1163,N_372,N_705);
and U1164 (N_1164,N_89,N_154);
and U1165 (N_1165,N_782,N_514);
and U1166 (N_1166,N_381,N_593);
and U1167 (N_1167,N_254,N_416);
and U1168 (N_1168,N_69,N_684);
nand U1169 (N_1169,N_869,N_305);
nor U1170 (N_1170,N_962,N_198);
nand U1171 (N_1171,N_436,N_930);
nor U1172 (N_1172,N_717,N_455);
nand U1173 (N_1173,N_488,N_938);
nor U1174 (N_1174,N_561,N_186);
nor U1175 (N_1175,N_588,N_136);
or U1176 (N_1176,N_925,N_969);
or U1177 (N_1177,N_418,N_941);
and U1178 (N_1178,N_384,N_161);
nand U1179 (N_1179,N_603,N_551);
or U1180 (N_1180,N_521,N_457);
or U1181 (N_1181,N_669,N_679);
and U1182 (N_1182,N_610,N_815);
nand U1183 (N_1183,N_507,N_169);
nand U1184 (N_1184,N_385,N_881);
or U1185 (N_1185,N_190,N_480);
nand U1186 (N_1186,N_470,N_989);
nand U1187 (N_1187,N_364,N_50);
nand U1188 (N_1188,N_467,N_387);
nor U1189 (N_1189,N_228,N_928);
and U1190 (N_1190,N_927,N_678);
and U1191 (N_1191,N_486,N_745);
or U1192 (N_1192,N_461,N_44);
or U1193 (N_1193,N_244,N_710);
nand U1194 (N_1194,N_689,N_916);
nand U1195 (N_1195,N_953,N_673);
or U1196 (N_1196,N_553,N_251);
or U1197 (N_1197,N_426,N_383);
and U1198 (N_1198,N_967,N_720);
or U1199 (N_1199,N_565,N_52);
nand U1200 (N_1200,N_574,N_157);
nor U1201 (N_1201,N_22,N_348);
nor U1202 (N_1202,N_965,N_351);
nand U1203 (N_1203,N_329,N_8);
nand U1204 (N_1204,N_590,N_413);
nand U1205 (N_1205,N_105,N_913);
nand U1206 (N_1206,N_20,N_960);
nor U1207 (N_1207,N_112,N_577);
and U1208 (N_1208,N_731,N_476);
nor U1209 (N_1209,N_598,N_174);
or U1210 (N_1210,N_714,N_772);
or U1211 (N_1211,N_25,N_183);
and U1212 (N_1212,N_296,N_670);
xnor U1213 (N_1213,N_214,N_39);
nor U1214 (N_1214,N_796,N_71);
and U1215 (N_1215,N_323,N_935);
nor U1216 (N_1216,N_838,N_390);
or U1217 (N_1217,N_181,N_166);
nor U1218 (N_1218,N_191,N_92);
nand U1219 (N_1219,N_331,N_824);
and U1220 (N_1220,N_641,N_430);
and U1221 (N_1221,N_995,N_238);
and U1222 (N_1222,N_604,N_320);
or U1223 (N_1223,N_216,N_905);
nor U1224 (N_1224,N_35,N_328);
nor U1225 (N_1225,N_26,N_681);
nand U1226 (N_1226,N_330,N_448);
nor U1227 (N_1227,N_687,N_327);
and U1228 (N_1228,N_981,N_243);
nor U1229 (N_1229,N_527,N_290);
nand U1230 (N_1230,N_495,N_196);
and U1231 (N_1231,N_279,N_977);
nor U1232 (N_1232,N_43,N_595);
and U1233 (N_1233,N_471,N_890);
and U1234 (N_1234,N_353,N_3);
or U1235 (N_1235,N_316,N_730);
nand U1236 (N_1236,N_644,N_452);
or U1237 (N_1237,N_473,N_803);
or U1238 (N_1238,N_910,N_15);
or U1239 (N_1239,N_819,N_352);
or U1240 (N_1240,N_172,N_975);
and U1241 (N_1241,N_639,N_343);
nor U1242 (N_1242,N_41,N_704);
nor U1243 (N_1243,N_636,N_676);
and U1244 (N_1244,N_175,N_281);
or U1245 (N_1245,N_862,N_100);
nand U1246 (N_1246,N_944,N_712);
nand U1247 (N_1247,N_224,N_871);
nand U1248 (N_1248,N_394,N_923);
nand U1249 (N_1249,N_59,N_379);
and U1250 (N_1250,N_698,N_277);
nand U1251 (N_1251,N_504,N_570);
and U1252 (N_1252,N_203,N_300);
xnor U1253 (N_1253,N_401,N_502);
nand U1254 (N_1254,N_949,N_863);
and U1255 (N_1255,N_185,N_753);
or U1256 (N_1256,N_716,N_63);
nor U1257 (N_1257,N_722,N_126);
or U1258 (N_1258,N_446,N_123);
nand U1259 (N_1259,N_306,N_686);
or U1260 (N_1260,N_611,N_36);
and U1261 (N_1261,N_398,N_42);
and U1262 (N_1262,N_215,N_820);
nand U1263 (N_1263,N_314,N_76);
nand U1264 (N_1264,N_886,N_764);
nand U1265 (N_1265,N_649,N_453);
nor U1266 (N_1266,N_46,N_65);
or U1267 (N_1267,N_355,N_635);
or U1268 (N_1268,N_48,N_267);
and U1269 (N_1269,N_94,N_347);
xnor U1270 (N_1270,N_509,N_748);
and U1271 (N_1271,N_475,N_806);
and U1272 (N_1272,N_655,N_359);
or U1273 (N_1273,N_342,N_261);
nor U1274 (N_1274,N_130,N_612);
or U1275 (N_1275,N_576,N_195);
and U1276 (N_1276,N_575,N_660);
and U1277 (N_1277,N_265,N_988);
and U1278 (N_1278,N_983,N_519);
and U1279 (N_1279,N_752,N_528);
nand U1280 (N_1280,N_117,N_23);
or U1281 (N_1281,N_903,N_219);
nand U1282 (N_1282,N_846,N_901);
nand U1283 (N_1283,N_97,N_259);
nor U1284 (N_1284,N_959,N_13);
or U1285 (N_1285,N_986,N_86);
or U1286 (N_1286,N_178,N_807);
nand U1287 (N_1287,N_365,N_421);
nand U1288 (N_1288,N_951,N_74);
or U1289 (N_1289,N_708,N_465);
and U1290 (N_1290,N_648,N_513);
or U1291 (N_1291,N_423,N_392);
or U1292 (N_1292,N_49,N_93);
or U1293 (N_1293,N_993,N_478);
and U1294 (N_1294,N_242,N_860);
or U1295 (N_1295,N_744,N_102);
or U1296 (N_1296,N_786,N_250);
and U1297 (N_1297,N_625,N_868);
nand U1298 (N_1298,N_867,N_707);
nor U1299 (N_1299,N_324,N_827);
and U1300 (N_1300,N_101,N_695);
or U1301 (N_1301,N_497,N_946);
nand U1302 (N_1302,N_419,N_839);
or U1303 (N_1303,N_462,N_692);
nand U1304 (N_1304,N_864,N_493);
nand U1305 (N_1305,N_270,N_524);
nand U1306 (N_1306,N_483,N_735);
and U1307 (N_1307,N_801,N_569);
and U1308 (N_1308,N_546,N_699);
and U1309 (N_1309,N_547,N_482);
nor U1310 (N_1310,N_376,N_240);
nor U1311 (N_1311,N_481,N_599);
or U1312 (N_1312,N_718,N_449);
and U1313 (N_1313,N_350,N_510);
and U1314 (N_1314,N_149,N_310);
nor U1315 (N_1315,N_623,N_840);
and U1316 (N_1316,N_817,N_889);
and U1317 (N_1317,N_223,N_618);
nand U1318 (N_1318,N_260,N_360);
and U1319 (N_1319,N_964,N_774);
or U1320 (N_1320,N_459,N_179);
nand U1321 (N_1321,N_942,N_128);
or U1322 (N_1322,N_765,N_734);
or U1323 (N_1323,N_741,N_53);
and U1324 (N_1324,N_345,N_737);
or U1325 (N_1325,N_784,N_506);
nor U1326 (N_1326,N_763,N_206);
xor U1327 (N_1327,N_432,N_273);
nor U1328 (N_1328,N_1,N_205);
nor U1329 (N_1329,N_790,N_586);
and U1330 (N_1330,N_368,N_129);
and U1331 (N_1331,N_12,N_29);
or U1332 (N_1332,N_773,N_832);
nand U1333 (N_1333,N_143,N_230);
and U1334 (N_1334,N_711,N_248);
nand U1335 (N_1335,N_918,N_932);
or U1336 (N_1336,N_412,N_568);
and U1337 (N_1337,N_106,N_947);
nor U1338 (N_1338,N_301,N_358);
or U1339 (N_1339,N_297,N_336);
nor U1340 (N_1340,N_252,N_621);
or U1341 (N_1341,N_266,N_841);
nand U1342 (N_1342,N_246,N_680);
nand U1343 (N_1343,N_998,N_18);
or U1344 (N_1344,N_854,N_548);
and U1345 (N_1345,N_313,N_88);
nand U1346 (N_1346,N_82,N_758);
and U1347 (N_1347,N_335,N_237);
nor U1348 (N_1348,N_943,N_276);
nand U1349 (N_1349,N_912,N_357);
nand U1350 (N_1350,N_268,N_887);
nor U1351 (N_1351,N_650,N_845);
nor U1352 (N_1352,N_165,N_60);
or U1353 (N_1353,N_319,N_374);
nand U1354 (N_1354,N_139,N_800);
nand U1355 (N_1355,N_836,N_898);
or U1356 (N_1356,N_958,N_798);
or U1357 (N_1357,N_47,N_640);
or U1358 (N_1358,N_538,N_945);
and U1359 (N_1359,N_872,N_996);
nor U1360 (N_1360,N_56,N_956);
nand U1361 (N_1361,N_879,N_234);
nor U1362 (N_1362,N_842,N_19);
nand U1363 (N_1363,N_464,N_728);
and U1364 (N_1364,N_232,N_738);
nand U1365 (N_1365,N_386,N_287);
nor U1366 (N_1366,N_435,N_715);
nand U1367 (N_1367,N_794,N_292);
nor U1368 (N_1368,N_515,N_578);
and U1369 (N_1369,N_541,N_110);
or U1370 (N_1370,N_978,N_442);
nand U1371 (N_1371,N_312,N_158);
and U1372 (N_1372,N_162,N_613);
xor U1373 (N_1373,N_38,N_597);
or U1374 (N_1374,N_396,N_425);
nand U1375 (N_1375,N_373,N_542);
and U1376 (N_1376,N_77,N_51);
nand U1377 (N_1377,N_325,N_666);
nor U1378 (N_1378,N_28,N_627);
or U1379 (N_1379,N_218,N_601);
and U1380 (N_1380,N_284,N_468);
and U1381 (N_1381,N_217,N_994);
nand U1382 (N_1382,N_67,N_567);
and U1383 (N_1383,N_992,N_120);
or U1384 (N_1384,N_701,N_835);
nand U1385 (N_1385,N_298,N_213);
or U1386 (N_1386,N_378,N_955);
nor U1387 (N_1387,N_518,N_229);
nand U1388 (N_1388,N_341,N_531);
nor U1389 (N_1389,N_629,N_674);
and U1390 (N_1390,N_403,N_333);
nand U1391 (N_1391,N_533,N_247);
nand U1392 (N_1392,N_587,N_477);
nor U1393 (N_1393,N_783,N_991);
or U1394 (N_1394,N_797,N_309);
xor U1395 (N_1395,N_902,N_498);
and U1396 (N_1396,N_440,N_55);
and U1397 (N_1397,N_919,N_257);
nand U1398 (N_1398,N_225,N_496);
xnor U1399 (N_1399,N_474,N_904);
nand U1400 (N_1400,N_900,N_828);
or U1401 (N_1401,N_469,N_878);
and U1402 (N_1402,N_235,N_127);
nor U1403 (N_1403,N_523,N_138);
nor U1404 (N_1404,N_870,N_626);
nand U1405 (N_1405,N_332,N_107);
nand U1406 (N_1406,N_236,N_199);
or U1407 (N_1407,N_966,N_207);
nor U1408 (N_1408,N_402,N_825);
nand U1409 (N_1409,N_194,N_443);
nand U1410 (N_1410,N_997,N_189);
nand U1411 (N_1411,N_103,N_536);
nor U1412 (N_1412,N_150,N_322);
nand U1413 (N_1413,N_388,N_494);
nand U1414 (N_1414,N_596,N_769);
and U1415 (N_1415,N_554,N_159);
nand U1416 (N_1416,N_608,N_14);
nor U1417 (N_1417,N_562,N_617);
and U1418 (N_1418,N_557,N_2);
nand U1419 (N_1419,N_929,N_968);
and U1420 (N_1420,N_853,N_202);
and U1421 (N_1421,N_361,N_661);
and U1422 (N_1422,N_182,N_160);
xnor U1423 (N_1423,N_231,N_233);
and U1424 (N_1424,N_522,N_934);
and U1425 (N_1425,N_572,N_814);
nor U1426 (N_1426,N_713,N_585);
or U1427 (N_1427,N_906,N_30);
or U1428 (N_1428,N_750,N_197);
nor U1429 (N_1429,N_646,N_11);
and U1430 (N_1430,N_104,N_788);
nor U1431 (N_1431,N_10,N_979);
and U1432 (N_1432,N_395,N_255);
and U1433 (N_1433,N_271,N_580);
nand U1434 (N_1434,N_822,N_501);
and U1435 (N_1435,N_84,N_638);
and U1436 (N_1436,N_985,N_980);
nand U1437 (N_1437,N_609,N_837);
and U1438 (N_1438,N_420,N_861);
nand U1439 (N_1439,N_339,N_917);
nand U1440 (N_1440,N_961,N_963);
nand U1441 (N_1441,N_875,N_658);
and U1442 (N_1442,N_517,N_410);
nor U1443 (N_1443,N_422,N_873);
nand U1444 (N_1444,N_558,N_85);
nor U1445 (N_1445,N_760,N_155);
nand U1446 (N_1446,N_241,N_406);
nand U1447 (N_1447,N_163,N_334);
and U1448 (N_1448,N_659,N_204);
and U1449 (N_1449,N_263,N_302);
and U1450 (N_1450,N_187,N_771);
and U1451 (N_1451,N_81,N_466);
and U1452 (N_1452,N_264,N_663);
or U1453 (N_1453,N_221,N_91);
or U1454 (N_1454,N_931,N_124);
or U1455 (N_1455,N_177,N_362);
or U1456 (N_1456,N_171,N_933);
nand U1457 (N_1457,N_274,N_589);
and U1458 (N_1458,N_552,N_921);
and U1459 (N_1459,N_210,N_132);
nand U1460 (N_1460,N_736,N_894);
and U1461 (N_1461,N_489,N_256);
nand U1462 (N_1462,N_703,N_802);
nand U1463 (N_1463,N_147,N_16);
nand U1464 (N_1464,N_115,N_781);
nand U1465 (N_1465,N_429,N_563);
nor U1466 (N_1466,N_500,N_858);
or U1467 (N_1467,N_757,N_982);
xor U1468 (N_1468,N_792,N_653);
nand U1469 (N_1469,N_831,N_209);
nand U1470 (N_1470,N_880,N_283);
and U1471 (N_1471,N_634,N_768);
and U1472 (N_1472,N_454,N_45);
and U1473 (N_1473,N_293,N_80);
and U1474 (N_1474,N_682,N_90);
and U1475 (N_1475,N_812,N_759);
nor U1476 (N_1476,N_530,N_114);
and U1477 (N_1477,N_813,N_984);
or U1478 (N_1478,N_665,N_193);
or U1479 (N_1479,N_970,N_688);
nand U1480 (N_1480,N_615,N_654);
nor U1481 (N_1481,N_779,N_754);
and U1482 (N_1482,N_407,N_957);
and U1483 (N_1483,N_411,N_382);
nand U1484 (N_1484,N_805,N_311);
and U1485 (N_1485,N_144,N_5);
nand U1486 (N_1486,N_78,N_532);
nor U1487 (N_1487,N_299,N_31);
or U1488 (N_1488,N_479,N_370);
nor U1489 (N_1489,N_520,N_291);
xor U1490 (N_1490,N_427,N_253);
and U1491 (N_1491,N_787,N_450);
or U1492 (N_1492,N_751,N_98);
xor U1493 (N_1493,N_795,N_843);
or U1494 (N_1494,N_693,N_437);
or U1495 (N_1495,N_79,N_637);
or U1496 (N_1496,N_672,N_721);
and U1497 (N_1497,N_64,N_141);
or U1498 (N_1498,N_393,N_516);
nor U1499 (N_1499,N_505,N_307);
nor U1500 (N_1500,N_150,N_783);
and U1501 (N_1501,N_731,N_516);
nand U1502 (N_1502,N_523,N_925);
or U1503 (N_1503,N_419,N_378);
nor U1504 (N_1504,N_369,N_212);
nand U1505 (N_1505,N_488,N_259);
nand U1506 (N_1506,N_28,N_754);
or U1507 (N_1507,N_456,N_965);
and U1508 (N_1508,N_883,N_869);
nor U1509 (N_1509,N_853,N_353);
nand U1510 (N_1510,N_24,N_915);
xor U1511 (N_1511,N_890,N_753);
nor U1512 (N_1512,N_743,N_350);
or U1513 (N_1513,N_963,N_817);
or U1514 (N_1514,N_147,N_817);
nand U1515 (N_1515,N_925,N_556);
or U1516 (N_1516,N_126,N_850);
nand U1517 (N_1517,N_335,N_434);
nand U1518 (N_1518,N_590,N_565);
nor U1519 (N_1519,N_920,N_798);
nand U1520 (N_1520,N_421,N_694);
and U1521 (N_1521,N_784,N_881);
nand U1522 (N_1522,N_86,N_373);
nand U1523 (N_1523,N_777,N_25);
or U1524 (N_1524,N_407,N_422);
nor U1525 (N_1525,N_599,N_656);
nand U1526 (N_1526,N_398,N_296);
or U1527 (N_1527,N_676,N_161);
nand U1528 (N_1528,N_981,N_990);
and U1529 (N_1529,N_885,N_939);
nor U1530 (N_1530,N_616,N_50);
and U1531 (N_1531,N_544,N_613);
or U1532 (N_1532,N_173,N_590);
nand U1533 (N_1533,N_634,N_170);
and U1534 (N_1534,N_440,N_840);
nand U1535 (N_1535,N_115,N_79);
nand U1536 (N_1536,N_172,N_978);
nor U1537 (N_1537,N_886,N_712);
or U1538 (N_1538,N_132,N_292);
or U1539 (N_1539,N_240,N_724);
nand U1540 (N_1540,N_88,N_548);
and U1541 (N_1541,N_941,N_64);
and U1542 (N_1542,N_535,N_253);
and U1543 (N_1543,N_834,N_22);
nand U1544 (N_1544,N_732,N_302);
nor U1545 (N_1545,N_515,N_557);
or U1546 (N_1546,N_184,N_349);
nand U1547 (N_1547,N_924,N_230);
nor U1548 (N_1548,N_653,N_531);
or U1549 (N_1549,N_214,N_425);
and U1550 (N_1550,N_377,N_168);
or U1551 (N_1551,N_189,N_869);
or U1552 (N_1552,N_577,N_443);
or U1553 (N_1553,N_725,N_694);
nand U1554 (N_1554,N_149,N_94);
and U1555 (N_1555,N_256,N_560);
nand U1556 (N_1556,N_697,N_124);
and U1557 (N_1557,N_659,N_194);
nor U1558 (N_1558,N_690,N_292);
nor U1559 (N_1559,N_907,N_271);
or U1560 (N_1560,N_147,N_596);
nand U1561 (N_1561,N_702,N_361);
nor U1562 (N_1562,N_970,N_246);
nand U1563 (N_1563,N_993,N_965);
or U1564 (N_1564,N_476,N_179);
nor U1565 (N_1565,N_976,N_778);
and U1566 (N_1566,N_634,N_227);
and U1567 (N_1567,N_391,N_556);
nor U1568 (N_1568,N_600,N_12);
and U1569 (N_1569,N_495,N_92);
or U1570 (N_1570,N_726,N_871);
nor U1571 (N_1571,N_875,N_70);
nand U1572 (N_1572,N_377,N_153);
and U1573 (N_1573,N_398,N_223);
and U1574 (N_1574,N_601,N_449);
nor U1575 (N_1575,N_619,N_620);
nor U1576 (N_1576,N_965,N_990);
nand U1577 (N_1577,N_290,N_316);
and U1578 (N_1578,N_642,N_979);
nor U1579 (N_1579,N_306,N_575);
nand U1580 (N_1580,N_626,N_101);
xor U1581 (N_1581,N_974,N_859);
nand U1582 (N_1582,N_769,N_77);
and U1583 (N_1583,N_341,N_474);
nand U1584 (N_1584,N_795,N_928);
or U1585 (N_1585,N_769,N_905);
nor U1586 (N_1586,N_631,N_646);
and U1587 (N_1587,N_221,N_581);
nand U1588 (N_1588,N_734,N_429);
and U1589 (N_1589,N_174,N_300);
nand U1590 (N_1590,N_625,N_532);
nand U1591 (N_1591,N_758,N_699);
and U1592 (N_1592,N_378,N_489);
and U1593 (N_1593,N_57,N_791);
nor U1594 (N_1594,N_305,N_737);
and U1595 (N_1595,N_589,N_29);
nor U1596 (N_1596,N_679,N_139);
nor U1597 (N_1597,N_131,N_947);
and U1598 (N_1598,N_350,N_233);
or U1599 (N_1599,N_328,N_213);
nor U1600 (N_1600,N_176,N_754);
nand U1601 (N_1601,N_187,N_555);
nand U1602 (N_1602,N_815,N_885);
and U1603 (N_1603,N_915,N_586);
nand U1604 (N_1604,N_860,N_171);
nand U1605 (N_1605,N_245,N_169);
or U1606 (N_1606,N_420,N_727);
nand U1607 (N_1607,N_259,N_770);
or U1608 (N_1608,N_497,N_321);
and U1609 (N_1609,N_463,N_154);
and U1610 (N_1610,N_838,N_441);
and U1611 (N_1611,N_702,N_103);
nand U1612 (N_1612,N_101,N_777);
nand U1613 (N_1613,N_391,N_637);
nand U1614 (N_1614,N_803,N_708);
nor U1615 (N_1615,N_362,N_787);
and U1616 (N_1616,N_880,N_971);
nor U1617 (N_1617,N_610,N_57);
nor U1618 (N_1618,N_845,N_392);
nor U1619 (N_1619,N_857,N_839);
and U1620 (N_1620,N_165,N_217);
and U1621 (N_1621,N_381,N_48);
or U1622 (N_1622,N_578,N_360);
nand U1623 (N_1623,N_871,N_99);
and U1624 (N_1624,N_547,N_127);
or U1625 (N_1625,N_877,N_715);
and U1626 (N_1626,N_988,N_982);
nor U1627 (N_1627,N_60,N_552);
nand U1628 (N_1628,N_190,N_643);
or U1629 (N_1629,N_99,N_147);
and U1630 (N_1630,N_524,N_611);
or U1631 (N_1631,N_66,N_970);
nor U1632 (N_1632,N_420,N_338);
nor U1633 (N_1633,N_618,N_9);
and U1634 (N_1634,N_11,N_343);
nand U1635 (N_1635,N_404,N_799);
xor U1636 (N_1636,N_979,N_975);
nor U1637 (N_1637,N_399,N_182);
or U1638 (N_1638,N_125,N_806);
or U1639 (N_1639,N_880,N_784);
and U1640 (N_1640,N_15,N_996);
nand U1641 (N_1641,N_920,N_873);
and U1642 (N_1642,N_731,N_863);
or U1643 (N_1643,N_692,N_624);
nand U1644 (N_1644,N_115,N_779);
nor U1645 (N_1645,N_83,N_59);
nand U1646 (N_1646,N_232,N_331);
nand U1647 (N_1647,N_696,N_542);
or U1648 (N_1648,N_588,N_905);
or U1649 (N_1649,N_78,N_920);
or U1650 (N_1650,N_157,N_915);
and U1651 (N_1651,N_208,N_641);
nor U1652 (N_1652,N_597,N_638);
nor U1653 (N_1653,N_704,N_758);
nand U1654 (N_1654,N_880,N_840);
and U1655 (N_1655,N_924,N_286);
and U1656 (N_1656,N_464,N_62);
nand U1657 (N_1657,N_359,N_798);
and U1658 (N_1658,N_820,N_699);
or U1659 (N_1659,N_285,N_325);
nor U1660 (N_1660,N_487,N_398);
or U1661 (N_1661,N_387,N_162);
or U1662 (N_1662,N_186,N_181);
nor U1663 (N_1663,N_290,N_128);
or U1664 (N_1664,N_471,N_782);
or U1665 (N_1665,N_844,N_58);
or U1666 (N_1666,N_213,N_343);
and U1667 (N_1667,N_766,N_381);
or U1668 (N_1668,N_383,N_435);
nor U1669 (N_1669,N_421,N_478);
or U1670 (N_1670,N_248,N_542);
and U1671 (N_1671,N_449,N_793);
nand U1672 (N_1672,N_752,N_570);
nor U1673 (N_1673,N_985,N_215);
nand U1674 (N_1674,N_429,N_185);
nor U1675 (N_1675,N_851,N_650);
or U1676 (N_1676,N_962,N_713);
or U1677 (N_1677,N_831,N_245);
and U1678 (N_1678,N_542,N_914);
nand U1679 (N_1679,N_789,N_339);
nor U1680 (N_1680,N_210,N_717);
nand U1681 (N_1681,N_791,N_179);
nor U1682 (N_1682,N_164,N_528);
or U1683 (N_1683,N_809,N_429);
nand U1684 (N_1684,N_465,N_929);
xnor U1685 (N_1685,N_200,N_563);
and U1686 (N_1686,N_785,N_413);
nor U1687 (N_1687,N_375,N_312);
and U1688 (N_1688,N_768,N_769);
and U1689 (N_1689,N_210,N_150);
nand U1690 (N_1690,N_516,N_411);
and U1691 (N_1691,N_479,N_780);
nand U1692 (N_1692,N_110,N_413);
nand U1693 (N_1693,N_976,N_723);
or U1694 (N_1694,N_908,N_668);
nor U1695 (N_1695,N_297,N_824);
and U1696 (N_1696,N_647,N_122);
or U1697 (N_1697,N_607,N_170);
and U1698 (N_1698,N_464,N_619);
nand U1699 (N_1699,N_975,N_797);
or U1700 (N_1700,N_437,N_949);
and U1701 (N_1701,N_557,N_417);
nor U1702 (N_1702,N_871,N_282);
and U1703 (N_1703,N_836,N_111);
nor U1704 (N_1704,N_514,N_119);
and U1705 (N_1705,N_935,N_13);
and U1706 (N_1706,N_102,N_442);
nand U1707 (N_1707,N_552,N_444);
nand U1708 (N_1708,N_401,N_713);
nand U1709 (N_1709,N_417,N_902);
nand U1710 (N_1710,N_389,N_53);
or U1711 (N_1711,N_376,N_968);
and U1712 (N_1712,N_813,N_369);
nand U1713 (N_1713,N_112,N_7);
nand U1714 (N_1714,N_121,N_153);
nand U1715 (N_1715,N_127,N_70);
nand U1716 (N_1716,N_871,N_672);
or U1717 (N_1717,N_127,N_225);
and U1718 (N_1718,N_296,N_534);
nand U1719 (N_1719,N_79,N_476);
and U1720 (N_1720,N_244,N_298);
and U1721 (N_1721,N_737,N_205);
nor U1722 (N_1722,N_687,N_654);
xnor U1723 (N_1723,N_169,N_982);
nor U1724 (N_1724,N_58,N_683);
and U1725 (N_1725,N_39,N_615);
nand U1726 (N_1726,N_747,N_190);
nor U1727 (N_1727,N_690,N_808);
or U1728 (N_1728,N_872,N_52);
and U1729 (N_1729,N_71,N_756);
and U1730 (N_1730,N_792,N_659);
and U1731 (N_1731,N_818,N_483);
nand U1732 (N_1732,N_615,N_131);
nor U1733 (N_1733,N_568,N_481);
and U1734 (N_1734,N_790,N_100);
nor U1735 (N_1735,N_646,N_813);
nor U1736 (N_1736,N_131,N_107);
nor U1737 (N_1737,N_242,N_902);
or U1738 (N_1738,N_459,N_501);
or U1739 (N_1739,N_96,N_818);
nor U1740 (N_1740,N_878,N_380);
and U1741 (N_1741,N_162,N_155);
and U1742 (N_1742,N_946,N_438);
or U1743 (N_1743,N_48,N_919);
nor U1744 (N_1744,N_919,N_37);
nand U1745 (N_1745,N_645,N_351);
and U1746 (N_1746,N_513,N_973);
nand U1747 (N_1747,N_268,N_742);
nor U1748 (N_1748,N_590,N_753);
nand U1749 (N_1749,N_415,N_856);
nor U1750 (N_1750,N_329,N_468);
nand U1751 (N_1751,N_883,N_725);
and U1752 (N_1752,N_527,N_626);
or U1753 (N_1753,N_889,N_565);
or U1754 (N_1754,N_267,N_223);
or U1755 (N_1755,N_821,N_402);
and U1756 (N_1756,N_425,N_222);
nand U1757 (N_1757,N_556,N_297);
or U1758 (N_1758,N_54,N_363);
nor U1759 (N_1759,N_941,N_416);
nand U1760 (N_1760,N_533,N_59);
nand U1761 (N_1761,N_753,N_742);
and U1762 (N_1762,N_993,N_215);
and U1763 (N_1763,N_25,N_227);
nor U1764 (N_1764,N_620,N_843);
nand U1765 (N_1765,N_505,N_84);
nand U1766 (N_1766,N_331,N_161);
nand U1767 (N_1767,N_731,N_478);
and U1768 (N_1768,N_249,N_643);
nor U1769 (N_1769,N_318,N_465);
and U1770 (N_1770,N_40,N_636);
nand U1771 (N_1771,N_369,N_844);
or U1772 (N_1772,N_338,N_136);
and U1773 (N_1773,N_272,N_267);
nand U1774 (N_1774,N_683,N_206);
nand U1775 (N_1775,N_816,N_955);
nand U1776 (N_1776,N_42,N_732);
nor U1777 (N_1777,N_358,N_83);
nor U1778 (N_1778,N_740,N_642);
and U1779 (N_1779,N_331,N_997);
or U1780 (N_1780,N_441,N_271);
or U1781 (N_1781,N_231,N_686);
and U1782 (N_1782,N_549,N_947);
nor U1783 (N_1783,N_731,N_723);
or U1784 (N_1784,N_567,N_969);
or U1785 (N_1785,N_373,N_196);
nor U1786 (N_1786,N_943,N_227);
and U1787 (N_1787,N_370,N_564);
or U1788 (N_1788,N_30,N_949);
and U1789 (N_1789,N_470,N_524);
nand U1790 (N_1790,N_288,N_60);
nand U1791 (N_1791,N_824,N_94);
nor U1792 (N_1792,N_651,N_847);
and U1793 (N_1793,N_855,N_20);
nand U1794 (N_1794,N_970,N_886);
and U1795 (N_1795,N_449,N_781);
nand U1796 (N_1796,N_30,N_882);
and U1797 (N_1797,N_873,N_939);
and U1798 (N_1798,N_405,N_198);
xnor U1799 (N_1799,N_769,N_100);
or U1800 (N_1800,N_634,N_479);
or U1801 (N_1801,N_373,N_956);
nor U1802 (N_1802,N_792,N_24);
nor U1803 (N_1803,N_125,N_963);
and U1804 (N_1804,N_496,N_42);
nor U1805 (N_1805,N_443,N_172);
or U1806 (N_1806,N_341,N_317);
nor U1807 (N_1807,N_644,N_125);
or U1808 (N_1808,N_383,N_877);
nor U1809 (N_1809,N_218,N_656);
nand U1810 (N_1810,N_367,N_297);
nand U1811 (N_1811,N_86,N_730);
nor U1812 (N_1812,N_125,N_892);
nor U1813 (N_1813,N_372,N_642);
nand U1814 (N_1814,N_878,N_941);
and U1815 (N_1815,N_358,N_408);
or U1816 (N_1816,N_519,N_490);
nor U1817 (N_1817,N_26,N_917);
and U1818 (N_1818,N_34,N_828);
nand U1819 (N_1819,N_866,N_242);
and U1820 (N_1820,N_938,N_62);
nand U1821 (N_1821,N_447,N_612);
nand U1822 (N_1822,N_640,N_883);
nor U1823 (N_1823,N_730,N_957);
or U1824 (N_1824,N_849,N_411);
and U1825 (N_1825,N_243,N_639);
nor U1826 (N_1826,N_924,N_85);
or U1827 (N_1827,N_763,N_131);
or U1828 (N_1828,N_892,N_983);
and U1829 (N_1829,N_868,N_643);
nand U1830 (N_1830,N_600,N_568);
and U1831 (N_1831,N_205,N_465);
xor U1832 (N_1832,N_399,N_491);
nand U1833 (N_1833,N_564,N_392);
nand U1834 (N_1834,N_244,N_327);
nand U1835 (N_1835,N_528,N_445);
nand U1836 (N_1836,N_268,N_618);
and U1837 (N_1837,N_547,N_916);
and U1838 (N_1838,N_19,N_828);
nand U1839 (N_1839,N_314,N_694);
nor U1840 (N_1840,N_103,N_914);
and U1841 (N_1841,N_803,N_415);
nand U1842 (N_1842,N_541,N_856);
xor U1843 (N_1843,N_131,N_355);
nand U1844 (N_1844,N_887,N_48);
or U1845 (N_1845,N_287,N_747);
and U1846 (N_1846,N_850,N_897);
nor U1847 (N_1847,N_254,N_788);
or U1848 (N_1848,N_654,N_439);
nand U1849 (N_1849,N_524,N_377);
nand U1850 (N_1850,N_12,N_468);
and U1851 (N_1851,N_980,N_141);
or U1852 (N_1852,N_854,N_107);
and U1853 (N_1853,N_250,N_904);
and U1854 (N_1854,N_46,N_438);
nor U1855 (N_1855,N_841,N_193);
nor U1856 (N_1856,N_442,N_494);
nand U1857 (N_1857,N_704,N_972);
and U1858 (N_1858,N_645,N_798);
or U1859 (N_1859,N_988,N_93);
nand U1860 (N_1860,N_140,N_404);
nor U1861 (N_1861,N_2,N_485);
and U1862 (N_1862,N_780,N_403);
or U1863 (N_1863,N_423,N_164);
or U1864 (N_1864,N_246,N_346);
nand U1865 (N_1865,N_206,N_370);
and U1866 (N_1866,N_112,N_490);
nor U1867 (N_1867,N_716,N_667);
and U1868 (N_1868,N_546,N_937);
nor U1869 (N_1869,N_54,N_274);
nor U1870 (N_1870,N_507,N_379);
nand U1871 (N_1871,N_807,N_270);
and U1872 (N_1872,N_869,N_687);
nand U1873 (N_1873,N_275,N_0);
nor U1874 (N_1874,N_675,N_589);
nor U1875 (N_1875,N_930,N_634);
xor U1876 (N_1876,N_997,N_143);
or U1877 (N_1877,N_914,N_601);
and U1878 (N_1878,N_918,N_791);
or U1879 (N_1879,N_412,N_413);
nand U1880 (N_1880,N_444,N_477);
nor U1881 (N_1881,N_738,N_87);
or U1882 (N_1882,N_515,N_97);
nand U1883 (N_1883,N_877,N_557);
xnor U1884 (N_1884,N_769,N_990);
xor U1885 (N_1885,N_358,N_233);
and U1886 (N_1886,N_223,N_530);
nand U1887 (N_1887,N_646,N_29);
nand U1888 (N_1888,N_606,N_921);
nor U1889 (N_1889,N_544,N_260);
or U1890 (N_1890,N_285,N_779);
or U1891 (N_1891,N_100,N_323);
nor U1892 (N_1892,N_966,N_408);
nor U1893 (N_1893,N_613,N_699);
nand U1894 (N_1894,N_975,N_669);
or U1895 (N_1895,N_694,N_140);
or U1896 (N_1896,N_128,N_259);
nand U1897 (N_1897,N_679,N_502);
or U1898 (N_1898,N_653,N_850);
nand U1899 (N_1899,N_716,N_665);
or U1900 (N_1900,N_92,N_626);
or U1901 (N_1901,N_189,N_550);
and U1902 (N_1902,N_342,N_770);
or U1903 (N_1903,N_726,N_452);
nor U1904 (N_1904,N_655,N_745);
and U1905 (N_1905,N_551,N_888);
or U1906 (N_1906,N_451,N_261);
nor U1907 (N_1907,N_341,N_977);
and U1908 (N_1908,N_632,N_347);
nor U1909 (N_1909,N_324,N_223);
or U1910 (N_1910,N_354,N_208);
nor U1911 (N_1911,N_366,N_286);
and U1912 (N_1912,N_848,N_369);
and U1913 (N_1913,N_542,N_90);
nand U1914 (N_1914,N_640,N_134);
nand U1915 (N_1915,N_689,N_326);
or U1916 (N_1916,N_116,N_747);
and U1917 (N_1917,N_772,N_230);
nor U1918 (N_1918,N_672,N_62);
or U1919 (N_1919,N_70,N_850);
or U1920 (N_1920,N_850,N_96);
or U1921 (N_1921,N_300,N_94);
nor U1922 (N_1922,N_473,N_716);
or U1923 (N_1923,N_364,N_20);
or U1924 (N_1924,N_40,N_391);
nor U1925 (N_1925,N_938,N_236);
or U1926 (N_1926,N_461,N_292);
and U1927 (N_1927,N_604,N_591);
nor U1928 (N_1928,N_704,N_691);
and U1929 (N_1929,N_896,N_936);
nor U1930 (N_1930,N_547,N_267);
nand U1931 (N_1931,N_61,N_346);
or U1932 (N_1932,N_112,N_376);
and U1933 (N_1933,N_668,N_187);
nand U1934 (N_1934,N_215,N_179);
nor U1935 (N_1935,N_292,N_330);
nor U1936 (N_1936,N_637,N_152);
or U1937 (N_1937,N_884,N_153);
nor U1938 (N_1938,N_450,N_785);
nand U1939 (N_1939,N_911,N_409);
and U1940 (N_1940,N_50,N_103);
and U1941 (N_1941,N_789,N_279);
nor U1942 (N_1942,N_757,N_279);
xnor U1943 (N_1943,N_111,N_320);
or U1944 (N_1944,N_313,N_248);
nand U1945 (N_1945,N_866,N_198);
or U1946 (N_1946,N_698,N_718);
and U1947 (N_1947,N_47,N_733);
nor U1948 (N_1948,N_705,N_736);
nor U1949 (N_1949,N_421,N_250);
or U1950 (N_1950,N_528,N_25);
nor U1951 (N_1951,N_163,N_282);
nor U1952 (N_1952,N_355,N_465);
and U1953 (N_1953,N_870,N_538);
nand U1954 (N_1954,N_887,N_945);
and U1955 (N_1955,N_116,N_573);
and U1956 (N_1956,N_280,N_492);
nor U1957 (N_1957,N_436,N_194);
nor U1958 (N_1958,N_357,N_733);
or U1959 (N_1959,N_331,N_155);
and U1960 (N_1960,N_31,N_672);
nand U1961 (N_1961,N_218,N_483);
or U1962 (N_1962,N_659,N_817);
nand U1963 (N_1963,N_645,N_931);
nor U1964 (N_1964,N_589,N_774);
nand U1965 (N_1965,N_163,N_900);
nand U1966 (N_1966,N_418,N_408);
nor U1967 (N_1967,N_845,N_132);
or U1968 (N_1968,N_220,N_486);
nand U1969 (N_1969,N_344,N_336);
or U1970 (N_1970,N_128,N_909);
nor U1971 (N_1971,N_32,N_197);
and U1972 (N_1972,N_928,N_490);
nor U1973 (N_1973,N_20,N_514);
and U1974 (N_1974,N_295,N_523);
and U1975 (N_1975,N_351,N_100);
or U1976 (N_1976,N_114,N_301);
nor U1977 (N_1977,N_191,N_590);
or U1978 (N_1978,N_968,N_961);
nor U1979 (N_1979,N_863,N_150);
nor U1980 (N_1980,N_77,N_763);
nand U1981 (N_1981,N_352,N_824);
or U1982 (N_1982,N_290,N_771);
nor U1983 (N_1983,N_978,N_832);
and U1984 (N_1984,N_738,N_116);
and U1985 (N_1985,N_747,N_264);
or U1986 (N_1986,N_826,N_873);
nor U1987 (N_1987,N_902,N_480);
or U1988 (N_1988,N_565,N_206);
and U1989 (N_1989,N_856,N_318);
nand U1990 (N_1990,N_586,N_712);
nor U1991 (N_1991,N_941,N_387);
and U1992 (N_1992,N_72,N_614);
and U1993 (N_1993,N_927,N_571);
nor U1994 (N_1994,N_607,N_850);
or U1995 (N_1995,N_919,N_638);
and U1996 (N_1996,N_644,N_594);
xor U1997 (N_1997,N_892,N_188);
nor U1998 (N_1998,N_438,N_207);
nand U1999 (N_1999,N_990,N_779);
and U2000 (N_2000,N_1051,N_1148);
or U2001 (N_2001,N_1065,N_1090);
or U2002 (N_2002,N_1158,N_1726);
nor U2003 (N_2003,N_1864,N_1178);
nand U2004 (N_2004,N_1219,N_1365);
nand U2005 (N_2005,N_1211,N_1594);
or U2006 (N_2006,N_1191,N_1984);
and U2007 (N_2007,N_1265,N_1913);
nand U2008 (N_2008,N_1624,N_1412);
nand U2009 (N_2009,N_1441,N_1427);
or U2010 (N_2010,N_1662,N_1709);
and U2011 (N_2011,N_1021,N_1223);
or U2012 (N_2012,N_1703,N_1194);
nand U2013 (N_2013,N_1399,N_1909);
and U2014 (N_2014,N_1453,N_1062);
and U2015 (N_2015,N_1487,N_1149);
nand U2016 (N_2016,N_1239,N_1401);
nand U2017 (N_2017,N_1436,N_1690);
and U2018 (N_2018,N_1004,N_1992);
or U2019 (N_2019,N_1147,N_1197);
nand U2020 (N_2020,N_1081,N_1146);
and U2021 (N_2021,N_1718,N_1664);
and U2022 (N_2022,N_1430,N_1565);
or U2023 (N_2023,N_1204,N_1267);
nor U2024 (N_2024,N_1393,N_1691);
and U2025 (N_2025,N_1126,N_1614);
or U2026 (N_2026,N_1829,N_1426);
or U2027 (N_2027,N_1716,N_1862);
nor U2028 (N_2028,N_1380,N_1776);
nand U2029 (N_2029,N_1564,N_1740);
nor U2030 (N_2030,N_1579,N_1446);
or U2031 (N_2031,N_1405,N_1171);
and U2032 (N_2032,N_1989,N_1605);
xnor U2033 (N_2033,N_1979,N_1230);
nand U2034 (N_2034,N_1654,N_1739);
and U2035 (N_2035,N_1530,N_1256);
or U2036 (N_2036,N_1082,N_1731);
nand U2037 (N_2037,N_1472,N_1429);
nand U2038 (N_2038,N_1708,N_1217);
or U2039 (N_2039,N_1272,N_1200);
and U2040 (N_2040,N_1074,N_1448);
nor U2041 (N_2041,N_1693,N_1033);
nand U2042 (N_2042,N_1028,N_1612);
or U2043 (N_2043,N_1023,N_1833);
nand U2044 (N_2044,N_1767,N_1069);
nand U2045 (N_2045,N_1712,N_1325);
xor U2046 (N_2046,N_1554,N_1407);
or U2047 (N_2047,N_1172,N_1159);
and U2048 (N_2048,N_1789,N_1155);
or U2049 (N_2049,N_1455,N_1356);
and U2050 (N_2050,N_1898,N_1536);
or U2051 (N_2051,N_1595,N_1611);
nand U2052 (N_2052,N_1641,N_1314);
and U2053 (N_2053,N_1971,N_1493);
nor U2054 (N_2054,N_1348,N_1344);
xnor U2055 (N_2055,N_1687,N_1319);
xor U2056 (N_2056,N_1680,N_1488);
nor U2057 (N_2057,N_1917,N_1904);
and U2058 (N_2058,N_1713,N_1918);
nand U2059 (N_2059,N_1830,N_1198);
or U2060 (N_2060,N_1506,N_1735);
or U2061 (N_2061,N_1338,N_1950);
and U2062 (N_2062,N_1258,N_1009);
and U2063 (N_2063,N_1832,N_1248);
nor U2064 (N_2064,N_1092,N_1805);
nor U2065 (N_2065,N_1632,N_1889);
or U2066 (N_2066,N_1125,N_1275);
or U2067 (N_2067,N_1865,N_1402);
and U2068 (N_2068,N_1041,N_1384);
and U2069 (N_2069,N_1428,N_1812);
nor U2070 (N_2070,N_1160,N_1145);
nor U2071 (N_2071,N_1867,N_1647);
xnor U2072 (N_2072,N_1414,N_1522);
nor U2073 (N_2073,N_1597,N_1018);
or U2074 (N_2074,N_1241,N_1880);
nor U2075 (N_2075,N_1855,N_1580);
nand U2076 (N_2076,N_1602,N_1860);
nor U2077 (N_2077,N_1086,N_1502);
xor U2078 (N_2078,N_1922,N_1759);
nand U2079 (N_2079,N_1001,N_1093);
nor U2080 (N_2080,N_1625,N_1127);
or U2081 (N_2081,N_1840,N_1841);
and U2082 (N_2082,N_1355,N_1471);
nor U2083 (N_2083,N_1755,N_1521);
nand U2084 (N_2084,N_1774,N_1507);
nor U2085 (N_2085,N_1704,N_1073);
nand U2086 (N_2086,N_1505,N_1834);
or U2087 (N_2087,N_1386,N_1391);
and U2088 (N_2088,N_1622,N_1036);
nor U2089 (N_2089,N_1788,N_1820);
and U2090 (N_2090,N_1328,N_1666);
or U2091 (N_2091,N_1295,N_1106);
nor U2092 (N_2092,N_1088,N_1469);
nand U2093 (N_2093,N_1431,N_1465);
or U2094 (N_2094,N_1977,N_1104);
nand U2095 (N_2095,N_1070,N_1555);
xnor U2096 (N_2096,N_1381,N_1362);
or U2097 (N_2097,N_1287,N_1944);
nor U2098 (N_2098,N_1993,N_1905);
and U2099 (N_2099,N_1615,N_1607);
and U2100 (N_2100,N_1091,N_1531);
or U2101 (N_2101,N_1445,N_1643);
nor U2102 (N_2102,N_1177,N_1161);
or U2103 (N_2103,N_1686,N_1285);
nand U2104 (N_2104,N_1960,N_1770);
or U2105 (N_2105,N_1875,N_1153);
nor U2106 (N_2106,N_1722,N_1806);
nor U2107 (N_2107,N_1667,N_1300);
and U2108 (N_2108,N_1137,N_1736);
nor U2109 (N_2109,N_1985,N_1173);
nor U2110 (N_2110,N_1183,N_1417);
nor U2111 (N_2111,N_1236,N_1911);
xnor U2112 (N_2112,N_1289,N_1079);
and U2113 (N_2113,N_1574,N_1273);
nand U2114 (N_2114,N_1863,N_1364);
nor U2115 (N_2115,N_1550,N_1347);
and U2116 (N_2116,N_1101,N_1180);
nand U2117 (N_2117,N_1665,N_1162);
nand U2118 (N_2118,N_1371,N_1283);
xnor U2119 (N_2119,N_1113,N_1901);
or U2120 (N_2120,N_1668,N_1475);
nor U2121 (N_2121,N_1930,N_1115);
or U2122 (N_2122,N_1752,N_1782);
and U2123 (N_2123,N_1120,N_1067);
or U2124 (N_2124,N_1608,N_1599);
nor U2125 (N_2125,N_1128,N_1938);
nor U2126 (N_2126,N_1591,N_1884);
nand U2127 (N_2127,N_1261,N_1886);
nand U2128 (N_2128,N_1872,N_1981);
and U2129 (N_2129,N_1123,N_1339);
nor U2130 (N_2130,N_1225,N_1354);
nor U2131 (N_2131,N_1111,N_1743);
and U2132 (N_2132,N_1439,N_1263);
nand U2133 (N_2133,N_1754,N_1682);
and U2134 (N_2134,N_1685,N_1166);
or U2135 (N_2135,N_1108,N_1621);
nand U2136 (N_2136,N_1022,N_1891);
or U2137 (N_2137,N_1728,N_1786);
and U2138 (N_2138,N_1819,N_1916);
and U2139 (N_2139,N_1485,N_1209);
nor U2140 (N_2140,N_1071,N_1213);
or U2141 (N_2141,N_1017,N_1560);
or U2142 (N_2142,N_1673,N_1228);
or U2143 (N_2143,N_1274,N_1363);
or U2144 (N_2144,N_1634,N_1481);
nor U2145 (N_2145,N_1970,N_1807);
or U2146 (N_2146,N_1698,N_1244);
or U2147 (N_2147,N_1633,N_1318);
or U2148 (N_2148,N_1185,N_1370);
or U2149 (N_2149,N_1112,N_1216);
nor U2150 (N_2150,N_1604,N_1656);
nand U2151 (N_2151,N_1031,N_1352);
nor U2152 (N_2152,N_1179,N_1672);
nand U2153 (N_2153,N_1498,N_1188);
and U2154 (N_2154,N_1503,N_1897);
or U2155 (N_2155,N_1497,N_1007);
nor U2156 (N_2156,N_1046,N_1936);
nand U2157 (N_2157,N_1327,N_1947);
and U2158 (N_2158,N_1233,N_1742);
nand U2159 (N_2159,N_1330,N_1231);
and U2160 (N_2160,N_1773,N_1764);
and U2161 (N_2161,N_1353,N_1978);
and U2162 (N_2162,N_1584,N_1114);
or U2163 (N_2163,N_1854,N_1098);
and U2164 (N_2164,N_1549,N_1677);
xnor U2165 (N_2165,N_1477,N_1110);
nand U2166 (N_2166,N_1868,N_1492);
nand U2167 (N_2167,N_1661,N_1598);
nor U2168 (N_2168,N_1286,N_1839);
or U2169 (N_2169,N_1249,N_1878);
nor U2170 (N_2170,N_1674,N_1824);
and U2171 (N_2171,N_1470,N_1271);
and U2172 (N_2172,N_1519,N_1077);
or U2173 (N_2173,N_1660,N_1652);
nor U2174 (N_2174,N_1545,N_1546);
or U2175 (N_2175,N_1190,N_1421);
or U2176 (N_2176,N_1730,N_1590);
nor U2177 (N_2177,N_1227,N_1450);
or U2178 (N_2178,N_1058,N_1606);
or U2179 (N_2179,N_1044,N_1721);
and U2180 (N_2180,N_1026,N_1281);
nor U2181 (N_2181,N_1395,N_1818);
nor U2182 (N_2182,N_1659,N_1746);
nand U2183 (N_2183,N_1954,N_1593);
nand U2184 (N_2184,N_1403,N_1030);
xor U2185 (N_2185,N_1826,N_1520);
nor U2186 (N_2186,N_1415,N_1939);
or U2187 (N_2187,N_1202,N_1557);
nand U2188 (N_2188,N_1468,N_1849);
nand U2189 (N_2189,N_1122,N_1929);
nand U2190 (N_2190,N_1055,N_1577);
nor U2191 (N_2191,N_1695,N_1684);
and U2192 (N_2192,N_1000,N_1534);
nor U2193 (N_2193,N_1511,N_1131);
nor U2194 (N_2194,N_1585,N_1424);
and U2195 (N_2195,N_1637,N_1252);
xnor U2196 (N_2196,N_1257,N_1940);
nor U2197 (N_2197,N_1164,N_1825);
or U2198 (N_2198,N_1053,N_1215);
xnor U2199 (N_2199,N_1156,N_1544);
nand U2200 (N_2200,N_1050,N_1116);
nor U2201 (N_2201,N_1847,N_1887);
and U2202 (N_2202,N_1696,N_1442);
nand U2203 (N_2203,N_1361,N_1956);
or U2204 (N_2204,N_1010,N_1836);
nor U2205 (N_2205,N_1459,N_1799);
or U2206 (N_2206,N_1397,N_1394);
or U2207 (N_2207,N_1121,N_1034);
and U2208 (N_2208,N_1254,N_1988);
xnor U2209 (N_2209,N_1206,N_1928);
nor U2210 (N_2210,N_1613,N_1946);
or U2211 (N_2211,N_1045,N_1943);
nand U2212 (N_2212,N_1547,N_1199);
nor U2213 (N_2213,N_1035,N_1890);
or U2214 (N_2214,N_1351,N_1738);
nand U2215 (N_2215,N_1303,N_1279);
or U2216 (N_2216,N_1298,N_1435);
or U2217 (N_2217,N_1229,N_1269);
and U2218 (N_2218,N_1676,N_1766);
nor U2219 (N_2219,N_1678,N_1136);
and U2220 (N_2220,N_1908,N_1080);
nor U2221 (N_2221,N_1107,N_1749);
and U2222 (N_2222,N_1389,N_1725);
or U2223 (N_2223,N_1013,N_1264);
nor U2224 (N_2224,N_1772,N_1804);
nor U2225 (N_2225,N_1959,N_1925);
and U2226 (N_2226,N_1334,N_1478);
nor U2227 (N_2227,N_1801,N_1657);
nor U2228 (N_2228,N_1496,N_1425);
and U2229 (N_2229,N_1484,N_1627);
nor U2230 (N_2230,N_1163,N_1130);
nor U2231 (N_2231,N_1785,N_1603);
and U2232 (N_2232,N_1433,N_1167);
or U2233 (N_2233,N_1902,N_1513);
nand U2234 (N_2234,N_1187,N_1175);
or U2235 (N_2235,N_1765,N_1638);
nand U2236 (N_2236,N_1095,N_1802);
or U2237 (N_2237,N_1320,N_1640);
nand U2238 (N_2238,N_1491,N_1259);
nand U2239 (N_2239,N_1192,N_1196);
nor U2240 (N_2240,N_1452,N_1941);
xor U2241 (N_2241,N_1336,N_1821);
nor U2242 (N_2242,N_1831,N_1124);
nor U2243 (N_2243,N_1420,N_1313);
or U2244 (N_2244,N_1135,N_1618);
and U2245 (N_2245,N_1998,N_1702);
or U2246 (N_2246,N_1942,N_1787);
and U2247 (N_2247,N_1623,N_1480);
or U2248 (N_2248,N_1170,N_1800);
nor U2249 (N_2249,N_1552,N_1078);
nand U2250 (N_2250,N_1518,N_1975);
nor U2251 (N_2251,N_1919,N_1692);
nand U2252 (N_2252,N_1588,N_1311);
nand U2253 (N_2253,N_1316,N_1870);
nor U2254 (N_2254,N_1490,N_1152);
nor U2255 (N_2255,N_1064,N_1845);
or U2256 (N_2256,N_1235,N_1655);
and U2257 (N_2257,N_1609,N_1043);
or U2258 (N_2258,N_1143,N_1768);
nor U2259 (N_2259,N_1012,N_1138);
or U2260 (N_2260,N_1457,N_1413);
nor U2261 (N_2261,N_1957,N_1208);
or U2262 (N_2262,N_1232,N_1063);
and U2263 (N_2263,N_1679,N_1842);
nor U2264 (N_2264,N_1541,N_1983);
nand U2265 (N_2265,N_1750,N_1935);
or U2266 (N_2266,N_1329,N_1587);
xnor U2267 (N_2267,N_1157,N_1504);
or U2268 (N_2268,N_1987,N_1008);
nand U2269 (N_2269,N_1990,N_1027);
and U2270 (N_2270,N_1482,N_1195);
and U2271 (N_2271,N_1129,N_1494);
or U2272 (N_2272,N_1011,N_1406);
nor U2273 (N_2273,N_1948,N_1630);
and U2274 (N_2274,N_1817,N_1463);
or U2275 (N_2275,N_1379,N_1489);
and U2276 (N_2276,N_1999,N_1974);
or U2277 (N_2277,N_1048,N_1284);
and U2278 (N_2278,N_1247,N_1601);
and U2279 (N_2279,N_1893,N_1461);
and U2280 (N_2280,N_1958,N_1649);
or U2281 (N_2281,N_1920,N_1432);
nor U2282 (N_2282,N_1853,N_1714);
and U2283 (N_2283,N_1301,N_1631);
and U2284 (N_2284,N_1270,N_1299);
nor U2285 (N_2285,N_1392,N_1462);
nor U2286 (N_2286,N_1575,N_1572);
and U2287 (N_2287,N_1539,N_1103);
nand U2288 (N_2288,N_1382,N_1210);
and U2289 (N_2289,N_1732,N_1510);
and U2290 (N_2290,N_1533,N_1951);
and U2291 (N_2291,N_1811,N_1097);
nand U2292 (N_2292,N_1671,N_1927);
nand U2293 (N_2293,N_1553,N_1385);
and U2294 (N_2294,N_1201,N_1059);
nand U2295 (N_2295,N_1892,N_1790);
and U2296 (N_2296,N_1085,N_1816);
nor U2297 (N_2297,N_1761,N_1896);
and U2298 (N_2298,N_1029,N_1296);
nand U2299 (N_2299,N_1047,N_1345);
nor U2300 (N_2300,N_1610,N_1038);
or U2301 (N_2301,N_1332,N_1322);
nor U2302 (N_2302,N_1002,N_1224);
nor U2303 (N_2303,N_1551,N_1877);
or U2304 (N_2304,N_1423,N_1873);
or U2305 (N_2305,N_1653,N_1566);
nand U2306 (N_2306,N_1856,N_1061);
nor U2307 (N_2307,N_1969,N_1844);
or U2308 (N_2308,N_1912,N_1858);
nand U2309 (N_2309,N_1084,N_1813);
and U2310 (N_2310,N_1105,N_1570);
nor U2311 (N_2311,N_1509,N_1744);
nand U2312 (N_2312,N_1723,N_1068);
or U2313 (N_2313,N_1616,N_1250);
nand U2314 (N_2314,N_1838,N_1784);
or U2315 (N_2315,N_1315,N_1537);
xnor U2316 (N_2316,N_1437,N_1524);
and U2317 (N_2317,N_1165,N_1052);
nand U2318 (N_2318,N_1447,N_1083);
nor U2319 (N_2319,N_1717,N_1791);
and U2320 (N_2320,N_1374,N_1952);
nor U2321 (N_2321,N_1532,N_1234);
xnor U2322 (N_2322,N_1184,N_1454);
and U2323 (N_2323,N_1760,N_1094);
nand U2324 (N_2324,N_1973,N_1543);
nand U2325 (N_2325,N_1751,N_1132);
nor U2326 (N_2326,N_1238,N_1343);
nand U2327 (N_2327,N_1317,N_1724);
nor U2328 (N_2328,N_1268,N_1240);
and U2329 (N_2329,N_1745,N_1823);
and U2330 (N_2330,N_1340,N_1561);
or U2331 (N_2331,N_1563,N_1848);
nand U2332 (N_2332,N_1049,N_1310);
nand U2333 (N_2333,N_1866,N_1358);
or U2334 (N_2334,N_1573,N_1769);
or U2335 (N_2335,N_1369,N_1843);
nor U2336 (N_2336,N_1562,N_1777);
or U2337 (N_2337,N_1367,N_1222);
nor U2338 (N_2338,N_1203,N_1168);
nor U2339 (N_2339,N_1473,N_1449);
and U2340 (N_2340,N_1357,N_1501);
nand U2341 (N_2341,N_1635,N_1133);
or U2342 (N_2342,N_1794,N_1458);
or U2343 (N_2343,N_1906,N_1378);
and U2344 (N_2344,N_1102,N_1715);
nor U2345 (N_2345,N_1582,N_1991);
and U2346 (N_2346,N_1278,N_1376);
xnor U2347 (N_2347,N_1057,N_1926);
or U2348 (N_2348,N_1408,N_1151);
nand U2349 (N_2349,N_1835,N_1576);
and U2350 (N_2350,N_1737,N_1780);
nor U2351 (N_2351,N_1705,N_1962);
nand U2352 (N_2352,N_1251,N_1953);
nand U2353 (N_2353,N_1410,N_1016);
and U2354 (N_2354,N_1218,N_1483);
nor U2355 (N_2355,N_1372,N_1174);
and U2356 (N_2356,N_1014,N_1072);
and U2357 (N_2357,N_1747,N_1400);
nand U2358 (N_2358,N_1879,N_1359);
nand U2359 (N_2359,N_1346,N_1099);
nand U2360 (N_2360,N_1663,N_1932);
nand U2361 (N_2361,N_1383,N_1689);
or U2362 (N_2362,N_1583,N_1337);
nand U2363 (N_2363,N_1109,N_1644);
nand U2364 (N_2364,N_1645,N_1523);
and U2365 (N_2365,N_1910,N_1642);
nor U2366 (N_2366,N_1419,N_1568);
and U2367 (N_2367,N_1792,N_1479);
and U2368 (N_2368,N_1388,N_1795);
or U2369 (N_2369,N_1629,N_1793);
or U2370 (N_2370,N_1054,N_1324);
and U2371 (N_2371,N_1683,N_1288);
nor U2372 (N_2372,N_1390,N_1538);
and U2373 (N_2373,N_1144,N_1476);
nand U2374 (N_2374,N_1894,N_1416);
nand U2375 (N_2375,N_1828,N_1592);
and U2376 (N_2376,N_1528,N_1142);
and U2377 (N_2377,N_1976,N_1422);
nor U2378 (N_2378,N_1277,N_1670);
nand U2379 (N_2379,N_1335,N_1741);
or U2380 (N_2380,N_1411,N_1967);
and U2381 (N_2381,N_1846,N_1700);
nor U2382 (N_2382,N_1945,N_1056);
nand U2383 (N_2383,N_1727,N_1596);
and U2384 (N_2384,N_1526,N_1965);
nand U2385 (N_2385,N_1815,N_1617);
nand U2386 (N_2386,N_1032,N_1681);
or U2387 (N_2387,N_1963,N_1720);
nand U2388 (N_2388,N_1852,N_1396);
nor U2389 (N_2389,N_1822,N_1207);
nor U2390 (N_2390,N_1719,N_1694);
nand U2391 (N_2391,N_1626,N_1972);
or U2392 (N_2392,N_1827,N_1669);
or U2393 (N_2393,N_1748,N_1753);
xor U2394 (N_2394,N_1189,N_1986);
nand U2395 (N_2395,N_1350,N_1193);
nor U2396 (N_2396,N_1140,N_1899);
nand U2397 (N_2397,N_1857,N_1443);
or U2398 (N_2398,N_1290,N_1467);
nand U2399 (N_2399,N_1141,N_1305);
nor U2400 (N_2400,N_1434,N_1375);
and U2401 (N_2401,N_1255,N_1486);
nor U2402 (N_2402,N_1808,N_1226);
nand U2403 (N_2403,N_1304,N_1349);
and U2404 (N_2404,N_1589,N_1262);
nand U2405 (N_2405,N_1581,N_1578);
nor U2406 (N_2406,N_1903,N_1451);
nand U2407 (N_2407,N_1331,N_1859);
nand U2408 (N_2408,N_1675,N_1874);
nor U2409 (N_2409,N_1096,N_1961);
nor U2410 (N_2410,N_1292,N_1763);
and U2411 (N_2411,N_1243,N_1688);
or U2412 (N_2412,N_1851,N_1924);
and U2413 (N_2413,N_1438,N_1024);
and U2414 (N_2414,N_1542,N_1150);
nand U2415 (N_2415,N_1307,N_1933);
nor U2416 (N_2416,N_1246,N_1139);
nor U2417 (N_2417,N_1186,N_1312);
and U2418 (N_2418,N_1810,N_1181);
or U2419 (N_2419,N_1237,N_1540);
nand U2420 (N_2420,N_1089,N_1075);
nand U2421 (N_2421,N_1282,N_1134);
nand U2422 (N_2422,N_1711,N_1914);
nand U2423 (N_2423,N_1326,N_1366);
nor U2424 (N_2424,N_1015,N_1444);
and U2425 (N_2425,N_1025,N_1517);
xor U2426 (N_2426,N_1636,N_1387);
or U2427 (N_2427,N_1321,N_1512);
nor U2428 (N_2428,N_1266,N_1559);
or U2429 (N_2429,N_1260,N_1797);
nand U2430 (N_2430,N_1734,N_1600);
nor U2431 (N_2431,N_1515,N_1418);
nand U2432 (N_2432,N_1076,N_1966);
nor U2433 (N_2433,N_1814,N_1876);
nand U2434 (N_2434,N_1205,N_1508);
nor U2435 (N_2435,N_1221,N_1620);
and U2436 (N_2436,N_1619,N_1360);
and U2437 (N_2437,N_1882,N_1119);
or U2438 (N_2438,N_1474,N_1323);
or U2439 (N_2439,N_1276,N_1850);
nor U2440 (N_2440,N_1100,N_1907);
or U2441 (N_2441,N_1558,N_1309);
nor U2442 (N_2442,N_1783,N_1756);
nand U2443 (N_2443,N_1658,N_1781);
and U2444 (N_2444,N_1569,N_1214);
or U2445 (N_2445,N_1567,N_1639);
and U2446 (N_2446,N_1293,N_1968);
nand U2447 (N_2447,N_1333,N_1900);
and U2448 (N_2448,N_1003,N_1466);
nand U2449 (N_2449,N_1861,N_1837);
nand U2450 (N_2450,N_1516,N_1499);
nor U2451 (N_2451,N_1005,N_1650);
and U2452 (N_2452,N_1341,N_1514);
nand U2453 (N_2453,N_1306,N_1994);
nand U2454 (N_2454,N_1242,N_1796);
nand U2455 (N_2455,N_1798,N_1280);
xnor U2456 (N_2456,N_1762,N_1373);
and U2457 (N_2457,N_1779,N_1803);
or U2458 (N_2458,N_1019,N_1571);
or U2459 (N_2459,N_1556,N_1809);
or U2460 (N_2460,N_1117,N_1701);
nand U2461 (N_2461,N_1087,N_1923);
nor U2462 (N_2462,N_1169,N_1377);
nor U2463 (N_2463,N_1154,N_1885);
nor U2464 (N_2464,N_1245,N_1495);
nor U2465 (N_2465,N_1342,N_1586);
or U2466 (N_2466,N_1404,N_1915);
nor U2467 (N_2467,N_1729,N_1398);
nor U2468 (N_2468,N_1757,N_1934);
nand U2469 (N_2469,N_1297,N_1037);
nand U2470 (N_2470,N_1883,N_1066);
nand U2471 (N_2471,N_1706,N_1464);
or U2472 (N_2472,N_1409,N_1648);
nand U2473 (N_2473,N_1699,N_1006);
nor U2474 (N_2474,N_1895,N_1040);
nor U2475 (N_2475,N_1997,N_1869);
nor U2476 (N_2476,N_1771,N_1651);
and U2477 (N_2477,N_1182,N_1982);
nor U2478 (N_2478,N_1697,N_1020);
or U2479 (N_2479,N_1881,N_1535);
nand U2480 (N_2480,N_1440,N_1042);
or U2481 (N_2481,N_1964,N_1060);
nor U2482 (N_2482,N_1996,N_1758);
and U2483 (N_2483,N_1253,N_1302);
nor U2484 (N_2484,N_1707,N_1888);
nand U2485 (N_2485,N_1628,N_1456);
and U2486 (N_2486,N_1039,N_1775);
nor U2487 (N_2487,N_1937,N_1291);
nor U2488 (N_2488,N_1871,N_1176);
nand U2489 (N_2489,N_1308,N_1529);
and U2490 (N_2490,N_1460,N_1118);
xor U2491 (N_2491,N_1368,N_1949);
and U2492 (N_2492,N_1646,N_1548);
nand U2493 (N_2493,N_1220,N_1525);
nor U2494 (N_2494,N_1995,N_1294);
or U2495 (N_2495,N_1921,N_1955);
and U2496 (N_2496,N_1778,N_1733);
and U2497 (N_2497,N_1931,N_1710);
nor U2498 (N_2498,N_1212,N_1527);
nand U2499 (N_2499,N_1980,N_1500);
and U2500 (N_2500,N_1522,N_1435);
and U2501 (N_2501,N_1678,N_1939);
nand U2502 (N_2502,N_1046,N_1522);
nand U2503 (N_2503,N_1402,N_1107);
nor U2504 (N_2504,N_1109,N_1478);
or U2505 (N_2505,N_1923,N_1778);
nor U2506 (N_2506,N_1301,N_1332);
and U2507 (N_2507,N_1406,N_1140);
nor U2508 (N_2508,N_1409,N_1456);
nor U2509 (N_2509,N_1871,N_1705);
nor U2510 (N_2510,N_1027,N_1731);
nor U2511 (N_2511,N_1699,N_1437);
or U2512 (N_2512,N_1518,N_1973);
and U2513 (N_2513,N_1409,N_1487);
nor U2514 (N_2514,N_1008,N_1909);
nand U2515 (N_2515,N_1413,N_1868);
and U2516 (N_2516,N_1830,N_1280);
or U2517 (N_2517,N_1113,N_1740);
or U2518 (N_2518,N_1033,N_1139);
nand U2519 (N_2519,N_1905,N_1138);
nand U2520 (N_2520,N_1966,N_1091);
nor U2521 (N_2521,N_1447,N_1359);
nor U2522 (N_2522,N_1354,N_1718);
nand U2523 (N_2523,N_1666,N_1133);
and U2524 (N_2524,N_1015,N_1944);
nand U2525 (N_2525,N_1230,N_1203);
nor U2526 (N_2526,N_1843,N_1364);
and U2527 (N_2527,N_1951,N_1014);
nand U2528 (N_2528,N_1257,N_1355);
or U2529 (N_2529,N_1154,N_1163);
and U2530 (N_2530,N_1518,N_1269);
nor U2531 (N_2531,N_1529,N_1468);
nor U2532 (N_2532,N_1438,N_1151);
nand U2533 (N_2533,N_1092,N_1579);
nor U2534 (N_2534,N_1829,N_1865);
nor U2535 (N_2535,N_1637,N_1479);
nand U2536 (N_2536,N_1371,N_1982);
xor U2537 (N_2537,N_1241,N_1194);
nand U2538 (N_2538,N_1299,N_1616);
or U2539 (N_2539,N_1573,N_1376);
and U2540 (N_2540,N_1995,N_1539);
or U2541 (N_2541,N_1100,N_1191);
nor U2542 (N_2542,N_1801,N_1332);
nor U2543 (N_2543,N_1462,N_1686);
nand U2544 (N_2544,N_1025,N_1063);
or U2545 (N_2545,N_1723,N_1980);
and U2546 (N_2546,N_1038,N_1379);
nor U2547 (N_2547,N_1621,N_1114);
nand U2548 (N_2548,N_1470,N_1063);
nor U2549 (N_2549,N_1590,N_1259);
nand U2550 (N_2550,N_1358,N_1558);
nand U2551 (N_2551,N_1262,N_1187);
or U2552 (N_2552,N_1809,N_1109);
nor U2553 (N_2553,N_1168,N_1115);
or U2554 (N_2554,N_1114,N_1463);
nand U2555 (N_2555,N_1582,N_1328);
nand U2556 (N_2556,N_1973,N_1169);
nand U2557 (N_2557,N_1745,N_1023);
nor U2558 (N_2558,N_1708,N_1538);
and U2559 (N_2559,N_1856,N_1210);
and U2560 (N_2560,N_1040,N_1201);
nor U2561 (N_2561,N_1616,N_1405);
nand U2562 (N_2562,N_1885,N_1554);
nand U2563 (N_2563,N_1863,N_1795);
and U2564 (N_2564,N_1347,N_1620);
and U2565 (N_2565,N_1506,N_1438);
nand U2566 (N_2566,N_1560,N_1309);
and U2567 (N_2567,N_1097,N_1939);
xnor U2568 (N_2568,N_1755,N_1540);
and U2569 (N_2569,N_1902,N_1751);
and U2570 (N_2570,N_1003,N_1234);
nor U2571 (N_2571,N_1434,N_1903);
xor U2572 (N_2572,N_1684,N_1705);
nor U2573 (N_2573,N_1017,N_1550);
nand U2574 (N_2574,N_1342,N_1289);
xor U2575 (N_2575,N_1390,N_1800);
or U2576 (N_2576,N_1306,N_1648);
nand U2577 (N_2577,N_1827,N_1894);
or U2578 (N_2578,N_1032,N_1622);
nor U2579 (N_2579,N_1962,N_1450);
and U2580 (N_2580,N_1521,N_1965);
nand U2581 (N_2581,N_1089,N_1344);
xor U2582 (N_2582,N_1832,N_1856);
nand U2583 (N_2583,N_1767,N_1864);
nor U2584 (N_2584,N_1207,N_1498);
or U2585 (N_2585,N_1464,N_1639);
nor U2586 (N_2586,N_1287,N_1314);
and U2587 (N_2587,N_1461,N_1648);
nand U2588 (N_2588,N_1533,N_1556);
nand U2589 (N_2589,N_1076,N_1996);
and U2590 (N_2590,N_1833,N_1080);
nor U2591 (N_2591,N_1760,N_1592);
or U2592 (N_2592,N_1695,N_1217);
nand U2593 (N_2593,N_1046,N_1166);
nor U2594 (N_2594,N_1472,N_1567);
nand U2595 (N_2595,N_1787,N_1531);
and U2596 (N_2596,N_1968,N_1973);
nand U2597 (N_2597,N_1543,N_1310);
nor U2598 (N_2598,N_1768,N_1062);
and U2599 (N_2599,N_1461,N_1244);
nor U2600 (N_2600,N_1496,N_1181);
xor U2601 (N_2601,N_1696,N_1390);
nor U2602 (N_2602,N_1470,N_1501);
nand U2603 (N_2603,N_1462,N_1494);
nor U2604 (N_2604,N_1340,N_1188);
and U2605 (N_2605,N_1205,N_1141);
or U2606 (N_2606,N_1125,N_1961);
and U2607 (N_2607,N_1946,N_1600);
nor U2608 (N_2608,N_1200,N_1148);
and U2609 (N_2609,N_1760,N_1778);
nand U2610 (N_2610,N_1296,N_1241);
nand U2611 (N_2611,N_1148,N_1828);
nor U2612 (N_2612,N_1262,N_1332);
and U2613 (N_2613,N_1677,N_1872);
or U2614 (N_2614,N_1189,N_1472);
or U2615 (N_2615,N_1828,N_1648);
and U2616 (N_2616,N_1199,N_1600);
nand U2617 (N_2617,N_1523,N_1192);
nor U2618 (N_2618,N_1109,N_1967);
nand U2619 (N_2619,N_1909,N_1206);
nand U2620 (N_2620,N_1370,N_1668);
or U2621 (N_2621,N_1396,N_1847);
nor U2622 (N_2622,N_1473,N_1176);
nor U2623 (N_2623,N_1079,N_1795);
or U2624 (N_2624,N_1831,N_1500);
nand U2625 (N_2625,N_1647,N_1735);
and U2626 (N_2626,N_1823,N_1194);
nand U2627 (N_2627,N_1384,N_1845);
nand U2628 (N_2628,N_1494,N_1205);
xor U2629 (N_2629,N_1575,N_1925);
and U2630 (N_2630,N_1136,N_1179);
or U2631 (N_2631,N_1496,N_1134);
or U2632 (N_2632,N_1191,N_1244);
or U2633 (N_2633,N_1763,N_1042);
or U2634 (N_2634,N_1773,N_1186);
or U2635 (N_2635,N_1427,N_1334);
nor U2636 (N_2636,N_1785,N_1912);
or U2637 (N_2637,N_1682,N_1278);
or U2638 (N_2638,N_1842,N_1002);
nand U2639 (N_2639,N_1725,N_1189);
and U2640 (N_2640,N_1289,N_1596);
or U2641 (N_2641,N_1918,N_1344);
xnor U2642 (N_2642,N_1047,N_1310);
and U2643 (N_2643,N_1308,N_1403);
nand U2644 (N_2644,N_1442,N_1165);
nand U2645 (N_2645,N_1506,N_1818);
nand U2646 (N_2646,N_1029,N_1689);
nand U2647 (N_2647,N_1677,N_1914);
or U2648 (N_2648,N_1927,N_1986);
and U2649 (N_2649,N_1291,N_1837);
nor U2650 (N_2650,N_1964,N_1897);
and U2651 (N_2651,N_1803,N_1368);
nor U2652 (N_2652,N_1325,N_1740);
nor U2653 (N_2653,N_1305,N_1403);
or U2654 (N_2654,N_1341,N_1411);
nand U2655 (N_2655,N_1607,N_1087);
nand U2656 (N_2656,N_1417,N_1866);
nor U2657 (N_2657,N_1666,N_1071);
nor U2658 (N_2658,N_1211,N_1177);
or U2659 (N_2659,N_1020,N_1009);
and U2660 (N_2660,N_1765,N_1520);
nor U2661 (N_2661,N_1871,N_1852);
and U2662 (N_2662,N_1790,N_1755);
nand U2663 (N_2663,N_1420,N_1190);
nand U2664 (N_2664,N_1388,N_1521);
or U2665 (N_2665,N_1000,N_1759);
nor U2666 (N_2666,N_1840,N_1577);
xor U2667 (N_2667,N_1199,N_1553);
and U2668 (N_2668,N_1549,N_1849);
and U2669 (N_2669,N_1121,N_1702);
nor U2670 (N_2670,N_1627,N_1535);
and U2671 (N_2671,N_1973,N_1794);
or U2672 (N_2672,N_1934,N_1272);
nand U2673 (N_2673,N_1839,N_1048);
nand U2674 (N_2674,N_1223,N_1133);
or U2675 (N_2675,N_1171,N_1733);
nor U2676 (N_2676,N_1285,N_1659);
or U2677 (N_2677,N_1247,N_1633);
or U2678 (N_2678,N_1201,N_1795);
nor U2679 (N_2679,N_1877,N_1897);
nor U2680 (N_2680,N_1695,N_1731);
nor U2681 (N_2681,N_1189,N_1364);
nor U2682 (N_2682,N_1275,N_1468);
nand U2683 (N_2683,N_1672,N_1573);
nand U2684 (N_2684,N_1452,N_1798);
nand U2685 (N_2685,N_1949,N_1917);
or U2686 (N_2686,N_1068,N_1229);
nor U2687 (N_2687,N_1365,N_1425);
and U2688 (N_2688,N_1294,N_1008);
or U2689 (N_2689,N_1444,N_1982);
nand U2690 (N_2690,N_1751,N_1429);
nor U2691 (N_2691,N_1733,N_1669);
and U2692 (N_2692,N_1490,N_1171);
nor U2693 (N_2693,N_1292,N_1271);
nand U2694 (N_2694,N_1769,N_1485);
or U2695 (N_2695,N_1866,N_1517);
nor U2696 (N_2696,N_1007,N_1127);
or U2697 (N_2697,N_1294,N_1442);
nor U2698 (N_2698,N_1650,N_1329);
nor U2699 (N_2699,N_1438,N_1016);
nor U2700 (N_2700,N_1809,N_1916);
nor U2701 (N_2701,N_1566,N_1658);
nand U2702 (N_2702,N_1150,N_1921);
and U2703 (N_2703,N_1324,N_1623);
or U2704 (N_2704,N_1436,N_1663);
nor U2705 (N_2705,N_1290,N_1272);
nor U2706 (N_2706,N_1522,N_1995);
or U2707 (N_2707,N_1962,N_1646);
and U2708 (N_2708,N_1526,N_1157);
nand U2709 (N_2709,N_1745,N_1270);
and U2710 (N_2710,N_1621,N_1589);
or U2711 (N_2711,N_1137,N_1655);
nor U2712 (N_2712,N_1951,N_1981);
and U2713 (N_2713,N_1741,N_1299);
nand U2714 (N_2714,N_1456,N_1104);
or U2715 (N_2715,N_1287,N_1422);
or U2716 (N_2716,N_1959,N_1768);
and U2717 (N_2717,N_1846,N_1788);
or U2718 (N_2718,N_1467,N_1140);
nand U2719 (N_2719,N_1966,N_1594);
and U2720 (N_2720,N_1381,N_1016);
and U2721 (N_2721,N_1637,N_1737);
nor U2722 (N_2722,N_1753,N_1584);
nor U2723 (N_2723,N_1198,N_1540);
and U2724 (N_2724,N_1964,N_1451);
nor U2725 (N_2725,N_1723,N_1580);
and U2726 (N_2726,N_1074,N_1539);
nand U2727 (N_2727,N_1162,N_1816);
and U2728 (N_2728,N_1164,N_1884);
or U2729 (N_2729,N_1847,N_1809);
or U2730 (N_2730,N_1007,N_1818);
and U2731 (N_2731,N_1205,N_1748);
nor U2732 (N_2732,N_1267,N_1259);
and U2733 (N_2733,N_1508,N_1080);
nor U2734 (N_2734,N_1648,N_1358);
and U2735 (N_2735,N_1769,N_1386);
nand U2736 (N_2736,N_1553,N_1405);
or U2737 (N_2737,N_1522,N_1576);
nand U2738 (N_2738,N_1091,N_1019);
nand U2739 (N_2739,N_1401,N_1898);
or U2740 (N_2740,N_1693,N_1434);
nand U2741 (N_2741,N_1145,N_1105);
xnor U2742 (N_2742,N_1877,N_1007);
and U2743 (N_2743,N_1219,N_1197);
and U2744 (N_2744,N_1675,N_1808);
nor U2745 (N_2745,N_1267,N_1561);
or U2746 (N_2746,N_1077,N_1318);
nor U2747 (N_2747,N_1858,N_1580);
and U2748 (N_2748,N_1712,N_1610);
and U2749 (N_2749,N_1295,N_1954);
nand U2750 (N_2750,N_1174,N_1693);
nand U2751 (N_2751,N_1855,N_1871);
nor U2752 (N_2752,N_1366,N_1819);
or U2753 (N_2753,N_1309,N_1137);
and U2754 (N_2754,N_1876,N_1788);
and U2755 (N_2755,N_1506,N_1228);
and U2756 (N_2756,N_1617,N_1609);
nor U2757 (N_2757,N_1387,N_1504);
and U2758 (N_2758,N_1594,N_1820);
nor U2759 (N_2759,N_1825,N_1545);
or U2760 (N_2760,N_1265,N_1895);
or U2761 (N_2761,N_1506,N_1979);
and U2762 (N_2762,N_1498,N_1094);
or U2763 (N_2763,N_1859,N_1108);
or U2764 (N_2764,N_1565,N_1063);
and U2765 (N_2765,N_1429,N_1796);
nand U2766 (N_2766,N_1656,N_1053);
and U2767 (N_2767,N_1096,N_1731);
nor U2768 (N_2768,N_1534,N_1096);
nand U2769 (N_2769,N_1913,N_1152);
nand U2770 (N_2770,N_1933,N_1567);
nor U2771 (N_2771,N_1882,N_1961);
and U2772 (N_2772,N_1687,N_1343);
nor U2773 (N_2773,N_1036,N_1104);
and U2774 (N_2774,N_1779,N_1331);
and U2775 (N_2775,N_1698,N_1763);
nand U2776 (N_2776,N_1976,N_1919);
nand U2777 (N_2777,N_1453,N_1547);
nor U2778 (N_2778,N_1551,N_1497);
and U2779 (N_2779,N_1461,N_1522);
or U2780 (N_2780,N_1369,N_1887);
nor U2781 (N_2781,N_1148,N_1500);
and U2782 (N_2782,N_1442,N_1148);
nor U2783 (N_2783,N_1799,N_1002);
and U2784 (N_2784,N_1646,N_1381);
or U2785 (N_2785,N_1691,N_1110);
and U2786 (N_2786,N_1563,N_1236);
nor U2787 (N_2787,N_1054,N_1094);
nor U2788 (N_2788,N_1328,N_1591);
nand U2789 (N_2789,N_1699,N_1180);
and U2790 (N_2790,N_1589,N_1489);
and U2791 (N_2791,N_1404,N_1287);
or U2792 (N_2792,N_1021,N_1965);
or U2793 (N_2793,N_1978,N_1990);
or U2794 (N_2794,N_1110,N_1604);
nor U2795 (N_2795,N_1943,N_1298);
and U2796 (N_2796,N_1230,N_1190);
and U2797 (N_2797,N_1249,N_1649);
and U2798 (N_2798,N_1361,N_1798);
nor U2799 (N_2799,N_1594,N_1229);
nand U2800 (N_2800,N_1381,N_1446);
and U2801 (N_2801,N_1501,N_1038);
xnor U2802 (N_2802,N_1750,N_1817);
or U2803 (N_2803,N_1897,N_1885);
or U2804 (N_2804,N_1571,N_1858);
nor U2805 (N_2805,N_1814,N_1277);
and U2806 (N_2806,N_1157,N_1079);
nand U2807 (N_2807,N_1195,N_1798);
and U2808 (N_2808,N_1431,N_1999);
or U2809 (N_2809,N_1210,N_1514);
and U2810 (N_2810,N_1771,N_1383);
and U2811 (N_2811,N_1750,N_1112);
nor U2812 (N_2812,N_1735,N_1486);
xor U2813 (N_2813,N_1507,N_1421);
or U2814 (N_2814,N_1652,N_1023);
nor U2815 (N_2815,N_1738,N_1460);
or U2816 (N_2816,N_1285,N_1761);
xor U2817 (N_2817,N_1447,N_1070);
or U2818 (N_2818,N_1628,N_1107);
nor U2819 (N_2819,N_1797,N_1815);
nand U2820 (N_2820,N_1250,N_1689);
nor U2821 (N_2821,N_1749,N_1900);
xnor U2822 (N_2822,N_1807,N_1030);
and U2823 (N_2823,N_1618,N_1083);
nor U2824 (N_2824,N_1250,N_1948);
nor U2825 (N_2825,N_1344,N_1748);
nand U2826 (N_2826,N_1875,N_1886);
nor U2827 (N_2827,N_1337,N_1766);
nand U2828 (N_2828,N_1527,N_1033);
nand U2829 (N_2829,N_1501,N_1025);
or U2830 (N_2830,N_1166,N_1446);
and U2831 (N_2831,N_1358,N_1529);
nand U2832 (N_2832,N_1739,N_1949);
nor U2833 (N_2833,N_1677,N_1964);
nand U2834 (N_2834,N_1170,N_1206);
nor U2835 (N_2835,N_1616,N_1312);
and U2836 (N_2836,N_1239,N_1841);
or U2837 (N_2837,N_1446,N_1733);
and U2838 (N_2838,N_1110,N_1223);
or U2839 (N_2839,N_1374,N_1317);
and U2840 (N_2840,N_1198,N_1227);
nand U2841 (N_2841,N_1532,N_1856);
or U2842 (N_2842,N_1726,N_1403);
and U2843 (N_2843,N_1766,N_1620);
nor U2844 (N_2844,N_1707,N_1233);
or U2845 (N_2845,N_1252,N_1095);
nand U2846 (N_2846,N_1189,N_1334);
nand U2847 (N_2847,N_1723,N_1636);
or U2848 (N_2848,N_1427,N_1660);
nand U2849 (N_2849,N_1418,N_1012);
and U2850 (N_2850,N_1111,N_1652);
nor U2851 (N_2851,N_1974,N_1143);
or U2852 (N_2852,N_1364,N_1191);
and U2853 (N_2853,N_1895,N_1622);
nand U2854 (N_2854,N_1389,N_1518);
or U2855 (N_2855,N_1087,N_1881);
or U2856 (N_2856,N_1879,N_1776);
nand U2857 (N_2857,N_1008,N_1862);
nand U2858 (N_2858,N_1111,N_1300);
or U2859 (N_2859,N_1117,N_1281);
nor U2860 (N_2860,N_1026,N_1961);
nand U2861 (N_2861,N_1216,N_1204);
and U2862 (N_2862,N_1771,N_1153);
or U2863 (N_2863,N_1119,N_1162);
nor U2864 (N_2864,N_1270,N_1832);
or U2865 (N_2865,N_1163,N_1504);
or U2866 (N_2866,N_1540,N_1497);
and U2867 (N_2867,N_1583,N_1397);
or U2868 (N_2868,N_1078,N_1922);
or U2869 (N_2869,N_1945,N_1112);
and U2870 (N_2870,N_1944,N_1376);
nand U2871 (N_2871,N_1739,N_1144);
nor U2872 (N_2872,N_1295,N_1030);
and U2873 (N_2873,N_1491,N_1216);
and U2874 (N_2874,N_1704,N_1932);
or U2875 (N_2875,N_1798,N_1069);
and U2876 (N_2876,N_1871,N_1359);
nand U2877 (N_2877,N_1490,N_1614);
nor U2878 (N_2878,N_1129,N_1119);
and U2879 (N_2879,N_1873,N_1259);
nor U2880 (N_2880,N_1082,N_1322);
nor U2881 (N_2881,N_1342,N_1807);
and U2882 (N_2882,N_1695,N_1092);
or U2883 (N_2883,N_1048,N_1846);
and U2884 (N_2884,N_1611,N_1479);
nand U2885 (N_2885,N_1491,N_1981);
nor U2886 (N_2886,N_1040,N_1082);
nand U2887 (N_2887,N_1456,N_1214);
or U2888 (N_2888,N_1029,N_1084);
nand U2889 (N_2889,N_1561,N_1741);
nor U2890 (N_2890,N_1815,N_1810);
nand U2891 (N_2891,N_1362,N_1400);
nor U2892 (N_2892,N_1865,N_1310);
or U2893 (N_2893,N_1959,N_1561);
nand U2894 (N_2894,N_1960,N_1580);
or U2895 (N_2895,N_1889,N_1887);
nor U2896 (N_2896,N_1768,N_1586);
nor U2897 (N_2897,N_1728,N_1795);
xor U2898 (N_2898,N_1193,N_1129);
nor U2899 (N_2899,N_1203,N_1797);
or U2900 (N_2900,N_1245,N_1258);
or U2901 (N_2901,N_1025,N_1915);
or U2902 (N_2902,N_1833,N_1930);
and U2903 (N_2903,N_1497,N_1467);
and U2904 (N_2904,N_1491,N_1784);
and U2905 (N_2905,N_1598,N_1057);
nand U2906 (N_2906,N_1276,N_1232);
nand U2907 (N_2907,N_1037,N_1533);
or U2908 (N_2908,N_1428,N_1786);
or U2909 (N_2909,N_1428,N_1966);
nand U2910 (N_2910,N_1474,N_1463);
and U2911 (N_2911,N_1524,N_1317);
and U2912 (N_2912,N_1723,N_1739);
or U2913 (N_2913,N_1563,N_1804);
and U2914 (N_2914,N_1751,N_1792);
and U2915 (N_2915,N_1071,N_1053);
nor U2916 (N_2916,N_1205,N_1076);
or U2917 (N_2917,N_1944,N_1752);
and U2918 (N_2918,N_1866,N_1221);
or U2919 (N_2919,N_1804,N_1571);
nand U2920 (N_2920,N_1820,N_1719);
and U2921 (N_2921,N_1916,N_1968);
or U2922 (N_2922,N_1428,N_1338);
nor U2923 (N_2923,N_1805,N_1924);
or U2924 (N_2924,N_1198,N_1457);
nor U2925 (N_2925,N_1764,N_1125);
nand U2926 (N_2926,N_1576,N_1073);
nand U2927 (N_2927,N_1819,N_1795);
and U2928 (N_2928,N_1353,N_1398);
nor U2929 (N_2929,N_1579,N_1986);
and U2930 (N_2930,N_1525,N_1601);
and U2931 (N_2931,N_1815,N_1785);
and U2932 (N_2932,N_1805,N_1722);
xor U2933 (N_2933,N_1373,N_1736);
and U2934 (N_2934,N_1850,N_1414);
and U2935 (N_2935,N_1318,N_1771);
and U2936 (N_2936,N_1685,N_1517);
nand U2937 (N_2937,N_1920,N_1484);
nand U2938 (N_2938,N_1958,N_1463);
or U2939 (N_2939,N_1321,N_1018);
and U2940 (N_2940,N_1664,N_1666);
or U2941 (N_2941,N_1913,N_1091);
xor U2942 (N_2942,N_1308,N_1524);
xor U2943 (N_2943,N_1472,N_1647);
nand U2944 (N_2944,N_1235,N_1024);
nor U2945 (N_2945,N_1578,N_1552);
or U2946 (N_2946,N_1622,N_1788);
nor U2947 (N_2947,N_1385,N_1230);
or U2948 (N_2948,N_1323,N_1019);
or U2949 (N_2949,N_1760,N_1426);
nand U2950 (N_2950,N_1359,N_1636);
nor U2951 (N_2951,N_1277,N_1519);
nand U2952 (N_2952,N_1969,N_1815);
or U2953 (N_2953,N_1108,N_1863);
nor U2954 (N_2954,N_1291,N_1715);
or U2955 (N_2955,N_1201,N_1562);
nand U2956 (N_2956,N_1356,N_1926);
nor U2957 (N_2957,N_1806,N_1787);
nand U2958 (N_2958,N_1816,N_1881);
or U2959 (N_2959,N_1595,N_1635);
or U2960 (N_2960,N_1960,N_1492);
nand U2961 (N_2961,N_1649,N_1377);
and U2962 (N_2962,N_1175,N_1391);
or U2963 (N_2963,N_1342,N_1820);
or U2964 (N_2964,N_1797,N_1962);
or U2965 (N_2965,N_1222,N_1523);
nand U2966 (N_2966,N_1357,N_1142);
nand U2967 (N_2967,N_1550,N_1660);
or U2968 (N_2968,N_1524,N_1266);
nor U2969 (N_2969,N_1313,N_1509);
or U2970 (N_2970,N_1345,N_1905);
nor U2971 (N_2971,N_1378,N_1020);
and U2972 (N_2972,N_1068,N_1352);
and U2973 (N_2973,N_1189,N_1088);
and U2974 (N_2974,N_1518,N_1356);
nand U2975 (N_2975,N_1463,N_1848);
nor U2976 (N_2976,N_1123,N_1393);
or U2977 (N_2977,N_1239,N_1556);
nand U2978 (N_2978,N_1243,N_1802);
nor U2979 (N_2979,N_1641,N_1115);
nand U2980 (N_2980,N_1765,N_1457);
or U2981 (N_2981,N_1288,N_1951);
nor U2982 (N_2982,N_1625,N_1952);
or U2983 (N_2983,N_1478,N_1185);
nor U2984 (N_2984,N_1975,N_1245);
nand U2985 (N_2985,N_1836,N_1936);
or U2986 (N_2986,N_1803,N_1305);
or U2987 (N_2987,N_1956,N_1838);
or U2988 (N_2988,N_1386,N_1081);
and U2989 (N_2989,N_1297,N_1959);
nand U2990 (N_2990,N_1942,N_1730);
nor U2991 (N_2991,N_1293,N_1151);
or U2992 (N_2992,N_1058,N_1270);
and U2993 (N_2993,N_1780,N_1530);
or U2994 (N_2994,N_1302,N_1584);
and U2995 (N_2995,N_1669,N_1991);
nand U2996 (N_2996,N_1630,N_1200);
nand U2997 (N_2997,N_1611,N_1171);
or U2998 (N_2998,N_1726,N_1490);
and U2999 (N_2999,N_1297,N_1225);
nor UO_0 (O_0,N_2685,N_2893);
nand UO_1 (O_1,N_2689,N_2872);
and UO_2 (O_2,N_2680,N_2942);
nand UO_3 (O_3,N_2849,N_2046);
and UO_4 (O_4,N_2793,N_2966);
or UO_5 (O_5,N_2246,N_2678);
or UO_6 (O_6,N_2317,N_2040);
nand UO_7 (O_7,N_2557,N_2479);
nor UO_8 (O_8,N_2665,N_2696);
nor UO_9 (O_9,N_2985,N_2164);
and UO_10 (O_10,N_2098,N_2178);
and UO_11 (O_11,N_2207,N_2537);
or UO_12 (O_12,N_2965,N_2387);
or UO_13 (O_13,N_2323,N_2854);
and UO_14 (O_14,N_2126,N_2371);
nand UO_15 (O_15,N_2429,N_2908);
or UO_16 (O_16,N_2605,N_2362);
and UO_17 (O_17,N_2023,N_2179);
or UO_18 (O_18,N_2891,N_2584);
and UO_19 (O_19,N_2386,N_2071);
nand UO_20 (O_20,N_2364,N_2654);
or UO_21 (O_21,N_2653,N_2233);
nor UO_22 (O_22,N_2290,N_2367);
and UO_23 (O_23,N_2080,N_2014);
nor UO_24 (O_24,N_2629,N_2964);
or UO_25 (O_25,N_2304,N_2572);
or UO_26 (O_26,N_2087,N_2644);
nand UO_27 (O_27,N_2796,N_2607);
nand UO_28 (O_28,N_2621,N_2863);
or UO_29 (O_29,N_2221,N_2694);
or UO_30 (O_30,N_2485,N_2769);
or UO_31 (O_31,N_2251,N_2292);
and UO_32 (O_32,N_2833,N_2216);
nand UO_33 (O_33,N_2556,N_2492);
and UO_34 (O_34,N_2036,N_2297);
and UO_35 (O_35,N_2512,N_2612);
nor UO_36 (O_36,N_2676,N_2899);
nor UO_37 (O_37,N_2748,N_2602);
or UO_38 (O_38,N_2747,N_2180);
or UO_39 (O_39,N_2016,N_2091);
or UO_40 (O_40,N_2493,N_2044);
nand UO_41 (O_41,N_2986,N_2523);
or UO_42 (O_42,N_2948,N_2397);
xor UO_43 (O_43,N_2874,N_2066);
and UO_44 (O_44,N_2093,N_2482);
or UO_45 (O_45,N_2941,N_2812);
or UO_46 (O_46,N_2618,N_2095);
and UO_47 (O_47,N_2967,N_2196);
nor UO_48 (O_48,N_2240,N_2341);
nand UO_49 (O_49,N_2634,N_2004);
nor UO_50 (O_50,N_2345,N_2003);
and UO_51 (O_51,N_2019,N_2760);
or UO_52 (O_52,N_2012,N_2610);
or UO_53 (O_53,N_2746,N_2472);
or UO_54 (O_54,N_2312,N_2218);
nand UO_55 (O_55,N_2960,N_2223);
or UO_56 (O_56,N_2477,N_2589);
or UO_57 (O_57,N_2754,N_2830);
and UO_58 (O_58,N_2474,N_2267);
xnor UO_59 (O_59,N_2068,N_2652);
and UO_60 (O_60,N_2463,N_2307);
nor UO_61 (O_61,N_2338,N_2327);
and UO_62 (O_62,N_2220,N_2745);
nand UO_63 (O_63,N_2279,N_2569);
and UO_64 (O_64,N_2790,N_2273);
nand UO_65 (O_65,N_2679,N_2766);
or UO_66 (O_66,N_2903,N_2757);
or UO_67 (O_67,N_2262,N_2383);
nor UO_68 (O_68,N_2856,N_2821);
nor UO_69 (O_69,N_2623,N_2291);
nor UO_70 (O_70,N_2910,N_2509);
or UO_71 (O_71,N_2843,N_2552);
or UO_72 (O_72,N_2845,N_2416);
nand UO_73 (O_73,N_2902,N_2263);
nor UO_74 (O_74,N_2088,N_2943);
nand UO_75 (O_75,N_2352,N_2256);
nor UO_76 (O_76,N_2033,N_2951);
nand UO_77 (O_77,N_2162,N_2441);
and UO_78 (O_78,N_2811,N_2320);
and UO_79 (O_79,N_2658,N_2593);
nor UO_80 (O_80,N_2912,N_2848);
and UO_81 (O_81,N_2978,N_2298);
and UO_82 (O_82,N_2002,N_2591);
nor UO_83 (O_83,N_2946,N_2513);
and UO_84 (O_84,N_2488,N_2968);
nor UO_85 (O_85,N_2466,N_2600);
or UO_86 (O_86,N_2663,N_2465);
nor UO_87 (O_87,N_2421,N_2773);
nor UO_88 (O_88,N_2732,N_2882);
or UO_89 (O_89,N_2542,N_2579);
nor UO_90 (O_90,N_2481,N_2794);
xnor UO_91 (O_91,N_2880,N_2245);
and UO_92 (O_92,N_2445,N_2299);
nand UO_93 (O_93,N_2423,N_2841);
or UO_94 (O_94,N_2063,N_2037);
and UO_95 (O_95,N_2737,N_2522);
nand UO_96 (O_96,N_2199,N_2138);
or UO_97 (O_97,N_2048,N_2917);
nor UO_98 (O_98,N_2081,N_2613);
and UO_99 (O_99,N_2209,N_2502);
nor UO_100 (O_100,N_2820,N_2375);
nand UO_101 (O_101,N_2639,N_2266);
or UO_102 (O_102,N_2759,N_2958);
nand UO_103 (O_103,N_2322,N_2484);
nor UO_104 (O_104,N_2301,N_2395);
or UO_105 (O_105,N_2527,N_2328);
and UO_106 (O_106,N_2982,N_2677);
and UO_107 (O_107,N_2483,N_2852);
nor UO_108 (O_108,N_2533,N_2420);
and UO_109 (O_109,N_2688,N_2624);
nand UO_110 (O_110,N_2107,N_2805);
nand UO_111 (O_111,N_2182,N_2718);
nor UO_112 (O_112,N_2619,N_2042);
or UO_113 (O_113,N_2189,N_2819);
nor UO_114 (O_114,N_2069,N_2907);
nor UO_115 (O_115,N_2120,N_2668);
nand UO_116 (O_116,N_2105,N_2149);
or UO_117 (O_117,N_2937,N_2271);
nand UO_118 (O_118,N_2708,N_2402);
nor UO_119 (O_119,N_2190,N_2456);
and UO_120 (O_120,N_2551,N_2562);
or UO_121 (O_121,N_2024,N_2581);
nand UO_122 (O_122,N_2406,N_2236);
nand UO_123 (O_123,N_2188,N_2661);
and UO_124 (O_124,N_2887,N_2800);
or UO_125 (O_125,N_2721,N_2728);
nor UO_126 (O_126,N_2075,N_2987);
nor UO_127 (O_127,N_2096,N_2727);
or UO_128 (O_128,N_2124,N_2510);
and UO_129 (O_129,N_2592,N_2158);
nor UO_130 (O_130,N_2735,N_2442);
nand UO_131 (O_131,N_2671,N_2803);
nor UO_132 (O_132,N_2807,N_2993);
nor UO_133 (O_133,N_2212,N_2278);
and UO_134 (O_134,N_2131,N_2909);
nor UO_135 (O_135,N_2580,N_2625);
and UO_136 (O_136,N_2544,N_2366);
or UO_137 (O_137,N_2167,N_2200);
or UO_138 (O_138,N_2077,N_2684);
and UO_139 (O_139,N_2422,N_2596);
nor UO_140 (O_140,N_2938,N_2775);
and UO_141 (O_141,N_2885,N_2136);
and UO_142 (O_142,N_2034,N_2026);
nand UO_143 (O_143,N_2761,N_2870);
nor UO_144 (O_144,N_2608,N_2940);
or UO_145 (O_145,N_2407,N_2869);
nor UO_146 (O_146,N_2376,N_2614);
nor UO_147 (O_147,N_2217,N_2576);
and UO_148 (O_148,N_2714,N_2999);
and UO_149 (O_149,N_2225,N_2115);
xnor UO_150 (O_150,N_2929,N_2249);
nor UO_151 (O_151,N_2662,N_2751);
and UO_152 (O_152,N_2097,N_2707);
nand UO_153 (O_153,N_2363,N_2815);
nand UO_154 (O_154,N_2112,N_2915);
nor UO_155 (O_155,N_2104,N_2187);
nor UO_156 (O_156,N_2140,N_2508);
or UO_157 (O_157,N_2117,N_2961);
nor UO_158 (O_158,N_2531,N_2191);
and UO_159 (O_159,N_2173,N_2720);
nand UO_160 (O_160,N_2637,N_2269);
or UO_161 (O_161,N_2393,N_2524);
nand UO_162 (O_162,N_2351,N_2532);
nor UO_163 (O_163,N_2275,N_2116);
nand UO_164 (O_164,N_2184,N_2823);
or UO_165 (O_165,N_2303,N_2308);
or UO_166 (O_166,N_2264,N_2094);
nand UO_167 (O_167,N_2950,N_2011);
and UO_168 (O_168,N_2148,N_2873);
nor UO_169 (O_169,N_2073,N_2704);
nor UO_170 (O_170,N_2563,N_2777);
and UO_171 (O_171,N_2875,N_2566);
nor UO_172 (O_172,N_2357,N_2074);
nand UO_173 (O_173,N_2930,N_2701);
nor UO_174 (O_174,N_2204,N_2391);
nor UO_175 (O_175,N_2226,N_2515);
nor UO_176 (O_176,N_2346,N_2467);
nor UO_177 (O_177,N_2260,N_2916);
nand UO_178 (O_178,N_2989,N_2729);
nand UO_179 (O_179,N_2529,N_2763);
xor UO_180 (O_180,N_2756,N_2744);
and UO_181 (O_181,N_2300,N_2213);
nor UO_182 (O_182,N_2868,N_2147);
or UO_183 (O_183,N_2065,N_2438);
or UO_184 (O_184,N_2851,N_2832);
nand UO_185 (O_185,N_2439,N_2770);
nor UO_186 (O_186,N_2546,N_2936);
nand UO_187 (O_187,N_2284,N_2996);
nand UO_188 (O_188,N_2924,N_2325);
and UO_189 (O_189,N_2876,N_2060);
nand UO_190 (O_190,N_2706,N_2137);
nor UO_191 (O_191,N_2287,N_2277);
nor UO_192 (O_192,N_2855,N_2038);
nor UO_193 (O_193,N_2548,N_2434);
nor UO_194 (O_194,N_2932,N_2448);
xor UO_195 (O_195,N_2501,N_2401);
nor UO_196 (O_196,N_2957,N_2558);
and UO_197 (O_197,N_2813,N_2555);
and UO_198 (O_198,N_2344,N_2716);
nand UO_199 (O_199,N_2450,N_2898);
or UO_200 (O_200,N_2920,N_2151);
nor UO_201 (O_201,N_2051,N_2831);
or UO_202 (O_202,N_2687,N_2155);
nor UO_203 (O_203,N_2324,N_2514);
nand UO_204 (O_204,N_2035,N_2645);
nand UO_205 (O_205,N_2500,N_2005);
xnor UO_206 (O_206,N_2041,N_2031);
or UO_207 (O_207,N_2417,N_2414);
xnor UO_208 (O_208,N_2254,N_2913);
and UO_209 (O_209,N_2486,N_2877);
or UO_210 (O_210,N_2468,N_2983);
or UO_211 (O_211,N_2517,N_2437);
or UO_212 (O_212,N_2403,N_2333);
and UO_213 (O_213,N_2926,N_2723);
nand UO_214 (O_214,N_2090,N_2296);
nor UO_215 (O_215,N_2740,N_2838);
and UO_216 (O_216,N_2586,N_2853);
or UO_217 (O_217,N_2419,N_2894);
nor UO_218 (O_218,N_2839,N_2409);
nand UO_219 (O_219,N_2358,N_2230);
nor UO_220 (O_220,N_2146,N_2521);
nand UO_221 (O_221,N_2862,N_2944);
nor UO_222 (O_222,N_2846,N_2519);
nor UO_223 (O_223,N_2997,N_2578);
nand UO_224 (O_224,N_2998,N_2145);
nand UO_225 (O_225,N_2836,N_2243);
nand UO_226 (O_226,N_2879,N_2971);
or UO_227 (O_227,N_2353,N_2415);
nor UO_228 (O_228,N_2110,N_2504);
nor UO_229 (O_229,N_2478,N_2092);
or UO_230 (O_230,N_2451,N_2847);
xnor UO_231 (O_231,N_2651,N_2128);
and UO_232 (O_232,N_2626,N_2959);
nor UO_233 (O_233,N_2118,N_2489);
nand UO_234 (O_234,N_2130,N_2791);
and UO_235 (O_235,N_2731,N_2144);
nand UO_236 (O_236,N_2281,N_2274);
and UO_237 (O_237,N_2412,N_2253);
nor UO_238 (O_238,N_2972,N_2354);
or UO_239 (O_239,N_2588,N_2310);
or UO_240 (O_240,N_2632,N_2878);
nor UO_241 (O_241,N_2963,N_2949);
and UO_242 (O_242,N_2647,N_2309);
nand UO_243 (O_243,N_2161,N_2881);
and UO_244 (O_244,N_2449,N_2683);
nand UO_245 (O_245,N_2890,N_2669);
xnor UO_246 (O_246,N_2954,N_2778);
and UO_247 (O_247,N_2106,N_2224);
nor UO_248 (O_248,N_2174,N_2435);
and UO_249 (O_249,N_2067,N_2459);
nor UO_250 (O_250,N_2049,N_2641);
and UO_251 (O_251,N_2139,N_2636);
or UO_252 (O_252,N_2767,N_2827);
or UO_253 (O_253,N_2886,N_2228);
nor UO_254 (O_254,N_2413,N_2674);
or UO_255 (O_255,N_2611,N_2313);
xor UO_256 (O_256,N_2302,N_2675);
nor UO_257 (O_257,N_2541,N_2165);
or UO_258 (O_258,N_2686,N_2446);
xor UO_259 (O_259,N_2134,N_2261);
nor UO_260 (O_260,N_2460,N_2705);
or UO_261 (O_261,N_2692,N_2762);
and UO_262 (O_262,N_2257,N_2765);
nor UO_263 (O_263,N_2782,N_2270);
nor UO_264 (O_264,N_2595,N_2994);
nor UO_265 (O_265,N_2540,N_2440);
or UO_266 (O_266,N_2742,N_2461);
or UO_267 (O_267,N_2750,N_2001);
or UO_268 (O_268,N_2657,N_2201);
or UO_269 (O_269,N_2113,N_2008);
xnor UO_270 (O_270,N_2724,N_2427);
nand UO_271 (O_271,N_2499,N_2824);
nand UO_272 (O_272,N_2753,N_2861);
and UO_273 (O_273,N_2168,N_2054);
nor UO_274 (O_274,N_2781,N_2939);
or UO_275 (O_275,N_2089,N_2469);
xor UO_276 (O_276,N_2785,N_2709);
nor UO_277 (O_277,N_2258,N_2470);
and UO_278 (O_278,N_2804,N_2047);
and UO_279 (O_279,N_2638,N_2617);
xor UO_280 (O_280,N_2057,N_2342);
nor UO_281 (O_281,N_2385,N_2028);
or UO_282 (O_282,N_2573,N_2177);
and UO_283 (O_283,N_2866,N_2480);
nor UO_284 (O_284,N_2006,N_2561);
nor UO_285 (O_285,N_2123,N_2802);
or UO_286 (O_286,N_2536,N_2698);
nand UO_287 (O_287,N_2356,N_2176);
nand UO_288 (O_288,N_2247,N_2945);
nor UO_289 (O_289,N_2897,N_2396);
or UO_290 (O_290,N_2293,N_2809);
or UO_291 (O_291,N_2382,N_2655);
nand UO_292 (O_292,N_2072,N_2976);
and UO_293 (O_293,N_2101,N_2547);
nor UO_294 (O_294,N_2305,N_2506);
or UO_295 (O_295,N_2494,N_2394);
or UO_296 (O_296,N_2222,N_2574);
and UO_297 (O_297,N_2717,N_2326);
nand UO_298 (O_298,N_2980,N_2122);
nand UO_299 (O_299,N_2330,N_2628);
nand UO_300 (O_300,N_2359,N_2922);
xor UO_301 (O_301,N_2534,N_2865);
or UO_302 (O_302,N_2447,N_2988);
nor UO_303 (O_303,N_2205,N_2336);
nand UO_304 (O_304,N_2681,N_2430);
nand UO_305 (O_305,N_2818,N_2009);
nor UO_306 (O_306,N_2210,N_2490);
or UO_307 (O_307,N_2214,N_2825);
xnor UO_308 (O_308,N_2864,N_2424);
or UO_309 (O_309,N_2433,N_2810);
and UO_310 (O_310,N_2082,N_2571);
nand UO_311 (O_311,N_2369,N_2377);
nor UO_312 (O_312,N_2892,N_2788);
nor UO_313 (O_313,N_2389,N_2952);
or UO_314 (O_314,N_2343,N_2025);
nor UO_315 (O_315,N_2193,N_2398);
and UO_316 (O_316,N_2232,N_2921);
or UO_317 (O_317,N_2829,N_2237);
nand UO_318 (O_318,N_2432,N_2064);
nand UO_319 (O_319,N_2736,N_2857);
and UO_320 (O_320,N_2858,N_2153);
nor UO_321 (O_321,N_2664,N_2039);
and UO_322 (O_322,N_2934,N_2911);
nand UO_323 (O_323,N_2660,N_2186);
nor UO_324 (O_324,N_2392,N_2814);
or UO_325 (O_325,N_2643,N_2102);
nor UO_326 (O_326,N_2587,N_2013);
nand UO_327 (O_327,N_2550,N_2565);
nand UO_328 (O_328,N_2022,N_2384);
nor UO_329 (O_329,N_2062,N_2076);
nor UO_330 (O_330,N_2764,N_2518);
nand UO_331 (O_331,N_2603,N_2283);
nor UO_332 (O_332,N_2808,N_2319);
or UO_333 (O_333,N_2443,N_2953);
xnor UO_334 (O_334,N_2919,N_2801);
and UO_335 (O_335,N_2666,N_2169);
nand UO_336 (O_336,N_2285,N_2295);
or UO_337 (O_337,N_2594,N_2462);
nor UO_338 (O_338,N_2935,N_2321);
or UO_339 (O_339,N_2871,N_2280);
and UO_340 (O_340,N_2837,N_2722);
nor UO_341 (O_341,N_2516,N_2776);
or UO_342 (O_342,N_2719,N_2198);
and UO_343 (O_343,N_2373,N_2826);
nand UO_344 (O_344,N_2365,N_2497);
or UO_345 (O_345,N_2288,N_2984);
nand UO_346 (O_346,N_2559,N_2337);
and UO_347 (O_347,N_2901,N_2306);
nor UO_348 (O_348,N_2368,N_2252);
or UO_349 (O_349,N_2318,N_2609);
or UO_350 (O_350,N_2635,N_2203);
or UO_351 (O_351,N_2156,N_2525);
and UO_352 (O_352,N_2713,N_2132);
and UO_353 (O_353,N_2646,N_2585);
nand UO_354 (O_354,N_2143,N_2693);
and UO_355 (O_355,N_2248,N_2454);
and UO_356 (O_356,N_2192,N_2741);
nand UO_357 (O_357,N_2969,N_2789);
or UO_358 (O_358,N_2234,N_2834);
nor UO_359 (O_359,N_2487,N_2331);
and UO_360 (O_360,N_2992,N_2734);
or UO_361 (O_361,N_2627,N_2553);
and UO_362 (O_362,N_2111,N_2170);
and UO_363 (O_363,N_2242,N_2206);
nor UO_364 (O_364,N_2015,N_2411);
and UO_365 (O_365,N_2642,N_2171);
or UO_366 (O_366,N_2361,N_2163);
and UO_367 (O_367,N_2505,N_2400);
nor UO_368 (O_368,N_2334,N_2202);
nor UO_369 (O_369,N_2241,N_2844);
nor UO_370 (O_370,N_2567,N_2582);
and UO_371 (O_371,N_2452,N_2606);
or UO_372 (O_372,N_2577,N_2520);
and UO_373 (O_373,N_2154,N_2730);
nor UO_374 (O_374,N_2768,N_2900);
or UO_375 (O_375,N_2604,N_2332);
nor UO_376 (O_376,N_2884,N_2700);
nor UO_377 (O_377,N_2141,N_2955);
or UO_378 (O_378,N_2119,N_2100);
nand UO_379 (O_379,N_2255,N_2656);
or UO_380 (O_380,N_2195,N_2029);
and UO_381 (O_381,N_2918,N_2215);
or UO_382 (O_382,N_2906,N_2990);
and UO_383 (O_383,N_2355,N_2828);
nand UO_384 (O_384,N_2822,N_2597);
and UO_385 (O_385,N_2455,N_2043);
and UO_386 (O_386,N_2099,N_2282);
nor UO_387 (O_387,N_2947,N_2329);
and UO_388 (O_388,N_2129,N_2208);
nand UO_389 (O_389,N_2360,N_2311);
and UO_390 (O_390,N_2272,N_2560);
or UO_391 (O_391,N_2491,N_2335);
nor UO_392 (O_392,N_2030,N_2712);
and UO_393 (O_393,N_2859,N_2710);
nand UO_394 (O_394,N_2150,N_2053);
nor UO_395 (O_395,N_2045,N_2250);
nand UO_396 (O_396,N_2640,N_2289);
or UO_397 (O_397,N_2511,N_2227);
or UO_398 (O_398,N_2599,N_2752);
nand UO_399 (O_399,N_2549,N_2058);
nor UO_400 (O_400,N_2539,N_2055);
nor UO_401 (O_401,N_2374,N_2780);
or UO_402 (O_402,N_2166,N_2904);
nor UO_403 (O_403,N_2498,N_2888);
or UO_404 (O_404,N_2121,N_2670);
nand UO_405 (O_405,N_2503,N_2349);
nand UO_406 (O_406,N_2598,N_2316);
nand UO_407 (O_407,N_2715,N_2183);
nand UO_408 (O_408,N_2061,N_2779);
and UO_409 (O_409,N_2127,N_2133);
nand UO_410 (O_410,N_2738,N_2370);
or UO_411 (O_411,N_2850,N_2530);
or UO_412 (O_412,N_2194,N_2294);
or UO_413 (O_413,N_2995,N_2755);
and UO_414 (O_414,N_2889,N_2795);
nor UO_415 (O_415,N_2649,N_2453);
nand UO_416 (O_416,N_2239,N_2883);
xnor UO_417 (O_417,N_2797,N_2032);
nor UO_418 (O_418,N_2973,N_2977);
or UO_419 (O_419,N_2380,N_2235);
or UO_420 (O_420,N_2339,N_2159);
or UO_421 (O_421,N_2372,N_2895);
nand UO_422 (O_422,N_2348,N_2925);
or UO_423 (O_423,N_2786,N_2601);
nor UO_424 (O_424,N_2615,N_2835);
nand UO_425 (O_425,N_2806,N_2000);
nor UO_426 (O_426,N_2458,N_2020);
and UO_427 (O_427,N_2630,N_2388);
and UO_428 (O_428,N_2404,N_2495);
or UO_429 (O_429,N_2981,N_2379);
nand UO_430 (O_430,N_2018,N_2390);
nor UO_431 (O_431,N_2428,N_2535);
and UO_432 (O_432,N_2905,N_2086);
xnor UO_433 (O_433,N_2431,N_2059);
nand UO_434 (O_434,N_2564,N_2538);
nor UO_435 (O_435,N_2787,N_2575);
or UO_436 (O_436,N_2157,N_2314);
and UO_437 (O_437,N_2238,N_2114);
or UO_438 (O_438,N_2211,N_2979);
and UO_439 (O_439,N_2476,N_2410);
or UO_440 (O_440,N_2528,N_2083);
and UO_441 (O_441,N_2816,N_2007);
or UO_442 (O_442,N_2231,N_2052);
or UO_443 (O_443,N_2672,N_2931);
nor UO_444 (O_444,N_2711,N_2928);
nand UO_445 (O_445,N_2444,N_2633);
or UO_446 (O_446,N_2347,N_2673);
and UO_447 (O_447,N_2350,N_2197);
or UO_448 (O_448,N_2695,N_2970);
and UO_449 (O_449,N_2991,N_2840);
xor UO_450 (O_450,N_2648,N_2017);
nor UO_451 (O_451,N_2962,N_2554);
or UO_452 (O_452,N_2070,N_2733);
or UO_453 (O_453,N_2697,N_2315);
or UO_454 (O_454,N_2078,N_2774);
nand UO_455 (O_455,N_2125,N_2771);
nand UO_456 (O_456,N_2244,N_2726);
and UO_457 (O_457,N_2842,N_2142);
nand UO_458 (O_458,N_2135,N_2473);
and UO_459 (O_459,N_2923,N_2739);
or UO_460 (O_460,N_2340,N_2725);
or UO_461 (O_461,N_2583,N_2974);
nand UO_462 (O_462,N_2405,N_2425);
or UO_463 (O_463,N_2914,N_2027);
xor UO_464 (O_464,N_2172,N_2175);
and UO_465 (O_465,N_2743,N_2010);
nor UO_466 (O_466,N_2956,N_2276);
xor UO_467 (O_467,N_2543,N_2084);
or UO_468 (O_468,N_2860,N_2021);
nand UO_469 (O_469,N_2160,N_2867);
nand UO_470 (O_470,N_2772,N_2185);
nor UO_471 (O_471,N_2817,N_2545);
and UO_472 (O_472,N_2702,N_2229);
xor UO_473 (O_473,N_2109,N_2457);
nor UO_474 (O_474,N_2056,N_2933);
or UO_475 (O_475,N_2268,N_2590);
nor UO_476 (O_476,N_2181,N_2631);
nor UO_477 (O_477,N_2616,N_2703);
nand UO_478 (O_478,N_2418,N_2378);
nor UO_479 (O_479,N_2103,N_2570);
and UO_480 (O_480,N_2471,N_2399);
and UO_481 (O_481,N_2152,N_2622);
and UO_482 (O_482,N_2682,N_2219);
or UO_483 (O_483,N_2286,N_2975);
and UO_484 (O_484,N_2691,N_2799);
or UO_485 (O_485,N_2659,N_2699);
nor UO_486 (O_486,N_2408,N_2381);
nor UO_487 (O_487,N_2526,N_2792);
and UO_488 (O_488,N_2108,N_2667);
or UO_489 (O_489,N_2464,N_2690);
nand UO_490 (O_490,N_2784,N_2507);
or UO_491 (O_491,N_2079,N_2475);
nor UO_492 (O_492,N_2798,N_2265);
nor UO_493 (O_493,N_2749,N_2085);
nor UO_494 (O_494,N_2620,N_2050);
or UO_495 (O_495,N_2896,N_2259);
or UO_496 (O_496,N_2783,N_2927);
nor UO_497 (O_497,N_2568,N_2426);
or UO_498 (O_498,N_2758,N_2650);
nand UO_499 (O_499,N_2436,N_2496);
endmodule