module basic_1500_15000_2000_10_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_1360,In_210);
nor U1 (N_1,In_1445,In_8);
or U2 (N_2,In_1218,In_755);
and U3 (N_3,In_179,In_1439);
nand U4 (N_4,In_1011,In_578);
nand U5 (N_5,In_1462,In_1494);
or U6 (N_6,In_165,In_1029);
or U7 (N_7,In_24,In_777);
nand U8 (N_8,In_698,In_899);
or U9 (N_9,In_1413,In_1231);
nand U10 (N_10,In_1422,In_617);
or U11 (N_11,In_923,In_985);
nor U12 (N_12,In_236,In_776);
xor U13 (N_13,In_61,In_237);
or U14 (N_14,In_412,In_1266);
or U15 (N_15,In_444,In_569);
and U16 (N_16,In_255,In_340);
nand U17 (N_17,In_957,In_1428);
nor U18 (N_18,In_737,In_97);
and U19 (N_19,In_726,In_290);
and U20 (N_20,In_835,In_645);
and U21 (N_21,In_298,In_954);
nor U22 (N_22,In_1290,In_1032);
or U23 (N_23,In_1034,In_631);
nand U24 (N_24,In_608,In_309);
xor U25 (N_25,In_79,In_1442);
or U26 (N_26,In_392,In_459);
xnor U27 (N_27,In_361,In_1305);
nor U28 (N_28,In_1424,In_612);
nor U29 (N_29,In_518,In_157);
nand U30 (N_30,In_1448,In_671);
nor U31 (N_31,In_979,In_1315);
nor U32 (N_32,In_377,In_821);
xnor U33 (N_33,In_370,In_1133);
and U34 (N_34,In_1477,In_843);
nand U35 (N_35,In_1320,In_874);
or U36 (N_36,In_545,In_1410);
xor U37 (N_37,In_1354,In_249);
nand U38 (N_38,In_485,In_567);
or U39 (N_39,In_50,In_222);
or U40 (N_40,In_568,In_891);
and U41 (N_41,In_1093,In_683);
or U42 (N_42,In_268,In_342);
nor U43 (N_43,In_1080,In_120);
nand U44 (N_44,In_173,In_563);
nor U45 (N_45,In_64,In_10);
and U46 (N_46,In_478,In_918);
nor U47 (N_47,In_1425,In_1040);
nand U48 (N_48,In_1476,In_1015);
xor U49 (N_49,In_376,In_372);
nor U50 (N_50,In_474,In_1308);
nand U51 (N_51,In_435,In_572);
nor U52 (N_52,In_928,In_615);
xor U53 (N_53,In_994,In_1267);
or U54 (N_54,In_1342,In_765);
and U55 (N_55,In_502,In_29);
nor U56 (N_56,In_1466,In_384);
and U57 (N_57,In_195,In_1152);
and U58 (N_58,In_281,In_774);
and U59 (N_59,In_834,In_215);
and U60 (N_60,In_1475,In_916);
nand U61 (N_61,In_481,In_152);
nor U62 (N_62,In_1082,In_225);
xnor U63 (N_63,In_1291,In_1028);
xor U64 (N_64,In_25,In_678);
and U65 (N_65,In_820,In_845);
xnor U66 (N_66,In_1274,In_497);
xor U67 (N_67,In_1008,In_1057);
nand U68 (N_68,In_118,In_814);
and U69 (N_69,In_308,In_987);
and U70 (N_70,In_1160,In_334);
and U71 (N_71,In_993,In_144);
nor U72 (N_72,In_410,In_1101);
or U73 (N_73,In_27,In_419);
nand U74 (N_74,In_1024,In_1416);
or U75 (N_75,In_798,In_443);
or U76 (N_76,In_712,In_905);
nand U77 (N_77,In_1210,In_694);
and U78 (N_78,In_790,In_1349);
xnor U79 (N_79,In_635,In_988);
and U80 (N_80,In_402,In_510);
or U81 (N_81,In_584,In_1199);
nor U82 (N_82,In_1255,In_853);
and U83 (N_83,In_270,In_368);
nor U84 (N_84,In_1429,In_894);
nand U85 (N_85,In_1285,In_764);
xnor U86 (N_86,In_445,In_101);
nand U87 (N_87,In_109,In_493);
or U88 (N_88,In_278,In_1155);
nor U89 (N_89,In_672,In_1336);
nor U90 (N_90,In_1184,In_1200);
xnor U91 (N_91,In_785,In_605);
xor U92 (N_92,In_437,In_411);
or U93 (N_93,In_525,In_1170);
nor U94 (N_94,In_665,In_257);
and U95 (N_95,In_1117,In_876);
and U96 (N_96,In_926,In_330);
and U97 (N_97,In_625,In_452);
xor U98 (N_98,In_286,In_86);
nand U99 (N_99,In_138,In_746);
nor U100 (N_100,In_1495,In_751);
and U101 (N_101,In_1118,In_620);
or U102 (N_102,In_646,In_576);
nand U103 (N_103,In_956,In_513);
nand U104 (N_104,In_1077,In_1149);
nor U105 (N_105,In_921,In_939);
nand U106 (N_106,In_111,In_495);
xor U107 (N_107,In_610,In_316);
and U108 (N_108,In_1414,In_1379);
or U109 (N_109,In_253,In_784);
nand U110 (N_110,In_1099,In_841);
nand U111 (N_111,In_149,In_583);
nor U112 (N_112,In_971,In_1039);
xnor U113 (N_113,In_69,In_1176);
nor U114 (N_114,In_1491,In_935);
nand U115 (N_115,In_686,In_33);
nand U116 (N_116,In_87,In_7);
nor U117 (N_117,In_1018,In_489);
or U118 (N_118,In_1196,In_1130);
nand U119 (N_119,In_828,In_103);
nand U120 (N_120,In_358,In_122);
nor U121 (N_121,In_657,In_1168);
xor U122 (N_122,In_1249,In_1206);
xor U123 (N_123,In_366,In_1020);
and U124 (N_124,In_1346,In_1131);
and U125 (N_125,In_648,In_1352);
or U126 (N_126,In_830,In_753);
xor U127 (N_127,In_702,In_1321);
nand U128 (N_128,In_732,In_554);
and U129 (N_129,In_1447,In_1453);
nor U130 (N_130,In_446,In_807);
nor U131 (N_131,In_775,In_388);
and U132 (N_132,In_1405,In_1229);
or U133 (N_133,In_362,In_571);
and U134 (N_134,In_184,In_863);
or U135 (N_135,In_1232,In_623);
nand U136 (N_136,In_1294,In_1211);
xor U137 (N_137,In_997,In_663);
xnor U138 (N_138,In_603,In_1132);
nand U139 (N_139,In_983,In_151);
or U140 (N_140,In_284,In_1022);
nand U141 (N_141,In_662,In_669);
nand U142 (N_142,In_818,In_48);
or U143 (N_143,In_1469,In_805);
and U144 (N_144,In_1393,In_1460);
xnor U145 (N_145,In_295,In_1191);
nand U146 (N_146,In_390,In_674);
xor U147 (N_147,In_604,In_889);
nand U148 (N_148,In_1060,In_104);
nor U149 (N_149,In_692,In_326);
or U150 (N_150,In_279,In_1182);
or U151 (N_151,In_1141,In_541);
and U152 (N_152,In_873,In_57);
or U153 (N_153,In_815,In_654);
or U154 (N_154,In_1279,In_310);
xor U155 (N_155,In_929,In_1483);
nor U156 (N_156,In_1383,In_629);
nor U157 (N_157,In_1450,In_901);
nor U158 (N_158,In_320,In_416);
nand U159 (N_159,In_154,In_323);
nor U160 (N_160,In_1202,In_1044);
xor U161 (N_161,In_356,In_1430);
xor U162 (N_162,In_1106,In_1071);
nor U163 (N_163,In_58,In_1356);
nor U164 (N_164,In_233,In_288);
or U165 (N_165,In_634,In_307);
and U166 (N_166,In_909,In_667);
or U167 (N_167,In_1151,In_429);
nand U168 (N_168,In_846,In_303);
and U169 (N_169,In_175,In_243);
nand U170 (N_170,In_950,In_1037);
and U171 (N_171,In_967,In_114);
nand U172 (N_172,In_90,In_272);
nor U173 (N_173,In_218,In_575);
nor U174 (N_174,In_738,In_117);
or U175 (N_175,In_728,In_1479);
nor U176 (N_176,In_884,In_81);
xor U177 (N_177,In_1474,In_407);
and U178 (N_178,In_581,In_482);
and U179 (N_179,In_761,In_214);
nor U180 (N_180,In_201,In_209);
xnor U181 (N_181,In_670,In_886);
xor U182 (N_182,In_464,In_391);
nor U183 (N_183,In_174,In_978);
xor U184 (N_184,In_325,In_773);
nor U185 (N_185,In_78,In_1197);
nor U186 (N_186,In_1454,In_1105);
xor U187 (N_187,In_508,In_1209);
and U188 (N_188,In_460,In_1282);
nor U189 (N_189,In_359,In_962);
or U190 (N_190,In_596,In_1396);
xnor U191 (N_191,In_658,In_529);
and U192 (N_192,In_1104,In_1338);
and U193 (N_193,In_1110,In_23);
nand U194 (N_194,In_992,In_748);
nand U195 (N_195,In_1280,In_386);
or U196 (N_196,In_703,In_46);
or U197 (N_197,In_1314,In_223);
xnor U198 (N_198,In_706,In_801);
nand U199 (N_199,In_216,In_153);
and U200 (N_200,In_852,In_877);
and U201 (N_201,In_251,In_20);
and U202 (N_202,In_491,In_102);
nand U203 (N_203,In_839,In_500);
nor U204 (N_204,In_26,In_135);
nand U205 (N_205,In_695,In_1481);
xor U206 (N_206,In_1156,In_709);
and U207 (N_207,In_1053,In_1056);
and U208 (N_208,In_1030,In_966);
or U209 (N_209,In_528,In_100);
or U210 (N_210,In_844,In_74);
nor U211 (N_211,In_1035,In_1108);
or U212 (N_212,In_1221,In_55);
and U213 (N_213,In_952,In_403);
and U214 (N_214,In_352,In_848);
or U215 (N_215,In_1389,In_1194);
nand U216 (N_216,In_531,In_463);
nand U217 (N_217,In_301,In_287);
and U218 (N_218,In_1323,In_364);
xor U219 (N_219,In_1400,In_250);
nor U220 (N_220,In_62,In_129);
or U221 (N_221,In_126,In_855);
and U222 (N_222,In_395,In_15);
and U223 (N_223,In_389,In_1432);
or U224 (N_224,In_740,In_1254);
nor U225 (N_225,In_782,In_958);
nor U226 (N_226,In_1162,In_1251);
and U227 (N_227,In_1302,In_82);
xnor U228 (N_228,In_548,In_742);
xor U229 (N_229,In_42,In_351);
nand U230 (N_230,In_1113,In_516);
xor U231 (N_231,In_507,In_275);
nand U232 (N_232,In_299,In_1041);
nor U233 (N_233,In_856,In_816);
or U234 (N_234,In_1187,In_809);
nand U235 (N_235,In_1148,In_727);
nor U236 (N_236,In_394,In_1487);
or U237 (N_237,In_494,In_1441);
and U238 (N_238,In_186,In_919);
xor U239 (N_239,In_1178,In_903);
xnor U240 (N_240,In_867,In_858);
xnor U241 (N_241,In_882,In_294);
xnor U242 (N_242,In_552,In_473);
and U243 (N_243,In_944,In_1373);
nand U244 (N_244,In_110,In_1241);
and U245 (N_245,In_312,In_1247);
nand U246 (N_246,In_514,In_1050);
and U247 (N_247,In_344,In_557);
and U248 (N_248,In_115,In_859);
nand U249 (N_249,In_1214,In_872);
xor U250 (N_250,In_1079,In_1137);
xor U251 (N_251,In_1066,In_611);
and U252 (N_252,In_527,In_199);
or U253 (N_253,In_191,In_976);
nand U254 (N_254,In_833,In_734);
nand U255 (N_255,In_1407,In_724);
nor U256 (N_256,In_185,In_558);
and U257 (N_257,In_1169,In_171);
and U258 (N_258,In_1318,In_1253);
and U259 (N_259,In_319,In_1122);
and U260 (N_260,In_397,In_458);
or U261 (N_261,In_550,In_613);
and U262 (N_262,In_1175,In_787);
nand U263 (N_263,In_1458,In_434);
nor U264 (N_264,In_984,In_649);
nand U265 (N_265,In_953,In_547);
nand U266 (N_266,In_1100,In_314);
nand U267 (N_267,In_83,In_32);
and U268 (N_268,In_1240,In_1488);
xnor U269 (N_269,In_1293,In_68);
or U270 (N_270,In_506,In_14);
or U271 (N_271,In_424,In_825);
xor U272 (N_272,In_520,In_769);
and U273 (N_273,In_586,In_1142);
nand U274 (N_274,In_1419,In_1343);
and U275 (N_275,In_744,In_684);
and U276 (N_276,In_895,In_139);
or U277 (N_277,In_826,In_333);
and U278 (N_278,In_213,In_1451);
nor U279 (N_279,In_1239,In_1486);
nand U280 (N_280,In_163,In_947);
or U281 (N_281,In_108,In_515);
xor U282 (N_282,In_675,In_41);
nor U283 (N_283,In_864,In_169);
and U284 (N_284,In_1192,In_143);
nand U285 (N_285,In_731,In_338);
and U286 (N_286,In_924,In_131);
nor U287 (N_287,In_1406,In_938);
and U288 (N_288,In_866,In_313);
xnor U289 (N_289,In_965,In_758);
or U290 (N_290,In_354,In_564);
or U291 (N_291,In_1382,In_1378);
and U292 (N_292,In_1374,In_1193);
nor U293 (N_293,In_1042,In_1046);
and U294 (N_294,In_1140,In_99);
nand U295 (N_295,In_94,In_677);
nand U296 (N_296,In_1112,In_741);
nor U297 (N_297,In_503,In_1499);
nand U298 (N_298,In_1456,In_246);
xor U299 (N_299,In_1361,In_133);
or U300 (N_300,In_360,In_1310);
xnor U301 (N_301,In_960,In_730);
or U302 (N_302,In_733,In_206);
nand U303 (N_303,In_704,In_1125);
or U304 (N_304,In_1337,In_804);
nor U305 (N_305,In_399,In_1370);
xnor U306 (N_306,In_974,In_1123);
and U307 (N_307,In_297,In_1440);
or U308 (N_308,In_824,In_881);
nand U309 (N_309,In_1036,In_140);
nor U310 (N_310,In_1283,In_451);
nor U311 (N_311,In_925,In_1468);
and U312 (N_312,In_418,In_207);
or U313 (N_313,In_1333,In_986);
and U314 (N_314,In_739,In_1412);
or U315 (N_315,In_779,In_888);
nor U316 (N_316,In_602,In_931);
xnor U317 (N_317,In_745,In_119);
nor U318 (N_318,In_311,In_262);
nand U319 (N_319,In_38,In_1078);
and U320 (N_320,In_523,In_1086);
and U321 (N_321,In_549,In_1183);
xnor U322 (N_322,In_1388,In_972);
xnor U323 (N_323,In_400,In_1497);
and U324 (N_324,In_1095,In_1208);
or U325 (N_325,In_865,In_291);
nand U326 (N_326,In_431,In_778);
or U327 (N_327,In_1212,In_722);
nor U328 (N_328,In_375,In_1173);
and U329 (N_329,In_9,In_639);
nor U330 (N_330,In_736,In_1449);
nand U331 (N_331,In_831,In_1284);
or U332 (N_332,In_229,In_1220);
or U333 (N_333,In_851,In_1401);
nor U334 (N_334,In_1059,In_760);
and U335 (N_335,In_1390,In_910);
or U336 (N_336,In_943,In_1074);
nand U337 (N_337,In_1496,In_107);
and U338 (N_338,In_720,In_806);
or U339 (N_339,In_1455,In_1147);
or U340 (N_340,In_168,In_341);
nand U341 (N_341,In_1097,In_1482);
xor U342 (N_342,In_105,In_182);
and U343 (N_343,In_651,In_1195);
nand U344 (N_344,In_1045,In_1435);
nand U345 (N_345,In_1426,In_193);
xnor U346 (N_346,In_1329,In_1129);
and U347 (N_347,In_355,In_1230);
nor U348 (N_348,In_1054,In_476);
and U349 (N_349,In_254,In_1252);
and U350 (N_350,In_1167,In_633);
xor U351 (N_351,In_1335,In_1242);
nand U352 (N_352,In_421,In_150);
and U353 (N_353,In_1437,In_296);
nand U354 (N_354,In_430,In_606);
xor U355 (N_355,In_43,In_932);
and U356 (N_356,In_879,In_212);
xnor U357 (N_357,In_791,In_475);
and U358 (N_358,In_227,In_945);
or U359 (N_359,In_335,In_77);
nand U360 (N_360,In_1480,In_1092);
or U361 (N_361,In_1418,In_1399);
xnor U362 (N_362,In_381,In_252);
nor U363 (N_363,In_98,In_630);
nor U364 (N_364,In_158,In_1325);
or U365 (N_365,In_1087,In_1157);
or U366 (N_366,In_729,In_276);
xnor U367 (N_367,In_4,In_1340);
xnor U368 (N_368,In_735,In_1052);
and U369 (N_369,In_220,In_1296);
or U370 (N_370,In_378,In_1359);
or U371 (N_371,In_180,In_699);
or U372 (N_372,In_754,In_123);
or U373 (N_373,In_1309,In_1444);
or U374 (N_374,In_1292,In_897);
nand U375 (N_375,In_1180,In_1019);
and U376 (N_376,In_537,In_1331);
nor U377 (N_377,In_1065,In_1004);
nand U378 (N_378,In_318,In_367);
or U379 (N_379,In_1070,In_1295);
nor U380 (N_380,In_1012,In_369);
or U381 (N_381,In_1213,In_1072);
nor U382 (N_382,In_887,In_264);
nand U383 (N_383,In_1402,In_680);
xnor U384 (N_384,In_991,In_1411);
xnor U385 (N_385,In_1471,In_788);
xor U386 (N_386,In_1225,In_382);
nor U387 (N_387,In_1243,In_585);
nor U388 (N_388,In_1286,In_221);
nor U389 (N_389,In_92,In_1386);
nand U390 (N_390,In_1387,In_1261);
xor U391 (N_391,In_1367,In_22);
nand U392 (N_392,In_89,In_679);
nand U393 (N_393,In_468,In_142);
and U394 (N_394,In_690,In_591);
nand U395 (N_395,In_668,In_203);
or U396 (N_396,In_810,In_1268);
and U397 (N_397,In_1236,In_462);
or U398 (N_398,In_5,In_1281);
nor U399 (N_399,In_1043,In_650);
nor U400 (N_400,In_426,In_836);
nand U401 (N_401,In_1385,In_1189);
xor U402 (N_402,In_878,In_1174);
and U403 (N_403,In_1490,In_717);
nor U404 (N_404,In_365,In_802);
nand U405 (N_405,In_1278,In_900);
nor U406 (N_406,In_1403,In_1300);
nand U407 (N_407,In_53,In_556);
nor U408 (N_408,In_172,In_159);
or U409 (N_409,In_1366,In_659);
or U410 (N_410,In_544,In_756);
or U411 (N_411,In_1250,In_39);
nor U412 (N_412,In_161,In_408);
xnor U413 (N_413,In_273,In_934);
nor U414 (N_414,In_1237,In_1391);
xnor U415 (N_415,In_534,In_19);
xnor U416 (N_416,In_1459,In_134);
and U417 (N_417,In_1047,In_282);
or U418 (N_418,In_155,In_618);
and U419 (N_419,In_1235,In_656);
xnor U420 (N_420,In_1478,In_817);
or U421 (N_421,In_823,In_31);
nor U422 (N_422,In_304,In_854);
and U423 (N_423,In_1364,In_1446);
xnor U424 (N_424,In_619,In_1145);
nand U425 (N_425,In_84,In_1215);
xor U426 (N_426,In_65,In_160);
nand U427 (N_427,In_850,In_234);
nor U428 (N_428,In_1381,In_1107);
nand U429 (N_429,In_1316,In_721);
nor U430 (N_430,In_1404,In_1324);
nand U431 (N_431,In_181,In_1114);
nor U432 (N_432,In_827,In_1326);
nor U433 (N_433,In_624,In_673);
nand U434 (N_434,In_484,In_425);
nor U435 (N_435,In_1088,In_1062);
xnor U436 (N_436,In_813,In_794);
nor U437 (N_437,In_1188,In_379);
xor U438 (N_438,In_1271,In_1089);
xor U439 (N_439,In_192,In_498);
nand U440 (N_440,In_1397,In_306);
nor U441 (N_441,In_398,In_1452);
and U442 (N_442,In_248,In_714);
nor U443 (N_443,In_1244,In_232);
nor U444 (N_444,In_1363,In_589);
xor U445 (N_445,In_1002,In_587);
nand U446 (N_446,In_1272,In_1238);
or U447 (N_447,In_439,In_1263);
nand U448 (N_448,In_91,In_592);
xor U449 (N_449,In_898,In_849);
nand U450 (N_450,In_167,In_936);
and U451 (N_451,In_691,In_146);
nand U452 (N_452,In_336,In_982);
and U453 (N_453,In_533,In_1465);
and U454 (N_454,In_949,In_1069);
or U455 (N_455,In_277,In_1368);
nand U456 (N_456,In_685,In_1298);
nand U457 (N_457,In_1126,In_488);
or U458 (N_458,In_196,In_3);
and U459 (N_459,In_870,In_188);
xor U460 (N_460,In_1222,In_1423);
and U461 (N_461,In_913,In_239);
and U462 (N_462,In_1023,In_36);
and U463 (N_463,In_136,In_847);
nor U464 (N_464,In_21,In_455);
and U465 (N_465,In_1408,In_561);
xnor U466 (N_466,In_1377,In_1223);
and U467 (N_467,In_404,In_247);
nor U468 (N_468,In_1365,In_472);
or U469 (N_469,In_436,In_505);
nand U470 (N_470,In_907,In_413);
nand U471 (N_471,In_1136,In_72);
nor U472 (N_472,In_1358,In_492);
nor U473 (N_473,In_579,In_697);
and U474 (N_474,In_346,In_707);
nor U475 (N_475,In_433,In_228);
xor U476 (N_476,In_980,In_1489);
nor U477 (N_477,In_1026,In_30);
xor U478 (N_478,In_509,In_540);
nand U479 (N_479,In_166,In_803);
nor U480 (N_480,In_1075,In_822);
nand U481 (N_481,In_70,In_955);
xnor U482 (N_482,In_705,In_127);
xor U483 (N_483,In_164,In_595);
nand U484 (N_484,In_593,In_566);
nand U485 (N_485,In_1103,In_1227);
or U486 (N_486,In_565,In_73);
or U487 (N_487,In_1203,In_911);
and U488 (N_488,In_1264,In_1417);
nand U489 (N_489,In_1154,In_970);
nor U490 (N_490,In_145,In_322);
nor U491 (N_491,In_496,In_197);
or U492 (N_492,In_543,In_819);
nor U493 (N_493,In_1013,In_868);
nor U494 (N_494,In_681,In_840);
nor U495 (N_495,In_1353,In_71);
or U496 (N_496,In_770,In_1007);
nand U497 (N_497,In_1461,In_644);
nor U498 (N_498,In_1205,In_1049);
nand U499 (N_499,In_52,In_1357);
nand U500 (N_500,In_260,In_1127);
nand U501 (N_501,In_661,In_1299);
and U502 (N_502,In_217,In_409);
nand U503 (N_503,In_0,In_265);
xor U504 (N_504,In_1025,In_438);
and U505 (N_505,In_914,In_536);
xnor U506 (N_506,In_1245,In_1415);
nor U507 (N_507,In_1084,In_1470);
and U508 (N_508,In_486,In_961);
xnor U509 (N_509,In_524,In_1306);
nor U510 (N_510,In_1322,In_883);
or U511 (N_511,In_573,In_176);
xnor U512 (N_512,In_501,In_280);
nand U513 (N_513,In_609,In_1031);
and U514 (N_514,In_1334,In_383);
nand U515 (N_515,In_121,In_1498);
or U516 (N_516,In_51,In_937);
xor U517 (N_517,In_292,In_371);
nor U518 (N_518,In_198,In_76);
nand U519 (N_519,In_973,In_1394);
xnor U520 (N_520,In_448,In_964);
nand U521 (N_521,In_1111,In_141);
and U522 (N_522,In_1128,In_555);
or U523 (N_523,In_601,In_240);
nand U524 (N_524,In_1017,In_688);
xnor U525 (N_525,In_1064,In_1143);
and U526 (N_526,In_522,In_652);
and U527 (N_527,In_600,In_17);
nor U528 (N_528,In_283,In_808);
and U529 (N_529,In_752,In_942);
or U530 (N_530,In_1219,In_1350);
nand U531 (N_531,In_1027,In_1472);
nor U532 (N_532,In_1006,In_130);
nand U533 (N_533,In_1181,In_45);
and U534 (N_534,In_1068,In_271);
xor U535 (N_535,In_1098,In_948);
xor U536 (N_536,In_653,In_759);
xnor U537 (N_537,In_772,In_194);
nand U538 (N_538,In_1438,In_1384);
nor U539 (N_539,In_1150,In_324);
xor U540 (N_540,In_345,In_908);
and U541 (N_541,In_628,In_829);
xor U542 (N_542,In_1433,In_551);
and U543 (N_543,In_1158,In_327);
xnor U544 (N_544,In_546,In_915);
or U545 (N_545,In_353,In_780);
nand U546 (N_546,In_80,In_93);
nor U547 (N_547,In_963,In_1380);
or U548 (N_548,In_37,In_968);
nor U549 (N_549,In_1427,In_1276);
xor U550 (N_550,In_267,In_1124);
xor U551 (N_551,In_427,In_1116);
and U552 (N_552,In_1345,In_259);
nand U553 (N_553,In_1304,In_1201);
nand U554 (N_554,In_420,In_693);
xnor U555 (N_555,In_838,In_1179);
and U556 (N_556,In_622,In_588);
xnor U557 (N_557,In_1275,In_289);
nand U558 (N_558,In_1146,In_162);
or U559 (N_559,In_170,In_795);
nor U560 (N_560,In_1090,In_116);
and U561 (N_561,In_499,In_263);
nor U562 (N_562,In_1207,In_457);
nand U563 (N_563,In_1277,In_469);
and U564 (N_564,In_1010,In_12);
xor U565 (N_565,In_747,In_542);
nand U566 (N_566,In_1339,In_700);
nor U567 (N_567,In_1372,In_1204);
xnor U568 (N_568,In_577,In_517);
nand U569 (N_569,In_621,In_454);
or U570 (N_570,In_238,In_996);
nor U571 (N_571,In_54,In_258);
or U572 (N_572,In_862,In_504);
xnor U573 (N_573,In_415,In_1217);
nor U574 (N_574,In_261,In_941);
and U575 (N_575,In_2,In_959);
and U576 (N_576,In_347,In_999);
nor U577 (N_577,In_401,In_580);
and U578 (N_578,In_1330,In_660);
xnor U579 (N_579,In_989,In_998);
nor U580 (N_580,In_11,In_1233);
nor U581 (N_581,In_442,In_532);
xnor U582 (N_582,In_1307,In_483);
xnor U583 (N_583,In_219,In_465);
nor U584 (N_584,In_453,In_927);
nor U585 (N_585,In_244,In_466);
or U586 (N_586,In_112,In_350);
or U587 (N_587,In_1409,In_1392);
nand U588 (N_588,In_655,In_871);
or U589 (N_589,In_1463,In_1467);
or U590 (N_590,In_1081,In_539);
or U591 (N_591,In_96,In_616);
or U592 (N_592,In_156,In_1164);
nor U593 (N_593,In_1256,In_1063);
nand U594 (N_594,In_594,In_242);
and U595 (N_595,In_857,In_642);
nor U596 (N_596,In_627,In_125);
and U597 (N_597,In_202,In_940);
xnor U598 (N_598,In_190,In_332);
nor U599 (N_599,In_480,In_1434);
and U600 (N_600,In_357,In_1260);
xnor U601 (N_601,In_456,In_44);
nor U602 (N_602,In_1347,In_1102);
nand U603 (N_603,In_590,In_560);
xor U604 (N_604,In_59,In_331);
and U605 (N_605,In_1073,In_869);
nand U606 (N_606,In_933,In_231);
and U607 (N_607,In_256,In_710);
xnor U608 (N_608,In_711,In_1058);
nand U609 (N_609,In_85,In_124);
or U610 (N_610,In_1186,In_471);
or U611 (N_611,In_470,In_904);
nor U612 (N_612,In_1270,In_1166);
nand U613 (N_613,In_1258,In_490);
nor U614 (N_614,In_896,In_423);
xor U615 (N_615,In_1038,In_6);
or U616 (N_616,In_1328,In_1055);
or U617 (N_617,In_1327,In_447);
xor U618 (N_618,In_230,In_177);
nand U619 (N_619,In_1190,In_718);
nor U620 (N_620,In_1139,In_205);
or U621 (N_621,In_1005,In_450);
nor U622 (N_622,In_1398,In_1493);
xnor U623 (N_623,In_1094,In_763);
nand U624 (N_624,In_641,In_1288);
and U625 (N_625,In_893,In_47);
xnor U626 (N_626,In_1135,In_467);
and U627 (N_627,In_638,In_1485);
xor U628 (N_628,In_329,In_1332);
xor U629 (N_629,In_792,In_1348);
xnor U630 (N_630,In_1171,In_63);
or U631 (N_631,In_348,In_1311);
nand U632 (N_632,In_1341,In_607);
xnor U633 (N_633,In_13,In_951);
xor U634 (N_634,In_1395,In_519);
nor U635 (N_635,In_373,In_113);
and U636 (N_636,In_428,In_178);
or U637 (N_637,In_837,In_538);
and U638 (N_638,In_1351,In_1091);
xor U639 (N_639,In_1312,In_95);
nand U640 (N_640,In_917,In_981);
nor U641 (N_641,In_1067,In_789);
nand U642 (N_642,In_1061,In_632);
or U643 (N_643,In_1120,In_990);
and U644 (N_644,In_106,In_374);
nand U645 (N_645,In_441,In_793);
nor U646 (N_646,In_771,In_1420);
xnor U647 (N_647,In_689,In_812);
or U648 (N_648,In_743,In_34);
and U649 (N_649,In_56,In_1319);
or U650 (N_650,In_701,In_1248);
nand U651 (N_651,In_1303,In_235);
nand U652 (N_652,In_892,In_969);
nand U653 (N_653,In_521,In_902);
nor U654 (N_654,In_1109,In_1138);
nand U655 (N_655,In_224,In_512);
or U656 (N_656,In_1115,In_339);
and U657 (N_657,In_245,In_640);
and U658 (N_658,In_713,In_875);
nand U659 (N_659,In_1134,In_1177);
or U660 (N_660,In_1262,In_266);
nor U661 (N_661,In_440,In_647);
or U662 (N_662,In_414,In_582);
nand U663 (N_663,In_396,In_1121);
nor U664 (N_664,In_922,In_1443);
and U665 (N_665,In_1083,In_1371);
nand U666 (N_666,In_559,In_60);
or U667 (N_667,In_626,In_137);
or U668 (N_668,In_598,In_796);
nor U669 (N_669,In_200,In_1376);
and U670 (N_670,In_574,In_148);
and U671 (N_671,In_67,In_1464);
nor U672 (N_672,In_553,In_28);
and U673 (N_673,In_783,In_811);
or U674 (N_674,In_725,In_1436);
nand U675 (N_675,In_406,In_1033);
nor U676 (N_676,In_1297,In_570);
nand U677 (N_677,In_1257,In_1431);
or U678 (N_678,In_226,In_1001);
xnor U679 (N_679,In_449,In_183);
xor U680 (N_680,In_343,In_189);
or U681 (N_681,In_530,In_293);
and U682 (N_682,In_535,In_1228);
xnor U683 (N_683,In_187,In_912);
or U684 (N_684,In_1,In_1003);
nor U685 (N_685,In_1198,In_487);
nor U686 (N_686,In_35,In_385);
nor U687 (N_687,In_766,In_302);
and U688 (N_688,In_664,In_781);
and U689 (N_689,In_387,In_716);
and U690 (N_690,In_1273,In_682);
nand U691 (N_691,In_666,In_1185);
and U692 (N_692,In_1246,In_1355);
xnor U693 (N_693,In_643,In_349);
nand U694 (N_694,In_1153,In_1289);
and U695 (N_695,In_1362,In_285);
nor U696 (N_696,In_211,In_16);
and U697 (N_697,In_1144,In_88);
or U698 (N_698,In_1085,In_1051);
xor U699 (N_699,In_363,In_1301);
nand U700 (N_700,In_562,In_1369);
and U701 (N_701,In_842,In_920);
nand U702 (N_702,In_1161,In_676);
nand U703 (N_703,In_417,In_1014);
xor U704 (N_704,In_930,In_597);
or U705 (N_705,In_405,In_757);
nor U706 (N_706,In_1009,In_511);
nor U707 (N_707,In_1224,In_786);
nor U708 (N_708,In_1313,In_1421);
xnor U709 (N_709,In_749,In_321);
and U710 (N_710,In_337,In_1016);
xor U711 (N_711,In_317,In_479);
nor U712 (N_712,In_1163,In_1317);
xnor U713 (N_713,In_274,In_75);
xnor U714 (N_714,In_49,In_1172);
or U715 (N_715,In_687,In_1484);
nand U716 (N_716,In_636,In_1165);
xnor U717 (N_717,In_1269,In_977);
nor U718 (N_718,In_477,In_1344);
or U719 (N_719,In_1096,In_40);
xnor U720 (N_720,In_696,In_380);
xnor U721 (N_721,In_305,In_526);
nor U722 (N_722,In_767,In_328);
or U723 (N_723,In_799,In_315);
or U724 (N_724,In_1159,In_208);
nand U725 (N_725,In_269,In_1375);
or U726 (N_726,In_147,In_723);
nor U727 (N_727,In_66,In_614);
and U728 (N_728,In_422,In_906);
and U729 (N_729,In_300,In_975);
xnor U730 (N_730,In_946,In_995);
nor U731 (N_731,In_1265,In_860);
xnor U732 (N_732,In_1457,In_1226);
or U733 (N_733,In_1000,In_708);
and U734 (N_734,In_128,In_1492);
nor U735 (N_735,In_1076,In_797);
nor U736 (N_736,In_18,In_1048);
xnor U737 (N_737,In_1216,In_885);
nand U738 (N_738,In_890,In_1287);
nand U739 (N_739,In_832,In_768);
nor U740 (N_740,In_1473,In_241);
nand U741 (N_741,In_1234,In_880);
nor U742 (N_742,In_637,In_432);
nor U743 (N_743,In_715,In_204);
xor U744 (N_744,In_599,In_762);
and U745 (N_745,In_132,In_461);
xnor U746 (N_746,In_1021,In_393);
nand U747 (N_747,In_861,In_1259);
xor U748 (N_748,In_750,In_719);
and U749 (N_749,In_800,In_1119);
nand U750 (N_750,In_775,In_1112);
xor U751 (N_751,In_449,In_1220);
nor U752 (N_752,In_1433,In_690);
nor U753 (N_753,In_1476,In_509);
nand U754 (N_754,In_720,In_796);
nand U755 (N_755,In_1089,In_956);
nand U756 (N_756,In_18,In_1429);
nor U757 (N_757,In_54,In_1381);
nand U758 (N_758,In_1110,In_44);
nand U759 (N_759,In_1492,In_731);
nand U760 (N_760,In_71,In_337);
xnor U761 (N_761,In_817,In_205);
and U762 (N_762,In_68,In_287);
nor U763 (N_763,In_1144,In_1270);
or U764 (N_764,In_644,In_68);
nor U765 (N_765,In_977,In_1101);
or U766 (N_766,In_593,In_401);
xor U767 (N_767,In_99,In_1351);
xor U768 (N_768,In_605,In_284);
and U769 (N_769,In_875,In_553);
nor U770 (N_770,In_1353,In_1013);
nor U771 (N_771,In_751,In_687);
xnor U772 (N_772,In_44,In_1280);
xor U773 (N_773,In_279,In_76);
nor U774 (N_774,In_38,In_860);
nor U775 (N_775,In_471,In_878);
and U776 (N_776,In_407,In_1236);
xnor U777 (N_777,In_1100,In_487);
nor U778 (N_778,In_1159,In_642);
or U779 (N_779,In_1134,In_886);
nor U780 (N_780,In_994,In_248);
nand U781 (N_781,In_631,In_268);
nand U782 (N_782,In_423,In_88);
xnor U783 (N_783,In_949,In_21);
xor U784 (N_784,In_457,In_687);
xor U785 (N_785,In_503,In_640);
and U786 (N_786,In_200,In_534);
nand U787 (N_787,In_1310,In_675);
or U788 (N_788,In_297,In_1389);
and U789 (N_789,In_1036,In_590);
nand U790 (N_790,In_863,In_683);
nor U791 (N_791,In_806,In_286);
and U792 (N_792,In_338,In_736);
nand U793 (N_793,In_364,In_1292);
nand U794 (N_794,In_603,In_632);
or U795 (N_795,In_965,In_1329);
and U796 (N_796,In_668,In_130);
xor U797 (N_797,In_1142,In_736);
or U798 (N_798,In_158,In_1293);
and U799 (N_799,In_124,In_158);
xnor U800 (N_800,In_269,In_1281);
and U801 (N_801,In_176,In_693);
and U802 (N_802,In_348,In_64);
or U803 (N_803,In_205,In_1114);
and U804 (N_804,In_98,In_772);
or U805 (N_805,In_536,In_1163);
nor U806 (N_806,In_1245,In_1462);
or U807 (N_807,In_8,In_940);
or U808 (N_808,In_1462,In_993);
xor U809 (N_809,In_1069,In_321);
or U810 (N_810,In_173,In_920);
nor U811 (N_811,In_649,In_98);
nor U812 (N_812,In_1279,In_818);
and U813 (N_813,In_743,In_677);
nor U814 (N_814,In_874,In_214);
nor U815 (N_815,In_200,In_381);
nor U816 (N_816,In_413,In_1434);
xor U817 (N_817,In_270,In_1077);
and U818 (N_818,In_263,In_1451);
and U819 (N_819,In_1085,In_429);
nand U820 (N_820,In_1412,In_101);
xor U821 (N_821,In_328,In_1203);
or U822 (N_822,In_1050,In_179);
nand U823 (N_823,In_1061,In_775);
xor U824 (N_824,In_687,In_639);
nand U825 (N_825,In_235,In_1092);
or U826 (N_826,In_1166,In_900);
nor U827 (N_827,In_1042,In_164);
xnor U828 (N_828,In_299,In_501);
or U829 (N_829,In_539,In_482);
xnor U830 (N_830,In_1394,In_960);
nand U831 (N_831,In_430,In_1474);
nor U832 (N_832,In_343,In_48);
and U833 (N_833,In_1108,In_753);
xnor U834 (N_834,In_1395,In_823);
nor U835 (N_835,In_1387,In_188);
and U836 (N_836,In_1309,In_1375);
nor U837 (N_837,In_456,In_572);
or U838 (N_838,In_417,In_1177);
or U839 (N_839,In_622,In_795);
xnor U840 (N_840,In_269,In_1160);
or U841 (N_841,In_862,In_277);
nand U842 (N_842,In_43,In_853);
or U843 (N_843,In_1457,In_1387);
nand U844 (N_844,In_914,In_1414);
xor U845 (N_845,In_1495,In_1490);
xor U846 (N_846,In_1167,In_191);
xnor U847 (N_847,In_381,In_1078);
nor U848 (N_848,In_72,In_30);
nand U849 (N_849,In_5,In_1403);
or U850 (N_850,In_1232,In_267);
nand U851 (N_851,In_1193,In_1338);
and U852 (N_852,In_157,In_1320);
nand U853 (N_853,In_725,In_108);
xor U854 (N_854,In_466,In_764);
xnor U855 (N_855,In_1080,In_981);
xnor U856 (N_856,In_479,In_1046);
or U857 (N_857,In_666,In_1098);
nor U858 (N_858,In_1031,In_959);
or U859 (N_859,In_679,In_771);
nand U860 (N_860,In_1314,In_409);
and U861 (N_861,In_1211,In_168);
and U862 (N_862,In_1401,In_261);
xor U863 (N_863,In_1223,In_238);
xor U864 (N_864,In_377,In_1178);
xor U865 (N_865,In_499,In_336);
nor U866 (N_866,In_523,In_611);
nand U867 (N_867,In_1423,In_811);
nor U868 (N_868,In_128,In_809);
nor U869 (N_869,In_364,In_721);
xor U870 (N_870,In_214,In_428);
nand U871 (N_871,In_708,In_898);
and U872 (N_872,In_1474,In_347);
nor U873 (N_873,In_269,In_1111);
and U874 (N_874,In_1060,In_188);
nor U875 (N_875,In_727,In_1058);
nor U876 (N_876,In_1061,In_517);
and U877 (N_877,In_1174,In_383);
nor U878 (N_878,In_331,In_236);
nand U879 (N_879,In_713,In_82);
nand U880 (N_880,In_550,In_800);
nor U881 (N_881,In_10,In_828);
and U882 (N_882,In_601,In_873);
or U883 (N_883,In_120,In_146);
xor U884 (N_884,In_938,In_1494);
nand U885 (N_885,In_587,In_452);
xnor U886 (N_886,In_1292,In_1444);
nor U887 (N_887,In_1233,In_423);
nand U888 (N_888,In_737,In_5);
or U889 (N_889,In_1415,In_615);
nor U890 (N_890,In_1441,In_773);
and U891 (N_891,In_256,In_497);
xor U892 (N_892,In_507,In_1346);
nor U893 (N_893,In_997,In_852);
nor U894 (N_894,In_1454,In_150);
nor U895 (N_895,In_923,In_505);
xor U896 (N_896,In_519,In_765);
xor U897 (N_897,In_536,In_143);
nor U898 (N_898,In_477,In_1404);
xor U899 (N_899,In_1402,In_675);
xor U900 (N_900,In_1090,In_1056);
or U901 (N_901,In_546,In_1061);
and U902 (N_902,In_500,In_168);
nand U903 (N_903,In_505,In_310);
and U904 (N_904,In_1089,In_164);
or U905 (N_905,In_449,In_172);
nand U906 (N_906,In_52,In_800);
xor U907 (N_907,In_1293,In_1276);
and U908 (N_908,In_1431,In_904);
nand U909 (N_909,In_1114,In_1311);
xnor U910 (N_910,In_1190,In_810);
xor U911 (N_911,In_964,In_316);
and U912 (N_912,In_946,In_1323);
nor U913 (N_913,In_1072,In_934);
nor U914 (N_914,In_790,In_1140);
nor U915 (N_915,In_308,In_267);
and U916 (N_916,In_78,In_209);
nand U917 (N_917,In_1115,In_699);
nand U918 (N_918,In_1229,In_345);
and U919 (N_919,In_301,In_1281);
and U920 (N_920,In_206,In_22);
nand U921 (N_921,In_1125,In_999);
xor U922 (N_922,In_303,In_417);
xnor U923 (N_923,In_1145,In_295);
nand U924 (N_924,In_1013,In_246);
and U925 (N_925,In_1428,In_710);
or U926 (N_926,In_989,In_681);
xnor U927 (N_927,In_837,In_973);
nor U928 (N_928,In_1250,In_526);
xor U929 (N_929,In_1151,In_1);
nand U930 (N_930,In_641,In_1112);
nand U931 (N_931,In_585,In_420);
xor U932 (N_932,In_1399,In_432);
xnor U933 (N_933,In_987,In_315);
xnor U934 (N_934,In_354,In_1381);
nor U935 (N_935,In_621,In_360);
nand U936 (N_936,In_0,In_927);
nor U937 (N_937,In_684,In_1129);
xnor U938 (N_938,In_356,In_507);
nand U939 (N_939,In_1033,In_305);
and U940 (N_940,In_1106,In_470);
xnor U941 (N_941,In_313,In_1323);
or U942 (N_942,In_685,In_636);
and U943 (N_943,In_101,In_216);
xnor U944 (N_944,In_1334,In_57);
nand U945 (N_945,In_1268,In_1145);
nand U946 (N_946,In_1494,In_650);
and U947 (N_947,In_650,In_1277);
or U948 (N_948,In_461,In_1316);
nand U949 (N_949,In_726,In_1402);
nor U950 (N_950,In_1426,In_1031);
xor U951 (N_951,In_1306,In_673);
nor U952 (N_952,In_514,In_570);
nor U953 (N_953,In_1214,In_116);
or U954 (N_954,In_846,In_1404);
nand U955 (N_955,In_319,In_869);
nand U956 (N_956,In_1079,In_1351);
xor U957 (N_957,In_751,In_402);
xor U958 (N_958,In_665,In_939);
and U959 (N_959,In_1192,In_1398);
xnor U960 (N_960,In_940,In_1380);
nor U961 (N_961,In_1190,In_290);
and U962 (N_962,In_991,In_600);
nor U963 (N_963,In_680,In_696);
xnor U964 (N_964,In_1385,In_1342);
or U965 (N_965,In_1327,In_837);
or U966 (N_966,In_994,In_139);
and U967 (N_967,In_520,In_747);
nor U968 (N_968,In_652,In_189);
or U969 (N_969,In_993,In_302);
nor U970 (N_970,In_123,In_187);
xor U971 (N_971,In_810,In_1359);
xnor U972 (N_972,In_989,In_25);
xor U973 (N_973,In_975,In_253);
or U974 (N_974,In_1488,In_1234);
nand U975 (N_975,In_757,In_1294);
nand U976 (N_976,In_1012,In_209);
or U977 (N_977,In_697,In_1133);
xor U978 (N_978,In_1035,In_1394);
nor U979 (N_979,In_1439,In_734);
nor U980 (N_980,In_815,In_155);
and U981 (N_981,In_1457,In_335);
nor U982 (N_982,In_4,In_189);
nand U983 (N_983,In_1136,In_569);
or U984 (N_984,In_116,In_1062);
nand U985 (N_985,In_881,In_217);
or U986 (N_986,In_196,In_173);
or U987 (N_987,In_112,In_205);
nor U988 (N_988,In_1181,In_570);
nand U989 (N_989,In_630,In_527);
nand U990 (N_990,In_116,In_682);
nor U991 (N_991,In_755,In_1184);
nand U992 (N_992,In_1344,In_18);
and U993 (N_993,In_471,In_1296);
or U994 (N_994,In_1217,In_1211);
nor U995 (N_995,In_1075,In_1081);
and U996 (N_996,In_738,In_1363);
nand U997 (N_997,In_1398,In_1134);
xnor U998 (N_998,In_908,In_417);
xnor U999 (N_999,In_223,In_464);
nand U1000 (N_1000,In_1420,In_1025);
nor U1001 (N_1001,In_811,In_887);
nand U1002 (N_1002,In_594,In_853);
or U1003 (N_1003,In_296,In_476);
nor U1004 (N_1004,In_1471,In_173);
nor U1005 (N_1005,In_752,In_1131);
and U1006 (N_1006,In_1430,In_774);
and U1007 (N_1007,In_1408,In_471);
and U1008 (N_1008,In_340,In_422);
nand U1009 (N_1009,In_123,In_68);
nand U1010 (N_1010,In_1328,In_281);
or U1011 (N_1011,In_1263,In_978);
or U1012 (N_1012,In_1098,In_1494);
xor U1013 (N_1013,In_164,In_855);
nor U1014 (N_1014,In_296,In_1467);
or U1015 (N_1015,In_631,In_701);
nor U1016 (N_1016,In_1432,In_147);
and U1017 (N_1017,In_1327,In_685);
nor U1018 (N_1018,In_91,In_1251);
nor U1019 (N_1019,In_38,In_1105);
and U1020 (N_1020,In_378,In_408);
and U1021 (N_1021,In_977,In_873);
or U1022 (N_1022,In_1474,In_207);
xnor U1023 (N_1023,In_1203,In_455);
nand U1024 (N_1024,In_658,In_311);
xnor U1025 (N_1025,In_6,In_1221);
and U1026 (N_1026,In_155,In_675);
xor U1027 (N_1027,In_571,In_338);
and U1028 (N_1028,In_550,In_487);
or U1029 (N_1029,In_907,In_646);
and U1030 (N_1030,In_728,In_903);
and U1031 (N_1031,In_1306,In_210);
nor U1032 (N_1032,In_894,In_1022);
nor U1033 (N_1033,In_814,In_105);
nand U1034 (N_1034,In_145,In_1117);
nor U1035 (N_1035,In_804,In_1376);
xnor U1036 (N_1036,In_849,In_42);
and U1037 (N_1037,In_451,In_945);
nor U1038 (N_1038,In_1365,In_36);
nor U1039 (N_1039,In_130,In_835);
or U1040 (N_1040,In_173,In_45);
xnor U1041 (N_1041,In_235,In_284);
or U1042 (N_1042,In_70,In_578);
and U1043 (N_1043,In_1428,In_414);
or U1044 (N_1044,In_333,In_1132);
nand U1045 (N_1045,In_1444,In_663);
nand U1046 (N_1046,In_441,In_729);
and U1047 (N_1047,In_880,In_1450);
xnor U1048 (N_1048,In_1066,In_1464);
and U1049 (N_1049,In_29,In_1201);
or U1050 (N_1050,In_880,In_417);
nand U1051 (N_1051,In_514,In_821);
or U1052 (N_1052,In_554,In_424);
xor U1053 (N_1053,In_174,In_1094);
nor U1054 (N_1054,In_1157,In_1409);
nor U1055 (N_1055,In_818,In_492);
nand U1056 (N_1056,In_1396,In_1052);
xnor U1057 (N_1057,In_1210,In_778);
or U1058 (N_1058,In_518,In_151);
nor U1059 (N_1059,In_1177,In_284);
and U1060 (N_1060,In_1179,In_391);
or U1061 (N_1061,In_15,In_338);
nand U1062 (N_1062,In_1404,In_1020);
xor U1063 (N_1063,In_278,In_1290);
xnor U1064 (N_1064,In_1138,In_851);
and U1065 (N_1065,In_425,In_955);
nor U1066 (N_1066,In_68,In_422);
xor U1067 (N_1067,In_918,In_1486);
nand U1068 (N_1068,In_32,In_1355);
or U1069 (N_1069,In_775,In_823);
xnor U1070 (N_1070,In_382,In_536);
nand U1071 (N_1071,In_520,In_1113);
nand U1072 (N_1072,In_922,In_115);
nor U1073 (N_1073,In_397,In_336);
nor U1074 (N_1074,In_698,In_51);
or U1075 (N_1075,In_659,In_814);
nor U1076 (N_1076,In_1401,In_138);
nor U1077 (N_1077,In_84,In_298);
and U1078 (N_1078,In_1454,In_1327);
nand U1079 (N_1079,In_114,In_233);
nand U1080 (N_1080,In_1492,In_1106);
and U1081 (N_1081,In_368,In_264);
nor U1082 (N_1082,In_1181,In_645);
nor U1083 (N_1083,In_336,In_1205);
or U1084 (N_1084,In_392,In_313);
or U1085 (N_1085,In_1431,In_29);
nand U1086 (N_1086,In_1314,In_624);
nor U1087 (N_1087,In_733,In_576);
nor U1088 (N_1088,In_461,In_1335);
nor U1089 (N_1089,In_711,In_1486);
nor U1090 (N_1090,In_941,In_513);
nand U1091 (N_1091,In_889,In_1131);
nor U1092 (N_1092,In_1498,In_78);
xor U1093 (N_1093,In_177,In_34);
and U1094 (N_1094,In_1465,In_405);
nand U1095 (N_1095,In_376,In_706);
or U1096 (N_1096,In_1028,In_1180);
nor U1097 (N_1097,In_190,In_1216);
nor U1098 (N_1098,In_453,In_114);
nor U1099 (N_1099,In_1016,In_1424);
nand U1100 (N_1100,In_1400,In_755);
nand U1101 (N_1101,In_1340,In_351);
nor U1102 (N_1102,In_1092,In_990);
nand U1103 (N_1103,In_677,In_854);
or U1104 (N_1104,In_772,In_1078);
and U1105 (N_1105,In_75,In_581);
and U1106 (N_1106,In_543,In_90);
and U1107 (N_1107,In_1402,In_1336);
nand U1108 (N_1108,In_426,In_1341);
and U1109 (N_1109,In_21,In_1343);
or U1110 (N_1110,In_763,In_1185);
and U1111 (N_1111,In_149,In_311);
or U1112 (N_1112,In_1231,In_821);
nand U1113 (N_1113,In_1127,In_984);
nand U1114 (N_1114,In_929,In_1370);
xnor U1115 (N_1115,In_207,In_347);
nor U1116 (N_1116,In_1456,In_1053);
xor U1117 (N_1117,In_1219,In_658);
xor U1118 (N_1118,In_720,In_664);
or U1119 (N_1119,In_1087,In_404);
xor U1120 (N_1120,In_1439,In_59);
and U1121 (N_1121,In_1330,In_752);
xor U1122 (N_1122,In_470,In_322);
or U1123 (N_1123,In_17,In_937);
nor U1124 (N_1124,In_284,In_572);
and U1125 (N_1125,In_2,In_1163);
xnor U1126 (N_1126,In_1225,In_364);
and U1127 (N_1127,In_374,In_1361);
nor U1128 (N_1128,In_1062,In_1206);
and U1129 (N_1129,In_666,In_1050);
xor U1130 (N_1130,In_18,In_1174);
nor U1131 (N_1131,In_654,In_1455);
nand U1132 (N_1132,In_64,In_486);
nor U1133 (N_1133,In_243,In_13);
xor U1134 (N_1134,In_1340,In_644);
xnor U1135 (N_1135,In_595,In_971);
xnor U1136 (N_1136,In_478,In_636);
xnor U1137 (N_1137,In_328,In_1327);
or U1138 (N_1138,In_1171,In_475);
nor U1139 (N_1139,In_44,In_228);
xor U1140 (N_1140,In_963,In_734);
xor U1141 (N_1141,In_61,In_815);
or U1142 (N_1142,In_1263,In_827);
or U1143 (N_1143,In_175,In_1336);
or U1144 (N_1144,In_1388,In_641);
nand U1145 (N_1145,In_1414,In_694);
or U1146 (N_1146,In_151,In_545);
nand U1147 (N_1147,In_1085,In_304);
xnor U1148 (N_1148,In_46,In_268);
xnor U1149 (N_1149,In_1156,In_888);
nor U1150 (N_1150,In_874,In_865);
and U1151 (N_1151,In_726,In_571);
xnor U1152 (N_1152,In_241,In_847);
nor U1153 (N_1153,In_916,In_908);
nand U1154 (N_1154,In_293,In_668);
nand U1155 (N_1155,In_825,In_151);
nand U1156 (N_1156,In_1180,In_1077);
nand U1157 (N_1157,In_682,In_774);
and U1158 (N_1158,In_252,In_859);
and U1159 (N_1159,In_704,In_120);
nand U1160 (N_1160,In_462,In_524);
nor U1161 (N_1161,In_367,In_632);
nor U1162 (N_1162,In_272,In_192);
xor U1163 (N_1163,In_473,In_929);
and U1164 (N_1164,In_719,In_111);
or U1165 (N_1165,In_1195,In_592);
nand U1166 (N_1166,In_337,In_990);
nor U1167 (N_1167,In_713,In_136);
and U1168 (N_1168,In_140,In_1122);
xnor U1169 (N_1169,In_718,In_1355);
xor U1170 (N_1170,In_950,In_1266);
and U1171 (N_1171,In_880,In_117);
nor U1172 (N_1172,In_169,In_645);
nor U1173 (N_1173,In_1008,In_1474);
xor U1174 (N_1174,In_653,In_583);
xnor U1175 (N_1175,In_1077,In_891);
xnor U1176 (N_1176,In_529,In_835);
or U1177 (N_1177,In_990,In_751);
xnor U1178 (N_1178,In_686,In_692);
and U1179 (N_1179,In_1450,In_685);
nand U1180 (N_1180,In_828,In_316);
or U1181 (N_1181,In_121,In_319);
nand U1182 (N_1182,In_765,In_1108);
xor U1183 (N_1183,In_64,In_1453);
nand U1184 (N_1184,In_646,In_219);
nand U1185 (N_1185,In_1084,In_1201);
nand U1186 (N_1186,In_1217,In_413);
nor U1187 (N_1187,In_232,In_480);
or U1188 (N_1188,In_471,In_972);
or U1189 (N_1189,In_175,In_1014);
xor U1190 (N_1190,In_788,In_386);
xor U1191 (N_1191,In_762,In_1051);
or U1192 (N_1192,In_444,In_1355);
nand U1193 (N_1193,In_290,In_485);
and U1194 (N_1194,In_1229,In_710);
and U1195 (N_1195,In_722,In_963);
xnor U1196 (N_1196,In_7,In_501);
nor U1197 (N_1197,In_864,In_1110);
and U1198 (N_1198,In_123,In_1149);
nand U1199 (N_1199,In_1448,In_966);
nor U1200 (N_1200,In_1079,In_1493);
xor U1201 (N_1201,In_866,In_229);
nand U1202 (N_1202,In_857,In_283);
nand U1203 (N_1203,In_382,In_151);
and U1204 (N_1204,In_960,In_753);
and U1205 (N_1205,In_1055,In_18);
xor U1206 (N_1206,In_1085,In_1427);
xor U1207 (N_1207,In_710,In_159);
and U1208 (N_1208,In_11,In_718);
nand U1209 (N_1209,In_1482,In_425);
xor U1210 (N_1210,In_368,In_56);
nor U1211 (N_1211,In_729,In_1456);
nor U1212 (N_1212,In_1035,In_1253);
xnor U1213 (N_1213,In_1091,In_461);
xor U1214 (N_1214,In_1411,In_166);
and U1215 (N_1215,In_1043,In_329);
nor U1216 (N_1216,In_578,In_1390);
or U1217 (N_1217,In_915,In_239);
nor U1218 (N_1218,In_741,In_1186);
nand U1219 (N_1219,In_1229,In_311);
nand U1220 (N_1220,In_758,In_1408);
nor U1221 (N_1221,In_428,In_847);
nor U1222 (N_1222,In_60,In_151);
nor U1223 (N_1223,In_31,In_1118);
xor U1224 (N_1224,In_238,In_520);
and U1225 (N_1225,In_1190,In_365);
nor U1226 (N_1226,In_1319,In_1244);
nand U1227 (N_1227,In_656,In_784);
or U1228 (N_1228,In_1474,In_1092);
nor U1229 (N_1229,In_606,In_766);
xor U1230 (N_1230,In_61,In_1040);
and U1231 (N_1231,In_1233,In_195);
nor U1232 (N_1232,In_419,In_1191);
nand U1233 (N_1233,In_167,In_129);
nand U1234 (N_1234,In_191,In_526);
xor U1235 (N_1235,In_849,In_996);
or U1236 (N_1236,In_585,In_794);
nand U1237 (N_1237,In_1038,In_177);
nand U1238 (N_1238,In_813,In_755);
xor U1239 (N_1239,In_507,In_479);
xor U1240 (N_1240,In_44,In_126);
nand U1241 (N_1241,In_1089,In_434);
xor U1242 (N_1242,In_649,In_525);
nor U1243 (N_1243,In_12,In_1142);
and U1244 (N_1244,In_1390,In_1068);
xor U1245 (N_1245,In_594,In_2);
or U1246 (N_1246,In_327,In_64);
xor U1247 (N_1247,In_25,In_949);
or U1248 (N_1248,In_1160,In_238);
nand U1249 (N_1249,In_253,In_802);
xnor U1250 (N_1250,In_1340,In_1415);
nand U1251 (N_1251,In_730,In_650);
or U1252 (N_1252,In_1463,In_1284);
nor U1253 (N_1253,In_1183,In_784);
and U1254 (N_1254,In_938,In_1193);
and U1255 (N_1255,In_978,In_1190);
nand U1256 (N_1256,In_304,In_159);
and U1257 (N_1257,In_75,In_349);
xnor U1258 (N_1258,In_988,In_69);
nand U1259 (N_1259,In_329,In_1403);
or U1260 (N_1260,In_125,In_907);
or U1261 (N_1261,In_1453,In_690);
xor U1262 (N_1262,In_719,In_346);
nand U1263 (N_1263,In_789,In_1120);
xnor U1264 (N_1264,In_257,In_1130);
xnor U1265 (N_1265,In_26,In_1494);
or U1266 (N_1266,In_716,In_275);
nand U1267 (N_1267,In_646,In_996);
nand U1268 (N_1268,In_1420,In_775);
xnor U1269 (N_1269,In_632,In_244);
nand U1270 (N_1270,In_403,In_1367);
and U1271 (N_1271,In_323,In_290);
or U1272 (N_1272,In_471,In_1086);
xnor U1273 (N_1273,In_15,In_741);
or U1274 (N_1274,In_387,In_1275);
and U1275 (N_1275,In_50,In_1289);
nor U1276 (N_1276,In_1296,In_963);
or U1277 (N_1277,In_151,In_1388);
and U1278 (N_1278,In_155,In_1145);
nand U1279 (N_1279,In_123,In_302);
nor U1280 (N_1280,In_153,In_277);
xor U1281 (N_1281,In_946,In_840);
nand U1282 (N_1282,In_232,In_818);
or U1283 (N_1283,In_538,In_856);
or U1284 (N_1284,In_442,In_137);
xor U1285 (N_1285,In_631,In_840);
or U1286 (N_1286,In_1377,In_311);
or U1287 (N_1287,In_1025,In_1126);
nand U1288 (N_1288,In_1080,In_652);
and U1289 (N_1289,In_943,In_449);
nor U1290 (N_1290,In_607,In_1411);
or U1291 (N_1291,In_897,In_989);
nand U1292 (N_1292,In_1343,In_1487);
xnor U1293 (N_1293,In_1437,In_83);
and U1294 (N_1294,In_655,In_1469);
nor U1295 (N_1295,In_514,In_445);
nor U1296 (N_1296,In_1411,In_1259);
nor U1297 (N_1297,In_1398,In_123);
or U1298 (N_1298,In_231,In_1427);
xor U1299 (N_1299,In_323,In_1165);
and U1300 (N_1300,In_775,In_781);
nand U1301 (N_1301,In_129,In_388);
nor U1302 (N_1302,In_1333,In_1103);
nor U1303 (N_1303,In_586,In_309);
and U1304 (N_1304,In_274,In_1448);
or U1305 (N_1305,In_1080,In_436);
xor U1306 (N_1306,In_1021,In_36);
and U1307 (N_1307,In_1011,In_210);
or U1308 (N_1308,In_1014,In_1089);
or U1309 (N_1309,In_336,In_678);
or U1310 (N_1310,In_538,In_928);
and U1311 (N_1311,In_295,In_1026);
nor U1312 (N_1312,In_481,In_163);
and U1313 (N_1313,In_416,In_243);
and U1314 (N_1314,In_931,In_1048);
nor U1315 (N_1315,In_281,In_796);
or U1316 (N_1316,In_43,In_725);
and U1317 (N_1317,In_590,In_431);
nor U1318 (N_1318,In_535,In_215);
xor U1319 (N_1319,In_1113,In_844);
nor U1320 (N_1320,In_719,In_1018);
xor U1321 (N_1321,In_1012,In_308);
nand U1322 (N_1322,In_557,In_946);
xor U1323 (N_1323,In_540,In_1044);
nand U1324 (N_1324,In_910,In_700);
and U1325 (N_1325,In_963,In_448);
and U1326 (N_1326,In_1231,In_1176);
nand U1327 (N_1327,In_1179,In_1135);
or U1328 (N_1328,In_656,In_1126);
and U1329 (N_1329,In_646,In_57);
and U1330 (N_1330,In_1034,In_970);
xor U1331 (N_1331,In_1021,In_753);
or U1332 (N_1332,In_1103,In_1269);
nand U1333 (N_1333,In_75,In_139);
or U1334 (N_1334,In_723,In_612);
or U1335 (N_1335,In_699,In_1238);
nor U1336 (N_1336,In_1442,In_1419);
and U1337 (N_1337,In_1143,In_1294);
and U1338 (N_1338,In_1490,In_545);
xnor U1339 (N_1339,In_917,In_1210);
nor U1340 (N_1340,In_546,In_1369);
nor U1341 (N_1341,In_983,In_2);
and U1342 (N_1342,In_582,In_491);
xnor U1343 (N_1343,In_115,In_1199);
and U1344 (N_1344,In_869,In_1196);
nor U1345 (N_1345,In_702,In_1081);
nor U1346 (N_1346,In_499,In_378);
xnor U1347 (N_1347,In_234,In_1147);
or U1348 (N_1348,In_1039,In_529);
and U1349 (N_1349,In_344,In_1207);
xor U1350 (N_1350,In_645,In_638);
or U1351 (N_1351,In_828,In_14);
nand U1352 (N_1352,In_91,In_1062);
nor U1353 (N_1353,In_1448,In_526);
xor U1354 (N_1354,In_529,In_114);
xor U1355 (N_1355,In_1285,In_1468);
xnor U1356 (N_1356,In_797,In_585);
nor U1357 (N_1357,In_1137,In_92);
and U1358 (N_1358,In_1114,In_390);
and U1359 (N_1359,In_248,In_165);
nand U1360 (N_1360,In_1450,In_169);
nand U1361 (N_1361,In_451,In_869);
xor U1362 (N_1362,In_223,In_700);
nor U1363 (N_1363,In_1071,In_650);
and U1364 (N_1364,In_108,In_1347);
xnor U1365 (N_1365,In_499,In_1053);
and U1366 (N_1366,In_554,In_1181);
or U1367 (N_1367,In_491,In_359);
xor U1368 (N_1368,In_1013,In_72);
or U1369 (N_1369,In_870,In_567);
nor U1370 (N_1370,In_138,In_1220);
nor U1371 (N_1371,In_448,In_1235);
or U1372 (N_1372,In_1389,In_1182);
xnor U1373 (N_1373,In_746,In_1091);
xnor U1374 (N_1374,In_1485,In_1020);
or U1375 (N_1375,In_230,In_1059);
and U1376 (N_1376,In_660,In_1134);
and U1377 (N_1377,In_737,In_122);
or U1378 (N_1378,In_1243,In_1250);
or U1379 (N_1379,In_1135,In_1419);
and U1380 (N_1380,In_1428,In_1281);
or U1381 (N_1381,In_1181,In_1482);
nor U1382 (N_1382,In_717,In_1032);
and U1383 (N_1383,In_120,In_440);
nor U1384 (N_1384,In_165,In_960);
nand U1385 (N_1385,In_1054,In_538);
nor U1386 (N_1386,In_1369,In_811);
nor U1387 (N_1387,In_1285,In_679);
nand U1388 (N_1388,In_284,In_849);
or U1389 (N_1389,In_1208,In_355);
and U1390 (N_1390,In_200,In_903);
or U1391 (N_1391,In_1007,In_1138);
nor U1392 (N_1392,In_375,In_123);
xor U1393 (N_1393,In_83,In_13);
xor U1394 (N_1394,In_486,In_728);
or U1395 (N_1395,In_1169,In_1461);
nor U1396 (N_1396,In_190,In_265);
and U1397 (N_1397,In_1477,In_134);
or U1398 (N_1398,In_1029,In_1404);
nor U1399 (N_1399,In_259,In_1389);
nand U1400 (N_1400,In_556,In_1279);
nand U1401 (N_1401,In_817,In_1177);
nand U1402 (N_1402,In_79,In_329);
nor U1403 (N_1403,In_855,In_1000);
or U1404 (N_1404,In_269,In_1227);
nand U1405 (N_1405,In_12,In_97);
and U1406 (N_1406,In_1053,In_1062);
or U1407 (N_1407,In_857,In_696);
xor U1408 (N_1408,In_645,In_927);
or U1409 (N_1409,In_578,In_1015);
nand U1410 (N_1410,In_1387,In_938);
or U1411 (N_1411,In_104,In_295);
xor U1412 (N_1412,In_584,In_740);
nor U1413 (N_1413,In_1411,In_616);
nor U1414 (N_1414,In_740,In_739);
xnor U1415 (N_1415,In_591,In_1345);
xnor U1416 (N_1416,In_1078,In_1184);
or U1417 (N_1417,In_502,In_383);
or U1418 (N_1418,In_1044,In_1053);
nor U1419 (N_1419,In_133,In_1257);
xnor U1420 (N_1420,In_965,In_1147);
nor U1421 (N_1421,In_84,In_1219);
or U1422 (N_1422,In_684,In_122);
and U1423 (N_1423,In_1086,In_984);
and U1424 (N_1424,In_1094,In_289);
nand U1425 (N_1425,In_640,In_1433);
xor U1426 (N_1426,In_1232,In_964);
or U1427 (N_1427,In_985,In_686);
xor U1428 (N_1428,In_257,In_152);
nand U1429 (N_1429,In_864,In_1350);
nand U1430 (N_1430,In_1144,In_1407);
nand U1431 (N_1431,In_1323,In_1146);
nand U1432 (N_1432,In_228,In_830);
nand U1433 (N_1433,In_923,In_324);
xor U1434 (N_1434,In_750,In_38);
nor U1435 (N_1435,In_948,In_912);
nand U1436 (N_1436,In_775,In_988);
nor U1437 (N_1437,In_397,In_1235);
or U1438 (N_1438,In_112,In_131);
nor U1439 (N_1439,In_779,In_1334);
or U1440 (N_1440,In_1475,In_998);
nor U1441 (N_1441,In_923,In_556);
nor U1442 (N_1442,In_1020,In_884);
xnor U1443 (N_1443,In_1160,In_563);
xor U1444 (N_1444,In_549,In_1139);
and U1445 (N_1445,In_1486,In_1343);
nand U1446 (N_1446,In_465,In_258);
and U1447 (N_1447,In_909,In_284);
xor U1448 (N_1448,In_1291,In_159);
or U1449 (N_1449,In_661,In_313);
and U1450 (N_1450,In_694,In_1303);
and U1451 (N_1451,In_134,In_916);
nor U1452 (N_1452,In_561,In_1237);
or U1453 (N_1453,In_504,In_987);
nand U1454 (N_1454,In_148,In_913);
nand U1455 (N_1455,In_344,In_476);
nand U1456 (N_1456,In_1444,In_808);
xnor U1457 (N_1457,In_788,In_25);
or U1458 (N_1458,In_213,In_1435);
nor U1459 (N_1459,In_613,In_202);
xor U1460 (N_1460,In_1015,In_237);
or U1461 (N_1461,In_1373,In_1208);
xnor U1462 (N_1462,In_1391,In_859);
or U1463 (N_1463,In_545,In_912);
and U1464 (N_1464,In_4,In_244);
and U1465 (N_1465,In_842,In_459);
nor U1466 (N_1466,In_1455,In_389);
nor U1467 (N_1467,In_1267,In_1140);
and U1468 (N_1468,In_547,In_1118);
xor U1469 (N_1469,In_924,In_757);
nor U1470 (N_1470,In_18,In_144);
nor U1471 (N_1471,In_968,In_1481);
and U1472 (N_1472,In_479,In_1169);
nand U1473 (N_1473,In_384,In_1462);
or U1474 (N_1474,In_813,In_349);
and U1475 (N_1475,In_80,In_60);
xor U1476 (N_1476,In_1119,In_1061);
or U1477 (N_1477,In_335,In_246);
nor U1478 (N_1478,In_395,In_444);
and U1479 (N_1479,In_728,In_599);
nor U1480 (N_1480,In_1136,In_383);
nand U1481 (N_1481,In_434,In_1462);
nand U1482 (N_1482,In_1465,In_410);
nor U1483 (N_1483,In_846,In_668);
nor U1484 (N_1484,In_267,In_146);
xor U1485 (N_1485,In_808,In_525);
xor U1486 (N_1486,In_967,In_24);
or U1487 (N_1487,In_580,In_225);
or U1488 (N_1488,In_592,In_1090);
xor U1489 (N_1489,In_641,In_601);
and U1490 (N_1490,In_429,In_548);
nor U1491 (N_1491,In_559,In_513);
and U1492 (N_1492,In_910,In_848);
nand U1493 (N_1493,In_358,In_125);
xnor U1494 (N_1494,In_435,In_727);
or U1495 (N_1495,In_1095,In_469);
xnor U1496 (N_1496,In_1316,In_998);
nand U1497 (N_1497,In_91,In_132);
xnor U1498 (N_1498,In_779,In_489);
and U1499 (N_1499,In_230,In_740);
nor U1500 (N_1500,N_812,N_1283);
nor U1501 (N_1501,N_621,N_42);
nand U1502 (N_1502,N_321,N_1316);
nand U1503 (N_1503,N_233,N_91);
nand U1504 (N_1504,N_1108,N_1498);
or U1505 (N_1505,N_238,N_4);
xnor U1506 (N_1506,N_225,N_404);
and U1507 (N_1507,N_1299,N_873);
nand U1508 (N_1508,N_1155,N_582);
nand U1509 (N_1509,N_577,N_364);
nand U1510 (N_1510,N_242,N_656);
nand U1511 (N_1511,N_882,N_203);
nor U1512 (N_1512,N_1091,N_1219);
xnor U1513 (N_1513,N_672,N_849);
nand U1514 (N_1514,N_900,N_778);
xor U1515 (N_1515,N_425,N_810);
or U1516 (N_1516,N_1371,N_642);
and U1517 (N_1517,N_1111,N_886);
and U1518 (N_1518,N_909,N_85);
and U1519 (N_1519,N_832,N_107);
and U1520 (N_1520,N_1172,N_722);
or U1521 (N_1521,N_517,N_1246);
nand U1522 (N_1522,N_219,N_498);
and U1523 (N_1523,N_714,N_950);
nor U1524 (N_1524,N_735,N_349);
xnor U1525 (N_1525,N_1495,N_495);
xor U1526 (N_1526,N_317,N_727);
or U1527 (N_1527,N_1477,N_981);
or U1528 (N_1528,N_890,N_1337);
and U1529 (N_1529,N_790,N_633);
xnor U1530 (N_1530,N_261,N_913);
or U1531 (N_1531,N_1385,N_1405);
nand U1532 (N_1532,N_824,N_77);
nor U1533 (N_1533,N_96,N_991);
or U1534 (N_1534,N_1325,N_1416);
and U1535 (N_1535,N_465,N_1234);
nor U1536 (N_1536,N_246,N_165);
nand U1537 (N_1537,N_1414,N_827);
nor U1538 (N_1538,N_996,N_1201);
nand U1539 (N_1539,N_34,N_82);
nor U1540 (N_1540,N_130,N_965);
xnor U1541 (N_1541,N_247,N_744);
xor U1542 (N_1542,N_289,N_401);
nand U1543 (N_1543,N_1157,N_1376);
nand U1544 (N_1544,N_1315,N_576);
or U1545 (N_1545,N_745,N_754);
or U1546 (N_1546,N_603,N_431);
or U1547 (N_1547,N_1398,N_734);
nor U1548 (N_1548,N_454,N_354);
and U1549 (N_1549,N_1152,N_568);
nand U1550 (N_1550,N_1318,N_1209);
and U1551 (N_1551,N_210,N_1175);
and U1552 (N_1552,N_40,N_19);
xnor U1553 (N_1553,N_1436,N_804);
nor U1554 (N_1554,N_555,N_1286);
nor U1555 (N_1555,N_845,N_867);
xnor U1556 (N_1556,N_707,N_716);
xor U1557 (N_1557,N_836,N_559);
nor U1558 (N_1558,N_1482,N_750);
xor U1559 (N_1559,N_1424,N_102);
or U1560 (N_1560,N_264,N_1162);
nand U1561 (N_1561,N_976,N_774);
xor U1562 (N_1562,N_433,N_1378);
or U1563 (N_1563,N_999,N_1345);
nor U1564 (N_1564,N_1227,N_418);
xnor U1565 (N_1565,N_1443,N_604);
or U1566 (N_1566,N_762,N_295);
nand U1567 (N_1567,N_647,N_236);
nand U1568 (N_1568,N_1431,N_737);
and U1569 (N_1569,N_769,N_232);
xnor U1570 (N_1570,N_541,N_327);
nor U1571 (N_1571,N_973,N_554);
or U1572 (N_1572,N_1381,N_516);
nor U1573 (N_1573,N_114,N_1139);
and U1574 (N_1574,N_718,N_291);
nor U1575 (N_1575,N_86,N_789);
xor U1576 (N_1576,N_314,N_1429);
or U1577 (N_1577,N_1154,N_690);
and U1578 (N_1578,N_752,N_667);
or U1579 (N_1579,N_300,N_1188);
nor U1580 (N_1580,N_837,N_685);
xor U1581 (N_1581,N_635,N_1061);
nor U1582 (N_1582,N_518,N_383);
or U1583 (N_1583,N_910,N_221);
or U1584 (N_1584,N_413,N_1425);
nand U1585 (N_1585,N_103,N_1189);
and U1586 (N_1586,N_521,N_509);
and U1587 (N_1587,N_339,N_343);
nor U1588 (N_1588,N_319,N_1390);
nand U1589 (N_1589,N_1455,N_970);
xnor U1590 (N_1590,N_713,N_1094);
xnor U1591 (N_1591,N_985,N_1462);
and U1592 (N_1592,N_868,N_285);
nor U1593 (N_1593,N_522,N_1133);
and U1594 (N_1594,N_1043,N_1497);
and U1595 (N_1595,N_1044,N_1237);
or U1596 (N_1596,N_1314,N_1352);
xnor U1597 (N_1597,N_760,N_453);
and U1598 (N_1598,N_456,N_833);
xnor U1599 (N_1599,N_175,N_535);
or U1600 (N_1600,N_829,N_1338);
and U1601 (N_1601,N_263,N_893);
and U1602 (N_1602,N_871,N_993);
nand U1603 (N_1603,N_29,N_583);
nand U1604 (N_1604,N_1127,N_1257);
and U1605 (N_1605,N_1469,N_146);
nor U1606 (N_1606,N_705,N_170);
or U1607 (N_1607,N_208,N_990);
xnor U1608 (N_1608,N_783,N_1432);
nand U1609 (N_1609,N_741,N_1271);
nand U1610 (N_1610,N_422,N_1323);
nor U1611 (N_1611,N_1202,N_126);
and U1612 (N_1612,N_174,N_703);
nand U1613 (N_1613,N_791,N_375);
xor U1614 (N_1614,N_255,N_1496);
and U1615 (N_1615,N_308,N_350);
xor U1616 (N_1616,N_792,N_207);
nand U1617 (N_1617,N_780,N_20);
nand U1618 (N_1618,N_90,N_854);
xor U1619 (N_1619,N_883,N_1366);
xnor U1620 (N_1620,N_200,N_65);
nand U1621 (N_1621,N_698,N_220);
xor U1622 (N_1622,N_1480,N_630);
nor U1623 (N_1623,N_117,N_1187);
or U1624 (N_1624,N_270,N_158);
nand U1625 (N_1625,N_1153,N_1330);
or U1626 (N_1626,N_793,N_898);
and U1627 (N_1627,N_556,N_1302);
xnor U1628 (N_1628,N_537,N_1456);
and U1629 (N_1629,N_1000,N_1065);
nand U1630 (N_1630,N_768,N_588);
xnor U1631 (N_1631,N_527,N_811);
nor U1632 (N_1632,N_52,N_275);
nand U1633 (N_1633,N_1274,N_58);
xor U1634 (N_1634,N_963,N_99);
nand U1635 (N_1635,N_1067,N_193);
xnor U1636 (N_1636,N_187,N_294);
and U1637 (N_1637,N_104,N_212);
xnor U1638 (N_1638,N_412,N_695);
or U1639 (N_1639,N_391,N_466);
xor U1640 (N_1640,N_427,N_875);
xor U1641 (N_1641,N_245,N_21);
xor U1642 (N_1642,N_1356,N_1453);
and U1643 (N_1643,N_1,N_13);
xor U1644 (N_1644,N_69,N_551);
and U1645 (N_1645,N_755,N_1001);
and U1646 (N_1646,N_310,N_277);
nor U1647 (N_1647,N_1132,N_1053);
and U1648 (N_1648,N_1342,N_926);
xor U1649 (N_1649,N_402,N_371);
or U1650 (N_1650,N_906,N_670);
xor U1651 (N_1651,N_1074,N_562);
nand U1652 (N_1652,N_1308,N_1492);
xor U1653 (N_1653,N_72,N_1420);
xor U1654 (N_1654,N_743,N_338);
or U1655 (N_1655,N_489,N_60);
nand U1656 (N_1656,N_1472,N_17);
nor U1657 (N_1657,N_335,N_533);
or U1658 (N_1658,N_152,N_631);
nor U1659 (N_1659,N_507,N_488);
xnor U1660 (N_1660,N_947,N_814);
xor U1661 (N_1661,N_194,N_896);
and U1662 (N_1662,N_885,N_997);
or U1663 (N_1663,N_988,N_70);
nor U1664 (N_1664,N_140,N_198);
and U1665 (N_1665,N_22,N_946);
nor U1666 (N_1666,N_346,N_729);
xor U1667 (N_1667,N_1300,N_680);
or U1668 (N_1668,N_1106,N_474);
xnor U1669 (N_1669,N_1276,N_566);
xnor U1670 (N_1670,N_1313,N_600);
or U1671 (N_1671,N_962,N_1236);
nor U1672 (N_1672,N_1422,N_110);
nor U1673 (N_1673,N_891,N_403);
or U1674 (N_1674,N_1176,N_197);
nor U1675 (N_1675,N_733,N_1251);
nand U1676 (N_1676,N_968,N_505);
and U1677 (N_1677,N_1489,N_76);
and U1678 (N_1678,N_185,N_1012);
or U1679 (N_1679,N_434,N_405);
xor U1680 (N_1680,N_1401,N_108);
or U1681 (N_1681,N_464,N_856);
xnor U1682 (N_1682,N_1297,N_1129);
xnor U1683 (N_1683,N_749,N_953);
or U1684 (N_1684,N_1451,N_312);
xnor U1685 (N_1685,N_468,N_1089);
and U1686 (N_1686,N_37,N_1428);
or U1687 (N_1687,N_919,N_1081);
nor U1688 (N_1688,N_437,N_131);
nor U1689 (N_1689,N_1193,N_663);
nor U1690 (N_1690,N_877,N_1470);
or U1691 (N_1691,N_715,N_282);
nand U1692 (N_1692,N_747,N_842);
nor U1693 (N_1693,N_138,N_662);
nand U1694 (N_1694,N_1389,N_1124);
or U1695 (N_1695,N_874,N_959);
xnor U1696 (N_1696,N_213,N_1367);
and U1697 (N_1697,N_1118,N_664);
nand U1698 (N_1698,N_572,N_884);
and U1699 (N_1699,N_540,N_98);
nor U1700 (N_1700,N_1382,N_441);
and U1701 (N_1701,N_11,N_1082);
or U1702 (N_1702,N_1364,N_803);
nand U1703 (N_1703,N_356,N_1442);
and U1704 (N_1704,N_846,N_1161);
nand U1705 (N_1705,N_513,N_1262);
nand U1706 (N_1706,N_111,N_591);
nor U1707 (N_1707,N_1407,N_1023);
nor U1708 (N_1708,N_1284,N_1239);
nor U1709 (N_1709,N_315,N_1281);
or U1710 (N_1710,N_799,N_1100);
xor U1711 (N_1711,N_1450,N_452);
nand U1712 (N_1712,N_1441,N_659);
nor U1713 (N_1713,N_1384,N_1215);
xor U1714 (N_1714,N_1164,N_665);
or U1715 (N_1715,N_843,N_616);
or U1716 (N_1716,N_153,N_1034);
or U1717 (N_1717,N_1038,N_660);
nand U1718 (N_1718,N_530,N_492);
nand U1719 (N_1719,N_1329,N_515);
nand U1720 (N_1720,N_237,N_243);
nor U1721 (N_1721,N_178,N_206);
nor U1722 (N_1722,N_368,N_655);
nor U1723 (N_1723,N_945,N_396);
xnor U1724 (N_1724,N_1213,N_1322);
or U1725 (N_1725,N_611,N_305);
and U1726 (N_1726,N_1458,N_1024);
nor U1727 (N_1727,N_1258,N_48);
nand U1728 (N_1728,N_1319,N_1208);
nor U1729 (N_1729,N_1479,N_798);
or U1730 (N_1730,N_1404,N_267);
or U1731 (N_1731,N_1008,N_1460);
and U1732 (N_1732,N_381,N_164);
xnor U1733 (N_1733,N_917,N_1334);
or U1734 (N_1734,N_190,N_1064);
or U1735 (N_1735,N_1349,N_1230);
or U1736 (N_1736,N_880,N_1007);
nand U1737 (N_1737,N_486,N_565);
nand U1738 (N_1738,N_1263,N_1475);
or U1739 (N_1739,N_124,N_142);
and U1740 (N_1740,N_1104,N_936);
xnor U1741 (N_1741,N_1415,N_1266);
nor U1742 (N_1742,N_306,N_1412);
xnor U1743 (N_1743,N_16,N_1174);
nor U1744 (N_1744,N_504,N_64);
or U1745 (N_1745,N_794,N_362);
xnor U1746 (N_1746,N_1306,N_378);
or U1747 (N_1747,N_1282,N_348);
and U1748 (N_1748,N_1427,N_1397);
nand U1749 (N_1749,N_1071,N_942);
nor U1750 (N_1750,N_95,N_1224);
nor U1751 (N_1751,N_1392,N_1273);
and U1752 (N_1752,N_15,N_1015);
nor U1753 (N_1753,N_1092,N_1052);
nor U1754 (N_1754,N_937,N_423);
xnor U1755 (N_1755,N_202,N_866);
nand U1756 (N_1756,N_809,N_392);
nand U1757 (N_1757,N_365,N_525);
nor U1758 (N_1758,N_214,N_1070);
and U1759 (N_1759,N_1212,N_217);
and U1760 (N_1760,N_1418,N_1448);
or U1761 (N_1761,N_644,N_84);
nand U1762 (N_1762,N_157,N_948);
and U1763 (N_1763,N_216,N_1093);
nor U1764 (N_1764,N_252,N_1003);
nand U1765 (N_1765,N_757,N_523);
xor U1766 (N_1766,N_748,N_271);
nand U1767 (N_1767,N_372,N_864);
or U1768 (N_1768,N_1056,N_544);
nand U1769 (N_1769,N_1370,N_341);
nand U1770 (N_1770,N_440,N_445);
and U1771 (N_1771,N_8,N_825);
nand U1772 (N_1772,N_1168,N_122);
nor U1773 (N_1773,N_1149,N_320);
and U1774 (N_1774,N_929,N_1310);
xor U1775 (N_1775,N_26,N_123);
nor U1776 (N_1776,N_696,N_1240);
or U1777 (N_1777,N_708,N_921);
and U1778 (N_1778,N_691,N_439);
or U1779 (N_1779,N_732,N_1333);
and U1780 (N_1780,N_1254,N_1085);
nand U1781 (N_1781,N_46,N_66);
and U1782 (N_1782,N_1447,N_1303);
or U1783 (N_1783,N_361,N_476);
nor U1784 (N_1784,N_668,N_1032);
nor U1785 (N_1785,N_738,N_987);
or U1786 (N_1786,N_419,N_834);
or U1787 (N_1787,N_905,N_595);
and U1788 (N_1788,N_1320,N_1090);
nand U1789 (N_1789,N_1046,N_719);
and U1790 (N_1790,N_746,N_1332);
or U1791 (N_1791,N_1277,N_395);
nor U1792 (N_1792,N_45,N_940);
or U1793 (N_1793,N_415,N_390);
nand U1794 (N_1794,N_1137,N_977);
xor U1795 (N_1795,N_380,N_761);
nor U1796 (N_1796,N_939,N_932);
and U1797 (N_1797,N_1244,N_795);
and U1798 (N_1798,N_673,N_1343);
xnor U1799 (N_1799,N_304,N_785);
nand U1800 (N_1800,N_370,N_1249);
nor U1801 (N_1801,N_1114,N_87);
or U1802 (N_1802,N_307,N_181);
nor U1803 (N_1803,N_1204,N_1413);
nand U1804 (N_1804,N_358,N_1134);
nand U1805 (N_1805,N_589,N_287);
and U1806 (N_1806,N_1233,N_1446);
and U1807 (N_1807,N_487,N_927);
nor U1808 (N_1808,N_624,N_1260);
xor U1809 (N_1809,N_1068,N_618);
nor U1810 (N_1810,N_1275,N_1242);
xor U1811 (N_1811,N_477,N_420);
nand U1812 (N_1812,N_1079,N_1148);
nor U1813 (N_1813,N_918,N_676);
nor U1814 (N_1814,N_1280,N_742);
or U1815 (N_1815,N_966,N_25);
nor U1816 (N_1816,N_1047,N_764);
or U1817 (N_1817,N_463,N_325);
and U1818 (N_1818,N_648,N_771);
xor U1819 (N_1819,N_775,N_32);
or U1820 (N_1820,N_1055,N_897);
and U1821 (N_1821,N_851,N_914);
or U1822 (N_1822,N_44,N_83);
or U1823 (N_1823,N_1099,N_168);
nor U1824 (N_1824,N_1130,N_112);
or U1825 (N_1825,N_1101,N_546);
nand U1826 (N_1826,N_1088,N_1484);
or U1827 (N_1827,N_351,N_134);
nand U1828 (N_1828,N_377,N_539);
xnor U1829 (N_1829,N_1380,N_1021);
nor U1830 (N_1830,N_1169,N_1011);
or U1831 (N_1831,N_710,N_192);
xnor U1832 (N_1832,N_593,N_1395);
nand U1833 (N_1833,N_272,N_1494);
nand U1834 (N_1834,N_1438,N_278);
or U1835 (N_1835,N_1362,N_93);
or U1836 (N_1836,N_532,N_1080);
or U1837 (N_1837,N_257,N_887);
xor U1838 (N_1838,N_1406,N_1221);
or U1839 (N_1839,N_435,N_643);
and U1840 (N_1840,N_81,N_1028);
or U1841 (N_1841,N_78,N_1009);
nand U1842 (N_1842,N_328,N_855);
nor U1843 (N_1843,N_596,N_1105);
and U1844 (N_1844,N_55,N_1336);
nand U1845 (N_1845,N_998,N_309);
or U1846 (N_1846,N_958,N_39);
and U1847 (N_1847,N_788,N_1321);
nor U1848 (N_1848,N_1177,N_979);
nor U1849 (N_1849,N_215,N_1151);
nor U1850 (N_1850,N_974,N_1487);
or U1851 (N_1851,N_1347,N_18);
nand U1852 (N_1852,N_1186,N_410);
nor U1853 (N_1853,N_485,N_961);
nand U1854 (N_1854,N_1304,N_201);
or U1855 (N_1855,N_1490,N_276);
or U1856 (N_1856,N_903,N_286);
and U1857 (N_1857,N_177,N_3);
nand U1858 (N_1858,N_1459,N_183);
nor U1859 (N_1859,N_1445,N_1307);
and U1860 (N_1860,N_1020,N_564);
and U1861 (N_1861,N_520,N_1241);
xor U1862 (N_1862,N_671,N_558);
nor U1863 (N_1863,N_901,N_1040);
nor U1864 (N_1864,N_571,N_1434);
and U1865 (N_1865,N_209,N_645);
and U1866 (N_1866,N_1409,N_1294);
nand U1867 (N_1867,N_189,N_1223);
or U1868 (N_1868,N_188,N_249);
or U1869 (N_1869,N_222,N_136);
or U1870 (N_1870,N_916,N_1196);
or U1871 (N_1871,N_53,N_911);
nand U1872 (N_1872,N_367,N_1076);
and U1873 (N_1873,N_751,N_273);
or U1874 (N_1874,N_759,N_169);
or U1875 (N_1875,N_613,N_557);
nand U1876 (N_1876,N_1373,N_574);
and U1877 (N_1877,N_137,N_928);
or U1878 (N_1878,N_145,N_704);
and U1879 (N_1879,N_1377,N_1194);
and U1880 (N_1880,N_167,N_241);
nand U1881 (N_1881,N_1268,N_865);
and U1882 (N_1882,N_720,N_1493);
xor U1883 (N_1883,N_1060,N_1440);
nand U1884 (N_1884,N_199,N_1125);
or U1885 (N_1885,N_1433,N_1402);
xnor U1886 (N_1886,N_61,N_89);
and U1887 (N_1887,N_560,N_382);
nor U1888 (N_1888,N_1195,N_1051);
or U1889 (N_1889,N_679,N_826);
nand U1890 (N_1890,N_781,N_975);
and U1891 (N_1891,N_1050,N_838);
and U1892 (N_1892,N_1305,N_610);
nor U1893 (N_1893,N_1328,N_924);
nor U1894 (N_1894,N_1348,N_1435);
or U1895 (N_1895,N_290,N_711);
and U1896 (N_1896,N_684,N_800);
and U1897 (N_1897,N_620,N_994);
nor U1898 (N_1898,N_1030,N_1063);
and U1899 (N_1899,N_1243,N_1339);
xnor U1900 (N_1900,N_756,N_779);
nor U1901 (N_1901,N_652,N_1340);
nor U1902 (N_1902,N_43,N_311);
xnor U1903 (N_1903,N_426,N_248);
nand U1904 (N_1904,N_231,N_347);
xnor U1905 (N_1905,N_863,N_649);
xnor U1906 (N_1906,N_1278,N_56);
nor U1907 (N_1907,N_862,N_360);
and U1908 (N_1908,N_374,N_949);
nor U1909 (N_1909,N_359,N_511);
xor U1910 (N_1910,N_739,N_943);
nand U1911 (N_1911,N_389,N_260);
nand U1912 (N_1912,N_859,N_1110);
or U1913 (N_1913,N_776,N_819);
or U1914 (N_1914,N_497,N_1410);
xnor U1915 (N_1915,N_1259,N_524);
xnor U1916 (N_1916,N_472,N_584);
xnor U1917 (N_1917,N_268,N_443);
xnor U1918 (N_1918,N_1374,N_1182);
nor U1919 (N_1919,N_561,N_1238);
xnor U1920 (N_1920,N_989,N_254);
or U1921 (N_1921,N_501,N_1466);
or U1922 (N_1922,N_702,N_133);
nand U1923 (N_1923,N_796,N_384);
and U1924 (N_1924,N_960,N_284);
xnor U1925 (N_1925,N_1086,N_1452);
and U1926 (N_1926,N_969,N_1031);
or U1927 (N_1927,N_575,N_1073);
and U1928 (N_1928,N_1017,N_606);
xnor U1929 (N_1929,N_409,N_545);
nand U1930 (N_1930,N_770,N_258);
and U1931 (N_1931,N_677,N_797);
and U1932 (N_1932,N_1203,N_447);
nand U1933 (N_1933,N_1383,N_653);
nor U1934 (N_1934,N_369,N_1198);
nand U1935 (N_1935,N_62,N_387);
xor U1936 (N_1936,N_33,N_1478);
xnor U1937 (N_1937,N_324,N_1476);
xor U1938 (N_1938,N_1312,N_68);
and U1939 (N_1939,N_160,N_787);
or U1940 (N_1940,N_92,N_609);
and U1941 (N_1941,N_262,N_1059);
nor U1942 (N_1942,N_97,N_646);
nand U1943 (N_1943,N_1199,N_478);
or U1944 (N_1944,N_196,N_666);
xnor U1945 (N_1945,N_101,N_1454);
nand U1946 (N_1946,N_329,N_28);
nand U1947 (N_1947,N_1045,N_1317);
or U1948 (N_1948,N_1181,N_1128);
or U1949 (N_1949,N_469,N_1368);
xnor U1950 (N_1950,N_38,N_1361);
nor U1951 (N_1951,N_470,N_129);
and U1952 (N_1952,N_528,N_1004);
xnor U1953 (N_1953,N_1235,N_920);
nand U1954 (N_1954,N_1375,N_817);
nor U1955 (N_1955,N_514,N_1115);
and U1956 (N_1956,N_550,N_573);
and U1957 (N_1957,N_166,N_784);
xor U1958 (N_1958,N_406,N_480);
nor U1959 (N_1959,N_923,N_964);
xnor U1960 (N_1960,N_602,N_1210);
or U1961 (N_1961,N_935,N_597);
and U1962 (N_1962,N_581,N_1341);
xor U1963 (N_1963,N_471,N_1077);
and U1964 (N_1964,N_491,N_23);
nand U1965 (N_1965,N_1192,N_1288);
and U1966 (N_1966,N_227,N_414);
nor U1967 (N_1967,N_1184,N_1491);
nand U1968 (N_1968,N_204,N_502);
and U1969 (N_1969,N_128,N_281);
or U1970 (N_1970,N_1036,N_661);
and U1971 (N_1971,N_179,N_899);
or U1972 (N_1972,N_113,N_1261);
nor U1973 (N_1973,N_1481,N_1013);
xnor U1974 (N_1974,N_1103,N_161);
xor U1975 (N_1975,N_1386,N_952);
xnor U1976 (N_1976,N_1353,N_1075);
xor U1977 (N_1977,N_1167,N_482);
and U1978 (N_1978,N_508,N_144);
or U1979 (N_1979,N_697,N_579);
nor U1980 (N_1980,N_205,N_1301);
nor U1981 (N_1981,N_637,N_63);
nand U1982 (N_1982,N_1387,N_1138);
xor U1983 (N_1983,N_1245,N_363);
xnor U1984 (N_1984,N_5,N_1488);
nand U1985 (N_1985,N_625,N_411);
and U1986 (N_1986,N_398,N_24);
and U1987 (N_1987,N_416,N_1109);
nor U1988 (N_1988,N_1107,N_1159);
nor U1989 (N_1989,N_318,N_1078);
and U1990 (N_1990,N_326,N_683);
and U1991 (N_1991,N_978,N_1019);
xnor U1992 (N_1992,N_570,N_869);
nand U1993 (N_1993,N_563,N_569);
nand U1994 (N_1994,N_176,N_1256);
nor U1995 (N_1995,N_1026,N_908);
and U1996 (N_1996,N_1253,N_1423);
nor U1997 (N_1997,N_590,N_462);
and U1998 (N_1998,N_458,N_585);
or U1999 (N_1999,N_1474,N_983);
nand U2000 (N_2000,N_640,N_27);
and U2001 (N_2001,N_682,N_878);
xnor U2002 (N_2002,N_116,N_1359);
or U2003 (N_2003,N_500,N_725);
nor U2004 (N_2004,N_650,N_186);
nand U2005 (N_2005,N_706,N_1014);
nand U2006 (N_2006,N_1123,N_345);
xor U2007 (N_2007,N_1369,N_1449);
nor U2008 (N_2008,N_408,N_1358);
or U2009 (N_2009,N_847,N_1140);
xor U2010 (N_2010,N_951,N_694);
and U2011 (N_2011,N_74,N_1272);
and U2012 (N_2012,N_279,N_429);
and U2013 (N_2013,N_322,N_1267);
nand U2014 (N_2014,N_740,N_1354);
nand U2015 (N_2015,N_1145,N_844);
and U2016 (N_2016,N_230,N_617);
nor U2017 (N_2017,N_1394,N_758);
and U2018 (N_2018,N_1185,N_155);
and U2019 (N_2019,N_1190,N_956);
nor U2020 (N_2020,N_1135,N_1486);
nor U2021 (N_2021,N_1005,N_1269);
nor U2022 (N_2022,N_266,N_31);
or U2023 (N_2023,N_228,N_1197);
nand U2024 (N_2024,N_280,N_1265);
nor U2025 (N_2025,N_1010,N_678);
xnor U2026 (N_2026,N_73,N_1039);
or U2027 (N_2027,N_1158,N_150);
or U2028 (N_2028,N_1116,N_805);
xor U2029 (N_2029,N_552,N_432);
nor U2030 (N_2030,N_506,N_1326);
or U2031 (N_2031,N_688,N_1057);
xor U2032 (N_2032,N_211,N_438);
nor U2033 (N_2033,N_1298,N_881);
nand U2034 (N_2034,N_1363,N_587);
and U2035 (N_2035,N_293,N_709);
xnor U2036 (N_2036,N_36,N_902);
nand U2037 (N_2037,N_858,N_954);
or U2038 (N_2038,N_930,N_182);
nand U2039 (N_2039,N_1220,N_115);
nor U2040 (N_2040,N_30,N_352);
nand U2041 (N_2041,N_1002,N_54);
xnor U2042 (N_2042,N_451,N_1098);
nor U2043 (N_2043,N_1121,N_1006);
and U2044 (N_2044,N_479,N_475);
and U2045 (N_2045,N_1218,N_657);
or U2046 (N_2046,N_344,N_995);
or U2047 (N_2047,N_407,N_461);
nor U2048 (N_2048,N_634,N_1165);
or U2049 (N_2049,N_444,N_728);
or U2050 (N_2050,N_786,N_283);
nor U2051 (N_2051,N_1357,N_1411);
xor U2052 (N_2052,N_481,N_1344);
nor U2053 (N_2053,N_376,N_9);
or U2054 (N_2054,N_173,N_6);
or U2055 (N_2055,N_1296,N_980);
or U2056 (N_2056,N_1084,N_712);
nand U2057 (N_2057,N_1166,N_578);
or U2058 (N_2058,N_417,N_689);
nor U2059 (N_2059,N_623,N_1285);
and U2060 (N_2060,N_1250,N_156);
or U2061 (N_2061,N_125,N_1225);
and U2062 (N_2062,N_421,N_536);
nand U2063 (N_2063,N_1066,N_542);
nor U2064 (N_2064,N_436,N_357);
nor U2065 (N_2065,N_1171,N_143);
nor U2066 (N_2066,N_355,N_674);
or U2067 (N_2067,N_490,N_14);
xor U2068 (N_2068,N_1292,N_636);
and U2069 (N_2069,N_1464,N_332);
or U2070 (N_2070,N_483,N_1437);
nor U2071 (N_2071,N_828,N_331);
nand U2072 (N_2072,N_118,N_1264);
xnor U2073 (N_2073,N_1200,N_724);
and U2074 (N_2074,N_473,N_1444);
or U2075 (N_2075,N_681,N_904);
nor U2076 (N_2076,N_388,N_457);
nand U2077 (N_2077,N_1141,N_1391);
nand U2078 (N_2078,N_1327,N_298);
or U2079 (N_2079,N_79,N_1016);
xnor U2080 (N_2080,N_967,N_1179);
nor U2081 (N_2081,N_822,N_109);
nor U2082 (N_2082,N_531,N_340);
nor U2083 (N_2083,N_1231,N_1205);
nand U2084 (N_2084,N_269,N_47);
xor U2085 (N_2085,N_1170,N_1287);
nand U2086 (N_2086,N_1350,N_669);
nor U2087 (N_2087,N_323,N_184);
nand U2088 (N_2088,N_1035,N_373);
nand U2089 (N_2089,N_753,N_41);
xnor U2090 (N_2090,N_1102,N_857);
nor U2091 (N_2091,N_627,N_922);
nand U2092 (N_2092,N_693,N_1120);
nor U2093 (N_2093,N_915,N_1247);
nand U2094 (N_2094,N_1360,N_818);
nor U2095 (N_2095,N_195,N_608);
nor U2096 (N_2096,N_1083,N_1467);
nand U2097 (N_2097,N_801,N_895);
or U2098 (N_2098,N_580,N_1222);
xnor U2099 (N_2099,N_639,N_229);
or U2100 (N_2100,N_159,N_105);
or U2101 (N_2101,N_1346,N_397);
nand U2102 (N_2102,N_393,N_1037);
nor U2103 (N_2103,N_1029,N_75);
or U2104 (N_2104,N_723,N_547);
nor U2105 (N_2105,N_615,N_88);
nand U2106 (N_2106,N_529,N_1049);
nand U2107 (N_2107,N_773,N_235);
and U2108 (N_2108,N_592,N_336);
xor U2109 (N_2109,N_629,N_1122);
nor U2110 (N_2110,N_1062,N_821);
xnor U2111 (N_2111,N_180,N_638);
nand U2112 (N_2112,N_605,N_288);
nand U2113 (N_2113,N_1087,N_944);
or U2114 (N_2114,N_984,N_467);
nand U2115 (N_2115,N_1097,N_1072);
and U2116 (N_2116,N_850,N_0);
and U2117 (N_2117,N_1293,N_459);
nand U2118 (N_2118,N_1335,N_1144);
and U2119 (N_2119,N_1207,N_687);
or U2120 (N_2120,N_1408,N_807);
or U2121 (N_2121,N_1041,N_1471);
nand U2122 (N_2122,N_1146,N_274);
or U2123 (N_2123,N_619,N_982);
nor U2124 (N_2124,N_1160,N_1142);
and U2125 (N_2125,N_839,N_424);
nand U2126 (N_2126,N_35,N_1499);
nand U2127 (N_2127,N_148,N_171);
nor U2128 (N_2128,N_399,N_1355);
nand U2129 (N_2129,N_50,N_1289);
and U2130 (N_2130,N_553,N_256);
and U2131 (N_2131,N_1150,N_815);
or U2132 (N_2132,N_594,N_806);
nor U2133 (N_2133,N_912,N_632);
or U2134 (N_2134,N_612,N_777);
nand U2135 (N_2135,N_1217,N_1485);
nand U2136 (N_2136,N_955,N_925);
or U2137 (N_2137,N_303,N_450);
nand U2138 (N_2138,N_654,N_934);
nand U2139 (N_2139,N_840,N_628);
and U2140 (N_2140,N_549,N_586);
and U2141 (N_2141,N_59,N_626);
xor U2142 (N_2142,N_1463,N_316);
nand U2143 (N_2143,N_333,N_599);
xor U2144 (N_2144,N_894,N_299);
nand U2145 (N_2145,N_567,N_510);
nor U2146 (N_2146,N_730,N_622);
and U2147 (N_2147,N_1180,N_1211);
xor U2148 (N_2148,N_933,N_296);
and U2149 (N_2149,N_394,N_446);
nor U2150 (N_2150,N_223,N_1372);
nand U2151 (N_2151,N_218,N_1119);
and U2152 (N_2152,N_12,N_1252);
or U2153 (N_2153,N_699,N_1379);
nor U2154 (N_2154,N_240,N_151);
nor U2155 (N_2155,N_139,N_512);
xor U2156 (N_2156,N_1226,N_1156);
and U2157 (N_2157,N_163,N_460);
xor U2158 (N_2158,N_841,N_860);
and U2159 (N_2159,N_1255,N_692);
or U2160 (N_2160,N_938,N_763);
and U2161 (N_2161,N_302,N_1095);
xnor U2162 (N_2162,N_1403,N_265);
nand U2163 (N_2163,N_701,N_1178);
xor U2164 (N_2164,N_1112,N_1473);
xor U2165 (N_2165,N_700,N_1291);
and U2166 (N_2166,N_870,N_71);
or U2167 (N_2167,N_848,N_1270);
xnor U2168 (N_2168,N_675,N_251);
and U2169 (N_2169,N_931,N_548);
nor U2170 (N_2170,N_7,N_1295);
xor U2171 (N_2171,N_1468,N_1430);
or U2172 (N_2172,N_889,N_1042);
and U2173 (N_2173,N_876,N_986);
and U2174 (N_2174,N_1228,N_337);
xnor U2175 (N_2175,N_766,N_686);
and U2176 (N_2176,N_499,N_853);
and U2177 (N_2177,N_721,N_802);
xnor U2178 (N_2178,N_538,N_641);
and U2179 (N_2179,N_1465,N_301);
xor U2180 (N_2180,N_1173,N_292);
nand U2181 (N_2181,N_1290,N_1393);
or U2182 (N_2182,N_1279,N_234);
xnor U2183 (N_2183,N_1419,N_244);
nand U2184 (N_2184,N_385,N_1022);
and U2185 (N_2185,N_651,N_1421);
nand U2186 (N_2186,N_1033,N_601);
nor U2187 (N_2187,N_484,N_49);
or U2188 (N_2188,N_149,N_141);
nor U2189 (N_2189,N_1417,N_226);
and U2190 (N_2190,N_813,N_1054);
nor U2191 (N_2191,N_162,N_57);
or U2192 (N_2192,N_428,N_1483);
xnor U2193 (N_2193,N_1113,N_259);
nand U2194 (N_2194,N_736,N_493);
nand U2195 (N_2195,N_253,N_154);
or U2196 (N_2196,N_879,N_51);
nand U2197 (N_2197,N_132,N_1439);
xor U2198 (N_2198,N_820,N_503);
xor U2199 (N_2199,N_1229,N_106);
or U2200 (N_2200,N_120,N_830);
and U2201 (N_2201,N_67,N_534);
and U2202 (N_2202,N_831,N_861);
xnor U2203 (N_2203,N_607,N_250);
and U2204 (N_2204,N_494,N_1331);
nand U2205 (N_2205,N_808,N_1131);
nor U2206 (N_2206,N_400,N_366);
or U2207 (N_2207,N_2,N_330);
or U2208 (N_2208,N_888,N_971);
nor U2209 (N_2209,N_100,N_386);
nor U2210 (N_2210,N_823,N_1309);
or U2211 (N_2211,N_658,N_430);
xnor U2212 (N_2212,N_1216,N_1311);
and U2213 (N_2213,N_772,N_816);
xor U2214 (N_2214,N_614,N_1351);
and U2215 (N_2215,N_1126,N_313);
and U2216 (N_2216,N_1399,N_835);
and U2217 (N_2217,N_147,N_1136);
nand U2218 (N_2218,N_765,N_767);
or U2219 (N_2219,N_442,N_941);
nand U2220 (N_2220,N_1025,N_1232);
nand U2221 (N_2221,N_957,N_726);
and U2222 (N_2222,N_1191,N_1147);
xor U2223 (N_2223,N_892,N_334);
nand U2224 (N_2224,N_80,N_342);
or U2225 (N_2225,N_1388,N_717);
nor U2226 (N_2226,N_1143,N_1457);
xnor U2227 (N_2227,N_94,N_496);
xnor U2228 (N_2228,N_449,N_1069);
and U2229 (N_2229,N_992,N_172);
xor U2230 (N_2230,N_1400,N_135);
nor U2231 (N_2231,N_239,N_1183);
nor U2232 (N_2232,N_119,N_1365);
or U2233 (N_2233,N_1117,N_1214);
nor U2234 (N_2234,N_448,N_598);
xor U2235 (N_2235,N_1248,N_1324);
xor U2236 (N_2236,N_907,N_1018);
nor U2237 (N_2237,N_1027,N_526);
nor U2238 (N_2238,N_10,N_1461);
nor U2239 (N_2239,N_127,N_379);
or U2240 (N_2240,N_121,N_1426);
nor U2241 (N_2241,N_353,N_782);
nor U2242 (N_2242,N_543,N_519);
xor U2243 (N_2243,N_1163,N_872);
and U2244 (N_2244,N_852,N_297);
nor U2245 (N_2245,N_972,N_1396);
nand U2246 (N_2246,N_1058,N_1206);
nor U2247 (N_2247,N_224,N_731);
xor U2248 (N_2248,N_1096,N_1048);
or U2249 (N_2249,N_455,N_191);
xor U2250 (N_2250,N_1050,N_1347);
nor U2251 (N_2251,N_698,N_165);
xor U2252 (N_2252,N_621,N_1219);
nand U2253 (N_2253,N_455,N_405);
xor U2254 (N_2254,N_397,N_329);
and U2255 (N_2255,N_1285,N_1381);
xnor U2256 (N_2256,N_630,N_273);
xor U2257 (N_2257,N_286,N_818);
xor U2258 (N_2258,N_173,N_1224);
nand U2259 (N_2259,N_1212,N_397);
nor U2260 (N_2260,N_1468,N_1380);
and U2261 (N_2261,N_118,N_95);
nand U2262 (N_2262,N_1002,N_855);
nor U2263 (N_2263,N_317,N_209);
nor U2264 (N_2264,N_952,N_809);
xor U2265 (N_2265,N_1020,N_592);
or U2266 (N_2266,N_133,N_1382);
and U2267 (N_2267,N_30,N_650);
nand U2268 (N_2268,N_1216,N_440);
and U2269 (N_2269,N_361,N_513);
nand U2270 (N_2270,N_1478,N_822);
or U2271 (N_2271,N_671,N_342);
xor U2272 (N_2272,N_139,N_1259);
xnor U2273 (N_2273,N_800,N_1380);
and U2274 (N_2274,N_962,N_794);
or U2275 (N_2275,N_140,N_344);
xor U2276 (N_2276,N_347,N_469);
or U2277 (N_2277,N_876,N_157);
and U2278 (N_2278,N_1336,N_568);
and U2279 (N_2279,N_1227,N_299);
nand U2280 (N_2280,N_121,N_67);
xor U2281 (N_2281,N_1383,N_407);
xnor U2282 (N_2282,N_891,N_215);
or U2283 (N_2283,N_121,N_1352);
xnor U2284 (N_2284,N_115,N_784);
xor U2285 (N_2285,N_686,N_252);
xnor U2286 (N_2286,N_703,N_504);
xnor U2287 (N_2287,N_748,N_437);
xor U2288 (N_2288,N_364,N_1090);
and U2289 (N_2289,N_173,N_585);
nand U2290 (N_2290,N_947,N_1399);
or U2291 (N_2291,N_256,N_504);
and U2292 (N_2292,N_1413,N_1042);
or U2293 (N_2293,N_994,N_665);
xor U2294 (N_2294,N_463,N_1315);
xor U2295 (N_2295,N_1236,N_231);
xor U2296 (N_2296,N_2,N_739);
and U2297 (N_2297,N_103,N_1164);
or U2298 (N_2298,N_456,N_1449);
nor U2299 (N_2299,N_1012,N_1428);
and U2300 (N_2300,N_1015,N_218);
or U2301 (N_2301,N_1289,N_1283);
and U2302 (N_2302,N_1437,N_670);
xor U2303 (N_2303,N_1437,N_1010);
nor U2304 (N_2304,N_1094,N_883);
xnor U2305 (N_2305,N_184,N_1070);
nand U2306 (N_2306,N_760,N_560);
xnor U2307 (N_2307,N_479,N_710);
or U2308 (N_2308,N_881,N_1449);
or U2309 (N_2309,N_850,N_543);
or U2310 (N_2310,N_360,N_524);
or U2311 (N_2311,N_115,N_1088);
or U2312 (N_2312,N_217,N_782);
nor U2313 (N_2313,N_795,N_353);
nor U2314 (N_2314,N_566,N_480);
and U2315 (N_2315,N_1369,N_32);
and U2316 (N_2316,N_613,N_61);
xnor U2317 (N_2317,N_1189,N_887);
nand U2318 (N_2318,N_1225,N_264);
nand U2319 (N_2319,N_1299,N_1245);
or U2320 (N_2320,N_1091,N_178);
or U2321 (N_2321,N_128,N_810);
and U2322 (N_2322,N_607,N_637);
nand U2323 (N_2323,N_670,N_1441);
nand U2324 (N_2324,N_1035,N_341);
or U2325 (N_2325,N_254,N_663);
or U2326 (N_2326,N_512,N_1286);
or U2327 (N_2327,N_1111,N_164);
xnor U2328 (N_2328,N_609,N_1455);
or U2329 (N_2329,N_205,N_493);
or U2330 (N_2330,N_1083,N_672);
xnor U2331 (N_2331,N_1427,N_938);
and U2332 (N_2332,N_1430,N_1325);
or U2333 (N_2333,N_103,N_1486);
nor U2334 (N_2334,N_99,N_84);
nor U2335 (N_2335,N_965,N_126);
and U2336 (N_2336,N_347,N_1364);
or U2337 (N_2337,N_315,N_913);
or U2338 (N_2338,N_1323,N_1454);
and U2339 (N_2339,N_903,N_531);
and U2340 (N_2340,N_1396,N_587);
nor U2341 (N_2341,N_1195,N_646);
xnor U2342 (N_2342,N_119,N_403);
or U2343 (N_2343,N_929,N_104);
nand U2344 (N_2344,N_32,N_233);
and U2345 (N_2345,N_1331,N_144);
nand U2346 (N_2346,N_940,N_204);
xor U2347 (N_2347,N_788,N_324);
xor U2348 (N_2348,N_1291,N_1206);
nor U2349 (N_2349,N_1427,N_1441);
xnor U2350 (N_2350,N_51,N_809);
xor U2351 (N_2351,N_734,N_640);
xnor U2352 (N_2352,N_748,N_535);
nand U2353 (N_2353,N_1039,N_272);
and U2354 (N_2354,N_1273,N_584);
nand U2355 (N_2355,N_315,N_1285);
and U2356 (N_2356,N_1132,N_339);
nand U2357 (N_2357,N_693,N_58);
nand U2358 (N_2358,N_1320,N_557);
nand U2359 (N_2359,N_1127,N_190);
nand U2360 (N_2360,N_1332,N_896);
or U2361 (N_2361,N_483,N_161);
and U2362 (N_2362,N_491,N_410);
and U2363 (N_2363,N_890,N_1383);
or U2364 (N_2364,N_1013,N_15);
xor U2365 (N_2365,N_1399,N_654);
nor U2366 (N_2366,N_1067,N_101);
nand U2367 (N_2367,N_189,N_254);
nand U2368 (N_2368,N_616,N_130);
nand U2369 (N_2369,N_1113,N_276);
or U2370 (N_2370,N_759,N_372);
nand U2371 (N_2371,N_1331,N_1184);
xor U2372 (N_2372,N_617,N_412);
and U2373 (N_2373,N_499,N_1291);
or U2374 (N_2374,N_1462,N_362);
nor U2375 (N_2375,N_147,N_296);
nor U2376 (N_2376,N_666,N_1452);
and U2377 (N_2377,N_1317,N_652);
nor U2378 (N_2378,N_252,N_229);
or U2379 (N_2379,N_377,N_753);
or U2380 (N_2380,N_148,N_1105);
or U2381 (N_2381,N_942,N_760);
or U2382 (N_2382,N_658,N_1005);
nand U2383 (N_2383,N_1077,N_648);
and U2384 (N_2384,N_205,N_1019);
and U2385 (N_2385,N_897,N_1051);
xnor U2386 (N_2386,N_966,N_1419);
and U2387 (N_2387,N_354,N_49);
xor U2388 (N_2388,N_827,N_775);
nor U2389 (N_2389,N_834,N_720);
nor U2390 (N_2390,N_1011,N_327);
xnor U2391 (N_2391,N_833,N_684);
or U2392 (N_2392,N_526,N_520);
nand U2393 (N_2393,N_214,N_636);
or U2394 (N_2394,N_1054,N_12);
or U2395 (N_2395,N_571,N_166);
nor U2396 (N_2396,N_824,N_913);
nand U2397 (N_2397,N_218,N_1128);
and U2398 (N_2398,N_1256,N_1048);
nand U2399 (N_2399,N_586,N_882);
or U2400 (N_2400,N_281,N_331);
nand U2401 (N_2401,N_63,N_1286);
nor U2402 (N_2402,N_232,N_1478);
and U2403 (N_2403,N_681,N_506);
or U2404 (N_2404,N_1478,N_1124);
xor U2405 (N_2405,N_1456,N_661);
and U2406 (N_2406,N_508,N_675);
nor U2407 (N_2407,N_330,N_7);
or U2408 (N_2408,N_1430,N_132);
xor U2409 (N_2409,N_1215,N_839);
nand U2410 (N_2410,N_854,N_322);
nand U2411 (N_2411,N_538,N_747);
and U2412 (N_2412,N_66,N_412);
xor U2413 (N_2413,N_907,N_1129);
or U2414 (N_2414,N_109,N_1121);
or U2415 (N_2415,N_1374,N_803);
nor U2416 (N_2416,N_26,N_951);
nand U2417 (N_2417,N_20,N_1018);
or U2418 (N_2418,N_398,N_314);
or U2419 (N_2419,N_1168,N_72);
xor U2420 (N_2420,N_478,N_838);
and U2421 (N_2421,N_119,N_50);
and U2422 (N_2422,N_1142,N_333);
and U2423 (N_2423,N_733,N_1448);
or U2424 (N_2424,N_1364,N_401);
nand U2425 (N_2425,N_853,N_508);
xnor U2426 (N_2426,N_1155,N_1464);
nand U2427 (N_2427,N_1080,N_366);
and U2428 (N_2428,N_441,N_1464);
nor U2429 (N_2429,N_120,N_1154);
and U2430 (N_2430,N_733,N_881);
xnor U2431 (N_2431,N_862,N_1314);
xor U2432 (N_2432,N_323,N_1211);
xor U2433 (N_2433,N_981,N_1422);
nand U2434 (N_2434,N_503,N_237);
xnor U2435 (N_2435,N_606,N_888);
xor U2436 (N_2436,N_103,N_153);
xnor U2437 (N_2437,N_698,N_681);
xor U2438 (N_2438,N_743,N_1052);
nand U2439 (N_2439,N_1122,N_500);
nand U2440 (N_2440,N_569,N_368);
or U2441 (N_2441,N_1156,N_1283);
nand U2442 (N_2442,N_192,N_510);
nand U2443 (N_2443,N_835,N_785);
xnor U2444 (N_2444,N_352,N_976);
or U2445 (N_2445,N_1353,N_1325);
nor U2446 (N_2446,N_987,N_1);
xor U2447 (N_2447,N_456,N_667);
nor U2448 (N_2448,N_369,N_331);
or U2449 (N_2449,N_632,N_39);
or U2450 (N_2450,N_643,N_362);
or U2451 (N_2451,N_535,N_1259);
xnor U2452 (N_2452,N_1296,N_635);
or U2453 (N_2453,N_760,N_1215);
nand U2454 (N_2454,N_541,N_249);
or U2455 (N_2455,N_303,N_1361);
nand U2456 (N_2456,N_1483,N_492);
nor U2457 (N_2457,N_1323,N_1376);
and U2458 (N_2458,N_969,N_1469);
nor U2459 (N_2459,N_1351,N_708);
and U2460 (N_2460,N_202,N_478);
nor U2461 (N_2461,N_781,N_1239);
and U2462 (N_2462,N_849,N_435);
xor U2463 (N_2463,N_426,N_493);
and U2464 (N_2464,N_104,N_391);
or U2465 (N_2465,N_284,N_793);
or U2466 (N_2466,N_378,N_1080);
or U2467 (N_2467,N_733,N_800);
nor U2468 (N_2468,N_143,N_957);
and U2469 (N_2469,N_934,N_1284);
and U2470 (N_2470,N_85,N_684);
nor U2471 (N_2471,N_945,N_538);
xor U2472 (N_2472,N_852,N_85);
and U2473 (N_2473,N_277,N_51);
or U2474 (N_2474,N_1051,N_655);
or U2475 (N_2475,N_1453,N_575);
xnor U2476 (N_2476,N_295,N_139);
xor U2477 (N_2477,N_1091,N_185);
or U2478 (N_2478,N_1057,N_341);
and U2479 (N_2479,N_89,N_916);
nor U2480 (N_2480,N_155,N_392);
nor U2481 (N_2481,N_1127,N_885);
and U2482 (N_2482,N_1383,N_1073);
nand U2483 (N_2483,N_349,N_308);
or U2484 (N_2484,N_445,N_11);
or U2485 (N_2485,N_230,N_1099);
xor U2486 (N_2486,N_500,N_65);
and U2487 (N_2487,N_902,N_283);
and U2488 (N_2488,N_231,N_307);
nand U2489 (N_2489,N_1106,N_1114);
xnor U2490 (N_2490,N_1256,N_815);
nor U2491 (N_2491,N_642,N_1037);
xnor U2492 (N_2492,N_1253,N_696);
xnor U2493 (N_2493,N_714,N_959);
nor U2494 (N_2494,N_535,N_1417);
and U2495 (N_2495,N_447,N_1121);
nand U2496 (N_2496,N_514,N_327);
xor U2497 (N_2497,N_119,N_941);
or U2498 (N_2498,N_1076,N_2);
or U2499 (N_2499,N_268,N_1317);
nand U2500 (N_2500,N_1336,N_533);
xor U2501 (N_2501,N_1141,N_1439);
nand U2502 (N_2502,N_90,N_253);
and U2503 (N_2503,N_62,N_470);
nor U2504 (N_2504,N_1430,N_1266);
or U2505 (N_2505,N_1009,N_526);
xor U2506 (N_2506,N_315,N_86);
nand U2507 (N_2507,N_1055,N_1134);
xnor U2508 (N_2508,N_1414,N_168);
or U2509 (N_2509,N_1095,N_340);
and U2510 (N_2510,N_541,N_747);
nand U2511 (N_2511,N_1232,N_447);
or U2512 (N_2512,N_1381,N_487);
xnor U2513 (N_2513,N_780,N_91);
xnor U2514 (N_2514,N_456,N_1027);
xor U2515 (N_2515,N_591,N_887);
and U2516 (N_2516,N_1352,N_807);
nand U2517 (N_2517,N_1008,N_1414);
and U2518 (N_2518,N_1251,N_141);
nor U2519 (N_2519,N_189,N_727);
and U2520 (N_2520,N_661,N_1041);
nor U2521 (N_2521,N_1179,N_1110);
or U2522 (N_2522,N_1430,N_932);
and U2523 (N_2523,N_1014,N_1152);
nor U2524 (N_2524,N_936,N_1226);
nand U2525 (N_2525,N_621,N_146);
nand U2526 (N_2526,N_1019,N_1217);
nor U2527 (N_2527,N_226,N_64);
nand U2528 (N_2528,N_1431,N_605);
nor U2529 (N_2529,N_832,N_878);
nor U2530 (N_2530,N_583,N_278);
nand U2531 (N_2531,N_159,N_1043);
nand U2532 (N_2532,N_1353,N_989);
xor U2533 (N_2533,N_1486,N_538);
or U2534 (N_2534,N_988,N_1203);
and U2535 (N_2535,N_923,N_108);
or U2536 (N_2536,N_467,N_399);
or U2537 (N_2537,N_279,N_222);
and U2538 (N_2538,N_1291,N_1417);
nand U2539 (N_2539,N_266,N_354);
and U2540 (N_2540,N_878,N_852);
xnor U2541 (N_2541,N_858,N_701);
nand U2542 (N_2542,N_1111,N_446);
and U2543 (N_2543,N_741,N_469);
nor U2544 (N_2544,N_1317,N_1068);
and U2545 (N_2545,N_875,N_1144);
nor U2546 (N_2546,N_691,N_1352);
and U2547 (N_2547,N_27,N_528);
nand U2548 (N_2548,N_766,N_202);
and U2549 (N_2549,N_768,N_1067);
nand U2550 (N_2550,N_425,N_1399);
xnor U2551 (N_2551,N_842,N_1161);
or U2552 (N_2552,N_408,N_588);
nor U2553 (N_2553,N_850,N_1120);
xnor U2554 (N_2554,N_852,N_687);
and U2555 (N_2555,N_1284,N_1051);
nor U2556 (N_2556,N_1002,N_1417);
and U2557 (N_2557,N_1360,N_1247);
and U2558 (N_2558,N_588,N_1297);
xnor U2559 (N_2559,N_998,N_491);
xnor U2560 (N_2560,N_131,N_1463);
nand U2561 (N_2561,N_716,N_563);
xnor U2562 (N_2562,N_1484,N_1168);
nor U2563 (N_2563,N_1090,N_553);
nand U2564 (N_2564,N_901,N_1365);
xnor U2565 (N_2565,N_412,N_1021);
nor U2566 (N_2566,N_665,N_1082);
or U2567 (N_2567,N_249,N_792);
or U2568 (N_2568,N_767,N_1344);
nor U2569 (N_2569,N_1483,N_511);
nor U2570 (N_2570,N_515,N_1032);
and U2571 (N_2571,N_121,N_365);
and U2572 (N_2572,N_463,N_592);
and U2573 (N_2573,N_1419,N_1270);
xnor U2574 (N_2574,N_536,N_1441);
or U2575 (N_2575,N_257,N_1090);
nor U2576 (N_2576,N_172,N_0);
or U2577 (N_2577,N_547,N_1056);
xor U2578 (N_2578,N_537,N_1226);
xor U2579 (N_2579,N_362,N_1105);
nor U2580 (N_2580,N_899,N_610);
or U2581 (N_2581,N_134,N_942);
nand U2582 (N_2582,N_866,N_1125);
or U2583 (N_2583,N_869,N_164);
nand U2584 (N_2584,N_1369,N_1306);
nand U2585 (N_2585,N_390,N_1430);
or U2586 (N_2586,N_325,N_695);
nand U2587 (N_2587,N_759,N_1326);
nand U2588 (N_2588,N_420,N_1276);
or U2589 (N_2589,N_531,N_875);
and U2590 (N_2590,N_31,N_890);
nor U2591 (N_2591,N_46,N_909);
nor U2592 (N_2592,N_373,N_501);
or U2593 (N_2593,N_1438,N_718);
or U2594 (N_2594,N_1101,N_289);
xor U2595 (N_2595,N_635,N_175);
and U2596 (N_2596,N_1381,N_1256);
or U2597 (N_2597,N_38,N_951);
nand U2598 (N_2598,N_1159,N_809);
or U2599 (N_2599,N_1214,N_83);
or U2600 (N_2600,N_69,N_1181);
nand U2601 (N_2601,N_102,N_498);
xnor U2602 (N_2602,N_1259,N_157);
and U2603 (N_2603,N_69,N_54);
and U2604 (N_2604,N_26,N_1452);
nand U2605 (N_2605,N_240,N_190);
xor U2606 (N_2606,N_471,N_879);
nand U2607 (N_2607,N_64,N_1373);
nand U2608 (N_2608,N_771,N_1359);
or U2609 (N_2609,N_130,N_291);
nand U2610 (N_2610,N_1408,N_887);
xor U2611 (N_2611,N_686,N_726);
or U2612 (N_2612,N_1097,N_47);
xor U2613 (N_2613,N_110,N_1441);
nor U2614 (N_2614,N_1005,N_1189);
xnor U2615 (N_2615,N_909,N_842);
and U2616 (N_2616,N_1053,N_40);
xor U2617 (N_2617,N_161,N_723);
nand U2618 (N_2618,N_982,N_1036);
xor U2619 (N_2619,N_159,N_1390);
xnor U2620 (N_2620,N_255,N_330);
or U2621 (N_2621,N_747,N_921);
nor U2622 (N_2622,N_738,N_816);
nand U2623 (N_2623,N_489,N_225);
or U2624 (N_2624,N_1472,N_1460);
and U2625 (N_2625,N_1432,N_223);
nor U2626 (N_2626,N_1382,N_740);
and U2627 (N_2627,N_265,N_343);
or U2628 (N_2628,N_1033,N_350);
nor U2629 (N_2629,N_703,N_238);
and U2630 (N_2630,N_953,N_190);
and U2631 (N_2631,N_834,N_312);
xnor U2632 (N_2632,N_1253,N_665);
nand U2633 (N_2633,N_480,N_700);
and U2634 (N_2634,N_195,N_1279);
nor U2635 (N_2635,N_915,N_791);
and U2636 (N_2636,N_372,N_1323);
and U2637 (N_2637,N_862,N_458);
and U2638 (N_2638,N_907,N_797);
and U2639 (N_2639,N_1060,N_277);
or U2640 (N_2640,N_1228,N_1475);
and U2641 (N_2641,N_256,N_1498);
nor U2642 (N_2642,N_900,N_41);
xor U2643 (N_2643,N_824,N_317);
xnor U2644 (N_2644,N_963,N_989);
or U2645 (N_2645,N_1321,N_833);
xnor U2646 (N_2646,N_1162,N_1230);
nor U2647 (N_2647,N_1423,N_557);
xnor U2648 (N_2648,N_126,N_655);
nor U2649 (N_2649,N_1213,N_1308);
or U2650 (N_2650,N_670,N_666);
and U2651 (N_2651,N_1000,N_709);
and U2652 (N_2652,N_179,N_1142);
xnor U2653 (N_2653,N_1139,N_153);
and U2654 (N_2654,N_607,N_31);
xor U2655 (N_2655,N_363,N_105);
nor U2656 (N_2656,N_634,N_293);
xor U2657 (N_2657,N_1018,N_1115);
xnor U2658 (N_2658,N_1036,N_391);
or U2659 (N_2659,N_1035,N_462);
xnor U2660 (N_2660,N_1373,N_1061);
nand U2661 (N_2661,N_1287,N_268);
and U2662 (N_2662,N_754,N_510);
or U2663 (N_2663,N_1380,N_216);
nand U2664 (N_2664,N_576,N_1223);
xnor U2665 (N_2665,N_585,N_1236);
or U2666 (N_2666,N_579,N_252);
and U2667 (N_2667,N_762,N_1486);
xor U2668 (N_2668,N_1464,N_490);
nor U2669 (N_2669,N_680,N_496);
and U2670 (N_2670,N_1405,N_156);
xor U2671 (N_2671,N_225,N_199);
and U2672 (N_2672,N_895,N_1383);
and U2673 (N_2673,N_1439,N_1432);
xor U2674 (N_2674,N_312,N_135);
xor U2675 (N_2675,N_1145,N_781);
and U2676 (N_2676,N_989,N_776);
and U2677 (N_2677,N_1141,N_1187);
and U2678 (N_2678,N_653,N_371);
nand U2679 (N_2679,N_927,N_1117);
xor U2680 (N_2680,N_631,N_160);
xor U2681 (N_2681,N_1114,N_7);
and U2682 (N_2682,N_1443,N_91);
nand U2683 (N_2683,N_589,N_784);
xor U2684 (N_2684,N_239,N_837);
or U2685 (N_2685,N_640,N_572);
and U2686 (N_2686,N_1029,N_333);
nand U2687 (N_2687,N_258,N_1482);
nor U2688 (N_2688,N_1431,N_1049);
nand U2689 (N_2689,N_476,N_1190);
and U2690 (N_2690,N_1184,N_69);
and U2691 (N_2691,N_1284,N_1347);
and U2692 (N_2692,N_1003,N_727);
nor U2693 (N_2693,N_502,N_776);
or U2694 (N_2694,N_1082,N_326);
xor U2695 (N_2695,N_760,N_725);
nor U2696 (N_2696,N_463,N_1232);
or U2697 (N_2697,N_1171,N_256);
xnor U2698 (N_2698,N_292,N_15);
nand U2699 (N_2699,N_1263,N_191);
nor U2700 (N_2700,N_1124,N_547);
nor U2701 (N_2701,N_324,N_532);
nand U2702 (N_2702,N_383,N_51);
nor U2703 (N_2703,N_186,N_59);
nor U2704 (N_2704,N_497,N_1016);
xnor U2705 (N_2705,N_518,N_1389);
nand U2706 (N_2706,N_901,N_776);
and U2707 (N_2707,N_78,N_1470);
and U2708 (N_2708,N_151,N_1180);
and U2709 (N_2709,N_308,N_1283);
or U2710 (N_2710,N_989,N_483);
xnor U2711 (N_2711,N_153,N_1357);
nand U2712 (N_2712,N_400,N_353);
and U2713 (N_2713,N_1070,N_545);
nor U2714 (N_2714,N_728,N_962);
or U2715 (N_2715,N_1305,N_604);
nor U2716 (N_2716,N_613,N_340);
nand U2717 (N_2717,N_411,N_41);
and U2718 (N_2718,N_1143,N_316);
or U2719 (N_2719,N_581,N_975);
and U2720 (N_2720,N_1451,N_147);
and U2721 (N_2721,N_1482,N_1494);
or U2722 (N_2722,N_1363,N_723);
xor U2723 (N_2723,N_935,N_861);
nand U2724 (N_2724,N_1293,N_812);
and U2725 (N_2725,N_1233,N_875);
nand U2726 (N_2726,N_889,N_366);
and U2727 (N_2727,N_28,N_386);
xnor U2728 (N_2728,N_1374,N_637);
or U2729 (N_2729,N_1493,N_1373);
and U2730 (N_2730,N_1356,N_380);
xor U2731 (N_2731,N_930,N_2);
xnor U2732 (N_2732,N_1483,N_1076);
nor U2733 (N_2733,N_1216,N_688);
nand U2734 (N_2734,N_76,N_731);
xnor U2735 (N_2735,N_805,N_286);
nor U2736 (N_2736,N_925,N_739);
nand U2737 (N_2737,N_1346,N_1095);
xnor U2738 (N_2738,N_1374,N_1012);
xor U2739 (N_2739,N_843,N_1469);
nand U2740 (N_2740,N_119,N_438);
or U2741 (N_2741,N_1495,N_1449);
and U2742 (N_2742,N_99,N_142);
nor U2743 (N_2743,N_977,N_720);
and U2744 (N_2744,N_732,N_588);
nand U2745 (N_2745,N_1425,N_751);
nor U2746 (N_2746,N_394,N_1329);
or U2747 (N_2747,N_373,N_471);
and U2748 (N_2748,N_581,N_703);
xnor U2749 (N_2749,N_154,N_1381);
and U2750 (N_2750,N_772,N_1331);
xor U2751 (N_2751,N_745,N_287);
nand U2752 (N_2752,N_29,N_204);
nand U2753 (N_2753,N_318,N_1200);
xnor U2754 (N_2754,N_268,N_766);
nor U2755 (N_2755,N_1479,N_935);
and U2756 (N_2756,N_777,N_2);
nor U2757 (N_2757,N_1096,N_630);
nand U2758 (N_2758,N_519,N_155);
xor U2759 (N_2759,N_831,N_596);
xor U2760 (N_2760,N_734,N_58);
or U2761 (N_2761,N_561,N_1173);
xor U2762 (N_2762,N_1269,N_870);
nand U2763 (N_2763,N_903,N_1283);
or U2764 (N_2764,N_129,N_773);
nor U2765 (N_2765,N_33,N_423);
xnor U2766 (N_2766,N_1037,N_1323);
nand U2767 (N_2767,N_1298,N_333);
or U2768 (N_2768,N_783,N_1152);
or U2769 (N_2769,N_144,N_792);
nand U2770 (N_2770,N_893,N_1108);
nor U2771 (N_2771,N_1221,N_803);
nand U2772 (N_2772,N_215,N_1450);
or U2773 (N_2773,N_524,N_820);
xor U2774 (N_2774,N_920,N_1368);
nand U2775 (N_2775,N_780,N_9);
or U2776 (N_2776,N_55,N_806);
xnor U2777 (N_2777,N_570,N_236);
nor U2778 (N_2778,N_1140,N_809);
nand U2779 (N_2779,N_900,N_974);
nand U2780 (N_2780,N_179,N_1304);
xor U2781 (N_2781,N_196,N_1113);
and U2782 (N_2782,N_96,N_1375);
or U2783 (N_2783,N_83,N_149);
xnor U2784 (N_2784,N_1480,N_641);
nand U2785 (N_2785,N_1409,N_904);
nor U2786 (N_2786,N_671,N_1339);
nand U2787 (N_2787,N_258,N_921);
nand U2788 (N_2788,N_179,N_689);
nand U2789 (N_2789,N_149,N_292);
xor U2790 (N_2790,N_749,N_1257);
or U2791 (N_2791,N_670,N_621);
or U2792 (N_2792,N_238,N_128);
and U2793 (N_2793,N_913,N_94);
and U2794 (N_2794,N_1349,N_920);
nand U2795 (N_2795,N_184,N_1243);
nor U2796 (N_2796,N_1194,N_86);
nor U2797 (N_2797,N_503,N_745);
nor U2798 (N_2798,N_48,N_780);
or U2799 (N_2799,N_890,N_1193);
xnor U2800 (N_2800,N_1041,N_700);
and U2801 (N_2801,N_1137,N_565);
nand U2802 (N_2802,N_1426,N_1154);
or U2803 (N_2803,N_125,N_888);
or U2804 (N_2804,N_464,N_465);
nor U2805 (N_2805,N_1243,N_447);
and U2806 (N_2806,N_449,N_1480);
and U2807 (N_2807,N_1445,N_138);
or U2808 (N_2808,N_690,N_555);
xor U2809 (N_2809,N_711,N_231);
nand U2810 (N_2810,N_698,N_1079);
nor U2811 (N_2811,N_318,N_253);
nor U2812 (N_2812,N_470,N_880);
nor U2813 (N_2813,N_134,N_496);
and U2814 (N_2814,N_392,N_1439);
or U2815 (N_2815,N_737,N_114);
or U2816 (N_2816,N_942,N_197);
xor U2817 (N_2817,N_131,N_13);
nand U2818 (N_2818,N_1193,N_72);
or U2819 (N_2819,N_256,N_218);
and U2820 (N_2820,N_1397,N_47);
or U2821 (N_2821,N_1389,N_786);
nand U2822 (N_2822,N_199,N_1017);
or U2823 (N_2823,N_1363,N_454);
xnor U2824 (N_2824,N_1299,N_34);
or U2825 (N_2825,N_428,N_1304);
and U2826 (N_2826,N_243,N_808);
xnor U2827 (N_2827,N_230,N_1263);
nand U2828 (N_2828,N_744,N_660);
nand U2829 (N_2829,N_968,N_790);
and U2830 (N_2830,N_464,N_1394);
xnor U2831 (N_2831,N_923,N_890);
and U2832 (N_2832,N_611,N_587);
nor U2833 (N_2833,N_1025,N_242);
xnor U2834 (N_2834,N_932,N_647);
xor U2835 (N_2835,N_658,N_1007);
and U2836 (N_2836,N_398,N_725);
or U2837 (N_2837,N_774,N_247);
nand U2838 (N_2838,N_1132,N_1011);
and U2839 (N_2839,N_1039,N_1266);
xnor U2840 (N_2840,N_1187,N_172);
and U2841 (N_2841,N_1234,N_972);
and U2842 (N_2842,N_175,N_1418);
nor U2843 (N_2843,N_1029,N_307);
or U2844 (N_2844,N_1270,N_1430);
and U2845 (N_2845,N_372,N_287);
xor U2846 (N_2846,N_793,N_576);
nand U2847 (N_2847,N_1338,N_28);
nor U2848 (N_2848,N_8,N_272);
nor U2849 (N_2849,N_1039,N_715);
nor U2850 (N_2850,N_205,N_618);
xnor U2851 (N_2851,N_459,N_354);
xor U2852 (N_2852,N_321,N_209);
and U2853 (N_2853,N_23,N_1156);
xor U2854 (N_2854,N_835,N_307);
and U2855 (N_2855,N_1421,N_1489);
nor U2856 (N_2856,N_1278,N_1256);
and U2857 (N_2857,N_332,N_117);
nand U2858 (N_2858,N_1098,N_130);
and U2859 (N_2859,N_1330,N_879);
and U2860 (N_2860,N_782,N_322);
xor U2861 (N_2861,N_774,N_738);
and U2862 (N_2862,N_318,N_1251);
nor U2863 (N_2863,N_1038,N_1213);
or U2864 (N_2864,N_327,N_98);
nand U2865 (N_2865,N_544,N_1203);
and U2866 (N_2866,N_1381,N_1401);
or U2867 (N_2867,N_469,N_1440);
and U2868 (N_2868,N_534,N_992);
and U2869 (N_2869,N_532,N_546);
nand U2870 (N_2870,N_770,N_91);
and U2871 (N_2871,N_220,N_562);
or U2872 (N_2872,N_120,N_805);
or U2873 (N_2873,N_16,N_783);
nand U2874 (N_2874,N_790,N_195);
and U2875 (N_2875,N_534,N_753);
xor U2876 (N_2876,N_1037,N_300);
nand U2877 (N_2877,N_502,N_778);
or U2878 (N_2878,N_1245,N_1415);
nor U2879 (N_2879,N_1093,N_1284);
or U2880 (N_2880,N_1240,N_1241);
nor U2881 (N_2881,N_69,N_1055);
nand U2882 (N_2882,N_1171,N_1435);
and U2883 (N_2883,N_1394,N_1473);
nor U2884 (N_2884,N_720,N_858);
or U2885 (N_2885,N_374,N_1082);
nand U2886 (N_2886,N_1104,N_435);
or U2887 (N_2887,N_658,N_495);
nor U2888 (N_2888,N_743,N_793);
nor U2889 (N_2889,N_1303,N_282);
and U2890 (N_2890,N_1254,N_731);
nand U2891 (N_2891,N_1109,N_1033);
or U2892 (N_2892,N_300,N_224);
xor U2893 (N_2893,N_799,N_1478);
nand U2894 (N_2894,N_522,N_211);
xnor U2895 (N_2895,N_1325,N_991);
xor U2896 (N_2896,N_1265,N_1109);
nor U2897 (N_2897,N_705,N_566);
xor U2898 (N_2898,N_1203,N_1222);
and U2899 (N_2899,N_504,N_438);
nand U2900 (N_2900,N_1171,N_849);
xnor U2901 (N_2901,N_185,N_1134);
nor U2902 (N_2902,N_154,N_1499);
or U2903 (N_2903,N_704,N_334);
nor U2904 (N_2904,N_281,N_354);
or U2905 (N_2905,N_643,N_579);
nand U2906 (N_2906,N_945,N_1150);
nor U2907 (N_2907,N_744,N_1174);
nor U2908 (N_2908,N_835,N_862);
nor U2909 (N_2909,N_166,N_756);
nand U2910 (N_2910,N_387,N_394);
and U2911 (N_2911,N_457,N_123);
nor U2912 (N_2912,N_334,N_990);
nor U2913 (N_2913,N_1170,N_991);
and U2914 (N_2914,N_28,N_716);
nor U2915 (N_2915,N_631,N_1261);
and U2916 (N_2916,N_761,N_728);
nor U2917 (N_2917,N_802,N_311);
xor U2918 (N_2918,N_911,N_582);
or U2919 (N_2919,N_418,N_1124);
nand U2920 (N_2920,N_1191,N_55);
nand U2921 (N_2921,N_17,N_72);
nand U2922 (N_2922,N_898,N_558);
and U2923 (N_2923,N_29,N_443);
xor U2924 (N_2924,N_271,N_877);
and U2925 (N_2925,N_1132,N_1086);
or U2926 (N_2926,N_877,N_509);
or U2927 (N_2927,N_438,N_29);
and U2928 (N_2928,N_337,N_406);
nor U2929 (N_2929,N_589,N_1354);
or U2930 (N_2930,N_1178,N_358);
and U2931 (N_2931,N_229,N_1322);
or U2932 (N_2932,N_1261,N_698);
xnor U2933 (N_2933,N_1236,N_116);
and U2934 (N_2934,N_1096,N_1480);
xnor U2935 (N_2935,N_1230,N_1091);
xnor U2936 (N_2936,N_962,N_1001);
and U2937 (N_2937,N_1213,N_880);
or U2938 (N_2938,N_1323,N_169);
and U2939 (N_2939,N_790,N_1275);
and U2940 (N_2940,N_306,N_903);
and U2941 (N_2941,N_132,N_1249);
nand U2942 (N_2942,N_645,N_1433);
nand U2943 (N_2943,N_1351,N_394);
or U2944 (N_2944,N_691,N_1068);
or U2945 (N_2945,N_1359,N_1380);
xnor U2946 (N_2946,N_1368,N_523);
or U2947 (N_2947,N_185,N_155);
and U2948 (N_2948,N_415,N_1255);
and U2949 (N_2949,N_828,N_581);
xor U2950 (N_2950,N_190,N_1492);
nor U2951 (N_2951,N_934,N_542);
and U2952 (N_2952,N_745,N_701);
and U2953 (N_2953,N_1074,N_688);
and U2954 (N_2954,N_721,N_833);
or U2955 (N_2955,N_759,N_611);
nand U2956 (N_2956,N_465,N_608);
nand U2957 (N_2957,N_716,N_561);
xor U2958 (N_2958,N_938,N_98);
or U2959 (N_2959,N_779,N_413);
xor U2960 (N_2960,N_429,N_148);
nor U2961 (N_2961,N_974,N_909);
xnor U2962 (N_2962,N_1446,N_714);
nor U2963 (N_2963,N_489,N_41);
or U2964 (N_2964,N_926,N_139);
nand U2965 (N_2965,N_1358,N_381);
and U2966 (N_2966,N_651,N_906);
or U2967 (N_2967,N_115,N_300);
nand U2968 (N_2968,N_913,N_478);
nor U2969 (N_2969,N_367,N_781);
nand U2970 (N_2970,N_1281,N_1054);
xnor U2971 (N_2971,N_1062,N_422);
nand U2972 (N_2972,N_1183,N_262);
nand U2973 (N_2973,N_874,N_363);
nor U2974 (N_2974,N_202,N_915);
nor U2975 (N_2975,N_881,N_974);
or U2976 (N_2976,N_1224,N_1046);
nor U2977 (N_2977,N_548,N_1369);
and U2978 (N_2978,N_1156,N_226);
and U2979 (N_2979,N_554,N_1342);
and U2980 (N_2980,N_668,N_587);
nand U2981 (N_2981,N_1135,N_1268);
nand U2982 (N_2982,N_512,N_1415);
xnor U2983 (N_2983,N_1469,N_300);
nand U2984 (N_2984,N_552,N_314);
xor U2985 (N_2985,N_880,N_818);
nor U2986 (N_2986,N_270,N_1262);
nand U2987 (N_2987,N_731,N_1214);
or U2988 (N_2988,N_451,N_801);
and U2989 (N_2989,N_1489,N_612);
and U2990 (N_2990,N_928,N_250);
and U2991 (N_2991,N_693,N_1460);
or U2992 (N_2992,N_1407,N_542);
xnor U2993 (N_2993,N_1307,N_436);
and U2994 (N_2994,N_1101,N_592);
xnor U2995 (N_2995,N_1071,N_1382);
or U2996 (N_2996,N_1156,N_300);
nor U2997 (N_2997,N_1330,N_578);
xor U2998 (N_2998,N_557,N_625);
and U2999 (N_2999,N_822,N_550);
xor U3000 (N_3000,N_1994,N_1883);
nor U3001 (N_3001,N_2444,N_2685);
and U3002 (N_3002,N_2747,N_2273);
and U3003 (N_3003,N_1795,N_2781);
xnor U3004 (N_3004,N_2011,N_2754);
nor U3005 (N_3005,N_1800,N_1873);
nor U3006 (N_3006,N_2723,N_1513);
nand U3007 (N_3007,N_2679,N_2043);
xnor U3008 (N_3008,N_2669,N_2980);
nand U3009 (N_3009,N_2154,N_2812);
nand U3010 (N_3010,N_1916,N_2144);
nor U3011 (N_3011,N_1984,N_1536);
xor U3012 (N_3012,N_2195,N_2831);
and U3013 (N_3013,N_2430,N_2921);
or U3014 (N_3014,N_2062,N_2982);
and U3015 (N_3015,N_2839,N_2339);
xor U3016 (N_3016,N_2010,N_1660);
xnor U3017 (N_3017,N_2616,N_2626);
xor U3018 (N_3018,N_2031,N_2354);
or U3019 (N_3019,N_2393,N_1540);
nor U3020 (N_3020,N_2032,N_1506);
or U3021 (N_3021,N_1977,N_1793);
or U3022 (N_3022,N_2186,N_2718);
xor U3023 (N_3023,N_1699,N_2618);
nand U3024 (N_3024,N_1673,N_1622);
nand U3025 (N_3025,N_2827,N_1568);
xnor U3026 (N_3026,N_2532,N_2058);
xor U3027 (N_3027,N_2145,N_2507);
or U3028 (N_3028,N_1954,N_2564);
nand U3029 (N_3029,N_2712,N_2651);
or U3030 (N_3030,N_2205,N_1970);
nor U3031 (N_3031,N_2592,N_1569);
or U3032 (N_3032,N_2080,N_2709);
xor U3033 (N_3033,N_2663,N_1767);
and U3034 (N_3034,N_2816,N_1841);
and U3035 (N_3035,N_2283,N_2544);
or U3036 (N_3036,N_2622,N_1700);
nor U3037 (N_3037,N_1606,N_2504);
nor U3038 (N_3038,N_2360,N_1556);
nor U3039 (N_3039,N_2732,N_1887);
and U3040 (N_3040,N_2837,N_1976);
xor U3041 (N_3041,N_1880,N_2192);
nand U3042 (N_3042,N_1871,N_1519);
or U3043 (N_3043,N_2127,N_2615);
and U3044 (N_3044,N_2091,N_1613);
nand U3045 (N_3045,N_2813,N_1683);
and U3046 (N_3046,N_2027,N_2920);
xnor U3047 (N_3047,N_2555,N_1902);
xnor U3048 (N_3048,N_2317,N_2560);
and U3049 (N_3049,N_2158,N_1624);
nand U3050 (N_3050,N_2017,N_2682);
and U3051 (N_3051,N_1864,N_2417);
xnor U3052 (N_3052,N_2316,N_2607);
or U3053 (N_3053,N_1741,N_2668);
nor U3054 (N_3054,N_2023,N_2968);
or U3055 (N_3055,N_1645,N_2635);
or U3056 (N_3056,N_1966,N_2940);
and U3057 (N_3057,N_2180,N_2092);
nor U3058 (N_3058,N_2614,N_1980);
nor U3059 (N_3059,N_1922,N_2101);
nand U3060 (N_3060,N_2434,N_2281);
nand U3061 (N_3061,N_2673,N_2882);
or U3062 (N_3062,N_1758,N_2196);
nand U3063 (N_3063,N_2600,N_2639);
or U3064 (N_3064,N_2647,N_2353);
xor U3065 (N_3065,N_2107,N_2655);
xnor U3066 (N_3066,N_2821,N_2586);
nor U3067 (N_3067,N_2112,N_2927);
or U3068 (N_3068,N_2806,N_2554);
and U3069 (N_3069,N_2719,N_2944);
or U3070 (N_3070,N_1670,N_1525);
nor U3071 (N_3071,N_1663,N_2495);
or U3072 (N_3072,N_2270,N_1773);
xnor U3073 (N_3073,N_2286,N_2585);
xor U3074 (N_3074,N_2276,N_2307);
nor U3075 (N_3075,N_2948,N_1579);
nor U3076 (N_3076,N_2213,N_2422);
nand U3077 (N_3077,N_2110,N_2476);
and U3078 (N_3078,N_2247,N_2876);
and U3079 (N_3079,N_2810,N_1859);
or U3080 (N_3080,N_2295,N_2318);
nor U3081 (N_3081,N_2451,N_1978);
nor U3082 (N_3082,N_2666,N_2922);
xor U3083 (N_3083,N_1739,N_2671);
nand U3084 (N_3084,N_1529,N_1655);
and U3085 (N_3085,N_1816,N_2960);
xnor U3086 (N_3086,N_2536,N_1761);
nor U3087 (N_3087,N_1627,N_2696);
nand U3088 (N_3088,N_1591,N_2202);
xor U3089 (N_3089,N_2184,N_2443);
and U3090 (N_3090,N_2603,N_1796);
nor U3091 (N_3091,N_2306,N_2082);
nand U3092 (N_3092,N_2912,N_1638);
nand U3093 (N_3093,N_2304,N_1596);
nand U3094 (N_3094,N_1913,N_1698);
nor U3095 (N_3095,N_1856,N_2249);
xor U3096 (N_3096,N_2363,N_1893);
and U3097 (N_3097,N_1764,N_2606);
xnor U3098 (N_3098,N_1675,N_2646);
and U3099 (N_3099,N_2569,N_2698);
or U3100 (N_3100,N_1840,N_1511);
nor U3101 (N_3101,N_1969,N_2266);
or U3102 (N_3102,N_2547,N_2338);
and U3103 (N_3103,N_2028,N_1528);
xnor U3104 (N_3104,N_2397,N_1690);
and U3105 (N_3105,N_2418,N_2431);
xnor U3106 (N_3106,N_2890,N_2764);
and U3107 (N_3107,N_2517,N_2176);
and U3108 (N_3108,N_2787,N_1743);
nand U3109 (N_3109,N_1892,N_2114);
and U3110 (N_3110,N_2975,N_2804);
xor U3111 (N_3111,N_1860,N_2456);
and U3112 (N_3112,N_2691,N_2420);
nor U3113 (N_3113,N_2264,N_2374);
xnor U3114 (N_3114,N_2933,N_2843);
or U3115 (N_3115,N_1659,N_1946);
xor U3116 (N_3116,N_2833,N_2542);
and U3117 (N_3117,N_2934,N_1787);
or U3118 (N_3118,N_2713,N_1538);
or U3119 (N_3119,N_2990,N_2825);
or U3120 (N_3120,N_2094,N_2343);
and U3121 (N_3121,N_1852,N_2983);
and U3122 (N_3122,N_2334,N_2391);
nor U3123 (N_3123,N_2593,N_1920);
nand U3124 (N_3124,N_2404,N_2278);
nor U3125 (N_3125,N_2897,N_2909);
and U3126 (N_3126,N_1714,N_2375);
and U3127 (N_3127,N_1881,N_2392);
nor U3128 (N_3128,N_2256,N_2178);
nand U3129 (N_3129,N_2893,N_2238);
and U3130 (N_3130,N_1935,N_2227);
nor U3131 (N_3131,N_2090,N_2520);
xnor U3132 (N_3132,N_1794,N_1983);
nor U3133 (N_3133,N_2974,N_1725);
xor U3134 (N_3134,N_1965,N_1708);
nor U3135 (N_3135,N_2291,N_2991);
xnor U3136 (N_3136,N_2182,N_2640);
and U3137 (N_3137,N_1592,N_2217);
nor U3138 (N_3138,N_2388,N_1680);
nand U3139 (N_3139,N_1771,N_2716);
nor U3140 (N_3140,N_1982,N_2401);
nor U3141 (N_3141,N_2779,N_2313);
nor U3142 (N_3142,N_2763,N_2570);
nand U3143 (N_3143,N_1737,N_1941);
xor U3144 (N_3144,N_1895,N_1792);
xnor U3145 (N_3145,N_2643,N_2026);
nand U3146 (N_3146,N_2997,N_2902);
xnor U3147 (N_3147,N_2051,N_2477);
and U3148 (N_3148,N_1598,N_2470);
and U3149 (N_3149,N_1918,N_2768);
or U3150 (N_3150,N_2595,N_2009);
or U3151 (N_3151,N_2487,N_1942);
and U3152 (N_3152,N_2598,N_1634);
or U3153 (N_3153,N_2840,N_2947);
nor U3154 (N_3154,N_2881,N_2059);
nand U3155 (N_3155,N_2147,N_2522);
nand U3156 (N_3156,N_1516,N_1582);
nand U3157 (N_3157,N_1843,N_2750);
nor U3158 (N_3158,N_1561,N_1998);
nand U3159 (N_3159,N_2057,N_1642);
or U3160 (N_3160,N_2644,N_2332);
xor U3161 (N_3161,N_1754,N_2138);
and U3162 (N_3162,N_2410,N_2419);
xor U3163 (N_3163,N_2796,N_2674);
xnor U3164 (N_3164,N_2539,N_2913);
and U3165 (N_3165,N_2736,N_2329);
nand U3166 (N_3166,N_2424,N_2302);
and U3167 (N_3167,N_1759,N_2442);
nand U3168 (N_3168,N_2856,N_1950);
or U3169 (N_3169,N_2282,N_2464);
or U3170 (N_3170,N_2686,N_2047);
nor U3171 (N_3171,N_1632,N_2244);
xor U3172 (N_3172,N_1697,N_2218);
nand U3173 (N_3173,N_1807,N_1594);
and U3174 (N_3174,N_2589,N_1502);
or U3175 (N_3175,N_1533,N_1952);
xnor U3176 (N_3176,N_2594,N_1581);
or U3177 (N_3177,N_1636,N_2061);
nor U3178 (N_3178,N_2002,N_1857);
xor U3179 (N_3179,N_1921,N_2926);
or U3180 (N_3180,N_2852,N_2908);
nor U3181 (N_3181,N_1701,N_2331);
nand U3182 (N_3182,N_2416,N_2402);
and U3183 (N_3183,N_1557,N_2848);
nor U3184 (N_3184,N_2650,N_2566);
xnor U3185 (N_3185,N_2753,N_1826);
nand U3186 (N_3186,N_2552,N_1580);
xnor U3187 (N_3187,N_1508,N_2224);
nand U3188 (N_3188,N_1957,N_2439);
xor U3189 (N_3189,N_2830,N_2008);
nand U3190 (N_3190,N_1571,N_2931);
nor U3191 (N_3191,N_1765,N_2194);
xnor U3192 (N_3192,N_1837,N_1629);
and U3193 (N_3193,N_2969,N_1710);
or U3194 (N_3194,N_2153,N_1786);
and U3195 (N_3195,N_1986,N_2999);
and U3196 (N_3196,N_1597,N_1832);
or U3197 (N_3197,N_1973,N_2398);
and U3198 (N_3198,N_2193,N_2540);
nor U3199 (N_3199,N_2269,N_1631);
nand U3200 (N_3200,N_1661,N_2183);
nand U3201 (N_3201,N_1809,N_2285);
xnor U3202 (N_3202,N_2054,N_2580);
and U3203 (N_3203,N_2007,N_1547);
xnor U3204 (N_3204,N_1886,N_2620);
nand U3205 (N_3205,N_1824,N_2628);
nand U3206 (N_3206,N_2099,N_2784);
nand U3207 (N_3207,N_2437,N_1707);
and U3208 (N_3208,N_2734,N_2708);
or U3209 (N_3209,N_2596,N_2248);
xor U3210 (N_3210,N_2314,N_2359);
and U3211 (N_3211,N_1963,N_2449);
or U3212 (N_3212,N_1929,N_2171);
xor U3213 (N_3213,N_1637,N_2945);
nand U3214 (N_3214,N_2019,N_2046);
xnor U3215 (N_3215,N_2219,N_2020);
nor U3216 (N_3216,N_1834,N_1926);
or U3217 (N_3217,N_2355,N_1992);
xnor U3218 (N_3218,N_2131,N_2978);
and U3219 (N_3219,N_1535,N_2150);
xor U3220 (N_3220,N_2220,N_2064);
nor U3221 (N_3221,N_2828,N_2799);
nand U3222 (N_3222,N_2661,N_2720);
xnor U3223 (N_3223,N_2457,N_2778);
or U3224 (N_3224,N_2413,N_2903);
nand U3225 (N_3225,N_2126,N_1900);
nor U3226 (N_3226,N_2526,N_1718);
and U3227 (N_3227,N_1885,N_2680);
and U3228 (N_3228,N_1563,N_2847);
and U3229 (N_3229,N_1940,N_2910);
xor U3230 (N_3230,N_1677,N_2040);
nand U3231 (N_3231,N_2930,N_1712);
or U3232 (N_3232,N_1818,N_2842);
nand U3233 (N_3233,N_2617,N_1811);
xor U3234 (N_3234,N_2965,N_2337);
nor U3235 (N_3235,N_2533,N_2148);
and U3236 (N_3236,N_1650,N_1762);
nand U3237 (N_3237,N_2993,N_2854);
xor U3238 (N_3238,N_2105,N_2130);
or U3239 (N_3239,N_2341,N_2369);
nor U3240 (N_3240,N_1932,N_1838);
nand U3241 (N_3241,N_1748,N_1769);
nand U3242 (N_3242,N_2385,N_2717);
or U3243 (N_3243,N_2645,N_1797);
or U3244 (N_3244,N_2488,N_1713);
and U3245 (N_3245,N_2116,N_1924);
xnor U3246 (N_3246,N_1740,N_2021);
nand U3247 (N_3247,N_2803,N_1602);
and U3248 (N_3248,N_2853,N_2378);
or U3249 (N_3249,N_2085,N_1831);
nor U3250 (N_3250,N_1609,N_2037);
and U3251 (N_3251,N_2395,N_2350);
and U3252 (N_3252,N_2067,N_2056);
and U3253 (N_3253,N_2177,N_2642);
xor U3254 (N_3254,N_2521,N_1968);
xnor U3255 (N_3255,N_1728,N_2272);
xor U3256 (N_3256,N_1651,N_2214);
xor U3257 (N_3257,N_2115,N_1835);
nand U3258 (N_3258,N_2946,N_2445);
nor U3259 (N_3259,N_2063,N_2845);
nor U3260 (N_3260,N_2469,N_1641);
nor U3261 (N_3261,N_2896,N_2299);
and U3262 (N_3262,N_2929,N_2838);
xnor U3263 (N_3263,N_2396,N_2376);
and U3264 (N_3264,N_1894,N_1515);
or U3265 (N_3265,N_2868,N_1925);
or U3266 (N_3266,N_2407,N_1665);
xnor U3267 (N_3267,N_2041,N_2265);
nand U3268 (N_3268,N_2044,N_2769);
nand U3269 (N_3269,N_1821,N_2458);
xnor U3270 (N_3270,N_2862,N_2260);
or U3271 (N_3271,N_2365,N_1991);
nand U3272 (N_3272,N_2473,N_1589);
nor U3273 (N_3273,N_2746,N_2344);
nor U3274 (N_3274,N_2489,N_1944);
nand U3275 (N_3275,N_2454,N_2400);
xor U3276 (N_3276,N_2918,N_2258);
and U3277 (N_3277,N_1791,N_2226);
nand U3278 (N_3278,N_1987,N_1640);
xor U3279 (N_3279,N_2478,N_2807);
and U3280 (N_3280,N_1676,N_2766);
xnor U3281 (N_3281,N_2321,N_2394);
nor U3282 (N_3282,N_2486,N_2894);
nor U3283 (N_3283,N_2887,N_1576);
nor U3284 (N_3284,N_2120,N_2137);
or U3285 (N_3285,N_2966,N_1827);
xnor U3286 (N_3286,N_2721,N_2572);
xnor U3287 (N_3287,N_2151,N_2652);
nand U3288 (N_3288,N_2704,N_1644);
or U3289 (N_3289,N_1679,N_2060);
and U3290 (N_3290,N_2514,N_2662);
nand U3291 (N_3291,N_2301,N_2914);
nand U3292 (N_3292,N_1825,N_1912);
or U3293 (N_3293,N_2867,N_2087);
xor U3294 (N_3294,N_2943,N_1903);
xnor U3295 (N_3295,N_2860,N_1964);
and U3296 (N_3296,N_1546,N_2294);
nand U3297 (N_3297,N_2878,N_2157);
or U3298 (N_3298,N_1779,N_1667);
xor U3299 (N_3299,N_2525,N_1847);
nand U3300 (N_3300,N_1879,N_2568);
xnor U3301 (N_3301,N_2911,N_1652);
nand U3302 (N_3302,N_2078,N_1653);
nor U3303 (N_3303,N_1620,N_2873);
xor U3304 (N_3304,N_2608,N_2098);
or U3305 (N_3305,N_1989,N_2271);
nor U3306 (N_3306,N_1774,N_2826);
and U3307 (N_3307,N_2069,N_2461);
and U3308 (N_3308,N_2004,N_2728);
and U3309 (N_3309,N_2726,N_2516);
and U3310 (N_3310,N_2700,N_1830);
xnor U3311 (N_3311,N_2233,N_1848);
xnor U3312 (N_3312,N_2875,N_2428);
or U3313 (N_3313,N_2795,N_1836);
xor U3314 (N_3314,N_2573,N_2072);
nand U3315 (N_3315,N_1789,N_1757);
xor U3316 (N_3316,N_2578,N_2328);
xor U3317 (N_3317,N_2528,N_2907);
nand U3318 (N_3318,N_2268,N_2279);
and U3319 (N_3319,N_2380,N_1874);
or U3320 (N_3320,N_2333,N_1906);
nor U3321 (N_3321,N_2379,N_2776);
nor U3322 (N_3322,N_2950,N_1972);
and U3323 (N_3323,N_1909,N_2001);
nor U3324 (N_3324,N_1822,N_2955);
xor U3325 (N_3325,N_2135,N_2971);
nand U3326 (N_3326,N_1806,N_1878);
xor U3327 (N_3327,N_1844,N_2591);
and U3328 (N_3328,N_2012,N_2710);
and U3329 (N_3329,N_2928,N_2924);
nor U3330 (N_3330,N_2935,N_1552);
nand U3331 (N_3331,N_2808,N_2039);
nor U3332 (N_3332,N_1975,N_1993);
xor U3333 (N_3333,N_2818,N_2246);
xor U3334 (N_3334,N_1749,N_1522);
nand U3335 (N_3335,N_1617,N_2427);
nand U3336 (N_3336,N_2221,N_2436);
or U3337 (N_3337,N_1805,N_1560);
or U3338 (N_3338,N_2203,N_1958);
nand U3339 (N_3339,N_2823,N_2822);
xor U3340 (N_3340,N_2311,N_2237);
and U3341 (N_3341,N_2494,N_2871);
or U3342 (N_3342,N_2888,N_2450);
and U3343 (N_3343,N_1599,N_1949);
nand U3344 (N_3344,N_2730,N_2013);
nand U3345 (N_3345,N_2267,N_2312);
nor U3346 (N_3346,N_2414,N_2179);
and U3347 (N_3347,N_2513,N_2065);
xor U3348 (N_3348,N_2096,N_2364);
or U3349 (N_3349,N_1514,N_2531);
nor U3350 (N_3350,N_1775,N_2932);
xor U3351 (N_3351,N_2741,N_2073);
nor U3352 (N_3352,N_2421,N_2623);
or U3353 (N_3353,N_2111,N_2289);
and U3354 (N_3354,N_2426,N_2462);
nor U3355 (N_3355,N_2979,N_1876);
nand U3356 (N_3356,N_2134,N_2780);
nand U3357 (N_3357,N_2467,N_2624);
nor U3358 (N_3358,N_2849,N_2706);
and U3359 (N_3359,N_2786,N_2234);
nand U3360 (N_3360,N_1961,N_2699);
xor U3361 (N_3361,N_2201,N_1584);
xnor U3362 (N_3362,N_1517,N_2738);
and U3363 (N_3363,N_2656,N_1565);
nand U3364 (N_3364,N_2015,N_1723);
xnor U3365 (N_3365,N_2174,N_1891);
nor U3366 (N_3366,N_2325,N_2599);
nor U3367 (N_3367,N_1782,N_1727);
and U3368 (N_3368,N_1829,N_1587);
xor U3369 (N_3369,N_2697,N_1541);
nand U3370 (N_3370,N_2297,N_1904);
xor U3371 (N_3371,N_1803,N_2481);
nand U3372 (N_3372,N_2370,N_2387);
nand U3373 (N_3373,N_2199,N_2155);
xor U3374 (N_3374,N_2565,N_2625);
nand U3375 (N_3375,N_1997,N_2025);
and U3376 (N_3376,N_1643,N_2200);
nand U3377 (N_3377,N_1567,N_2366);
xnor U3378 (N_3378,N_2794,N_2883);
and U3379 (N_3379,N_2904,N_2100);
or U3380 (N_3380,N_1823,N_2739);
nand U3381 (N_3381,N_2801,N_2242);
and U3382 (N_3382,N_2485,N_2949);
or U3383 (N_3383,N_2143,N_2895);
and U3384 (N_3384,N_1619,N_2745);
nor U3385 (N_3385,N_1687,N_2084);
nand U3386 (N_3386,N_2089,N_2851);
or U3387 (N_3387,N_2558,N_1890);
nand U3388 (N_3388,N_2384,N_1988);
nand U3389 (N_3389,N_1504,N_2638);
and U3390 (N_3390,N_2440,N_2511);
xnor U3391 (N_3391,N_1751,N_2479);
xnor U3392 (N_3392,N_2140,N_1910);
xor U3393 (N_3393,N_2164,N_1635);
and U3394 (N_3394,N_1649,N_2172);
or U3395 (N_3395,N_2577,N_2232);
nand U3396 (N_3396,N_2406,N_2253);
or U3397 (N_3397,N_1731,N_2231);
nand U3398 (N_3398,N_1745,N_1744);
and U3399 (N_3399,N_2777,N_1575);
or U3400 (N_3400,N_2129,N_2024);
or U3401 (N_3401,N_2689,N_2800);
or U3402 (N_3402,N_1586,N_2029);
xor U3403 (N_3403,N_2841,N_1542);
nor U3404 (N_3404,N_2235,N_2748);
xnor U3405 (N_3405,N_2447,N_2453);
or U3406 (N_3406,N_2412,N_2052);
nor U3407 (N_3407,N_2798,N_1889);
or U3408 (N_3408,N_1500,N_1730);
nor U3409 (N_3409,N_1842,N_2973);
or U3410 (N_3410,N_2760,N_1877);
nand U3411 (N_3411,N_2405,N_2954);
and U3412 (N_3412,N_2670,N_2582);
or U3413 (N_3413,N_1526,N_2866);
nand U3414 (N_3414,N_2208,N_2659);
nand U3415 (N_3415,N_2225,N_2240);
and U3416 (N_3416,N_2634,N_1742);
or U3417 (N_3417,N_2347,N_1870);
or U3418 (N_3418,N_2538,N_1604);
xnor U3419 (N_3419,N_1593,N_2071);
and U3420 (N_3420,N_1603,N_2688);
xor U3421 (N_3421,N_2744,N_1947);
xnor U3422 (N_3422,N_2381,N_2229);
and U3423 (N_3423,N_1899,N_1763);
nand U3424 (N_3424,N_2335,N_2465);
or U3425 (N_3425,N_2601,N_2702);
nor U3426 (N_3426,N_1555,N_2508);
nor U3427 (N_3427,N_2677,N_1548);
or U3428 (N_3428,N_1549,N_2588);
nand U3429 (N_3429,N_2373,N_1756);
xor U3430 (N_3430,N_1945,N_2916);
and U3431 (N_3431,N_1768,N_2937);
xnor U3432 (N_3432,N_2168,N_2658);
or U3433 (N_3433,N_2499,N_1608);
nor U3434 (N_3434,N_2315,N_2128);
or U3435 (N_3435,N_2792,N_1884);
xor U3436 (N_3436,N_2117,N_1573);
xor U3437 (N_3437,N_2549,N_1717);
nand U3438 (N_3438,N_2079,N_1734);
or U3439 (N_3439,N_1553,N_1674);
nand U3440 (N_3440,N_2348,N_2006);
or U3441 (N_3441,N_2602,N_2259);
and U3442 (N_3442,N_2684,N_1705);
xor U3443 (N_3443,N_1990,N_1703);
xnor U3444 (N_3444,N_2263,N_1785);
nand U3445 (N_3445,N_2774,N_1908);
nor U3446 (N_3446,N_2579,N_2492);
xor U3447 (N_3447,N_2132,N_2113);
nor U3448 (N_3448,N_2257,N_1951);
nor U3449 (N_3449,N_2610,N_2701);
and U3450 (N_3450,N_1539,N_2563);
nor U3451 (N_3451,N_2613,N_2038);
xor U3452 (N_3452,N_2254,N_1915);
nor U3453 (N_3453,N_1766,N_2068);
or U3454 (N_3454,N_2125,N_2676);
nand U3455 (N_3455,N_2305,N_1815);
xnor U3456 (N_3456,N_2362,N_2022);
xor U3457 (N_3457,N_2575,N_2915);
and U3458 (N_3458,N_2802,N_2829);
and U3459 (N_3459,N_1578,N_1999);
or U3460 (N_3460,N_2767,N_1657);
and U3461 (N_3461,N_1696,N_1760);
nor U3462 (N_3462,N_1671,N_2995);
or U3463 (N_3463,N_1865,N_2290);
nor U3464 (N_3464,N_1817,N_2501);
nand U3465 (N_3465,N_2204,N_1928);
nand U3466 (N_3466,N_2751,N_1543);
and U3467 (N_3467,N_2733,N_2743);
and U3468 (N_3468,N_2793,N_1595);
xnor U3469 (N_3469,N_2118,N_2463);
nand U3470 (N_3470,N_2740,N_1778);
nor U3471 (N_3471,N_1798,N_1570);
xnor U3472 (N_3472,N_2389,N_1802);
nand U3473 (N_3473,N_2493,N_1666);
nand U3474 (N_3474,N_2874,N_2055);
or U3475 (N_3475,N_1882,N_1981);
nand U3476 (N_3476,N_2216,N_2844);
nor U3477 (N_3477,N_2729,N_1611);
nor U3478 (N_3478,N_2324,N_2455);
xor U3479 (N_3479,N_1733,N_1623);
nand U3480 (N_3480,N_2210,N_2857);
xnor U3481 (N_3481,N_2992,N_1931);
nor U3482 (N_3482,N_2711,N_2088);
nand U3483 (N_3483,N_2503,N_2496);
and U3484 (N_3484,N_2277,N_1588);
and U3485 (N_3485,N_2858,N_1804);
nor U3486 (N_3486,N_2095,N_2432);
nand U3487 (N_3487,N_2797,N_2681);
nor U3488 (N_3488,N_2475,N_2102);
nand U3489 (N_3489,N_2835,N_2707);
and U3490 (N_3490,N_2925,N_2251);
or U3491 (N_3491,N_1985,N_2597);
nand U3492 (N_3492,N_2206,N_2322);
xor U3493 (N_3493,N_2149,N_1783);
and U3494 (N_3494,N_2988,N_2274);
xnor U3495 (N_3495,N_2292,N_2901);
and U3496 (N_3496,N_1505,N_2399);
nor U3497 (N_3497,N_1618,N_2212);
and U3498 (N_3498,N_1849,N_2627);
nor U3499 (N_3499,N_1692,N_2611);
xnor U3500 (N_3500,N_2466,N_2529);
or U3501 (N_3501,N_2109,N_2692);
or U3502 (N_3502,N_2497,N_2790);
nor U3503 (N_3503,N_2003,N_2211);
nand U3504 (N_3504,N_2411,N_1639);
xnor U3505 (N_3505,N_2587,N_2941);
nor U3506 (N_3506,N_1685,N_2959);
nand U3507 (N_3507,N_1858,N_1550);
and U3508 (N_3508,N_2961,N_2124);
xnor U3509 (N_3509,N_1704,N_1735);
xnor U3510 (N_3510,N_2619,N_2425);
and U3511 (N_3511,N_1559,N_2243);
nand U3512 (N_3512,N_2996,N_2185);
xor U3513 (N_3513,N_2288,N_1810);
nand U3514 (N_3514,N_2345,N_2571);
nor U3515 (N_3515,N_1566,N_1715);
nor U3516 (N_3516,N_1750,N_1630);
or U3517 (N_3517,N_2275,N_1562);
xnor U3518 (N_3518,N_2715,N_2879);
nor U3519 (N_3519,N_1537,N_1583);
nor U3520 (N_3520,N_2141,N_2584);
xor U3521 (N_3521,N_2498,N_1753);
nor U3522 (N_3522,N_2678,N_2724);
nand U3523 (N_3523,N_2782,N_2320);
xnor U3524 (N_3524,N_1672,N_2000);
xnor U3525 (N_3525,N_2574,N_2173);
nand U3526 (N_3526,N_2252,N_1719);
nand U3527 (N_3527,N_2632,N_2358);
xnor U3528 (N_3528,N_2905,N_1846);
or U3529 (N_3529,N_2817,N_2972);
or U3530 (N_3530,N_2484,N_1558);
and U3531 (N_3531,N_2885,N_2994);
or U3532 (N_3532,N_1610,N_2984);
or U3533 (N_3533,N_1694,N_2326);
nor U3534 (N_3534,N_2880,N_2770);
nand U3535 (N_3535,N_1654,N_2198);
nand U3536 (N_3536,N_2014,N_1996);
nand U3537 (N_3537,N_1626,N_1682);
xor U3538 (N_3538,N_2005,N_2703);
xnor U3539 (N_3539,N_2438,N_2296);
xor U3540 (N_3540,N_1691,N_1788);
or U3541 (N_3541,N_2284,N_2308);
xor U3542 (N_3542,N_1646,N_2725);
xnor U3543 (N_3543,N_2609,N_2761);
nor U3544 (N_3544,N_2156,N_2472);
or U3545 (N_3545,N_2048,N_2519);
or U3546 (N_3546,N_1633,N_1720);
nand U3547 (N_3547,N_2383,N_2742);
or U3548 (N_3548,N_2665,N_1601);
and U3549 (N_3549,N_2053,N_2239);
nor U3550 (N_3550,N_2367,N_1554);
or U3551 (N_3551,N_2811,N_1564);
nand U3552 (N_3552,N_2865,N_1861);
and U3553 (N_3553,N_2352,N_2884);
nor U3554 (N_3554,N_2323,N_2336);
nor U3555 (N_3555,N_2783,N_2737);
xor U3556 (N_3556,N_1868,N_2919);
or U3557 (N_3557,N_2429,N_1572);
nand U3558 (N_3558,N_1510,N_2900);
nor U3559 (N_3559,N_1875,N_2550);
and U3560 (N_3560,N_2649,N_2523);
nand U3561 (N_3561,N_1668,N_2474);
nor U3562 (N_3562,N_2448,N_2557);
or U3563 (N_3563,N_2809,N_2361);
and U3564 (N_3564,N_1948,N_1896);
nand U3565 (N_3565,N_1784,N_2951);
nor U3566 (N_3566,N_2690,N_1702);
nor U3567 (N_3567,N_1960,N_1722);
nor U3568 (N_3568,N_2500,N_1907);
xnor U3569 (N_3569,N_2408,N_1656);
nor U3570 (N_3570,N_2403,N_2163);
nand U3571 (N_3571,N_1585,N_2104);
and U3572 (N_3572,N_2106,N_2446);
or U3573 (N_3573,N_2788,N_1509);
and U3574 (N_3574,N_2505,N_2899);
xnor U3575 (N_3575,N_2319,N_1616);
nand U3576 (N_3576,N_2819,N_2967);
and U3577 (N_3577,N_2162,N_2491);
nor U3578 (N_3578,N_2667,N_2166);
and U3579 (N_3579,N_2018,N_2832);
and U3580 (N_3580,N_1914,N_2938);
and U3581 (N_3581,N_2820,N_2357);
nand U3582 (N_3582,N_1937,N_2789);
nor U3583 (N_3583,N_1738,N_2191);
or U3584 (N_3584,N_2340,N_2382);
or U3585 (N_3585,N_1854,N_2121);
nand U3586 (N_3586,N_2309,N_2836);
xnor U3587 (N_3587,N_1607,N_1869);
nor U3588 (N_3588,N_1621,N_1979);
xnor U3589 (N_3589,N_2834,N_2752);
nand U3590 (N_3590,N_2872,N_1962);
or U3591 (N_3591,N_2633,N_2970);
xor U3592 (N_3592,N_1664,N_2963);
nand U3593 (N_3593,N_1647,N_2654);
nor U3594 (N_3594,N_1724,N_2016);
and U3595 (N_3595,N_1901,N_2714);
and U3596 (N_3596,N_2527,N_2985);
and U3597 (N_3597,N_2765,N_2330);
or U3598 (N_3598,N_1897,N_2327);
xor U3599 (N_3599,N_1855,N_2035);
or U3600 (N_3600,N_1706,N_2502);
xor U3601 (N_3601,N_2230,N_2228);
and U3602 (N_3602,N_2386,N_2189);
and U3603 (N_3603,N_1551,N_2371);
nor U3604 (N_3604,N_2349,N_2906);
nand U3605 (N_3605,N_2197,N_1689);
and U3606 (N_3606,N_2553,N_2705);
nor U3607 (N_3607,N_2641,N_1612);
xnor U3608 (N_3608,N_1726,N_2310);
or U3609 (N_3609,N_1938,N_2683);
nand U3610 (N_3610,N_2562,N_2863);
nand U3611 (N_3611,N_2898,N_2877);
and U3612 (N_3612,N_2621,N_2460);
nand U3613 (N_3613,N_2964,N_2952);
xor U3614 (N_3614,N_2303,N_1781);
or U3615 (N_3615,N_1801,N_2824);
nor U3616 (N_3616,N_2986,N_2524);
nor U3617 (N_3617,N_1820,N_2280);
xnor U3618 (N_3618,N_1930,N_1772);
nor U3619 (N_3619,N_1845,N_2561);
xor U3620 (N_3620,N_1605,N_2356);
xnor U3621 (N_3621,N_2660,N_1863);
nor U3622 (N_3622,N_1524,N_1736);
or U3623 (N_3623,N_1780,N_1956);
nor U3624 (N_3624,N_2987,N_2695);
and U3625 (N_3625,N_2409,N_2490);
and U3626 (N_3626,N_1628,N_1531);
xor U3627 (N_3627,N_1799,N_2583);
or U3628 (N_3628,N_1839,N_2042);
nand U3629 (N_3629,N_2546,N_1967);
or U3630 (N_3630,N_1658,N_2033);
nor U3631 (N_3631,N_2423,N_2815);
nor U3632 (N_3632,N_2142,N_2075);
nor U3633 (N_3633,N_2771,N_1648);
nor U3634 (N_3634,N_2605,N_2859);
xor U3635 (N_3635,N_2630,N_2441);
xor U3636 (N_3636,N_1919,N_2515);
nor U3637 (N_3637,N_1933,N_2636);
xnor U3638 (N_3638,N_1833,N_2604);
or U3639 (N_3639,N_2590,N_2083);
and U3640 (N_3640,N_2187,N_2772);
xnor U3641 (N_3641,N_2977,N_1732);
xnor U3642 (N_3642,N_2510,N_1974);
or U3643 (N_3643,N_2170,N_1577);
or U3644 (N_3644,N_2215,N_2942);
nand U3645 (N_3645,N_2159,N_2372);
nand U3646 (N_3646,N_2509,N_2755);
nor U3647 (N_3647,N_2958,N_2245);
nor U3648 (N_3648,N_1716,N_1888);
xor U3649 (N_3649,N_2030,N_2637);
or U3650 (N_3650,N_2165,N_2103);
nor U3651 (N_3651,N_2188,N_1681);
nor U3652 (N_3652,N_1615,N_2482);
and U3653 (N_3653,N_2086,N_1953);
nand U3654 (N_3654,N_2548,N_2066);
nand U3655 (N_3655,N_2675,N_1532);
or U3656 (N_3656,N_2175,N_1614);
xor U3657 (N_3657,N_1625,N_2433);
and U3658 (N_3658,N_1711,N_2814);
or U3659 (N_3659,N_2864,N_1662);
nand U3660 (N_3660,N_2119,N_2756);
nand U3661 (N_3661,N_2076,N_1943);
nand U3662 (N_3662,N_1521,N_1695);
nand U3663 (N_3663,N_1911,N_2850);
nand U3664 (N_3664,N_1923,N_2506);
nor U3665 (N_3665,N_2435,N_2889);
xor U3666 (N_3666,N_2537,N_1693);
and U3667 (N_3667,N_2222,N_2886);
nor U3668 (N_3668,N_2209,N_1867);
and U3669 (N_3669,N_1721,N_2541);
xnor U3670 (N_3670,N_1523,N_1819);
nand U3671 (N_3671,N_2250,N_1936);
nor U3672 (N_3672,N_2368,N_2459);
and U3673 (N_3673,N_2693,N_2545);
xor U3674 (N_3674,N_2390,N_2181);
nand U3675 (N_3675,N_1971,N_1777);
nand U3676 (N_3676,N_2050,N_2559);
xor U3677 (N_3677,N_2846,N_2581);
and U3678 (N_3678,N_2300,N_2664);
and U3679 (N_3679,N_2223,N_2108);
nor U3680 (N_3680,N_1955,N_2262);
and U3681 (N_3681,N_2512,N_2791);
nor U3682 (N_3682,N_1853,N_2731);
xnor U3683 (N_3683,N_1828,N_1862);
xnor U3684 (N_3684,N_2190,N_1747);
nor U3685 (N_3685,N_2727,N_2346);
and U3686 (N_3686,N_2480,N_1995);
and U3687 (N_3687,N_2122,N_2535);
or U3688 (N_3688,N_1770,N_1746);
nand U3689 (N_3689,N_2070,N_1501);
or U3690 (N_3690,N_2483,N_2152);
nor U3691 (N_3691,N_1850,N_2074);
nor U3692 (N_3692,N_2758,N_2762);
nor U3693 (N_3693,N_1813,N_2093);
and U3694 (N_3694,N_2293,N_2939);
nand U3695 (N_3695,N_2161,N_1534);
nand U3696 (N_3696,N_1518,N_1814);
nand U3697 (N_3697,N_2870,N_2998);
or U3698 (N_3698,N_1959,N_2133);
xor U3699 (N_3699,N_2631,N_1507);
nor U3700 (N_3700,N_1808,N_2146);
xnor U3701 (N_3701,N_2518,N_1927);
and U3702 (N_3702,N_1600,N_1851);
nor U3703 (N_3703,N_2160,N_1544);
or U3704 (N_3704,N_2081,N_2236);
and U3705 (N_3705,N_2169,N_2773);
xor U3706 (N_3706,N_2936,N_2036);
xnor U3707 (N_3707,N_1527,N_2298);
and U3708 (N_3708,N_1866,N_2471);
nand U3709 (N_3709,N_1669,N_2377);
and U3710 (N_3710,N_2759,N_2749);
nor U3711 (N_3711,N_2468,N_2045);
nand U3712 (N_3712,N_1790,N_2657);
nand U3713 (N_3713,N_1898,N_2989);
xnor U3714 (N_3714,N_2287,N_2556);
or U3715 (N_3715,N_2452,N_2891);
or U3716 (N_3716,N_2722,N_1686);
nor U3717 (N_3717,N_2049,N_2855);
or U3718 (N_3718,N_2775,N_1939);
or U3719 (N_3719,N_2342,N_1684);
or U3720 (N_3720,N_2139,N_1530);
nand U3721 (N_3721,N_1590,N_2534);
and U3722 (N_3722,N_2123,N_2077);
nand U3723 (N_3723,N_2861,N_1872);
nor U3724 (N_3724,N_2785,N_2957);
nor U3725 (N_3725,N_1917,N_2976);
or U3726 (N_3726,N_2097,N_1812);
nand U3727 (N_3727,N_2892,N_2917);
nor U3728 (N_3728,N_1755,N_2415);
or U3729 (N_3729,N_1678,N_2034);
and U3730 (N_3730,N_1729,N_2735);
and U3731 (N_3731,N_2981,N_1905);
nand U3732 (N_3732,N_2953,N_2261);
and U3733 (N_3733,N_2672,N_1776);
nand U3734 (N_3734,N_2956,N_1512);
xnor U3735 (N_3735,N_1574,N_2567);
and U3736 (N_3736,N_2653,N_2612);
and U3737 (N_3737,N_2241,N_1688);
nand U3738 (N_3738,N_2648,N_2869);
and U3739 (N_3739,N_2757,N_2687);
and U3740 (N_3740,N_2629,N_2551);
nor U3741 (N_3741,N_1503,N_2136);
nor U3742 (N_3742,N_2962,N_2351);
or U3743 (N_3743,N_2805,N_1709);
nand U3744 (N_3744,N_1520,N_2255);
xor U3745 (N_3745,N_2167,N_2543);
xor U3746 (N_3746,N_2207,N_2530);
or U3747 (N_3747,N_2923,N_1752);
nand U3748 (N_3748,N_2576,N_1545);
or U3749 (N_3749,N_1934,N_2694);
xor U3750 (N_3750,N_2767,N_1716);
nor U3751 (N_3751,N_2612,N_2614);
nor U3752 (N_3752,N_2491,N_2719);
or U3753 (N_3753,N_2162,N_2723);
nor U3754 (N_3754,N_2796,N_2628);
xor U3755 (N_3755,N_2484,N_2786);
and U3756 (N_3756,N_1739,N_2772);
nor U3757 (N_3757,N_2482,N_2052);
xor U3758 (N_3758,N_2090,N_2368);
or U3759 (N_3759,N_1896,N_2272);
or U3760 (N_3760,N_1911,N_2293);
or U3761 (N_3761,N_2019,N_2244);
nor U3762 (N_3762,N_2233,N_2407);
and U3763 (N_3763,N_2733,N_1731);
or U3764 (N_3764,N_1821,N_1852);
xor U3765 (N_3765,N_1650,N_2079);
xor U3766 (N_3766,N_2435,N_2914);
or U3767 (N_3767,N_2858,N_1852);
and U3768 (N_3768,N_1644,N_2263);
nor U3769 (N_3769,N_2963,N_2925);
or U3770 (N_3770,N_1791,N_1970);
and U3771 (N_3771,N_2351,N_2008);
or U3772 (N_3772,N_2048,N_2018);
xor U3773 (N_3773,N_2657,N_2896);
xor U3774 (N_3774,N_2017,N_1618);
nand U3775 (N_3775,N_2275,N_2161);
and U3776 (N_3776,N_1761,N_1653);
xnor U3777 (N_3777,N_1720,N_1624);
and U3778 (N_3778,N_2739,N_2864);
nand U3779 (N_3779,N_1697,N_2175);
or U3780 (N_3780,N_1925,N_1540);
nor U3781 (N_3781,N_2116,N_1723);
or U3782 (N_3782,N_2280,N_1900);
nor U3783 (N_3783,N_1505,N_2641);
nand U3784 (N_3784,N_2366,N_1774);
and U3785 (N_3785,N_1743,N_2798);
nand U3786 (N_3786,N_1553,N_2661);
or U3787 (N_3787,N_2593,N_2019);
nor U3788 (N_3788,N_2821,N_2075);
nor U3789 (N_3789,N_1507,N_2574);
xnor U3790 (N_3790,N_1729,N_1658);
nor U3791 (N_3791,N_1508,N_1639);
and U3792 (N_3792,N_1882,N_2327);
nand U3793 (N_3793,N_2848,N_2190);
or U3794 (N_3794,N_1795,N_2037);
nand U3795 (N_3795,N_2377,N_2848);
nor U3796 (N_3796,N_1916,N_1561);
xor U3797 (N_3797,N_2161,N_2043);
nor U3798 (N_3798,N_2344,N_2995);
and U3799 (N_3799,N_1804,N_1583);
nor U3800 (N_3800,N_2085,N_1761);
nor U3801 (N_3801,N_2024,N_2833);
or U3802 (N_3802,N_2927,N_1648);
nand U3803 (N_3803,N_2917,N_2576);
nor U3804 (N_3804,N_2411,N_1838);
and U3805 (N_3805,N_1698,N_1625);
nor U3806 (N_3806,N_2794,N_1631);
nor U3807 (N_3807,N_2715,N_2682);
nor U3808 (N_3808,N_2251,N_1690);
xor U3809 (N_3809,N_1677,N_1997);
nor U3810 (N_3810,N_1548,N_2629);
nand U3811 (N_3811,N_2380,N_2948);
nor U3812 (N_3812,N_2477,N_2431);
nor U3813 (N_3813,N_1580,N_1628);
xnor U3814 (N_3814,N_2552,N_2835);
nor U3815 (N_3815,N_2739,N_1931);
nor U3816 (N_3816,N_2522,N_1568);
nor U3817 (N_3817,N_1734,N_2051);
or U3818 (N_3818,N_2277,N_2293);
nand U3819 (N_3819,N_2892,N_2870);
nand U3820 (N_3820,N_2957,N_2441);
xor U3821 (N_3821,N_1787,N_1830);
nand U3822 (N_3822,N_2949,N_2251);
nor U3823 (N_3823,N_2080,N_2554);
nand U3824 (N_3824,N_2772,N_2157);
and U3825 (N_3825,N_2793,N_2318);
nor U3826 (N_3826,N_2505,N_2807);
nand U3827 (N_3827,N_2489,N_2375);
nor U3828 (N_3828,N_2446,N_2560);
nand U3829 (N_3829,N_2029,N_2289);
xnor U3830 (N_3830,N_2226,N_2596);
and U3831 (N_3831,N_2652,N_1691);
xor U3832 (N_3832,N_1550,N_2290);
or U3833 (N_3833,N_2432,N_2475);
nor U3834 (N_3834,N_2224,N_2103);
nand U3835 (N_3835,N_2407,N_2935);
nand U3836 (N_3836,N_1881,N_1718);
nor U3837 (N_3837,N_2504,N_2446);
nor U3838 (N_3838,N_2716,N_2592);
and U3839 (N_3839,N_2091,N_1845);
nand U3840 (N_3840,N_1762,N_1862);
nand U3841 (N_3841,N_2085,N_2038);
nand U3842 (N_3842,N_1537,N_2949);
or U3843 (N_3843,N_2972,N_2874);
nand U3844 (N_3844,N_2688,N_1976);
xor U3845 (N_3845,N_2663,N_2601);
or U3846 (N_3846,N_2534,N_2384);
or U3847 (N_3847,N_2956,N_2225);
or U3848 (N_3848,N_2504,N_1509);
nor U3849 (N_3849,N_2214,N_2063);
nand U3850 (N_3850,N_2713,N_1890);
nor U3851 (N_3851,N_2746,N_2078);
nor U3852 (N_3852,N_2117,N_2174);
nand U3853 (N_3853,N_2177,N_1509);
nor U3854 (N_3854,N_2506,N_2730);
nor U3855 (N_3855,N_1753,N_1533);
xor U3856 (N_3856,N_1663,N_2628);
or U3857 (N_3857,N_2115,N_1694);
or U3858 (N_3858,N_2564,N_2159);
and U3859 (N_3859,N_1909,N_2645);
and U3860 (N_3860,N_1719,N_1933);
nand U3861 (N_3861,N_2675,N_2271);
or U3862 (N_3862,N_2974,N_1733);
xnor U3863 (N_3863,N_2439,N_2992);
nand U3864 (N_3864,N_2253,N_2797);
or U3865 (N_3865,N_1750,N_2252);
nor U3866 (N_3866,N_2060,N_2061);
nor U3867 (N_3867,N_1530,N_2477);
nor U3868 (N_3868,N_2721,N_1662);
xor U3869 (N_3869,N_1602,N_1579);
nand U3870 (N_3870,N_1805,N_2902);
or U3871 (N_3871,N_2548,N_2079);
and U3872 (N_3872,N_2285,N_2143);
nand U3873 (N_3873,N_2016,N_2079);
or U3874 (N_3874,N_1663,N_2423);
xor U3875 (N_3875,N_2451,N_2757);
nor U3876 (N_3876,N_2961,N_2316);
nand U3877 (N_3877,N_2909,N_2232);
nand U3878 (N_3878,N_1667,N_2193);
and U3879 (N_3879,N_2362,N_2591);
or U3880 (N_3880,N_2737,N_1805);
nor U3881 (N_3881,N_1820,N_1934);
xnor U3882 (N_3882,N_1681,N_2896);
xnor U3883 (N_3883,N_2199,N_2299);
nand U3884 (N_3884,N_2076,N_1521);
or U3885 (N_3885,N_2830,N_1644);
nand U3886 (N_3886,N_1838,N_1509);
nand U3887 (N_3887,N_2636,N_1563);
xor U3888 (N_3888,N_2726,N_2796);
nor U3889 (N_3889,N_1860,N_2511);
nand U3890 (N_3890,N_2499,N_2972);
nor U3891 (N_3891,N_2276,N_2944);
and U3892 (N_3892,N_1644,N_2581);
nand U3893 (N_3893,N_2272,N_1965);
or U3894 (N_3894,N_1545,N_2531);
or U3895 (N_3895,N_2370,N_2571);
xnor U3896 (N_3896,N_1677,N_2491);
and U3897 (N_3897,N_1823,N_2575);
nor U3898 (N_3898,N_1962,N_1928);
or U3899 (N_3899,N_2125,N_1767);
and U3900 (N_3900,N_1991,N_1923);
nand U3901 (N_3901,N_1611,N_2089);
nor U3902 (N_3902,N_1611,N_1793);
or U3903 (N_3903,N_2109,N_2251);
nor U3904 (N_3904,N_1873,N_1931);
xor U3905 (N_3905,N_1827,N_1591);
and U3906 (N_3906,N_2435,N_2811);
nor U3907 (N_3907,N_2454,N_2386);
nor U3908 (N_3908,N_1913,N_2269);
nand U3909 (N_3909,N_2657,N_2993);
nor U3910 (N_3910,N_2091,N_1756);
nand U3911 (N_3911,N_2522,N_2276);
nand U3912 (N_3912,N_1619,N_2461);
and U3913 (N_3913,N_2095,N_2421);
nor U3914 (N_3914,N_1821,N_2677);
nor U3915 (N_3915,N_2235,N_1693);
and U3916 (N_3916,N_1529,N_1734);
and U3917 (N_3917,N_2446,N_2285);
xor U3918 (N_3918,N_2513,N_1695);
and U3919 (N_3919,N_1614,N_2669);
and U3920 (N_3920,N_2652,N_1559);
and U3921 (N_3921,N_1534,N_2570);
or U3922 (N_3922,N_2309,N_2333);
or U3923 (N_3923,N_1774,N_1950);
or U3924 (N_3924,N_1988,N_2165);
nor U3925 (N_3925,N_2668,N_2231);
xnor U3926 (N_3926,N_1536,N_1712);
and U3927 (N_3927,N_1595,N_2549);
xnor U3928 (N_3928,N_2376,N_2100);
nand U3929 (N_3929,N_1922,N_2240);
xor U3930 (N_3930,N_2394,N_2209);
or U3931 (N_3931,N_1684,N_2148);
nor U3932 (N_3932,N_1810,N_1984);
nor U3933 (N_3933,N_2917,N_2313);
or U3934 (N_3934,N_2620,N_2963);
and U3935 (N_3935,N_1917,N_2126);
or U3936 (N_3936,N_2794,N_2544);
nor U3937 (N_3937,N_2026,N_2108);
xor U3938 (N_3938,N_2126,N_2719);
xnor U3939 (N_3939,N_1772,N_1950);
and U3940 (N_3940,N_2314,N_2530);
xnor U3941 (N_3941,N_2811,N_2515);
nand U3942 (N_3942,N_2055,N_2121);
nand U3943 (N_3943,N_2381,N_2244);
nand U3944 (N_3944,N_1686,N_2968);
xor U3945 (N_3945,N_2609,N_1704);
nor U3946 (N_3946,N_2251,N_1842);
and U3947 (N_3947,N_1532,N_2694);
xor U3948 (N_3948,N_2893,N_1652);
and U3949 (N_3949,N_2905,N_2753);
nor U3950 (N_3950,N_2596,N_1820);
xor U3951 (N_3951,N_2760,N_2453);
and U3952 (N_3952,N_2072,N_2043);
nor U3953 (N_3953,N_1714,N_1948);
nand U3954 (N_3954,N_2375,N_2295);
or U3955 (N_3955,N_2933,N_2813);
nand U3956 (N_3956,N_2637,N_2499);
nand U3957 (N_3957,N_2937,N_1775);
nor U3958 (N_3958,N_1866,N_2084);
nor U3959 (N_3959,N_2338,N_2428);
nor U3960 (N_3960,N_2387,N_2908);
nand U3961 (N_3961,N_2901,N_2844);
or U3962 (N_3962,N_2946,N_2534);
or U3963 (N_3963,N_2434,N_1924);
or U3964 (N_3964,N_2763,N_2683);
nand U3965 (N_3965,N_1921,N_2994);
or U3966 (N_3966,N_2572,N_2990);
and U3967 (N_3967,N_2836,N_2475);
and U3968 (N_3968,N_2119,N_2744);
nand U3969 (N_3969,N_2350,N_1510);
nor U3970 (N_3970,N_2989,N_2869);
or U3971 (N_3971,N_1724,N_2172);
and U3972 (N_3972,N_1532,N_2338);
nor U3973 (N_3973,N_2409,N_2741);
nor U3974 (N_3974,N_2986,N_2213);
and U3975 (N_3975,N_1651,N_2079);
xnor U3976 (N_3976,N_2553,N_2587);
and U3977 (N_3977,N_1802,N_2217);
and U3978 (N_3978,N_2890,N_1537);
xor U3979 (N_3979,N_1763,N_2063);
and U3980 (N_3980,N_2323,N_1552);
nor U3981 (N_3981,N_1962,N_1992);
nand U3982 (N_3982,N_1578,N_2562);
and U3983 (N_3983,N_1618,N_2960);
and U3984 (N_3984,N_2810,N_2663);
and U3985 (N_3985,N_2908,N_2452);
nor U3986 (N_3986,N_1950,N_1717);
nand U3987 (N_3987,N_2645,N_1902);
xor U3988 (N_3988,N_1872,N_2730);
nand U3989 (N_3989,N_2423,N_2982);
nor U3990 (N_3990,N_2130,N_2662);
and U3991 (N_3991,N_2293,N_1686);
nand U3992 (N_3992,N_2308,N_2110);
and U3993 (N_3993,N_1978,N_1719);
xor U3994 (N_3994,N_2010,N_2185);
xnor U3995 (N_3995,N_2119,N_1754);
xor U3996 (N_3996,N_2436,N_2371);
and U3997 (N_3997,N_2555,N_2217);
nand U3998 (N_3998,N_1713,N_2236);
or U3999 (N_3999,N_2565,N_2132);
and U4000 (N_4000,N_1567,N_2978);
xnor U4001 (N_4001,N_2657,N_2315);
nand U4002 (N_4002,N_2428,N_2794);
xor U4003 (N_4003,N_2729,N_1651);
nand U4004 (N_4004,N_2231,N_1891);
xor U4005 (N_4005,N_1739,N_1831);
nand U4006 (N_4006,N_1525,N_2861);
xnor U4007 (N_4007,N_1635,N_2491);
xnor U4008 (N_4008,N_1806,N_2679);
or U4009 (N_4009,N_2754,N_2093);
or U4010 (N_4010,N_1769,N_2449);
xnor U4011 (N_4011,N_2849,N_1673);
nor U4012 (N_4012,N_2925,N_2947);
nand U4013 (N_4013,N_2277,N_1704);
nand U4014 (N_4014,N_2112,N_1647);
or U4015 (N_4015,N_2207,N_2554);
or U4016 (N_4016,N_2022,N_2232);
and U4017 (N_4017,N_2196,N_2207);
or U4018 (N_4018,N_2562,N_1709);
nor U4019 (N_4019,N_2558,N_2708);
nand U4020 (N_4020,N_1598,N_2801);
or U4021 (N_4021,N_1993,N_2515);
or U4022 (N_4022,N_2288,N_2618);
xnor U4023 (N_4023,N_1625,N_2349);
nand U4024 (N_4024,N_2333,N_1870);
nand U4025 (N_4025,N_2640,N_2424);
or U4026 (N_4026,N_2255,N_1935);
xnor U4027 (N_4027,N_2175,N_2467);
nand U4028 (N_4028,N_1838,N_1574);
nor U4029 (N_4029,N_1801,N_1785);
nand U4030 (N_4030,N_2649,N_1691);
nand U4031 (N_4031,N_2611,N_2351);
nor U4032 (N_4032,N_1587,N_2922);
nand U4033 (N_4033,N_1669,N_2203);
xnor U4034 (N_4034,N_2832,N_2457);
or U4035 (N_4035,N_1755,N_2731);
nor U4036 (N_4036,N_2933,N_2486);
nor U4037 (N_4037,N_2477,N_1784);
xnor U4038 (N_4038,N_2578,N_2693);
or U4039 (N_4039,N_2571,N_2772);
and U4040 (N_4040,N_1809,N_1739);
or U4041 (N_4041,N_2262,N_1596);
and U4042 (N_4042,N_1881,N_2483);
and U4043 (N_4043,N_1807,N_2946);
and U4044 (N_4044,N_2360,N_2905);
and U4045 (N_4045,N_2053,N_2618);
nand U4046 (N_4046,N_2570,N_2342);
nand U4047 (N_4047,N_1898,N_2992);
nor U4048 (N_4048,N_2399,N_2767);
xor U4049 (N_4049,N_1638,N_1608);
nand U4050 (N_4050,N_2135,N_2974);
xnor U4051 (N_4051,N_1697,N_2610);
and U4052 (N_4052,N_2188,N_2916);
xnor U4053 (N_4053,N_2214,N_2837);
nand U4054 (N_4054,N_1724,N_2322);
xor U4055 (N_4055,N_2045,N_2463);
xnor U4056 (N_4056,N_2045,N_1742);
xor U4057 (N_4057,N_2698,N_1708);
nor U4058 (N_4058,N_2358,N_2885);
nor U4059 (N_4059,N_1702,N_2591);
nor U4060 (N_4060,N_2397,N_1823);
xor U4061 (N_4061,N_2472,N_2884);
xnor U4062 (N_4062,N_2705,N_1724);
nand U4063 (N_4063,N_1868,N_2344);
or U4064 (N_4064,N_2651,N_2548);
xnor U4065 (N_4065,N_2854,N_2666);
and U4066 (N_4066,N_2005,N_1938);
nor U4067 (N_4067,N_2405,N_1729);
xnor U4068 (N_4068,N_1592,N_2213);
or U4069 (N_4069,N_1931,N_2853);
nand U4070 (N_4070,N_2269,N_2746);
nor U4071 (N_4071,N_1921,N_2047);
and U4072 (N_4072,N_1545,N_2501);
or U4073 (N_4073,N_2241,N_1710);
nand U4074 (N_4074,N_2579,N_2881);
nand U4075 (N_4075,N_1788,N_2028);
and U4076 (N_4076,N_1982,N_2820);
nor U4077 (N_4077,N_2822,N_2492);
nand U4078 (N_4078,N_2435,N_2021);
or U4079 (N_4079,N_2783,N_1586);
or U4080 (N_4080,N_2502,N_2134);
xor U4081 (N_4081,N_2788,N_1557);
or U4082 (N_4082,N_2196,N_2914);
and U4083 (N_4083,N_2864,N_2403);
or U4084 (N_4084,N_2786,N_2424);
nand U4085 (N_4085,N_2870,N_2203);
xor U4086 (N_4086,N_2701,N_2502);
and U4087 (N_4087,N_2842,N_1752);
or U4088 (N_4088,N_2496,N_2233);
and U4089 (N_4089,N_2569,N_1955);
xor U4090 (N_4090,N_2459,N_2366);
and U4091 (N_4091,N_2654,N_2203);
xor U4092 (N_4092,N_2762,N_2461);
and U4093 (N_4093,N_2809,N_1652);
and U4094 (N_4094,N_1675,N_1729);
or U4095 (N_4095,N_1605,N_2964);
or U4096 (N_4096,N_1549,N_1856);
and U4097 (N_4097,N_1558,N_1589);
nor U4098 (N_4098,N_2115,N_2801);
nor U4099 (N_4099,N_2793,N_2118);
and U4100 (N_4100,N_2560,N_2379);
nand U4101 (N_4101,N_2576,N_1990);
and U4102 (N_4102,N_1847,N_1991);
and U4103 (N_4103,N_1838,N_2324);
or U4104 (N_4104,N_1751,N_1569);
or U4105 (N_4105,N_2798,N_1653);
xnor U4106 (N_4106,N_2757,N_2889);
nor U4107 (N_4107,N_2070,N_2593);
and U4108 (N_4108,N_2674,N_2280);
or U4109 (N_4109,N_2711,N_2029);
or U4110 (N_4110,N_2982,N_2809);
nor U4111 (N_4111,N_2778,N_2182);
xnor U4112 (N_4112,N_2930,N_2349);
nand U4113 (N_4113,N_2021,N_2774);
and U4114 (N_4114,N_1691,N_2911);
and U4115 (N_4115,N_2969,N_1552);
nand U4116 (N_4116,N_2843,N_2421);
or U4117 (N_4117,N_1871,N_2726);
and U4118 (N_4118,N_2402,N_2396);
nand U4119 (N_4119,N_1862,N_2455);
and U4120 (N_4120,N_1694,N_1850);
nor U4121 (N_4121,N_2857,N_2891);
or U4122 (N_4122,N_2585,N_2664);
nor U4123 (N_4123,N_1778,N_2692);
nor U4124 (N_4124,N_2605,N_2000);
nand U4125 (N_4125,N_1655,N_2096);
and U4126 (N_4126,N_2414,N_2109);
nor U4127 (N_4127,N_2495,N_1797);
or U4128 (N_4128,N_2848,N_2821);
or U4129 (N_4129,N_1879,N_1932);
and U4130 (N_4130,N_2833,N_1954);
nand U4131 (N_4131,N_1720,N_2411);
xnor U4132 (N_4132,N_1829,N_2318);
and U4133 (N_4133,N_2944,N_1985);
and U4134 (N_4134,N_2844,N_2214);
or U4135 (N_4135,N_1527,N_1547);
or U4136 (N_4136,N_1905,N_1763);
and U4137 (N_4137,N_2587,N_1888);
xor U4138 (N_4138,N_2678,N_2346);
nand U4139 (N_4139,N_2153,N_1558);
nand U4140 (N_4140,N_2570,N_2991);
and U4141 (N_4141,N_2806,N_2695);
nor U4142 (N_4142,N_2262,N_1817);
nor U4143 (N_4143,N_1862,N_2382);
or U4144 (N_4144,N_2630,N_2350);
xnor U4145 (N_4145,N_1635,N_2501);
nand U4146 (N_4146,N_2234,N_2544);
xnor U4147 (N_4147,N_2234,N_2547);
nor U4148 (N_4148,N_2852,N_2105);
or U4149 (N_4149,N_2200,N_1589);
and U4150 (N_4150,N_2593,N_1695);
nand U4151 (N_4151,N_1977,N_1523);
nand U4152 (N_4152,N_2209,N_1994);
nor U4153 (N_4153,N_1832,N_1617);
or U4154 (N_4154,N_1508,N_2318);
nor U4155 (N_4155,N_2125,N_2669);
xnor U4156 (N_4156,N_2336,N_1832);
xnor U4157 (N_4157,N_2011,N_2617);
and U4158 (N_4158,N_2291,N_2978);
xor U4159 (N_4159,N_2125,N_2914);
nor U4160 (N_4160,N_2865,N_2155);
or U4161 (N_4161,N_1881,N_2482);
or U4162 (N_4162,N_2420,N_2961);
nor U4163 (N_4163,N_2271,N_1950);
or U4164 (N_4164,N_1786,N_2006);
nor U4165 (N_4165,N_2895,N_2608);
or U4166 (N_4166,N_2086,N_1767);
or U4167 (N_4167,N_1568,N_2634);
nor U4168 (N_4168,N_2203,N_2883);
nand U4169 (N_4169,N_2406,N_2648);
nand U4170 (N_4170,N_1765,N_1797);
nor U4171 (N_4171,N_1853,N_2237);
nand U4172 (N_4172,N_1939,N_2641);
or U4173 (N_4173,N_2566,N_2922);
and U4174 (N_4174,N_1942,N_2127);
or U4175 (N_4175,N_1936,N_2821);
or U4176 (N_4176,N_2948,N_2960);
and U4177 (N_4177,N_2729,N_2478);
nor U4178 (N_4178,N_1939,N_2623);
xor U4179 (N_4179,N_1851,N_1730);
nand U4180 (N_4180,N_2965,N_2474);
and U4181 (N_4181,N_2849,N_1758);
or U4182 (N_4182,N_2920,N_2006);
and U4183 (N_4183,N_1519,N_1796);
nor U4184 (N_4184,N_1764,N_2489);
or U4185 (N_4185,N_2326,N_2193);
and U4186 (N_4186,N_1684,N_2759);
nor U4187 (N_4187,N_1794,N_2041);
xor U4188 (N_4188,N_2314,N_2012);
or U4189 (N_4189,N_1908,N_1870);
or U4190 (N_4190,N_2034,N_2928);
xnor U4191 (N_4191,N_2003,N_2259);
and U4192 (N_4192,N_2202,N_2762);
nand U4193 (N_4193,N_2176,N_1630);
xor U4194 (N_4194,N_2674,N_2652);
nand U4195 (N_4195,N_2067,N_1820);
xnor U4196 (N_4196,N_1517,N_1513);
nand U4197 (N_4197,N_1836,N_1501);
nand U4198 (N_4198,N_1773,N_2686);
or U4199 (N_4199,N_1813,N_1861);
nor U4200 (N_4200,N_2120,N_2700);
nor U4201 (N_4201,N_2823,N_2336);
xnor U4202 (N_4202,N_1969,N_2472);
xor U4203 (N_4203,N_2412,N_2039);
or U4204 (N_4204,N_2117,N_2634);
nor U4205 (N_4205,N_2817,N_2062);
nor U4206 (N_4206,N_1721,N_2641);
xor U4207 (N_4207,N_2946,N_2107);
nor U4208 (N_4208,N_1676,N_2936);
nor U4209 (N_4209,N_2588,N_2695);
or U4210 (N_4210,N_2327,N_2393);
and U4211 (N_4211,N_2698,N_1525);
or U4212 (N_4212,N_2474,N_2163);
xor U4213 (N_4213,N_2704,N_1626);
or U4214 (N_4214,N_2303,N_1678);
nor U4215 (N_4215,N_2802,N_2139);
xor U4216 (N_4216,N_2811,N_2775);
nand U4217 (N_4217,N_2258,N_1611);
and U4218 (N_4218,N_2859,N_2714);
or U4219 (N_4219,N_2347,N_1616);
and U4220 (N_4220,N_2169,N_1909);
or U4221 (N_4221,N_1516,N_2662);
nand U4222 (N_4222,N_2404,N_2083);
xnor U4223 (N_4223,N_2637,N_1812);
nor U4224 (N_4224,N_2968,N_2754);
or U4225 (N_4225,N_1839,N_1504);
nand U4226 (N_4226,N_2885,N_1622);
nand U4227 (N_4227,N_2440,N_1914);
nand U4228 (N_4228,N_2854,N_2844);
or U4229 (N_4229,N_2339,N_2945);
and U4230 (N_4230,N_1671,N_2212);
or U4231 (N_4231,N_2685,N_2287);
xnor U4232 (N_4232,N_2933,N_2935);
or U4233 (N_4233,N_1870,N_1896);
nor U4234 (N_4234,N_2059,N_2692);
nand U4235 (N_4235,N_2103,N_2845);
nor U4236 (N_4236,N_1807,N_2714);
or U4237 (N_4237,N_2548,N_2364);
and U4238 (N_4238,N_2867,N_2070);
and U4239 (N_4239,N_2778,N_2753);
xnor U4240 (N_4240,N_2125,N_2795);
or U4241 (N_4241,N_1708,N_2708);
nor U4242 (N_4242,N_2030,N_1910);
and U4243 (N_4243,N_2926,N_2917);
or U4244 (N_4244,N_1761,N_2161);
or U4245 (N_4245,N_1572,N_2056);
xnor U4246 (N_4246,N_2374,N_1518);
nor U4247 (N_4247,N_1558,N_2360);
and U4248 (N_4248,N_1833,N_1531);
or U4249 (N_4249,N_1932,N_2376);
nor U4250 (N_4250,N_2894,N_1837);
nand U4251 (N_4251,N_2568,N_1980);
and U4252 (N_4252,N_2321,N_2312);
nand U4253 (N_4253,N_2757,N_1643);
or U4254 (N_4254,N_2563,N_2203);
or U4255 (N_4255,N_2538,N_2254);
xnor U4256 (N_4256,N_1665,N_2667);
xor U4257 (N_4257,N_2897,N_1891);
xor U4258 (N_4258,N_2393,N_1993);
or U4259 (N_4259,N_1610,N_2559);
nand U4260 (N_4260,N_2932,N_2541);
nor U4261 (N_4261,N_1573,N_1959);
nor U4262 (N_4262,N_2936,N_1726);
nand U4263 (N_4263,N_2362,N_2306);
xnor U4264 (N_4264,N_2206,N_1857);
nand U4265 (N_4265,N_2383,N_1554);
or U4266 (N_4266,N_2918,N_2155);
nand U4267 (N_4267,N_2050,N_2092);
nor U4268 (N_4268,N_1702,N_2652);
xor U4269 (N_4269,N_1593,N_1968);
and U4270 (N_4270,N_2465,N_2449);
or U4271 (N_4271,N_2956,N_2541);
nor U4272 (N_4272,N_1775,N_2128);
and U4273 (N_4273,N_1739,N_2770);
nor U4274 (N_4274,N_2814,N_1898);
nor U4275 (N_4275,N_2268,N_1919);
or U4276 (N_4276,N_2985,N_2798);
and U4277 (N_4277,N_1915,N_2739);
nand U4278 (N_4278,N_2900,N_1809);
nand U4279 (N_4279,N_2718,N_2863);
and U4280 (N_4280,N_1781,N_2450);
or U4281 (N_4281,N_2975,N_1996);
or U4282 (N_4282,N_2765,N_2944);
nand U4283 (N_4283,N_2072,N_2921);
or U4284 (N_4284,N_2192,N_2755);
or U4285 (N_4285,N_2053,N_2784);
xor U4286 (N_4286,N_2296,N_1641);
or U4287 (N_4287,N_2585,N_1805);
xor U4288 (N_4288,N_2499,N_2140);
or U4289 (N_4289,N_2022,N_1688);
nand U4290 (N_4290,N_2599,N_2481);
or U4291 (N_4291,N_2745,N_1691);
and U4292 (N_4292,N_2034,N_1515);
or U4293 (N_4293,N_2790,N_2582);
nand U4294 (N_4294,N_2547,N_1865);
and U4295 (N_4295,N_1651,N_1659);
nand U4296 (N_4296,N_2290,N_2011);
and U4297 (N_4297,N_2123,N_2354);
and U4298 (N_4298,N_2497,N_2486);
xor U4299 (N_4299,N_1898,N_2253);
or U4300 (N_4300,N_2742,N_1722);
nand U4301 (N_4301,N_1970,N_2466);
nor U4302 (N_4302,N_1565,N_2937);
nand U4303 (N_4303,N_1595,N_2652);
nand U4304 (N_4304,N_1557,N_2655);
nor U4305 (N_4305,N_2192,N_2088);
xnor U4306 (N_4306,N_2309,N_2782);
and U4307 (N_4307,N_1557,N_1696);
nand U4308 (N_4308,N_1793,N_1829);
nand U4309 (N_4309,N_2553,N_1730);
xor U4310 (N_4310,N_2986,N_1833);
nor U4311 (N_4311,N_1896,N_2409);
or U4312 (N_4312,N_2594,N_2354);
and U4313 (N_4313,N_1958,N_2231);
or U4314 (N_4314,N_2408,N_1909);
and U4315 (N_4315,N_2696,N_2399);
xor U4316 (N_4316,N_1699,N_2117);
nand U4317 (N_4317,N_1538,N_2205);
nand U4318 (N_4318,N_1748,N_1521);
and U4319 (N_4319,N_2949,N_1682);
or U4320 (N_4320,N_2426,N_2870);
xor U4321 (N_4321,N_2944,N_2086);
and U4322 (N_4322,N_2985,N_2524);
nand U4323 (N_4323,N_2235,N_2731);
nand U4324 (N_4324,N_1805,N_1896);
xor U4325 (N_4325,N_2615,N_1895);
and U4326 (N_4326,N_1739,N_2851);
nand U4327 (N_4327,N_2528,N_2090);
nor U4328 (N_4328,N_2198,N_2393);
xor U4329 (N_4329,N_2269,N_2251);
xnor U4330 (N_4330,N_2535,N_2167);
xor U4331 (N_4331,N_2641,N_1999);
and U4332 (N_4332,N_2187,N_1501);
xnor U4333 (N_4333,N_1568,N_1888);
or U4334 (N_4334,N_1507,N_2436);
nor U4335 (N_4335,N_2885,N_1710);
and U4336 (N_4336,N_2607,N_2492);
xor U4337 (N_4337,N_2919,N_1517);
xor U4338 (N_4338,N_2206,N_2943);
nor U4339 (N_4339,N_1789,N_2802);
or U4340 (N_4340,N_2312,N_2440);
xor U4341 (N_4341,N_1851,N_2599);
or U4342 (N_4342,N_2369,N_1977);
xor U4343 (N_4343,N_2476,N_2212);
nor U4344 (N_4344,N_2521,N_1664);
nor U4345 (N_4345,N_1990,N_2142);
and U4346 (N_4346,N_2482,N_2544);
or U4347 (N_4347,N_2382,N_2187);
nand U4348 (N_4348,N_2840,N_2352);
and U4349 (N_4349,N_2462,N_2508);
or U4350 (N_4350,N_2693,N_2256);
nor U4351 (N_4351,N_1570,N_1775);
nor U4352 (N_4352,N_1530,N_1669);
and U4353 (N_4353,N_2936,N_2170);
nor U4354 (N_4354,N_2883,N_2284);
nor U4355 (N_4355,N_2215,N_2203);
and U4356 (N_4356,N_2219,N_2636);
nand U4357 (N_4357,N_2176,N_2922);
nor U4358 (N_4358,N_2647,N_1737);
xor U4359 (N_4359,N_1837,N_2365);
xnor U4360 (N_4360,N_1798,N_2270);
or U4361 (N_4361,N_2631,N_1878);
nand U4362 (N_4362,N_1902,N_2703);
and U4363 (N_4363,N_2875,N_1849);
nor U4364 (N_4364,N_2111,N_2754);
nand U4365 (N_4365,N_2905,N_1733);
nor U4366 (N_4366,N_2468,N_2014);
xor U4367 (N_4367,N_1628,N_2436);
nor U4368 (N_4368,N_2825,N_1843);
and U4369 (N_4369,N_2835,N_2192);
nand U4370 (N_4370,N_2607,N_2347);
nand U4371 (N_4371,N_2409,N_2022);
xor U4372 (N_4372,N_2304,N_1856);
or U4373 (N_4373,N_1996,N_1944);
nor U4374 (N_4374,N_1674,N_1847);
nor U4375 (N_4375,N_2305,N_2757);
nor U4376 (N_4376,N_2535,N_2458);
nand U4377 (N_4377,N_1564,N_2575);
and U4378 (N_4378,N_1788,N_2452);
nand U4379 (N_4379,N_2157,N_1812);
xnor U4380 (N_4380,N_2966,N_2691);
nor U4381 (N_4381,N_2515,N_2665);
or U4382 (N_4382,N_2056,N_2920);
and U4383 (N_4383,N_2590,N_1887);
or U4384 (N_4384,N_2711,N_2765);
and U4385 (N_4385,N_2326,N_2032);
or U4386 (N_4386,N_2216,N_2350);
and U4387 (N_4387,N_2641,N_2632);
nor U4388 (N_4388,N_1831,N_1656);
nor U4389 (N_4389,N_2071,N_2206);
nor U4390 (N_4390,N_1938,N_2214);
or U4391 (N_4391,N_2615,N_2703);
nand U4392 (N_4392,N_2331,N_2567);
nand U4393 (N_4393,N_2623,N_1976);
xor U4394 (N_4394,N_2956,N_2479);
or U4395 (N_4395,N_2321,N_1786);
nand U4396 (N_4396,N_2431,N_2809);
nand U4397 (N_4397,N_2115,N_2334);
or U4398 (N_4398,N_2337,N_2219);
nand U4399 (N_4399,N_1647,N_2994);
or U4400 (N_4400,N_2042,N_1947);
or U4401 (N_4401,N_2399,N_1708);
nand U4402 (N_4402,N_2071,N_2162);
nor U4403 (N_4403,N_2117,N_2988);
nand U4404 (N_4404,N_2488,N_2061);
and U4405 (N_4405,N_2509,N_2641);
nand U4406 (N_4406,N_2669,N_1919);
nor U4407 (N_4407,N_2120,N_1628);
nor U4408 (N_4408,N_2899,N_2194);
xnor U4409 (N_4409,N_1573,N_1761);
nand U4410 (N_4410,N_1808,N_2458);
and U4411 (N_4411,N_2117,N_1864);
nand U4412 (N_4412,N_2231,N_1860);
and U4413 (N_4413,N_2960,N_2711);
or U4414 (N_4414,N_2071,N_1618);
or U4415 (N_4415,N_2812,N_2640);
nor U4416 (N_4416,N_1866,N_2738);
and U4417 (N_4417,N_2243,N_1900);
or U4418 (N_4418,N_2207,N_1645);
or U4419 (N_4419,N_2154,N_2593);
or U4420 (N_4420,N_1726,N_1865);
xor U4421 (N_4421,N_2674,N_1942);
xor U4422 (N_4422,N_1808,N_1955);
nor U4423 (N_4423,N_2325,N_2489);
and U4424 (N_4424,N_2639,N_1782);
nor U4425 (N_4425,N_2804,N_2820);
nor U4426 (N_4426,N_2043,N_2789);
xor U4427 (N_4427,N_1641,N_2333);
and U4428 (N_4428,N_2764,N_1779);
and U4429 (N_4429,N_1908,N_1682);
or U4430 (N_4430,N_2710,N_2222);
nand U4431 (N_4431,N_1503,N_2105);
xor U4432 (N_4432,N_2127,N_2654);
or U4433 (N_4433,N_2821,N_1532);
nand U4434 (N_4434,N_1597,N_1992);
xnor U4435 (N_4435,N_1926,N_1789);
nor U4436 (N_4436,N_2213,N_2970);
nor U4437 (N_4437,N_1656,N_1904);
nand U4438 (N_4438,N_1854,N_2460);
nor U4439 (N_4439,N_1654,N_1738);
or U4440 (N_4440,N_1575,N_2657);
nand U4441 (N_4441,N_1798,N_2840);
nor U4442 (N_4442,N_2803,N_2667);
xnor U4443 (N_4443,N_2666,N_1518);
nand U4444 (N_4444,N_2273,N_1939);
and U4445 (N_4445,N_2751,N_2544);
and U4446 (N_4446,N_2582,N_2249);
and U4447 (N_4447,N_2247,N_2809);
or U4448 (N_4448,N_2856,N_2961);
xor U4449 (N_4449,N_1556,N_2223);
and U4450 (N_4450,N_2087,N_2127);
nand U4451 (N_4451,N_2467,N_2061);
and U4452 (N_4452,N_2972,N_1700);
or U4453 (N_4453,N_2133,N_2878);
nor U4454 (N_4454,N_1563,N_2124);
and U4455 (N_4455,N_2976,N_2311);
nand U4456 (N_4456,N_2716,N_2933);
or U4457 (N_4457,N_2834,N_1829);
or U4458 (N_4458,N_2114,N_2752);
nor U4459 (N_4459,N_1789,N_2745);
or U4460 (N_4460,N_2570,N_2273);
nand U4461 (N_4461,N_2718,N_2238);
nand U4462 (N_4462,N_2674,N_2858);
nor U4463 (N_4463,N_1844,N_2307);
nor U4464 (N_4464,N_1814,N_2691);
nand U4465 (N_4465,N_1787,N_2028);
or U4466 (N_4466,N_1964,N_2911);
nand U4467 (N_4467,N_1747,N_1991);
nor U4468 (N_4468,N_1532,N_1675);
nand U4469 (N_4469,N_1548,N_1706);
and U4470 (N_4470,N_2744,N_2285);
nand U4471 (N_4471,N_2215,N_1706);
xnor U4472 (N_4472,N_1861,N_1720);
nand U4473 (N_4473,N_1954,N_1966);
nand U4474 (N_4474,N_1793,N_2418);
or U4475 (N_4475,N_2458,N_2983);
or U4476 (N_4476,N_2692,N_1619);
and U4477 (N_4477,N_2390,N_1650);
nor U4478 (N_4478,N_1757,N_2213);
nand U4479 (N_4479,N_2301,N_2093);
nand U4480 (N_4480,N_1872,N_2446);
xor U4481 (N_4481,N_2751,N_2464);
nand U4482 (N_4482,N_1658,N_2987);
nor U4483 (N_4483,N_2705,N_1754);
nor U4484 (N_4484,N_2377,N_2504);
nand U4485 (N_4485,N_1898,N_2302);
and U4486 (N_4486,N_1731,N_2379);
nor U4487 (N_4487,N_1591,N_1638);
xor U4488 (N_4488,N_2670,N_2586);
xor U4489 (N_4489,N_2295,N_2798);
nor U4490 (N_4490,N_1781,N_1899);
xnor U4491 (N_4491,N_1985,N_1582);
and U4492 (N_4492,N_2421,N_1902);
or U4493 (N_4493,N_2151,N_2323);
nor U4494 (N_4494,N_1870,N_1561);
or U4495 (N_4495,N_1992,N_2349);
nor U4496 (N_4496,N_2512,N_2524);
and U4497 (N_4497,N_2488,N_2625);
xnor U4498 (N_4498,N_2748,N_1546);
or U4499 (N_4499,N_2548,N_2049);
nand U4500 (N_4500,N_3308,N_4128);
xnor U4501 (N_4501,N_4462,N_4029);
nand U4502 (N_4502,N_4368,N_4136);
xor U4503 (N_4503,N_3083,N_4240);
nor U4504 (N_4504,N_4168,N_3655);
nand U4505 (N_4505,N_3850,N_3679);
or U4506 (N_4506,N_4272,N_3234);
nor U4507 (N_4507,N_3390,N_4409);
or U4508 (N_4508,N_3082,N_3859);
or U4509 (N_4509,N_4092,N_3558);
nor U4510 (N_4510,N_3989,N_3452);
nand U4511 (N_4511,N_3907,N_3775);
and U4512 (N_4512,N_4487,N_3335);
and U4513 (N_4513,N_3355,N_3835);
and U4514 (N_4514,N_3577,N_3170);
and U4515 (N_4515,N_4347,N_3372);
or U4516 (N_4516,N_3641,N_3579);
nand U4517 (N_4517,N_4359,N_3305);
and U4518 (N_4518,N_3793,N_3794);
nand U4519 (N_4519,N_4423,N_3988);
or U4520 (N_4520,N_3976,N_3779);
xnor U4521 (N_4521,N_3387,N_3936);
xnor U4522 (N_4522,N_4155,N_3391);
nand U4523 (N_4523,N_3683,N_4179);
nand U4524 (N_4524,N_3913,N_3172);
nor U4525 (N_4525,N_4342,N_3499);
or U4526 (N_4526,N_3445,N_3951);
xnor U4527 (N_4527,N_4331,N_4356);
nor U4528 (N_4528,N_3408,N_3104);
nor U4529 (N_4529,N_3118,N_3857);
and U4530 (N_4530,N_3903,N_3381);
nor U4531 (N_4531,N_3868,N_3155);
nor U4532 (N_4532,N_3882,N_3266);
xnor U4533 (N_4533,N_3371,N_3418);
and U4534 (N_4534,N_3311,N_4332);
xnor U4535 (N_4535,N_4123,N_4137);
nand U4536 (N_4536,N_3941,N_3776);
nand U4537 (N_4537,N_3502,N_3191);
xor U4538 (N_4538,N_3316,N_4183);
xor U4539 (N_4539,N_4420,N_3331);
xor U4540 (N_4540,N_3040,N_3759);
and U4541 (N_4541,N_3484,N_3497);
nand U4542 (N_4542,N_3001,N_4158);
nand U4543 (N_4543,N_3678,N_3132);
and U4544 (N_4544,N_3275,N_3545);
xor U4545 (N_4545,N_3238,N_3341);
or U4546 (N_4546,N_3627,N_3127);
xnor U4547 (N_4547,N_3973,N_3550);
nand U4548 (N_4548,N_4387,N_3872);
nor U4549 (N_4549,N_4341,N_3726);
xor U4550 (N_4550,N_4232,N_4204);
nand U4551 (N_4551,N_4460,N_4153);
or U4552 (N_4552,N_3061,N_3760);
nor U4553 (N_4553,N_4004,N_3405);
nand U4554 (N_4554,N_3221,N_3450);
or U4555 (N_4555,N_3303,N_3855);
or U4556 (N_4556,N_3599,N_3350);
xnor U4557 (N_4557,N_3301,N_3232);
and U4558 (N_4558,N_3620,N_3159);
nand U4559 (N_4559,N_3917,N_3531);
or U4560 (N_4560,N_3516,N_3644);
and U4561 (N_4561,N_3729,N_3832);
nand U4562 (N_4562,N_3697,N_4126);
and U4563 (N_4563,N_4038,N_3789);
nand U4564 (N_4564,N_4060,N_3330);
or U4565 (N_4565,N_4122,N_4378);
nand U4566 (N_4566,N_3160,N_3097);
xnor U4567 (N_4567,N_4262,N_3542);
nor U4568 (N_4568,N_4250,N_3431);
or U4569 (N_4569,N_3648,N_3087);
nand U4570 (N_4570,N_3947,N_3465);
and U4571 (N_4571,N_3652,N_3970);
and U4572 (N_4572,N_3909,N_3777);
and U4573 (N_4573,N_3313,N_3685);
nor U4574 (N_4574,N_3753,N_3161);
nor U4575 (N_4575,N_4100,N_3660);
xor U4576 (N_4576,N_3119,N_3805);
or U4577 (N_4577,N_3203,N_3126);
nand U4578 (N_4578,N_3877,N_4256);
or U4579 (N_4579,N_4129,N_3990);
nor U4580 (N_4580,N_3011,N_4241);
xor U4581 (N_4581,N_3133,N_3716);
and U4582 (N_4582,N_4434,N_4018);
nor U4583 (N_4583,N_4468,N_3862);
xnor U4584 (N_4584,N_4292,N_4380);
or U4585 (N_4585,N_3427,N_4353);
xor U4586 (N_4586,N_4303,N_3441);
or U4587 (N_4587,N_3731,N_3264);
nand U4588 (N_4588,N_3458,N_4194);
nand U4589 (N_4589,N_3763,N_4216);
xnor U4590 (N_4590,N_3267,N_4473);
nor U4591 (N_4591,N_4389,N_3103);
and U4592 (N_4592,N_4152,N_4217);
or U4593 (N_4593,N_4480,N_3404);
nor U4594 (N_4594,N_4317,N_3704);
nor U4595 (N_4595,N_3256,N_3826);
and U4596 (N_4596,N_3538,N_3927);
or U4597 (N_4597,N_3676,N_3474);
and U4598 (N_4598,N_3819,N_4455);
xor U4599 (N_4599,N_3412,N_4329);
and U4600 (N_4600,N_3028,N_3639);
or U4601 (N_4601,N_3874,N_3743);
or U4602 (N_4602,N_3437,N_3601);
xor U4603 (N_4603,N_3252,N_3230);
xnor U4604 (N_4604,N_4138,N_4308);
nand U4605 (N_4605,N_3320,N_4497);
and U4606 (N_4606,N_4145,N_3629);
and U4607 (N_4607,N_3810,N_4211);
nand U4608 (N_4608,N_4311,N_3987);
xor U4609 (N_4609,N_3722,N_3288);
xor U4610 (N_4610,N_4463,N_4139);
nand U4611 (N_4611,N_3756,N_3143);
xor U4612 (N_4612,N_3837,N_3281);
nand U4613 (N_4613,N_3672,N_3841);
xnor U4614 (N_4614,N_3044,N_3183);
xor U4615 (N_4615,N_3135,N_3370);
and U4616 (N_4616,N_4323,N_4316);
nor U4617 (N_4617,N_3585,N_4307);
nand U4618 (N_4618,N_3449,N_3858);
nand U4619 (N_4619,N_3442,N_3154);
nor U4620 (N_4620,N_3840,N_3235);
nand U4621 (N_4621,N_4336,N_3491);
or U4622 (N_4622,N_3261,N_3719);
nand U4623 (N_4623,N_3559,N_4478);
or U4624 (N_4624,N_3684,N_3942);
or U4625 (N_4625,N_3269,N_3345);
nor U4626 (N_4626,N_4391,N_3124);
or U4627 (N_4627,N_4255,N_4124);
and U4628 (N_4628,N_3401,N_3626);
nor U4629 (N_4629,N_4432,N_3764);
nor U4630 (N_4630,N_3781,N_4258);
and U4631 (N_4631,N_4374,N_3247);
or U4632 (N_4632,N_3204,N_4279);
xor U4633 (N_4633,N_4056,N_3661);
nand U4634 (N_4634,N_4392,N_3327);
xor U4635 (N_4635,N_3461,N_3851);
and U4636 (N_4636,N_4361,N_4452);
nor U4637 (N_4637,N_4094,N_4025);
nor U4638 (N_4638,N_3169,N_3470);
and U4639 (N_4639,N_3512,N_3354);
nand U4640 (N_4640,N_4039,N_4020);
nand U4641 (N_4641,N_3227,N_3333);
and U4642 (N_4642,N_3236,N_3710);
nand U4643 (N_4643,N_3633,N_4388);
xnor U4644 (N_4644,N_3416,N_3768);
or U4645 (N_4645,N_3807,N_3062);
xnor U4646 (N_4646,N_3507,N_4458);
or U4647 (N_4647,N_4352,N_3259);
and U4648 (N_4648,N_4416,N_4456);
nor U4649 (N_4649,N_3934,N_3834);
nor U4650 (N_4650,N_4333,N_3323);
xor U4651 (N_4651,N_3896,N_3617);
nand U4652 (N_4652,N_4221,N_3965);
and U4653 (N_4653,N_3482,N_3034);
xor U4654 (N_4654,N_4161,N_3572);
or U4655 (N_4655,N_4111,N_4435);
and U4656 (N_4656,N_4231,N_4453);
nor U4657 (N_4657,N_3194,N_3060);
xnor U4658 (N_4658,N_3243,N_4101);
xor U4659 (N_4659,N_3564,N_4437);
xor U4660 (N_4660,N_4367,N_3214);
nor U4661 (N_4661,N_4411,N_3215);
nor U4662 (N_4662,N_4436,N_3640);
and U4663 (N_4663,N_3166,N_4309);
nor U4664 (N_4664,N_4091,N_3220);
and U4665 (N_4665,N_3889,N_3102);
and U4666 (N_4666,N_3031,N_3552);
xnor U4667 (N_4667,N_4181,N_3048);
or U4668 (N_4668,N_3425,N_3517);
or U4669 (N_4669,N_4069,N_3935);
and U4670 (N_4670,N_3718,N_4083);
and U4671 (N_4671,N_3513,N_3636);
or U4672 (N_4672,N_3492,N_4287);
and U4673 (N_4673,N_3049,N_4234);
nor U4674 (N_4674,N_4220,N_3885);
nand U4675 (N_4675,N_3285,N_3150);
nand U4676 (N_4676,N_4470,N_3940);
xnor U4677 (N_4677,N_4189,N_4228);
nand U4678 (N_4678,N_3351,N_3078);
and U4679 (N_4679,N_4031,N_3076);
and U4680 (N_4680,N_4439,N_3613);
and U4681 (N_4681,N_3042,N_3010);
nand U4682 (N_4682,N_3747,N_3438);
xnor U4683 (N_4683,N_4270,N_4426);
nor U4684 (N_4684,N_4298,N_4113);
or U4685 (N_4685,N_4047,N_4070);
or U4686 (N_4686,N_3195,N_3244);
nor U4687 (N_4687,N_4427,N_3532);
xnor U4688 (N_4688,N_3975,N_3846);
xnor U4689 (N_4689,N_4163,N_4397);
and U4690 (N_4690,N_4053,N_3762);
and U4691 (N_4691,N_3598,N_4088);
nor U4692 (N_4692,N_3200,N_3299);
nand U4693 (N_4693,N_3117,N_3039);
nand U4694 (N_4694,N_3712,N_3095);
and U4695 (N_4695,N_3820,N_3436);
and U4696 (N_4696,N_4097,N_3346);
nand U4697 (N_4697,N_3758,N_3528);
nor U4698 (N_4698,N_3567,N_4003);
nand U4699 (N_4699,N_3337,N_3737);
xnor U4700 (N_4700,N_3925,N_3177);
or U4701 (N_4701,N_3123,N_3421);
and U4702 (N_4702,N_3892,N_3239);
xnor U4703 (N_4703,N_3145,N_3326);
nand U4704 (N_4704,N_3242,N_3847);
and U4705 (N_4705,N_3945,N_3356);
or U4706 (N_4706,N_4193,N_3251);
nand U4707 (N_4707,N_4477,N_4115);
xnor U4708 (N_4708,N_4265,N_3540);
nand U4709 (N_4709,N_3991,N_3179);
nor U4710 (N_4710,N_3094,N_4087);
and U4711 (N_4711,N_4132,N_3268);
nand U4712 (N_4712,N_3506,N_3895);
nor U4713 (N_4713,N_4045,N_3074);
xor U4714 (N_4714,N_3570,N_4283);
or U4715 (N_4715,N_3706,N_3724);
nor U4716 (N_4716,N_3817,N_4402);
nand U4717 (N_4717,N_4251,N_3799);
nand U4718 (N_4718,N_3486,N_3803);
nand U4719 (N_4719,N_3526,N_4268);
nor U4720 (N_4720,N_3995,N_3787);
nor U4721 (N_4721,N_3795,N_3900);
xor U4722 (N_4722,N_3589,N_4035);
xor U4723 (N_4723,N_3573,N_3035);
and U4724 (N_4724,N_3385,N_3361);
xnor U4725 (N_4725,N_3920,N_3304);
or U4726 (N_4726,N_3955,N_4379);
nor U4727 (N_4727,N_4269,N_3714);
or U4728 (N_4728,N_4103,N_3199);
xnor U4729 (N_4729,N_3216,N_4229);
or U4730 (N_4730,N_3016,N_3595);
nand U4731 (N_4731,N_3373,N_4202);
xnor U4732 (N_4732,N_4167,N_3692);
or U4733 (N_4733,N_4260,N_3348);
nand U4734 (N_4734,N_4222,N_3070);
xnor U4735 (N_4735,N_3015,N_3854);
nand U4736 (N_4736,N_3129,N_3402);
nor U4737 (N_4737,N_3377,N_4118);
and U4738 (N_4738,N_3201,N_3911);
xnor U4739 (N_4739,N_4233,N_4339);
or U4740 (N_4740,N_3422,N_3481);
xor U4741 (N_4741,N_3761,N_4475);
xnor U4742 (N_4742,N_3165,N_4005);
and U4743 (N_4743,N_3656,N_3434);
xor U4744 (N_4744,N_3157,N_4418);
or U4745 (N_4745,N_3100,N_4146);
nor U4746 (N_4746,N_3443,N_3563);
or U4747 (N_4747,N_3510,N_4030);
and U4748 (N_4748,N_3770,N_3833);
or U4749 (N_4749,N_3876,N_4294);
nand U4750 (N_4750,N_3398,N_3977);
and U4751 (N_4751,N_3957,N_3671);
nand U4752 (N_4752,N_3018,N_3265);
xnor U4753 (N_4753,N_3680,N_4357);
or U4754 (N_4754,N_3568,N_4178);
nor U4755 (N_4755,N_4280,N_3698);
nor U4756 (N_4756,N_3845,N_3852);
and U4757 (N_4757,N_4198,N_3005);
or U4758 (N_4758,N_3196,N_3116);
or U4759 (N_4759,N_3397,N_3565);
nor U4760 (N_4760,N_3677,N_3428);
and U4761 (N_4761,N_4071,N_3312);
or U4762 (N_4762,N_3602,N_4469);
nand U4763 (N_4763,N_4383,N_4358);
nor U4764 (N_4764,N_4344,N_3536);
or U4765 (N_4765,N_3417,N_4274);
nor U4766 (N_4766,N_4174,N_4396);
nand U4767 (N_4767,N_4444,N_3733);
or U4768 (N_4768,N_3555,N_4160);
xnor U4769 (N_4769,N_4290,N_4102);
nor U4770 (N_4770,N_3258,N_4114);
nand U4771 (N_4771,N_4313,N_4385);
and U4772 (N_4772,N_3745,N_3273);
nor U4773 (N_4773,N_3784,N_3184);
or U4774 (N_4774,N_4065,N_3149);
or U4775 (N_4775,N_4325,N_3349);
or U4776 (N_4776,N_4142,N_3147);
and U4777 (N_4777,N_3836,N_3212);
nand U4778 (N_4778,N_3144,N_4300);
or U4779 (N_4779,N_3537,N_3021);
xor U4780 (N_4780,N_3241,N_3113);
and U4781 (N_4781,N_4019,N_3072);
or U4782 (N_4782,N_4377,N_4017);
nand U4783 (N_4783,N_4442,N_4225);
nor U4784 (N_4784,N_3686,N_3751);
or U4785 (N_4785,N_4041,N_4008);
nor U4786 (N_4786,N_3396,N_4172);
and U4787 (N_4787,N_4408,N_3332);
and U4788 (N_4788,N_3918,N_4213);
or U4789 (N_4789,N_4354,N_3115);
or U4790 (N_4790,N_4147,N_3700);
nand U4791 (N_4791,N_3077,N_4295);
xnor U4792 (N_4792,N_3651,N_4401);
nor U4793 (N_4793,N_4485,N_3785);
nand U4794 (N_4794,N_4276,N_3109);
and U4795 (N_4795,N_3664,N_4150);
and U4796 (N_4796,N_3981,N_4495);
nand U4797 (N_4797,N_4296,N_4464);
or U4798 (N_4798,N_3295,N_4127);
or U4799 (N_4799,N_3358,N_3209);
or U4800 (N_4800,N_4390,N_3720);
nand U4801 (N_4801,N_3860,N_4043);
nand U4802 (N_4802,N_3400,N_3253);
and U4803 (N_4803,N_3831,N_3734);
xor U4804 (N_4804,N_3923,N_4382);
nor U4805 (N_4805,N_3052,N_3090);
xor U4806 (N_4806,N_3142,N_4483);
nand U4807 (N_4807,N_3271,N_3456);
and U4808 (N_4808,N_4471,N_3013);
xnor U4809 (N_4809,N_3689,N_3891);
or U4810 (N_4810,N_3612,N_3732);
xnor U4811 (N_4811,N_4214,N_3823);
and U4812 (N_4812,N_3494,N_3000);
xor U4813 (N_4813,N_3926,N_4200);
nand U4814 (N_4814,N_3739,N_3921);
xnor U4815 (N_4815,N_3992,N_4159);
or U4816 (N_4816,N_3435,N_3725);
nand U4817 (N_4817,N_3219,N_3472);
and U4818 (N_4818,N_3974,N_4184);
nand U4819 (N_4819,N_3596,N_4445);
nor U4820 (N_4820,N_3883,N_3959);
and U4821 (N_4821,N_3999,N_3814);
nor U4822 (N_4822,N_4499,N_3294);
and U4823 (N_4823,N_4218,N_3571);
xor U4824 (N_4824,N_3014,N_4494);
nand U4825 (N_4825,N_4170,N_3696);
and U4826 (N_4826,N_3757,N_4196);
xor U4827 (N_4827,N_4491,N_4496);
nand U4828 (N_4828,N_3856,N_3389);
or U4829 (N_4829,N_3575,N_3274);
xnor U4830 (N_4830,N_3222,N_4376);
and U4831 (N_4831,N_3500,N_3827);
xnor U4832 (N_4832,N_3364,N_3755);
nor U4833 (N_4833,N_3688,N_3105);
and U4834 (N_4834,N_3319,N_3064);
or U4835 (N_4835,N_3594,N_3255);
and U4836 (N_4836,N_4033,N_3736);
nor U4837 (N_4837,N_4125,N_3340);
xor U4838 (N_4838,N_3673,N_4051);
and U4839 (N_4839,N_3296,N_3058);
nor U4840 (N_4840,N_3270,N_4177);
xor U4841 (N_4841,N_4165,N_4350);
nand U4842 (N_4842,N_4073,N_4082);
xor U4843 (N_4843,N_4346,N_4375);
nor U4844 (N_4844,N_4117,N_3302);
xnor U4845 (N_4845,N_4281,N_3873);
and U4846 (N_4846,N_3705,N_4093);
xnor U4847 (N_4847,N_3384,N_3004);
nor U4848 (N_4848,N_4299,N_3284);
nor U4849 (N_4849,N_3985,N_3276);
nand U4850 (N_4850,N_3659,N_3468);
nand U4851 (N_4851,N_3409,N_3631);
nor U4852 (N_4852,N_4037,N_3210);
and U4853 (N_4853,N_4121,N_3742);
or U4854 (N_4854,N_3539,N_3190);
and U4855 (N_4855,N_3444,N_3628);
or U4856 (N_4856,N_3168,N_3167);
or U4857 (N_4857,N_4348,N_3560);
nand U4858 (N_4858,N_4048,N_3272);
xor U4859 (N_4859,N_3518,N_3307);
nor U4860 (N_4860,N_4106,N_4244);
nor U4861 (N_4861,N_4291,N_3393);
nand U4862 (N_4862,N_3250,N_4238);
and U4863 (N_4863,N_3454,N_3662);
xnor U4864 (N_4864,N_4286,N_3125);
nand U4865 (N_4865,N_3534,N_4252);
xnor U4866 (N_4866,N_4484,N_3012);
xnor U4867 (N_4867,N_4143,N_3410);
nand U4868 (N_4868,N_3081,N_3344);
nand U4869 (N_4869,N_4373,N_4448);
xnor U4870 (N_4870,N_3114,N_4058);
xnor U4871 (N_4871,N_3453,N_3600);
and U4872 (N_4872,N_3546,N_3708);
nor U4873 (N_4873,N_4314,N_3735);
nand U4874 (N_4874,N_3681,N_3246);
or U4875 (N_4875,N_3549,N_3792);
xnor U4876 (N_4876,N_4355,N_4064);
nor U4877 (N_4877,N_3801,N_4199);
xnor U4878 (N_4878,N_3023,N_4407);
or U4879 (N_4879,N_3146,N_3309);
or U4880 (N_4880,N_3488,N_3625);
nor U4881 (N_4881,N_3096,N_3156);
nand U4882 (N_4882,N_4078,N_3623);
or U4883 (N_4883,N_3324,N_4000);
nor U4884 (N_4884,N_4012,N_3809);
and U4885 (N_4885,N_3533,N_3137);
xor U4886 (N_4886,N_3707,N_3561);
nand U4887 (N_4887,N_3475,N_3979);
and U4888 (N_4888,N_3033,N_3535);
xnor U4889 (N_4889,N_3949,N_3003);
and U4890 (N_4890,N_4130,N_4187);
or U4891 (N_4891,N_3587,N_3178);
and U4892 (N_4892,N_3611,N_3830);
or U4893 (N_4893,N_3298,N_3511);
or U4894 (N_4894,N_3131,N_3174);
xor U4895 (N_4895,N_3961,N_3411);
nand U4896 (N_4896,N_3026,N_3228);
xor U4897 (N_4897,N_3110,N_4372);
nand U4898 (N_4898,N_4243,N_3483);
nand U4899 (N_4899,N_3007,N_3056);
xor U4900 (N_4900,N_3812,N_3842);
nor U4901 (N_4901,N_3347,N_3771);
nand U4902 (N_4902,N_3036,N_3937);
and U4903 (N_4903,N_3495,N_3863);
nor U4904 (N_4904,N_3399,N_3413);
nor U4905 (N_4905,N_3861,N_4107);
nand U4906 (N_4906,N_3694,N_3046);
nor U4907 (N_4907,N_3924,N_4072);
xnor U4908 (N_4908,N_4148,N_3588);
nor U4909 (N_4909,N_3352,N_3933);
or U4910 (N_4910,N_4266,N_4277);
nor U4911 (N_4911,N_3931,N_4320);
xnor U4912 (N_4912,N_3485,N_3884);
nand U4913 (N_4913,N_4176,N_4016);
nand U4914 (N_4914,N_3592,N_3780);
xor U4915 (N_4915,N_3515,N_3916);
or U4916 (N_4916,N_3279,N_3017);
xnor U4917 (N_4917,N_4074,N_4186);
nor U4918 (N_4918,N_3980,N_3501);
nand U4919 (N_4919,N_3654,N_4247);
nand U4920 (N_4920,N_4109,N_3765);
nand U4921 (N_4921,N_3429,N_4242);
xor U4922 (N_4922,N_4212,N_3525);
and U4923 (N_4923,N_3618,N_4013);
nand U4924 (N_4924,N_3815,N_3967);
xnor U4925 (N_4925,N_3291,N_3782);
xor U4926 (N_4926,N_3637,N_3120);
xnor U4927 (N_4927,N_4306,N_3375);
nor U4928 (N_4928,N_3257,N_4040);
nor U4929 (N_4929,N_4403,N_3093);
or U4930 (N_4930,N_4318,N_4371);
or U4931 (N_4931,N_4324,N_4034);
nor U4932 (N_4932,N_3141,N_3176);
nor U4933 (N_4933,N_3140,N_3727);
and U4934 (N_4934,N_4430,N_4479);
or U4935 (N_4935,N_3695,N_4340);
and U4936 (N_4936,N_3392,N_4068);
and U4937 (N_4937,N_3634,N_4112);
xor U4938 (N_4938,N_3188,N_4075);
xnor U4939 (N_4939,N_4149,N_4027);
nor U4940 (N_4940,N_4322,N_3158);
xor U4941 (N_4941,N_3630,N_3217);
or U4942 (N_4942,N_4438,N_3521);
or U4943 (N_4943,N_3293,N_4364);
and U4944 (N_4944,N_4466,N_3800);
and U4945 (N_4945,N_4141,N_4044);
or U4946 (N_4946,N_4046,N_3569);
nor U4947 (N_4947,N_3173,N_3202);
or U4948 (N_4948,N_3946,N_3604);
xnor U4949 (N_4949,N_3211,N_3063);
nor U4950 (N_4950,N_3480,N_3658);
nand U4951 (N_4951,N_3362,N_3994);
or U4952 (N_4952,N_4089,N_3055);
xor U4953 (N_4953,N_3426,N_4425);
or U4954 (N_4954,N_3287,N_3466);
and U4955 (N_4955,N_4334,N_3646);
nor U4956 (N_4956,N_4289,N_4486);
and U4957 (N_4957,N_3122,N_3906);
and U4958 (N_4958,N_3136,N_4345);
or U4959 (N_4959,N_3963,N_3740);
or U4960 (N_4960,N_4063,N_3766);
nor U4961 (N_4961,N_4096,N_4208);
and U4962 (N_4962,N_3621,N_4282);
nor U4963 (N_4963,N_3290,N_4011);
nand U4964 (N_4964,N_3690,N_4398);
and U4965 (N_4965,N_3419,N_3477);
nand U4966 (N_4966,N_3164,N_3774);
nor U4967 (N_4967,N_3447,N_3079);
and U4968 (N_4968,N_4195,N_3008);
xnor U4969 (N_4969,N_3059,N_4237);
and U4970 (N_4970,N_3053,N_3439);
or U4971 (N_4971,N_4328,N_4498);
xor U4972 (N_4972,N_3189,N_3952);
nor U4973 (N_4973,N_3024,N_3469);
nand U4974 (N_4974,N_3687,N_4024);
or U4975 (N_4975,N_3328,N_3881);
nor U4976 (N_4976,N_3138,N_4349);
nand U4977 (N_4977,N_3233,N_3867);
or U4978 (N_4978,N_3134,N_3489);
nor U4979 (N_4979,N_4055,N_4433);
or U4980 (N_4980,N_3607,N_3353);
or U4981 (N_4981,N_3245,N_4067);
nand U4982 (N_4982,N_4415,N_4338);
and U4983 (N_4983,N_3825,N_3574);
xor U4984 (N_4984,N_3289,N_3365);
xor U4985 (N_4985,N_3186,N_3582);
xnor U4986 (N_4986,N_3329,N_4171);
and U4987 (N_4987,N_4386,N_3193);
xnor U4988 (N_4988,N_4086,N_3121);
or U4989 (N_4989,N_4482,N_3905);
or U4990 (N_4990,N_3610,N_3380);
or U4991 (N_4991,N_3032,N_4363);
xor U4992 (N_4992,N_4014,N_3325);
or U4993 (N_4993,N_4273,N_4443);
and U4994 (N_4994,N_3054,N_3092);
or U4995 (N_4995,N_3386,N_4366);
xor U4996 (N_4996,N_3045,N_4370);
nand U4997 (N_4997,N_4059,N_3964);
or U4998 (N_4998,N_4081,N_4006);
nor U4999 (N_4999,N_3703,N_3663);
xnor U5000 (N_5000,N_4007,N_3300);
nand U5001 (N_5001,N_4085,N_4288);
or U5002 (N_5002,N_3566,N_3608);
and U5003 (N_5003,N_4330,N_3796);
nand U5004 (N_5004,N_3954,N_3606);
and U5005 (N_5005,N_3379,N_3783);
xor U5006 (N_5006,N_3414,N_3711);
nor U5007 (N_5007,N_3806,N_3670);
nand U5008 (N_5008,N_4028,N_3998);
nor U5009 (N_5009,N_3647,N_3019);
and U5010 (N_5010,N_4015,N_3226);
nand U5011 (N_5011,N_3128,N_4226);
and U5012 (N_5012,N_3557,N_4151);
xor U5013 (N_5013,N_3616,N_3773);
nor U5014 (N_5014,N_4465,N_3897);
xor U5015 (N_5015,N_3919,N_3730);
or U5016 (N_5016,N_3187,N_3904);
and U5017 (N_5017,N_3175,N_3382);
or U5018 (N_5018,N_4343,N_3778);
xnor U5019 (N_5019,N_3767,N_3106);
nand U5020 (N_5020,N_3972,N_3752);
or U5021 (N_5021,N_3948,N_4406);
or U5022 (N_5022,N_3148,N_3050);
or U5023 (N_5023,N_3009,N_4077);
nor U5024 (N_5024,N_3130,N_3180);
nand U5025 (N_5025,N_4488,N_3471);
or U5026 (N_5026,N_4095,N_3721);
nand U5027 (N_5027,N_3624,N_3888);
or U5028 (N_5028,N_4492,N_3151);
nand U5029 (N_5029,N_4278,N_3182);
xnor U5030 (N_5030,N_3619,N_4321);
nor U5031 (N_5031,N_4413,N_3359);
and U5032 (N_5032,N_3459,N_4032);
and U5033 (N_5033,N_3880,N_4054);
and U5034 (N_5034,N_4451,N_3950);
nor U5035 (N_5035,N_3723,N_4134);
or U5036 (N_5036,N_4429,N_3938);
and U5037 (N_5037,N_4454,N_3038);
nor U5038 (N_5038,N_3075,N_3682);
nor U5039 (N_5039,N_4175,N_4284);
xnor U5040 (N_5040,N_3263,N_3614);
nor U5041 (N_5041,N_4360,N_4140);
xor U5042 (N_5042,N_4428,N_4417);
and U5043 (N_5043,N_3225,N_3519);
and U5044 (N_5044,N_4062,N_4410);
or U5045 (N_5045,N_3336,N_4057);
nor U5046 (N_5046,N_3966,N_3467);
or U5047 (N_5047,N_4061,N_3152);
or U5048 (N_5048,N_3929,N_3638);
or U5049 (N_5049,N_3984,N_3657);
or U5050 (N_5050,N_4084,N_3828);
xnor U5051 (N_5051,N_4180,N_3645);
nor U5052 (N_5052,N_4144,N_3591);
nor U5053 (N_5053,N_4021,N_3207);
and U5054 (N_5054,N_4305,N_3181);
nor U5055 (N_5055,N_3597,N_3818);
or U5056 (N_5056,N_3527,N_3584);
nor U5057 (N_5057,N_3675,N_3249);
and U5058 (N_5058,N_3986,N_4099);
xor U5059 (N_5059,N_4337,N_3338);
xnor U5060 (N_5060,N_4481,N_4154);
or U5061 (N_5061,N_4365,N_3635);
nor U5062 (N_5062,N_3811,N_3609);
xor U5063 (N_5063,N_4245,N_4412);
nor U5064 (N_5064,N_3824,N_3254);
nand U5065 (N_5065,N_3073,N_3821);
or U5066 (N_5066,N_4210,N_3479);
or U5067 (N_5067,N_3543,N_3030);
nand U5068 (N_5068,N_3524,N_4302);
and U5069 (N_5069,N_4105,N_4248);
nor U5070 (N_5070,N_4310,N_3367);
and U5071 (N_5071,N_3544,N_3339);
xnor U5072 (N_5072,N_4440,N_3369);
nand U5073 (N_5073,N_3192,N_4166);
nand U5074 (N_5074,N_3522,N_3509);
xnor U5075 (N_5075,N_3523,N_3887);
nand U5076 (N_5076,N_3260,N_4191);
nand U5077 (N_5077,N_3292,N_3668);
and U5078 (N_5078,N_4472,N_3983);
nand U5079 (N_5079,N_4457,N_4190);
and U5080 (N_5080,N_3530,N_4450);
or U5081 (N_5081,N_4400,N_3996);
xnor U5082 (N_5082,N_3112,N_3407);
nor U5083 (N_5083,N_4327,N_4493);
and U5084 (N_5084,N_4253,N_3928);
and U5085 (N_5085,N_3932,N_3487);
nor U5086 (N_5086,N_4449,N_3041);
nand U5087 (N_5087,N_3699,N_3871);
or U5088 (N_5088,N_3088,N_3237);
and U5089 (N_5089,N_3171,N_3153);
or U5090 (N_5090,N_3576,N_4162);
xor U5091 (N_5091,N_3915,N_3898);
nor U5092 (N_5092,N_3693,N_3581);
nand U5093 (N_5093,N_3875,N_3368);
and U5094 (N_5094,N_3224,N_4459);
and U5095 (N_5095,N_3318,N_3098);
nor U5096 (N_5096,N_3069,N_3971);
and U5097 (N_5097,N_4080,N_4236);
xnor U5098 (N_5098,N_3378,N_3902);
nand U5099 (N_5099,N_4010,N_3430);
nor U5100 (N_5100,N_3798,N_3958);
nor U5101 (N_5101,N_3043,N_3843);
nand U5102 (N_5102,N_3020,N_3772);
xor U5103 (N_5103,N_3334,N_3490);
nor U5104 (N_5104,N_3748,N_3769);
and U5105 (N_5105,N_4271,N_3669);
xnor U5106 (N_5106,N_3813,N_3360);
nand U5107 (N_5107,N_3029,N_4192);
nand U5108 (N_5108,N_3797,N_3101);
nor U5109 (N_5109,N_4393,N_3071);
nand U5110 (N_5110,N_4395,N_4009);
xnor U5111 (N_5111,N_4404,N_3464);
and U5112 (N_5112,N_3248,N_4297);
and U5113 (N_5113,N_3432,N_3702);
nand U5114 (N_5114,N_3822,N_3930);
nor U5115 (N_5115,N_4131,N_3162);
xnor U5116 (N_5116,N_3869,N_3548);
and U5117 (N_5117,N_4050,N_3786);
nor U5118 (N_5118,N_3460,N_3057);
and U5119 (N_5119,N_4164,N_3498);
and U5120 (N_5120,N_4235,N_4224);
xor U5121 (N_5121,N_3068,N_3593);
and U5122 (N_5122,N_3508,N_4446);
nor U5123 (N_5123,N_4135,N_4381);
xor U5124 (N_5124,N_4173,N_3982);
nand U5125 (N_5125,N_3586,N_3912);
or U5126 (N_5126,N_4419,N_4489);
and U5127 (N_5127,N_3870,N_3366);
xor U5128 (N_5128,N_3701,N_3890);
or U5129 (N_5129,N_4384,N_4249);
or U5130 (N_5130,N_3650,N_4405);
xor U5131 (N_5131,N_3969,N_3943);
or U5132 (N_5132,N_3848,N_3750);
nor U5133 (N_5133,N_4319,N_4267);
and U5134 (N_5134,N_3580,N_3374);
or U5135 (N_5135,N_3163,N_3229);
nand U5136 (N_5136,N_4182,N_3643);
nand U5137 (N_5137,N_3099,N_3462);
nor U5138 (N_5138,N_3738,N_3423);
nand U5139 (N_5139,N_3886,N_3741);
xor U5140 (N_5140,N_3002,N_3864);
xnor U5141 (N_5141,N_3403,N_3642);
or U5142 (N_5142,N_3849,N_3632);
or U5143 (N_5143,N_3080,N_3893);
nand U5144 (N_5144,N_3715,N_3006);
nand U5145 (N_5145,N_3415,N_3853);
nor U5146 (N_5146,N_3901,N_3051);
and U5147 (N_5147,N_4156,N_4185);
nor U5148 (N_5148,N_3968,N_4023);
xnor U5149 (N_5149,N_3107,N_3838);
nand U5150 (N_5150,N_3406,N_3551);
xnor U5151 (N_5151,N_4215,N_3085);
nand U5152 (N_5152,N_3463,N_3908);
nor U5153 (N_5153,N_4206,N_4157);
nor U5154 (N_5154,N_3944,N_4490);
nand U5155 (N_5155,N_3067,N_3622);
or U5156 (N_5156,N_4326,N_3476);
nor U5157 (N_5157,N_3816,N_4254);
xor U5158 (N_5158,N_4120,N_3022);
nor U5159 (N_5159,N_3388,N_3914);
xor U5160 (N_5160,N_3306,N_3514);
nor U5161 (N_5161,N_3865,N_3839);
xnor U5162 (N_5162,N_3717,N_4002);
xor U5163 (N_5163,N_3788,N_3280);
nor U5164 (N_5164,N_3286,N_3278);
and U5165 (N_5165,N_4036,N_3037);
or U5166 (N_5166,N_3804,N_3108);
and U5167 (N_5167,N_3315,N_4209);
nand U5168 (N_5168,N_3197,N_3894);
xnor U5169 (N_5169,N_3529,N_3065);
or U5170 (N_5170,N_4304,N_4026);
and U5171 (N_5171,N_3383,N_4312);
and U5172 (N_5172,N_3844,N_3605);
nand U5173 (N_5173,N_3922,N_3583);
and U5174 (N_5174,N_4066,N_3746);
and U5175 (N_5175,N_4476,N_3866);
or U5176 (N_5176,N_3556,N_4261);
and U5177 (N_5177,N_3111,N_4223);
nand U5178 (N_5178,N_3939,N_3503);
nor U5179 (N_5179,N_3139,N_4301);
nand U5180 (N_5180,N_3440,N_4090);
xnor U5181 (N_5181,N_4133,N_3198);
and U5182 (N_5182,N_4227,N_3446);
or U5183 (N_5183,N_4467,N_3086);
or U5184 (N_5184,N_4351,N_4022);
nand U5185 (N_5185,N_3653,N_4205);
nand U5186 (N_5186,N_3185,N_3473);
or U5187 (N_5187,N_4079,N_3342);
and U5188 (N_5188,N_3205,N_4441);
nand U5189 (N_5189,N_3240,N_3603);
and U5190 (N_5190,N_4076,N_3277);
xor U5191 (N_5191,N_4108,N_3231);
and U5192 (N_5192,N_3910,N_3343);
or U5193 (N_5193,N_3376,N_4049);
and U5194 (N_5194,N_4201,N_4259);
and U5195 (N_5195,N_3674,N_3047);
nor U5196 (N_5196,N_3091,N_3394);
and U5197 (N_5197,N_4001,N_3208);
and U5198 (N_5198,N_3317,N_3027);
xnor U5199 (N_5199,N_3322,N_4335);
and U5200 (N_5200,N_3691,N_3790);
nor U5201 (N_5201,N_3505,N_4285);
nand U5202 (N_5202,N_3218,N_3562);
nand U5203 (N_5203,N_3749,N_3420);
and U5204 (N_5204,N_3808,N_4399);
nor U5205 (N_5205,N_4042,N_3713);
and U5206 (N_5206,N_3084,N_4424);
and U5207 (N_5207,N_4431,N_3802);
and U5208 (N_5208,N_4414,N_4230);
nand U5209 (N_5209,N_3357,N_3206);
and U5210 (N_5210,N_4116,N_3496);
and U5211 (N_5211,N_3978,N_3666);
or U5212 (N_5212,N_3455,N_4246);
xor U5213 (N_5213,N_3960,N_3297);
and U5214 (N_5214,N_3066,N_3956);
nand U5215 (N_5215,N_3541,N_3962);
xnor U5216 (N_5216,N_4098,N_3451);
and U5217 (N_5217,N_3754,N_3547);
nor U5218 (N_5218,N_3878,N_3448);
nand U5219 (N_5219,N_3953,N_4422);
or U5220 (N_5220,N_3993,N_3578);
xor U5221 (N_5221,N_4110,N_3433);
nand U5222 (N_5222,N_3314,N_4104);
nand U5223 (N_5223,N_3089,N_3649);
xnor U5224 (N_5224,N_4264,N_3262);
and U5225 (N_5225,N_3829,N_3520);
nand U5226 (N_5226,N_3709,N_3554);
nand U5227 (N_5227,N_4315,N_4263);
nor U5228 (N_5228,N_3310,N_3363);
nor U5229 (N_5229,N_3899,N_3424);
xor U5230 (N_5230,N_4362,N_4197);
and U5231 (N_5231,N_3879,N_4461);
or U5232 (N_5232,N_3493,N_4188);
or U5233 (N_5233,N_3667,N_4421);
nor U5234 (N_5234,N_4169,N_4394);
and U5235 (N_5235,N_4119,N_3997);
xor U5236 (N_5236,N_4447,N_3213);
xor U5237 (N_5237,N_3553,N_3395);
and U5238 (N_5238,N_3457,N_4052);
nand U5239 (N_5239,N_3321,N_4293);
xor U5240 (N_5240,N_4275,N_4207);
nor U5241 (N_5241,N_3025,N_4369);
nand U5242 (N_5242,N_3590,N_4219);
and U5243 (N_5243,N_3615,N_3791);
and U5244 (N_5244,N_4257,N_3282);
nor U5245 (N_5245,N_3728,N_3283);
or U5246 (N_5246,N_3223,N_4474);
or U5247 (N_5247,N_3504,N_3478);
xor U5248 (N_5248,N_3744,N_3665);
nor U5249 (N_5249,N_4203,N_4239);
or U5250 (N_5250,N_3580,N_3417);
xnor U5251 (N_5251,N_4361,N_4078);
nand U5252 (N_5252,N_4133,N_3780);
or U5253 (N_5253,N_3377,N_4055);
nor U5254 (N_5254,N_4451,N_3944);
and U5255 (N_5255,N_3119,N_3451);
nor U5256 (N_5256,N_4029,N_3785);
xnor U5257 (N_5257,N_4377,N_3367);
nor U5258 (N_5258,N_4107,N_3150);
nand U5259 (N_5259,N_3361,N_3608);
or U5260 (N_5260,N_3962,N_3425);
and U5261 (N_5261,N_3975,N_3099);
or U5262 (N_5262,N_4054,N_3810);
and U5263 (N_5263,N_4172,N_3739);
xor U5264 (N_5264,N_3977,N_3229);
nor U5265 (N_5265,N_4060,N_4056);
or U5266 (N_5266,N_3692,N_4144);
nand U5267 (N_5267,N_3289,N_4394);
nor U5268 (N_5268,N_3744,N_4001);
nand U5269 (N_5269,N_4443,N_3636);
xnor U5270 (N_5270,N_3579,N_4384);
and U5271 (N_5271,N_3381,N_3230);
and U5272 (N_5272,N_4390,N_4418);
nor U5273 (N_5273,N_3290,N_3099);
xor U5274 (N_5274,N_3317,N_3849);
nand U5275 (N_5275,N_3678,N_3884);
xnor U5276 (N_5276,N_4116,N_3704);
xnor U5277 (N_5277,N_3840,N_3487);
nor U5278 (N_5278,N_3101,N_4248);
nand U5279 (N_5279,N_4440,N_3808);
or U5280 (N_5280,N_3527,N_3161);
nand U5281 (N_5281,N_4319,N_3843);
or U5282 (N_5282,N_3511,N_3726);
xnor U5283 (N_5283,N_3150,N_3988);
xnor U5284 (N_5284,N_3786,N_4494);
xor U5285 (N_5285,N_3358,N_3469);
nand U5286 (N_5286,N_4353,N_3622);
xnor U5287 (N_5287,N_3723,N_3146);
xnor U5288 (N_5288,N_3383,N_4214);
xor U5289 (N_5289,N_3216,N_4396);
xnor U5290 (N_5290,N_4227,N_3012);
xnor U5291 (N_5291,N_4293,N_3042);
and U5292 (N_5292,N_3984,N_3404);
xor U5293 (N_5293,N_3188,N_3322);
nand U5294 (N_5294,N_3287,N_4104);
or U5295 (N_5295,N_3313,N_3052);
xnor U5296 (N_5296,N_3734,N_3263);
or U5297 (N_5297,N_3112,N_3713);
nor U5298 (N_5298,N_3193,N_3705);
nand U5299 (N_5299,N_4053,N_4062);
nor U5300 (N_5300,N_4299,N_3782);
xor U5301 (N_5301,N_4339,N_3545);
nor U5302 (N_5302,N_4283,N_4180);
xor U5303 (N_5303,N_4429,N_3546);
xnor U5304 (N_5304,N_3099,N_3988);
and U5305 (N_5305,N_3213,N_3040);
nand U5306 (N_5306,N_3423,N_4181);
xor U5307 (N_5307,N_3518,N_4205);
xor U5308 (N_5308,N_3256,N_3840);
or U5309 (N_5309,N_3566,N_3994);
nand U5310 (N_5310,N_4345,N_4452);
nor U5311 (N_5311,N_4160,N_3646);
nor U5312 (N_5312,N_4455,N_3786);
and U5313 (N_5313,N_4052,N_4072);
and U5314 (N_5314,N_4220,N_3553);
or U5315 (N_5315,N_4307,N_3050);
or U5316 (N_5316,N_3784,N_3452);
and U5317 (N_5317,N_3074,N_4357);
and U5318 (N_5318,N_4487,N_3925);
xnor U5319 (N_5319,N_3496,N_4119);
and U5320 (N_5320,N_3334,N_3002);
nand U5321 (N_5321,N_4495,N_3559);
or U5322 (N_5322,N_3711,N_3780);
xor U5323 (N_5323,N_4003,N_4000);
nor U5324 (N_5324,N_3734,N_4137);
nand U5325 (N_5325,N_3720,N_3914);
xnor U5326 (N_5326,N_4401,N_3409);
xnor U5327 (N_5327,N_4349,N_4058);
xnor U5328 (N_5328,N_3938,N_3193);
xor U5329 (N_5329,N_4465,N_3360);
nor U5330 (N_5330,N_4231,N_3803);
or U5331 (N_5331,N_4014,N_4032);
nand U5332 (N_5332,N_3879,N_4361);
or U5333 (N_5333,N_3232,N_3557);
nor U5334 (N_5334,N_3147,N_4104);
nor U5335 (N_5335,N_4282,N_3725);
or U5336 (N_5336,N_3013,N_4328);
and U5337 (N_5337,N_4469,N_3746);
or U5338 (N_5338,N_4066,N_3913);
nor U5339 (N_5339,N_3863,N_4429);
or U5340 (N_5340,N_3381,N_3261);
nor U5341 (N_5341,N_4208,N_3538);
xnor U5342 (N_5342,N_3445,N_3897);
nand U5343 (N_5343,N_3816,N_4087);
xor U5344 (N_5344,N_4329,N_4207);
and U5345 (N_5345,N_3881,N_3209);
or U5346 (N_5346,N_3753,N_4355);
or U5347 (N_5347,N_3011,N_3093);
and U5348 (N_5348,N_3664,N_3208);
xor U5349 (N_5349,N_3048,N_4461);
nor U5350 (N_5350,N_3808,N_4087);
nor U5351 (N_5351,N_3898,N_3971);
and U5352 (N_5352,N_3109,N_3073);
nand U5353 (N_5353,N_3539,N_3505);
and U5354 (N_5354,N_4428,N_4379);
xor U5355 (N_5355,N_3495,N_3315);
nand U5356 (N_5356,N_3006,N_4328);
nor U5357 (N_5357,N_3221,N_3310);
nor U5358 (N_5358,N_3953,N_4287);
nor U5359 (N_5359,N_3160,N_3355);
and U5360 (N_5360,N_3754,N_3193);
nor U5361 (N_5361,N_3577,N_3974);
and U5362 (N_5362,N_3727,N_3855);
or U5363 (N_5363,N_3521,N_3211);
or U5364 (N_5364,N_3268,N_3126);
xnor U5365 (N_5365,N_3619,N_3373);
or U5366 (N_5366,N_3179,N_3542);
xnor U5367 (N_5367,N_3092,N_3029);
xor U5368 (N_5368,N_3464,N_4430);
and U5369 (N_5369,N_4489,N_3561);
nand U5370 (N_5370,N_3597,N_3392);
xnor U5371 (N_5371,N_3236,N_3952);
and U5372 (N_5372,N_3220,N_3947);
nand U5373 (N_5373,N_4473,N_3694);
or U5374 (N_5374,N_3927,N_3035);
xnor U5375 (N_5375,N_3992,N_3837);
or U5376 (N_5376,N_3041,N_4281);
or U5377 (N_5377,N_3394,N_4185);
and U5378 (N_5378,N_4113,N_4399);
and U5379 (N_5379,N_3552,N_4429);
or U5380 (N_5380,N_3334,N_3783);
xnor U5381 (N_5381,N_3723,N_4055);
and U5382 (N_5382,N_3098,N_4194);
xor U5383 (N_5383,N_3066,N_3127);
and U5384 (N_5384,N_3800,N_3725);
nor U5385 (N_5385,N_3226,N_4113);
nand U5386 (N_5386,N_3266,N_3121);
nor U5387 (N_5387,N_3198,N_3493);
nand U5388 (N_5388,N_3537,N_3012);
nand U5389 (N_5389,N_4341,N_3237);
nor U5390 (N_5390,N_4208,N_4413);
and U5391 (N_5391,N_4425,N_3295);
nor U5392 (N_5392,N_4285,N_4428);
nand U5393 (N_5393,N_3852,N_3258);
or U5394 (N_5394,N_3139,N_3376);
xor U5395 (N_5395,N_4316,N_4060);
or U5396 (N_5396,N_4426,N_4238);
and U5397 (N_5397,N_3157,N_3491);
nor U5398 (N_5398,N_3950,N_3005);
xnor U5399 (N_5399,N_3393,N_3944);
nand U5400 (N_5400,N_3563,N_3914);
or U5401 (N_5401,N_4072,N_3916);
nand U5402 (N_5402,N_4248,N_3695);
xnor U5403 (N_5403,N_3995,N_3434);
nand U5404 (N_5404,N_3377,N_3552);
xnor U5405 (N_5405,N_3612,N_3703);
xor U5406 (N_5406,N_3515,N_3410);
xnor U5407 (N_5407,N_3276,N_4173);
and U5408 (N_5408,N_3045,N_3198);
nor U5409 (N_5409,N_3056,N_3136);
and U5410 (N_5410,N_4109,N_3102);
nand U5411 (N_5411,N_4213,N_3036);
xnor U5412 (N_5412,N_3173,N_4284);
xor U5413 (N_5413,N_3216,N_3640);
nor U5414 (N_5414,N_3564,N_3311);
nand U5415 (N_5415,N_3365,N_3740);
nor U5416 (N_5416,N_3292,N_3303);
nor U5417 (N_5417,N_3025,N_3027);
nand U5418 (N_5418,N_4404,N_4321);
xnor U5419 (N_5419,N_3700,N_4468);
nor U5420 (N_5420,N_4030,N_3272);
and U5421 (N_5421,N_3646,N_3217);
nor U5422 (N_5422,N_3914,N_4344);
nand U5423 (N_5423,N_3823,N_3668);
nor U5424 (N_5424,N_3196,N_3658);
nor U5425 (N_5425,N_4070,N_4028);
nand U5426 (N_5426,N_3467,N_3164);
nor U5427 (N_5427,N_4015,N_3460);
or U5428 (N_5428,N_3399,N_3472);
nand U5429 (N_5429,N_4405,N_3603);
and U5430 (N_5430,N_3548,N_3822);
nand U5431 (N_5431,N_4383,N_3985);
xnor U5432 (N_5432,N_3790,N_4228);
or U5433 (N_5433,N_4345,N_4041);
nand U5434 (N_5434,N_3666,N_3571);
or U5435 (N_5435,N_3648,N_3732);
nor U5436 (N_5436,N_3714,N_3945);
or U5437 (N_5437,N_4053,N_3152);
and U5438 (N_5438,N_3552,N_4263);
nor U5439 (N_5439,N_3643,N_3493);
or U5440 (N_5440,N_3075,N_4378);
nor U5441 (N_5441,N_3006,N_3682);
nand U5442 (N_5442,N_3168,N_3703);
nand U5443 (N_5443,N_3861,N_3530);
nor U5444 (N_5444,N_3892,N_3163);
nand U5445 (N_5445,N_3323,N_3942);
xnor U5446 (N_5446,N_4249,N_3180);
xor U5447 (N_5447,N_4338,N_3404);
or U5448 (N_5448,N_4278,N_4099);
nand U5449 (N_5449,N_3250,N_3353);
nor U5450 (N_5450,N_4384,N_4380);
nor U5451 (N_5451,N_3357,N_3954);
nand U5452 (N_5452,N_4458,N_3186);
nand U5453 (N_5453,N_3443,N_3352);
nand U5454 (N_5454,N_4449,N_3133);
nand U5455 (N_5455,N_3228,N_4136);
and U5456 (N_5456,N_3698,N_3470);
nor U5457 (N_5457,N_3479,N_3338);
xnor U5458 (N_5458,N_3896,N_3812);
nor U5459 (N_5459,N_3861,N_3133);
nor U5460 (N_5460,N_3255,N_4037);
and U5461 (N_5461,N_4002,N_4202);
and U5462 (N_5462,N_3811,N_3403);
and U5463 (N_5463,N_4375,N_3261);
nand U5464 (N_5464,N_3757,N_4371);
and U5465 (N_5465,N_3966,N_3301);
xor U5466 (N_5466,N_3908,N_4214);
xor U5467 (N_5467,N_3915,N_4337);
nor U5468 (N_5468,N_4189,N_3552);
xor U5469 (N_5469,N_4248,N_3969);
xnor U5470 (N_5470,N_3767,N_3437);
or U5471 (N_5471,N_4495,N_3216);
nor U5472 (N_5472,N_4168,N_3190);
or U5473 (N_5473,N_3330,N_3323);
nor U5474 (N_5474,N_3015,N_4373);
nor U5475 (N_5475,N_3930,N_4460);
and U5476 (N_5476,N_3510,N_3555);
or U5477 (N_5477,N_3416,N_3563);
xnor U5478 (N_5478,N_3803,N_4398);
and U5479 (N_5479,N_3087,N_3625);
and U5480 (N_5480,N_3247,N_3767);
xor U5481 (N_5481,N_4168,N_3867);
nor U5482 (N_5482,N_3285,N_3588);
nor U5483 (N_5483,N_3014,N_3013);
xnor U5484 (N_5484,N_3778,N_4486);
or U5485 (N_5485,N_3693,N_3457);
and U5486 (N_5486,N_3820,N_3837);
xnor U5487 (N_5487,N_3678,N_3894);
nand U5488 (N_5488,N_3895,N_3081);
nand U5489 (N_5489,N_3046,N_3055);
xor U5490 (N_5490,N_3695,N_4245);
nand U5491 (N_5491,N_4327,N_3909);
nor U5492 (N_5492,N_4316,N_3193);
and U5493 (N_5493,N_3804,N_3597);
nor U5494 (N_5494,N_4027,N_4470);
or U5495 (N_5495,N_4477,N_3004);
or U5496 (N_5496,N_3532,N_3425);
or U5497 (N_5497,N_3408,N_3407);
and U5498 (N_5498,N_3383,N_3050);
xnor U5499 (N_5499,N_3484,N_3382);
nand U5500 (N_5500,N_4290,N_4093);
nor U5501 (N_5501,N_3848,N_3064);
and U5502 (N_5502,N_3063,N_3339);
xnor U5503 (N_5503,N_3108,N_3514);
nor U5504 (N_5504,N_3614,N_3212);
or U5505 (N_5505,N_4063,N_3387);
and U5506 (N_5506,N_4440,N_4361);
nor U5507 (N_5507,N_3505,N_3326);
and U5508 (N_5508,N_4130,N_4398);
and U5509 (N_5509,N_3818,N_4422);
and U5510 (N_5510,N_4009,N_4371);
nand U5511 (N_5511,N_3859,N_3149);
nand U5512 (N_5512,N_3820,N_3475);
and U5513 (N_5513,N_3978,N_3690);
or U5514 (N_5514,N_3015,N_3367);
xnor U5515 (N_5515,N_3378,N_4377);
nor U5516 (N_5516,N_4155,N_3771);
and U5517 (N_5517,N_4109,N_3480);
and U5518 (N_5518,N_3674,N_4470);
or U5519 (N_5519,N_4110,N_3799);
nor U5520 (N_5520,N_3193,N_4311);
nor U5521 (N_5521,N_4234,N_4274);
or U5522 (N_5522,N_3734,N_3781);
xnor U5523 (N_5523,N_3462,N_4276);
and U5524 (N_5524,N_3783,N_4241);
or U5525 (N_5525,N_3474,N_4314);
nor U5526 (N_5526,N_3548,N_4085);
xor U5527 (N_5527,N_3345,N_3334);
nand U5528 (N_5528,N_3498,N_4091);
nand U5529 (N_5529,N_3994,N_3286);
nand U5530 (N_5530,N_4073,N_3075);
or U5531 (N_5531,N_3661,N_4020);
xnor U5532 (N_5532,N_3383,N_4487);
nor U5533 (N_5533,N_4117,N_3330);
nand U5534 (N_5534,N_4288,N_3181);
or U5535 (N_5535,N_3122,N_3833);
and U5536 (N_5536,N_3628,N_3215);
nor U5537 (N_5537,N_3233,N_4121);
xor U5538 (N_5538,N_3821,N_3722);
nand U5539 (N_5539,N_4445,N_3753);
or U5540 (N_5540,N_3226,N_3865);
xnor U5541 (N_5541,N_3667,N_3069);
xor U5542 (N_5542,N_4389,N_3591);
nor U5543 (N_5543,N_4122,N_3423);
xnor U5544 (N_5544,N_4135,N_3643);
xor U5545 (N_5545,N_3386,N_3465);
or U5546 (N_5546,N_3630,N_4051);
nor U5547 (N_5547,N_3944,N_4099);
nand U5548 (N_5548,N_3972,N_3146);
and U5549 (N_5549,N_4430,N_3179);
and U5550 (N_5550,N_3880,N_3478);
nor U5551 (N_5551,N_3844,N_4001);
and U5552 (N_5552,N_3796,N_3742);
and U5553 (N_5553,N_3734,N_3183);
nand U5554 (N_5554,N_3081,N_4261);
or U5555 (N_5555,N_3886,N_4065);
and U5556 (N_5556,N_3296,N_3388);
or U5557 (N_5557,N_3898,N_3885);
xor U5558 (N_5558,N_3586,N_3407);
or U5559 (N_5559,N_3133,N_4353);
nand U5560 (N_5560,N_3104,N_3080);
or U5561 (N_5561,N_4083,N_3856);
or U5562 (N_5562,N_3499,N_3311);
nor U5563 (N_5563,N_3468,N_4078);
and U5564 (N_5564,N_4489,N_3165);
xor U5565 (N_5565,N_3742,N_4300);
or U5566 (N_5566,N_4331,N_4025);
nor U5567 (N_5567,N_4057,N_3988);
nand U5568 (N_5568,N_3359,N_3530);
and U5569 (N_5569,N_4240,N_3049);
or U5570 (N_5570,N_3299,N_3003);
xnor U5571 (N_5571,N_3781,N_3823);
xnor U5572 (N_5572,N_3495,N_4284);
or U5573 (N_5573,N_4452,N_3092);
nor U5574 (N_5574,N_4046,N_4357);
nand U5575 (N_5575,N_3209,N_3180);
or U5576 (N_5576,N_3972,N_4220);
xnor U5577 (N_5577,N_3370,N_3825);
nor U5578 (N_5578,N_4282,N_3849);
nand U5579 (N_5579,N_4369,N_3705);
or U5580 (N_5580,N_4468,N_3688);
nor U5581 (N_5581,N_3602,N_4353);
nor U5582 (N_5582,N_3439,N_3760);
or U5583 (N_5583,N_3946,N_3592);
and U5584 (N_5584,N_4021,N_4209);
or U5585 (N_5585,N_4178,N_4066);
xnor U5586 (N_5586,N_3446,N_3643);
nor U5587 (N_5587,N_3864,N_3741);
or U5588 (N_5588,N_3379,N_3993);
and U5589 (N_5589,N_3604,N_3074);
and U5590 (N_5590,N_3182,N_3274);
nor U5591 (N_5591,N_3004,N_4224);
or U5592 (N_5592,N_3690,N_3913);
nand U5593 (N_5593,N_4053,N_4350);
xnor U5594 (N_5594,N_3131,N_3041);
nand U5595 (N_5595,N_3920,N_4378);
nand U5596 (N_5596,N_3073,N_3689);
nor U5597 (N_5597,N_3173,N_4017);
or U5598 (N_5598,N_3303,N_3731);
xor U5599 (N_5599,N_4194,N_4214);
or U5600 (N_5600,N_3870,N_3672);
xnor U5601 (N_5601,N_3350,N_3048);
nor U5602 (N_5602,N_4440,N_3525);
nand U5603 (N_5603,N_3101,N_4192);
nor U5604 (N_5604,N_3257,N_3373);
xor U5605 (N_5605,N_3598,N_3332);
and U5606 (N_5606,N_3621,N_4178);
and U5607 (N_5607,N_4101,N_3882);
xor U5608 (N_5608,N_3812,N_3860);
and U5609 (N_5609,N_3659,N_3792);
nand U5610 (N_5610,N_4309,N_4430);
nand U5611 (N_5611,N_4389,N_4210);
xnor U5612 (N_5612,N_3937,N_4152);
or U5613 (N_5613,N_3783,N_3552);
xnor U5614 (N_5614,N_4460,N_3661);
or U5615 (N_5615,N_3300,N_3392);
or U5616 (N_5616,N_3995,N_4229);
nor U5617 (N_5617,N_3547,N_4407);
xnor U5618 (N_5618,N_4444,N_3434);
nor U5619 (N_5619,N_4466,N_3873);
xnor U5620 (N_5620,N_4381,N_3098);
nand U5621 (N_5621,N_3227,N_3058);
nand U5622 (N_5622,N_3413,N_4430);
and U5623 (N_5623,N_4414,N_3966);
or U5624 (N_5624,N_4006,N_3876);
and U5625 (N_5625,N_3579,N_3865);
or U5626 (N_5626,N_3356,N_3193);
or U5627 (N_5627,N_4439,N_4361);
nor U5628 (N_5628,N_3221,N_3261);
or U5629 (N_5629,N_4062,N_3759);
or U5630 (N_5630,N_4334,N_4063);
and U5631 (N_5631,N_3493,N_4099);
xnor U5632 (N_5632,N_3293,N_4405);
or U5633 (N_5633,N_3260,N_3262);
or U5634 (N_5634,N_4285,N_4188);
and U5635 (N_5635,N_3151,N_4012);
xor U5636 (N_5636,N_3531,N_3695);
xnor U5637 (N_5637,N_3705,N_3218);
xnor U5638 (N_5638,N_3867,N_3673);
nor U5639 (N_5639,N_3216,N_3877);
nor U5640 (N_5640,N_4326,N_4205);
xor U5641 (N_5641,N_3922,N_4209);
nor U5642 (N_5642,N_3544,N_3465);
and U5643 (N_5643,N_4080,N_3043);
nand U5644 (N_5644,N_3912,N_3250);
nand U5645 (N_5645,N_3701,N_3147);
nand U5646 (N_5646,N_4022,N_3330);
and U5647 (N_5647,N_4430,N_3896);
and U5648 (N_5648,N_4377,N_3761);
nor U5649 (N_5649,N_3509,N_3315);
or U5650 (N_5650,N_4411,N_4258);
nand U5651 (N_5651,N_3125,N_4004);
and U5652 (N_5652,N_3327,N_3678);
nor U5653 (N_5653,N_4166,N_3962);
or U5654 (N_5654,N_3004,N_4074);
and U5655 (N_5655,N_4180,N_3034);
and U5656 (N_5656,N_4434,N_3571);
nand U5657 (N_5657,N_3472,N_3031);
nor U5658 (N_5658,N_3121,N_4342);
and U5659 (N_5659,N_3537,N_3682);
xnor U5660 (N_5660,N_3559,N_3541);
nor U5661 (N_5661,N_3673,N_3742);
nand U5662 (N_5662,N_3925,N_3551);
xor U5663 (N_5663,N_3611,N_3878);
and U5664 (N_5664,N_3470,N_3887);
nor U5665 (N_5665,N_3519,N_3467);
xor U5666 (N_5666,N_3052,N_3274);
and U5667 (N_5667,N_4243,N_4277);
nand U5668 (N_5668,N_4265,N_3937);
xnor U5669 (N_5669,N_3764,N_4261);
and U5670 (N_5670,N_4098,N_3959);
xnor U5671 (N_5671,N_4005,N_3435);
nor U5672 (N_5672,N_3702,N_4140);
and U5673 (N_5673,N_3063,N_3361);
or U5674 (N_5674,N_4172,N_4070);
and U5675 (N_5675,N_4314,N_3595);
and U5676 (N_5676,N_3954,N_3360);
and U5677 (N_5677,N_3692,N_3933);
and U5678 (N_5678,N_3521,N_3871);
and U5679 (N_5679,N_3986,N_4236);
and U5680 (N_5680,N_3230,N_3372);
and U5681 (N_5681,N_3029,N_4476);
nand U5682 (N_5682,N_4004,N_4374);
and U5683 (N_5683,N_4409,N_4270);
and U5684 (N_5684,N_4283,N_4297);
and U5685 (N_5685,N_3364,N_4224);
nor U5686 (N_5686,N_3341,N_3662);
nand U5687 (N_5687,N_3395,N_3501);
xnor U5688 (N_5688,N_4166,N_3441);
or U5689 (N_5689,N_4274,N_3775);
or U5690 (N_5690,N_3732,N_3746);
or U5691 (N_5691,N_3281,N_3879);
nand U5692 (N_5692,N_4356,N_3517);
nor U5693 (N_5693,N_3915,N_4141);
xnor U5694 (N_5694,N_4339,N_4069);
and U5695 (N_5695,N_3131,N_3909);
nand U5696 (N_5696,N_3100,N_3186);
xnor U5697 (N_5697,N_3475,N_3121);
or U5698 (N_5698,N_3016,N_3581);
and U5699 (N_5699,N_3853,N_3862);
nor U5700 (N_5700,N_3488,N_4053);
and U5701 (N_5701,N_3813,N_3117);
or U5702 (N_5702,N_3341,N_3419);
xor U5703 (N_5703,N_3536,N_4130);
and U5704 (N_5704,N_3431,N_3669);
and U5705 (N_5705,N_3851,N_4080);
and U5706 (N_5706,N_3017,N_3392);
and U5707 (N_5707,N_3855,N_3664);
xnor U5708 (N_5708,N_4044,N_3744);
xnor U5709 (N_5709,N_4237,N_3604);
or U5710 (N_5710,N_3866,N_3742);
nor U5711 (N_5711,N_3103,N_3777);
nor U5712 (N_5712,N_4245,N_4082);
or U5713 (N_5713,N_3867,N_3993);
xor U5714 (N_5714,N_4186,N_3194);
and U5715 (N_5715,N_3443,N_4275);
xnor U5716 (N_5716,N_3207,N_3843);
or U5717 (N_5717,N_3139,N_4066);
nand U5718 (N_5718,N_3160,N_3555);
and U5719 (N_5719,N_4221,N_3809);
and U5720 (N_5720,N_3932,N_3467);
nand U5721 (N_5721,N_4395,N_3613);
nor U5722 (N_5722,N_3487,N_3709);
or U5723 (N_5723,N_3455,N_3807);
and U5724 (N_5724,N_3491,N_4229);
xnor U5725 (N_5725,N_3993,N_3954);
and U5726 (N_5726,N_3085,N_4111);
or U5727 (N_5727,N_4030,N_3516);
and U5728 (N_5728,N_4332,N_3194);
xnor U5729 (N_5729,N_3906,N_3367);
xnor U5730 (N_5730,N_4114,N_4257);
nand U5731 (N_5731,N_3069,N_4019);
or U5732 (N_5732,N_3414,N_4342);
nor U5733 (N_5733,N_3404,N_4425);
xor U5734 (N_5734,N_3043,N_4485);
and U5735 (N_5735,N_3807,N_3572);
nor U5736 (N_5736,N_3458,N_3410);
nand U5737 (N_5737,N_3558,N_4349);
nor U5738 (N_5738,N_4225,N_4053);
xor U5739 (N_5739,N_4105,N_3269);
nor U5740 (N_5740,N_3371,N_3388);
nand U5741 (N_5741,N_3443,N_3505);
nor U5742 (N_5742,N_4178,N_3864);
nor U5743 (N_5743,N_3693,N_3549);
nor U5744 (N_5744,N_4477,N_4100);
or U5745 (N_5745,N_3013,N_4118);
xor U5746 (N_5746,N_4170,N_3761);
xor U5747 (N_5747,N_3208,N_4353);
or U5748 (N_5748,N_3997,N_3988);
xor U5749 (N_5749,N_3411,N_3690);
or U5750 (N_5750,N_3495,N_3980);
xor U5751 (N_5751,N_4490,N_4014);
nor U5752 (N_5752,N_3924,N_4451);
xor U5753 (N_5753,N_3839,N_3268);
xnor U5754 (N_5754,N_4108,N_3865);
and U5755 (N_5755,N_3090,N_3064);
nand U5756 (N_5756,N_3241,N_3096);
or U5757 (N_5757,N_4364,N_4427);
nand U5758 (N_5758,N_3146,N_3584);
or U5759 (N_5759,N_3732,N_4064);
nand U5760 (N_5760,N_4230,N_3561);
or U5761 (N_5761,N_3363,N_4195);
or U5762 (N_5762,N_3412,N_4099);
and U5763 (N_5763,N_3563,N_3350);
nand U5764 (N_5764,N_4410,N_3841);
and U5765 (N_5765,N_4193,N_3991);
nand U5766 (N_5766,N_4286,N_3953);
or U5767 (N_5767,N_3512,N_4383);
and U5768 (N_5768,N_3347,N_3677);
xnor U5769 (N_5769,N_3842,N_3747);
nor U5770 (N_5770,N_4379,N_3742);
nor U5771 (N_5771,N_4489,N_3551);
or U5772 (N_5772,N_3505,N_3347);
or U5773 (N_5773,N_3289,N_4409);
and U5774 (N_5774,N_3199,N_3873);
xor U5775 (N_5775,N_4338,N_3536);
xnor U5776 (N_5776,N_3605,N_3848);
xor U5777 (N_5777,N_3232,N_3541);
xor U5778 (N_5778,N_4285,N_3364);
and U5779 (N_5779,N_4160,N_4070);
or U5780 (N_5780,N_3138,N_3223);
or U5781 (N_5781,N_3291,N_3801);
nor U5782 (N_5782,N_4221,N_3138);
nand U5783 (N_5783,N_3317,N_4082);
or U5784 (N_5784,N_3279,N_4473);
nand U5785 (N_5785,N_4033,N_4494);
and U5786 (N_5786,N_4495,N_3341);
and U5787 (N_5787,N_4320,N_3008);
or U5788 (N_5788,N_3311,N_4481);
or U5789 (N_5789,N_3064,N_3305);
xnor U5790 (N_5790,N_4455,N_3643);
or U5791 (N_5791,N_3393,N_3078);
nor U5792 (N_5792,N_3750,N_3506);
nand U5793 (N_5793,N_4490,N_4359);
nand U5794 (N_5794,N_3077,N_3865);
or U5795 (N_5795,N_3316,N_3964);
nand U5796 (N_5796,N_3551,N_3082);
or U5797 (N_5797,N_3683,N_3888);
xor U5798 (N_5798,N_4383,N_3753);
and U5799 (N_5799,N_3594,N_3716);
nand U5800 (N_5800,N_3882,N_3497);
nor U5801 (N_5801,N_3157,N_3414);
nand U5802 (N_5802,N_3410,N_4114);
xor U5803 (N_5803,N_3615,N_3215);
and U5804 (N_5804,N_3965,N_3454);
and U5805 (N_5805,N_4164,N_4370);
nor U5806 (N_5806,N_4032,N_4024);
and U5807 (N_5807,N_4238,N_4480);
xnor U5808 (N_5808,N_3193,N_4329);
xnor U5809 (N_5809,N_4240,N_4229);
nand U5810 (N_5810,N_3940,N_3651);
or U5811 (N_5811,N_3868,N_3485);
xnor U5812 (N_5812,N_3330,N_4072);
or U5813 (N_5813,N_4126,N_3512);
nor U5814 (N_5814,N_4346,N_3401);
or U5815 (N_5815,N_3529,N_3239);
or U5816 (N_5816,N_3238,N_3962);
and U5817 (N_5817,N_4086,N_3467);
xnor U5818 (N_5818,N_3849,N_4269);
nor U5819 (N_5819,N_3146,N_3631);
nand U5820 (N_5820,N_3041,N_4438);
and U5821 (N_5821,N_4255,N_3054);
nand U5822 (N_5822,N_3783,N_3048);
nor U5823 (N_5823,N_3398,N_3214);
nor U5824 (N_5824,N_4418,N_4082);
nor U5825 (N_5825,N_3386,N_3171);
nor U5826 (N_5826,N_4285,N_3113);
or U5827 (N_5827,N_3371,N_3136);
xor U5828 (N_5828,N_4310,N_4045);
or U5829 (N_5829,N_3718,N_3285);
and U5830 (N_5830,N_4427,N_4323);
nand U5831 (N_5831,N_4122,N_3331);
xnor U5832 (N_5832,N_3586,N_4106);
nand U5833 (N_5833,N_3898,N_4320);
nor U5834 (N_5834,N_4390,N_4104);
nand U5835 (N_5835,N_3020,N_4185);
xor U5836 (N_5836,N_3788,N_4389);
xor U5837 (N_5837,N_4204,N_3838);
nor U5838 (N_5838,N_3066,N_3227);
xnor U5839 (N_5839,N_3809,N_3683);
nand U5840 (N_5840,N_3319,N_3024);
and U5841 (N_5841,N_3668,N_4251);
and U5842 (N_5842,N_4097,N_4135);
or U5843 (N_5843,N_3479,N_3781);
nand U5844 (N_5844,N_4440,N_4065);
xor U5845 (N_5845,N_3032,N_4469);
or U5846 (N_5846,N_4436,N_3053);
or U5847 (N_5847,N_4313,N_3323);
nor U5848 (N_5848,N_3720,N_3409);
and U5849 (N_5849,N_3011,N_3316);
or U5850 (N_5850,N_4419,N_3991);
or U5851 (N_5851,N_3849,N_3137);
xor U5852 (N_5852,N_4435,N_3727);
and U5853 (N_5853,N_3673,N_3450);
nand U5854 (N_5854,N_3148,N_3596);
nor U5855 (N_5855,N_3159,N_3716);
nor U5856 (N_5856,N_4445,N_4297);
and U5857 (N_5857,N_4211,N_3295);
xor U5858 (N_5858,N_3709,N_3356);
nand U5859 (N_5859,N_3681,N_3805);
nand U5860 (N_5860,N_3888,N_3405);
nor U5861 (N_5861,N_3803,N_3485);
nand U5862 (N_5862,N_3480,N_3517);
xnor U5863 (N_5863,N_3923,N_4205);
nor U5864 (N_5864,N_3095,N_4319);
nand U5865 (N_5865,N_4371,N_3845);
nor U5866 (N_5866,N_3152,N_3224);
xnor U5867 (N_5867,N_4293,N_3592);
and U5868 (N_5868,N_3958,N_3632);
xnor U5869 (N_5869,N_3716,N_3268);
and U5870 (N_5870,N_3273,N_4081);
nor U5871 (N_5871,N_3383,N_3220);
or U5872 (N_5872,N_4434,N_3206);
xor U5873 (N_5873,N_4079,N_3876);
nor U5874 (N_5874,N_4457,N_3629);
and U5875 (N_5875,N_3401,N_4386);
nand U5876 (N_5876,N_3222,N_4027);
nor U5877 (N_5877,N_4287,N_4496);
or U5878 (N_5878,N_3514,N_4430);
or U5879 (N_5879,N_3688,N_3189);
or U5880 (N_5880,N_3490,N_4122);
and U5881 (N_5881,N_3548,N_3500);
or U5882 (N_5882,N_3490,N_3902);
or U5883 (N_5883,N_3252,N_3364);
and U5884 (N_5884,N_3078,N_4119);
and U5885 (N_5885,N_4036,N_3712);
xnor U5886 (N_5886,N_3095,N_3070);
nand U5887 (N_5887,N_3366,N_3148);
and U5888 (N_5888,N_4440,N_3932);
nand U5889 (N_5889,N_3682,N_4054);
nand U5890 (N_5890,N_3068,N_4395);
nand U5891 (N_5891,N_4266,N_3934);
xor U5892 (N_5892,N_4208,N_3690);
or U5893 (N_5893,N_3562,N_3585);
xnor U5894 (N_5894,N_3581,N_3965);
nand U5895 (N_5895,N_4321,N_3138);
nor U5896 (N_5896,N_4178,N_3922);
and U5897 (N_5897,N_4180,N_3641);
and U5898 (N_5898,N_4074,N_4256);
nand U5899 (N_5899,N_4007,N_3372);
nand U5900 (N_5900,N_4372,N_4178);
nor U5901 (N_5901,N_3810,N_3967);
and U5902 (N_5902,N_4170,N_4153);
or U5903 (N_5903,N_3952,N_3849);
xor U5904 (N_5904,N_3298,N_3227);
xor U5905 (N_5905,N_3377,N_3595);
or U5906 (N_5906,N_3268,N_4265);
and U5907 (N_5907,N_4298,N_4495);
nand U5908 (N_5908,N_3891,N_3788);
nor U5909 (N_5909,N_3780,N_4276);
or U5910 (N_5910,N_3457,N_3873);
or U5911 (N_5911,N_3520,N_4137);
and U5912 (N_5912,N_4453,N_3802);
nand U5913 (N_5913,N_3040,N_3096);
nor U5914 (N_5914,N_3917,N_3973);
or U5915 (N_5915,N_4063,N_3863);
nand U5916 (N_5916,N_3413,N_4119);
and U5917 (N_5917,N_3320,N_3449);
and U5918 (N_5918,N_3410,N_4003);
or U5919 (N_5919,N_3301,N_4116);
xor U5920 (N_5920,N_3638,N_3269);
nor U5921 (N_5921,N_4319,N_4424);
and U5922 (N_5922,N_4373,N_3822);
nand U5923 (N_5923,N_3519,N_4454);
xnor U5924 (N_5924,N_4286,N_3629);
or U5925 (N_5925,N_3109,N_3015);
or U5926 (N_5926,N_3271,N_3594);
xnor U5927 (N_5927,N_3978,N_3125);
nor U5928 (N_5928,N_4402,N_3283);
and U5929 (N_5929,N_3815,N_3653);
xnor U5930 (N_5930,N_3931,N_3737);
nand U5931 (N_5931,N_4211,N_3213);
nand U5932 (N_5932,N_4344,N_3927);
nand U5933 (N_5933,N_3658,N_3324);
xor U5934 (N_5934,N_3012,N_3029);
and U5935 (N_5935,N_3793,N_3226);
nand U5936 (N_5936,N_3693,N_3883);
and U5937 (N_5937,N_3140,N_4338);
xor U5938 (N_5938,N_3850,N_3900);
nand U5939 (N_5939,N_4141,N_4320);
xor U5940 (N_5940,N_3020,N_4395);
or U5941 (N_5941,N_4244,N_3263);
or U5942 (N_5942,N_3175,N_3533);
xnor U5943 (N_5943,N_4178,N_4142);
nand U5944 (N_5944,N_3581,N_3730);
or U5945 (N_5945,N_3495,N_3965);
or U5946 (N_5946,N_4058,N_3554);
or U5947 (N_5947,N_4263,N_3674);
nand U5948 (N_5948,N_4426,N_3933);
nand U5949 (N_5949,N_3904,N_4062);
xnor U5950 (N_5950,N_3188,N_3767);
xor U5951 (N_5951,N_4363,N_3619);
xnor U5952 (N_5952,N_4469,N_4087);
nor U5953 (N_5953,N_3432,N_3010);
nor U5954 (N_5954,N_3850,N_3281);
nor U5955 (N_5955,N_3214,N_3675);
and U5956 (N_5956,N_3379,N_4134);
nand U5957 (N_5957,N_4343,N_4051);
nand U5958 (N_5958,N_3696,N_4188);
or U5959 (N_5959,N_3360,N_4182);
or U5960 (N_5960,N_3910,N_4178);
and U5961 (N_5961,N_4468,N_4066);
or U5962 (N_5962,N_3653,N_4267);
or U5963 (N_5963,N_3736,N_3429);
or U5964 (N_5964,N_3365,N_3719);
xor U5965 (N_5965,N_4159,N_4476);
or U5966 (N_5966,N_3187,N_3032);
nand U5967 (N_5967,N_3586,N_4451);
or U5968 (N_5968,N_3264,N_4138);
and U5969 (N_5969,N_3525,N_3155);
nor U5970 (N_5970,N_3841,N_3647);
or U5971 (N_5971,N_3870,N_3058);
nand U5972 (N_5972,N_3640,N_3748);
nor U5973 (N_5973,N_3535,N_3500);
xor U5974 (N_5974,N_4477,N_4393);
xnor U5975 (N_5975,N_3386,N_4272);
or U5976 (N_5976,N_3349,N_3951);
nor U5977 (N_5977,N_3967,N_3755);
xor U5978 (N_5978,N_3586,N_3716);
xnor U5979 (N_5979,N_3730,N_4144);
xor U5980 (N_5980,N_3596,N_3317);
and U5981 (N_5981,N_3010,N_3712);
or U5982 (N_5982,N_3587,N_3646);
and U5983 (N_5983,N_3506,N_4320);
nand U5984 (N_5984,N_3296,N_3616);
nand U5985 (N_5985,N_3764,N_3467);
and U5986 (N_5986,N_4203,N_4328);
and U5987 (N_5987,N_3964,N_3825);
and U5988 (N_5988,N_3657,N_4059);
and U5989 (N_5989,N_3871,N_3770);
or U5990 (N_5990,N_3940,N_4348);
or U5991 (N_5991,N_3666,N_3753);
xnor U5992 (N_5992,N_4205,N_3535);
and U5993 (N_5993,N_3060,N_3684);
or U5994 (N_5994,N_3498,N_3837);
and U5995 (N_5995,N_3109,N_3241);
xor U5996 (N_5996,N_3946,N_3827);
nor U5997 (N_5997,N_3325,N_3536);
nor U5998 (N_5998,N_3730,N_4497);
nor U5999 (N_5999,N_3882,N_4130);
or U6000 (N_6000,N_4858,N_5739);
nor U6001 (N_6001,N_4679,N_5467);
and U6002 (N_6002,N_5128,N_5170);
xor U6003 (N_6003,N_5534,N_5951);
and U6004 (N_6004,N_5440,N_5411);
nand U6005 (N_6005,N_5610,N_5949);
and U6006 (N_6006,N_5186,N_4928);
and U6007 (N_6007,N_4519,N_4933);
and U6008 (N_6008,N_5259,N_5395);
and U6009 (N_6009,N_5831,N_5102);
and U6010 (N_6010,N_5914,N_5133);
nor U6011 (N_6011,N_5086,N_4775);
nor U6012 (N_6012,N_5427,N_5942);
xor U6013 (N_6013,N_4937,N_5357);
nor U6014 (N_6014,N_5268,N_5124);
and U6015 (N_6015,N_5125,N_4972);
and U6016 (N_6016,N_5466,N_4605);
or U6017 (N_6017,N_5381,N_5185);
and U6018 (N_6018,N_5382,N_5639);
xor U6019 (N_6019,N_5583,N_5813);
nand U6020 (N_6020,N_5296,N_4820);
or U6021 (N_6021,N_5001,N_5577);
xor U6022 (N_6022,N_5607,N_5389);
xnor U6023 (N_6023,N_5498,N_4923);
nor U6024 (N_6024,N_5622,N_5488);
or U6025 (N_6025,N_5580,N_5812);
nand U6026 (N_6026,N_4709,N_4719);
and U6027 (N_6027,N_5334,N_5116);
xnor U6028 (N_6028,N_4506,N_5762);
or U6029 (N_6029,N_5800,N_5645);
xnor U6030 (N_6030,N_4753,N_5307);
nand U6031 (N_6031,N_4992,N_4536);
nand U6032 (N_6032,N_4705,N_5325);
nand U6033 (N_6033,N_4723,N_4703);
and U6034 (N_6034,N_4978,N_4504);
and U6035 (N_6035,N_4843,N_4558);
xor U6036 (N_6036,N_5464,N_4762);
nor U6037 (N_6037,N_4916,N_4982);
and U6038 (N_6038,N_4784,N_4989);
xnor U6039 (N_6039,N_4689,N_4921);
nor U6040 (N_6040,N_5505,N_4793);
nand U6041 (N_6041,N_5141,N_5954);
nor U6042 (N_6042,N_5712,N_5655);
nor U6043 (N_6043,N_4773,N_5683);
or U6044 (N_6044,N_5687,N_4875);
xor U6045 (N_6045,N_5302,N_5794);
nand U6046 (N_6046,N_4897,N_4765);
and U6047 (N_6047,N_4665,N_5333);
or U6048 (N_6048,N_5079,N_5053);
and U6049 (N_6049,N_5595,N_5851);
or U6050 (N_6050,N_5693,N_5659);
nand U6051 (N_6051,N_4654,N_5074);
nand U6052 (N_6052,N_4635,N_5815);
xor U6053 (N_6053,N_5682,N_4850);
nand U6054 (N_6054,N_4788,N_5470);
xnor U6055 (N_6055,N_4701,N_5866);
or U6056 (N_6056,N_5569,N_5448);
nand U6057 (N_6057,N_5088,N_4633);
or U6058 (N_6058,N_4999,N_5328);
or U6059 (N_6059,N_5859,N_5646);
nand U6060 (N_6060,N_5066,N_5450);
nand U6061 (N_6061,N_5413,N_5924);
and U6062 (N_6062,N_4970,N_5153);
nand U6063 (N_6063,N_5211,N_4587);
xor U6064 (N_6064,N_5849,N_5894);
and U6065 (N_6065,N_4981,N_4881);
nor U6066 (N_6066,N_5008,N_4721);
and U6067 (N_6067,N_5027,N_4518);
xor U6068 (N_6068,N_5918,N_4692);
or U6069 (N_6069,N_4706,N_5176);
or U6070 (N_6070,N_5679,N_5308);
nor U6071 (N_6071,N_4994,N_5095);
or U6072 (N_6072,N_4581,N_5516);
xor U6073 (N_6073,N_5403,N_4620);
nor U6074 (N_6074,N_5043,N_4533);
and U6075 (N_6075,N_5675,N_4849);
nor U6076 (N_6076,N_5987,N_4732);
and U6077 (N_6077,N_5097,N_5070);
or U6078 (N_6078,N_4625,N_5255);
xnor U6079 (N_6079,N_4939,N_5637);
and U6080 (N_6080,N_5156,N_5549);
and U6081 (N_6081,N_4597,N_4568);
nand U6082 (N_6082,N_5888,N_4915);
nor U6083 (N_6083,N_5239,N_5269);
nor U6084 (N_6084,N_4935,N_5321);
and U6085 (N_6085,N_5198,N_5537);
and U6086 (N_6086,N_5520,N_5226);
nor U6087 (N_6087,N_5232,N_4895);
and U6088 (N_6088,N_5991,N_5662);
nand U6089 (N_6089,N_5099,N_4754);
xor U6090 (N_6090,N_5768,N_5338);
and U6091 (N_6091,N_5291,N_4808);
xor U6092 (N_6092,N_4799,N_5953);
and U6093 (N_6093,N_4616,N_5451);
xnor U6094 (N_6094,N_5227,N_4795);
nor U6095 (N_6095,N_4546,N_5618);
xor U6096 (N_6096,N_4936,N_5278);
nand U6097 (N_6097,N_4543,N_5028);
xnor U6098 (N_6098,N_5509,N_5363);
xor U6099 (N_6099,N_4867,N_4641);
nor U6100 (N_6100,N_4940,N_5871);
nor U6101 (N_6101,N_5998,N_5624);
xnor U6102 (N_6102,N_4686,N_5472);
xor U6103 (N_6103,N_5779,N_5788);
and U6104 (N_6104,N_4718,N_5643);
xnor U6105 (N_6105,N_4583,N_5592);
or U6106 (N_6106,N_5602,N_5559);
xnor U6107 (N_6107,N_5674,N_5006);
nand U6108 (N_6108,N_4797,N_5535);
xor U6109 (N_6109,N_5290,N_4783);
or U6110 (N_6110,N_5838,N_5658);
nand U6111 (N_6111,N_5225,N_5911);
or U6112 (N_6112,N_5890,N_5260);
nand U6113 (N_6113,N_5140,N_5587);
xnor U6114 (N_6114,N_4963,N_5630);
and U6115 (N_6115,N_5319,N_5243);
nand U6116 (N_6116,N_5927,N_4645);
xor U6117 (N_6117,N_5635,N_4621);
and U6118 (N_6118,N_5702,N_4697);
and U6119 (N_6119,N_5756,N_5523);
nor U6120 (N_6120,N_4555,N_4863);
xnor U6121 (N_6121,N_4856,N_4591);
xor U6122 (N_6122,N_5808,N_5173);
and U6123 (N_6123,N_4685,N_5664);
nor U6124 (N_6124,N_5103,N_4845);
and U6125 (N_6125,N_5500,N_5995);
or U6126 (N_6126,N_5570,N_5294);
nand U6127 (N_6127,N_5874,N_4780);
and U6128 (N_6128,N_5044,N_5390);
nor U6129 (N_6129,N_4903,N_5596);
xnor U6130 (N_6130,N_5482,N_4725);
nand U6131 (N_6131,N_5201,N_5692);
nor U6132 (N_6132,N_5576,N_5743);
or U6133 (N_6133,N_5165,N_5904);
xnor U6134 (N_6134,N_5069,N_5881);
and U6135 (N_6135,N_5256,N_5879);
nand U6136 (N_6136,N_5989,N_4854);
nand U6137 (N_6137,N_4741,N_4855);
nand U6138 (N_6138,N_5555,N_5852);
and U6139 (N_6139,N_4639,N_4510);
nand U6140 (N_6140,N_5356,N_4567);
xor U6141 (N_6141,N_5059,N_5025);
nor U6142 (N_6142,N_5318,N_4693);
nor U6143 (N_6143,N_5967,N_4926);
nor U6144 (N_6144,N_4714,N_5311);
and U6145 (N_6145,N_4729,N_5604);
and U6146 (N_6146,N_5301,N_5912);
nor U6147 (N_6147,N_4914,N_5892);
and U6148 (N_6148,N_5417,N_5016);
or U6149 (N_6149,N_5986,N_5612);
and U6150 (N_6150,N_4660,N_5358);
nand U6151 (N_6151,N_5917,N_4734);
nand U6152 (N_6152,N_4929,N_5522);
nand U6153 (N_6153,N_5137,N_5891);
and U6154 (N_6154,N_5840,N_4826);
and U6155 (N_6155,N_5160,N_5832);
nor U6156 (N_6156,N_4515,N_5210);
xnor U6157 (N_6157,N_5538,N_5617);
and U6158 (N_6158,N_5003,N_5663);
and U6159 (N_6159,N_5494,N_5396);
or U6160 (N_6160,N_4707,N_5309);
nor U6161 (N_6161,N_5588,N_5366);
nand U6162 (N_6162,N_5770,N_4545);
nand U6163 (N_6163,N_5452,N_4526);
nor U6164 (N_6164,N_5551,N_5857);
or U6165 (N_6165,N_5684,N_5741);
nor U6166 (N_6166,N_5340,N_4873);
and U6167 (N_6167,N_5531,N_5856);
nand U6168 (N_6168,N_5910,N_4861);
and U6169 (N_6169,N_4758,N_4987);
xor U6170 (N_6170,N_5429,N_4918);
and U6171 (N_6171,N_5096,N_5067);
or U6172 (N_6172,N_5332,N_5005);
and U6173 (N_6173,N_5957,N_5694);
nor U6174 (N_6174,N_5872,N_4742);
and U6175 (N_6175,N_5385,N_4727);
and U6176 (N_6176,N_5771,N_5354);
xor U6177 (N_6177,N_5816,N_5039);
nor U6178 (N_6178,N_5335,N_5804);
nand U6179 (N_6179,N_5324,N_5401);
nand U6180 (N_6180,N_4737,N_5169);
nand U6181 (N_6181,N_5937,N_5966);
or U6182 (N_6182,N_4521,N_4925);
nand U6183 (N_6183,N_5886,N_4818);
xnor U6184 (N_6184,N_4930,N_5492);
nor U6185 (N_6185,N_5697,N_5152);
and U6186 (N_6186,N_4927,N_5218);
nor U6187 (N_6187,N_5721,N_4954);
or U6188 (N_6188,N_5188,N_5080);
nand U6189 (N_6189,N_5248,N_4640);
nor U6190 (N_6190,N_4576,N_5519);
or U6191 (N_6191,N_4817,N_5458);
nor U6192 (N_6192,N_4604,N_5187);
nand U6193 (N_6193,N_5971,N_5252);
or U6194 (N_6194,N_5347,N_4595);
or U6195 (N_6195,N_5719,N_4752);
nor U6196 (N_6196,N_4547,N_5030);
xor U6197 (N_6197,N_5056,N_5035);
nor U6198 (N_6198,N_5359,N_4827);
nand U6199 (N_6199,N_4539,N_5199);
xor U6200 (N_6200,N_5154,N_4893);
and U6201 (N_6201,N_5566,N_5364);
xor U6202 (N_6202,N_5980,N_5548);
nor U6203 (N_6203,N_4919,N_4749);
and U6204 (N_6204,N_5757,N_5705);
or U6205 (N_6205,N_4699,N_5192);
xor U6206 (N_6206,N_4938,N_4663);
nor U6207 (N_6207,N_5456,N_4892);
nor U6208 (N_6208,N_4866,N_5484);
nor U6209 (N_6209,N_5718,N_5327);
nor U6210 (N_6210,N_5072,N_4674);
and U6211 (N_6211,N_4672,N_5700);
nand U6212 (N_6212,N_4606,N_5959);
xor U6213 (N_6213,N_5541,N_4636);
or U6214 (N_6214,N_4659,N_5446);
nor U6215 (N_6215,N_4608,N_4713);
or U6216 (N_6216,N_5497,N_5399);
xor U6217 (N_6217,N_5809,N_5796);
xnor U6218 (N_6218,N_5501,N_4750);
or U6219 (N_6219,N_4891,N_5207);
xnor U6220 (N_6220,N_5214,N_5597);
nor U6221 (N_6221,N_5283,N_5078);
nand U6222 (N_6222,N_5323,N_4957);
and U6223 (N_6223,N_5932,N_5825);
or U6224 (N_6224,N_5392,N_4744);
xnor U6225 (N_6225,N_5341,N_4973);
nand U6226 (N_6226,N_5454,N_5530);
or U6227 (N_6227,N_5860,N_5121);
nor U6228 (N_6228,N_5626,N_5021);
nor U6229 (N_6229,N_5876,N_4680);
and U6230 (N_6230,N_4804,N_5644);
nand U6231 (N_6231,N_5415,N_4724);
or U6232 (N_6232,N_4759,N_5046);
nor U6233 (N_6233,N_4614,N_5163);
xor U6234 (N_6234,N_4968,N_5715);
and U6235 (N_6235,N_5270,N_4800);
nor U6236 (N_6236,N_4880,N_5913);
and U6237 (N_6237,N_5230,N_5921);
xnor U6238 (N_6238,N_5142,N_5640);
nand U6239 (N_6239,N_5360,N_5887);
nand U6240 (N_6240,N_5704,N_5854);
xnor U6241 (N_6241,N_5556,N_4556);
nor U6242 (N_6242,N_5634,N_4810);
and U6243 (N_6243,N_5579,N_5691);
or U6244 (N_6244,N_5985,N_5714);
nor U6245 (N_6245,N_4986,N_4971);
xnor U6246 (N_6246,N_5571,N_4998);
or U6247 (N_6247,N_4888,N_4805);
or U6248 (N_6248,N_4761,N_5463);
nand U6249 (N_6249,N_5155,N_4691);
nand U6250 (N_6250,N_4535,N_5666);
nand U6251 (N_6251,N_5740,N_5112);
nor U6252 (N_6252,N_4600,N_5736);
and U6253 (N_6253,N_5013,N_5065);
and U6254 (N_6254,N_5614,N_4711);
or U6255 (N_6255,N_5233,N_5349);
nor U6256 (N_6256,N_4523,N_5981);
xnor U6257 (N_6257,N_5436,N_5996);
and U6258 (N_6258,N_5062,N_5204);
or U6259 (N_6259,N_5805,N_5814);
nor U6260 (N_6260,N_5249,N_5508);
nand U6261 (N_6261,N_5561,N_5212);
xor U6262 (N_6262,N_5157,N_5903);
or U6263 (N_6263,N_5976,N_5055);
xor U6264 (N_6264,N_5336,N_5082);
nor U6265 (N_6265,N_5843,N_4630);
xor U6266 (N_6266,N_4859,N_5940);
and U6267 (N_6267,N_5772,N_5421);
xor U6268 (N_6268,N_5798,N_5222);
nor U6269 (N_6269,N_5136,N_5973);
nor U6270 (N_6270,N_5897,N_4842);
or U6271 (N_6271,N_4599,N_4760);
or U6272 (N_6272,N_5629,N_5761);
nor U6273 (N_6273,N_5869,N_5650);
xnor U6274 (N_6274,N_4648,N_5784);
nand U6275 (N_6275,N_5706,N_5305);
or U6276 (N_6276,N_5513,N_4733);
and U6277 (N_6277,N_5134,N_5480);
and U6278 (N_6278,N_5900,N_5829);
and U6279 (N_6279,N_4561,N_4509);
nor U6280 (N_6280,N_4746,N_5628);
and U6281 (N_6281,N_5208,N_5696);
nor U6282 (N_6282,N_5594,N_5581);
xnor U6283 (N_6283,N_5443,N_5707);
xor U6284 (N_6284,N_5999,N_5130);
xor U6285 (N_6285,N_4534,N_5827);
nand U6286 (N_6286,N_5111,N_5060);
and U6287 (N_6287,N_5101,N_5958);
nor U6288 (N_6288,N_5388,N_5532);
xnor U6289 (N_6289,N_4979,N_5368);
nand U6290 (N_6290,N_4774,N_4670);
nand U6291 (N_6291,N_5909,N_5320);
nor U6292 (N_6292,N_4769,N_5179);
nor U6293 (N_6293,N_4990,N_5282);
or U6294 (N_6294,N_4934,N_5884);
nor U6295 (N_6295,N_4531,N_5115);
xor U6296 (N_6296,N_4965,N_5084);
and U6297 (N_6297,N_4823,N_5286);
nand U6298 (N_6298,N_5708,N_5284);
or U6299 (N_6299,N_4794,N_4988);
or U6300 (N_6300,N_5135,N_4557);
and U6301 (N_6301,N_5605,N_5203);
xor U6302 (N_6302,N_5022,N_5750);
xor U6303 (N_6303,N_5017,N_5713);
xnor U6304 (N_6304,N_5978,N_4951);
xnor U6305 (N_6305,N_5783,N_4768);
nand U6306 (N_6306,N_4624,N_5939);
xor U6307 (N_6307,N_5168,N_5455);
and U6308 (N_6308,N_4688,N_5058);
xnor U6309 (N_6309,N_5528,N_5002);
nand U6310 (N_6310,N_5337,N_5342);
or U6311 (N_6311,N_5235,N_4816);
nand U6312 (N_6312,N_5710,N_5240);
nand U6313 (N_6313,N_5882,N_5351);
xor U6314 (N_6314,N_4920,N_5582);
or U6315 (N_6315,N_5295,N_5004);
nor U6316 (N_6316,N_5469,N_4590);
xnor U6317 (N_6317,N_5507,N_5041);
nand U6318 (N_6318,N_5398,N_4564);
or U6319 (N_6319,N_4739,N_4887);
nand U6320 (N_6320,N_5310,N_4646);
nand U6321 (N_6321,N_5853,N_4908);
and U6322 (N_6322,N_4682,N_5150);
xnor U6323 (N_6323,N_5251,N_4618);
nor U6324 (N_6324,N_5375,N_5438);
xor U6325 (N_6325,N_4767,N_5386);
or U6326 (N_6326,N_5730,N_5114);
nor U6327 (N_6327,N_4772,N_5754);
and U6328 (N_6328,N_5083,N_5547);
xnor U6329 (N_6329,N_5638,N_5842);
or U6330 (N_6330,N_5174,N_5956);
nand U6331 (N_6331,N_5824,N_5720);
and U6332 (N_6332,N_5405,N_5120);
xnor U6333 (N_6333,N_4868,N_5619);
and U6334 (N_6334,N_5493,N_5304);
nor U6335 (N_6335,N_5071,N_4851);
and U6336 (N_6336,N_5274,N_4985);
or U6337 (N_6337,N_5425,N_5540);
or U6338 (N_6338,N_5032,N_5938);
or U6339 (N_6339,N_4809,N_5416);
nand U6340 (N_6340,N_5830,N_4550);
xor U6341 (N_6341,N_4796,N_5117);
nor U6342 (N_6342,N_5428,N_4596);
or U6343 (N_6343,N_5807,N_5355);
or U6344 (N_6344,N_5262,N_5974);
xor U6345 (N_6345,N_4756,N_4650);
or U6346 (N_6346,N_4694,N_5961);
or U6347 (N_6347,N_5503,N_4637);
nand U6348 (N_6348,N_5131,N_5919);
xor U6349 (N_6349,N_4704,N_5045);
nand U6350 (N_6350,N_5544,N_4528);
or U6351 (N_6351,N_4601,N_5733);
or U6352 (N_6352,N_4955,N_4983);
and U6353 (N_6353,N_4502,N_5975);
and U6354 (N_6354,N_4984,N_5196);
nand U6355 (N_6355,N_4513,N_4511);
nand U6356 (N_6356,N_5620,N_4906);
nand U6357 (N_6357,N_4743,N_4722);
or U6358 (N_6358,N_5652,N_4589);
and U6359 (N_6359,N_5246,N_4898);
nand U6360 (N_6360,N_5087,N_4785);
nand U6361 (N_6361,N_4993,N_4664);
nor U6362 (N_6362,N_5007,N_5667);
nor U6363 (N_6363,N_4837,N_5747);
nand U6364 (N_6364,N_5015,N_5344);
xor U6365 (N_6365,N_5977,N_5461);
nand U6366 (N_6366,N_4948,N_5799);
and U6367 (N_6367,N_5526,N_5864);
nand U6368 (N_6368,N_5611,N_5312);
nand U6369 (N_6369,N_5834,N_5093);
nand U6370 (N_6370,N_5433,N_5345);
or U6371 (N_6371,N_5901,N_4889);
nand U6372 (N_6372,N_5616,N_5791);
and U6373 (N_6373,N_5431,N_5209);
nor U6374 (N_6374,N_4966,N_4819);
xnor U6375 (N_6375,N_5510,N_4871);
nor U6376 (N_6376,N_5326,N_5313);
xor U6377 (N_6377,N_5376,N_5647);
nor U6378 (N_6378,N_5786,N_5902);
and U6379 (N_6379,N_4671,N_5092);
and U6380 (N_6380,N_5023,N_5264);
nor U6381 (N_6381,N_5293,N_5589);
and U6382 (N_6382,N_4755,N_4501);
and U6383 (N_6383,N_4735,N_5042);
nand U6384 (N_6384,N_5515,N_5627);
nor U6385 (N_6385,N_4790,N_5374);
nand U6386 (N_6386,N_5877,N_5603);
and U6387 (N_6387,N_5499,N_5393);
nand U6388 (N_6388,N_5495,N_5823);
nand U6389 (N_6389,N_5346,N_5898);
nor U6390 (N_6390,N_5766,N_5839);
nor U6391 (N_6391,N_4952,N_4628);
and U6392 (N_6392,N_5167,N_5370);
xor U6393 (N_6393,N_4668,N_4976);
and U6394 (N_6394,N_5126,N_4570);
nand U6395 (N_6395,N_5184,N_4537);
nand U6396 (N_6396,N_4500,N_5723);
nor U6397 (N_6397,N_5936,N_5468);
and U6398 (N_6398,N_5931,N_4922);
or U6399 (N_6399,N_5946,N_5190);
nand U6400 (N_6400,N_5514,N_5699);
nor U6401 (N_6401,N_5565,N_5965);
xnor U6402 (N_6402,N_4638,N_5631);
xor U6403 (N_6403,N_5298,N_4977);
and U6404 (N_6404,N_5933,N_5845);
xor U6405 (N_6405,N_4840,N_5752);
xor U6406 (N_6406,N_4807,N_4830);
nand U6407 (N_6407,N_4559,N_5238);
nand U6408 (N_6408,N_5867,N_5462);
nor U6409 (N_6409,N_5836,N_5297);
and U6410 (N_6410,N_5279,N_4588);
and U6411 (N_6411,N_4740,N_5024);
and U6412 (N_6412,N_5223,N_5362);
nand U6413 (N_6413,N_5600,N_4931);
and U6414 (N_6414,N_4812,N_4996);
nor U6415 (N_6415,N_4777,N_5195);
nor U6416 (N_6416,N_4757,N_5123);
nand U6417 (N_6417,N_5292,N_4514);
and U6418 (N_6418,N_5474,N_5726);
or U6419 (N_6419,N_5010,N_5929);
nor U6420 (N_6420,N_5317,N_4806);
xor U6421 (N_6421,N_5018,N_5599);
xor U6422 (N_6422,N_5460,N_4832);
nand U6423 (N_6423,N_5764,N_5780);
nor U6424 (N_6424,N_4690,N_5907);
nor U6425 (N_6425,N_4852,N_4609);
or U6426 (N_6426,N_4626,N_5844);
nand U6427 (N_6427,N_5916,N_5506);
or U6428 (N_6428,N_4698,N_4870);
xor U6429 (N_6429,N_5748,N_4932);
or U6430 (N_6430,N_4838,N_4874);
and U6431 (N_6431,N_4766,N_5435);
nand U6432 (N_6432,N_5709,N_5502);
xnor U6433 (N_6433,N_5486,N_5878);
and U6434 (N_6434,N_4508,N_4560);
xnor U6435 (N_6435,N_5855,N_5406);
xnor U6436 (N_6436,N_5552,N_5928);
xor U6437 (N_6437,N_5012,N_5266);
nor U6438 (N_6438,N_5068,N_5533);
nand U6439 (N_6439,N_4909,N_5331);
nand U6440 (N_6440,N_5491,N_5686);
or U6441 (N_6441,N_5963,N_5811);
nand U6442 (N_6442,N_5665,N_5343);
nand U6443 (N_6443,N_4789,N_4779);
and U6444 (N_6444,N_4945,N_4611);
nor U6445 (N_6445,N_5109,N_5820);
or U6446 (N_6446,N_5833,N_5972);
nor U6447 (N_6447,N_4613,N_5930);
and U6448 (N_6448,N_4771,N_5690);
nor U6449 (N_6449,N_5171,N_5127);
or U6450 (N_6450,N_5081,N_5288);
nand U6451 (N_6451,N_5402,N_5689);
or U6452 (N_6452,N_5164,N_4894);
xor U6453 (N_6453,N_5372,N_5100);
nor U6454 (N_6454,N_4554,N_5162);
and U6455 (N_6455,N_4846,N_5329);
nor U6456 (N_6456,N_4917,N_4549);
nand U6457 (N_6457,N_4708,N_5870);
or U6458 (N_6458,N_5899,N_5228);
nand U6459 (N_6459,N_5383,N_5773);
or U6460 (N_6460,N_5553,N_5229);
nand U6461 (N_6461,N_5738,N_5414);
xnor U6462 (N_6462,N_5822,N_4553);
or U6463 (N_6463,N_5019,N_4520);
nor U6464 (N_6464,N_5057,N_5189);
and U6465 (N_6465,N_4666,N_5968);
xnor U6466 (N_6466,N_4675,N_5680);
and U6467 (N_6467,N_5471,N_5089);
and U6468 (N_6468,N_5273,N_4726);
xnor U6469 (N_6469,N_5848,N_5982);
xor U6470 (N_6470,N_5789,N_4667);
nor U6471 (N_6471,N_5219,N_5090);
nand U6472 (N_6472,N_4833,N_5180);
and U6473 (N_6473,N_4786,N_5560);
nor U6474 (N_6474,N_4730,N_5423);
xor U6475 (N_6475,N_5653,N_5785);
xor U6476 (N_6476,N_4728,N_5161);
or U6477 (N_6477,N_5145,N_5642);
and U6478 (N_6478,N_5847,N_5512);
xnor U6479 (N_6479,N_5200,N_5182);
or U6480 (N_6480,N_5765,N_4622);
nand U6481 (N_6481,N_5479,N_4619);
nor U6482 (N_6482,N_5073,N_4731);
nand U6483 (N_6483,N_4839,N_4967);
nor U6484 (N_6484,N_4864,N_5197);
xor U6485 (N_6485,N_4824,N_5177);
xnor U6486 (N_6486,N_5420,N_5969);
nor U6487 (N_6487,N_4695,N_4944);
nand U6488 (N_6488,N_4592,N_4673);
nand U6489 (N_6489,N_5782,N_4647);
nand U6490 (N_6490,N_5330,N_5988);
nor U6491 (N_6491,N_5749,N_4853);
and U6492 (N_6492,N_5430,N_5496);
xor U6493 (N_6493,N_5670,N_4907);
and U6494 (N_6494,N_5801,N_4814);
and U6495 (N_6495,N_4503,N_5118);
xnor U6496 (N_6496,N_5194,N_4649);
or U6497 (N_6497,N_5408,N_5862);
xor U6498 (N_6498,N_4676,N_4995);
xnor U6499 (N_6499,N_5792,N_5826);
nand U6500 (N_6500,N_5545,N_4947);
nor U6501 (N_6501,N_5806,N_5483);
nor U6502 (N_6502,N_5418,N_5660);
xnor U6503 (N_6503,N_5525,N_4538);
xor U6504 (N_6504,N_4569,N_4763);
xor U6505 (N_6505,N_4551,N_5945);
nor U6506 (N_6506,N_5668,N_4961);
nand U6507 (N_6507,N_4904,N_5992);
nor U6508 (N_6508,N_5955,N_5373);
nand U6509 (N_6509,N_5960,N_5557);
nor U6510 (N_6510,N_4634,N_4530);
xnor U6511 (N_6511,N_4662,N_4844);
nand U6512 (N_6512,N_5465,N_5567);
nand U6513 (N_6513,N_5703,N_5191);
xor U6514 (N_6514,N_4629,N_4958);
nand U6515 (N_6515,N_5776,N_5231);
or U6516 (N_6516,N_5352,N_5026);
nand U6517 (N_6517,N_5701,N_5573);
or U6518 (N_6518,N_5850,N_5224);
and U6519 (N_6519,N_5014,N_5106);
or U6520 (N_6520,N_4542,N_4571);
and U6521 (N_6521,N_4862,N_5104);
and U6522 (N_6522,N_4885,N_5529);
xnor U6523 (N_6523,N_5064,N_5220);
nand U6524 (N_6524,N_5289,N_5367);
and U6525 (N_6525,N_5034,N_5148);
nand U6526 (N_6526,N_5656,N_5725);
nand U6527 (N_6527,N_5205,N_5263);
nand U6528 (N_6528,N_5094,N_4677);
or U6529 (N_6529,N_4798,N_5077);
nand U6530 (N_6530,N_5558,N_4716);
and U6531 (N_6531,N_4577,N_5281);
or U6532 (N_6532,N_4525,N_5795);
and U6533 (N_6533,N_5299,N_4524);
nor U6534 (N_6534,N_5361,N_5432);
nand U6535 (N_6535,N_4835,N_4575);
nand U6536 (N_6536,N_5202,N_4579);
nand U6537 (N_6537,N_5050,N_5818);
xnor U6538 (N_6538,N_5950,N_4529);
xnor U6539 (N_6539,N_4782,N_4747);
xnor U6540 (N_6540,N_5477,N_5242);
nand U6541 (N_6541,N_4941,N_5758);
xnor U6542 (N_6542,N_5457,N_5138);
xnor U6543 (N_6543,N_5377,N_5896);
and U6544 (N_6544,N_5893,N_4738);
and U6545 (N_6545,N_5728,N_4953);
and U6546 (N_6546,N_5217,N_5731);
xor U6547 (N_6547,N_5445,N_4610);
nand U6548 (N_6548,N_5672,N_5300);
nand U6549 (N_6549,N_5915,N_4959);
and U6550 (N_6550,N_5441,N_4623);
and U6551 (N_6551,N_5206,N_4834);
and U6552 (N_6552,N_4803,N_5265);
xor U6553 (N_6553,N_4651,N_5245);
or U6554 (N_6554,N_5371,N_4578);
and U6555 (N_6555,N_5504,N_5817);
nor U6556 (N_6556,N_4653,N_5623);
or U6557 (N_6557,N_4710,N_5122);
xnor U6558 (N_6558,N_4778,N_5048);
nor U6559 (N_6559,N_5271,N_4681);
or U6560 (N_6560,N_4631,N_4602);
xnor U6561 (N_6561,N_5178,N_5407);
nor U6562 (N_6562,N_5810,N_4687);
xor U6563 (N_6563,N_5287,N_5669);
xnor U6564 (N_6564,N_5119,N_5984);
and U6565 (N_6565,N_5047,N_5033);
nor U6566 (N_6566,N_5895,N_5397);
nand U6567 (N_6567,N_5625,N_4912);
xnor U6568 (N_6568,N_5722,N_5585);
nor U6569 (N_6569,N_5316,N_5979);
xnor U6570 (N_6570,N_5803,N_5753);
or U6571 (N_6571,N_4975,N_4900);
xor U6572 (N_6572,N_4905,N_4882);
nand U6573 (N_6573,N_5517,N_4962);
and U6574 (N_6574,N_5846,N_4960);
nand U6575 (N_6575,N_5020,N_5651);
nand U6576 (N_6576,N_4715,N_5964);
or U6577 (N_6577,N_5146,N_5254);
nor U6578 (N_6578,N_5590,N_5213);
or U6579 (N_6579,N_4828,N_5598);
xnor U6580 (N_6580,N_5378,N_5875);
nor U6581 (N_6581,N_5241,N_5654);
xnor U6582 (N_6582,N_5926,N_5554);
and U6583 (N_6583,N_5944,N_5661);
nand U6584 (N_6584,N_5419,N_5036);
or U6585 (N_6585,N_4522,N_4632);
nor U6586 (N_6586,N_5948,N_4781);
nand U6587 (N_6587,N_5485,N_5920);
xor U6588 (N_6588,N_4517,N_4787);
or U6589 (N_6589,N_4573,N_5863);
or U6590 (N_6590,N_5835,N_5437);
and U6591 (N_6591,N_5609,N_5993);
nand U6592 (N_6592,N_5139,N_4815);
nor U6593 (N_6593,N_5166,N_4548);
nor U6594 (N_6594,N_5657,N_4644);
nand U6595 (N_6595,N_5105,N_5673);
or U6596 (N_6596,N_4607,N_5524);
nand U6597 (N_6597,N_5970,N_4831);
xnor U6598 (N_6598,N_5601,N_4910);
xnor U6599 (N_6599,N_5676,N_5075);
xor U6600 (N_6600,N_5280,N_5449);
xnor U6601 (N_6601,N_4764,N_5369);
or U6602 (N_6602,N_5621,N_5574);
xnor U6603 (N_6603,N_5108,N_5434);
and U6604 (N_6604,N_4980,N_5444);
nor U6605 (N_6605,N_5787,N_4883);
nand U6606 (N_6606,N_5221,N_5775);
or U6607 (N_6607,N_4776,N_4642);
and U6608 (N_6608,N_5732,N_5935);
nor U6609 (N_6609,N_5841,N_5591);
nor U6610 (N_6610,N_5129,N_4997);
and U6611 (N_6611,N_4745,N_5883);
and U6612 (N_6612,N_5459,N_5677);
nand U6613 (N_6613,N_4655,N_5353);
xor U6614 (N_6614,N_5038,N_5040);
nand U6615 (N_6615,N_5681,N_5257);
or U6616 (N_6616,N_5404,N_5426);
xor U6617 (N_6617,N_5481,N_5439);
nand U6618 (N_6618,N_5442,N_5678);
xnor U6619 (N_6619,N_4552,N_5511);
nor U6620 (N_6620,N_5215,N_5098);
nor U6621 (N_6621,N_4678,N_5061);
or U6622 (N_6622,N_5906,N_4991);
nor U6623 (N_6623,N_5339,N_5054);
or U6624 (N_6624,N_4857,N_4562);
nor U6625 (N_6625,N_5608,N_4507);
and U6626 (N_6626,N_4791,N_4949);
nand U6627 (N_6627,N_5085,N_5615);
or U6628 (N_6628,N_5158,N_5037);
xor U6629 (N_6629,N_5941,N_5518);
and U6630 (N_6630,N_5063,N_4911);
or U6631 (N_6631,N_4901,N_5267);
xnor U6632 (N_6632,N_5350,N_5724);
or U6633 (N_6633,N_4913,N_4748);
xor U6634 (N_6634,N_5997,N_5143);
nand U6635 (N_6635,N_5234,N_4878);
or U6636 (N_6636,N_5751,N_5029);
nor U6637 (N_6637,N_5943,N_5922);
nand U6638 (N_6638,N_4702,N_4860);
nor U6639 (N_6639,N_5536,N_4802);
nand U6640 (N_6640,N_4540,N_5322);
and U6641 (N_6641,N_5905,N_5760);
nor U6642 (N_6642,N_5315,N_4505);
xor U6643 (N_6643,N_5688,N_5737);
nand U6644 (N_6644,N_5778,N_5990);
nor U6645 (N_6645,N_5563,N_5181);
xnor U6646 (N_6646,N_5562,N_5542);
xnor U6647 (N_6647,N_5584,N_5698);
nor U6648 (N_6648,N_5729,N_5755);
and U6649 (N_6649,N_4544,N_5193);
xor U6650 (N_6650,N_5889,N_5384);
and U6651 (N_6651,N_5543,N_4879);
nor U6652 (N_6652,N_5572,N_5671);
and U6653 (N_6653,N_5285,N_5952);
xor U6654 (N_6654,N_4736,N_5648);
nor U6655 (N_6655,N_5606,N_5476);
nor U6656 (N_6656,N_4683,N_4574);
xor U6657 (N_6657,N_5880,N_4751);
nand U6658 (N_6658,N_5409,N_4884);
and U6659 (N_6659,N_4829,N_5447);
nand U6660 (N_6660,N_5769,N_5633);
xor U6661 (N_6661,N_5641,N_5632);
or U6662 (N_6662,N_4956,N_5873);
nor U6663 (N_6663,N_5487,N_4684);
xnor U6664 (N_6664,N_4974,N_4964);
nand U6665 (N_6665,N_5000,N_5868);
and U6666 (N_6666,N_5424,N_5717);
xor U6667 (N_6667,N_4872,N_5781);
nand U6668 (N_6668,N_5746,N_5236);
nand U6669 (N_6669,N_5858,N_4661);
nand U6670 (N_6670,N_4586,N_4627);
nand U6671 (N_6671,N_4847,N_4594);
xor U6672 (N_6672,N_4617,N_4792);
xor U6673 (N_6673,N_5253,N_5151);
xnor U6674 (N_6674,N_5716,N_5790);
or U6675 (N_6675,N_5303,N_5802);
nor U6676 (N_6676,N_4582,N_5400);
nand U6677 (N_6677,N_4565,N_5819);
and U6678 (N_6678,N_5489,N_4822);
and U6679 (N_6679,N_5091,N_5276);
nand U6680 (N_6680,N_4696,N_4532);
nor U6681 (N_6681,N_5149,N_4700);
and U6682 (N_6682,N_5272,N_4886);
nand U6683 (N_6683,N_5183,N_5478);
xor U6684 (N_6684,N_5261,N_4821);
nand U6685 (N_6685,N_5237,N_5742);
and U6686 (N_6686,N_4811,N_4669);
nand U6687 (N_6687,N_4876,N_4652);
or U6688 (N_6688,N_5379,N_4598);
and U6689 (N_6689,N_5410,N_5394);
or U6690 (N_6690,N_5113,N_5777);
xor U6691 (N_6691,N_4585,N_5132);
and U6692 (N_6692,N_5216,N_4896);
nand U6693 (N_6693,N_5076,N_5051);
and U6694 (N_6694,N_5348,N_4712);
xor U6695 (N_6695,N_4836,N_4657);
nand U6696 (N_6696,N_5797,N_5962);
nor U6697 (N_6697,N_5147,N_5247);
or U6698 (N_6698,N_5052,N_5412);
nand U6699 (N_6699,N_5277,N_4825);
xor U6700 (N_6700,N_4572,N_4943);
nor U6701 (N_6701,N_5110,N_4877);
xnor U6702 (N_6702,N_4516,N_5711);
nor U6703 (N_6703,N_4841,N_4584);
and U6704 (N_6704,N_4899,N_4946);
xor U6705 (N_6705,N_5527,N_5885);
nor U6706 (N_6706,N_5865,N_5244);
xor U6707 (N_6707,N_5821,N_5774);
xnor U6708 (N_6708,N_5763,N_5314);
nor U6709 (N_6709,N_5994,N_5745);
or U6710 (N_6710,N_5172,N_5793);
xnor U6711 (N_6711,N_5490,N_5744);
xnor U6712 (N_6712,N_5049,N_5009);
xnor U6713 (N_6713,N_4869,N_5387);
nor U6714 (N_6714,N_4612,N_5250);
or U6715 (N_6715,N_4902,N_5275);
nand U6716 (N_6716,N_5031,N_5695);
nand U6717 (N_6717,N_5011,N_5828);
nor U6718 (N_6718,N_5947,N_5306);
and U6719 (N_6719,N_5391,N_4658);
xnor U6720 (N_6720,N_4580,N_5578);
or U6721 (N_6721,N_5759,N_4603);
nand U6722 (N_6722,N_4813,N_5473);
and U6723 (N_6723,N_4527,N_5107);
or U6724 (N_6724,N_4656,N_5586);
or U6725 (N_6725,N_4770,N_5380);
and U6726 (N_6726,N_5685,N_5923);
or U6727 (N_6727,N_5908,N_5539);
or U6728 (N_6728,N_5546,N_4890);
and U6729 (N_6729,N_4563,N_5521);
and U6730 (N_6730,N_4848,N_5144);
nor U6731 (N_6731,N_4942,N_5649);
and U6732 (N_6732,N_5613,N_5550);
nand U6733 (N_6733,N_4865,N_5734);
or U6734 (N_6734,N_5735,N_5727);
and U6735 (N_6735,N_5175,N_5568);
nor U6736 (N_6736,N_5453,N_4720);
nand U6737 (N_6737,N_4950,N_5475);
xnor U6738 (N_6738,N_5365,N_5159);
or U6739 (N_6739,N_5837,N_5767);
and U6740 (N_6740,N_4512,N_4593);
or U6741 (N_6741,N_5422,N_4566);
nand U6742 (N_6742,N_5861,N_5636);
xor U6743 (N_6743,N_4969,N_4643);
or U6744 (N_6744,N_5564,N_5925);
or U6745 (N_6745,N_5934,N_5593);
xnor U6746 (N_6746,N_5258,N_4924);
nand U6747 (N_6747,N_4717,N_4615);
nor U6748 (N_6748,N_4801,N_5983);
nand U6749 (N_6749,N_5575,N_4541);
or U6750 (N_6750,N_5616,N_5396);
nor U6751 (N_6751,N_5339,N_4577);
xnor U6752 (N_6752,N_5968,N_5007);
xnor U6753 (N_6753,N_4594,N_5956);
or U6754 (N_6754,N_5773,N_5175);
nor U6755 (N_6755,N_5174,N_5371);
or U6756 (N_6756,N_4711,N_4962);
or U6757 (N_6757,N_5237,N_4788);
nand U6758 (N_6758,N_4593,N_5729);
nand U6759 (N_6759,N_5022,N_4823);
nand U6760 (N_6760,N_4833,N_5071);
nand U6761 (N_6761,N_5340,N_5910);
nand U6762 (N_6762,N_5755,N_5221);
xnor U6763 (N_6763,N_4812,N_5140);
xor U6764 (N_6764,N_5936,N_5786);
nand U6765 (N_6765,N_5260,N_5510);
nand U6766 (N_6766,N_5530,N_5219);
nand U6767 (N_6767,N_5997,N_5337);
xnor U6768 (N_6768,N_5818,N_5826);
nand U6769 (N_6769,N_5836,N_5056);
nand U6770 (N_6770,N_5933,N_5148);
nand U6771 (N_6771,N_4966,N_4737);
and U6772 (N_6772,N_4659,N_5465);
or U6773 (N_6773,N_5174,N_4551);
and U6774 (N_6774,N_4641,N_5451);
nor U6775 (N_6775,N_5251,N_4510);
and U6776 (N_6776,N_5117,N_4623);
xnor U6777 (N_6777,N_5132,N_5442);
nand U6778 (N_6778,N_4815,N_5415);
and U6779 (N_6779,N_5203,N_5396);
nor U6780 (N_6780,N_4788,N_4895);
nor U6781 (N_6781,N_4925,N_4899);
nand U6782 (N_6782,N_5526,N_4723);
nor U6783 (N_6783,N_5565,N_4928);
and U6784 (N_6784,N_5438,N_4761);
or U6785 (N_6785,N_4811,N_5568);
or U6786 (N_6786,N_4992,N_5154);
nor U6787 (N_6787,N_5407,N_5666);
nand U6788 (N_6788,N_5408,N_5700);
nand U6789 (N_6789,N_5516,N_5795);
nor U6790 (N_6790,N_4593,N_4950);
xnor U6791 (N_6791,N_5440,N_4595);
and U6792 (N_6792,N_4658,N_5566);
nor U6793 (N_6793,N_5992,N_5963);
nor U6794 (N_6794,N_5905,N_4822);
nor U6795 (N_6795,N_5096,N_5126);
nor U6796 (N_6796,N_5535,N_5762);
xnor U6797 (N_6797,N_5323,N_5626);
or U6798 (N_6798,N_5346,N_5590);
nand U6799 (N_6799,N_5546,N_5034);
or U6800 (N_6800,N_4541,N_4818);
nor U6801 (N_6801,N_5026,N_5039);
nand U6802 (N_6802,N_4521,N_4718);
nor U6803 (N_6803,N_4721,N_4506);
nand U6804 (N_6804,N_5322,N_4521);
nand U6805 (N_6805,N_4899,N_5185);
xnor U6806 (N_6806,N_4804,N_4681);
xor U6807 (N_6807,N_5249,N_5729);
xnor U6808 (N_6808,N_5763,N_5206);
xnor U6809 (N_6809,N_4621,N_5703);
or U6810 (N_6810,N_4754,N_4953);
nor U6811 (N_6811,N_5230,N_4904);
xor U6812 (N_6812,N_4807,N_5639);
nand U6813 (N_6813,N_5413,N_5338);
and U6814 (N_6814,N_5228,N_4554);
nand U6815 (N_6815,N_5411,N_4598);
or U6816 (N_6816,N_5869,N_4828);
nand U6817 (N_6817,N_5886,N_5550);
nor U6818 (N_6818,N_4899,N_5393);
nor U6819 (N_6819,N_4923,N_4500);
xnor U6820 (N_6820,N_4579,N_5368);
nor U6821 (N_6821,N_5030,N_5446);
or U6822 (N_6822,N_4795,N_4780);
xor U6823 (N_6823,N_5830,N_5307);
nor U6824 (N_6824,N_5231,N_4862);
or U6825 (N_6825,N_5106,N_5227);
xor U6826 (N_6826,N_5870,N_4672);
nor U6827 (N_6827,N_5752,N_5989);
nand U6828 (N_6828,N_5431,N_5160);
nand U6829 (N_6829,N_4870,N_4964);
nor U6830 (N_6830,N_5901,N_5017);
and U6831 (N_6831,N_5471,N_5000);
xor U6832 (N_6832,N_5237,N_5405);
nand U6833 (N_6833,N_5777,N_5501);
nand U6834 (N_6834,N_5390,N_4647);
xor U6835 (N_6835,N_4563,N_5397);
nor U6836 (N_6836,N_5746,N_5118);
nand U6837 (N_6837,N_5005,N_5741);
nor U6838 (N_6838,N_5164,N_5083);
xnor U6839 (N_6839,N_4729,N_4918);
nand U6840 (N_6840,N_4773,N_5675);
nor U6841 (N_6841,N_5874,N_5000);
or U6842 (N_6842,N_5330,N_4772);
and U6843 (N_6843,N_5166,N_4831);
nor U6844 (N_6844,N_5647,N_4847);
nand U6845 (N_6845,N_5590,N_5741);
and U6846 (N_6846,N_5701,N_4764);
xor U6847 (N_6847,N_4855,N_4622);
nor U6848 (N_6848,N_5106,N_4672);
and U6849 (N_6849,N_4533,N_5027);
and U6850 (N_6850,N_5328,N_5142);
nand U6851 (N_6851,N_5679,N_5222);
nand U6852 (N_6852,N_5358,N_5103);
or U6853 (N_6853,N_5399,N_5390);
xor U6854 (N_6854,N_5884,N_4827);
nor U6855 (N_6855,N_5844,N_5686);
and U6856 (N_6856,N_5171,N_4605);
nand U6857 (N_6857,N_5659,N_4971);
xnor U6858 (N_6858,N_4681,N_5844);
nand U6859 (N_6859,N_5216,N_5634);
nand U6860 (N_6860,N_5831,N_4689);
nor U6861 (N_6861,N_4751,N_5263);
or U6862 (N_6862,N_5807,N_5806);
and U6863 (N_6863,N_4656,N_5827);
and U6864 (N_6864,N_4775,N_4596);
xnor U6865 (N_6865,N_5438,N_5988);
and U6866 (N_6866,N_4948,N_4772);
and U6867 (N_6867,N_5755,N_5804);
nor U6868 (N_6868,N_4947,N_5569);
or U6869 (N_6869,N_4758,N_5997);
or U6870 (N_6870,N_5368,N_5240);
nand U6871 (N_6871,N_5803,N_5214);
xnor U6872 (N_6872,N_4723,N_4782);
xnor U6873 (N_6873,N_5458,N_4979);
and U6874 (N_6874,N_5361,N_5220);
nand U6875 (N_6875,N_5193,N_5723);
and U6876 (N_6876,N_5697,N_5185);
xnor U6877 (N_6877,N_5737,N_5467);
nor U6878 (N_6878,N_5270,N_5696);
nor U6879 (N_6879,N_5169,N_5191);
and U6880 (N_6880,N_4550,N_5991);
nor U6881 (N_6881,N_4556,N_4571);
nor U6882 (N_6882,N_4965,N_5398);
nand U6883 (N_6883,N_4810,N_5168);
nor U6884 (N_6884,N_5734,N_5182);
nor U6885 (N_6885,N_5199,N_4693);
nor U6886 (N_6886,N_4652,N_5967);
and U6887 (N_6887,N_4638,N_4985);
nand U6888 (N_6888,N_5620,N_4925);
xnor U6889 (N_6889,N_5433,N_5151);
and U6890 (N_6890,N_5803,N_5844);
or U6891 (N_6891,N_4532,N_5514);
xor U6892 (N_6892,N_4783,N_5473);
xnor U6893 (N_6893,N_4879,N_5052);
xor U6894 (N_6894,N_5911,N_4934);
and U6895 (N_6895,N_5016,N_5711);
or U6896 (N_6896,N_5451,N_4993);
or U6897 (N_6897,N_5311,N_5724);
and U6898 (N_6898,N_5252,N_5832);
or U6899 (N_6899,N_5281,N_4995);
nand U6900 (N_6900,N_4759,N_4593);
nor U6901 (N_6901,N_5406,N_5795);
nand U6902 (N_6902,N_5373,N_4575);
nand U6903 (N_6903,N_5996,N_4633);
or U6904 (N_6904,N_5187,N_5099);
nor U6905 (N_6905,N_5095,N_5565);
nor U6906 (N_6906,N_5108,N_5936);
nand U6907 (N_6907,N_4647,N_4826);
nand U6908 (N_6908,N_4747,N_5089);
xor U6909 (N_6909,N_5839,N_4763);
nand U6910 (N_6910,N_5620,N_5985);
nor U6911 (N_6911,N_5039,N_5866);
nor U6912 (N_6912,N_4872,N_5339);
and U6913 (N_6913,N_4913,N_4557);
nor U6914 (N_6914,N_5392,N_5826);
xnor U6915 (N_6915,N_5013,N_5125);
or U6916 (N_6916,N_5795,N_5235);
xor U6917 (N_6917,N_5451,N_5368);
xor U6918 (N_6918,N_4628,N_5592);
and U6919 (N_6919,N_4617,N_4969);
or U6920 (N_6920,N_4583,N_4855);
and U6921 (N_6921,N_4589,N_4692);
nor U6922 (N_6922,N_5184,N_5269);
and U6923 (N_6923,N_5469,N_5809);
nand U6924 (N_6924,N_5377,N_5060);
or U6925 (N_6925,N_4913,N_4812);
nand U6926 (N_6926,N_4528,N_5442);
xnor U6927 (N_6927,N_5021,N_5329);
nor U6928 (N_6928,N_5569,N_5557);
nand U6929 (N_6929,N_5202,N_5753);
and U6930 (N_6930,N_4625,N_4567);
nand U6931 (N_6931,N_5631,N_5805);
xor U6932 (N_6932,N_4842,N_5833);
nor U6933 (N_6933,N_5365,N_5701);
nand U6934 (N_6934,N_5636,N_5801);
and U6935 (N_6935,N_5112,N_5691);
nor U6936 (N_6936,N_5710,N_5502);
and U6937 (N_6937,N_5373,N_4996);
nand U6938 (N_6938,N_5789,N_5697);
xor U6939 (N_6939,N_5416,N_5037);
nand U6940 (N_6940,N_5835,N_4904);
or U6941 (N_6941,N_4817,N_5500);
nand U6942 (N_6942,N_5162,N_4560);
and U6943 (N_6943,N_4674,N_4844);
nor U6944 (N_6944,N_5449,N_5764);
nand U6945 (N_6945,N_4859,N_5925);
or U6946 (N_6946,N_5155,N_4827);
nand U6947 (N_6947,N_5764,N_5286);
and U6948 (N_6948,N_5122,N_5037);
or U6949 (N_6949,N_5351,N_5461);
nand U6950 (N_6950,N_5890,N_5625);
and U6951 (N_6951,N_5550,N_5820);
nor U6952 (N_6952,N_5097,N_5980);
or U6953 (N_6953,N_5446,N_4930);
and U6954 (N_6954,N_5050,N_5232);
and U6955 (N_6955,N_5109,N_5358);
nor U6956 (N_6956,N_5078,N_5054);
or U6957 (N_6957,N_4520,N_5046);
or U6958 (N_6958,N_5100,N_5909);
nand U6959 (N_6959,N_5264,N_5853);
nor U6960 (N_6960,N_5548,N_5943);
nor U6961 (N_6961,N_5957,N_5930);
nand U6962 (N_6962,N_4935,N_5477);
or U6963 (N_6963,N_5135,N_5981);
xor U6964 (N_6964,N_4815,N_5342);
nor U6965 (N_6965,N_5908,N_4529);
nand U6966 (N_6966,N_5032,N_4979);
nor U6967 (N_6967,N_5361,N_5810);
nand U6968 (N_6968,N_5505,N_5955);
xor U6969 (N_6969,N_5214,N_5067);
and U6970 (N_6970,N_5269,N_4918);
xor U6971 (N_6971,N_5561,N_5306);
and U6972 (N_6972,N_5034,N_5641);
xor U6973 (N_6973,N_5424,N_5029);
nand U6974 (N_6974,N_5482,N_5203);
xor U6975 (N_6975,N_5080,N_4954);
nand U6976 (N_6976,N_4629,N_5858);
or U6977 (N_6977,N_5425,N_4668);
or U6978 (N_6978,N_5976,N_5829);
nand U6979 (N_6979,N_5666,N_5711);
and U6980 (N_6980,N_5310,N_5261);
nand U6981 (N_6981,N_5931,N_5514);
nor U6982 (N_6982,N_4676,N_5173);
nor U6983 (N_6983,N_4729,N_5966);
xor U6984 (N_6984,N_5921,N_4758);
nand U6985 (N_6985,N_5704,N_5973);
nand U6986 (N_6986,N_4749,N_5799);
xor U6987 (N_6987,N_5001,N_4625);
nor U6988 (N_6988,N_5622,N_5580);
nand U6989 (N_6989,N_5694,N_5052);
and U6990 (N_6990,N_5512,N_5087);
nor U6991 (N_6991,N_4849,N_5848);
or U6992 (N_6992,N_5210,N_5299);
and U6993 (N_6993,N_5552,N_4583);
or U6994 (N_6994,N_5856,N_5421);
nand U6995 (N_6995,N_4630,N_4721);
or U6996 (N_6996,N_5090,N_5375);
nand U6997 (N_6997,N_5983,N_4828);
and U6998 (N_6998,N_4515,N_4715);
nand U6999 (N_6999,N_5414,N_4994);
and U7000 (N_7000,N_4651,N_5391);
nor U7001 (N_7001,N_5333,N_4738);
xnor U7002 (N_7002,N_5477,N_5683);
nand U7003 (N_7003,N_5551,N_5920);
nor U7004 (N_7004,N_5650,N_5126);
and U7005 (N_7005,N_5941,N_5062);
nand U7006 (N_7006,N_4816,N_4530);
xor U7007 (N_7007,N_5857,N_4624);
and U7008 (N_7008,N_5017,N_5604);
or U7009 (N_7009,N_4880,N_4562);
nand U7010 (N_7010,N_5669,N_5798);
xor U7011 (N_7011,N_5554,N_4674);
nand U7012 (N_7012,N_5443,N_4765);
or U7013 (N_7013,N_5581,N_5613);
nand U7014 (N_7014,N_5272,N_5369);
nor U7015 (N_7015,N_5812,N_4901);
and U7016 (N_7016,N_5259,N_5648);
xnor U7017 (N_7017,N_4712,N_4921);
and U7018 (N_7018,N_4942,N_5844);
and U7019 (N_7019,N_4521,N_5739);
xor U7020 (N_7020,N_5214,N_4540);
xnor U7021 (N_7021,N_5573,N_5877);
or U7022 (N_7022,N_4504,N_4934);
xor U7023 (N_7023,N_4769,N_5726);
nand U7024 (N_7024,N_5814,N_5706);
nand U7025 (N_7025,N_5311,N_4810);
nand U7026 (N_7026,N_5740,N_4915);
xor U7027 (N_7027,N_5856,N_5989);
nor U7028 (N_7028,N_4872,N_4847);
nor U7029 (N_7029,N_4901,N_5317);
or U7030 (N_7030,N_5577,N_5168);
or U7031 (N_7031,N_4990,N_5339);
or U7032 (N_7032,N_4837,N_5768);
or U7033 (N_7033,N_5985,N_4942);
nor U7034 (N_7034,N_4832,N_4773);
xor U7035 (N_7035,N_4504,N_4726);
nor U7036 (N_7036,N_4846,N_4931);
nand U7037 (N_7037,N_5822,N_4705);
or U7038 (N_7038,N_5280,N_4875);
xor U7039 (N_7039,N_4924,N_5406);
or U7040 (N_7040,N_5723,N_5181);
xor U7041 (N_7041,N_5205,N_5323);
and U7042 (N_7042,N_4801,N_4961);
or U7043 (N_7043,N_5537,N_4628);
and U7044 (N_7044,N_4795,N_5329);
and U7045 (N_7045,N_5961,N_5724);
xor U7046 (N_7046,N_5460,N_5837);
or U7047 (N_7047,N_5003,N_5759);
and U7048 (N_7048,N_5055,N_4581);
nand U7049 (N_7049,N_5105,N_5987);
or U7050 (N_7050,N_4696,N_4760);
xnor U7051 (N_7051,N_5453,N_5550);
and U7052 (N_7052,N_5644,N_5591);
nand U7053 (N_7053,N_5509,N_5219);
xnor U7054 (N_7054,N_5894,N_4552);
nor U7055 (N_7055,N_4949,N_5077);
xor U7056 (N_7056,N_5660,N_5384);
or U7057 (N_7057,N_4660,N_5372);
nand U7058 (N_7058,N_5786,N_4631);
or U7059 (N_7059,N_5677,N_5872);
xor U7060 (N_7060,N_5616,N_4662);
or U7061 (N_7061,N_5831,N_5903);
nand U7062 (N_7062,N_4796,N_5113);
or U7063 (N_7063,N_5981,N_4859);
xor U7064 (N_7064,N_4673,N_5166);
xor U7065 (N_7065,N_5780,N_5236);
or U7066 (N_7066,N_5764,N_5371);
nor U7067 (N_7067,N_4753,N_4878);
nor U7068 (N_7068,N_5058,N_4924);
nand U7069 (N_7069,N_4894,N_4688);
nand U7070 (N_7070,N_4546,N_5082);
xor U7071 (N_7071,N_5118,N_4509);
nor U7072 (N_7072,N_4997,N_4573);
and U7073 (N_7073,N_5707,N_4720);
xor U7074 (N_7074,N_4677,N_5103);
or U7075 (N_7075,N_5182,N_5349);
or U7076 (N_7076,N_5073,N_5895);
xnor U7077 (N_7077,N_4535,N_5673);
nand U7078 (N_7078,N_5697,N_4900);
xor U7079 (N_7079,N_5565,N_5849);
or U7080 (N_7080,N_5984,N_5111);
nand U7081 (N_7081,N_5784,N_5229);
or U7082 (N_7082,N_5236,N_4665);
nor U7083 (N_7083,N_5295,N_5017);
nand U7084 (N_7084,N_5757,N_5944);
and U7085 (N_7085,N_5981,N_5113);
nand U7086 (N_7086,N_5387,N_5175);
nand U7087 (N_7087,N_5391,N_5814);
xor U7088 (N_7088,N_5873,N_5673);
xor U7089 (N_7089,N_4702,N_5609);
xnor U7090 (N_7090,N_5956,N_5432);
and U7091 (N_7091,N_5468,N_4718);
nor U7092 (N_7092,N_4657,N_5144);
or U7093 (N_7093,N_5512,N_5388);
nand U7094 (N_7094,N_5742,N_4963);
and U7095 (N_7095,N_5662,N_5595);
xnor U7096 (N_7096,N_5122,N_4869);
and U7097 (N_7097,N_5058,N_4754);
nand U7098 (N_7098,N_5835,N_4595);
xor U7099 (N_7099,N_5356,N_4793);
nand U7100 (N_7100,N_5289,N_5164);
nor U7101 (N_7101,N_4576,N_4717);
xor U7102 (N_7102,N_5206,N_5132);
or U7103 (N_7103,N_5055,N_5748);
or U7104 (N_7104,N_5696,N_4675);
and U7105 (N_7105,N_5803,N_5392);
or U7106 (N_7106,N_4903,N_5536);
nand U7107 (N_7107,N_5505,N_5921);
nand U7108 (N_7108,N_5039,N_4843);
and U7109 (N_7109,N_5001,N_4586);
xor U7110 (N_7110,N_5774,N_4938);
and U7111 (N_7111,N_5022,N_4835);
nor U7112 (N_7112,N_5437,N_5874);
xor U7113 (N_7113,N_4644,N_5505);
xor U7114 (N_7114,N_4951,N_5115);
xor U7115 (N_7115,N_5728,N_5813);
or U7116 (N_7116,N_5510,N_5018);
nand U7117 (N_7117,N_5468,N_5198);
nand U7118 (N_7118,N_5894,N_4874);
and U7119 (N_7119,N_4667,N_5974);
or U7120 (N_7120,N_5948,N_4782);
xnor U7121 (N_7121,N_5504,N_4787);
nor U7122 (N_7122,N_4549,N_5187);
nor U7123 (N_7123,N_4685,N_5147);
xnor U7124 (N_7124,N_5070,N_5699);
or U7125 (N_7125,N_5905,N_5177);
nand U7126 (N_7126,N_5003,N_5155);
or U7127 (N_7127,N_5674,N_5527);
xnor U7128 (N_7128,N_5058,N_5988);
or U7129 (N_7129,N_5897,N_5643);
nor U7130 (N_7130,N_5966,N_5872);
nor U7131 (N_7131,N_5051,N_5391);
or U7132 (N_7132,N_5132,N_4706);
nor U7133 (N_7133,N_4655,N_5834);
and U7134 (N_7134,N_5540,N_5049);
nor U7135 (N_7135,N_5563,N_5320);
nand U7136 (N_7136,N_5267,N_4545);
nor U7137 (N_7137,N_4617,N_4794);
or U7138 (N_7138,N_4786,N_4711);
nor U7139 (N_7139,N_5401,N_5371);
and U7140 (N_7140,N_5724,N_5682);
nand U7141 (N_7141,N_5995,N_5357);
or U7142 (N_7142,N_4554,N_4914);
nor U7143 (N_7143,N_5922,N_5338);
and U7144 (N_7144,N_5520,N_4661);
or U7145 (N_7145,N_4877,N_5673);
nor U7146 (N_7146,N_5824,N_4727);
and U7147 (N_7147,N_4945,N_4691);
and U7148 (N_7148,N_5052,N_5808);
nor U7149 (N_7149,N_5810,N_4779);
nor U7150 (N_7150,N_5521,N_5480);
and U7151 (N_7151,N_5357,N_5801);
xnor U7152 (N_7152,N_4967,N_4939);
or U7153 (N_7153,N_4967,N_5114);
or U7154 (N_7154,N_5160,N_5569);
nor U7155 (N_7155,N_5073,N_4814);
xnor U7156 (N_7156,N_4553,N_5536);
nand U7157 (N_7157,N_4625,N_4860);
and U7158 (N_7158,N_5271,N_4988);
or U7159 (N_7159,N_5984,N_4655);
or U7160 (N_7160,N_5983,N_4763);
nor U7161 (N_7161,N_5938,N_5243);
nand U7162 (N_7162,N_4794,N_4808);
and U7163 (N_7163,N_4894,N_4546);
or U7164 (N_7164,N_5232,N_5228);
nand U7165 (N_7165,N_4811,N_5852);
and U7166 (N_7166,N_5973,N_5205);
xnor U7167 (N_7167,N_4714,N_4855);
nor U7168 (N_7168,N_4503,N_5653);
xor U7169 (N_7169,N_5883,N_5300);
and U7170 (N_7170,N_5495,N_5069);
xor U7171 (N_7171,N_5045,N_4623);
or U7172 (N_7172,N_5269,N_5505);
and U7173 (N_7173,N_4809,N_4895);
xnor U7174 (N_7174,N_5444,N_4884);
nor U7175 (N_7175,N_5302,N_5715);
nor U7176 (N_7176,N_4502,N_5594);
nand U7177 (N_7177,N_5430,N_4900);
nor U7178 (N_7178,N_5216,N_4610);
nand U7179 (N_7179,N_5252,N_5042);
or U7180 (N_7180,N_5705,N_4557);
and U7181 (N_7181,N_5015,N_5300);
nand U7182 (N_7182,N_5500,N_5863);
nor U7183 (N_7183,N_5673,N_4641);
xor U7184 (N_7184,N_5501,N_5349);
nor U7185 (N_7185,N_5155,N_5829);
xnor U7186 (N_7186,N_5385,N_5243);
xor U7187 (N_7187,N_5684,N_4791);
nand U7188 (N_7188,N_5076,N_5893);
nor U7189 (N_7189,N_4739,N_5461);
or U7190 (N_7190,N_5589,N_4923);
or U7191 (N_7191,N_5314,N_4624);
or U7192 (N_7192,N_5736,N_5605);
nand U7193 (N_7193,N_5124,N_5291);
xor U7194 (N_7194,N_5903,N_5791);
or U7195 (N_7195,N_5849,N_5834);
nor U7196 (N_7196,N_4527,N_5102);
nor U7197 (N_7197,N_4511,N_5993);
xor U7198 (N_7198,N_4773,N_4585);
nand U7199 (N_7199,N_5546,N_5311);
xnor U7200 (N_7200,N_5266,N_5879);
xor U7201 (N_7201,N_5710,N_5379);
nand U7202 (N_7202,N_5727,N_4914);
nor U7203 (N_7203,N_5357,N_5244);
and U7204 (N_7204,N_5045,N_5688);
xnor U7205 (N_7205,N_4842,N_5252);
xnor U7206 (N_7206,N_4632,N_4977);
nand U7207 (N_7207,N_5095,N_5163);
nand U7208 (N_7208,N_4603,N_5454);
nor U7209 (N_7209,N_5586,N_5231);
nor U7210 (N_7210,N_5049,N_5885);
or U7211 (N_7211,N_4623,N_4919);
xnor U7212 (N_7212,N_4839,N_5789);
xor U7213 (N_7213,N_4749,N_5159);
nor U7214 (N_7214,N_4645,N_4618);
nor U7215 (N_7215,N_5547,N_5744);
and U7216 (N_7216,N_5635,N_5009);
or U7217 (N_7217,N_5606,N_5366);
nor U7218 (N_7218,N_5120,N_5051);
nand U7219 (N_7219,N_4572,N_4904);
xnor U7220 (N_7220,N_4641,N_5506);
xnor U7221 (N_7221,N_5884,N_4578);
or U7222 (N_7222,N_5721,N_5294);
xor U7223 (N_7223,N_5572,N_4947);
xor U7224 (N_7224,N_5568,N_4650);
xor U7225 (N_7225,N_5711,N_4543);
nor U7226 (N_7226,N_5252,N_5698);
or U7227 (N_7227,N_5083,N_5322);
xor U7228 (N_7228,N_5077,N_5188);
nor U7229 (N_7229,N_5297,N_5244);
nand U7230 (N_7230,N_4915,N_5128);
xor U7231 (N_7231,N_5499,N_5239);
nand U7232 (N_7232,N_5143,N_5927);
or U7233 (N_7233,N_5325,N_5009);
nand U7234 (N_7234,N_5126,N_4854);
nor U7235 (N_7235,N_5427,N_4790);
or U7236 (N_7236,N_5704,N_5897);
or U7237 (N_7237,N_4978,N_4752);
or U7238 (N_7238,N_4500,N_4934);
or U7239 (N_7239,N_4855,N_4736);
nor U7240 (N_7240,N_4693,N_4737);
nor U7241 (N_7241,N_4845,N_4668);
nand U7242 (N_7242,N_5497,N_4730);
or U7243 (N_7243,N_4536,N_4535);
or U7244 (N_7244,N_5788,N_5777);
nor U7245 (N_7245,N_4962,N_5163);
or U7246 (N_7246,N_5830,N_5464);
or U7247 (N_7247,N_5843,N_4756);
or U7248 (N_7248,N_4828,N_5571);
and U7249 (N_7249,N_5367,N_5795);
nand U7250 (N_7250,N_5467,N_5049);
or U7251 (N_7251,N_5024,N_5161);
nor U7252 (N_7252,N_5257,N_5420);
nand U7253 (N_7253,N_5916,N_5734);
and U7254 (N_7254,N_5468,N_5870);
or U7255 (N_7255,N_4699,N_4622);
nor U7256 (N_7256,N_4598,N_4613);
and U7257 (N_7257,N_5799,N_4614);
xor U7258 (N_7258,N_4596,N_5627);
nand U7259 (N_7259,N_5860,N_5996);
nor U7260 (N_7260,N_5781,N_4673);
nor U7261 (N_7261,N_4672,N_5919);
and U7262 (N_7262,N_5666,N_4905);
and U7263 (N_7263,N_4930,N_5973);
nor U7264 (N_7264,N_4831,N_4623);
xor U7265 (N_7265,N_5915,N_5542);
and U7266 (N_7266,N_5692,N_5326);
or U7267 (N_7267,N_5625,N_5035);
nor U7268 (N_7268,N_5367,N_5479);
and U7269 (N_7269,N_4672,N_5750);
or U7270 (N_7270,N_4809,N_5617);
nand U7271 (N_7271,N_4567,N_5746);
nand U7272 (N_7272,N_5792,N_5363);
nand U7273 (N_7273,N_5077,N_5294);
or U7274 (N_7274,N_5092,N_4862);
and U7275 (N_7275,N_4977,N_5410);
or U7276 (N_7276,N_5518,N_5668);
and U7277 (N_7277,N_5844,N_5264);
and U7278 (N_7278,N_5396,N_4776);
nand U7279 (N_7279,N_4679,N_5503);
and U7280 (N_7280,N_5928,N_5180);
nand U7281 (N_7281,N_5021,N_5449);
nand U7282 (N_7282,N_5464,N_5616);
nor U7283 (N_7283,N_5038,N_5845);
xor U7284 (N_7284,N_4866,N_5954);
nand U7285 (N_7285,N_5741,N_5115);
nor U7286 (N_7286,N_5275,N_5723);
xnor U7287 (N_7287,N_5896,N_4841);
xnor U7288 (N_7288,N_5295,N_5855);
xor U7289 (N_7289,N_5793,N_4993);
nor U7290 (N_7290,N_4546,N_5178);
nor U7291 (N_7291,N_5410,N_5494);
nand U7292 (N_7292,N_5713,N_5095);
or U7293 (N_7293,N_5838,N_4875);
and U7294 (N_7294,N_5832,N_5673);
xnor U7295 (N_7295,N_5380,N_5404);
and U7296 (N_7296,N_5814,N_4521);
xnor U7297 (N_7297,N_4933,N_5936);
xnor U7298 (N_7298,N_5067,N_5052);
or U7299 (N_7299,N_5874,N_4544);
or U7300 (N_7300,N_5744,N_4600);
xnor U7301 (N_7301,N_4947,N_5294);
nand U7302 (N_7302,N_4577,N_5190);
nor U7303 (N_7303,N_4998,N_5834);
xnor U7304 (N_7304,N_5307,N_4600);
nand U7305 (N_7305,N_5598,N_5100);
and U7306 (N_7306,N_5935,N_4687);
or U7307 (N_7307,N_4666,N_4705);
xnor U7308 (N_7308,N_5163,N_5382);
xnor U7309 (N_7309,N_5129,N_5729);
nand U7310 (N_7310,N_4898,N_5785);
and U7311 (N_7311,N_5317,N_5892);
nand U7312 (N_7312,N_5065,N_4570);
nand U7313 (N_7313,N_5380,N_5034);
nor U7314 (N_7314,N_4798,N_5849);
or U7315 (N_7315,N_5069,N_4807);
nor U7316 (N_7316,N_4768,N_5471);
nor U7317 (N_7317,N_4791,N_4977);
nor U7318 (N_7318,N_5719,N_5410);
xnor U7319 (N_7319,N_5020,N_5500);
nand U7320 (N_7320,N_5033,N_4811);
xnor U7321 (N_7321,N_4885,N_4830);
nand U7322 (N_7322,N_5129,N_4507);
nand U7323 (N_7323,N_5374,N_4689);
and U7324 (N_7324,N_5667,N_5263);
nand U7325 (N_7325,N_4691,N_5049);
xnor U7326 (N_7326,N_4947,N_5807);
and U7327 (N_7327,N_5104,N_4669);
or U7328 (N_7328,N_5561,N_5702);
xor U7329 (N_7329,N_5483,N_5923);
or U7330 (N_7330,N_5572,N_5745);
xor U7331 (N_7331,N_4521,N_5036);
or U7332 (N_7332,N_4946,N_4752);
xor U7333 (N_7333,N_4544,N_5438);
xnor U7334 (N_7334,N_5461,N_5590);
and U7335 (N_7335,N_5476,N_5876);
and U7336 (N_7336,N_5579,N_5569);
nor U7337 (N_7337,N_5123,N_5396);
xnor U7338 (N_7338,N_5763,N_4603);
xnor U7339 (N_7339,N_5614,N_5604);
xor U7340 (N_7340,N_4677,N_4669);
or U7341 (N_7341,N_4662,N_4581);
or U7342 (N_7342,N_5391,N_5498);
or U7343 (N_7343,N_5856,N_4594);
nor U7344 (N_7344,N_4854,N_5774);
nand U7345 (N_7345,N_5032,N_4708);
xor U7346 (N_7346,N_5093,N_4514);
xnor U7347 (N_7347,N_5089,N_4744);
nor U7348 (N_7348,N_4507,N_5255);
xnor U7349 (N_7349,N_5988,N_5654);
or U7350 (N_7350,N_4537,N_5908);
nand U7351 (N_7351,N_5596,N_4754);
nor U7352 (N_7352,N_5589,N_4669);
xnor U7353 (N_7353,N_5576,N_5846);
nand U7354 (N_7354,N_5046,N_5725);
and U7355 (N_7355,N_5346,N_5609);
nor U7356 (N_7356,N_4886,N_5543);
xnor U7357 (N_7357,N_4851,N_5499);
xnor U7358 (N_7358,N_5844,N_5690);
nand U7359 (N_7359,N_5372,N_4599);
nand U7360 (N_7360,N_4521,N_5642);
xor U7361 (N_7361,N_4993,N_5079);
nand U7362 (N_7362,N_4807,N_4689);
xnor U7363 (N_7363,N_4807,N_5617);
or U7364 (N_7364,N_5286,N_5360);
nor U7365 (N_7365,N_5938,N_4679);
and U7366 (N_7366,N_5966,N_5953);
and U7367 (N_7367,N_4529,N_5161);
or U7368 (N_7368,N_5006,N_4642);
nand U7369 (N_7369,N_5066,N_4896);
nor U7370 (N_7370,N_5345,N_5343);
nor U7371 (N_7371,N_4506,N_4989);
or U7372 (N_7372,N_5565,N_5848);
nand U7373 (N_7373,N_4645,N_4891);
nor U7374 (N_7374,N_5703,N_4846);
xor U7375 (N_7375,N_4636,N_5951);
xor U7376 (N_7376,N_4949,N_4620);
nor U7377 (N_7377,N_5709,N_4876);
nand U7378 (N_7378,N_5817,N_4871);
and U7379 (N_7379,N_5651,N_5266);
nand U7380 (N_7380,N_5783,N_5880);
or U7381 (N_7381,N_5222,N_4861);
nor U7382 (N_7382,N_5905,N_5965);
or U7383 (N_7383,N_4754,N_5874);
nand U7384 (N_7384,N_5166,N_5314);
nand U7385 (N_7385,N_4955,N_4957);
or U7386 (N_7386,N_5947,N_4945);
or U7387 (N_7387,N_4823,N_5274);
and U7388 (N_7388,N_5876,N_4548);
and U7389 (N_7389,N_5275,N_4587);
and U7390 (N_7390,N_4539,N_5388);
and U7391 (N_7391,N_5159,N_4633);
or U7392 (N_7392,N_5073,N_5448);
nor U7393 (N_7393,N_5818,N_4594);
nor U7394 (N_7394,N_5641,N_5011);
nand U7395 (N_7395,N_5045,N_4929);
xnor U7396 (N_7396,N_5180,N_4938);
or U7397 (N_7397,N_5419,N_5794);
nor U7398 (N_7398,N_4638,N_4577);
and U7399 (N_7399,N_4795,N_4952);
or U7400 (N_7400,N_5595,N_5651);
xnor U7401 (N_7401,N_5061,N_5906);
nand U7402 (N_7402,N_5937,N_4849);
and U7403 (N_7403,N_4994,N_4985);
or U7404 (N_7404,N_5109,N_4677);
and U7405 (N_7405,N_5888,N_4806);
nor U7406 (N_7406,N_5474,N_5048);
nand U7407 (N_7407,N_5642,N_4703);
or U7408 (N_7408,N_4777,N_5404);
nor U7409 (N_7409,N_5170,N_5905);
and U7410 (N_7410,N_5439,N_5271);
nor U7411 (N_7411,N_4910,N_5523);
nand U7412 (N_7412,N_5462,N_4632);
and U7413 (N_7413,N_4836,N_4712);
or U7414 (N_7414,N_4852,N_5790);
and U7415 (N_7415,N_5419,N_5154);
nand U7416 (N_7416,N_5739,N_4800);
nand U7417 (N_7417,N_5809,N_5510);
or U7418 (N_7418,N_5469,N_4897);
xnor U7419 (N_7419,N_5507,N_4577);
and U7420 (N_7420,N_5098,N_4629);
xor U7421 (N_7421,N_5965,N_5985);
nor U7422 (N_7422,N_4567,N_5814);
nand U7423 (N_7423,N_5359,N_5247);
xnor U7424 (N_7424,N_4926,N_5085);
nor U7425 (N_7425,N_4631,N_5608);
or U7426 (N_7426,N_5082,N_5390);
and U7427 (N_7427,N_5796,N_5986);
or U7428 (N_7428,N_5682,N_5271);
nor U7429 (N_7429,N_5540,N_5289);
nand U7430 (N_7430,N_5346,N_5593);
nor U7431 (N_7431,N_4574,N_5473);
and U7432 (N_7432,N_5234,N_4674);
nor U7433 (N_7433,N_5587,N_4800);
or U7434 (N_7434,N_4525,N_4795);
nand U7435 (N_7435,N_5828,N_5485);
nor U7436 (N_7436,N_5775,N_5909);
nor U7437 (N_7437,N_4714,N_5774);
xnor U7438 (N_7438,N_4897,N_5297);
nor U7439 (N_7439,N_5650,N_5017);
or U7440 (N_7440,N_5884,N_5815);
xor U7441 (N_7441,N_5494,N_5288);
nor U7442 (N_7442,N_5849,N_4862);
xor U7443 (N_7443,N_5959,N_4515);
xnor U7444 (N_7444,N_5861,N_4863);
or U7445 (N_7445,N_5228,N_5610);
nor U7446 (N_7446,N_5366,N_5992);
nor U7447 (N_7447,N_5681,N_4505);
or U7448 (N_7448,N_5738,N_5788);
and U7449 (N_7449,N_4549,N_4760);
xnor U7450 (N_7450,N_5591,N_5336);
nand U7451 (N_7451,N_4876,N_5553);
and U7452 (N_7452,N_4518,N_4530);
or U7453 (N_7453,N_5727,N_5180);
nor U7454 (N_7454,N_5660,N_5196);
nor U7455 (N_7455,N_5067,N_5053);
nand U7456 (N_7456,N_5326,N_4846);
nor U7457 (N_7457,N_5895,N_4712);
nor U7458 (N_7458,N_5670,N_5048);
or U7459 (N_7459,N_5992,N_5973);
xor U7460 (N_7460,N_4621,N_5296);
or U7461 (N_7461,N_5027,N_4785);
nor U7462 (N_7462,N_5432,N_4659);
and U7463 (N_7463,N_4980,N_5248);
and U7464 (N_7464,N_5023,N_5322);
nand U7465 (N_7465,N_5139,N_5364);
nand U7466 (N_7466,N_4741,N_4707);
nand U7467 (N_7467,N_4817,N_5511);
nand U7468 (N_7468,N_5074,N_5328);
nor U7469 (N_7469,N_5704,N_4526);
xor U7470 (N_7470,N_5832,N_4668);
or U7471 (N_7471,N_5660,N_4737);
nor U7472 (N_7472,N_4695,N_5353);
nor U7473 (N_7473,N_4523,N_5337);
and U7474 (N_7474,N_5735,N_5488);
xnor U7475 (N_7475,N_4999,N_5930);
nor U7476 (N_7476,N_5627,N_5830);
nor U7477 (N_7477,N_4637,N_5153);
and U7478 (N_7478,N_5715,N_5515);
nand U7479 (N_7479,N_4756,N_5086);
xor U7480 (N_7480,N_5531,N_5455);
nand U7481 (N_7481,N_5312,N_5969);
or U7482 (N_7482,N_4897,N_5614);
nor U7483 (N_7483,N_5115,N_5791);
nor U7484 (N_7484,N_5265,N_4747);
or U7485 (N_7485,N_5464,N_4682);
nor U7486 (N_7486,N_4849,N_5742);
or U7487 (N_7487,N_5140,N_5023);
xor U7488 (N_7488,N_5529,N_5287);
and U7489 (N_7489,N_5222,N_4986);
or U7490 (N_7490,N_5999,N_5611);
and U7491 (N_7491,N_5319,N_5317);
xor U7492 (N_7492,N_4986,N_4938);
or U7493 (N_7493,N_5354,N_4540);
or U7494 (N_7494,N_5324,N_5218);
xnor U7495 (N_7495,N_4894,N_4919);
nor U7496 (N_7496,N_4510,N_5501);
nand U7497 (N_7497,N_4735,N_5984);
xor U7498 (N_7498,N_5005,N_5699);
and U7499 (N_7499,N_4592,N_5329);
or U7500 (N_7500,N_6314,N_6462);
and U7501 (N_7501,N_6699,N_6642);
nor U7502 (N_7502,N_7004,N_7001);
or U7503 (N_7503,N_6159,N_6329);
nor U7504 (N_7504,N_7209,N_6971);
nand U7505 (N_7505,N_6029,N_6361);
nor U7506 (N_7506,N_7311,N_6498);
or U7507 (N_7507,N_6485,N_6725);
and U7508 (N_7508,N_7218,N_6575);
nor U7509 (N_7509,N_6786,N_6011);
and U7510 (N_7510,N_6936,N_7281);
nor U7511 (N_7511,N_6331,N_6750);
xnor U7512 (N_7512,N_6760,N_6705);
xor U7513 (N_7513,N_6647,N_6256);
nor U7514 (N_7514,N_6567,N_6694);
and U7515 (N_7515,N_6319,N_6248);
and U7516 (N_7516,N_7419,N_6906);
nor U7517 (N_7517,N_6904,N_6215);
xor U7518 (N_7518,N_6925,N_6003);
nor U7519 (N_7519,N_6438,N_7245);
xnor U7520 (N_7520,N_6338,N_7081);
nand U7521 (N_7521,N_7136,N_7280);
or U7522 (N_7522,N_7264,N_7201);
and U7523 (N_7523,N_6006,N_6747);
nand U7524 (N_7524,N_6278,N_7456);
nand U7525 (N_7525,N_7086,N_7040);
nand U7526 (N_7526,N_6288,N_6665);
and U7527 (N_7527,N_7338,N_6561);
xor U7528 (N_7528,N_6882,N_6210);
or U7529 (N_7529,N_6590,N_6229);
and U7530 (N_7530,N_7015,N_6231);
and U7531 (N_7531,N_6174,N_6086);
nor U7532 (N_7532,N_6082,N_6764);
nand U7533 (N_7533,N_7157,N_7309);
nor U7534 (N_7534,N_6578,N_6626);
and U7535 (N_7535,N_6352,N_7296);
and U7536 (N_7536,N_7232,N_6163);
and U7537 (N_7537,N_7066,N_6240);
nand U7538 (N_7538,N_6509,N_7165);
nor U7539 (N_7539,N_6475,N_7110);
or U7540 (N_7540,N_6744,N_7315);
xor U7541 (N_7541,N_7133,N_6680);
nor U7542 (N_7542,N_6600,N_6966);
or U7543 (N_7543,N_6834,N_7016);
or U7544 (N_7544,N_7047,N_6991);
or U7545 (N_7545,N_6650,N_7484);
and U7546 (N_7546,N_7400,N_6242);
and U7547 (N_7547,N_6563,N_6099);
or U7548 (N_7548,N_6782,N_6207);
or U7549 (N_7549,N_7424,N_6377);
and U7550 (N_7550,N_6459,N_6281);
nor U7551 (N_7551,N_6609,N_6209);
xor U7552 (N_7552,N_7073,N_6374);
nand U7553 (N_7553,N_6681,N_7046);
and U7554 (N_7554,N_7444,N_6506);
nor U7555 (N_7555,N_6817,N_6870);
nand U7556 (N_7556,N_6812,N_6565);
xnor U7557 (N_7557,N_7101,N_7342);
xnor U7558 (N_7558,N_6426,N_7149);
nand U7559 (N_7559,N_6917,N_6039);
xor U7560 (N_7560,N_6689,N_6214);
nor U7561 (N_7561,N_6739,N_7297);
xnor U7562 (N_7562,N_7359,N_6171);
xor U7563 (N_7563,N_6830,N_6101);
nand U7564 (N_7564,N_6604,N_6837);
nor U7565 (N_7565,N_7399,N_6063);
nor U7566 (N_7566,N_7117,N_6525);
or U7567 (N_7567,N_6037,N_6810);
or U7568 (N_7568,N_6083,N_7222);
and U7569 (N_7569,N_6342,N_6829);
nand U7570 (N_7570,N_6613,N_7446);
nand U7571 (N_7571,N_6058,N_6606);
nand U7572 (N_7572,N_6838,N_7403);
nor U7573 (N_7573,N_6419,N_6191);
nor U7574 (N_7574,N_7486,N_6913);
and U7575 (N_7575,N_6467,N_7119);
and U7576 (N_7576,N_7471,N_6129);
nor U7577 (N_7577,N_6218,N_6683);
and U7578 (N_7578,N_6146,N_6894);
and U7579 (N_7579,N_7491,N_6045);
nand U7580 (N_7580,N_7352,N_6597);
and U7581 (N_7581,N_7289,N_7158);
and U7582 (N_7582,N_6335,N_7294);
and U7583 (N_7583,N_6857,N_6616);
and U7584 (N_7584,N_7048,N_6263);
or U7585 (N_7585,N_7061,N_6056);
nand U7586 (N_7586,N_6260,N_6555);
or U7587 (N_7587,N_7435,N_7454);
xnor U7588 (N_7588,N_6236,N_6763);
nand U7589 (N_7589,N_6127,N_7227);
nor U7590 (N_7590,N_6283,N_6005);
and U7591 (N_7591,N_7021,N_6435);
or U7592 (N_7592,N_6295,N_6748);
and U7593 (N_7593,N_6398,N_7215);
xor U7594 (N_7594,N_6638,N_6022);
or U7595 (N_7595,N_6270,N_7335);
or U7596 (N_7596,N_6866,N_6441);
nor U7597 (N_7597,N_6357,N_6570);
or U7598 (N_7598,N_6098,N_7205);
and U7599 (N_7599,N_6652,N_6144);
xnor U7600 (N_7600,N_7022,N_6967);
nand U7601 (N_7601,N_6976,N_6093);
nand U7602 (N_7602,N_6534,N_6385);
xnor U7603 (N_7603,N_7060,N_7429);
xor U7604 (N_7604,N_6696,N_6275);
xnor U7605 (N_7605,N_6131,N_6300);
or U7606 (N_7606,N_6784,N_6585);
nor U7607 (N_7607,N_6334,N_7235);
or U7608 (N_7608,N_6852,N_7287);
nor U7609 (N_7609,N_6995,N_6420);
or U7610 (N_7610,N_6389,N_6228);
nand U7611 (N_7611,N_7090,N_6767);
and U7612 (N_7612,N_7260,N_6495);
nand U7613 (N_7613,N_6137,N_6019);
and U7614 (N_7614,N_6494,N_7188);
and U7615 (N_7615,N_6775,N_6051);
and U7616 (N_7616,N_6250,N_6823);
or U7617 (N_7617,N_6956,N_6518);
nor U7618 (N_7618,N_6010,N_6623);
or U7619 (N_7619,N_6414,N_6199);
or U7620 (N_7620,N_6094,N_6486);
nand U7621 (N_7621,N_7416,N_7452);
xor U7622 (N_7622,N_7139,N_6713);
xnor U7623 (N_7623,N_6688,N_6977);
xor U7624 (N_7624,N_6589,N_6772);
or U7625 (N_7625,N_6035,N_6999);
nand U7626 (N_7626,N_6566,N_6150);
nand U7627 (N_7627,N_6751,N_6611);
nor U7628 (N_7628,N_6679,N_7255);
or U7629 (N_7629,N_6203,N_6911);
nand U7630 (N_7630,N_6643,N_6235);
and U7631 (N_7631,N_6928,N_6660);
nor U7632 (N_7632,N_6571,N_7483);
or U7633 (N_7633,N_6164,N_7380);
and U7634 (N_7634,N_6880,N_7387);
nor U7635 (N_7635,N_7316,N_7396);
and U7636 (N_7636,N_7208,N_6173);
or U7637 (N_7637,N_6392,N_7310);
xnor U7638 (N_7638,N_6266,N_7358);
xnor U7639 (N_7639,N_6141,N_6187);
nand U7640 (N_7640,N_7293,N_6104);
and U7641 (N_7641,N_6631,N_6493);
xor U7642 (N_7642,N_6644,N_7192);
and U7643 (N_7643,N_6265,N_7497);
nand U7644 (N_7644,N_6864,N_6992);
or U7645 (N_7645,N_6983,N_6395);
nor U7646 (N_7646,N_6794,N_6701);
or U7647 (N_7647,N_6607,N_6793);
and U7648 (N_7648,N_6412,N_6196);
and U7649 (N_7649,N_6769,N_6773);
xor U7650 (N_7650,N_7198,N_6023);
nor U7651 (N_7651,N_6602,N_6997);
and U7652 (N_7652,N_6289,N_7443);
nor U7653 (N_7653,N_6456,N_6798);
and U7654 (N_7654,N_6076,N_7002);
or U7655 (N_7655,N_7050,N_6321);
nor U7656 (N_7656,N_6861,N_6349);
nand U7657 (N_7657,N_7327,N_6080);
nand U7658 (N_7658,N_7499,N_7204);
or U7659 (N_7659,N_6253,N_6247);
nand U7660 (N_7660,N_6788,N_7112);
nor U7661 (N_7661,N_6167,N_7391);
nor U7662 (N_7662,N_6869,N_6111);
and U7663 (N_7663,N_6517,N_7160);
and U7664 (N_7664,N_7250,N_7346);
xnor U7665 (N_7665,N_7434,N_6519);
nand U7666 (N_7666,N_7091,N_6286);
nor U7667 (N_7667,N_7175,N_6312);
xnor U7668 (N_7668,N_7372,N_6016);
and U7669 (N_7669,N_7489,N_6282);
nor U7670 (N_7670,N_6536,N_7465);
and U7671 (N_7671,N_7357,N_6139);
and U7672 (N_7672,N_6117,N_7064);
xnor U7673 (N_7673,N_6478,N_6133);
and U7674 (N_7674,N_7267,N_6376);
nor U7675 (N_7675,N_6386,N_6640);
and U7676 (N_7676,N_6558,N_6854);
or U7677 (N_7677,N_7003,N_6630);
or U7678 (N_7678,N_6937,N_6178);
xor U7679 (N_7679,N_6007,N_7492);
and U7680 (N_7680,N_7174,N_7355);
and U7681 (N_7681,N_7082,N_6716);
or U7682 (N_7682,N_6900,N_6136);
nand U7683 (N_7683,N_6635,N_7168);
nand U7684 (N_7684,N_7238,N_6065);
nor U7685 (N_7685,N_7448,N_6390);
nand U7686 (N_7686,N_7284,N_6557);
and U7687 (N_7687,N_6388,N_6934);
xor U7688 (N_7688,N_6732,N_6401);
and U7689 (N_7689,N_6340,N_7071);
nand U7690 (N_7690,N_6789,N_7373);
nor U7691 (N_7691,N_6531,N_7303);
nand U7692 (N_7692,N_6828,N_6027);
and U7693 (N_7693,N_6610,N_6918);
xnor U7694 (N_7694,N_7286,N_6128);
xnor U7695 (N_7695,N_7412,N_6706);
nor U7696 (N_7696,N_7195,N_7045);
xnor U7697 (N_7697,N_7487,N_7422);
and U7698 (N_7698,N_6726,N_6134);
xor U7699 (N_7699,N_6985,N_7244);
and U7700 (N_7700,N_6439,N_7010);
xor U7701 (N_7701,N_6048,N_7383);
nor U7702 (N_7702,N_6826,N_6119);
and U7703 (N_7703,N_7051,N_6803);
and U7704 (N_7704,N_6427,N_6077);
and U7705 (N_7705,N_6227,N_7056);
nor U7706 (N_7706,N_6473,N_7037);
nor U7707 (N_7707,N_6158,N_6107);
nand U7708 (N_7708,N_6960,N_7441);
nor U7709 (N_7709,N_6415,N_6755);
nand U7710 (N_7710,N_6059,N_7231);
xnor U7711 (N_7711,N_7087,N_6238);
xnor U7712 (N_7712,N_6592,N_6050);
nand U7713 (N_7713,N_7191,N_7254);
nor U7714 (N_7714,N_6587,N_7299);
xnor U7715 (N_7715,N_6115,N_6064);
nand U7716 (N_7716,N_6806,N_6280);
or U7717 (N_7717,N_7320,N_7089);
nand U7718 (N_7718,N_6285,N_6922);
and U7719 (N_7719,N_6690,N_7365);
nand U7720 (N_7720,N_7367,N_6695);
nand U7721 (N_7721,N_6516,N_7318);
nor U7722 (N_7722,N_7324,N_6827);
nand U7723 (N_7723,N_6206,N_6332);
xor U7724 (N_7724,N_6096,N_6118);
xor U7725 (N_7725,N_6397,N_7242);
nor U7726 (N_7726,N_6195,N_6483);
xnor U7727 (N_7727,N_6916,N_6959);
nand U7728 (N_7728,N_6299,N_6943);
nand U7729 (N_7729,N_6440,N_6497);
nor U7730 (N_7730,N_6108,N_7239);
nor U7731 (N_7731,N_6919,N_6477);
and U7732 (N_7732,N_7233,N_6912);
or U7733 (N_7733,N_6267,N_6004);
xnor U7734 (N_7734,N_7183,N_6879);
xor U7735 (N_7735,N_7362,N_6243);
or U7736 (N_7736,N_7433,N_7025);
nor U7737 (N_7737,N_7138,N_7478);
or U7738 (N_7738,N_6968,N_7169);
or U7739 (N_7739,N_7151,N_7179);
and U7740 (N_7740,N_6994,N_7241);
nor U7741 (N_7741,N_6182,N_6370);
or U7742 (N_7742,N_6043,N_6898);
or U7743 (N_7743,N_6860,N_6054);
or U7744 (N_7744,N_6831,N_7333);
or U7745 (N_7745,N_6514,N_6084);
xnor U7746 (N_7746,N_7361,N_7044);
or U7747 (N_7747,N_6758,N_6205);
or U7748 (N_7748,N_7099,N_6948);
nand U7749 (N_7749,N_6875,N_6757);
nand U7750 (N_7750,N_6453,N_6072);
or U7751 (N_7751,N_6718,N_6279);
nor U7752 (N_7752,N_6686,N_7214);
xnor U7753 (N_7753,N_7115,N_6770);
or U7754 (N_7754,N_6805,N_6756);
nor U7755 (N_7755,N_6989,N_6868);
nor U7756 (N_7756,N_6742,N_6221);
nand U7757 (N_7757,N_6637,N_6871);
or U7758 (N_7758,N_6383,N_6520);
nor U7759 (N_7759,N_7414,N_6669);
nor U7760 (N_7760,N_7180,N_6268);
or U7761 (N_7761,N_6733,N_7273);
nor U7762 (N_7762,N_6208,N_7439);
nor U7763 (N_7763,N_6172,N_6403);
or U7764 (N_7764,N_6526,N_6399);
and U7765 (N_7765,N_6507,N_7413);
nand U7766 (N_7766,N_6554,N_6293);
or U7767 (N_7767,N_7295,N_6539);
nor U7768 (N_7768,N_7152,N_6400);
xnor U7769 (N_7769,N_7417,N_7085);
nor U7770 (N_7770,N_6302,N_6836);
nand U7771 (N_7771,N_6548,N_6169);
nor U7772 (N_7772,N_6892,N_6581);
or U7773 (N_7773,N_7109,N_7421);
xor U7774 (N_7774,N_6450,N_6382);
and U7775 (N_7775,N_6044,N_6457);
xor U7776 (N_7776,N_6620,N_6365);
nor U7777 (N_7777,N_6672,N_6797);
xnor U7778 (N_7778,N_6639,N_6940);
xor U7779 (N_7779,N_6819,N_6160);
or U7780 (N_7780,N_6200,N_7011);
nor U7781 (N_7781,N_6336,N_6847);
xnor U7782 (N_7782,N_6622,N_7172);
nor U7783 (N_7783,N_6292,N_7438);
or U7784 (N_7784,N_7059,N_7142);
and U7785 (N_7785,N_6474,N_6381);
or U7786 (N_7786,N_7332,N_7114);
nor U7787 (N_7787,N_6470,N_6327);
or U7788 (N_7788,N_6255,N_6724);
xor U7789 (N_7789,N_7164,N_6523);
or U7790 (N_7790,N_6931,N_6901);
or U7791 (N_7791,N_7312,N_6413);
and U7792 (N_7792,N_6425,N_7272);
or U7793 (N_7793,N_6344,N_7212);
or U7794 (N_7794,N_6655,N_6042);
nand U7795 (N_7795,N_6120,N_6198);
nor U7796 (N_7796,N_7098,N_6738);
xnor U7797 (N_7797,N_6612,N_6380);
or U7798 (N_7798,N_6728,N_7156);
and U7799 (N_7799,N_6012,N_6351);
xor U7800 (N_7800,N_7018,N_7418);
and U7801 (N_7801,N_6816,N_6708);
and U7802 (N_7802,N_6941,N_6379);
or U7803 (N_7803,N_6217,N_6416);
nor U7804 (N_7804,N_7307,N_7005);
nor U7805 (N_7805,N_6853,N_6147);
nand U7806 (N_7806,N_6779,N_7432);
nor U7807 (N_7807,N_6923,N_6091);
xor U7808 (N_7808,N_6030,N_7058);
and U7809 (N_7809,N_6674,N_7240);
xor U7810 (N_7810,N_6804,N_6168);
nor U7811 (N_7811,N_6957,N_7135);
nand U7812 (N_7812,N_7124,N_7290);
nor U7813 (N_7813,N_6862,N_7145);
nor U7814 (N_7814,N_6360,N_6262);
xor U7815 (N_7815,N_6213,N_7469);
and U7816 (N_7816,N_6355,N_6987);
nor U7817 (N_7817,N_7182,N_7030);
nor U7818 (N_7818,N_6276,N_7243);
and U7819 (N_7819,N_7268,N_6492);
or U7820 (N_7820,N_7331,N_7450);
nand U7821 (N_7821,N_6109,N_6277);
nand U7822 (N_7822,N_7467,N_7033);
or U7823 (N_7823,N_6835,N_6036);
xnor U7824 (N_7824,N_7265,N_7302);
nand U7825 (N_7825,N_6723,N_6888);
and U7826 (N_7826,N_6149,N_6194);
or U7827 (N_7827,N_7269,N_6244);
nor U7828 (N_7828,N_7477,N_6246);
or U7829 (N_7829,N_6795,N_6541);
or U7830 (N_7830,N_6855,N_7213);
nand U7831 (N_7831,N_6654,N_6691);
nor U7832 (N_7832,N_6990,N_7282);
or U7833 (N_7833,N_6832,N_6678);
nor U7834 (N_7834,N_6740,N_6627);
nor U7835 (N_7835,N_6323,N_6181);
nor U7836 (N_7836,N_7340,N_7148);
xor U7837 (N_7837,N_7249,N_6095);
nor U7838 (N_7838,N_6152,N_6040);
nor U7839 (N_7839,N_6009,N_6387);
nor U7840 (N_7840,N_6547,N_6501);
xnor U7841 (N_7841,N_7088,N_6165);
and U7842 (N_7842,N_7384,N_7473);
and U7843 (N_7843,N_7146,N_7027);
xnor U7844 (N_7844,N_6132,N_6887);
or U7845 (N_7845,N_6053,N_6431);
nor U7846 (N_7846,N_7415,N_6996);
xnor U7847 (N_7847,N_6116,N_7493);
nand U7848 (N_7848,N_6014,N_7186);
nand U7849 (N_7849,N_6313,N_6648);
xor U7850 (N_7850,N_6406,N_6649);
and U7851 (N_7851,N_7217,N_6890);
nor U7852 (N_7852,N_6752,N_6297);
nor U7853 (N_7853,N_7379,N_6156);
and U7854 (N_7854,N_6993,N_6496);
or U7855 (N_7855,N_6304,N_6226);
or U7856 (N_7856,N_6068,N_6472);
or U7857 (N_7857,N_6384,N_6897);
nand U7858 (N_7858,N_7262,N_7470);
and U7859 (N_7859,N_6433,N_6722);
or U7860 (N_7860,N_6926,N_7451);
or U7861 (N_7861,N_7274,N_6841);
xor U7862 (N_7862,N_7095,N_6443);
or U7863 (N_7863,N_6807,N_7330);
nand U7864 (N_7864,N_6867,N_7102);
nor U7865 (N_7865,N_6749,N_7364);
xnor U7866 (N_7866,N_6814,N_6503);
xnor U7867 (N_7867,N_7032,N_6322);
nand U7868 (N_7868,N_6687,N_7143);
nand U7869 (N_7869,N_6211,N_6330);
xnor U7870 (N_7870,N_6833,N_7278);
nor U7871 (N_7871,N_6252,N_6598);
or U7872 (N_7872,N_6130,N_7258);
or U7873 (N_7873,N_6527,N_7389);
nor U7874 (N_7874,N_6505,N_7189);
or U7875 (N_7875,N_7225,N_7490);
or U7876 (N_7876,N_6759,N_6067);
xor U7877 (N_7877,N_6907,N_6444);
or U7878 (N_7878,N_6801,N_6930);
and U7879 (N_7879,N_6446,N_6538);
xnor U7880 (N_7880,N_6820,N_7371);
nand U7881 (N_7881,N_7084,N_6809);
xor U7882 (N_7882,N_7053,N_7147);
nand U7883 (N_7883,N_6666,N_6092);
or U7884 (N_7884,N_7106,N_6677);
and U7885 (N_7885,N_6488,N_6145);
nand U7886 (N_7886,N_6469,N_7453);
nor U7887 (N_7887,N_7052,N_7236);
nand U7888 (N_7888,N_7035,N_6069);
and U7889 (N_7889,N_6032,N_6362);
or U7890 (N_7890,N_6151,N_7121);
nor U7891 (N_7891,N_6633,N_6052);
xor U7892 (N_7892,N_6761,N_7356);
or U7893 (N_7893,N_6811,N_6974);
nor U7894 (N_7894,N_6729,N_6410);
xor U7895 (N_7895,N_7194,N_6646);
xnor U7896 (N_7896,N_6078,N_6730);
or U7897 (N_7897,N_6434,N_6693);
or U7898 (N_7898,N_7130,N_7430);
nor U7899 (N_7899,N_6000,N_6341);
or U7900 (N_7900,N_6998,N_7495);
nand U7901 (N_7901,N_6813,N_7251);
and U7902 (N_7902,N_6143,N_7128);
or U7903 (N_7903,N_7075,N_6303);
and U7904 (N_7904,N_6239,N_6549);
nand U7905 (N_7905,N_6668,N_7488);
nor U7906 (N_7906,N_6721,N_6202);
nor U7907 (N_7907,N_6808,N_7184);
or U7908 (N_7908,N_7402,N_6294);
and U7909 (N_7909,N_6588,N_7068);
nand U7910 (N_7910,N_6929,N_6185);
nand U7911 (N_7911,N_6251,N_6367);
nand U7912 (N_7912,N_6359,N_7393);
nor U7913 (N_7913,N_7049,N_7398);
or U7914 (N_7914,N_7036,N_6110);
or U7915 (N_7915,N_6942,N_6596);
or U7916 (N_7916,N_6714,N_6296);
nor U7917 (N_7917,N_7425,N_6924);
xor U7918 (N_7918,N_7083,N_7008);
xor U7919 (N_7919,N_6796,N_6580);
nor U7920 (N_7920,N_6114,N_6778);
nand U7921 (N_7921,N_6423,N_7374);
nor U7922 (N_7922,N_7237,N_6073);
nand U7923 (N_7923,N_7141,N_6938);
nand U7924 (N_7924,N_6951,N_6465);
xnor U7925 (N_7925,N_6225,N_7079);
or U7926 (N_7926,N_6245,N_6468);
xor U7927 (N_7927,N_6736,N_7459);
nor U7928 (N_7928,N_7038,N_6715);
nand U7929 (N_7929,N_6945,N_6081);
nand U7930 (N_7930,N_7074,N_6645);
xnor U7931 (N_7931,N_6272,N_6316);
nor U7932 (N_7932,N_6568,N_6982);
nor U7933 (N_7933,N_6102,N_6259);
or U7934 (N_7934,N_6121,N_7283);
and U7935 (N_7935,N_7449,N_6676);
or U7936 (N_7936,N_7013,N_7031);
nand U7937 (N_7937,N_6700,N_6290);
and U7938 (N_7938,N_7420,N_6920);
xnor U7939 (N_7939,N_6845,N_6621);
nor U7940 (N_7940,N_6792,N_6510);
and U7941 (N_7941,N_7020,N_6318);
and U7942 (N_7942,N_6891,N_7210);
xor U7943 (N_7943,N_6219,N_6155);
xnor U7944 (N_7944,N_6126,N_6947);
or U7945 (N_7945,N_6261,N_6842);
and U7946 (N_7946,N_6448,N_7140);
xnor U7947 (N_7947,N_7256,N_6463);
or U7948 (N_7948,N_6562,N_6902);
and U7949 (N_7949,N_6464,N_6656);
nor U7950 (N_7950,N_6958,N_6532);
xnor U7951 (N_7951,N_7261,N_6489);
nor U7952 (N_7952,N_6766,N_6573);
xor U7953 (N_7953,N_6768,N_7461);
or U7954 (N_7954,N_6024,N_7131);
nor U7955 (N_7955,N_6320,N_6641);
and U7956 (N_7956,N_7474,N_6932);
and U7957 (N_7957,N_6428,N_6582);
and U7958 (N_7958,N_6513,N_6927);
and U7959 (N_7959,N_7024,N_7171);
or U7960 (N_7960,N_6579,N_7328);
nand U7961 (N_7961,N_6935,N_6154);
nor U7962 (N_7962,N_7270,N_6552);
xor U7963 (N_7963,N_7325,N_6949);
and U7964 (N_7964,N_7369,N_6524);
nand U7965 (N_7965,N_6372,N_6720);
nor U7966 (N_7966,N_6905,N_6908);
nand U7967 (N_7967,N_7494,N_6100);
or U7968 (N_7968,N_6572,N_6339);
xnor U7969 (N_7969,N_6241,N_6311);
nor U7970 (N_7970,N_6305,N_7029);
xnor U7971 (N_7971,N_7203,N_6970);
nor U7972 (N_7972,N_6673,N_6087);
nand U7973 (N_7973,N_7313,N_6170);
xnor U7974 (N_7974,N_6363,N_6577);
xnor U7975 (N_7975,N_7344,N_6103);
nor U7976 (N_7976,N_7132,N_6148);
or U7977 (N_7977,N_6543,N_6821);
and U7978 (N_7978,N_6986,N_6881);
xor U7979 (N_7979,N_6553,N_6484);
and U7980 (N_7980,N_6675,N_7190);
or U7981 (N_7981,N_6089,N_6333);
xnor U7982 (N_7982,N_6972,N_6017);
nor U7983 (N_7983,N_6530,N_6124);
nand U7984 (N_7984,N_7481,N_6368);
xor U7985 (N_7985,N_7034,N_6802);
nor U7986 (N_7986,N_6224,N_6634);
xor U7987 (N_7987,N_6106,N_7159);
xor U7988 (N_7988,N_7196,N_6015);
xnor U7989 (N_7989,N_6780,N_6480);
and U7990 (N_7990,N_6364,N_7322);
or U7991 (N_7991,N_7308,N_6186);
nor U7992 (N_7992,N_6734,N_7063);
nor U7993 (N_7993,N_6046,N_7126);
nor U7994 (N_7994,N_6661,N_7291);
nor U7995 (N_7995,N_6085,N_6455);
nand U7996 (N_7996,N_7304,N_6326);
xnor U7997 (N_7997,N_7298,N_6033);
or U7998 (N_7998,N_6049,N_7226);
xnor U7999 (N_7999,N_7054,N_7431);
xnor U8000 (N_8000,N_6402,N_6981);
nand U8001 (N_8001,N_7436,N_6746);
or U8002 (N_8002,N_7197,N_6878);
nand U8003 (N_8003,N_6437,N_7426);
nor U8004 (N_8004,N_6090,N_6964);
and U8005 (N_8005,N_6430,N_7276);
or U8006 (N_8006,N_6021,N_7348);
and U8007 (N_8007,N_6201,N_6777);
and U8008 (N_8008,N_6741,N_7353);
nand U8009 (N_8009,N_6061,N_7317);
or U8010 (N_8010,N_6896,N_6946);
xor U8011 (N_8011,N_6317,N_7211);
nand U8012 (N_8012,N_6850,N_6391);
or U8013 (N_8013,N_6608,N_6140);
or U8014 (N_8014,N_7167,N_7097);
and U8015 (N_8015,N_7078,N_7462);
xor U8016 (N_8016,N_7234,N_6432);
xor U8017 (N_8017,N_6776,N_7207);
nor U8018 (N_8018,N_6535,N_6002);
or U8019 (N_8019,N_7428,N_6347);
and U8020 (N_8020,N_7153,N_6112);
nand U8021 (N_8021,N_6569,N_7014);
nand U8022 (N_8022,N_7103,N_7343);
and U8023 (N_8023,N_6233,N_6618);
or U8024 (N_8024,N_7404,N_6984);
nor U8025 (N_8025,N_7230,N_6550);
xor U8026 (N_8026,N_6237,N_7386);
nor U8027 (N_8027,N_7163,N_7155);
xor U8028 (N_8028,N_7041,N_6157);
nand U8029 (N_8029,N_7319,N_6704);
or U8030 (N_8030,N_6369,N_7166);
and U8031 (N_8031,N_7017,N_7277);
xnor U8032 (N_8032,N_6020,N_6066);
nand U8033 (N_8033,N_7080,N_7375);
nand U8034 (N_8034,N_6424,N_6914);
nor U8035 (N_8035,N_6719,N_6849);
and U8036 (N_8036,N_6952,N_6479);
and U8037 (N_8037,N_6843,N_6559);
or U8038 (N_8038,N_6404,N_6954);
or U8039 (N_8039,N_6153,N_6088);
and U8040 (N_8040,N_7437,N_7200);
xnor U8041 (N_8041,N_6702,N_6765);
nand U8042 (N_8042,N_6624,N_7445);
xor U8043 (N_8043,N_6487,N_7458);
nor U8044 (N_8044,N_7223,N_7382);
xnor U8045 (N_8045,N_6176,N_6013);
and U8046 (N_8046,N_6576,N_6405);
xnor U8047 (N_8047,N_6230,N_6545);
and U8048 (N_8048,N_6447,N_7039);
and U8049 (N_8049,N_7134,N_6461);
xor U8050 (N_8050,N_6605,N_7026);
or U8051 (N_8051,N_7127,N_6418);
and U8052 (N_8052,N_6122,N_6458);
and U8053 (N_8053,N_7007,N_7329);
nor U8054 (N_8054,N_6599,N_6865);
or U8055 (N_8055,N_7410,N_7457);
xnor U8056 (N_8056,N_6396,N_6232);
and U8057 (N_8057,N_6625,N_6197);
or U8058 (N_8058,N_7409,N_6583);
or U8059 (N_8059,N_6979,N_7275);
nand U8060 (N_8060,N_7176,N_6781);
nand U8061 (N_8061,N_6711,N_7069);
or U8062 (N_8062,N_7118,N_6574);
xor U8063 (N_8063,N_6762,N_6975);
and U8064 (N_8064,N_6408,N_6846);
nor U8065 (N_8065,N_7475,N_6522);
or U8066 (N_8066,N_6223,N_6308);
and U8067 (N_8067,N_6371,N_7094);
and U8068 (N_8068,N_7122,N_7178);
and U8069 (N_8069,N_6070,N_6791);
or U8070 (N_8070,N_6883,N_6502);
xor U8071 (N_8071,N_6234,N_7055);
nor U8072 (N_8072,N_7193,N_6698);
xor U8073 (N_8073,N_7257,N_7228);
or U8074 (N_8074,N_6358,N_6774);
and U8075 (N_8075,N_6075,N_6560);
nor U8076 (N_8076,N_6899,N_6452);
and U8077 (N_8077,N_7247,N_6595);
nor U8078 (N_8078,N_6851,N_6521);
nand U8079 (N_8079,N_6499,N_6269);
nand U8080 (N_8080,N_6378,N_7440);
xnor U8081 (N_8081,N_6682,N_6460);
and U8082 (N_8082,N_7394,N_6703);
nand U8083 (N_8083,N_6790,N_6544);
xor U8084 (N_8084,N_6771,N_7070);
nor U8085 (N_8085,N_7259,N_6712);
nand U8086 (N_8086,N_6177,N_6515);
xnor U8087 (N_8087,N_7113,N_7472);
or U8088 (N_8088,N_7408,N_6872);
or U8089 (N_8089,N_7363,N_6658);
nor U8090 (N_8090,N_7170,N_6615);
or U8091 (N_8091,N_7405,N_6031);
and U8092 (N_8092,N_7076,N_7305);
xor U8093 (N_8093,N_6192,N_6353);
xor U8094 (N_8094,N_6707,N_7181);
and U8095 (N_8095,N_6636,N_6657);
nand U8096 (N_8096,N_6629,N_7381);
and U8097 (N_8097,N_7390,N_6466);
nor U8098 (N_8098,N_6257,N_6074);
nand U8099 (N_8099,N_6047,N_6863);
nand U8100 (N_8100,N_6034,N_7455);
nand U8101 (N_8101,N_7496,N_6753);
and U8102 (N_8102,N_7339,N_6204);
or U8103 (N_8103,N_7423,N_7401);
nor U8104 (N_8104,N_6886,N_7221);
xnor U8105 (N_8105,N_7154,N_6667);
and U8106 (N_8106,N_7185,N_7411);
nor U8107 (N_8107,N_6895,N_6944);
nand U8108 (N_8108,N_6511,N_6884);
xnor U8109 (N_8109,N_7009,N_7012);
or U8110 (N_8110,N_7463,N_6490);
and U8111 (N_8111,N_7351,N_7111);
nor U8112 (N_8112,N_6529,N_6138);
nand U8113 (N_8113,N_6476,N_7388);
nor U8114 (N_8114,N_6653,N_6953);
and U8115 (N_8115,N_6350,N_7271);
nor U8116 (N_8116,N_6785,N_6315);
or U8117 (N_8117,N_6662,N_6041);
nor U8118 (N_8118,N_6393,N_6026);
xnor U8119 (N_8119,N_6939,N_6858);
xnor U8120 (N_8120,N_6745,N_6893);
and U8121 (N_8121,N_6481,N_6743);
nor U8122 (N_8122,N_7392,N_6619);
xnor U8123 (N_8123,N_6345,N_6617);
and U8124 (N_8124,N_6584,N_6603);
nand U8125 (N_8125,N_6542,N_7376);
or U8126 (N_8126,N_6445,N_6471);
xnor U8127 (N_8127,N_6135,N_7028);
and U8128 (N_8128,N_6659,N_6962);
nor U8129 (N_8129,N_6429,N_7466);
or U8130 (N_8130,N_6025,N_6008);
and U8131 (N_8131,N_6727,N_7334);
and U8132 (N_8132,N_6216,N_7460);
xnor U8133 (N_8133,N_6551,N_6787);
nand U8134 (N_8134,N_7263,N_6512);
nor U8135 (N_8135,N_6844,N_7485);
nor U8136 (N_8136,N_7144,N_7368);
or U8137 (N_8137,N_6105,N_6356);
and U8138 (N_8138,N_7266,N_6079);
and U8139 (N_8139,N_6001,N_7406);
nand U8140 (N_8140,N_7202,N_7161);
or U8141 (N_8141,N_6909,N_7468);
and U8142 (N_8142,N_6783,N_6540);
and U8143 (N_8143,N_6822,N_7370);
xor U8144 (N_8144,N_7366,N_6885);
nand U8145 (N_8145,N_6586,N_6411);
nor U8146 (N_8146,N_7123,N_7077);
or U8147 (N_8147,N_7006,N_6212);
nand U8148 (N_8148,N_6876,N_6298);
xor U8149 (N_8149,N_6533,N_7220);
xor U8150 (N_8150,N_7224,N_6028);
xor U8151 (N_8151,N_7464,N_6179);
nand U8152 (N_8152,N_6306,N_6337);
nor U8153 (N_8153,N_6988,N_6856);
or U8154 (N_8154,N_7067,N_6632);
xnor U8155 (N_8155,N_6799,N_6818);
nor U8156 (N_8156,N_6528,N_6697);
and U8157 (N_8157,N_6537,N_6407);
nand U8158 (N_8158,N_7252,N_6057);
and U8159 (N_8159,N_6889,N_6055);
nand U8160 (N_8160,N_7285,N_6564);
xor U8161 (N_8161,N_6546,N_6717);
and U8162 (N_8162,N_6628,N_7301);
nor U8163 (N_8163,N_6166,N_6188);
nor U8164 (N_8164,N_6436,N_6183);
nand U8165 (N_8165,N_6254,N_6451);
and U8166 (N_8166,N_6491,N_7321);
xnor U8167 (N_8167,N_7377,N_6504);
and U8168 (N_8168,N_6973,N_6417);
and U8169 (N_8169,N_7341,N_7105);
nand U8170 (N_8170,N_6731,N_6184);
nor U8171 (N_8171,N_6309,N_6800);
xor U8172 (N_8172,N_6593,N_7378);
and U8173 (N_8173,N_6978,N_7043);
and U8174 (N_8174,N_6220,N_6454);
and U8175 (N_8175,N_7397,N_7104);
and U8176 (N_8176,N_7107,N_6018);
nand U8177 (N_8177,N_7093,N_7288);
or U8178 (N_8178,N_7229,N_6685);
or U8179 (N_8179,N_6189,N_7000);
or U8180 (N_8180,N_6190,N_7326);
xor U8181 (N_8181,N_6980,N_7072);
and U8182 (N_8182,N_7057,N_7306);
nor U8183 (N_8183,N_6366,N_6060);
xnor U8184 (N_8184,N_6348,N_6825);
nor U8185 (N_8185,N_6754,N_7407);
and U8186 (N_8186,N_6343,N_6955);
nor U8187 (N_8187,N_7442,N_7108);
nand U8188 (N_8188,N_6670,N_6394);
and U8189 (N_8189,N_6449,N_6735);
or U8190 (N_8190,N_6824,N_6921);
nand U8191 (N_8191,N_6346,N_7023);
or U8192 (N_8192,N_7292,N_6307);
and U8193 (N_8193,N_6193,N_6222);
or U8194 (N_8194,N_6873,N_6161);
or U8195 (N_8195,N_6591,N_7100);
xor U8196 (N_8196,N_7479,N_6614);
xnor U8197 (N_8197,N_6663,N_6815);
nor U8198 (N_8198,N_6324,N_6038);
or U8199 (N_8199,N_6142,N_6651);
nor U8200 (N_8200,N_6175,N_6500);
xnor U8201 (N_8201,N_7137,N_6874);
nor U8202 (N_8202,N_6482,N_6123);
or U8203 (N_8203,N_6125,N_7395);
nand U8204 (N_8204,N_6950,N_6601);
xnor U8205 (N_8205,N_6373,N_6664);
and U8206 (N_8206,N_7125,N_7385);
and U8207 (N_8207,N_6709,N_6274);
nor U8208 (N_8208,N_6839,N_7427);
and U8209 (N_8209,N_6062,N_6969);
and U8210 (N_8210,N_7349,N_6442);
nand U8211 (N_8211,N_6284,N_7116);
xnor U8212 (N_8212,N_7120,N_7447);
nor U8213 (N_8213,N_7177,N_6180);
and U8214 (N_8214,N_7187,N_6287);
or U8215 (N_8215,N_6422,N_7350);
and U8216 (N_8216,N_6301,N_7173);
or U8217 (N_8217,N_7300,N_7323);
nand U8218 (N_8218,N_6840,N_7092);
nand U8219 (N_8219,N_6375,N_6097);
nor U8220 (N_8220,N_6071,N_6848);
xor U8221 (N_8221,N_7065,N_6291);
nor U8222 (N_8222,N_6877,N_6903);
and U8223 (N_8223,N_7279,N_6249);
and U8224 (N_8224,N_6963,N_7498);
nor U8225 (N_8225,N_7219,N_7246);
and U8226 (N_8226,N_6162,N_6933);
nand U8227 (N_8227,N_6271,N_7096);
or U8228 (N_8228,N_7337,N_7019);
and U8229 (N_8229,N_7253,N_6258);
nand U8230 (N_8230,N_7206,N_6910);
xor U8231 (N_8231,N_7482,N_6354);
nand U8232 (N_8232,N_6409,N_6113);
or U8233 (N_8233,N_6325,N_7199);
and U8234 (N_8234,N_6737,N_7480);
or U8235 (N_8235,N_6508,N_6273);
xnor U8236 (N_8236,N_7129,N_6710);
nand U8237 (N_8237,N_6556,N_6859);
nand U8238 (N_8238,N_6328,N_6421);
xor U8239 (N_8239,N_6965,N_6692);
or U8240 (N_8240,N_7360,N_7042);
or U8241 (N_8241,N_6684,N_6310);
nand U8242 (N_8242,N_7354,N_7476);
xor U8243 (N_8243,N_7314,N_6915);
or U8244 (N_8244,N_7216,N_7248);
and U8245 (N_8245,N_7162,N_6264);
and U8246 (N_8246,N_7347,N_7150);
and U8247 (N_8247,N_7345,N_7062);
xor U8248 (N_8248,N_6594,N_6671);
and U8249 (N_8249,N_7336,N_6961);
and U8250 (N_8250,N_7469,N_6861);
nand U8251 (N_8251,N_6928,N_7217);
nand U8252 (N_8252,N_6517,N_6770);
and U8253 (N_8253,N_6248,N_6830);
or U8254 (N_8254,N_6307,N_6810);
or U8255 (N_8255,N_6543,N_6904);
xor U8256 (N_8256,N_6054,N_6316);
xnor U8257 (N_8257,N_6580,N_6413);
nand U8258 (N_8258,N_6985,N_7432);
or U8259 (N_8259,N_7297,N_6704);
or U8260 (N_8260,N_6303,N_6191);
xnor U8261 (N_8261,N_7273,N_6690);
nand U8262 (N_8262,N_6189,N_6826);
and U8263 (N_8263,N_7013,N_6977);
nand U8264 (N_8264,N_6289,N_7340);
and U8265 (N_8265,N_7098,N_6289);
or U8266 (N_8266,N_6004,N_6282);
nand U8267 (N_8267,N_6845,N_6699);
and U8268 (N_8268,N_7363,N_6974);
xor U8269 (N_8269,N_6408,N_6963);
xnor U8270 (N_8270,N_6970,N_6913);
nor U8271 (N_8271,N_7158,N_6949);
or U8272 (N_8272,N_7376,N_6308);
or U8273 (N_8273,N_7296,N_6170);
nand U8274 (N_8274,N_7289,N_6767);
and U8275 (N_8275,N_6024,N_7336);
xnor U8276 (N_8276,N_6948,N_6509);
or U8277 (N_8277,N_6719,N_6447);
xor U8278 (N_8278,N_6061,N_6916);
or U8279 (N_8279,N_6242,N_6883);
xnor U8280 (N_8280,N_6892,N_6696);
and U8281 (N_8281,N_6920,N_6796);
nand U8282 (N_8282,N_6959,N_6870);
xnor U8283 (N_8283,N_6185,N_6820);
nand U8284 (N_8284,N_6251,N_6014);
nand U8285 (N_8285,N_6776,N_6685);
xor U8286 (N_8286,N_6986,N_6919);
nand U8287 (N_8287,N_6368,N_6765);
nand U8288 (N_8288,N_6642,N_7131);
nor U8289 (N_8289,N_7139,N_6543);
xnor U8290 (N_8290,N_6186,N_7135);
and U8291 (N_8291,N_6993,N_7019);
nand U8292 (N_8292,N_6937,N_7095);
and U8293 (N_8293,N_6266,N_7335);
nand U8294 (N_8294,N_7453,N_7228);
xnor U8295 (N_8295,N_6364,N_7294);
nor U8296 (N_8296,N_6932,N_6873);
nand U8297 (N_8297,N_6197,N_7240);
xnor U8298 (N_8298,N_6200,N_6163);
xnor U8299 (N_8299,N_7292,N_6889);
or U8300 (N_8300,N_6981,N_6704);
nand U8301 (N_8301,N_6442,N_6352);
nor U8302 (N_8302,N_6211,N_7190);
nor U8303 (N_8303,N_6289,N_6118);
nand U8304 (N_8304,N_7436,N_7062);
nand U8305 (N_8305,N_7054,N_7253);
and U8306 (N_8306,N_7217,N_6551);
or U8307 (N_8307,N_7429,N_6013);
nand U8308 (N_8308,N_6069,N_6846);
nand U8309 (N_8309,N_6213,N_7131);
and U8310 (N_8310,N_6881,N_6454);
nand U8311 (N_8311,N_6428,N_7102);
nor U8312 (N_8312,N_6269,N_6803);
xnor U8313 (N_8313,N_7196,N_6487);
or U8314 (N_8314,N_7185,N_6076);
and U8315 (N_8315,N_7475,N_6311);
and U8316 (N_8316,N_6732,N_6863);
and U8317 (N_8317,N_7450,N_6642);
nor U8318 (N_8318,N_7098,N_6824);
or U8319 (N_8319,N_6949,N_6782);
and U8320 (N_8320,N_7304,N_6285);
or U8321 (N_8321,N_7119,N_6366);
and U8322 (N_8322,N_6465,N_7316);
nor U8323 (N_8323,N_7393,N_6848);
and U8324 (N_8324,N_6776,N_6521);
nand U8325 (N_8325,N_7296,N_6249);
and U8326 (N_8326,N_6346,N_7438);
and U8327 (N_8327,N_7009,N_7002);
or U8328 (N_8328,N_6492,N_6255);
xnor U8329 (N_8329,N_6182,N_6931);
nor U8330 (N_8330,N_6245,N_6392);
xnor U8331 (N_8331,N_6917,N_7443);
xnor U8332 (N_8332,N_7334,N_7411);
nor U8333 (N_8333,N_6329,N_6431);
nand U8334 (N_8334,N_7465,N_6584);
and U8335 (N_8335,N_7156,N_6899);
or U8336 (N_8336,N_7194,N_6658);
nand U8337 (N_8337,N_6892,N_6158);
and U8338 (N_8338,N_6682,N_7497);
and U8339 (N_8339,N_6821,N_6294);
and U8340 (N_8340,N_6124,N_6431);
or U8341 (N_8341,N_6883,N_6132);
or U8342 (N_8342,N_6312,N_6139);
or U8343 (N_8343,N_6245,N_6146);
nand U8344 (N_8344,N_6623,N_6979);
nand U8345 (N_8345,N_7379,N_6590);
or U8346 (N_8346,N_7095,N_7275);
nor U8347 (N_8347,N_7428,N_6528);
or U8348 (N_8348,N_7157,N_7067);
or U8349 (N_8349,N_6857,N_6293);
nand U8350 (N_8350,N_7115,N_6452);
nor U8351 (N_8351,N_7101,N_6122);
xnor U8352 (N_8352,N_6862,N_6133);
nor U8353 (N_8353,N_6062,N_7020);
nor U8354 (N_8354,N_6135,N_7201);
and U8355 (N_8355,N_7270,N_6058);
and U8356 (N_8356,N_7155,N_6704);
nand U8357 (N_8357,N_6110,N_6243);
xor U8358 (N_8358,N_6965,N_6330);
xnor U8359 (N_8359,N_6359,N_7252);
nand U8360 (N_8360,N_6963,N_7411);
nor U8361 (N_8361,N_6833,N_6769);
nand U8362 (N_8362,N_6176,N_6834);
and U8363 (N_8363,N_6241,N_7325);
xor U8364 (N_8364,N_6408,N_7084);
and U8365 (N_8365,N_6989,N_6679);
nor U8366 (N_8366,N_6692,N_6474);
nor U8367 (N_8367,N_6665,N_7254);
and U8368 (N_8368,N_6480,N_6259);
xor U8369 (N_8369,N_6205,N_7400);
xor U8370 (N_8370,N_6678,N_7093);
and U8371 (N_8371,N_6911,N_7237);
nand U8372 (N_8372,N_7007,N_6280);
and U8373 (N_8373,N_7436,N_6482);
or U8374 (N_8374,N_7241,N_6853);
and U8375 (N_8375,N_6936,N_6372);
nor U8376 (N_8376,N_6286,N_7460);
xor U8377 (N_8377,N_7295,N_7338);
or U8378 (N_8378,N_7407,N_6230);
nand U8379 (N_8379,N_7359,N_6099);
or U8380 (N_8380,N_6190,N_7373);
and U8381 (N_8381,N_6603,N_7219);
nand U8382 (N_8382,N_6746,N_6803);
nor U8383 (N_8383,N_7185,N_6522);
or U8384 (N_8384,N_7011,N_6005);
nor U8385 (N_8385,N_6864,N_6814);
nand U8386 (N_8386,N_6581,N_6030);
or U8387 (N_8387,N_6419,N_7180);
nand U8388 (N_8388,N_6739,N_7371);
and U8389 (N_8389,N_6679,N_6297);
nand U8390 (N_8390,N_7163,N_7145);
and U8391 (N_8391,N_7332,N_6213);
and U8392 (N_8392,N_6880,N_6676);
and U8393 (N_8393,N_7330,N_7115);
xor U8394 (N_8394,N_6371,N_7112);
and U8395 (N_8395,N_7390,N_6290);
and U8396 (N_8396,N_6998,N_6595);
and U8397 (N_8397,N_7224,N_7135);
and U8398 (N_8398,N_6273,N_6308);
and U8399 (N_8399,N_6263,N_7447);
and U8400 (N_8400,N_6906,N_6172);
nand U8401 (N_8401,N_6400,N_7036);
nor U8402 (N_8402,N_7236,N_7484);
nor U8403 (N_8403,N_6196,N_7119);
nor U8404 (N_8404,N_7326,N_6828);
nand U8405 (N_8405,N_6938,N_7440);
and U8406 (N_8406,N_6528,N_7174);
or U8407 (N_8407,N_7420,N_6501);
nor U8408 (N_8408,N_6181,N_6039);
nor U8409 (N_8409,N_6435,N_7205);
or U8410 (N_8410,N_7306,N_7222);
nor U8411 (N_8411,N_7494,N_7292);
nor U8412 (N_8412,N_7016,N_7020);
and U8413 (N_8413,N_6610,N_6475);
or U8414 (N_8414,N_6864,N_7282);
or U8415 (N_8415,N_6309,N_7367);
nor U8416 (N_8416,N_7009,N_6314);
xor U8417 (N_8417,N_7035,N_7317);
nor U8418 (N_8418,N_6881,N_6562);
xor U8419 (N_8419,N_6592,N_7025);
nand U8420 (N_8420,N_7400,N_6371);
or U8421 (N_8421,N_6168,N_6994);
nand U8422 (N_8422,N_6109,N_6414);
or U8423 (N_8423,N_6125,N_6394);
nand U8424 (N_8424,N_7010,N_6454);
nand U8425 (N_8425,N_6173,N_6806);
nand U8426 (N_8426,N_7065,N_7193);
and U8427 (N_8427,N_7343,N_7123);
nand U8428 (N_8428,N_7470,N_7479);
or U8429 (N_8429,N_7135,N_7221);
nor U8430 (N_8430,N_7296,N_6252);
or U8431 (N_8431,N_6180,N_6029);
or U8432 (N_8432,N_6148,N_7361);
nand U8433 (N_8433,N_6111,N_6737);
or U8434 (N_8434,N_7308,N_6843);
nand U8435 (N_8435,N_7341,N_6597);
or U8436 (N_8436,N_6096,N_6296);
or U8437 (N_8437,N_6953,N_6210);
nor U8438 (N_8438,N_7099,N_7066);
xor U8439 (N_8439,N_7366,N_6756);
nand U8440 (N_8440,N_6190,N_6422);
nand U8441 (N_8441,N_6409,N_6487);
xor U8442 (N_8442,N_7401,N_7209);
nor U8443 (N_8443,N_6039,N_6946);
xnor U8444 (N_8444,N_7234,N_7073);
nor U8445 (N_8445,N_6899,N_6901);
nor U8446 (N_8446,N_6752,N_6142);
nand U8447 (N_8447,N_7485,N_6579);
and U8448 (N_8448,N_6831,N_6462);
nor U8449 (N_8449,N_6430,N_7328);
and U8450 (N_8450,N_6379,N_7302);
nand U8451 (N_8451,N_6608,N_7237);
nand U8452 (N_8452,N_6568,N_6924);
or U8453 (N_8453,N_7012,N_7112);
nand U8454 (N_8454,N_6324,N_6364);
nor U8455 (N_8455,N_7121,N_6723);
xor U8456 (N_8456,N_6513,N_7455);
nand U8457 (N_8457,N_7078,N_6453);
nor U8458 (N_8458,N_6575,N_7355);
nand U8459 (N_8459,N_6239,N_7403);
nor U8460 (N_8460,N_6713,N_6345);
or U8461 (N_8461,N_6916,N_6375);
and U8462 (N_8462,N_7448,N_6631);
nor U8463 (N_8463,N_7003,N_6238);
or U8464 (N_8464,N_7025,N_6323);
xnor U8465 (N_8465,N_6620,N_6389);
or U8466 (N_8466,N_6871,N_6791);
nor U8467 (N_8467,N_6608,N_7067);
or U8468 (N_8468,N_6144,N_7284);
xor U8469 (N_8469,N_6044,N_7144);
nor U8470 (N_8470,N_6517,N_6502);
nand U8471 (N_8471,N_6582,N_6416);
nor U8472 (N_8472,N_6898,N_7232);
nor U8473 (N_8473,N_7356,N_6213);
and U8474 (N_8474,N_7428,N_7413);
and U8475 (N_8475,N_6888,N_6034);
nor U8476 (N_8476,N_6797,N_6805);
nor U8477 (N_8477,N_6964,N_7077);
xor U8478 (N_8478,N_6462,N_6681);
nor U8479 (N_8479,N_7214,N_6237);
nand U8480 (N_8480,N_6583,N_6796);
and U8481 (N_8481,N_6329,N_7091);
nand U8482 (N_8482,N_7055,N_6562);
nand U8483 (N_8483,N_6524,N_6592);
xor U8484 (N_8484,N_6235,N_7285);
nand U8485 (N_8485,N_6437,N_7051);
nand U8486 (N_8486,N_6796,N_6595);
nand U8487 (N_8487,N_6781,N_7002);
or U8488 (N_8488,N_7296,N_6995);
and U8489 (N_8489,N_6289,N_7326);
nor U8490 (N_8490,N_6443,N_6436);
or U8491 (N_8491,N_6423,N_7316);
nand U8492 (N_8492,N_6081,N_7325);
or U8493 (N_8493,N_6809,N_7484);
or U8494 (N_8494,N_7317,N_6472);
or U8495 (N_8495,N_6417,N_6385);
and U8496 (N_8496,N_6359,N_7229);
nand U8497 (N_8497,N_6972,N_6309);
nand U8498 (N_8498,N_6847,N_6430);
nor U8499 (N_8499,N_7090,N_6739);
xnor U8500 (N_8500,N_6259,N_6710);
or U8501 (N_8501,N_6713,N_6684);
nand U8502 (N_8502,N_6846,N_7360);
xnor U8503 (N_8503,N_7249,N_6011);
and U8504 (N_8504,N_6097,N_7308);
nor U8505 (N_8505,N_6369,N_6448);
nand U8506 (N_8506,N_7011,N_6139);
and U8507 (N_8507,N_6445,N_7056);
and U8508 (N_8508,N_6209,N_6665);
nand U8509 (N_8509,N_6498,N_6325);
and U8510 (N_8510,N_6171,N_6578);
nor U8511 (N_8511,N_6288,N_7397);
xnor U8512 (N_8512,N_6631,N_7059);
nand U8513 (N_8513,N_7123,N_7257);
nor U8514 (N_8514,N_6967,N_6554);
nor U8515 (N_8515,N_6760,N_6085);
nor U8516 (N_8516,N_6625,N_6894);
and U8517 (N_8517,N_6073,N_6295);
xor U8518 (N_8518,N_7278,N_7110);
and U8519 (N_8519,N_7262,N_6178);
nand U8520 (N_8520,N_6639,N_6418);
and U8521 (N_8521,N_6413,N_6881);
and U8522 (N_8522,N_6509,N_6693);
nand U8523 (N_8523,N_6881,N_6470);
nor U8524 (N_8524,N_7171,N_7071);
xnor U8525 (N_8525,N_7011,N_6471);
nand U8526 (N_8526,N_7099,N_7063);
nor U8527 (N_8527,N_6625,N_6104);
and U8528 (N_8528,N_6653,N_7474);
or U8529 (N_8529,N_7228,N_6596);
and U8530 (N_8530,N_6207,N_6757);
xnor U8531 (N_8531,N_7055,N_6187);
nand U8532 (N_8532,N_7029,N_6637);
and U8533 (N_8533,N_6010,N_6956);
nand U8534 (N_8534,N_7421,N_6728);
xor U8535 (N_8535,N_7144,N_6172);
and U8536 (N_8536,N_7089,N_7369);
nand U8537 (N_8537,N_7379,N_6267);
and U8538 (N_8538,N_6812,N_6171);
or U8539 (N_8539,N_7368,N_7241);
xor U8540 (N_8540,N_7445,N_6271);
xor U8541 (N_8541,N_6661,N_6297);
or U8542 (N_8542,N_6544,N_7065);
or U8543 (N_8543,N_7077,N_7416);
and U8544 (N_8544,N_6196,N_6097);
nand U8545 (N_8545,N_6487,N_7411);
nor U8546 (N_8546,N_6973,N_7239);
nand U8547 (N_8547,N_7014,N_6512);
nand U8548 (N_8548,N_6403,N_6578);
and U8549 (N_8549,N_6430,N_6366);
nand U8550 (N_8550,N_7084,N_6984);
nor U8551 (N_8551,N_7260,N_6634);
or U8552 (N_8552,N_7046,N_7116);
or U8553 (N_8553,N_6753,N_6411);
nor U8554 (N_8554,N_6272,N_7477);
or U8555 (N_8555,N_7288,N_6206);
nor U8556 (N_8556,N_7072,N_6701);
nor U8557 (N_8557,N_6605,N_6508);
and U8558 (N_8558,N_6146,N_6639);
nor U8559 (N_8559,N_7259,N_7105);
xor U8560 (N_8560,N_6191,N_7299);
nand U8561 (N_8561,N_6873,N_6586);
or U8562 (N_8562,N_7093,N_7324);
or U8563 (N_8563,N_6141,N_6127);
nand U8564 (N_8564,N_6547,N_6222);
nor U8565 (N_8565,N_6314,N_6919);
or U8566 (N_8566,N_6564,N_6747);
or U8567 (N_8567,N_6605,N_6507);
nor U8568 (N_8568,N_6132,N_6268);
xor U8569 (N_8569,N_6765,N_7496);
nand U8570 (N_8570,N_7014,N_7428);
xor U8571 (N_8571,N_6075,N_6836);
xnor U8572 (N_8572,N_6748,N_6079);
nor U8573 (N_8573,N_7276,N_7302);
nand U8574 (N_8574,N_7005,N_6694);
or U8575 (N_8575,N_6766,N_6091);
and U8576 (N_8576,N_6868,N_6152);
nor U8577 (N_8577,N_6745,N_6281);
xnor U8578 (N_8578,N_6755,N_7111);
xnor U8579 (N_8579,N_6628,N_7214);
and U8580 (N_8580,N_6793,N_6181);
xor U8581 (N_8581,N_7373,N_6964);
or U8582 (N_8582,N_7381,N_7020);
and U8583 (N_8583,N_6713,N_7246);
nand U8584 (N_8584,N_7259,N_6876);
nand U8585 (N_8585,N_6429,N_7188);
xnor U8586 (N_8586,N_7431,N_6508);
nand U8587 (N_8587,N_7405,N_7270);
nand U8588 (N_8588,N_6685,N_6431);
nor U8589 (N_8589,N_6952,N_6414);
or U8590 (N_8590,N_7014,N_7007);
and U8591 (N_8591,N_6180,N_6401);
nand U8592 (N_8592,N_6015,N_6698);
and U8593 (N_8593,N_6662,N_6533);
and U8594 (N_8594,N_7281,N_6677);
xor U8595 (N_8595,N_6983,N_6864);
nand U8596 (N_8596,N_7423,N_6140);
and U8597 (N_8597,N_6985,N_7451);
xnor U8598 (N_8598,N_6908,N_6505);
or U8599 (N_8599,N_6740,N_6149);
and U8600 (N_8600,N_6957,N_7343);
or U8601 (N_8601,N_6651,N_7402);
or U8602 (N_8602,N_7267,N_6375);
xnor U8603 (N_8603,N_7003,N_6298);
nor U8604 (N_8604,N_7329,N_6948);
xnor U8605 (N_8605,N_6510,N_6391);
xor U8606 (N_8606,N_6416,N_7424);
xnor U8607 (N_8607,N_6430,N_7001);
xor U8608 (N_8608,N_6018,N_6516);
nand U8609 (N_8609,N_7468,N_7459);
nand U8610 (N_8610,N_7453,N_6913);
xor U8611 (N_8611,N_6835,N_7332);
or U8612 (N_8612,N_7362,N_6155);
and U8613 (N_8613,N_6267,N_7012);
xor U8614 (N_8614,N_6243,N_6196);
and U8615 (N_8615,N_6236,N_6004);
nor U8616 (N_8616,N_6981,N_6203);
and U8617 (N_8617,N_6161,N_7358);
xnor U8618 (N_8618,N_7108,N_7346);
or U8619 (N_8619,N_6616,N_6017);
nor U8620 (N_8620,N_7167,N_6551);
nand U8621 (N_8621,N_6626,N_6877);
nor U8622 (N_8622,N_6753,N_7445);
xnor U8623 (N_8623,N_6276,N_6102);
nand U8624 (N_8624,N_6729,N_6326);
xnor U8625 (N_8625,N_7042,N_7125);
or U8626 (N_8626,N_7322,N_6311);
nor U8627 (N_8627,N_6560,N_6298);
xnor U8628 (N_8628,N_6688,N_6867);
nor U8629 (N_8629,N_6649,N_7390);
or U8630 (N_8630,N_7012,N_6930);
xnor U8631 (N_8631,N_6211,N_6551);
nor U8632 (N_8632,N_6418,N_6367);
nand U8633 (N_8633,N_7309,N_6392);
nor U8634 (N_8634,N_7329,N_6722);
nand U8635 (N_8635,N_6738,N_6329);
or U8636 (N_8636,N_6879,N_6729);
nand U8637 (N_8637,N_7460,N_7094);
or U8638 (N_8638,N_6790,N_7091);
and U8639 (N_8639,N_6725,N_6649);
and U8640 (N_8640,N_7428,N_7185);
or U8641 (N_8641,N_6354,N_7462);
nand U8642 (N_8642,N_6624,N_7112);
nor U8643 (N_8643,N_6106,N_6001);
and U8644 (N_8644,N_6476,N_6509);
or U8645 (N_8645,N_6153,N_6027);
and U8646 (N_8646,N_6820,N_6602);
nand U8647 (N_8647,N_6383,N_6241);
xor U8648 (N_8648,N_7345,N_6481);
or U8649 (N_8649,N_6439,N_6338);
nand U8650 (N_8650,N_6824,N_6267);
nand U8651 (N_8651,N_6198,N_6883);
nand U8652 (N_8652,N_6260,N_6817);
and U8653 (N_8653,N_7107,N_7200);
nor U8654 (N_8654,N_6929,N_6909);
xnor U8655 (N_8655,N_6102,N_6514);
nand U8656 (N_8656,N_7148,N_7398);
or U8657 (N_8657,N_6268,N_6289);
xnor U8658 (N_8658,N_6140,N_6671);
and U8659 (N_8659,N_6818,N_7426);
xor U8660 (N_8660,N_6409,N_7261);
nor U8661 (N_8661,N_6490,N_6726);
or U8662 (N_8662,N_7361,N_6583);
nand U8663 (N_8663,N_7409,N_7225);
or U8664 (N_8664,N_6422,N_6983);
and U8665 (N_8665,N_7081,N_6707);
or U8666 (N_8666,N_6584,N_6868);
nor U8667 (N_8667,N_6731,N_6912);
nor U8668 (N_8668,N_6038,N_6157);
or U8669 (N_8669,N_7253,N_7308);
and U8670 (N_8670,N_6570,N_7276);
and U8671 (N_8671,N_6720,N_6322);
or U8672 (N_8672,N_6663,N_6189);
nor U8673 (N_8673,N_6967,N_7307);
nor U8674 (N_8674,N_6339,N_7290);
and U8675 (N_8675,N_6905,N_6562);
xnor U8676 (N_8676,N_6002,N_6080);
or U8677 (N_8677,N_7263,N_6019);
xnor U8678 (N_8678,N_6291,N_6646);
nor U8679 (N_8679,N_6987,N_6649);
and U8680 (N_8680,N_6128,N_6354);
xnor U8681 (N_8681,N_6619,N_7084);
xnor U8682 (N_8682,N_7147,N_6522);
and U8683 (N_8683,N_6945,N_6708);
or U8684 (N_8684,N_7196,N_6291);
or U8685 (N_8685,N_6919,N_6242);
and U8686 (N_8686,N_7017,N_6024);
nand U8687 (N_8687,N_6043,N_6528);
xnor U8688 (N_8688,N_7023,N_7285);
nand U8689 (N_8689,N_6276,N_7115);
nand U8690 (N_8690,N_6248,N_6388);
and U8691 (N_8691,N_6412,N_7246);
and U8692 (N_8692,N_6644,N_6016);
xor U8693 (N_8693,N_7048,N_6138);
nor U8694 (N_8694,N_6571,N_6747);
and U8695 (N_8695,N_6036,N_7256);
nand U8696 (N_8696,N_6313,N_6155);
or U8697 (N_8697,N_7475,N_6701);
and U8698 (N_8698,N_7407,N_6414);
nand U8699 (N_8699,N_6220,N_7490);
and U8700 (N_8700,N_6451,N_6414);
xnor U8701 (N_8701,N_6814,N_7210);
nor U8702 (N_8702,N_6174,N_6021);
nand U8703 (N_8703,N_6340,N_6832);
or U8704 (N_8704,N_6852,N_6920);
or U8705 (N_8705,N_7475,N_6615);
nor U8706 (N_8706,N_6083,N_6949);
or U8707 (N_8707,N_6038,N_6426);
nor U8708 (N_8708,N_6849,N_6056);
nand U8709 (N_8709,N_6991,N_6696);
xor U8710 (N_8710,N_6479,N_7385);
xnor U8711 (N_8711,N_7042,N_6540);
and U8712 (N_8712,N_7150,N_6018);
nand U8713 (N_8713,N_7271,N_7169);
nor U8714 (N_8714,N_7389,N_6724);
nor U8715 (N_8715,N_6504,N_6875);
nor U8716 (N_8716,N_7373,N_6936);
and U8717 (N_8717,N_6855,N_6981);
xor U8718 (N_8718,N_7263,N_6371);
xnor U8719 (N_8719,N_6205,N_6984);
or U8720 (N_8720,N_7370,N_6039);
nor U8721 (N_8721,N_7384,N_6945);
or U8722 (N_8722,N_6991,N_6863);
nand U8723 (N_8723,N_6321,N_6829);
xnor U8724 (N_8724,N_6468,N_7380);
xnor U8725 (N_8725,N_6154,N_7230);
xor U8726 (N_8726,N_6965,N_7421);
xnor U8727 (N_8727,N_6024,N_6866);
nand U8728 (N_8728,N_6909,N_6890);
and U8729 (N_8729,N_6373,N_7353);
nand U8730 (N_8730,N_6867,N_6791);
xor U8731 (N_8731,N_7433,N_7046);
xnor U8732 (N_8732,N_7157,N_7475);
and U8733 (N_8733,N_6031,N_6328);
or U8734 (N_8734,N_6851,N_7120);
xor U8735 (N_8735,N_7329,N_7029);
xnor U8736 (N_8736,N_7262,N_6463);
nand U8737 (N_8737,N_7119,N_7223);
nor U8738 (N_8738,N_6807,N_6790);
nor U8739 (N_8739,N_6203,N_7006);
nor U8740 (N_8740,N_6680,N_6247);
xor U8741 (N_8741,N_6360,N_6073);
nor U8742 (N_8742,N_6432,N_7205);
xnor U8743 (N_8743,N_6616,N_6938);
xnor U8744 (N_8744,N_6859,N_6520);
xnor U8745 (N_8745,N_7248,N_6960);
nor U8746 (N_8746,N_6336,N_7207);
xor U8747 (N_8747,N_7446,N_6800);
nand U8748 (N_8748,N_6513,N_7388);
or U8749 (N_8749,N_6094,N_6392);
nand U8750 (N_8750,N_6400,N_6666);
and U8751 (N_8751,N_7294,N_6483);
xor U8752 (N_8752,N_6458,N_6218);
or U8753 (N_8753,N_7012,N_7320);
nand U8754 (N_8754,N_6833,N_6548);
nand U8755 (N_8755,N_6264,N_7208);
nor U8756 (N_8756,N_6783,N_6897);
or U8757 (N_8757,N_7264,N_6310);
nor U8758 (N_8758,N_7020,N_7337);
nand U8759 (N_8759,N_6877,N_6078);
nor U8760 (N_8760,N_6947,N_6278);
and U8761 (N_8761,N_6778,N_6549);
nand U8762 (N_8762,N_6421,N_7121);
and U8763 (N_8763,N_7339,N_6380);
or U8764 (N_8764,N_6621,N_6695);
or U8765 (N_8765,N_6502,N_6560);
and U8766 (N_8766,N_6181,N_6208);
nor U8767 (N_8767,N_6528,N_7218);
nor U8768 (N_8768,N_6229,N_7096);
xor U8769 (N_8769,N_6169,N_7094);
xor U8770 (N_8770,N_7461,N_6053);
and U8771 (N_8771,N_6728,N_6939);
nor U8772 (N_8772,N_6553,N_6944);
xnor U8773 (N_8773,N_6211,N_6970);
xor U8774 (N_8774,N_7110,N_6023);
nor U8775 (N_8775,N_6632,N_6289);
or U8776 (N_8776,N_6034,N_7153);
and U8777 (N_8777,N_6485,N_6251);
or U8778 (N_8778,N_6092,N_7391);
nor U8779 (N_8779,N_7382,N_6282);
or U8780 (N_8780,N_6488,N_6046);
nand U8781 (N_8781,N_6893,N_6662);
and U8782 (N_8782,N_6690,N_7459);
nor U8783 (N_8783,N_6682,N_6859);
and U8784 (N_8784,N_6020,N_6958);
nor U8785 (N_8785,N_6344,N_6081);
and U8786 (N_8786,N_6492,N_7359);
or U8787 (N_8787,N_7261,N_6750);
nand U8788 (N_8788,N_7296,N_7121);
xor U8789 (N_8789,N_7068,N_6397);
or U8790 (N_8790,N_7082,N_7326);
or U8791 (N_8791,N_6491,N_6336);
nand U8792 (N_8792,N_6998,N_7359);
nor U8793 (N_8793,N_6213,N_7182);
nand U8794 (N_8794,N_7214,N_6391);
nor U8795 (N_8795,N_6236,N_7152);
or U8796 (N_8796,N_6242,N_6186);
nand U8797 (N_8797,N_7097,N_6079);
or U8798 (N_8798,N_7339,N_6933);
and U8799 (N_8799,N_7281,N_6560);
or U8800 (N_8800,N_6049,N_6377);
nor U8801 (N_8801,N_6251,N_7279);
or U8802 (N_8802,N_6802,N_6589);
or U8803 (N_8803,N_6162,N_7126);
or U8804 (N_8804,N_6115,N_7022);
nand U8805 (N_8805,N_7372,N_7390);
and U8806 (N_8806,N_6780,N_7480);
nor U8807 (N_8807,N_7147,N_7334);
or U8808 (N_8808,N_6694,N_6785);
nor U8809 (N_8809,N_6333,N_6485);
or U8810 (N_8810,N_6410,N_6714);
or U8811 (N_8811,N_7410,N_6971);
nand U8812 (N_8812,N_7393,N_7002);
xor U8813 (N_8813,N_6319,N_6987);
xnor U8814 (N_8814,N_7404,N_6980);
nor U8815 (N_8815,N_7192,N_6325);
nand U8816 (N_8816,N_6860,N_7364);
nor U8817 (N_8817,N_6369,N_6211);
nand U8818 (N_8818,N_7380,N_6636);
xnor U8819 (N_8819,N_6536,N_7232);
nor U8820 (N_8820,N_7376,N_7404);
and U8821 (N_8821,N_6100,N_6836);
nand U8822 (N_8822,N_6249,N_6876);
nand U8823 (N_8823,N_6444,N_6463);
nor U8824 (N_8824,N_6955,N_6454);
xnor U8825 (N_8825,N_6803,N_7222);
and U8826 (N_8826,N_6540,N_6100);
or U8827 (N_8827,N_6533,N_6544);
xor U8828 (N_8828,N_6281,N_6997);
or U8829 (N_8829,N_6039,N_7468);
and U8830 (N_8830,N_7160,N_6327);
nor U8831 (N_8831,N_7253,N_7131);
xnor U8832 (N_8832,N_6304,N_6073);
and U8833 (N_8833,N_6022,N_7322);
nor U8834 (N_8834,N_7143,N_7183);
or U8835 (N_8835,N_6299,N_7242);
and U8836 (N_8836,N_7462,N_6006);
xor U8837 (N_8837,N_7254,N_6044);
and U8838 (N_8838,N_6324,N_7413);
or U8839 (N_8839,N_6812,N_7348);
xnor U8840 (N_8840,N_7437,N_6766);
nand U8841 (N_8841,N_6099,N_7425);
nand U8842 (N_8842,N_7427,N_6548);
nand U8843 (N_8843,N_6886,N_6642);
nor U8844 (N_8844,N_6650,N_6589);
xor U8845 (N_8845,N_6764,N_6514);
nand U8846 (N_8846,N_7074,N_6720);
nand U8847 (N_8847,N_7048,N_6662);
xnor U8848 (N_8848,N_6320,N_6807);
nor U8849 (N_8849,N_6172,N_6660);
or U8850 (N_8850,N_6494,N_6138);
nor U8851 (N_8851,N_7123,N_6330);
or U8852 (N_8852,N_7057,N_6718);
nand U8853 (N_8853,N_6893,N_6980);
nand U8854 (N_8854,N_7050,N_7441);
nand U8855 (N_8855,N_6444,N_7093);
nand U8856 (N_8856,N_6579,N_6267);
and U8857 (N_8857,N_7093,N_6628);
nand U8858 (N_8858,N_7207,N_6523);
xnor U8859 (N_8859,N_6021,N_7196);
nand U8860 (N_8860,N_7211,N_6606);
nand U8861 (N_8861,N_6023,N_6745);
and U8862 (N_8862,N_6252,N_6735);
nor U8863 (N_8863,N_6504,N_6481);
or U8864 (N_8864,N_6414,N_6637);
and U8865 (N_8865,N_7244,N_6799);
and U8866 (N_8866,N_7338,N_6029);
and U8867 (N_8867,N_7482,N_7060);
or U8868 (N_8868,N_6833,N_6146);
and U8869 (N_8869,N_7342,N_7352);
or U8870 (N_8870,N_6827,N_6388);
nor U8871 (N_8871,N_6183,N_6273);
and U8872 (N_8872,N_6294,N_6844);
nor U8873 (N_8873,N_7053,N_6595);
xnor U8874 (N_8874,N_7239,N_6097);
nand U8875 (N_8875,N_7265,N_7333);
or U8876 (N_8876,N_7205,N_6292);
and U8877 (N_8877,N_6524,N_7430);
and U8878 (N_8878,N_7477,N_6039);
and U8879 (N_8879,N_7062,N_6067);
or U8880 (N_8880,N_6404,N_7068);
xor U8881 (N_8881,N_6871,N_7152);
nor U8882 (N_8882,N_6617,N_6632);
nand U8883 (N_8883,N_6903,N_6930);
xor U8884 (N_8884,N_7204,N_7474);
nor U8885 (N_8885,N_6101,N_7003);
xnor U8886 (N_8886,N_6181,N_6915);
xnor U8887 (N_8887,N_6579,N_7222);
or U8888 (N_8888,N_7355,N_7074);
nor U8889 (N_8889,N_7181,N_7146);
nand U8890 (N_8890,N_6024,N_6389);
xor U8891 (N_8891,N_7018,N_6701);
nor U8892 (N_8892,N_6159,N_6518);
or U8893 (N_8893,N_7050,N_7022);
nor U8894 (N_8894,N_6807,N_6302);
nand U8895 (N_8895,N_6912,N_6687);
or U8896 (N_8896,N_6632,N_7166);
nand U8897 (N_8897,N_6897,N_7193);
xor U8898 (N_8898,N_6985,N_6945);
xnor U8899 (N_8899,N_6728,N_6410);
or U8900 (N_8900,N_6908,N_6705);
xnor U8901 (N_8901,N_6725,N_7238);
xnor U8902 (N_8902,N_6445,N_6991);
or U8903 (N_8903,N_7105,N_7284);
or U8904 (N_8904,N_7278,N_6530);
xor U8905 (N_8905,N_6424,N_6093);
or U8906 (N_8906,N_6553,N_7184);
nor U8907 (N_8907,N_7193,N_6585);
xor U8908 (N_8908,N_7458,N_7182);
nor U8909 (N_8909,N_6321,N_6839);
nor U8910 (N_8910,N_7472,N_7389);
nand U8911 (N_8911,N_6551,N_6636);
nand U8912 (N_8912,N_7034,N_7385);
and U8913 (N_8913,N_6995,N_6425);
nand U8914 (N_8914,N_6187,N_6560);
xnor U8915 (N_8915,N_6325,N_6009);
or U8916 (N_8916,N_6994,N_7118);
or U8917 (N_8917,N_7092,N_6707);
nor U8918 (N_8918,N_7095,N_6535);
xnor U8919 (N_8919,N_6571,N_7191);
nand U8920 (N_8920,N_6535,N_6178);
xor U8921 (N_8921,N_6101,N_6685);
xnor U8922 (N_8922,N_6979,N_6013);
and U8923 (N_8923,N_7388,N_7482);
xor U8924 (N_8924,N_6513,N_6448);
nor U8925 (N_8925,N_6823,N_6611);
nor U8926 (N_8926,N_6581,N_7272);
nand U8927 (N_8927,N_6014,N_7035);
nor U8928 (N_8928,N_7314,N_6519);
and U8929 (N_8929,N_6617,N_6544);
xnor U8930 (N_8930,N_7476,N_7006);
xnor U8931 (N_8931,N_7437,N_7332);
xor U8932 (N_8932,N_7428,N_7399);
or U8933 (N_8933,N_7324,N_7221);
and U8934 (N_8934,N_6418,N_6280);
nand U8935 (N_8935,N_7429,N_7015);
nand U8936 (N_8936,N_6358,N_6198);
xor U8937 (N_8937,N_6609,N_6332);
xnor U8938 (N_8938,N_7282,N_6679);
nor U8939 (N_8939,N_6368,N_6605);
nor U8940 (N_8940,N_7425,N_6523);
nand U8941 (N_8941,N_7429,N_6632);
and U8942 (N_8942,N_6036,N_7335);
or U8943 (N_8943,N_7084,N_6864);
nand U8944 (N_8944,N_6202,N_6950);
nand U8945 (N_8945,N_6681,N_6018);
nand U8946 (N_8946,N_6658,N_6282);
and U8947 (N_8947,N_7123,N_6350);
xor U8948 (N_8948,N_6827,N_6900);
or U8949 (N_8949,N_6777,N_6279);
or U8950 (N_8950,N_6141,N_7043);
and U8951 (N_8951,N_6767,N_7306);
nand U8952 (N_8952,N_7417,N_7434);
nand U8953 (N_8953,N_6651,N_7387);
or U8954 (N_8954,N_6815,N_6427);
or U8955 (N_8955,N_6636,N_7462);
or U8956 (N_8956,N_6224,N_6626);
xor U8957 (N_8957,N_6211,N_6101);
or U8958 (N_8958,N_7369,N_6043);
or U8959 (N_8959,N_7305,N_6644);
xnor U8960 (N_8960,N_6257,N_6209);
xnor U8961 (N_8961,N_6551,N_6688);
nor U8962 (N_8962,N_6994,N_7354);
nor U8963 (N_8963,N_6597,N_6668);
nand U8964 (N_8964,N_6301,N_6816);
xnor U8965 (N_8965,N_6586,N_7118);
nor U8966 (N_8966,N_6816,N_6204);
or U8967 (N_8967,N_6421,N_7271);
nand U8968 (N_8968,N_7087,N_6177);
xor U8969 (N_8969,N_6414,N_6422);
and U8970 (N_8970,N_6805,N_6474);
or U8971 (N_8971,N_6725,N_6574);
nand U8972 (N_8972,N_6989,N_6522);
nand U8973 (N_8973,N_6931,N_6991);
nand U8974 (N_8974,N_6249,N_7082);
and U8975 (N_8975,N_6420,N_7471);
xor U8976 (N_8976,N_6677,N_7220);
nor U8977 (N_8977,N_6749,N_6446);
nor U8978 (N_8978,N_6888,N_7401);
and U8979 (N_8979,N_6609,N_6910);
or U8980 (N_8980,N_6325,N_7474);
nand U8981 (N_8981,N_6202,N_7050);
and U8982 (N_8982,N_6337,N_7401);
xnor U8983 (N_8983,N_6523,N_7258);
nand U8984 (N_8984,N_6346,N_6251);
and U8985 (N_8985,N_7058,N_6256);
nand U8986 (N_8986,N_7193,N_6733);
or U8987 (N_8987,N_6849,N_6895);
and U8988 (N_8988,N_7272,N_6710);
or U8989 (N_8989,N_7102,N_6651);
xnor U8990 (N_8990,N_7092,N_7426);
and U8991 (N_8991,N_7172,N_7360);
and U8992 (N_8992,N_7077,N_7176);
and U8993 (N_8993,N_6636,N_6695);
and U8994 (N_8994,N_6789,N_6975);
and U8995 (N_8995,N_6743,N_7495);
and U8996 (N_8996,N_7165,N_6327);
nand U8997 (N_8997,N_7148,N_6815);
xor U8998 (N_8998,N_6388,N_6345);
nand U8999 (N_8999,N_6415,N_7215);
xor U9000 (N_9000,N_7954,N_8957);
xor U9001 (N_9001,N_7889,N_7965);
and U9002 (N_9002,N_7600,N_8244);
nand U9003 (N_9003,N_7761,N_8804);
and U9004 (N_9004,N_7816,N_8519);
xnor U9005 (N_9005,N_7564,N_8882);
nand U9006 (N_9006,N_8399,N_7859);
nor U9007 (N_9007,N_7651,N_8313);
xnor U9008 (N_9008,N_7676,N_7738);
xnor U9009 (N_9009,N_8910,N_8366);
xor U9010 (N_9010,N_8018,N_8294);
nand U9011 (N_9011,N_8765,N_7991);
and U9012 (N_9012,N_8738,N_7573);
nand U9013 (N_9013,N_7733,N_7681);
nor U9014 (N_9014,N_8101,N_7969);
or U9015 (N_9015,N_7932,N_7848);
or U9016 (N_9016,N_8229,N_8601);
or U9017 (N_9017,N_8243,N_8044);
or U9018 (N_9018,N_8794,N_8387);
or U9019 (N_9019,N_7522,N_7687);
and U9020 (N_9020,N_8016,N_7524);
xor U9021 (N_9021,N_7638,N_7942);
nor U9022 (N_9022,N_8041,N_7831);
nand U9023 (N_9023,N_7604,N_7941);
or U9024 (N_9024,N_7565,N_8763);
nand U9025 (N_9025,N_8344,N_7553);
xor U9026 (N_9026,N_8599,N_7963);
and U9027 (N_9027,N_7987,N_7996);
xor U9028 (N_9028,N_8784,N_8972);
nor U9029 (N_9029,N_8071,N_7542);
nor U9030 (N_9030,N_8603,N_8120);
and U9031 (N_9031,N_8452,N_7702);
and U9032 (N_9032,N_7888,N_8797);
or U9033 (N_9033,N_8065,N_8187);
xnor U9034 (N_9034,N_8395,N_8915);
xnor U9035 (N_9035,N_8689,N_8935);
nor U9036 (N_9036,N_8312,N_8571);
xor U9037 (N_9037,N_7914,N_7850);
or U9038 (N_9038,N_7791,N_7578);
xnor U9039 (N_9039,N_7902,N_8131);
and U9040 (N_9040,N_7915,N_8236);
nor U9041 (N_9041,N_8698,N_8655);
nor U9042 (N_9042,N_8114,N_8653);
nor U9043 (N_9043,N_8898,N_8839);
nand U9044 (N_9044,N_8844,N_8221);
xnor U9045 (N_9045,N_8859,N_8628);
or U9046 (N_9046,N_8146,N_7558);
nor U9047 (N_9047,N_8151,N_7627);
nor U9048 (N_9048,N_8752,N_8803);
xnor U9049 (N_9049,N_7943,N_8363);
and U9050 (N_9050,N_8194,N_8122);
nor U9051 (N_9051,N_8412,N_8157);
nand U9052 (N_9052,N_7898,N_8608);
nor U9053 (N_9053,N_7879,N_7547);
nand U9054 (N_9054,N_8212,N_8899);
nand U9055 (N_9055,N_7612,N_8554);
or U9056 (N_9056,N_7555,N_7784);
nand U9057 (N_9057,N_7514,N_8751);
and U9058 (N_9058,N_8549,N_7855);
or U9059 (N_9059,N_8333,N_8838);
or U9060 (N_9060,N_8799,N_7793);
nor U9061 (N_9061,N_7998,N_8465);
nor U9062 (N_9062,N_8654,N_7803);
or U9063 (N_9063,N_8250,N_7680);
xnor U9064 (N_9064,N_8798,N_8248);
xor U9065 (N_9065,N_8315,N_7532);
nor U9066 (N_9066,N_8423,N_8287);
or U9067 (N_9067,N_8460,N_8130);
or U9068 (N_9068,N_8572,N_8106);
xor U9069 (N_9069,N_7725,N_8938);
nor U9070 (N_9070,N_7587,N_7517);
xnor U9071 (N_9071,N_8768,N_7504);
nand U9072 (N_9072,N_8463,N_8953);
nor U9073 (N_9073,N_8304,N_7701);
xor U9074 (N_9074,N_8156,N_7607);
or U9075 (N_9075,N_7974,N_8822);
nand U9076 (N_9076,N_8680,N_8357);
or U9077 (N_9077,N_8781,N_8612);
nand U9078 (N_9078,N_8918,N_8977);
or U9079 (N_9079,N_7823,N_8725);
or U9080 (N_9080,N_8657,N_7561);
and U9081 (N_9081,N_8871,N_7846);
and U9082 (N_9082,N_8547,N_8591);
nand U9083 (N_9083,N_8185,N_7637);
xnor U9084 (N_9084,N_8389,N_8636);
xnor U9085 (N_9085,N_7628,N_8046);
nor U9086 (N_9086,N_8284,N_8192);
or U9087 (N_9087,N_7623,N_7506);
or U9088 (N_9088,N_8514,N_7598);
nand U9089 (N_9089,N_8881,N_8233);
and U9090 (N_9090,N_7636,N_7770);
xnor U9091 (N_9091,N_7775,N_8235);
nor U9092 (N_9092,N_8474,N_8339);
nor U9093 (N_9093,N_8761,N_8638);
nor U9094 (N_9094,N_8802,N_7854);
nor U9095 (N_9095,N_7824,N_8677);
nand U9096 (N_9096,N_8732,N_8334);
xor U9097 (N_9097,N_8620,N_7679);
or U9098 (N_9098,N_8014,N_8265);
nand U9099 (N_9099,N_7834,N_7646);
nand U9100 (N_9100,N_8133,N_7984);
and U9101 (N_9101,N_8548,N_7906);
or U9102 (N_9102,N_8231,N_8806);
nor U9103 (N_9103,N_8714,N_7952);
or U9104 (N_9104,N_7669,N_8783);
or U9105 (N_9105,N_7557,N_7698);
nor U9106 (N_9106,N_8791,N_8617);
xnor U9107 (N_9107,N_8427,N_8511);
and U9108 (N_9108,N_8756,N_7938);
and U9109 (N_9109,N_8553,N_8573);
or U9110 (N_9110,N_8490,N_7625);
and U9111 (N_9111,N_7986,N_8729);
and U9112 (N_9112,N_8793,N_8568);
nor U9113 (N_9113,N_7527,N_7655);
xor U9114 (N_9114,N_8629,N_8922);
nor U9115 (N_9115,N_8393,N_7617);
nand U9116 (N_9116,N_7560,N_8533);
and U9117 (N_9117,N_8285,N_8588);
or U9118 (N_9118,N_8652,N_8809);
nor U9119 (N_9119,N_8613,N_8811);
nor U9120 (N_9120,N_8104,N_7516);
nand U9121 (N_9121,N_8430,N_8015);
xnor U9122 (N_9122,N_8475,N_8593);
and U9123 (N_9123,N_8434,N_7559);
xor U9124 (N_9124,N_8209,N_7836);
xnor U9125 (N_9125,N_8162,N_8414);
nor U9126 (N_9126,N_8085,N_8109);
nand U9127 (N_9127,N_8834,N_7933);
nor U9128 (N_9128,N_7830,N_8346);
nand U9129 (N_9129,N_8905,N_7597);
and U9130 (N_9130,N_7609,N_8940);
nor U9131 (N_9131,N_8525,N_8604);
and U9132 (N_9132,N_8999,N_8679);
xor U9133 (N_9133,N_7767,N_8088);
nand U9134 (N_9134,N_8945,N_8497);
and U9135 (N_9135,N_7614,N_8606);
nand U9136 (N_9136,N_8320,N_7556);
nand U9137 (N_9137,N_8245,N_7853);
nor U9138 (N_9138,N_8073,N_7537);
nand U9139 (N_9139,N_8520,N_7758);
nor U9140 (N_9140,N_7962,N_8358);
or U9141 (N_9141,N_8372,N_8993);
nand U9142 (N_9142,N_8111,N_7501);
nand U9143 (N_9143,N_8931,N_7842);
or U9144 (N_9144,N_7878,N_8832);
xor U9145 (N_9145,N_8627,N_8754);
nor U9146 (N_9146,N_7575,N_8730);
nand U9147 (N_9147,N_8521,N_8687);
and U9148 (N_9148,N_8555,N_8824);
or U9149 (N_9149,N_7774,N_8305);
xnor U9150 (N_9150,N_8966,N_7533);
xnor U9151 (N_9151,N_8685,N_8830);
nand U9152 (N_9152,N_7893,N_8842);
and U9153 (N_9153,N_7961,N_8928);
or U9154 (N_9154,N_8155,N_8326);
and U9155 (N_9155,N_7534,N_7549);
or U9156 (N_9156,N_8818,N_8869);
or U9157 (N_9157,N_7925,N_8113);
or U9158 (N_9158,N_8787,N_8904);
nor U9159 (N_9159,N_8665,N_8924);
nand U9160 (N_9160,N_7876,N_8976);
and U9161 (N_9161,N_8420,N_8186);
and U9162 (N_9162,N_8926,N_7599);
and U9163 (N_9163,N_8951,N_7781);
xor U9164 (N_9164,N_8552,N_7502);
nand U9165 (N_9165,N_7838,N_8664);
and U9166 (N_9166,N_8856,N_7905);
and U9167 (N_9167,N_8433,N_7696);
and U9168 (N_9168,N_8805,N_8188);
and U9169 (N_9169,N_8397,N_8039);
xor U9170 (N_9170,N_7935,N_8402);
and U9171 (N_9171,N_8293,N_8254);
or U9172 (N_9172,N_8585,N_8075);
nor U9173 (N_9173,N_8239,N_8322);
nor U9174 (N_9174,N_8263,N_7845);
xnor U9175 (N_9175,N_8051,N_8328);
nand U9176 (N_9176,N_7685,N_8369);
and U9177 (N_9177,N_8772,N_7511);
xor U9178 (N_9178,N_8643,N_8646);
xor U9179 (N_9179,N_8789,N_8163);
or U9180 (N_9180,N_8973,N_7708);
and U9181 (N_9181,N_8963,N_8353);
and U9182 (N_9182,N_8579,N_8974);
and U9183 (N_9183,N_8063,N_8735);
xor U9184 (N_9184,N_7688,N_7923);
xor U9185 (N_9185,N_8991,N_8962);
xnor U9186 (N_9186,N_8534,N_8598);
xor U9187 (N_9187,N_8650,N_8894);
nor U9188 (N_9188,N_8211,N_8117);
or U9189 (N_9189,N_7541,N_8639);
and U9190 (N_9190,N_8062,N_7610);
nand U9191 (N_9191,N_8508,N_8539);
and U9192 (N_9192,N_8149,N_8990);
nand U9193 (N_9193,N_8589,N_8790);
and U9194 (N_9194,N_8868,N_8171);
and U9195 (N_9195,N_7880,N_8054);
xor U9196 (N_9196,N_7968,N_8703);
nand U9197 (N_9197,N_8129,N_8906);
and U9198 (N_9198,N_7783,N_8503);
nor U9199 (N_9199,N_7668,N_8934);
nand U9200 (N_9200,N_7785,N_8726);
and U9201 (N_9201,N_8406,N_7572);
and U9202 (N_9202,N_8029,N_7677);
nand U9203 (N_9203,N_7819,N_7722);
nand U9204 (N_9204,N_8174,N_8220);
nor U9205 (N_9205,N_8847,N_8795);
nand U9206 (N_9206,N_8377,N_8878);
nand U9207 (N_9207,N_7920,N_8828);
nand U9208 (N_9208,N_8008,N_7795);
nand U9209 (N_9209,N_8777,N_8865);
nand U9210 (N_9210,N_8505,N_8032);
and U9211 (N_9211,N_8574,N_7822);
nand U9212 (N_9212,N_8202,N_7500);
nor U9213 (N_9213,N_7828,N_7727);
and U9214 (N_9214,N_8307,N_8764);
nand U9215 (N_9215,N_8676,N_8561);
nand U9216 (N_9216,N_8693,N_7869);
and U9217 (N_9217,N_8038,N_8979);
xnor U9218 (N_9218,N_8241,N_7631);
nor U9219 (N_9219,N_7659,N_8482);
or U9220 (N_9220,N_8686,N_8127);
and U9221 (N_9221,N_7981,N_8031);
nand U9222 (N_9222,N_7664,N_8558);
nor U9223 (N_9223,N_8647,N_8464);
and U9224 (N_9224,N_7595,N_8443);
nor U9225 (N_9225,N_7912,N_7526);
nor U9226 (N_9226,N_7994,N_8296);
or U9227 (N_9227,N_8670,N_7874);
xnor U9228 (N_9228,N_8440,N_8769);
xor U9229 (N_9229,N_8086,N_8700);
nor U9230 (N_9230,N_8902,N_8289);
nand U9231 (N_9231,N_8242,N_8150);
or U9232 (N_9232,N_8094,N_8341);
or U9233 (N_9233,N_7521,N_7922);
nand U9234 (N_9234,N_7579,N_8323);
xor U9235 (N_9235,N_8669,N_8701);
or U9236 (N_9236,N_7972,N_7678);
xor U9237 (N_9237,N_8874,N_8959);
and U9238 (N_9238,N_8416,N_7800);
and U9239 (N_9239,N_8718,N_8897);
or U9240 (N_9240,N_7613,N_7691);
nand U9241 (N_9241,N_8064,N_8067);
nor U9242 (N_9242,N_8578,N_8141);
xor U9243 (N_9243,N_8500,N_7886);
nor U9244 (N_9244,N_8089,N_7666);
or U9245 (N_9245,N_8237,N_8501);
and U9246 (N_9246,N_7723,N_8043);
and U9247 (N_9247,N_8815,N_8238);
nor U9248 (N_9248,N_7960,N_8858);
xnor U9249 (N_9249,N_7776,N_8340);
nor U9250 (N_9250,N_8978,N_8742);
nor U9251 (N_9251,N_8849,N_7799);
and U9252 (N_9252,N_8596,N_8033);
or U9253 (N_9253,N_8223,N_8564);
nor U9254 (N_9254,N_8052,N_8139);
nand U9255 (N_9255,N_8213,N_7630);
and U9256 (N_9256,N_8609,N_8078);
nor U9257 (N_9257,N_8895,N_7635);
xor U9258 (N_9258,N_7763,N_7820);
or U9259 (N_9259,N_8813,N_8425);
and U9260 (N_9260,N_8401,N_8800);
nor U9261 (N_9261,N_8445,N_7772);
nor U9262 (N_9262,N_7946,N_8513);
or U9263 (N_9263,N_8386,N_8485);
nand U9264 (N_9264,N_8364,N_8690);
nor U9265 (N_9265,N_7538,N_8193);
xnor U9266 (N_9266,N_8295,N_8424);
xnor U9267 (N_9267,N_8634,N_8587);
or U9268 (N_9268,N_7643,N_8747);
nand U9269 (N_9269,N_8626,N_7529);
or U9270 (N_9270,N_7990,N_8496);
nand U9271 (N_9271,N_8177,N_8350);
or U9272 (N_9272,N_8255,N_7779);
nand U9273 (N_9273,N_7588,N_8217);
nor U9274 (N_9274,N_7736,N_7971);
nand U9275 (N_9275,N_8359,N_7596);
nand U9276 (N_9276,N_8477,N_8215);
nand U9277 (N_9277,N_8739,N_8913);
nor U9278 (N_9278,N_7832,N_8731);
nor U9279 (N_9279,N_8884,N_8442);
or U9280 (N_9280,N_8290,N_7647);
nand U9281 (N_9281,N_7699,N_8891);
nor U9282 (N_9282,N_7642,N_8218);
xor U9283 (N_9283,N_8232,N_7985);
xnor U9284 (N_9284,N_8835,N_7528);
or U9285 (N_9285,N_8699,N_7782);
xnor U9286 (N_9286,N_8337,N_7882);
nand U9287 (N_9287,N_7551,N_8506);
nor U9288 (N_9288,N_7903,N_7901);
nand U9289 (N_9289,N_8180,N_7827);
nand U9290 (N_9290,N_7868,N_8706);
nor U9291 (N_9291,N_8541,N_8097);
xor U9292 (N_9292,N_8674,N_8392);
nand U9293 (N_9293,N_8743,N_8026);
nand U9294 (N_9294,N_8631,N_8348);
nor U9295 (N_9295,N_8361,N_7732);
and U9296 (N_9296,N_7980,N_8240);
xnor U9297 (N_9297,N_7860,N_8059);
or U9298 (N_9298,N_8321,N_8275);
or U9299 (N_9299,N_7540,N_7835);
xor U9300 (N_9300,N_8493,N_7519);
and U9301 (N_9301,N_7843,N_8786);
nand U9302 (N_9302,N_7752,N_8551);
nand U9303 (N_9303,N_7620,N_8126);
nor U9304 (N_9304,N_7520,N_7590);
nor U9305 (N_9305,N_8538,N_8417);
nor U9306 (N_9306,N_8096,N_7826);
nor U9307 (N_9307,N_8352,N_8444);
nor U9308 (N_9308,N_8583,N_8258);
xnor U9309 (N_9309,N_8354,N_8074);
nand U9310 (N_9310,N_8331,N_8741);
and U9311 (N_9311,N_7746,N_7881);
or U9312 (N_9312,N_8013,N_7536);
or U9313 (N_9313,N_8035,N_7861);
nor U9314 (N_9314,N_8093,N_7592);
nand U9315 (N_9315,N_8695,N_8855);
xor U9316 (N_9316,N_7858,N_8374);
or U9317 (N_9317,N_7773,N_7694);
nand U9318 (N_9318,N_8975,N_7802);
or U9319 (N_9319,N_8582,N_8873);
nand U9320 (N_9320,N_8715,N_8812);
nand U9321 (N_9321,N_8079,N_7703);
or U9322 (N_9322,N_8300,N_7750);
nor U9323 (N_9323,N_8770,N_7851);
and U9324 (N_9324,N_8886,N_8995);
nor U9325 (N_9325,N_8208,N_8261);
or U9326 (N_9326,N_8264,N_8370);
nor U9327 (N_9327,N_7711,N_8484);
nand U9328 (N_9328,N_8137,N_7717);
nand U9329 (N_9329,N_8622,N_7726);
nand U9330 (N_9330,N_7945,N_8489);
nor U9331 (N_9331,N_7966,N_7576);
nand U9332 (N_9332,N_8776,N_7734);
nor U9333 (N_9333,N_8458,N_7747);
xnor U9334 (N_9334,N_8145,N_8624);
nor U9335 (N_9335,N_7619,N_8068);
nand U9336 (N_9336,N_8970,N_8021);
nor U9337 (N_9337,N_8119,N_8537);
and U9338 (N_9338,N_8138,N_7766);
and U9339 (N_9339,N_7909,N_8825);
nand U9340 (N_9340,N_7715,N_8204);
and U9341 (N_9341,N_8376,N_8597);
nor U9342 (N_9342,N_7856,N_8001);
or U9343 (N_9343,N_7992,N_8382);
or U9344 (N_9344,N_7515,N_8843);
or U9345 (N_9345,N_7639,N_7801);
nor U9346 (N_9346,N_7967,N_8413);
or U9347 (N_9347,N_8755,N_7875);
xor U9348 (N_9348,N_8708,N_8170);
xnor U9349 (N_9349,N_7554,N_8981);
or U9350 (N_9350,N_7917,N_7955);
nor U9351 (N_9351,N_8396,N_8228);
and U9352 (N_9352,N_8084,N_8892);
nand U9353 (N_9353,N_7672,N_8867);
xor U9354 (N_9354,N_8470,N_8814);
xnor U9355 (N_9355,N_8022,N_7505);
or U9356 (N_9356,N_8877,N_7661);
and U9357 (N_9357,N_7741,N_7825);
xor U9358 (N_9358,N_8398,N_8118);
nand U9359 (N_9359,N_8632,N_7810);
or U9360 (N_9360,N_8190,N_8125);
xor U9361 (N_9361,N_8378,N_8550);
nor U9362 (N_9362,N_7837,N_7887);
and U9363 (N_9363,N_7787,N_8532);
and U9364 (N_9364,N_8020,N_8441);
nor U9365 (N_9365,N_8965,N_7754);
or U9366 (N_9366,N_8559,N_8887);
or U9367 (N_9367,N_7908,N_8176);
nand U9368 (N_9368,N_8487,N_8851);
nand U9369 (N_9369,N_7751,N_7704);
or U9370 (N_9370,N_7977,N_7608);
nand U9371 (N_9371,N_8429,N_7740);
xnor U9372 (N_9372,N_7671,N_8581);
xor U9373 (N_9373,N_7927,N_8012);
nand U9374 (N_9374,N_8003,N_8941);
xor U9375 (N_9375,N_8488,N_8419);
or U9376 (N_9376,N_7545,N_7550);
or U9377 (N_9377,N_8908,N_8411);
xnor U9378 (N_9378,N_7720,N_7899);
or U9379 (N_9379,N_8826,N_7663);
and U9380 (N_9380,N_7916,N_8450);
and U9381 (N_9381,N_8112,N_8727);
and U9382 (N_9382,N_8019,N_8270);
nor U9383 (N_9383,N_7697,N_8980);
xnor U9384 (N_9384,N_7921,N_7583);
nand U9385 (N_9385,N_7870,N_8227);
or U9386 (N_9386,N_8437,N_8421);
and U9387 (N_9387,N_8697,N_8030);
xnor U9388 (N_9388,N_8036,N_8457);
and U9389 (N_9389,N_8316,N_7602);
nor U9390 (N_9390,N_8943,N_8509);
and U9391 (N_9391,N_8527,N_8821);
nand U9392 (N_9392,N_8324,N_8050);
nand U9393 (N_9393,N_7947,N_7546);
nor U9394 (N_9394,N_8775,N_7673);
nor U9395 (N_9395,N_8077,N_8862);
and U9396 (N_9396,N_8375,N_8345);
xnor U9397 (N_9397,N_8586,N_7806);
nand U9398 (N_9398,N_8649,N_8148);
and U9399 (N_9399,N_8724,N_7807);
nand U9400 (N_9400,N_8381,N_8658);
and U9401 (N_9401,N_8810,N_8956);
xnor U9402 (N_9402,N_8297,N_8455);
or U9403 (N_9403,N_8136,N_8308);
and U9404 (N_9404,N_8251,N_8753);
and U9405 (N_9405,N_8584,N_8594);
and U9406 (N_9406,N_7719,N_8932);
xor U9407 (N_9407,N_8335,N_8347);
xor U9408 (N_9408,N_7805,N_7798);
and U9409 (N_9409,N_8214,N_8183);
nor U9410 (N_9410,N_8845,N_8694);
and U9411 (N_9411,N_7731,N_8197);
xor U9412 (N_9412,N_8422,N_8034);
or U9413 (N_9413,N_7562,N_7919);
xnor U9414 (N_9414,N_8355,N_7518);
nand U9415 (N_9415,N_8577,N_7706);
and U9416 (N_9416,N_8723,N_7924);
nor U9417 (N_9417,N_8023,N_8901);
nand U9418 (N_9418,N_7937,N_8985);
or U9419 (N_9419,N_8403,N_8318);
and U9420 (N_9420,N_8746,N_8529);
or U9421 (N_9421,N_8462,N_8486);
nor U9422 (N_9422,N_8216,N_8563);
nor U9423 (N_9423,N_7512,N_7895);
or U9424 (N_9424,N_8545,N_8860);
nor U9425 (N_9425,N_8515,N_8576);
and U9426 (N_9426,N_8124,N_8668);
xnor U9427 (N_9427,N_7568,N_8092);
and U9428 (N_9428,N_8605,N_8385);
and U9429 (N_9429,N_7762,N_7716);
nand U9430 (N_9430,N_7821,N_8557);
or U9431 (N_9431,N_7891,N_8997);
or U9432 (N_9432,N_8744,N_8282);
or U9433 (N_9433,N_8817,N_8528);
or U9434 (N_9434,N_7648,N_8268);
nor U9435 (N_9435,N_8792,N_7897);
nor U9436 (N_9436,N_8049,N_8053);
and U9437 (N_9437,N_7794,N_8807);
nor U9438 (N_9438,N_8404,N_7667);
or U9439 (N_9439,N_8274,N_8410);
xor U9440 (N_9440,N_8121,N_8667);
or U9441 (N_9441,N_8671,N_7867);
or U9442 (N_9442,N_8841,N_7778);
and U9443 (N_9443,N_8566,N_8659);
nand U9444 (N_9444,N_7653,N_8160);
and U9445 (N_9445,N_8616,N_8749);
xor U9446 (N_9446,N_7654,N_8967);
and U9447 (N_9447,N_7936,N_8454);
xnor U9448 (N_9448,N_8750,N_7970);
nor U9449 (N_9449,N_8889,N_8954);
nand U9450 (N_9450,N_8095,N_7983);
xnor U9451 (N_9451,N_8291,N_7624);
xnor U9452 (N_9452,N_8949,N_8950);
nor U9453 (N_9453,N_8536,N_8154);
nand U9454 (N_9454,N_8143,N_7650);
xnor U9455 (N_9455,N_8516,N_7594);
nor U9456 (N_9456,N_7928,N_7633);
or U9457 (N_9457,N_8681,N_7973);
nor U9458 (N_9458,N_8716,N_8081);
xnor U9459 (N_9459,N_7713,N_7989);
nand U9460 (N_9460,N_8279,N_8142);
nor U9461 (N_9461,N_8611,N_8936);
nand U9462 (N_9462,N_7813,N_8483);
xnor U9463 (N_9463,N_8929,N_7675);
and U9464 (N_9464,N_8785,N_8994);
and U9465 (N_9465,N_8875,N_8702);
or U9466 (N_9466,N_7622,N_8580);
nor U9467 (N_9467,N_7616,N_8303);
nor U9468 (N_9468,N_8432,N_8249);
nor U9469 (N_9469,N_8651,N_8002);
nor U9470 (N_9470,N_8569,N_8134);
nand U9471 (N_9471,N_8682,N_7712);
and U9472 (N_9472,N_8182,N_8060);
and U9473 (N_9473,N_8848,N_8319);
or U9474 (N_9474,N_8327,N_7566);
or U9475 (N_9475,N_8927,N_8916);
or U9476 (N_9476,N_8083,N_8467);
or U9477 (N_9477,N_8854,N_8921);
and U9478 (N_9478,N_8618,N_8788);
or U9479 (N_9479,N_8846,N_8480);
or U9480 (N_9480,N_7883,N_8510);
nand U9481 (N_9481,N_7913,N_7904);
nor U9482 (N_9482,N_8736,N_8201);
xor U9483 (N_9483,N_7640,N_8115);
nor U9484 (N_9484,N_8801,N_7611);
and U9485 (N_9485,N_8923,N_8526);
or U9486 (N_9486,N_8384,N_8688);
nor U9487 (N_9487,N_8435,N_7581);
and U9488 (N_9488,N_7847,N_8098);
xor U9489 (N_9489,N_7605,N_8481);
xor U9490 (N_9490,N_8592,N_7657);
nor U9491 (N_9491,N_8301,N_7690);
nand U9492 (N_9492,N_7705,N_8925);
xnor U9493 (N_9493,N_7764,N_7755);
nor U9494 (N_9494,N_8234,N_8367);
xnor U9495 (N_9495,N_8773,N_7753);
or U9496 (N_9496,N_8893,N_8969);
nand U9497 (N_9497,N_8879,N_7863);
or U9498 (N_9498,N_8017,N_7593);
nand U9499 (N_9499,N_8644,N_8710);
nand U9500 (N_9500,N_7840,N_7729);
nand U9501 (N_9501,N_8310,N_8989);
nor U9502 (N_9502,N_7601,N_8329);
or U9503 (N_9503,N_7714,N_8253);
nand U9504 (N_9504,N_8349,N_8819);
nand U9505 (N_9505,N_8011,N_7615);
nand U9506 (N_9506,N_8757,N_8070);
or U9507 (N_9507,N_7748,N_8090);
or U9508 (N_9508,N_8544,N_8332);
and U9509 (N_9509,N_8418,N_8946);
nor U9510 (N_9510,N_7780,N_8368);
nor U9511 (N_9511,N_8436,N_8317);
and U9512 (N_9512,N_7577,N_8451);
or U9513 (N_9513,N_8273,N_8257);
xnor U9514 (N_9514,N_8311,N_8836);
or U9515 (N_9515,N_8494,N_8448);
or U9516 (N_9516,N_8625,N_7890);
nand U9517 (N_9517,N_7896,N_8968);
xor U9518 (N_9518,N_8720,N_8161);
or U9519 (N_9519,N_7982,N_8502);
or U9520 (N_9520,N_7949,N_7724);
xor U9521 (N_9521,N_8276,N_8734);
and U9522 (N_9522,N_8178,N_8010);
and U9523 (N_9523,N_8123,N_8379);
xnor U9524 (N_9524,N_8745,N_7884);
nand U9525 (N_9525,N_8888,N_8567);
and U9526 (N_9526,N_8206,N_7814);
nand U9527 (N_9527,N_8542,N_8356);
and U9528 (N_9528,N_8939,N_8152);
nand U9529 (N_9529,N_7809,N_8391);
nor U9530 (N_9530,N_7585,N_8663);
and U9531 (N_9531,N_8140,N_8779);
and U9532 (N_9532,N_7833,N_8495);
nor U9533 (N_9533,N_7569,N_8000);
and U9534 (N_9534,N_8116,N_7790);
xnor U9535 (N_9535,N_8907,N_8837);
or U9536 (N_9536,N_7939,N_7841);
and U9537 (N_9537,N_8930,N_8602);
nor U9538 (N_9538,N_8759,N_8225);
nand U9539 (N_9539,N_7877,N_7811);
and U9540 (N_9540,N_8944,N_8595);
and U9541 (N_9541,N_7975,N_7808);
or U9542 (N_9542,N_8048,N_8105);
and U9543 (N_9543,N_7743,N_8314);
nand U9544 (N_9544,N_8863,N_8796);
nand U9545 (N_9545,N_7689,N_8523);
nor U9546 (N_9546,N_8299,N_8640);
nand U9547 (N_9547,N_7700,N_8748);
and U9548 (N_9548,N_8292,N_7777);
or U9549 (N_9549,N_8492,N_8222);
and U9550 (N_9550,N_8040,N_8342);
xnor U9551 (N_9551,N_7730,N_8740);
nor U9552 (N_9552,N_8996,N_8857);
and U9553 (N_9553,N_8415,N_8172);
or U9554 (N_9554,N_7812,N_8132);
xnor U9555 (N_9555,N_7603,N_8256);
xnor U9556 (N_9556,N_8728,N_8645);
xnor U9557 (N_9557,N_8343,N_7530);
nand U9558 (N_9558,N_8230,N_8167);
xor U9559 (N_9559,N_8272,N_7817);
xor U9560 (N_9560,N_8351,N_8535);
and U9561 (N_9561,N_7523,N_8883);
and U9562 (N_9562,N_8983,N_8683);
nor U9563 (N_9563,N_7995,N_8298);
or U9564 (N_9564,N_8082,N_8271);
nand U9565 (N_9565,N_7931,N_8909);
or U9566 (N_9566,N_8191,N_8405);
and U9567 (N_9567,N_8135,N_8546);
xor U9568 (N_9568,N_7944,N_7662);
and U9569 (N_9569,N_8524,N_7934);
nor U9570 (N_9570,N_8961,N_8866);
or U9571 (N_9571,N_7760,N_7976);
xnor U9572 (N_9572,N_8309,N_8266);
nor U9573 (N_9573,N_8365,N_7797);
nor U9574 (N_9574,N_8277,N_8512);
xor U9575 (N_9575,N_8478,N_8189);
or U9576 (N_9576,N_8360,N_8590);
nor U9577 (N_9577,N_7692,N_7641);
and U9578 (N_9578,N_8147,N_8760);
xnor U9579 (N_9579,N_8110,N_8173);
nor U9580 (N_9580,N_8153,N_8614);
nand U9581 (N_9581,N_8864,N_8948);
nand U9582 (N_9582,N_8621,N_8100);
nor U9583 (N_9583,N_8246,N_8556);
nor U9584 (N_9584,N_8704,N_8600);
or U9585 (N_9585,N_7645,N_7957);
or U9586 (N_9586,N_7660,N_7993);
nand U9587 (N_9587,N_8072,N_8660);
and U9588 (N_9588,N_8472,N_8517);
or U9589 (N_9589,N_7768,N_7829);
and U9590 (N_9590,N_8207,N_8986);
nand U9591 (N_9591,N_7815,N_7910);
nor U9592 (N_9592,N_8984,N_8453);
xnor U9593 (N_9593,N_8428,N_8633);
and U9594 (N_9594,N_7503,N_8371);
and U9595 (N_9595,N_8325,N_7513);
or U9596 (N_9596,N_8388,N_8338);
nor U9597 (N_9597,N_7872,N_8840);
nand U9598 (N_9598,N_7759,N_8827);
and U9599 (N_9599,N_7658,N_8900);
or U9600 (N_9600,N_7852,N_7999);
nand U9601 (N_9601,N_8707,N_8200);
or U9602 (N_9602,N_7606,N_8169);
xor U9603 (N_9603,N_8400,N_8852);
nand U9604 (N_9604,N_8733,N_7563);
or U9605 (N_9605,N_8007,N_8880);
nor U9606 (N_9606,N_7737,N_7629);
xnor U9607 (N_9607,N_8224,N_8540);
xor U9608 (N_9608,N_8988,N_8607);
or U9609 (N_9609,N_8306,N_8247);
nor U9610 (N_9610,N_7892,N_8992);
and U9611 (N_9611,N_7510,N_8461);
xor U9612 (N_9612,N_8128,N_7988);
and U9613 (N_9613,N_7792,N_8833);
or U9614 (N_9614,N_7948,N_8158);
or U9615 (N_9615,N_8914,N_8184);
nand U9616 (N_9616,N_8637,N_8782);
nand U9617 (N_9617,N_7634,N_8491);
and U9618 (N_9618,N_8168,N_8226);
xor U9619 (N_9619,N_8850,N_8175);
nand U9620 (N_9620,N_8853,N_8937);
nand U9621 (N_9621,N_8971,N_8447);
xor U9622 (N_9622,N_8767,N_8648);
nor U9623 (N_9623,N_8562,N_8661);
xor U9624 (N_9624,N_8766,N_7525);
nand U9625 (N_9625,N_8942,N_7745);
xnor U9626 (N_9626,N_8047,N_8219);
and U9627 (N_9627,N_8198,N_8252);
and U9628 (N_9628,N_8565,N_8964);
or U9629 (N_9629,N_8570,N_8426);
nand U9630 (N_9630,N_8006,N_8717);
or U9631 (N_9631,N_8870,N_7739);
nand U9632 (N_9632,N_7507,N_7757);
nand U9633 (N_9633,N_7940,N_7735);
xor U9634 (N_9634,N_7552,N_8431);
nor U9635 (N_9635,N_7978,N_7586);
nand U9636 (N_9636,N_8861,N_7632);
or U9637 (N_9637,N_7570,N_8890);
nand U9638 (N_9638,N_8678,N_8056);
nand U9639 (N_9639,N_8911,N_8283);
or U9640 (N_9640,N_7670,N_8456);
nor U9641 (N_9641,N_8820,N_8076);
or U9642 (N_9642,N_8199,N_8196);
or U9643 (N_9643,N_7907,N_8610);
nand U9644 (N_9644,N_8711,N_8919);
xor U9645 (N_9645,N_7786,N_8987);
and U9646 (N_9646,N_7709,N_8045);
nor U9647 (N_9647,N_8302,N_7871);
or U9648 (N_9648,N_7580,N_7710);
nand U9649 (N_9649,N_7589,N_7964);
nor U9650 (N_9650,N_7864,N_8666);
or U9651 (N_9651,N_7959,N_7626);
nand U9652 (N_9652,N_7894,N_7818);
xor U9653 (N_9653,N_7958,N_8762);
xor U9654 (N_9654,N_8960,N_8037);
and U9655 (N_9655,N_7951,N_8476);
and U9656 (N_9656,N_7644,N_7718);
or U9657 (N_9657,N_7844,N_8498);
and U9658 (N_9658,N_8560,N_8091);
xor U9659 (N_9659,N_7539,N_8955);
nand U9660 (N_9660,N_8195,N_7652);
or U9661 (N_9661,N_8933,N_8408);
or U9662 (N_9662,N_8635,N_8719);
or U9663 (N_9663,N_8662,N_8713);
nand U9664 (N_9664,N_7862,N_8473);
nor U9665 (N_9665,N_8912,N_7544);
or U9666 (N_9666,N_7548,N_7567);
nor U9667 (N_9667,N_8816,N_8780);
xnor U9668 (N_9668,N_8099,N_7918);
and U9669 (N_9669,N_7543,N_7926);
nor U9670 (N_9670,N_8439,N_7997);
nand U9671 (N_9671,N_8982,N_8896);
and U9672 (N_9672,N_8144,N_8831);
nor U9673 (N_9673,N_7956,N_8920);
nor U9674 (N_9674,N_7571,N_8623);
nand U9675 (N_9675,N_7930,N_8705);
and U9676 (N_9676,N_8057,N_8469);
or U9677 (N_9677,N_8058,N_7885);
and U9678 (N_9678,N_8409,N_8952);
or U9679 (N_9679,N_7788,N_8380);
nand U9680 (N_9680,N_8009,N_8210);
or U9681 (N_9681,N_8885,N_7649);
or U9682 (N_9682,N_8466,N_8164);
or U9683 (N_9683,N_8107,N_8575);
xnor U9684 (N_9684,N_7771,N_8642);
or U9685 (N_9685,N_7756,N_8269);
nor U9686 (N_9686,N_7591,N_8055);
or U9687 (N_9687,N_8630,N_7804);
and U9688 (N_9688,N_8543,N_8696);
nand U9689 (N_9689,N_8181,N_7582);
nand U9690 (N_9690,N_8446,N_8518);
or U9691 (N_9691,N_8692,N_8267);
or U9692 (N_9692,N_8278,N_8286);
nand U9693 (N_9693,N_7665,N_8774);
xor U9694 (N_9694,N_7911,N_8205);
nor U9695 (N_9695,N_8691,N_8722);
nor U9696 (N_9696,N_8390,N_8876);
nor U9697 (N_9697,N_8712,N_8108);
nor U9698 (N_9698,N_8531,N_8080);
and U9699 (N_9699,N_7744,N_8042);
or U9700 (N_9700,N_8102,N_7929);
or U9701 (N_9701,N_8383,N_7839);
nor U9702 (N_9702,N_7742,N_8471);
nand U9703 (N_9703,N_8259,N_8027);
nor U9704 (N_9704,N_8684,N_7979);
xnor U9705 (N_9705,N_8737,N_8025);
nor U9706 (N_9706,N_8479,N_8028);
xnor U9707 (N_9707,N_7693,N_7849);
and U9708 (N_9708,N_8165,N_8829);
and U9709 (N_9709,N_8066,N_8159);
nor U9710 (N_9710,N_8947,N_8641);
or U9711 (N_9711,N_8407,N_7674);
nand U9712 (N_9712,N_7683,N_7789);
xor U9713 (N_9713,N_8672,N_8721);
nand U9714 (N_9714,N_8808,N_7749);
nand U9715 (N_9715,N_8004,N_8203);
nor U9716 (N_9716,N_8362,N_8499);
or U9717 (N_9717,N_7509,N_7769);
or U9718 (N_9718,N_8288,N_8005);
and U9719 (N_9719,N_8778,N_8061);
xnor U9720 (N_9720,N_8872,N_8758);
or U9721 (N_9721,N_7508,N_8522);
or U9722 (N_9722,N_7796,N_8903);
xnor U9723 (N_9723,N_8330,N_7728);
nand U9724 (N_9724,N_8103,N_8438);
nor U9725 (N_9725,N_8917,N_8673);
xnor U9726 (N_9726,N_8656,N_7686);
xor U9727 (N_9727,N_8771,N_7765);
nand U9728 (N_9728,N_8373,N_8281);
nor U9729 (N_9729,N_7574,N_8675);
or U9730 (N_9730,N_8507,N_8262);
nand U9731 (N_9731,N_7865,N_7656);
or U9732 (N_9732,N_8069,N_8336);
or U9733 (N_9733,N_8530,N_8179);
nor U9734 (N_9734,N_8166,N_8459);
xnor U9735 (N_9735,N_8998,N_7618);
nor U9736 (N_9736,N_8468,N_7621);
and U9737 (N_9737,N_8449,N_7584);
and U9738 (N_9738,N_7531,N_7953);
nand U9739 (N_9739,N_8709,N_7857);
or U9740 (N_9740,N_8615,N_8823);
nor U9741 (N_9741,N_7707,N_8024);
and U9742 (N_9742,N_7682,N_7866);
and U9743 (N_9743,N_8280,N_8504);
nand U9744 (N_9744,N_7873,N_8394);
nand U9745 (N_9745,N_7721,N_7535);
nand U9746 (N_9746,N_8958,N_7684);
and U9747 (N_9747,N_8087,N_8619);
or U9748 (N_9748,N_7900,N_7950);
nand U9749 (N_9749,N_7695,N_8260);
xor U9750 (N_9750,N_8038,N_8663);
nand U9751 (N_9751,N_8860,N_8032);
and U9752 (N_9752,N_8623,N_7924);
nand U9753 (N_9753,N_8277,N_8495);
nand U9754 (N_9754,N_8504,N_7695);
nor U9755 (N_9755,N_8984,N_8351);
xnor U9756 (N_9756,N_7836,N_7960);
xnor U9757 (N_9757,N_8718,N_8208);
xor U9758 (N_9758,N_8085,N_7928);
xor U9759 (N_9759,N_7722,N_8940);
or U9760 (N_9760,N_7545,N_8728);
and U9761 (N_9761,N_7514,N_8757);
nor U9762 (N_9762,N_8167,N_8229);
nand U9763 (N_9763,N_8422,N_8081);
and U9764 (N_9764,N_7809,N_8929);
or U9765 (N_9765,N_8795,N_8529);
or U9766 (N_9766,N_7768,N_8593);
or U9767 (N_9767,N_8093,N_8806);
nand U9768 (N_9768,N_7779,N_7950);
nand U9769 (N_9769,N_8988,N_8484);
xnor U9770 (N_9770,N_7852,N_8063);
xor U9771 (N_9771,N_8857,N_7507);
or U9772 (N_9772,N_7552,N_8287);
and U9773 (N_9773,N_7868,N_8812);
xor U9774 (N_9774,N_8269,N_7840);
nor U9775 (N_9775,N_7586,N_8662);
nor U9776 (N_9776,N_8312,N_7737);
xor U9777 (N_9777,N_7750,N_8565);
or U9778 (N_9778,N_8679,N_8968);
xor U9779 (N_9779,N_8177,N_7517);
nor U9780 (N_9780,N_8190,N_8031);
xnor U9781 (N_9781,N_7626,N_7732);
and U9782 (N_9782,N_8088,N_7924);
nor U9783 (N_9783,N_8003,N_8367);
nor U9784 (N_9784,N_8426,N_8549);
nand U9785 (N_9785,N_8108,N_8121);
or U9786 (N_9786,N_8353,N_7934);
and U9787 (N_9787,N_8444,N_8671);
or U9788 (N_9788,N_8598,N_8149);
nand U9789 (N_9789,N_7958,N_7705);
and U9790 (N_9790,N_8177,N_7566);
or U9791 (N_9791,N_8863,N_7536);
or U9792 (N_9792,N_8536,N_8449);
or U9793 (N_9793,N_8346,N_8772);
nor U9794 (N_9794,N_7558,N_7890);
xor U9795 (N_9795,N_7989,N_8457);
xor U9796 (N_9796,N_8920,N_8805);
or U9797 (N_9797,N_8837,N_8645);
nand U9798 (N_9798,N_7747,N_8966);
and U9799 (N_9799,N_7801,N_8531);
nor U9800 (N_9800,N_8134,N_8726);
nand U9801 (N_9801,N_8234,N_8920);
xor U9802 (N_9802,N_7659,N_8414);
nand U9803 (N_9803,N_8545,N_7632);
or U9804 (N_9804,N_8235,N_7620);
nand U9805 (N_9805,N_7700,N_8099);
nand U9806 (N_9806,N_8079,N_8464);
nand U9807 (N_9807,N_7863,N_8771);
or U9808 (N_9808,N_8866,N_8501);
xnor U9809 (N_9809,N_8135,N_8729);
nand U9810 (N_9810,N_7638,N_8341);
nand U9811 (N_9811,N_8193,N_8435);
nand U9812 (N_9812,N_8766,N_7813);
or U9813 (N_9813,N_8877,N_7830);
nor U9814 (N_9814,N_7981,N_8534);
or U9815 (N_9815,N_7959,N_7537);
or U9816 (N_9816,N_7521,N_8263);
nand U9817 (N_9817,N_8523,N_7754);
and U9818 (N_9818,N_8793,N_8885);
or U9819 (N_9819,N_7767,N_7650);
xnor U9820 (N_9820,N_8774,N_8402);
nand U9821 (N_9821,N_8328,N_7809);
xnor U9822 (N_9822,N_7772,N_7578);
and U9823 (N_9823,N_8380,N_8116);
or U9824 (N_9824,N_8069,N_7791);
xnor U9825 (N_9825,N_8856,N_8629);
and U9826 (N_9826,N_8187,N_8777);
xnor U9827 (N_9827,N_8097,N_8506);
and U9828 (N_9828,N_8209,N_8983);
nand U9829 (N_9829,N_8929,N_8383);
or U9830 (N_9830,N_8208,N_8950);
nor U9831 (N_9831,N_8918,N_7661);
or U9832 (N_9832,N_8504,N_8082);
or U9833 (N_9833,N_8426,N_7998);
nor U9834 (N_9834,N_7532,N_8152);
xnor U9835 (N_9835,N_7958,N_7538);
nand U9836 (N_9836,N_7765,N_8388);
xnor U9837 (N_9837,N_8343,N_8619);
nor U9838 (N_9838,N_7632,N_8324);
xnor U9839 (N_9839,N_8962,N_7922);
and U9840 (N_9840,N_8849,N_7508);
nand U9841 (N_9841,N_8653,N_8230);
nor U9842 (N_9842,N_8023,N_8575);
xor U9843 (N_9843,N_7750,N_8433);
xnor U9844 (N_9844,N_8260,N_8148);
and U9845 (N_9845,N_7834,N_8043);
nor U9846 (N_9846,N_7844,N_7679);
or U9847 (N_9847,N_8021,N_8532);
nand U9848 (N_9848,N_7529,N_7609);
nand U9849 (N_9849,N_7722,N_8207);
or U9850 (N_9850,N_7530,N_7646);
nor U9851 (N_9851,N_8973,N_7838);
nor U9852 (N_9852,N_8965,N_8969);
nor U9853 (N_9853,N_8328,N_8985);
and U9854 (N_9854,N_8330,N_7535);
xnor U9855 (N_9855,N_7920,N_8140);
or U9856 (N_9856,N_7704,N_8460);
and U9857 (N_9857,N_8329,N_7910);
xor U9858 (N_9858,N_8739,N_7695);
xor U9859 (N_9859,N_8756,N_7683);
nor U9860 (N_9860,N_8768,N_7553);
nor U9861 (N_9861,N_8581,N_8798);
xor U9862 (N_9862,N_8692,N_8392);
xnor U9863 (N_9863,N_7515,N_8478);
and U9864 (N_9864,N_8019,N_8087);
or U9865 (N_9865,N_8148,N_8129);
nor U9866 (N_9866,N_8949,N_8934);
xor U9867 (N_9867,N_8579,N_8371);
and U9868 (N_9868,N_7926,N_7713);
or U9869 (N_9869,N_7660,N_7572);
and U9870 (N_9870,N_8501,N_8275);
and U9871 (N_9871,N_7677,N_7780);
xor U9872 (N_9872,N_8354,N_8952);
and U9873 (N_9873,N_8644,N_7850);
and U9874 (N_9874,N_8918,N_7707);
nor U9875 (N_9875,N_8214,N_8587);
nand U9876 (N_9876,N_7519,N_7611);
or U9877 (N_9877,N_8176,N_7770);
or U9878 (N_9878,N_8301,N_8370);
nand U9879 (N_9879,N_7632,N_8633);
nand U9880 (N_9880,N_8543,N_7643);
xor U9881 (N_9881,N_7678,N_7851);
and U9882 (N_9882,N_8148,N_7728);
or U9883 (N_9883,N_8915,N_7776);
and U9884 (N_9884,N_7545,N_7743);
or U9885 (N_9885,N_7602,N_7581);
nor U9886 (N_9886,N_8693,N_7570);
nor U9887 (N_9887,N_7975,N_8096);
or U9888 (N_9888,N_7897,N_8875);
or U9889 (N_9889,N_7596,N_8062);
and U9890 (N_9890,N_8207,N_8364);
or U9891 (N_9891,N_7687,N_7574);
or U9892 (N_9892,N_8883,N_7628);
and U9893 (N_9893,N_7641,N_7652);
and U9894 (N_9894,N_8911,N_8720);
nand U9895 (N_9895,N_8663,N_8305);
xor U9896 (N_9896,N_7560,N_7648);
xor U9897 (N_9897,N_7841,N_7621);
nand U9898 (N_9898,N_8513,N_8700);
or U9899 (N_9899,N_8294,N_8908);
xor U9900 (N_9900,N_8662,N_8010);
or U9901 (N_9901,N_7956,N_7569);
nor U9902 (N_9902,N_8113,N_8988);
nor U9903 (N_9903,N_7984,N_8778);
and U9904 (N_9904,N_8289,N_8530);
and U9905 (N_9905,N_7526,N_7929);
or U9906 (N_9906,N_8163,N_7636);
nor U9907 (N_9907,N_8782,N_7987);
xnor U9908 (N_9908,N_8322,N_8705);
or U9909 (N_9909,N_8525,N_8893);
and U9910 (N_9910,N_7813,N_8856);
nand U9911 (N_9911,N_7513,N_8780);
nor U9912 (N_9912,N_7615,N_7600);
and U9913 (N_9913,N_8549,N_7868);
and U9914 (N_9914,N_8005,N_7861);
xnor U9915 (N_9915,N_8283,N_8186);
and U9916 (N_9916,N_8617,N_8857);
or U9917 (N_9917,N_8839,N_8021);
xnor U9918 (N_9918,N_8313,N_8620);
nor U9919 (N_9919,N_7644,N_8016);
or U9920 (N_9920,N_8515,N_7592);
nand U9921 (N_9921,N_7879,N_8484);
or U9922 (N_9922,N_8454,N_8068);
nor U9923 (N_9923,N_7723,N_8672);
and U9924 (N_9924,N_8897,N_8708);
xnor U9925 (N_9925,N_7681,N_8953);
xnor U9926 (N_9926,N_8539,N_7740);
or U9927 (N_9927,N_8562,N_8079);
nand U9928 (N_9928,N_8460,N_7700);
xor U9929 (N_9929,N_8514,N_8563);
xor U9930 (N_9930,N_8178,N_8850);
or U9931 (N_9931,N_7829,N_7620);
xor U9932 (N_9932,N_7515,N_8584);
nor U9933 (N_9933,N_8445,N_8000);
nand U9934 (N_9934,N_8024,N_8411);
nor U9935 (N_9935,N_8101,N_8561);
xnor U9936 (N_9936,N_8893,N_8828);
and U9937 (N_9937,N_8646,N_7601);
or U9938 (N_9938,N_7558,N_8169);
and U9939 (N_9939,N_7551,N_7744);
or U9940 (N_9940,N_8359,N_8819);
nor U9941 (N_9941,N_7994,N_8897);
nor U9942 (N_9942,N_8751,N_8982);
xnor U9943 (N_9943,N_7575,N_8944);
and U9944 (N_9944,N_7716,N_8121);
xnor U9945 (N_9945,N_7879,N_8052);
or U9946 (N_9946,N_8165,N_7985);
xnor U9947 (N_9947,N_8778,N_8707);
or U9948 (N_9948,N_8120,N_8198);
xor U9949 (N_9949,N_8059,N_8999);
or U9950 (N_9950,N_7704,N_8911);
and U9951 (N_9951,N_8800,N_8896);
or U9952 (N_9952,N_8530,N_8783);
or U9953 (N_9953,N_8780,N_7576);
and U9954 (N_9954,N_7920,N_8270);
nor U9955 (N_9955,N_7871,N_8665);
and U9956 (N_9956,N_7642,N_8010);
or U9957 (N_9957,N_8868,N_8264);
xor U9958 (N_9958,N_7677,N_8003);
xnor U9959 (N_9959,N_8598,N_8086);
and U9960 (N_9960,N_8367,N_8596);
and U9961 (N_9961,N_7932,N_8019);
xor U9962 (N_9962,N_7577,N_8539);
nor U9963 (N_9963,N_7985,N_8820);
nand U9964 (N_9964,N_8904,N_8484);
nand U9965 (N_9965,N_8698,N_8751);
xor U9966 (N_9966,N_8988,N_8852);
nor U9967 (N_9967,N_7913,N_8697);
nor U9968 (N_9968,N_8927,N_7542);
and U9969 (N_9969,N_8116,N_7802);
and U9970 (N_9970,N_8416,N_7501);
or U9971 (N_9971,N_8057,N_8163);
xnor U9972 (N_9972,N_8355,N_8459);
or U9973 (N_9973,N_7846,N_7681);
and U9974 (N_9974,N_7708,N_8518);
or U9975 (N_9975,N_8821,N_7799);
or U9976 (N_9976,N_8688,N_8037);
or U9977 (N_9977,N_8603,N_8936);
or U9978 (N_9978,N_8626,N_8697);
or U9979 (N_9979,N_7645,N_7593);
nor U9980 (N_9980,N_8427,N_8155);
xnor U9981 (N_9981,N_8825,N_8142);
or U9982 (N_9982,N_8643,N_7587);
xor U9983 (N_9983,N_8122,N_7973);
and U9984 (N_9984,N_8506,N_8187);
and U9985 (N_9985,N_8757,N_7991);
nor U9986 (N_9986,N_8091,N_8545);
nor U9987 (N_9987,N_8175,N_8184);
or U9988 (N_9988,N_8933,N_8512);
xor U9989 (N_9989,N_7755,N_8409);
nand U9990 (N_9990,N_7511,N_8325);
or U9991 (N_9991,N_8793,N_8388);
or U9992 (N_9992,N_8537,N_8987);
nand U9993 (N_9993,N_8968,N_7863);
xnor U9994 (N_9994,N_8999,N_8681);
or U9995 (N_9995,N_8052,N_8822);
nor U9996 (N_9996,N_7854,N_8262);
xnor U9997 (N_9997,N_8791,N_7956);
nand U9998 (N_9998,N_8390,N_8215);
or U9999 (N_9999,N_8291,N_7681);
and U10000 (N_10000,N_8236,N_8338);
and U10001 (N_10001,N_8168,N_7911);
nand U10002 (N_10002,N_7910,N_8446);
nor U10003 (N_10003,N_7675,N_7528);
and U10004 (N_10004,N_7507,N_8494);
nand U10005 (N_10005,N_8114,N_8175);
nor U10006 (N_10006,N_7625,N_8161);
nand U10007 (N_10007,N_8859,N_7706);
or U10008 (N_10008,N_8980,N_7542);
nand U10009 (N_10009,N_8829,N_7616);
and U10010 (N_10010,N_8173,N_8625);
or U10011 (N_10011,N_8783,N_8488);
xor U10012 (N_10012,N_8930,N_8253);
and U10013 (N_10013,N_8048,N_8049);
and U10014 (N_10014,N_8282,N_8975);
nand U10015 (N_10015,N_7611,N_8265);
xor U10016 (N_10016,N_8892,N_8570);
and U10017 (N_10017,N_7745,N_8898);
and U10018 (N_10018,N_8092,N_7854);
xor U10019 (N_10019,N_8395,N_8325);
xor U10020 (N_10020,N_8981,N_8242);
or U10021 (N_10021,N_8656,N_8097);
and U10022 (N_10022,N_7568,N_7613);
and U10023 (N_10023,N_8470,N_8780);
or U10024 (N_10024,N_8058,N_7949);
and U10025 (N_10025,N_8702,N_7632);
nand U10026 (N_10026,N_7592,N_8701);
xnor U10027 (N_10027,N_8733,N_8232);
or U10028 (N_10028,N_7774,N_7874);
and U10029 (N_10029,N_8230,N_8492);
or U10030 (N_10030,N_8845,N_7778);
and U10031 (N_10031,N_7940,N_8527);
nor U10032 (N_10032,N_8068,N_8870);
xnor U10033 (N_10033,N_7940,N_8698);
or U10034 (N_10034,N_7795,N_8667);
and U10035 (N_10035,N_8643,N_7822);
or U10036 (N_10036,N_8330,N_7760);
xnor U10037 (N_10037,N_8589,N_8189);
xor U10038 (N_10038,N_7555,N_8791);
nand U10039 (N_10039,N_8942,N_8785);
or U10040 (N_10040,N_8699,N_8553);
nor U10041 (N_10041,N_8437,N_8817);
nand U10042 (N_10042,N_8092,N_8200);
or U10043 (N_10043,N_7663,N_8086);
nor U10044 (N_10044,N_7632,N_8712);
or U10045 (N_10045,N_7821,N_8317);
xor U10046 (N_10046,N_8316,N_8293);
nor U10047 (N_10047,N_8220,N_8669);
xor U10048 (N_10048,N_8884,N_8867);
or U10049 (N_10049,N_8920,N_8839);
nor U10050 (N_10050,N_8360,N_8068);
nor U10051 (N_10051,N_8687,N_8752);
or U10052 (N_10052,N_7865,N_7913);
nand U10053 (N_10053,N_7605,N_7734);
and U10054 (N_10054,N_8317,N_7947);
nor U10055 (N_10055,N_8067,N_7503);
xor U10056 (N_10056,N_8212,N_7659);
nand U10057 (N_10057,N_8781,N_8233);
nand U10058 (N_10058,N_7800,N_8629);
or U10059 (N_10059,N_7529,N_7915);
nor U10060 (N_10060,N_7879,N_8245);
nand U10061 (N_10061,N_8296,N_8406);
nor U10062 (N_10062,N_8468,N_8393);
and U10063 (N_10063,N_8236,N_7530);
xor U10064 (N_10064,N_7839,N_8175);
or U10065 (N_10065,N_7661,N_8680);
nor U10066 (N_10066,N_8595,N_8637);
xnor U10067 (N_10067,N_8185,N_7766);
or U10068 (N_10068,N_7877,N_8675);
nand U10069 (N_10069,N_8263,N_8635);
or U10070 (N_10070,N_8592,N_8995);
nor U10071 (N_10071,N_8334,N_8473);
xnor U10072 (N_10072,N_7602,N_8415);
nand U10073 (N_10073,N_8222,N_8981);
and U10074 (N_10074,N_7792,N_8104);
xnor U10075 (N_10075,N_8787,N_8647);
and U10076 (N_10076,N_8600,N_8005);
nor U10077 (N_10077,N_8436,N_7776);
and U10078 (N_10078,N_8310,N_8858);
or U10079 (N_10079,N_7671,N_8360);
xnor U10080 (N_10080,N_8710,N_8265);
or U10081 (N_10081,N_7533,N_7517);
nor U10082 (N_10082,N_8696,N_8358);
nor U10083 (N_10083,N_7858,N_7640);
nor U10084 (N_10084,N_8856,N_7699);
xnor U10085 (N_10085,N_8699,N_8779);
nor U10086 (N_10086,N_8264,N_8725);
and U10087 (N_10087,N_8875,N_8426);
xnor U10088 (N_10088,N_8644,N_8871);
xnor U10089 (N_10089,N_7852,N_8368);
and U10090 (N_10090,N_8370,N_7955);
nand U10091 (N_10091,N_7831,N_8295);
and U10092 (N_10092,N_7630,N_8784);
or U10093 (N_10093,N_7697,N_8686);
or U10094 (N_10094,N_8644,N_7681);
or U10095 (N_10095,N_8827,N_7622);
or U10096 (N_10096,N_7823,N_8035);
nand U10097 (N_10097,N_8793,N_8916);
and U10098 (N_10098,N_7861,N_8839);
xnor U10099 (N_10099,N_8585,N_8171);
xnor U10100 (N_10100,N_8827,N_8790);
or U10101 (N_10101,N_8202,N_7805);
nor U10102 (N_10102,N_7614,N_7949);
nand U10103 (N_10103,N_8827,N_7702);
nor U10104 (N_10104,N_7936,N_8111);
nand U10105 (N_10105,N_7835,N_8362);
nor U10106 (N_10106,N_7695,N_8312);
xor U10107 (N_10107,N_7549,N_8203);
or U10108 (N_10108,N_8946,N_7615);
or U10109 (N_10109,N_8904,N_7793);
and U10110 (N_10110,N_7657,N_7915);
nor U10111 (N_10111,N_8008,N_8554);
nand U10112 (N_10112,N_7566,N_7638);
nand U10113 (N_10113,N_8267,N_7601);
and U10114 (N_10114,N_7656,N_7516);
and U10115 (N_10115,N_7705,N_8738);
nor U10116 (N_10116,N_7689,N_8906);
xor U10117 (N_10117,N_7894,N_8331);
nor U10118 (N_10118,N_8626,N_8957);
or U10119 (N_10119,N_8889,N_7869);
nor U10120 (N_10120,N_8270,N_8015);
nand U10121 (N_10121,N_8776,N_7779);
nand U10122 (N_10122,N_8425,N_8101);
xnor U10123 (N_10123,N_8883,N_8394);
or U10124 (N_10124,N_8392,N_8633);
and U10125 (N_10125,N_7522,N_7971);
nor U10126 (N_10126,N_8176,N_7840);
or U10127 (N_10127,N_8292,N_7699);
xnor U10128 (N_10128,N_8741,N_7901);
nor U10129 (N_10129,N_8257,N_8210);
xor U10130 (N_10130,N_8412,N_8608);
nand U10131 (N_10131,N_8745,N_8650);
nand U10132 (N_10132,N_7935,N_8427);
and U10133 (N_10133,N_8370,N_7867);
or U10134 (N_10134,N_8832,N_8276);
or U10135 (N_10135,N_8739,N_7533);
nor U10136 (N_10136,N_7563,N_8016);
or U10137 (N_10137,N_8469,N_8761);
or U10138 (N_10138,N_8404,N_8954);
xor U10139 (N_10139,N_8467,N_7725);
or U10140 (N_10140,N_8649,N_8111);
nand U10141 (N_10141,N_8042,N_7613);
nor U10142 (N_10142,N_8105,N_8233);
or U10143 (N_10143,N_8783,N_7778);
and U10144 (N_10144,N_8751,N_8761);
xnor U10145 (N_10145,N_8642,N_8698);
and U10146 (N_10146,N_8766,N_7938);
nor U10147 (N_10147,N_8726,N_7556);
xnor U10148 (N_10148,N_7733,N_7941);
and U10149 (N_10149,N_7792,N_7951);
xor U10150 (N_10150,N_8176,N_8265);
nand U10151 (N_10151,N_7513,N_8236);
or U10152 (N_10152,N_8349,N_7815);
or U10153 (N_10153,N_8653,N_8744);
nand U10154 (N_10154,N_7933,N_8725);
or U10155 (N_10155,N_7900,N_8264);
nand U10156 (N_10156,N_8927,N_7909);
nor U10157 (N_10157,N_8335,N_8290);
nor U10158 (N_10158,N_7818,N_8252);
nand U10159 (N_10159,N_7978,N_8544);
xnor U10160 (N_10160,N_7629,N_7627);
xnor U10161 (N_10161,N_8757,N_8539);
or U10162 (N_10162,N_8241,N_8629);
and U10163 (N_10163,N_8216,N_8388);
nand U10164 (N_10164,N_8181,N_8781);
nor U10165 (N_10165,N_7784,N_8084);
nor U10166 (N_10166,N_7669,N_8135);
and U10167 (N_10167,N_8183,N_8864);
or U10168 (N_10168,N_7588,N_8575);
or U10169 (N_10169,N_8340,N_7955);
or U10170 (N_10170,N_8200,N_8273);
nor U10171 (N_10171,N_8957,N_8486);
and U10172 (N_10172,N_7963,N_8624);
nor U10173 (N_10173,N_8708,N_8348);
or U10174 (N_10174,N_8620,N_8838);
and U10175 (N_10175,N_7854,N_8243);
xor U10176 (N_10176,N_8320,N_8895);
nand U10177 (N_10177,N_8236,N_8826);
or U10178 (N_10178,N_7541,N_8856);
xnor U10179 (N_10179,N_8787,N_7830);
nand U10180 (N_10180,N_7597,N_8848);
nand U10181 (N_10181,N_8568,N_8377);
or U10182 (N_10182,N_7667,N_7542);
nor U10183 (N_10183,N_8473,N_8880);
nand U10184 (N_10184,N_8966,N_8424);
nand U10185 (N_10185,N_8422,N_7994);
and U10186 (N_10186,N_8479,N_7900);
or U10187 (N_10187,N_7882,N_7887);
nor U10188 (N_10188,N_7929,N_8836);
nor U10189 (N_10189,N_7569,N_7775);
or U10190 (N_10190,N_8341,N_7572);
nor U10191 (N_10191,N_7975,N_8686);
nand U10192 (N_10192,N_8297,N_8738);
nand U10193 (N_10193,N_7759,N_8051);
nor U10194 (N_10194,N_8267,N_8495);
or U10195 (N_10195,N_8318,N_7505);
or U10196 (N_10196,N_8479,N_8284);
and U10197 (N_10197,N_7560,N_8755);
and U10198 (N_10198,N_8611,N_7564);
xor U10199 (N_10199,N_8728,N_8563);
and U10200 (N_10200,N_7984,N_8362);
xnor U10201 (N_10201,N_7598,N_8105);
and U10202 (N_10202,N_8222,N_7779);
and U10203 (N_10203,N_8733,N_8983);
xor U10204 (N_10204,N_8926,N_8478);
nand U10205 (N_10205,N_8569,N_8880);
and U10206 (N_10206,N_8456,N_8948);
nor U10207 (N_10207,N_7931,N_7821);
or U10208 (N_10208,N_8234,N_7901);
or U10209 (N_10209,N_7661,N_7816);
nor U10210 (N_10210,N_7857,N_7579);
or U10211 (N_10211,N_7698,N_8953);
and U10212 (N_10212,N_7871,N_7969);
xor U10213 (N_10213,N_8852,N_8426);
or U10214 (N_10214,N_7927,N_8961);
nor U10215 (N_10215,N_7922,N_7747);
xor U10216 (N_10216,N_8510,N_7855);
nand U10217 (N_10217,N_7822,N_8205);
xnor U10218 (N_10218,N_7544,N_8684);
nand U10219 (N_10219,N_8217,N_7762);
nor U10220 (N_10220,N_8559,N_8504);
xor U10221 (N_10221,N_8205,N_7565);
nor U10222 (N_10222,N_8394,N_7747);
or U10223 (N_10223,N_8964,N_7723);
xnor U10224 (N_10224,N_7966,N_8758);
xnor U10225 (N_10225,N_8556,N_8237);
or U10226 (N_10226,N_7767,N_8545);
nand U10227 (N_10227,N_7849,N_8599);
or U10228 (N_10228,N_7916,N_8031);
and U10229 (N_10229,N_8239,N_8535);
or U10230 (N_10230,N_8409,N_8343);
xnor U10231 (N_10231,N_7574,N_8304);
nor U10232 (N_10232,N_8916,N_8120);
nor U10233 (N_10233,N_8395,N_8447);
and U10234 (N_10234,N_8815,N_7714);
nor U10235 (N_10235,N_8999,N_7762);
or U10236 (N_10236,N_8580,N_8056);
nor U10237 (N_10237,N_8946,N_8321);
xnor U10238 (N_10238,N_8435,N_8763);
nand U10239 (N_10239,N_8735,N_8242);
nand U10240 (N_10240,N_8355,N_8297);
xnor U10241 (N_10241,N_7882,N_8477);
nor U10242 (N_10242,N_7547,N_8801);
nand U10243 (N_10243,N_8220,N_8005);
nand U10244 (N_10244,N_7558,N_7622);
nand U10245 (N_10245,N_7596,N_7697);
xor U10246 (N_10246,N_8087,N_8080);
or U10247 (N_10247,N_7816,N_8008);
nor U10248 (N_10248,N_7580,N_8645);
xor U10249 (N_10249,N_8413,N_8176);
nand U10250 (N_10250,N_7707,N_7901);
and U10251 (N_10251,N_8180,N_8360);
or U10252 (N_10252,N_8322,N_7555);
xor U10253 (N_10253,N_8308,N_8385);
and U10254 (N_10254,N_7780,N_8774);
nand U10255 (N_10255,N_7524,N_8038);
nand U10256 (N_10256,N_8170,N_8437);
or U10257 (N_10257,N_8312,N_7754);
or U10258 (N_10258,N_7776,N_7563);
xor U10259 (N_10259,N_7957,N_8576);
xnor U10260 (N_10260,N_8598,N_7516);
and U10261 (N_10261,N_8937,N_7535);
and U10262 (N_10262,N_8934,N_7915);
nand U10263 (N_10263,N_8094,N_8566);
xor U10264 (N_10264,N_8324,N_8557);
nand U10265 (N_10265,N_8412,N_8658);
and U10266 (N_10266,N_8419,N_8939);
or U10267 (N_10267,N_7511,N_7553);
or U10268 (N_10268,N_7791,N_8109);
nand U10269 (N_10269,N_7633,N_8250);
or U10270 (N_10270,N_8582,N_8377);
or U10271 (N_10271,N_7956,N_8727);
or U10272 (N_10272,N_8247,N_7748);
nor U10273 (N_10273,N_8694,N_8314);
or U10274 (N_10274,N_7650,N_8984);
nor U10275 (N_10275,N_7876,N_8985);
nor U10276 (N_10276,N_8850,N_8713);
nor U10277 (N_10277,N_7789,N_8378);
nand U10278 (N_10278,N_8799,N_7653);
nand U10279 (N_10279,N_8984,N_8132);
xnor U10280 (N_10280,N_8350,N_8216);
nand U10281 (N_10281,N_7802,N_8944);
nor U10282 (N_10282,N_7920,N_8168);
or U10283 (N_10283,N_8626,N_8365);
or U10284 (N_10284,N_8615,N_8624);
nor U10285 (N_10285,N_8287,N_8357);
nand U10286 (N_10286,N_7890,N_7809);
and U10287 (N_10287,N_8302,N_7741);
nor U10288 (N_10288,N_8959,N_8230);
and U10289 (N_10289,N_8232,N_8356);
nand U10290 (N_10290,N_7743,N_7610);
and U10291 (N_10291,N_8487,N_7589);
and U10292 (N_10292,N_7507,N_8962);
or U10293 (N_10293,N_7734,N_8158);
and U10294 (N_10294,N_8243,N_8104);
or U10295 (N_10295,N_7695,N_8785);
nand U10296 (N_10296,N_7574,N_7622);
or U10297 (N_10297,N_7787,N_8392);
and U10298 (N_10298,N_7718,N_8017);
nor U10299 (N_10299,N_8720,N_7877);
xor U10300 (N_10300,N_8925,N_8091);
xnor U10301 (N_10301,N_8876,N_7729);
nand U10302 (N_10302,N_8310,N_8776);
or U10303 (N_10303,N_8080,N_7840);
xor U10304 (N_10304,N_8216,N_8693);
or U10305 (N_10305,N_8885,N_7586);
or U10306 (N_10306,N_7775,N_8367);
nor U10307 (N_10307,N_7829,N_8085);
nor U10308 (N_10308,N_8843,N_8198);
nor U10309 (N_10309,N_8924,N_8294);
or U10310 (N_10310,N_8219,N_8009);
nand U10311 (N_10311,N_8271,N_8985);
nand U10312 (N_10312,N_8892,N_8190);
nand U10313 (N_10313,N_8348,N_7715);
or U10314 (N_10314,N_7634,N_8040);
nand U10315 (N_10315,N_7581,N_7876);
and U10316 (N_10316,N_7867,N_8696);
xor U10317 (N_10317,N_7954,N_8412);
xor U10318 (N_10318,N_8783,N_8349);
nor U10319 (N_10319,N_7732,N_8145);
nand U10320 (N_10320,N_7687,N_8424);
nand U10321 (N_10321,N_8169,N_8185);
or U10322 (N_10322,N_8304,N_8020);
nand U10323 (N_10323,N_8768,N_8950);
or U10324 (N_10324,N_8943,N_7756);
nor U10325 (N_10325,N_8201,N_7934);
nor U10326 (N_10326,N_8735,N_8910);
and U10327 (N_10327,N_7562,N_8396);
and U10328 (N_10328,N_8717,N_7982);
nor U10329 (N_10329,N_7750,N_8960);
nand U10330 (N_10330,N_8809,N_7527);
nand U10331 (N_10331,N_8064,N_7784);
xnor U10332 (N_10332,N_8917,N_8550);
or U10333 (N_10333,N_7709,N_7958);
xor U10334 (N_10334,N_8651,N_7950);
nor U10335 (N_10335,N_7618,N_8176);
nor U10336 (N_10336,N_8695,N_8717);
and U10337 (N_10337,N_8777,N_8031);
xor U10338 (N_10338,N_8465,N_8784);
or U10339 (N_10339,N_7894,N_8282);
or U10340 (N_10340,N_8550,N_7984);
xor U10341 (N_10341,N_7831,N_8967);
nor U10342 (N_10342,N_8752,N_8067);
and U10343 (N_10343,N_8350,N_8069);
nand U10344 (N_10344,N_7654,N_7526);
or U10345 (N_10345,N_8341,N_7736);
and U10346 (N_10346,N_7869,N_8781);
nor U10347 (N_10347,N_7522,N_8629);
or U10348 (N_10348,N_8256,N_8089);
or U10349 (N_10349,N_7915,N_8235);
xor U10350 (N_10350,N_7690,N_8798);
and U10351 (N_10351,N_8021,N_7759);
or U10352 (N_10352,N_7825,N_7960);
xor U10353 (N_10353,N_7616,N_7597);
nand U10354 (N_10354,N_8245,N_7846);
nand U10355 (N_10355,N_8104,N_7946);
or U10356 (N_10356,N_8676,N_7811);
xor U10357 (N_10357,N_8090,N_8873);
nor U10358 (N_10358,N_7793,N_7961);
nand U10359 (N_10359,N_8490,N_8244);
nand U10360 (N_10360,N_8601,N_8117);
or U10361 (N_10361,N_7949,N_7912);
nand U10362 (N_10362,N_7615,N_8717);
and U10363 (N_10363,N_8266,N_7568);
nor U10364 (N_10364,N_7569,N_7789);
and U10365 (N_10365,N_7781,N_7701);
xnor U10366 (N_10366,N_8595,N_8177);
nor U10367 (N_10367,N_7917,N_8034);
or U10368 (N_10368,N_8649,N_8985);
nand U10369 (N_10369,N_7577,N_7744);
and U10370 (N_10370,N_8286,N_7680);
or U10371 (N_10371,N_7749,N_8621);
or U10372 (N_10372,N_8393,N_8960);
xor U10373 (N_10373,N_8117,N_8284);
and U10374 (N_10374,N_8476,N_8153);
xnor U10375 (N_10375,N_7904,N_7899);
xor U10376 (N_10376,N_7500,N_8066);
nand U10377 (N_10377,N_7511,N_7515);
nor U10378 (N_10378,N_7832,N_8979);
nor U10379 (N_10379,N_8938,N_7879);
nor U10380 (N_10380,N_7714,N_8059);
and U10381 (N_10381,N_8471,N_8313);
nand U10382 (N_10382,N_7702,N_8158);
and U10383 (N_10383,N_8141,N_7613);
xnor U10384 (N_10384,N_8371,N_8991);
xnor U10385 (N_10385,N_8850,N_8156);
nor U10386 (N_10386,N_7501,N_7664);
nor U10387 (N_10387,N_8383,N_8428);
xor U10388 (N_10388,N_7547,N_8313);
nor U10389 (N_10389,N_7662,N_8535);
nor U10390 (N_10390,N_8964,N_7632);
xor U10391 (N_10391,N_8973,N_8990);
nand U10392 (N_10392,N_8705,N_8419);
xor U10393 (N_10393,N_7938,N_8284);
xor U10394 (N_10394,N_7660,N_7634);
or U10395 (N_10395,N_8858,N_8495);
and U10396 (N_10396,N_8769,N_8884);
nor U10397 (N_10397,N_8510,N_7738);
xnor U10398 (N_10398,N_7851,N_8642);
nand U10399 (N_10399,N_8547,N_8231);
nand U10400 (N_10400,N_8614,N_8669);
xnor U10401 (N_10401,N_7553,N_7649);
xnor U10402 (N_10402,N_8179,N_8466);
nand U10403 (N_10403,N_8843,N_8193);
or U10404 (N_10404,N_7963,N_8713);
nand U10405 (N_10405,N_8605,N_7561);
or U10406 (N_10406,N_8969,N_7924);
nand U10407 (N_10407,N_7622,N_7562);
nor U10408 (N_10408,N_8899,N_8408);
nor U10409 (N_10409,N_8302,N_7594);
nor U10410 (N_10410,N_7518,N_7544);
nand U10411 (N_10411,N_7729,N_8619);
nand U10412 (N_10412,N_8785,N_8652);
nand U10413 (N_10413,N_8675,N_8437);
nand U10414 (N_10414,N_7894,N_8831);
nor U10415 (N_10415,N_8835,N_8335);
xnor U10416 (N_10416,N_8322,N_7981);
nand U10417 (N_10417,N_7602,N_8390);
and U10418 (N_10418,N_8154,N_7552);
nand U10419 (N_10419,N_8450,N_8163);
or U10420 (N_10420,N_7574,N_7521);
or U10421 (N_10421,N_8118,N_8462);
nor U10422 (N_10422,N_8990,N_7911);
or U10423 (N_10423,N_8005,N_8653);
or U10424 (N_10424,N_7620,N_8511);
xor U10425 (N_10425,N_8735,N_7666);
nand U10426 (N_10426,N_8149,N_8123);
xor U10427 (N_10427,N_7622,N_7748);
nand U10428 (N_10428,N_8952,N_7515);
and U10429 (N_10429,N_8887,N_8676);
or U10430 (N_10430,N_7839,N_7580);
xor U10431 (N_10431,N_8055,N_8322);
xnor U10432 (N_10432,N_8676,N_8368);
xor U10433 (N_10433,N_8103,N_8658);
nand U10434 (N_10434,N_7804,N_7862);
xnor U10435 (N_10435,N_7807,N_8122);
nor U10436 (N_10436,N_8761,N_7982);
or U10437 (N_10437,N_8881,N_8932);
or U10438 (N_10438,N_8670,N_8185);
and U10439 (N_10439,N_8592,N_8935);
nor U10440 (N_10440,N_8174,N_8425);
or U10441 (N_10441,N_7972,N_7642);
and U10442 (N_10442,N_8306,N_8352);
nor U10443 (N_10443,N_8275,N_8473);
nor U10444 (N_10444,N_7861,N_7539);
nor U10445 (N_10445,N_8036,N_8028);
nand U10446 (N_10446,N_7811,N_8905);
nor U10447 (N_10447,N_8830,N_8602);
or U10448 (N_10448,N_8606,N_8387);
xnor U10449 (N_10449,N_8431,N_7807);
nand U10450 (N_10450,N_8876,N_8921);
xor U10451 (N_10451,N_8332,N_7631);
and U10452 (N_10452,N_8626,N_8782);
xor U10453 (N_10453,N_7905,N_7705);
xnor U10454 (N_10454,N_8562,N_8225);
or U10455 (N_10455,N_8728,N_8245);
or U10456 (N_10456,N_7901,N_8331);
nand U10457 (N_10457,N_8368,N_8844);
and U10458 (N_10458,N_8254,N_8496);
xnor U10459 (N_10459,N_7802,N_8960);
nor U10460 (N_10460,N_8087,N_8681);
and U10461 (N_10461,N_8727,N_7507);
nor U10462 (N_10462,N_8689,N_8957);
nor U10463 (N_10463,N_8207,N_8952);
and U10464 (N_10464,N_7523,N_8588);
and U10465 (N_10465,N_8314,N_8817);
nor U10466 (N_10466,N_7568,N_7817);
and U10467 (N_10467,N_8439,N_7917);
and U10468 (N_10468,N_8253,N_8014);
xor U10469 (N_10469,N_7825,N_8614);
and U10470 (N_10470,N_8798,N_8055);
xnor U10471 (N_10471,N_8478,N_8438);
xnor U10472 (N_10472,N_7870,N_8620);
and U10473 (N_10473,N_8636,N_8296);
nor U10474 (N_10474,N_8727,N_8641);
nand U10475 (N_10475,N_8454,N_8936);
and U10476 (N_10476,N_7898,N_7807);
and U10477 (N_10477,N_7875,N_7703);
nor U10478 (N_10478,N_8547,N_7711);
xnor U10479 (N_10479,N_8997,N_8538);
and U10480 (N_10480,N_7917,N_8469);
nor U10481 (N_10481,N_7838,N_8032);
and U10482 (N_10482,N_8631,N_7516);
or U10483 (N_10483,N_7635,N_8083);
or U10484 (N_10484,N_8825,N_8115);
nor U10485 (N_10485,N_7983,N_7763);
xor U10486 (N_10486,N_8920,N_8987);
or U10487 (N_10487,N_8112,N_7554);
xor U10488 (N_10488,N_8892,N_8248);
or U10489 (N_10489,N_7716,N_7555);
nor U10490 (N_10490,N_8194,N_7801);
or U10491 (N_10491,N_7724,N_8857);
nand U10492 (N_10492,N_8821,N_8402);
and U10493 (N_10493,N_8943,N_8309);
and U10494 (N_10494,N_7752,N_7946);
nand U10495 (N_10495,N_8826,N_8904);
or U10496 (N_10496,N_7624,N_7500);
and U10497 (N_10497,N_7844,N_8133);
xor U10498 (N_10498,N_8394,N_8085);
or U10499 (N_10499,N_8297,N_8304);
and U10500 (N_10500,N_9211,N_9588);
or U10501 (N_10501,N_10445,N_9248);
and U10502 (N_10502,N_10014,N_10027);
or U10503 (N_10503,N_10345,N_9142);
nor U10504 (N_10504,N_9400,N_10354);
xor U10505 (N_10505,N_9589,N_9693);
nor U10506 (N_10506,N_10149,N_10444);
nor U10507 (N_10507,N_10464,N_9104);
or U10508 (N_10508,N_9125,N_9455);
and U10509 (N_10509,N_9658,N_10315);
nor U10510 (N_10510,N_9661,N_9164);
and U10511 (N_10511,N_9408,N_9791);
nand U10512 (N_10512,N_10299,N_9637);
nand U10513 (N_10513,N_10408,N_9959);
nor U10514 (N_10514,N_9702,N_10333);
nand U10515 (N_10515,N_9007,N_9941);
or U10516 (N_10516,N_9134,N_9127);
and U10517 (N_10517,N_10317,N_10339);
nand U10518 (N_10518,N_9648,N_9472);
nor U10519 (N_10519,N_9535,N_10072);
xor U10520 (N_10520,N_9691,N_9527);
xnor U10521 (N_10521,N_9572,N_9521);
nand U10522 (N_10522,N_9253,N_9234);
or U10523 (N_10523,N_9875,N_9516);
xor U10524 (N_10524,N_9450,N_9943);
nand U10525 (N_10525,N_9321,N_9093);
and U10526 (N_10526,N_9448,N_9124);
or U10527 (N_10527,N_9928,N_9157);
or U10528 (N_10528,N_9641,N_9984);
nand U10529 (N_10529,N_9267,N_9489);
nand U10530 (N_10530,N_9368,N_10024);
nor U10531 (N_10531,N_10092,N_9704);
or U10532 (N_10532,N_10214,N_10434);
and U10533 (N_10533,N_10300,N_9401);
nor U10534 (N_10534,N_9505,N_9882);
xnor U10535 (N_10535,N_10261,N_10351);
or U10536 (N_10536,N_9039,N_10277);
nand U10537 (N_10537,N_9915,N_9445);
or U10538 (N_10538,N_10053,N_9366);
xor U10539 (N_10539,N_9724,N_10198);
or U10540 (N_10540,N_9814,N_9813);
xor U10541 (N_10541,N_9195,N_10468);
or U10542 (N_10542,N_9439,N_10347);
xor U10543 (N_10543,N_9676,N_10302);
nand U10544 (N_10544,N_9895,N_9912);
nor U10545 (N_10545,N_10303,N_9871);
or U10546 (N_10546,N_9189,N_9683);
nand U10547 (N_10547,N_9059,N_10242);
and U10548 (N_10548,N_9259,N_10356);
xor U10549 (N_10549,N_10078,N_9162);
xor U10550 (N_10550,N_9126,N_9907);
or U10551 (N_10551,N_10153,N_9832);
or U10552 (N_10552,N_9014,N_9231);
nor U10553 (N_10553,N_10297,N_9414);
and U10554 (N_10554,N_9388,N_10268);
and U10555 (N_10555,N_9734,N_9640);
nand U10556 (N_10556,N_10201,N_9772);
and U10557 (N_10557,N_9046,N_9602);
or U10558 (N_10558,N_10113,N_10022);
nor U10559 (N_10559,N_10013,N_10428);
and U10560 (N_10560,N_9333,N_9056);
xor U10561 (N_10561,N_9733,N_9203);
or U10562 (N_10562,N_10115,N_10382);
xor U10563 (N_10563,N_9787,N_9083);
nor U10564 (N_10564,N_9576,N_9753);
xnor U10565 (N_10565,N_9365,N_10417);
xnor U10566 (N_10566,N_10017,N_10295);
or U10567 (N_10567,N_9156,N_9770);
xnor U10568 (N_10568,N_9725,N_9543);
xor U10569 (N_10569,N_10367,N_9235);
nand U10570 (N_10570,N_9573,N_10344);
and U10571 (N_10571,N_10025,N_10184);
and U10572 (N_10572,N_10070,N_9533);
nand U10573 (N_10573,N_10392,N_9993);
and U10574 (N_10574,N_9372,N_9990);
or U10575 (N_10575,N_9577,N_9247);
nor U10576 (N_10576,N_9120,N_9161);
xnor U10577 (N_10577,N_9062,N_9567);
or U10578 (N_10578,N_9828,N_9740);
and U10579 (N_10579,N_9902,N_9611);
and U10580 (N_10580,N_9181,N_9051);
or U10581 (N_10581,N_10438,N_10418);
xor U10582 (N_10582,N_9668,N_9284);
nor U10583 (N_10583,N_10177,N_9979);
and U10584 (N_10584,N_9595,N_9122);
and U10585 (N_10585,N_9716,N_10056);
nor U10586 (N_10586,N_9881,N_9295);
and U10587 (N_10587,N_10081,N_10101);
or U10588 (N_10588,N_9252,N_9242);
xor U10589 (N_10589,N_9584,N_10217);
and U10590 (N_10590,N_9262,N_10135);
and U10591 (N_10591,N_9416,N_9530);
or U10592 (N_10592,N_9382,N_10485);
xnor U10593 (N_10593,N_10439,N_9158);
and U10594 (N_10594,N_10038,N_10362);
xor U10595 (N_10595,N_9592,N_9167);
xnor U10596 (N_10596,N_9954,N_9698);
xnor U10597 (N_10597,N_9723,N_9280);
xnor U10598 (N_10598,N_9310,N_9481);
or U10599 (N_10599,N_9047,N_9425);
xor U10600 (N_10600,N_9298,N_9623);
and U10601 (N_10601,N_9876,N_9249);
or U10602 (N_10602,N_9088,N_9901);
or U10603 (N_10603,N_9357,N_10009);
nor U10604 (N_10604,N_9410,N_10373);
and U10605 (N_10605,N_9739,N_9620);
nor U10606 (N_10606,N_9258,N_9309);
nor U10607 (N_10607,N_9290,N_10194);
and U10608 (N_10608,N_9135,N_10257);
and U10609 (N_10609,N_9672,N_10465);
nor U10610 (N_10610,N_9475,N_9370);
and U10611 (N_10611,N_9524,N_9349);
nor U10612 (N_10612,N_10415,N_9340);
nor U10613 (N_10613,N_9557,N_9735);
or U10614 (N_10614,N_9462,N_9392);
or U10615 (N_10615,N_9794,N_9376);
and U10616 (N_10616,N_9112,N_9515);
or U10617 (N_10617,N_9497,N_10309);
xor U10618 (N_10618,N_10323,N_10479);
nor U10619 (N_10619,N_9810,N_9699);
nor U10620 (N_10620,N_9304,N_10091);
nor U10621 (N_10621,N_9800,N_9100);
and U10622 (N_10622,N_9453,N_9465);
nand U10623 (N_10623,N_9168,N_9706);
nor U10624 (N_10624,N_9916,N_9406);
or U10625 (N_10625,N_9621,N_10100);
nor U10626 (N_10626,N_9237,N_9694);
xnor U10627 (N_10627,N_9331,N_9049);
nand U10628 (N_10628,N_9525,N_9351);
nand U10629 (N_10629,N_9456,N_9469);
xnor U10630 (N_10630,N_10394,N_9415);
and U10631 (N_10631,N_10493,N_9170);
xnor U10632 (N_10632,N_9457,N_9685);
nand U10633 (N_10633,N_9487,N_10316);
nand U10634 (N_10634,N_10234,N_10168);
nand U10635 (N_10635,N_9485,N_10369);
xor U10636 (N_10636,N_10384,N_10290);
and U10637 (N_10637,N_9617,N_9279);
xnor U10638 (N_10638,N_10232,N_9562);
and U10639 (N_10639,N_10086,N_10121);
xor U10640 (N_10640,N_9356,N_10429);
nor U10641 (N_10641,N_10243,N_10364);
and U10642 (N_10642,N_9609,N_9643);
nor U10643 (N_10643,N_10377,N_9380);
xnor U10644 (N_10644,N_10080,N_10007);
and U10645 (N_10645,N_9675,N_9674);
and U10646 (N_10646,N_9982,N_10338);
nor U10647 (N_10647,N_9361,N_9980);
nand U10648 (N_10648,N_9728,N_9950);
and U10649 (N_10649,N_9520,N_9085);
nor U10650 (N_10650,N_9801,N_9574);
nand U10651 (N_10651,N_10467,N_9468);
nand U10652 (N_10652,N_9452,N_10123);
nor U10653 (N_10653,N_10361,N_10008);
or U10654 (N_10654,N_10205,N_9583);
nand U10655 (N_10655,N_9552,N_10348);
or U10656 (N_10656,N_9549,N_10402);
and U10657 (N_10657,N_10156,N_10193);
and U10658 (N_10658,N_9116,N_9955);
nor U10659 (N_10659,N_9246,N_9829);
or U10660 (N_10660,N_9146,N_9075);
xnor U10661 (N_10661,N_9834,N_9068);
nor U10662 (N_10662,N_10462,N_9710);
xnor U10663 (N_10663,N_9782,N_10474);
and U10664 (N_10664,N_9656,N_10167);
or U10665 (N_10665,N_9303,N_9273);
nor U10666 (N_10666,N_10137,N_9846);
nand U10667 (N_10667,N_10125,N_9581);
nor U10668 (N_10668,N_10222,N_10179);
or U10669 (N_10669,N_10108,N_10247);
and U10670 (N_10670,N_9276,N_9073);
or U10671 (N_10671,N_9060,N_10142);
nand U10672 (N_10672,N_9934,N_10074);
nor U10673 (N_10673,N_9551,N_9287);
xor U10674 (N_10674,N_9250,N_9722);
or U10675 (N_10675,N_9300,N_9080);
and U10676 (N_10676,N_10237,N_9783);
nand U10677 (N_10677,N_9216,N_9914);
xor U10678 (N_10678,N_10202,N_9850);
nor U10679 (N_10679,N_9117,N_9936);
xor U10680 (N_10680,N_9910,N_10158);
or U10681 (N_10681,N_9807,N_9865);
nor U10682 (N_10682,N_9764,N_9681);
nand U10683 (N_10683,N_9671,N_9888);
and U10684 (N_10684,N_9923,N_10131);
and U10685 (N_10685,N_9076,N_10006);
nor U10686 (N_10686,N_10099,N_9669);
xor U10687 (N_10687,N_9209,N_9411);
or U10688 (N_10688,N_9449,N_9114);
nand U10689 (N_10689,N_10151,N_10058);
or U10690 (N_10690,N_9346,N_10094);
nand U10691 (N_10691,N_9695,N_9045);
nor U10692 (N_10692,N_10269,N_9148);
nand U10693 (N_10693,N_9792,N_10204);
and U10694 (N_10694,N_10016,N_9441);
nor U10695 (N_10695,N_10355,N_9678);
nand U10696 (N_10696,N_9731,N_9002);
and U10697 (N_10697,N_9839,N_9514);
nor U10698 (N_10698,N_10319,N_10190);
or U10699 (N_10699,N_9989,N_9956);
or U10700 (N_10700,N_9442,N_9541);
nand U10701 (N_10701,N_10207,N_9610);
and U10702 (N_10702,N_9337,N_9129);
xnor U10703 (N_10703,N_9329,N_10241);
nor U10704 (N_10704,N_9526,N_10145);
nor U10705 (N_10705,N_9155,N_9625);
or U10706 (N_10706,N_10410,N_9556);
nand U10707 (N_10707,N_10189,N_9412);
xor U10708 (N_10708,N_10305,N_9052);
nand U10709 (N_10709,N_9359,N_9585);
nand U10710 (N_10710,N_9296,N_9467);
nand U10711 (N_10711,N_9999,N_10256);
xnor U10712 (N_10712,N_10046,N_10456);
and U10713 (N_10713,N_9808,N_9291);
or U10714 (N_10714,N_9214,N_10229);
or U10715 (N_10715,N_9212,N_9277);
nand U10716 (N_10716,N_9074,N_10065);
nor U10717 (N_10717,N_9221,N_9429);
nor U10718 (N_10718,N_10353,N_9174);
and U10719 (N_10719,N_9024,N_10117);
and U10720 (N_10720,N_9634,N_10152);
xnor U10721 (N_10721,N_10096,N_9599);
and U10722 (N_10722,N_9379,N_9795);
nor U10723 (N_10723,N_9289,N_9391);
nand U10724 (N_10724,N_9496,N_9005);
xor U10725 (N_10725,N_9348,N_10021);
and U10726 (N_10726,N_9630,N_10320);
or U10727 (N_10727,N_9743,N_10363);
nand U10728 (N_10728,N_9664,N_10118);
nor U10729 (N_10729,N_9930,N_9145);
nand U10730 (N_10730,N_9756,N_9210);
xor U10731 (N_10731,N_10488,N_9078);
nor U10732 (N_10732,N_9763,N_10063);
and U10733 (N_10733,N_10276,N_9421);
nand U10734 (N_10734,N_10250,N_9077);
nand U10735 (N_10735,N_10172,N_9711);
or U10736 (N_10736,N_9729,N_10087);
or U10737 (N_10737,N_10228,N_9490);
and U10738 (N_10738,N_9719,N_9872);
or U10739 (N_10739,N_10425,N_9709);
or U10740 (N_10740,N_9926,N_10230);
nor U10741 (N_10741,N_9942,N_9822);
nor U10742 (N_10742,N_9482,N_9089);
nand U10743 (N_10743,N_10448,N_10048);
and U10744 (N_10744,N_9190,N_9427);
and U10745 (N_10745,N_9477,N_9555);
xnor U10746 (N_10746,N_10255,N_9301);
xnor U10747 (N_10747,N_10374,N_10440);
nand U10748 (N_10748,N_9413,N_9447);
or U10749 (N_10749,N_9636,N_9745);
nor U10750 (N_10750,N_9179,N_9435);
or U10751 (N_10751,N_9771,N_10365);
and U10752 (N_10752,N_9633,N_9545);
nor U10753 (N_10753,N_9136,N_10171);
and U10754 (N_10754,N_9084,N_9874);
xnor U10755 (N_10755,N_10358,N_9504);
nor U10756 (N_10756,N_9696,N_10378);
nor U10757 (N_10757,N_9818,N_9920);
nand U10758 (N_10758,N_9517,N_10352);
nor U10759 (N_10759,N_9464,N_9050);
or U10760 (N_10760,N_9799,N_9961);
xor U10761 (N_10761,N_9420,N_10102);
and U10762 (N_10762,N_9629,N_10141);
and U10763 (N_10763,N_9804,N_10258);
xnor U10764 (N_10764,N_9966,N_9500);
nand U10765 (N_10765,N_9809,N_9570);
nand U10766 (N_10766,N_10129,N_9540);
nand U10767 (N_10767,N_10213,N_9236);
and U10768 (N_10768,N_9779,N_9431);
or U10769 (N_10769,N_9836,N_9502);
and U10770 (N_10770,N_10181,N_9879);
nor U10771 (N_10771,N_9697,N_9402);
nand U10772 (N_10772,N_10280,N_9741);
xnor U10773 (N_10773,N_9363,N_9758);
nand U10774 (N_10774,N_9434,N_9529);
or U10775 (N_10775,N_10327,N_9407);
nand U10776 (N_10776,N_9843,N_9451);
nor U10777 (N_10777,N_10238,N_9471);
and U10778 (N_10778,N_9269,N_9578);
xor U10779 (N_10779,N_9769,N_10267);
nand U10780 (N_10780,N_9017,N_9981);
or U10781 (N_10781,N_9048,N_9868);
nor U10782 (N_10782,N_9816,N_9513);
nor U10783 (N_10783,N_9713,N_9384);
nor U10784 (N_10784,N_9043,N_9436);
nor U10785 (N_10785,N_10112,N_9001);
nor U10786 (N_10786,N_9332,N_9659);
nor U10787 (N_10787,N_9183,N_9548);
or U10788 (N_10788,N_10098,N_9624);
xnor U10789 (N_10789,N_9193,N_10029);
xor U10790 (N_10790,N_10391,N_10416);
nor U10791 (N_10791,N_9326,N_9742);
nand U10792 (N_10792,N_9110,N_9369);
nor U10793 (N_10793,N_10340,N_10042);
nand U10794 (N_10794,N_9215,N_9622);
xor U10795 (N_10795,N_10262,N_9564);
or U10796 (N_10796,N_9185,N_9367);
or U10797 (N_10797,N_10043,N_9230);
or U10798 (N_10798,N_9103,N_10388);
nor U10799 (N_10799,N_10155,N_9652);
and U10800 (N_10800,N_9776,N_9393);
and U10801 (N_10801,N_9064,N_9662);
or U10802 (N_10802,N_9948,N_9108);
xnor U10803 (N_10803,N_9243,N_9478);
xor U10804 (N_10804,N_10306,N_9889);
xor U10805 (N_10805,N_9314,N_10076);
or U10806 (N_10806,N_9123,N_10011);
or U10807 (N_10807,N_9880,N_9755);
nor U10808 (N_10808,N_9315,N_9820);
xnor U10809 (N_10809,N_9483,N_10187);
xnor U10810 (N_10810,N_9328,N_9152);
and U10811 (N_10811,N_10265,N_10421);
and U10812 (N_10812,N_9495,N_9650);
nor U10813 (N_10813,N_10055,N_9967);
or U10814 (N_10814,N_10393,N_10329);
and U10815 (N_10815,N_9812,N_10195);
and U10816 (N_10816,N_9786,N_10330);
nand U10817 (N_10817,N_10067,N_9443);
xor U10818 (N_10818,N_10466,N_9878);
or U10819 (N_10819,N_9041,N_9492);
and U10820 (N_10820,N_10138,N_9690);
nor U10821 (N_10821,N_9823,N_9245);
nand U10822 (N_10822,N_9528,N_9021);
or U10823 (N_10823,N_9974,N_9579);
xnor U10824 (N_10824,N_9184,N_9151);
and U10825 (N_10825,N_9618,N_10107);
and U10826 (N_10826,N_10469,N_9983);
or U10827 (N_10827,N_9638,N_10482);
xor U10828 (N_10828,N_10089,N_9859);
or U10829 (N_10829,N_9035,N_9006);
and U10830 (N_10830,N_9373,N_9857);
nor U10831 (N_10831,N_9113,N_9860);
xor U10832 (N_10832,N_9949,N_9774);
xnor U10833 (N_10833,N_9793,N_9946);
nand U10834 (N_10834,N_9199,N_10103);
or U10835 (N_10835,N_9649,N_9119);
and U10836 (N_10836,N_9811,N_9327);
nor U10837 (N_10837,N_9030,N_9225);
or U10838 (N_10838,N_10035,N_9440);
and U10839 (N_10839,N_9261,N_9347);
nor U10840 (N_10840,N_9015,N_9616);
or U10841 (N_10841,N_9299,N_9509);
and U10842 (N_10842,N_9342,N_10490);
or U10843 (N_10843,N_9819,N_9272);
nor U10844 (N_10844,N_9798,N_10331);
or U10845 (N_10845,N_10039,N_9665);
and U10846 (N_10846,N_10463,N_10454);
nand U10847 (N_10847,N_9397,N_10461);
nand U10848 (N_10848,N_9917,N_10165);
or U10849 (N_10849,N_9132,N_9852);
xor U10850 (N_10850,N_9849,N_10475);
and U10851 (N_10851,N_9866,N_10289);
nand U10852 (N_10852,N_9121,N_9603);
or U10853 (N_10853,N_10341,N_9666);
and U10854 (N_10854,N_9994,N_10497);
xnor U10855 (N_10855,N_9985,N_9667);
nand U10856 (N_10856,N_9292,N_10212);
and U10857 (N_10857,N_9969,N_9430);
xnor U10858 (N_10858,N_9647,N_9069);
or U10859 (N_10859,N_9886,N_9682);
xor U10860 (N_10860,N_10307,N_9560);
nor U10861 (N_10861,N_9466,N_10322);
nand U10862 (N_10862,N_9657,N_9925);
or U10863 (N_10863,N_10275,N_9635);
nand U10864 (N_10864,N_9877,N_10128);
and U10865 (N_10865,N_9937,N_9598);
xnor U10866 (N_10866,N_10215,N_9590);
nor U10867 (N_10867,N_9508,N_9172);
xor U10868 (N_10868,N_9751,N_9510);
nand U10869 (N_10869,N_9854,N_10054);
nor U10870 (N_10870,N_9011,N_9867);
nor U10871 (N_10871,N_10376,N_10263);
nand U10872 (N_10872,N_9227,N_10003);
and U10873 (N_10873,N_10208,N_9817);
nand U10874 (N_10874,N_10359,N_9263);
xnor U10875 (N_10875,N_9396,N_9884);
and U10876 (N_10876,N_10431,N_10380);
and U10877 (N_10877,N_10036,N_9345);
and U10878 (N_10878,N_10409,N_9470);
nand U10879 (N_10879,N_10430,N_10426);
nor U10880 (N_10880,N_9824,N_10166);
xor U10881 (N_10881,N_9343,N_10335);
nor U10882 (N_10882,N_10396,N_10203);
or U10883 (N_10883,N_9746,N_10105);
or U10884 (N_10884,N_10270,N_9087);
nand U10885 (N_10885,N_9714,N_10337);
and U10886 (N_10886,N_9547,N_9099);
nand U10887 (N_10887,N_9264,N_9383);
or U10888 (N_10888,N_9257,N_10235);
xor U10889 (N_10889,N_9358,N_10447);
and U10890 (N_10890,N_10032,N_10005);
nor U10891 (N_10891,N_9730,N_10271);
and U10892 (N_10892,N_9270,N_10028);
nand U10893 (N_10893,N_9308,N_9239);
nor U10894 (N_10894,N_9458,N_9196);
or U10895 (N_10895,N_9232,N_9364);
or U10896 (N_10896,N_9686,N_10104);
nand U10897 (N_10897,N_9438,N_9858);
xnor U10898 (N_10898,N_9677,N_9016);
nor U10899 (N_10899,N_9830,N_9405);
nand U10900 (N_10900,N_9921,N_9374);
nor U10901 (N_10901,N_10130,N_9831);
and U10902 (N_10902,N_9175,N_9053);
nor U10903 (N_10903,N_9197,N_10085);
xor U10904 (N_10904,N_9171,N_10150);
and U10905 (N_10905,N_9612,N_9848);
xnor U10906 (N_10906,N_10372,N_9718);
nor U10907 (N_10907,N_9480,N_10071);
xor U10908 (N_10908,N_9484,N_9238);
nor U10909 (N_10909,N_9944,N_9163);
nand U10910 (N_10910,N_9202,N_9098);
or U10911 (N_10911,N_9766,N_9957);
nor U10912 (N_10912,N_9684,N_10209);
nand U10913 (N_10913,N_9097,N_9389);
or U10914 (N_10914,N_9042,N_10383);
and U10915 (N_10915,N_10326,N_9204);
and U10916 (N_10916,N_10147,N_9626);
or U10917 (N_10917,N_10293,N_10459);
or U10918 (N_10918,N_9821,N_9072);
and U10919 (N_10919,N_9815,N_9748);
or U10920 (N_10920,N_9128,N_9404);
or U10921 (N_10921,N_9320,N_10436);
or U10922 (N_10922,N_10225,N_9773);
nor U10923 (N_10923,N_10248,N_9842);
and U10924 (N_10924,N_10231,N_9534);
or U10925 (N_10925,N_10350,N_9803);
and U10926 (N_10926,N_9207,N_9627);
or U10927 (N_10927,N_10489,N_10346);
or U10928 (N_10928,N_10336,N_9101);
and U10929 (N_10929,N_9133,N_10484);
nor U10930 (N_10930,N_9251,N_10492);
nor U10931 (N_10931,N_9997,N_9226);
and U10932 (N_10932,N_9775,N_9992);
or U10933 (N_10933,N_9316,N_10266);
or U10934 (N_10934,N_10292,N_9424);
xor U10935 (N_10935,N_9987,N_10239);
or U10936 (N_10936,N_9687,N_9071);
nor U10937 (N_10937,N_9512,N_9282);
or U10938 (N_10938,N_10012,N_10360);
nand U10939 (N_10939,N_9067,N_9118);
nand U10940 (N_10940,N_9350,N_10278);
or U10941 (N_10941,N_10174,N_9318);
or U10942 (N_10942,N_10274,N_9031);
xor U10943 (N_10943,N_10260,N_10398);
nand U10944 (N_10944,N_9386,N_10134);
nand U10945 (N_10945,N_10496,N_10191);
xnor U10946 (N_10946,N_9939,N_9330);
and U10947 (N_10947,N_9352,N_10127);
or U10948 (N_10948,N_10452,N_10311);
xnor U10949 (N_10949,N_9606,N_10218);
or U10950 (N_10950,N_10045,N_9619);
or U10951 (N_10951,N_10090,N_9628);
or U10952 (N_10952,N_10455,N_9522);
and U10953 (N_10953,N_9856,N_10437);
nor U10954 (N_10954,N_10414,N_10478);
nand U10955 (N_10955,N_9220,N_9154);
and U10956 (N_10956,N_9417,N_10291);
xnor U10957 (N_10957,N_9266,N_9887);
nand U10958 (N_10958,N_9762,N_10403);
or U10959 (N_10959,N_10298,N_9371);
nor U10960 (N_10960,N_9692,N_9173);
or U10961 (N_10961,N_9600,N_10233);
nand U10962 (N_10962,N_9805,N_9519);
or U10963 (N_10963,N_9707,N_9660);
and U10964 (N_10964,N_9399,N_9240);
nor U10965 (N_10965,N_9027,N_10139);
and U10966 (N_10966,N_9908,N_9255);
and U10967 (N_10967,N_9845,N_9023);
and U10968 (N_10968,N_9094,N_9559);
nor U10969 (N_10969,N_9631,N_10349);
nor U10970 (N_10970,N_9594,N_10050);
or U10971 (N_10971,N_10062,N_9968);
or U10972 (N_10972,N_9507,N_9546);
nand U10973 (N_10973,N_10004,N_9651);
or U10974 (N_10974,N_10216,N_10088);
nor U10975 (N_10975,N_9180,N_10140);
nand U10976 (N_10976,N_9463,N_10057);
nor U10977 (N_10977,N_9286,N_10473);
xor U10978 (N_10978,N_10313,N_10284);
nand U10979 (N_10979,N_10160,N_10318);
and U10980 (N_10980,N_10084,N_9544);
or U10981 (N_10981,N_9198,N_9532);
and U10982 (N_10982,N_10321,N_9288);
xnor U10983 (N_10983,N_9717,N_10126);
xor U10984 (N_10984,N_9040,N_9044);
xor U10985 (N_10985,N_10023,N_9446);
nand U10986 (N_10986,N_9566,N_10109);
or U10987 (N_10987,N_10264,N_9569);
and U10988 (N_10988,N_10471,N_9977);
nand U10989 (N_10989,N_9003,N_9274);
nand U10990 (N_10990,N_9026,N_9903);
xnor U10991 (N_10991,N_9851,N_9760);
or U10992 (N_10992,N_10325,N_10272);
xnor U10993 (N_10993,N_10114,N_9057);
nand U10994 (N_10994,N_9554,N_9837);
xor U10995 (N_10995,N_10064,N_9028);
xnor U10996 (N_10996,N_9864,N_10357);
nand U10997 (N_10997,N_10051,N_9986);
nor U10998 (N_10998,N_9354,N_9614);
xor U10999 (N_10999,N_9847,N_9285);
or U11000 (N_11000,N_9281,N_9825);
nand U11001 (N_11001,N_10221,N_9790);
nor U11002 (N_11002,N_9863,N_9038);
nor U11003 (N_11003,N_9422,N_9780);
nand U11004 (N_11004,N_9323,N_9861);
and U11005 (N_11005,N_10163,N_9106);
or U11006 (N_11006,N_9297,N_10296);
and U11007 (N_11007,N_9377,N_9498);
and U11008 (N_11008,N_10283,N_9796);
nor U11009 (N_11009,N_10449,N_10371);
nor U11010 (N_11010,N_10154,N_9065);
and U11011 (N_11011,N_9474,N_10143);
or U11012 (N_11012,N_9096,N_10192);
nand U11013 (N_11013,N_9082,N_9423);
nand U11014 (N_11014,N_9605,N_9655);
nor U11015 (N_11015,N_9176,N_9344);
xnor U11016 (N_11016,N_10162,N_10132);
or U11017 (N_11017,N_9063,N_9575);
nor U11018 (N_11018,N_9991,N_10487);
nor U11019 (N_11019,N_9141,N_9971);
xnor U11020 (N_11020,N_10161,N_9904);
nand U11021 (N_11021,N_10049,N_9213);
and U11022 (N_11022,N_9918,N_9964);
nand U11023 (N_11023,N_9275,N_9165);
nor U11024 (N_11024,N_10173,N_10495);
or U11025 (N_11025,N_9341,N_10185);
or U11026 (N_11026,N_10068,N_9437);
nor U11027 (N_11027,N_9222,N_10411);
or U11028 (N_11028,N_9645,N_10423);
and U11029 (N_11029,N_10304,N_9913);
xnor U11030 (N_11030,N_10075,N_9767);
xor U11031 (N_11031,N_9192,N_10059);
xnor U11032 (N_11032,N_9454,N_9894);
xnor U11033 (N_11033,N_9066,N_9924);
nand U11034 (N_11034,N_9147,N_10457);
or U11035 (N_11035,N_9311,N_10460);
and U11036 (N_11036,N_9689,N_9680);
or U11037 (N_11037,N_10389,N_10476);
nor U11038 (N_11038,N_10407,N_10079);
nand U11039 (N_11039,N_9459,N_10390);
xor U11040 (N_11040,N_9217,N_9563);
xnor U11041 (N_11041,N_9976,N_9757);
or U11042 (N_11042,N_9107,N_9008);
xnor U11043 (N_11043,N_9900,N_10220);
nand U11044 (N_11044,N_9278,N_9538);
nor U11045 (N_11045,N_10015,N_9754);
and U11046 (N_11046,N_10106,N_9109);
nor U11047 (N_11047,N_9150,N_9111);
nand U11048 (N_11048,N_9586,N_10406);
nor U11049 (N_11049,N_9394,N_9550);
xnor U11050 (N_11050,N_9873,N_10294);
nand U11051 (N_11051,N_10066,N_10249);
and U11052 (N_11052,N_9870,N_10470);
and U11053 (N_11053,N_9353,N_9582);
and U11054 (N_11054,N_10001,N_9700);
or U11055 (N_11055,N_9833,N_9885);
nand U11056 (N_11056,N_10196,N_9159);
nand U11057 (N_11057,N_10385,N_9788);
or U11058 (N_11058,N_9102,N_9187);
nand U11059 (N_11059,N_9138,N_9254);
and U11060 (N_11060,N_10176,N_10111);
nand U11061 (N_11061,N_9091,N_9523);
and U11062 (N_11062,N_9476,N_9945);
xor U11063 (N_11063,N_9841,N_9744);
nand U11064 (N_11064,N_9978,N_10110);
or U11065 (N_11065,N_10427,N_9607);
or U11066 (N_11066,N_9688,N_9897);
xnor U11067 (N_11067,N_9494,N_9553);
and U11068 (N_11068,N_9149,N_9293);
and U11069 (N_11069,N_9130,N_9844);
or U11070 (N_11070,N_9428,N_10120);
or U11071 (N_11071,N_9036,N_9777);
nor U11072 (N_11072,N_9896,N_9105);
and U11073 (N_11073,N_10169,N_9206);
and U11074 (N_11074,N_9539,N_9952);
nand U11075 (N_11075,N_10446,N_9604);
and U11076 (N_11076,N_9398,N_9632);
xor U11077 (N_11077,N_9228,N_10031);
and U11078 (N_11078,N_10312,N_10486);
or U11079 (N_11079,N_9395,N_9998);
and U11080 (N_11080,N_10381,N_10133);
xor U11081 (N_11081,N_10122,N_10424);
and U11082 (N_11082,N_9177,N_10259);
nand U11083 (N_11083,N_9765,N_9970);
xnor U11084 (N_11084,N_9784,N_9869);
nand U11085 (N_11085,N_9838,N_10060);
and U11086 (N_11086,N_9705,N_9639);
nor U11087 (N_11087,N_9009,N_9018);
nand U11088 (N_11088,N_10397,N_9644);
nor U11089 (N_11089,N_9542,N_10301);
nor U11090 (N_11090,N_9186,N_9208);
nor U11091 (N_11091,N_10412,N_10286);
nand U11092 (N_11092,N_9892,N_10401);
and U11093 (N_11093,N_9962,N_9591);
and U11094 (N_11094,N_9260,N_10443);
and U11095 (N_11095,N_9378,N_10206);
or U11096 (N_11096,N_10040,N_9486);
nand U11097 (N_11097,N_9339,N_9079);
nor U11098 (N_11098,N_9721,N_10273);
xnor U11099 (N_11099,N_10246,N_10314);
or U11100 (N_11100,N_9283,N_9360);
xnor U11101 (N_11101,N_10375,N_9418);
and U11102 (N_11102,N_10093,N_10368);
nor U11103 (N_11103,N_10387,N_9218);
nand U11104 (N_11104,N_9390,N_9893);
and U11105 (N_11105,N_9140,N_10188);
and U11106 (N_11106,N_9511,N_9086);
xor U11107 (N_11107,N_9090,N_9899);
or U11108 (N_11108,N_9568,N_10052);
xor U11109 (N_11109,N_9827,N_10047);
and U11110 (N_11110,N_10472,N_10148);
and U11111 (N_11111,N_9013,N_9409);
xnor U11112 (N_11112,N_9444,N_9200);
xnor U11113 (N_11113,N_10186,N_9375);
and U11114 (N_11114,N_10287,N_9294);
xor U11115 (N_11115,N_9385,N_9432);
and U11116 (N_11116,N_10413,N_9010);
xnor U11117 (N_11117,N_9032,N_10095);
xnor U11118 (N_11118,N_10044,N_9840);
nor U11119 (N_11119,N_9905,N_9781);
nor U11120 (N_11120,N_9426,N_9419);
and U11121 (N_11121,N_9324,N_9256);
xnor U11122 (N_11122,N_9265,N_9313);
nor U11123 (N_11123,N_9597,N_9160);
xor U11124 (N_11124,N_9191,N_9679);
nand U11125 (N_11125,N_9473,N_9081);
xnor U11126 (N_11126,N_10223,N_10180);
or U11127 (N_11127,N_9749,N_9491);
nand U11128 (N_11128,N_9571,N_9797);
nor U11129 (N_11129,N_10342,N_10433);
and U11130 (N_11130,N_9960,N_9806);
and U11131 (N_11131,N_9608,N_10450);
xor U11132 (N_11132,N_10254,N_9488);
and U11133 (N_11133,N_9166,N_9975);
nand U11134 (N_11134,N_9931,N_10178);
nor U11135 (N_11135,N_9312,N_10386);
and U11136 (N_11136,N_9736,N_10175);
nor U11137 (N_11137,N_10310,N_9034);
or U11138 (N_11138,N_10419,N_9726);
nor U11139 (N_11139,N_9933,N_9229);
xor U11140 (N_11140,N_9593,N_9201);
or U11141 (N_11141,N_10251,N_9501);
or U11142 (N_11142,N_9670,N_9750);
or U11143 (N_11143,N_10144,N_10200);
xor U11144 (N_11144,N_9890,N_9000);
nor U11145 (N_11145,N_9953,N_9715);
nand U11146 (N_11146,N_9642,N_9708);
nand U11147 (N_11147,N_9387,N_9862);
and U11148 (N_11148,N_9194,N_9938);
or U11149 (N_11149,N_9929,N_9927);
nand U11150 (N_11150,N_10334,N_9703);
nand U11151 (N_11151,N_9188,N_9004);
nand U11152 (N_11152,N_10210,N_10308);
and U11153 (N_11153,N_9460,N_9919);
nand U11154 (N_11154,N_10379,N_9898);
and U11155 (N_11155,N_9070,N_10030);
or U11156 (N_11156,N_10159,N_10405);
and U11157 (N_11157,N_10483,N_9531);
nand U11158 (N_11158,N_9025,N_9565);
and U11159 (N_11159,N_9587,N_10282);
nand U11160 (N_11160,N_10432,N_9536);
xnor U11161 (N_11161,N_9561,N_9663);
nor U11162 (N_11162,N_9355,N_9307);
and U11163 (N_11163,N_9493,N_9835);
and U11164 (N_11164,N_10480,N_9712);
and U11165 (N_11165,N_9271,N_10083);
nor U11166 (N_11166,N_9319,N_9325);
xor U11167 (N_11167,N_9855,N_10002);
or U11168 (N_11168,N_9653,N_10018);
xnor U11169 (N_11169,N_10197,N_9241);
or U11170 (N_11170,N_10253,N_10000);
and U11171 (N_11171,N_10116,N_9759);
xnor U11172 (N_11172,N_9205,N_9362);
nor U11173 (N_11173,N_9789,N_10451);
and U11174 (N_11174,N_9022,N_9732);
nor U11175 (N_11175,N_9029,N_9761);
nand U11176 (N_11176,N_10182,N_9988);
nand U11177 (N_11177,N_10498,N_10324);
or U11178 (N_11178,N_9947,N_9499);
nand U11179 (N_11179,N_10164,N_9143);
nand U11180 (N_11180,N_10245,N_10370);
nor U11181 (N_11181,N_9139,N_10288);
nor U11182 (N_11182,N_9305,N_9131);
nor U11183 (N_11183,N_10010,N_10211);
xnor U11184 (N_11184,N_10199,N_9095);
or U11185 (N_11185,N_10219,N_9433);
nor U11186 (N_11186,N_9596,N_9958);
xor U11187 (N_11187,N_9720,N_9853);
or U11188 (N_11188,N_10285,N_10119);
and U11189 (N_11189,N_10034,N_9058);
nand U11190 (N_11190,N_10252,N_10477);
and U11191 (N_11191,N_10435,N_10157);
or U11192 (N_11192,N_9826,N_9778);
nor U11193 (N_11193,N_9768,N_10136);
or U11194 (N_11194,N_9996,N_9503);
and U11195 (N_11195,N_10026,N_10481);
nand U11196 (N_11196,N_9306,N_10404);
or U11197 (N_11197,N_9322,N_9334);
nor U11198 (N_11198,N_10422,N_10124);
nor U11199 (N_11199,N_9654,N_9268);
or U11200 (N_11200,N_10400,N_9335);
and U11201 (N_11201,N_10224,N_9506);
and U11202 (N_11202,N_9940,N_9244);
nor U11203 (N_11203,N_9169,N_10328);
or U11204 (N_11204,N_9233,N_10146);
xnor U11205 (N_11205,N_9911,N_9302);
or U11206 (N_11206,N_10226,N_9144);
xnor U11207 (N_11207,N_10019,N_10366);
or U11208 (N_11208,N_10069,N_10020);
or U11209 (N_11209,N_10332,N_9932);
or U11210 (N_11210,N_9737,N_10236);
nand U11211 (N_11211,N_9092,N_9518);
and U11212 (N_11212,N_9061,N_9558);
nand U11213 (N_11213,N_9012,N_10183);
nor U11214 (N_11214,N_10073,N_10441);
nor U11215 (N_11215,N_9580,N_9802);
xnor U11216 (N_11216,N_9613,N_10399);
or U11217 (N_11217,N_9673,N_9338);
nor U11218 (N_11218,N_9701,N_10240);
and U11219 (N_11219,N_9906,N_9403);
or U11220 (N_11220,N_10279,N_9965);
xnor U11221 (N_11221,N_9537,N_10499);
nor U11222 (N_11222,N_9115,N_9646);
nor U11223 (N_11223,N_10442,N_9479);
and U11224 (N_11224,N_9178,N_10343);
nand U11225 (N_11225,N_10097,N_9336);
or U11226 (N_11226,N_9785,N_10281);
nor U11227 (N_11227,N_9963,N_10170);
nor U11228 (N_11228,N_9223,N_9054);
xor U11229 (N_11229,N_10077,N_9891);
xnor U11230 (N_11230,N_9752,N_10037);
or U11231 (N_11231,N_10420,N_9219);
nor U11232 (N_11232,N_9615,N_9935);
and U11233 (N_11233,N_10082,N_9020);
and U11234 (N_11234,N_10453,N_10244);
and U11235 (N_11235,N_9601,N_9055);
or U11236 (N_11236,N_9033,N_10395);
nor U11237 (N_11237,N_10033,N_10494);
nor U11238 (N_11238,N_9883,N_9037);
nor U11239 (N_11239,N_10458,N_9973);
and U11240 (N_11240,N_9972,N_9381);
xor U11241 (N_11241,N_10041,N_9922);
xnor U11242 (N_11242,N_9153,N_9738);
xor U11243 (N_11243,N_9747,N_9461);
or U11244 (N_11244,N_9317,N_9909);
xor U11245 (N_11245,N_9727,N_9995);
and U11246 (N_11246,N_10491,N_10061);
and U11247 (N_11247,N_9137,N_9019);
nand U11248 (N_11248,N_10227,N_9224);
xor U11249 (N_11249,N_9951,N_9182);
and U11250 (N_11250,N_9185,N_9148);
nor U11251 (N_11251,N_10008,N_9069);
nor U11252 (N_11252,N_9134,N_10132);
nand U11253 (N_11253,N_9165,N_9815);
nor U11254 (N_11254,N_9848,N_10122);
xnor U11255 (N_11255,N_10236,N_9444);
or U11256 (N_11256,N_9757,N_9127);
nand U11257 (N_11257,N_9343,N_9191);
nand U11258 (N_11258,N_9017,N_10323);
and U11259 (N_11259,N_9825,N_9740);
or U11260 (N_11260,N_10055,N_10433);
nor U11261 (N_11261,N_9660,N_10264);
and U11262 (N_11262,N_10065,N_10105);
or U11263 (N_11263,N_10395,N_9277);
or U11264 (N_11264,N_9499,N_9445);
or U11265 (N_11265,N_10383,N_10229);
nand U11266 (N_11266,N_10426,N_9240);
and U11267 (N_11267,N_9378,N_9581);
nand U11268 (N_11268,N_9161,N_9764);
or U11269 (N_11269,N_9186,N_9172);
or U11270 (N_11270,N_10257,N_9661);
nor U11271 (N_11271,N_9478,N_10375);
nand U11272 (N_11272,N_10065,N_9374);
and U11273 (N_11273,N_10454,N_10055);
nand U11274 (N_11274,N_10129,N_9750);
nand U11275 (N_11275,N_9525,N_10004);
and U11276 (N_11276,N_9079,N_9065);
nor U11277 (N_11277,N_10096,N_10056);
nand U11278 (N_11278,N_9165,N_9960);
xnor U11279 (N_11279,N_9298,N_9591);
and U11280 (N_11280,N_9118,N_9862);
and U11281 (N_11281,N_9117,N_9759);
nor U11282 (N_11282,N_9155,N_10106);
nor U11283 (N_11283,N_9527,N_9733);
and U11284 (N_11284,N_9655,N_10354);
or U11285 (N_11285,N_9882,N_10248);
xnor U11286 (N_11286,N_9237,N_9994);
nor U11287 (N_11287,N_10351,N_9714);
nand U11288 (N_11288,N_10239,N_9662);
and U11289 (N_11289,N_9906,N_9617);
and U11290 (N_11290,N_9525,N_10352);
xnor U11291 (N_11291,N_9157,N_9078);
xnor U11292 (N_11292,N_9084,N_9042);
nor U11293 (N_11293,N_10074,N_9203);
and U11294 (N_11294,N_9826,N_10186);
or U11295 (N_11295,N_9395,N_9045);
nor U11296 (N_11296,N_9987,N_10414);
xor U11297 (N_11297,N_9763,N_10159);
xnor U11298 (N_11298,N_9184,N_9072);
nor U11299 (N_11299,N_10395,N_9270);
xnor U11300 (N_11300,N_10120,N_10228);
nor U11301 (N_11301,N_9254,N_10314);
nand U11302 (N_11302,N_10180,N_9933);
nand U11303 (N_11303,N_9407,N_9186);
nor U11304 (N_11304,N_10445,N_9076);
nor U11305 (N_11305,N_9163,N_9957);
nor U11306 (N_11306,N_9603,N_9358);
or U11307 (N_11307,N_9165,N_9623);
nand U11308 (N_11308,N_9533,N_10252);
or U11309 (N_11309,N_10387,N_9516);
or U11310 (N_11310,N_9782,N_9278);
nor U11311 (N_11311,N_9411,N_10178);
nor U11312 (N_11312,N_10479,N_10385);
or U11313 (N_11313,N_9682,N_9796);
or U11314 (N_11314,N_10240,N_9495);
or U11315 (N_11315,N_9881,N_10061);
or U11316 (N_11316,N_9826,N_9898);
nor U11317 (N_11317,N_10342,N_9499);
or U11318 (N_11318,N_9076,N_10104);
xor U11319 (N_11319,N_9104,N_9809);
nor U11320 (N_11320,N_10134,N_9052);
or U11321 (N_11321,N_9154,N_9407);
and U11322 (N_11322,N_10111,N_10068);
xor U11323 (N_11323,N_9494,N_9236);
and U11324 (N_11324,N_9527,N_9703);
xor U11325 (N_11325,N_9797,N_9543);
and U11326 (N_11326,N_10204,N_9891);
nor U11327 (N_11327,N_9689,N_9665);
or U11328 (N_11328,N_9015,N_10399);
nor U11329 (N_11329,N_9936,N_9911);
or U11330 (N_11330,N_9123,N_9806);
and U11331 (N_11331,N_9277,N_9077);
or U11332 (N_11332,N_9403,N_9760);
xor U11333 (N_11333,N_9856,N_9818);
nand U11334 (N_11334,N_9951,N_9381);
nor U11335 (N_11335,N_9030,N_9020);
and U11336 (N_11336,N_9448,N_10313);
nand U11337 (N_11337,N_9629,N_9877);
and U11338 (N_11338,N_9888,N_9214);
xnor U11339 (N_11339,N_9639,N_9108);
xnor U11340 (N_11340,N_9011,N_9220);
xnor U11341 (N_11341,N_9019,N_10344);
nand U11342 (N_11342,N_10080,N_9471);
and U11343 (N_11343,N_10267,N_9964);
xnor U11344 (N_11344,N_9884,N_9591);
nand U11345 (N_11345,N_10036,N_9850);
nor U11346 (N_11346,N_9833,N_9089);
and U11347 (N_11347,N_9195,N_9427);
xnor U11348 (N_11348,N_9258,N_9118);
or U11349 (N_11349,N_9783,N_9992);
xor U11350 (N_11350,N_10356,N_10205);
xnor U11351 (N_11351,N_9476,N_9761);
or U11352 (N_11352,N_9689,N_9042);
and U11353 (N_11353,N_9348,N_9565);
nor U11354 (N_11354,N_9176,N_9317);
or U11355 (N_11355,N_10275,N_9738);
nor U11356 (N_11356,N_10012,N_9763);
nor U11357 (N_11357,N_10149,N_9968);
xnor U11358 (N_11358,N_10462,N_10397);
and U11359 (N_11359,N_9402,N_9714);
or U11360 (N_11360,N_10473,N_9948);
or U11361 (N_11361,N_9206,N_9115);
and U11362 (N_11362,N_10462,N_9416);
and U11363 (N_11363,N_10082,N_10409);
nand U11364 (N_11364,N_10483,N_9908);
nand U11365 (N_11365,N_10365,N_9922);
or U11366 (N_11366,N_9578,N_9296);
or U11367 (N_11367,N_9293,N_9014);
nand U11368 (N_11368,N_9328,N_9586);
xor U11369 (N_11369,N_10164,N_9888);
nor U11370 (N_11370,N_9542,N_9469);
nor U11371 (N_11371,N_9538,N_9416);
or U11372 (N_11372,N_9514,N_9663);
nor U11373 (N_11373,N_10327,N_10223);
xor U11374 (N_11374,N_10348,N_9110);
nand U11375 (N_11375,N_9988,N_9314);
nor U11376 (N_11376,N_10445,N_10312);
nor U11377 (N_11377,N_9506,N_10410);
nand U11378 (N_11378,N_9108,N_9049);
nand U11379 (N_11379,N_10438,N_9459);
nor U11380 (N_11380,N_10268,N_10103);
nand U11381 (N_11381,N_9706,N_9595);
xor U11382 (N_11382,N_9552,N_9184);
and U11383 (N_11383,N_10459,N_10212);
or U11384 (N_11384,N_9724,N_9084);
nand U11385 (N_11385,N_10308,N_10194);
and U11386 (N_11386,N_10061,N_9504);
nand U11387 (N_11387,N_10268,N_9453);
nor U11388 (N_11388,N_10459,N_10158);
nor U11389 (N_11389,N_9257,N_9206);
and U11390 (N_11390,N_9849,N_9701);
and U11391 (N_11391,N_9184,N_9948);
nand U11392 (N_11392,N_10085,N_10019);
and U11393 (N_11393,N_9430,N_9873);
nand U11394 (N_11394,N_9249,N_10431);
and U11395 (N_11395,N_9716,N_9330);
xor U11396 (N_11396,N_10443,N_9733);
xor U11397 (N_11397,N_9740,N_9442);
nor U11398 (N_11398,N_10377,N_10324);
nor U11399 (N_11399,N_10301,N_10032);
or U11400 (N_11400,N_9643,N_9433);
nand U11401 (N_11401,N_10083,N_10263);
nor U11402 (N_11402,N_9757,N_10433);
xor U11403 (N_11403,N_10311,N_10355);
xnor U11404 (N_11404,N_10201,N_10063);
nor U11405 (N_11405,N_9640,N_9936);
and U11406 (N_11406,N_9293,N_9710);
nand U11407 (N_11407,N_10268,N_10043);
nand U11408 (N_11408,N_10155,N_9581);
and U11409 (N_11409,N_9306,N_10157);
xor U11410 (N_11410,N_9256,N_9280);
or U11411 (N_11411,N_10351,N_9260);
nand U11412 (N_11412,N_9202,N_10235);
or U11413 (N_11413,N_10165,N_10263);
or U11414 (N_11414,N_9697,N_10210);
nand U11415 (N_11415,N_9300,N_10143);
nand U11416 (N_11416,N_10333,N_9822);
nor U11417 (N_11417,N_9959,N_9592);
nand U11418 (N_11418,N_10225,N_9563);
xor U11419 (N_11419,N_9141,N_9446);
and U11420 (N_11420,N_9311,N_10183);
nor U11421 (N_11421,N_9081,N_9113);
nor U11422 (N_11422,N_9944,N_10290);
xnor U11423 (N_11423,N_9931,N_9690);
nand U11424 (N_11424,N_9724,N_9457);
nand U11425 (N_11425,N_9920,N_9333);
xnor U11426 (N_11426,N_10225,N_9258);
nand U11427 (N_11427,N_9929,N_9588);
xnor U11428 (N_11428,N_10477,N_9801);
or U11429 (N_11429,N_9841,N_9500);
or U11430 (N_11430,N_10495,N_10029);
and U11431 (N_11431,N_10475,N_9749);
and U11432 (N_11432,N_10137,N_9076);
xor U11433 (N_11433,N_10236,N_9230);
nand U11434 (N_11434,N_9126,N_10435);
or U11435 (N_11435,N_9033,N_9393);
nor U11436 (N_11436,N_9785,N_10172);
and U11437 (N_11437,N_10107,N_9502);
nor U11438 (N_11438,N_9360,N_9889);
nand U11439 (N_11439,N_9770,N_10187);
or U11440 (N_11440,N_10175,N_10180);
and U11441 (N_11441,N_9748,N_9143);
or U11442 (N_11442,N_9442,N_9181);
xor U11443 (N_11443,N_10306,N_9273);
xnor U11444 (N_11444,N_9352,N_9808);
or U11445 (N_11445,N_10491,N_9030);
and U11446 (N_11446,N_9998,N_9977);
or U11447 (N_11447,N_10229,N_9309);
nand U11448 (N_11448,N_9744,N_9168);
nor U11449 (N_11449,N_9496,N_9331);
nand U11450 (N_11450,N_9419,N_9509);
nor U11451 (N_11451,N_10168,N_9323);
or U11452 (N_11452,N_9591,N_9676);
or U11453 (N_11453,N_9091,N_9253);
nand U11454 (N_11454,N_10133,N_9180);
and U11455 (N_11455,N_9184,N_9882);
xor U11456 (N_11456,N_9428,N_9615);
xor U11457 (N_11457,N_10456,N_9249);
xnor U11458 (N_11458,N_10251,N_9358);
nand U11459 (N_11459,N_10422,N_9440);
xnor U11460 (N_11460,N_9123,N_10248);
nor U11461 (N_11461,N_9297,N_9390);
and U11462 (N_11462,N_9116,N_10434);
and U11463 (N_11463,N_9257,N_9875);
and U11464 (N_11464,N_9384,N_9029);
nor U11465 (N_11465,N_9722,N_9154);
nand U11466 (N_11466,N_9574,N_10209);
nand U11467 (N_11467,N_9109,N_9302);
xnor U11468 (N_11468,N_9912,N_9399);
nor U11469 (N_11469,N_9905,N_10387);
nand U11470 (N_11470,N_9802,N_9891);
nand U11471 (N_11471,N_10178,N_9510);
xnor U11472 (N_11472,N_10431,N_9283);
nand U11473 (N_11473,N_9659,N_9908);
or U11474 (N_11474,N_9045,N_10225);
nand U11475 (N_11475,N_9114,N_9398);
nor U11476 (N_11476,N_10342,N_9835);
and U11477 (N_11477,N_10255,N_9945);
xor U11478 (N_11478,N_10293,N_9019);
or U11479 (N_11479,N_9302,N_9623);
xor U11480 (N_11480,N_10439,N_9638);
and U11481 (N_11481,N_9562,N_9285);
or U11482 (N_11482,N_9214,N_9612);
xnor U11483 (N_11483,N_10048,N_9615);
xnor U11484 (N_11484,N_9525,N_10255);
and U11485 (N_11485,N_9021,N_9309);
nand U11486 (N_11486,N_9559,N_10352);
xor U11487 (N_11487,N_9864,N_9145);
nor U11488 (N_11488,N_9112,N_10478);
nand U11489 (N_11489,N_9242,N_10402);
nor U11490 (N_11490,N_9249,N_10306);
nor U11491 (N_11491,N_10442,N_10482);
or U11492 (N_11492,N_9453,N_10183);
nor U11493 (N_11493,N_9684,N_10010);
or U11494 (N_11494,N_9649,N_10042);
nand U11495 (N_11495,N_9086,N_9514);
nor U11496 (N_11496,N_9036,N_10457);
xnor U11497 (N_11497,N_9859,N_9720);
nand U11498 (N_11498,N_10211,N_9384);
and U11499 (N_11499,N_9391,N_9080);
nor U11500 (N_11500,N_10269,N_10489);
xnor U11501 (N_11501,N_10084,N_9407);
and U11502 (N_11502,N_9552,N_9864);
xnor U11503 (N_11503,N_10312,N_10263);
or U11504 (N_11504,N_9997,N_9363);
and U11505 (N_11505,N_9614,N_9829);
nand U11506 (N_11506,N_9917,N_9003);
nor U11507 (N_11507,N_10053,N_10206);
and U11508 (N_11508,N_9170,N_9357);
and U11509 (N_11509,N_9256,N_10482);
or U11510 (N_11510,N_9252,N_10479);
xor U11511 (N_11511,N_9130,N_9418);
or U11512 (N_11512,N_9096,N_9690);
and U11513 (N_11513,N_9969,N_10312);
or U11514 (N_11514,N_10370,N_9385);
or U11515 (N_11515,N_9708,N_10197);
xor U11516 (N_11516,N_9097,N_10095);
nor U11517 (N_11517,N_10025,N_9994);
and U11518 (N_11518,N_9410,N_9296);
and U11519 (N_11519,N_9625,N_9376);
xor U11520 (N_11520,N_9009,N_9970);
xor U11521 (N_11521,N_10419,N_10016);
nand U11522 (N_11522,N_9167,N_10472);
nor U11523 (N_11523,N_9498,N_9666);
nor U11524 (N_11524,N_9172,N_9003);
or U11525 (N_11525,N_9074,N_10007);
xor U11526 (N_11526,N_9629,N_9825);
and U11527 (N_11527,N_9426,N_9970);
and U11528 (N_11528,N_10300,N_10301);
or U11529 (N_11529,N_10012,N_9699);
nor U11530 (N_11530,N_9751,N_9427);
nand U11531 (N_11531,N_10042,N_9699);
or U11532 (N_11532,N_10043,N_10059);
nor U11533 (N_11533,N_10029,N_9125);
and U11534 (N_11534,N_10300,N_9288);
or U11535 (N_11535,N_10156,N_10056);
nor U11536 (N_11536,N_9959,N_9671);
nand U11537 (N_11537,N_10386,N_9467);
or U11538 (N_11538,N_10464,N_9436);
and U11539 (N_11539,N_9027,N_9278);
or U11540 (N_11540,N_9720,N_9602);
nand U11541 (N_11541,N_9317,N_10396);
xnor U11542 (N_11542,N_9345,N_9337);
xor U11543 (N_11543,N_9436,N_9284);
or U11544 (N_11544,N_9516,N_9633);
nor U11545 (N_11545,N_9164,N_9433);
nor U11546 (N_11546,N_9847,N_9410);
nor U11547 (N_11547,N_9721,N_9655);
and U11548 (N_11548,N_10096,N_9364);
xnor U11549 (N_11549,N_10086,N_9670);
and U11550 (N_11550,N_10107,N_9821);
xor U11551 (N_11551,N_9641,N_9563);
xor U11552 (N_11552,N_9713,N_9274);
or U11553 (N_11553,N_9461,N_10100);
nor U11554 (N_11554,N_9325,N_9666);
nand U11555 (N_11555,N_9520,N_9029);
nand U11556 (N_11556,N_9455,N_10255);
or U11557 (N_11557,N_9901,N_10441);
xor U11558 (N_11558,N_10165,N_9737);
xor U11559 (N_11559,N_9016,N_10435);
or U11560 (N_11560,N_10362,N_10194);
nand U11561 (N_11561,N_9388,N_10133);
or U11562 (N_11562,N_9783,N_9321);
and U11563 (N_11563,N_10202,N_10441);
and U11564 (N_11564,N_9091,N_9264);
nand U11565 (N_11565,N_9639,N_9372);
xor U11566 (N_11566,N_9653,N_9818);
xor U11567 (N_11567,N_10038,N_9565);
xor U11568 (N_11568,N_9532,N_9278);
nand U11569 (N_11569,N_9639,N_9002);
xor U11570 (N_11570,N_9021,N_10423);
or U11571 (N_11571,N_9841,N_10130);
or U11572 (N_11572,N_10297,N_9544);
and U11573 (N_11573,N_10054,N_9435);
and U11574 (N_11574,N_9432,N_10104);
nand U11575 (N_11575,N_10485,N_9038);
or U11576 (N_11576,N_10090,N_9578);
or U11577 (N_11577,N_9836,N_9004);
xor U11578 (N_11578,N_9457,N_9526);
xor U11579 (N_11579,N_9945,N_10469);
or U11580 (N_11580,N_10274,N_10052);
and U11581 (N_11581,N_9124,N_9119);
xnor U11582 (N_11582,N_10054,N_9736);
nor U11583 (N_11583,N_10070,N_10498);
nand U11584 (N_11584,N_10325,N_9740);
and U11585 (N_11585,N_9640,N_9698);
nand U11586 (N_11586,N_9279,N_9433);
xor U11587 (N_11587,N_9226,N_10462);
or U11588 (N_11588,N_9976,N_9936);
and U11589 (N_11589,N_10198,N_9193);
xor U11590 (N_11590,N_9441,N_9571);
or U11591 (N_11591,N_9550,N_10056);
xor U11592 (N_11592,N_9151,N_10214);
or U11593 (N_11593,N_9782,N_9807);
nand U11594 (N_11594,N_10081,N_9740);
nor U11595 (N_11595,N_9750,N_10273);
nor U11596 (N_11596,N_10426,N_9299);
xnor U11597 (N_11597,N_10471,N_9022);
and U11598 (N_11598,N_10417,N_10299);
nor U11599 (N_11599,N_9772,N_10362);
and U11600 (N_11600,N_9092,N_9903);
and U11601 (N_11601,N_9513,N_10183);
nand U11602 (N_11602,N_9670,N_9719);
and U11603 (N_11603,N_9611,N_10424);
and U11604 (N_11604,N_9416,N_9976);
and U11605 (N_11605,N_9889,N_9551);
and U11606 (N_11606,N_9377,N_10004);
xnor U11607 (N_11607,N_10139,N_10429);
and U11608 (N_11608,N_9269,N_9073);
and U11609 (N_11609,N_10442,N_9028);
xor U11610 (N_11610,N_10387,N_9893);
or U11611 (N_11611,N_10156,N_9964);
and U11612 (N_11612,N_9620,N_9793);
xnor U11613 (N_11613,N_9047,N_9055);
nor U11614 (N_11614,N_9300,N_10006);
xnor U11615 (N_11615,N_10111,N_9116);
nand U11616 (N_11616,N_9958,N_9919);
nor U11617 (N_11617,N_10167,N_10291);
xor U11618 (N_11618,N_9660,N_10290);
and U11619 (N_11619,N_10099,N_10268);
xor U11620 (N_11620,N_10240,N_9954);
and U11621 (N_11621,N_9603,N_9730);
nor U11622 (N_11622,N_9574,N_10175);
nor U11623 (N_11623,N_9053,N_9951);
or U11624 (N_11624,N_9520,N_9861);
nor U11625 (N_11625,N_10098,N_9297);
nand U11626 (N_11626,N_10156,N_10472);
and U11627 (N_11627,N_10388,N_10250);
or U11628 (N_11628,N_9833,N_9920);
nand U11629 (N_11629,N_9879,N_9385);
nand U11630 (N_11630,N_9243,N_10192);
or U11631 (N_11631,N_10095,N_10252);
and U11632 (N_11632,N_10433,N_10093);
or U11633 (N_11633,N_10227,N_9774);
or U11634 (N_11634,N_10035,N_10369);
nor U11635 (N_11635,N_9657,N_9923);
and U11636 (N_11636,N_9935,N_9749);
xor U11637 (N_11637,N_9550,N_10352);
xnor U11638 (N_11638,N_9300,N_9506);
and U11639 (N_11639,N_10172,N_9028);
xor U11640 (N_11640,N_9438,N_9025);
nand U11641 (N_11641,N_9603,N_9770);
and U11642 (N_11642,N_9003,N_10481);
xnor U11643 (N_11643,N_9379,N_10097);
xnor U11644 (N_11644,N_9636,N_10454);
nor U11645 (N_11645,N_9368,N_9340);
nor U11646 (N_11646,N_10283,N_9985);
nand U11647 (N_11647,N_9489,N_9349);
xnor U11648 (N_11648,N_9982,N_10467);
or U11649 (N_11649,N_9153,N_9428);
or U11650 (N_11650,N_9220,N_9288);
nor U11651 (N_11651,N_10397,N_10071);
xnor U11652 (N_11652,N_10463,N_10192);
and U11653 (N_11653,N_9154,N_10414);
and U11654 (N_11654,N_9379,N_9630);
and U11655 (N_11655,N_9800,N_10113);
nor U11656 (N_11656,N_9765,N_9339);
or U11657 (N_11657,N_9886,N_10224);
and U11658 (N_11658,N_10078,N_9774);
nor U11659 (N_11659,N_9390,N_9344);
xor U11660 (N_11660,N_10489,N_9792);
or U11661 (N_11661,N_10438,N_9807);
or U11662 (N_11662,N_9012,N_9040);
xor U11663 (N_11663,N_9339,N_9327);
xor U11664 (N_11664,N_9158,N_9753);
nand U11665 (N_11665,N_9979,N_10386);
nor U11666 (N_11666,N_9712,N_9402);
and U11667 (N_11667,N_9901,N_9971);
nor U11668 (N_11668,N_9389,N_9288);
xnor U11669 (N_11669,N_9964,N_10170);
or U11670 (N_11670,N_9712,N_10119);
xnor U11671 (N_11671,N_9882,N_10066);
and U11672 (N_11672,N_9951,N_10356);
nor U11673 (N_11673,N_9939,N_9415);
or U11674 (N_11674,N_9786,N_9683);
nor U11675 (N_11675,N_9338,N_9393);
nand U11676 (N_11676,N_10263,N_9081);
xnor U11677 (N_11677,N_10200,N_9378);
nor U11678 (N_11678,N_9903,N_9762);
xnor U11679 (N_11679,N_9028,N_9820);
xor U11680 (N_11680,N_9209,N_9908);
nor U11681 (N_11681,N_9902,N_9113);
nand U11682 (N_11682,N_9019,N_10282);
and U11683 (N_11683,N_9369,N_10430);
nor U11684 (N_11684,N_10156,N_9637);
xnor U11685 (N_11685,N_9791,N_10317);
or U11686 (N_11686,N_9432,N_9274);
and U11687 (N_11687,N_10137,N_9869);
xor U11688 (N_11688,N_10071,N_9747);
or U11689 (N_11689,N_9022,N_9921);
or U11690 (N_11690,N_9389,N_10361);
or U11691 (N_11691,N_9913,N_10195);
nor U11692 (N_11692,N_10472,N_9339);
nand U11693 (N_11693,N_9914,N_9459);
nand U11694 (N_11694,N_9694,N_9479);
xnor U11695 (N_11695,N_10099,N_10481);
xnor U11696 (N_11696,N_9785,N_9840);
or U11697 (N_11697,N_9042,N_9119);
nor U11698 (N_11698,N_9663,N_10310);
and U11699 (N_11699,N_9000,N_9788);
nor U11700 (N_11700,N_10057,N_9304);
nor U11701 (N_11701,N_9091,N_9737);
xor U11702 (N_11702,N_9879,N_9084);
nand U11703 (N_11703,N_10067,N_10387);
xnor U11704 (N_11704,N_10180,N_9804);
nand U11705 (N_11705,N_9638,N_9890);
xnor U11706 (N_11706,N_9287,N_9930);
nand U11707 (N_11707,N_10434,N_10046);
xor U11708 (N_11708,N_9612,N_9909);
xor U11709 (N_11709,N_9668,N_9568);
xnor U11710 (N_11710,N_9802,N_9660);
nor U11711 (N_11711,N_10251,N_9913);
and U11712 (N_11712,N_10072,N_9834);
or U11713 (N_11713,N_9139,N_9189);
nor U11714 (N_11714,N_9193,N_9606);
nand U11715 (N_11715,N_9648,N_9510);
nand U11716 (N_11716,N_9197,N_9681);
nor U11717 (N_11717,N_9842,N_9215);
and U11718 (N_11718,N_9747,N_9116);
nand U11719 (N_11719,N_10179,N_9333);
xor U11720 (N_11720,N_9425,N_9500);
nor U11721 (N_11721,N_9752,N_10125);
and U11722 (N_11722,N_9116,N_10219);
nor U11723 (N_11723,N_9149,N_9840);
xnor U11724 (N_11724,N_9500,N_9951);
nand U11725 (N_11725,N_9270,N_9277);
nand U11726 (N_11726,N_9312,N_9173);
nor U11727 (N_11727,N_9971,N_9704);
and U11728 (N_11728,N_10100,N_9078);
and U11729 (N_11729,N_10232,N_9144);
nand U11730 (N_11730,N_10241,N_10080);
xnor U11731 (N_11731,N_10136,N_9323);
or U11732 (N_11732,N_9210,N_10343);
and U11733 (N_11733,N_10472,N_9161);
or U11734 (N_11734,N_9814,N_9948);
nor U11735 (N_11735,N_9647,N_9856);
and U11736 (N_11736,N_10050,N_10392);
nor U11737 (N_11737,N_9617,N_9461);
and U11738 (N_11738,N_10330,N_9318);
nand U11739 (N_11739,N_9988,N_10064);
xnor U11740 (N_11740,N_10197,N_9477);
and U11741 (N_11741,N_9242,N_10386);
nand U11742 (N_11742,N_9610,N_9569);
nor U11743 (N_11743,N_9374,N_9384);
nor U11744 (N_11744,N_10396,N_10265);
nand U11745 (N_11745,N_9206,N_9754);
and U11746 (N_11746,N_9379,N_9248);
or U11747 (N_11747,N_9712,N_10172);
nand U11748 (N_11748,N_9393,N_9537);
or U11749 (N_11749,N_10222,N_10290);
xnor U11750 (N_11750,N_10129,N_10424);
nand U11751 (N_11751,N_9178,N_9762);
nor U11752 (N_11752,N_9222,N_10378);
nand U11753 (N_11753,N_9208,N_10235);
xor U11754 (N_11754,N_10180,N_9139);
nor U11755 (N_11755,N_10345,N_10134);
nor U11756 (N_11756,N_10420,N_9575);
nand U11757 (N_11757,N_10160,N_9985);
and U11758 (N_11758,N_10092,N_9949);
nor U11759 (N_11759,N_9452,N_10205);
or U11760 (N_11760,N_10259,N_9162);
and U11761 (N_11761,N_9379,N_10300);
or U11762 (N_11762,N_9791,N_9255);
xnor U11763 (N_11763,N_9943,N_9198);
nor U11764 (N_11764,N_9257,N_10452);
nand U11765 (N_11765,N_10351,N_9339);
nor U11766 (N_11766,N_9313,N_10055);
or U11767 (N_11767,N_10087,N_9451);
and U11768 (N_11768,N_9427,N_9780);
and U11769 (N_11769,N_9580,N_9374);
nor U11770 (N_11770,N_9015,N_9773);
nor U11771 (N_11771,N_9594,N_9831);
or U11772 (N_11772,N_9454,N_9526);
or U11773 (N_11773,N_9476,N_9187);
or U11774 (N_11774,N_10281,N_9981);
and U11775 (N_11775,N_9645,N_9198);
or U11776 (N_11776,N_10412,N_10065);
nand U11777 (N_11777,N_9249,N_9422);
or U11778 (N_11778,N_10004,N_9301);
or U11779 (N_11779,N_9245,N_10255);
nand U11780 (N_11780,N_10351,N_9132);
nand U11781 (N_11781,N_9629,N_9321);
xor U11782 (N_11782,N_9506,N_9399);
nand U11783 (N_11783,N_9048,N_9320);
or U11784 (N_11784,N_10151,N_9240);
nor U11785 (N_11785,N_10488,N_10122);
and U11786 (N_11786,N_9511,N_9179);
and U11787 (N_11787,N_9274,N_9371);
and U11788 (N_11788,N_9709,N_10499);
nor U11789 (N_11789,N_10493,N_10230);
and U11790 (N_11790,N_9171,N_10427);
or U11791 (N_11791,N_10182,N_9193);
xor U11792 (N_11792,N_9759,N_9453);
or U11793 (N_11793,N_9073,N_10467);
nor U11794 (N_11794,N_9656,N_10444);
nor U11795 (N_11795,N_9623,N_9292);
nor U11796 (N_11796,N_9065,N_9560);
nand U11797 (N_11797,N_10358,N_10438);
or U11798 (N_11798,N_9148,N_9237);
and U11799 (N_11799,N_9530,N_10387);
nor U11800 (N_11800,N_9187,N_10265);
xor U11801 (N_11801,N_10153,N_9839);
xor U11802 (N_11802,N_9875,N_9077);
and U11803 (N_11803,N_9909,N_9967);
or U11804 (N_11804,N_9337,N_9877);
and U11805 (N_11805,N_9611,N_9780);
or U11806 (N_11806,N_9533,N_10216);
nor U11807 (N_11807,N_9839,N_9622);
nand U11808 (N_11808,N_10233,N_10244);
nand U11809 (N_11809,N_10190,N_10422);
nand U11810 (N_11810,N_9903,N_10303);
and U11811 (N_11811,N_9326,N_9102);
xnor U11812 (N_11812,N_9272,N_10107);
xnor U11813 (N_11813,N_9896,N_9296);
nand U11814 (N_11814,N_9881,N_9761);
xor U11815 (N_11815,N_9271,N_9539);
nand U11816 (N_11816,N_10346,N_10425);
nor U11817 (N_11817,N_9045,N_9194);
nor U11818 (N_11818,N_9551,N_9175);
or U11819 (N_11819,N_9906,N_9216);
nand U11820 (N_11820,N_9673,N_10150);
and U11821 (N_11821,N_10263,N_9177);
nand U11822 (N_11822,N_9675,N_10335);
nor U11823 (N_11823,N_10147,N_10293);
nand U11824 (N_11824,N_9685,N_9044);
or U11825 (N_11825,N_9870,N_10156);
nor U11826 (N_11826,N_9337,N_9796);
and U11827 (N_11827,N_9909,N_9478);
xor U11828 (N_11828,N_10449,N_10271);
nand U11829 (N_11829,N_9385,N_9112);
xnor U11830 (N_11830,N_9818,N_9946);
nor U11831 (N_11831,N_9418,N_10490);
xnor U11832 (N_11832,N_9433,N_10250);
nor U11833 (N_11833,N_10323,N_9963);
nand U11834 (N_11834,N_10250,N_9919);
xnor U11835 (N_11835,N_9731,N_9576);
and U11836 (N_11836,N_10452,N_9016);
nor U11837 (N_11837,N_10256,N_9593);
and U11838 (N_11838,N_9031,N_9263);
xor U11839 (N_11839,N_10300,N_9822);
xor U11840 (N_11840,N_9363,N_9941);
or U11841 (N_11841,N_9643,N_10075);
nor U11842 (N_11842,N_10008,N_10442);
and U11843 (N_11843,N_10056,N_10276);
nand U11844 (N_11844,N_10276,N_9460);
or U11845 (N_11845,N_9819,N_9297);
or U11846 (N_11846,N_9116,N_9547);
or U11847 (N_11847,N_10139,N_10401);
xor U11848 (N_11848,N_9109,N_9970);
and U11849 (N_11849,N_9837,N_10138);
or U11850 (N_11850,N_10496,N_10056);
xnor U11851 (N_11851,N_9585,N_9346);
and U11852 (N_11852,N_10399,N_9701);
nor U11853 (N_11853,N_9508,N_10265);
or U11854 (N_11854,N_9386,N_9875);
xnor U11855 (N_11855,N_10407,N_9705);
nand U11856 (N_11856,N_9987,N_9772);
nand U11857 (N_11857,N_9198,N_9097);
nor U11858 (N_11858,N_9353,N_9248);
nand U11859 (N_11859,N_9709,N_9040);
xor U11860 (N_11860,N_10099,N_9906);
nor U11861 (N_11861,N_10002,N_9717);
or U11862 (N_11862,N_9273,N_10494);
nand U11863 (N_11863,N_9648,N_9078);
or U11864 (N_11864,N_10000,N_9944);
and U11865 (N_11865,N_10283,N_10441);
nor U11866 (N_11866,N_9431,N_10044);
nor U11867 (N_11867,N_10200,N_9856);
nor U11868 (N_11868,N_9790,N_9154);
or U11869 (N_11869,N_9491,N_9955);
and U11870 (N_11870,N_9874,N_9506);
nand U11871 (N_11871,N_10245,N_9975);
or U11872 (N_11872,N_9764,N_10151);
nor U11873 (N_11873,N_10330,N_9954);
nand U11874 (N_11874,N_9055,N_9016);
or U11875 (N_11875,N_9001,N_9678);
and U11876 (N_11876,N_10429,N_10394);
and U11877 (N_11877,N_9670,N_9850);
nor U11878 (N_11878,N_9282,N_9310);
or U11879 (N_11879,N_10231,N_9677);
and U11880 (N_11880,N_9203,N_10313);
or U11881 (N_11881,N_9307,N_10467);
nand U11882 (N_11882,N_9789,N_9733);
xnor U11883 (N_11883,N_10044,N_9235);
nand U11884 (N_11884,N_9342,N_9826);
or U11885 (N_11885,N_10360,N_9369);
nor U11886 (N_11886,N_9264,N_9481);
xor U11887 (N_11887,N_10085,N_9962);
xor U11888 (N_11888,N_10337,N_10122);
nand U11889 (N_11889,N_9023,N_9695);
nor U11890 (N_11890,N_9184,N_9571);
nor U11891 (N_11891,N_9689,N_9169);
and U11892 (N_11892,N_10288,N_10419);
and U11893 (N_11893,N_9487,N_9531);
and U11894 (N_11894,N_9405,N_10343);
nor U11895 (N_11895,N_9146,N_9442);
xor U11896 (N_11896,N_10351,N_9520);
and U11897 (N_11897,N_9034,N_9596);
xor U11898 (N_11898,N_9517,N_10066);
and U11899 (N_11899,N_9318,N_9256);
xnor U11900 (N_11900,N_9003,N_9555);
xor U11901 (N_11901,N_9664,N_9631);
nand U11902 (N_11902,N_9382,N_10307);
nor U11903 (N_11903,N_10139,N_9398);
xnor U11904 (N_11904,N_10360,N_10071);
xor U11905 (N_11905,N_9325,N_9810);
or U11906 (N_11906,N_9287,N_10182);
nor U11907 (N_11907,N_10395,N_10237);
or U11908 (N_11908,N_9570,N_9762);
and U11909 (N_11909,N_9803,N_9614);
and U11910 (N_11910,N_10064,N_9527);
or U11911 (N_11911,N_9803,N_9993);
or U11912 (N_11912,N_9704,N_9745);
xor U11913 (N_11913,N_9289,N_9442);
nand U11914 (N_11914,N_9129,N_9874);
nor U11915 (N_11915,N_10307,N_9078);
xnor U11916 (N_11916,N_10260,N_9960);
and U11917 (N_11917,N_9540,N_10322);
nand U11918 (N_11918,N_10315,N_10277);
or U11919 (N_11919,N_9679,N_9475);
or U11920 (N_11920,N_9148,N_9813);
nand U11921 (N_11921,N_9146,N_10328);
nor U11922 (N_11922,N_9416,N_10195);
nor U11923 (N_11923,N_10364,N_9828);
or U11924 (N_11924,N_10241,N_9462);
nand U11925 (N_11925,N_10233,N_10017);
nor U11926 (N_11926,N_10199,N_9988);
nand U11927 (N_11927,N_9306,N_9004);
nand U11928 (N_11928,N_10160,N_9986);
nand U11929 (N_11929,N_10306,N_10170);
nand U11930 (N_11930,N_10130,N_9772);
and U11931 (N_11931,N_10403,N_9378);
nand U11932 (N_11932,N_10437,N_9678);
xor U11933 (N_11933,N_9823,N_10131);
or U11934 (N_11934,N_9485,N_9525);
or U11935 (N_11935,N_9900,N_9098);
or U11936 (N_11936,N_9772,N_9907);
nand U11937 (N_11937,N_10407,N_9112);
or U11938 (N_11938,N_9704,N_9997);
nor U11939 (N_11939,N_9817,N_10290);
xor U11940 (N_11940,N_10233,N_10212);
and U11941 (N_11941,N_9198,N_10182);
nand U11942 (N_11942,N_9054,N_10082);
nor U11943 (N_11943,N_9888,N_9653);
or U11944 (N_11944,N_10402,N_9309);
and U11945 (N_11945,N_9520,N_9535);
xnor U11946 (N_11946,N_10155,N_10283);
xnor U11947 (N_11947,N_9597,N_9421);
or U11948 (N_11948,N_9101,N_10462);
nor U11949 (N_11949,N_9711,N_9753);
xor U11950 (N_11950,N_9707,N_9336);
and U11951 (N_11951,N_9910,N_9331);
nand U11952 (N_11952,N_9353,N_9237);
and U11953 (N_11953,N_9209,N_10470);
xnor U11954 (N_11954,N_10259,N_9164);
and U11955 (N_11955,N_10071,N_10287);
xor U11956 (N_11956,N_9818,N_10389);
or U11957 (N_11957,N_10355,N_9936);
nor U11958 (N_11958,N_9879,N_10236);
or U11959 (N_11959,N_10475,N_10387);
and U11960 (N_11960,N_9810,N_10440);
xor U11961 (N_11961,N_9013,N_10153);
and U11962 (N_11962,N_9492,N_9925);
and U11963 (N_11963,N_9138,N_10050);
nor U11964 (N_11964,N_9139,N_9272);
nor U11965 (N_11965,N_9480,N_9515);
nand U11966 (N_11966,N_10167,N_9857);
xor U11967 (N_11967,N_10037,N_9988);
nand U11968 (N_11968,N_9563,N_9323);
xor U11969 (N_11969,N_9917,N_9289);
nand U11970 (N_11970,N_9630,N_9883);
and U11971 (N_11971,N_10226,N_9065);
xor U11972 (N_11972,N_10192,N_10168);
and U11973 (N_11973,N_10203,N_9413);
and U11974 (N_11974,N_9545,N_9699);
and U11975 (N_11975,N_9037,N_9401);
and U11976 (N_11976,N_10150,N_10427);
or U11977 (N_11977,N_9235,N_10096);
nand U11978 (N_11978,N_10475,N_9425);
nor U11979 (N_11979,N_9974,N_9264);
and U11980 (N_11980,N_10252,N_9157);
xnor U11981 (N_11981,N_10447,N_9233);
nor U11982 (N_11982,N_9405,N_9323);
or U11983 (N_11983,N_9934,N_9473);
and U11984 (N_11984,N_9093,N_9224);
or U11985 (N_11985,N_9835,N_10349);
and U11986 (N_11986,N_9614,N_10187);
and U11987 (N_11987,N_9938,N_9450);
xnor U11988 (N_11988,N_10123,N_9773);
or U11989 (N_11989,N_10010,N_9906);
nand U11990 (N_11990,N_9285,N_10290);
nand U11991 (N_11991,N_9992,N_9144);
and U11992 (N_11992,N_9601,N_9353);
nor U11993 (N_11993,N_9006,N_9499);
nor U11994 (N_11994,N_10083,N_9682);
xor U11995 (N_11995,N_9270,N_9645);
and U11996 (N_11996,N_9431,N_9368);
nand U11997 (N_11997,N_10404,N_9569);
nand U11998 (N_11998,N_10483,N_9078);
or U11999 (N_11999,N_9591,N_9306);
nor U12000 (N_12000,N_10961,N_11714);
or U12001 (N_12001,N_11241,N_11441);
xnor U12002 (N_12002,N_11504,N_10861);
and U12003 (N_12003,N_11567,N_10851);
nand U12004 (N_12004,N_11332,N_10729);
xor U12005 (N_12005,N_11793,N_11067);
or U12006 (N_12006,N_11640,N_11113);
nand U12007 (N_12007,N_10658,N_11650);
xor U12008 (N_12008,N_11514,N_11179);
nor U12009 (N_12009,N_11999,N_11828);
or U12010 (N_12010,N_11340,N_10684);
nand U12011 (N_12011,N_10556,N_11289);
nor U12012 (N_12012,N_11226,N_11552);
nand U12013 (N_12013,N_11304,N_11287);
nand U12014 (N_12014,N_10832,N_11173);
nand U12015 (N_12015,N_11358,N_10847);
or U12016 (N_12016,N_10512,N_11328);
xnor U12017 (N_12017,N_11543,N_11291);
or U12018 (N_12018,N_10764,N_11591);
nand U12019 (N_12019,N_11360,N_11326);
nor U12020 (N_12020,N_10824,N_10790);
or U12021 (N_12021,N_11570,N_10965);
xnor U12022 (N_12022,N_10649,N_10676);
xor U12023 (N_12023,N_11166,N_11622);
and U12024 (N_12024,N_10741,N_11833);
nor U12025 (N_12025,N_11485,N_11100);
nor U12026 (N_12026,N_11996,N_10924);
nand U12027 (N_12027,N_11525,N_11672);
and U12028 (N_12028,N_11503,N_11598);
or U12029 (N_12029,N_11080,N_11991);
xnor U12030 (N_12030,N_11721,N_11435);
nor U12031 (N_12031,N_11314,N_11666);
or U12032 (N_12032,N_10756,N_11933);
nor U12033 (N_12033,N_10980,N_11269);
nor U12034 (N_12034,N_10501,N_11183);
and U12035 (N_12035,N_10542,N_10648);
and U12036 (N_12036,N_11406,N_10683);
or U12037 (N_12037,N_11741,N_11042);
or U12038 (N_12038,N_11097,N_11807);
xor U12039 (N_12039,N_11271,N_11362);
nand U12040 (N_12040,N_10738,N_10918);
xnor U12041 (N_12041,N_10629,N_11123);
and U12042 (N_12042,N_11024,N_11238);
xor U12043 (N_12043,N_10695,N_11161);
xnor U12044 (N_12044,N_10560,N_11397);
nor U12045 (N_12045,N_11506,N_10569);
nand U12046 (N_12046,N_10717,N_11253);
nand U12047 (N_12047,N_11225,N_11861);
and U12048 (N_12048,N_11391,N_11477);
nand U12049 (N_12049,N_11605,N_11261);
nor U12050 (N_12050,N_11856,N_11973);
or U12051 (N_12051,N_11330,N_11323);
nand U12052 (N_12052,N_11408,N_10731);
and U12053 (N_12053,N_11122,N_11223);
xor U12054 (N_12054,N_11842,N_11559);
xnor U12055 (N_12055,N_11965,N_11583);
xor U12056 (N_12056,N_11727,N_10757);
or U12057 (N_12057,N_11799,N_11202);
and U12058 (N_12058,N_10660,N_11715);
and U12059 (N_12059,N_11544,N_11027);
or U12060 (N_12060,N_11617,N_10645);
or U12061 (N_12061,N_10674,N_11722);
nand U12062 (N_12062,N_11438,N_11930);
or U12063 (N_12063,N_11609,N_11811);
and U12064 (N_12064,N_11245,N_10713);
nand U12065 (N_12065,N_10547,N_10807);
or U12066 (N_12066,N_11150,N_11974);
xnor U12067 (N_12067,N_11732,N_11781);
xnor U12068 (N_12068,N_10769,N_10815);
and U12069 (N_12069,N_11127,N_11275);
nand U12070 (N_12070,N_10604,N_11257);
xnor U12071 (N_12071,N_10899,N_10936);
and U12072 (N_12072,N_10510,N_10829);
xor U12073 (N_12073,N_11213,N_11849);
nand U12074 (N_12074,N_10709,N_11294);
or U12075 (N_12075,N_11001,N_10794);
nand U12076 (N_12076,N_11553,N_10849);
nor U12077 (N_12077,N_11451,N_11639);
and U12078 (N_12078,N_11034,N_11797);
nor U12079 (N_12079,N_11248,N_11465);
xnor U12080 (N_12080,N_11051,N_10827);
or U12081 (N_12081,N_11554,N_11449);
nor U12082 (N_12082,N_11073,N_10916);
nand U12083 (N_12083,N_11897,N_10758);
xnor U12084 (N_12084,N_10608,N_11731);
xnor U12085 (N_12085,N_11911,N_11835);
and U12086 (N_12086,N_11433,N_11091);
or U12087 (N_12087,N_11535,N_10932);
nand U12088 (N_12088,N_11702,N_11082);
or U12089 (N_12089,N_11129,N_11874);
or U12090 (N_12090,N_10876,N_11987);
nand U12091 (N_12091,N_10969,N_10549);
or U12092 (N_12092,N_11376,N_11062);
and U12093 (N_12093,N_11203,N_11879);
nor U12094 (N_12094,N_10766,N_10503);
nor U12095 (N_12095,N_11063,N_10831);
nand U12096 (N_12096,N_10740,N_10810);
and U12097 (N_12097,N_11832,N_11555);
nor U12098 (N_12098,N_11379,N_11690);
nand U12099 (N_12099,N_10908,N_10571);
and U12100 (N_12100,N_11252,N_11300);
nor U12101 (N_12101,N_11475,N_11547);
nand U12102 (N_12102,N_11802,N_10811);
xor U12103 (N_12103,N_11986,N_11568);
xor U12104 (N_12104,N_10785,N_10643);
nor U12105 (N_12105,N_11762,N_11366);
and U12106 (N_12106,N_10545,N_11194);
and U12107 (N_12107,N_11794,N_11000);
or U12108 (N_12108,N_11751,N_11657);
nor U12109 (N_12109,N_11590,N_10987);
nand U12110 (N_12110,N_11560,N_10947);
xor U12111 (N_12111,N_10825,N_11284);
nor U12112 (N_12112,N_10808,N_11906);
xor U12113 (N_12113,N_10647,N_11395);
nor U12114 (N_12114,N_10983,N_11199);
and U12115 (N_12115,N_10664,N_11997);
and U12116 (N_12116,N_10621,N_10591);
and U12117 (N_12117,N_11821,N_11789);
and U12118 (N_12118,N_10711,N_11884);
nand U12119 (N_12119,N_10948,N_10665);
or U12120 (N_12120,N_11264,N_10972);
or U12121 (N_12121,N_11921,N_11882);
nand U12122 (N_12122,N_10784,N_11681);
xnor U12123 (N_12123,N_10506,N_10630);
xor U12124 (N_12124,N_11613,N_10990);
nor U12125 (N_12125,N_11317,N_10742);
nor U12126 (N_12126,N_11759,N_10791);
xor U12127 (N_12127,N_10973,N_11780);
nand U12128 (N_12128,N_11411,N_10715);
nand U12129 (N_12129,N_11356,N_10786);
or U12130 (N_12130,N_10511,N_11324);
nor U12131 (N_12131,N_10737,N_11233);
nor U12132 (N_12132,N_10687,N_10735);
nand U12133 (N_12133,N_11370,N_10920);
or U12134 (N_12134,N_11197,N_10537);
nor U12135 (N_12135,N_10736,N_11392);
nor U12136 (N_12136,N_11019,N_11888);
or U12137 (N_12137,N_10652,N_10610);
nor U12138 (N_12138,N_11185,N_11153);
or U12139 (N_12139,N_10619,N_11131);
or U12140 (N_12140,N_11703,N_11581);
xor U12141 (N_12141,N_11147,N_11154);
nor U12142 (N_12142,N_10733,N_11803);
nor U12143 (N_12143,N_10612,N_11499);
or U12144 (N_12144,N_11577,N_11306);
and U12145 (N_12145,N_10580,N_10699);
nor U12146 (N_12146,N_11212,N_11028);
nand U12147 (N_12147,N_11162,N_11716);
and U12148 (N_12148,N_11148,N_10890);
xnor U12149 (N_12149,N_11094,N_11787);
or U12150 (N_12150,N_11293,N_11976);
nor U12151 (N_12151,N_11769,N_11557);
or U12152 (N_12152,N_11218,N_11662);
or U12153 (N_12153,N_11563,N_11130);
xnor U12154 (N_12154,N_10934,N_11854);
xor U12155 (N_12155,N_11195,N_10703);
xor U12156 (N_12156,N_11184,N_11462);
and U12157 (N_12157,N_11669,N_11817);
nor U12158 (N_12158,N_11335,N_10767);
xor U12159 (N_12159,N_11527,N_10595);
and U12160 (N_12160,N_11457,N_10869);
nor U12161 (N_12161,N_10917,N_11984);
nor U12162 (N_12162,N_11423,N_10989);
or U12163 (N_12163,N_10639,N_11536);
nand U12164 (N_12164,N_11501,N_11198);
nand U12165 (N_12165,N_11818,N_10531);
and U12166 (N_12166,N_11945,N_10780);
or U12167 (N_12167,N_11822,N_10698);
or U12168 (N_12168,N_11894,N_11924);
or U12169 (N_12169,N_10602,N_11163);
or U12170 (N_12170,N_11117,N_11415);
nand U12171 (N_12171,N_11603,N_10586);
nand U12172 (N_12172,N_11421,N_10966);
xor U12173 (N_12173,N_11417,N_10759);
nand U12174 (N_12174,N_10776,N_11045);
nor U12175 (N_12175,N_11813,N_11493);
or U12176 (N_12176,N_10789,N_10615);
nor U12177 (N_12177,N_11419,N_10685);
and U12178 (N_12178,N_11352,N_11982);
and U12179 (N_12179,N_11315,N_11954);
nand U12180 (N_12180,N_11827,N_11929);
or U12181 (N_12181,N_11160,N_10730);
xor U12182 (N_12182,N_10535,N_11685);
nand U12183 (N_12183,N_11054,N_11021);
or U12184 (N_12184,N_10605,N_10992);
and U12185 (N_12185,N_11420,N_11846);
and U12186 (N_12186,N_10541,N_10804);
xnor U12187 (N_12187,N_11491,N_11508);
or U12188 (N_12188,N_11180,N_11737);
or U12189 (N_12189,N_10568,N_10835);
nand U12190 (N_12190,N_11642,N_11146);
and U12191 (N_12191,N_11579,N_11636);
xor U12192 (N_12192,N_10878,N_11013);
nor U12193 (N_12193,N_11592,N_10889);
nor U12194 (N_12194,N_11061,N_10977);
nand U12195 (N_12195,N_10912,N_11215);
xor U12196 (N_12196,N_11249,N_11318);
xnor U12197 (N_12197,N_11187,N_11096);
nor U12198 (N_12198,N_11600,N_11172);
nand U12199 (N_12199,N_11711,N_11643);
nor U12200 (N_12200,N_11389,N_11628);
or U12201 (N_12201,N_10819,N_11677);
or U12202 (N_12202,N_11492,N_11740);
or U12203 (N_12203,N_11339,N_11145);
and U12204 (N_12204,N_11255,N_10734);
nor U12205 (N_12205,N_11890,N_11608);
nor U12206 (N_12206,N_11667,N_11035);
and U12207 (N_12207,N_10840,N_11396);
nor U12208 (N_12208,N_11734,N_11490);
xnor U12209 (N_12209,N_11513,N_11437);
nand U12210 (N_12210,N_10588,N_10644);
or U12211 (N_12211,N_10671,N_10892);
or U12212 (N_12212,N_11967,N_10529);
nand U12213 (N_12213,N_11717,N_10507);
nor U12214 (N_12214,N_11192,N_10944);
xor U12215 (N_12215,N_11009,N_11791);
and U12216 (N_12216,N_11134,N_11847);
xnor U12217 (N_12217,N_11784,N_11645);
nor U12218 (N_12218,N_11586,N_10986);
xnor U12219 (N_12219,N_11774,N_11786);
nor U12220 (N_12220,N_11938,N_11268);
nand U12221 (N_12221,N_11654,N_11334);
nand U12222 (N_12222,N_10561,N_10651);
nor U12223 (N_12223,N_11521,N_11103);
and U12224 (N_12224,N_11319,N_11047);
and U12225 (N_12225,N_11414,N_11723);
or U12226 (N_12226,N_10637,N_11355);
and U12227 (N_12227,N_11534,N_11664);
nand U12228 (N_12228,N_11707,N_10628);
and U12229 (N_12229,N_11469,N_11305);
xor U12230 (N_12230,N_11008,N_11140);
or U12231 (N_12231,N_10566,N_10500);
or U12232 (N_12232,N_11452,N_11016);
and U12233 (N_12233,N_11267,N_10668);
nand U12234 (N_12234,N_11671,N_10617);
xor U12235 (N_12235,N_11222,N_10792);
and U12236 (N_12236,N_11804,N_11281);
nor U12237 (N_12237,N_11038,N_11824);
or U12238 (N_12238,N_11597,N_10865);
xor U12239 (N_12239,N_11750,N_10576);
nand U12240 (N_12240,N_11602,N_10999);
xnor U12241 (N_12241,N_10783,N_11151);
and U12242 (N_12242,N_11770,N_10739);
nor U12243 (N_12243,N_10853,N_11312);
xor U12244 (N_12244,N_11668,N_10875);
nand U12245 (N_12245,N_10521,N_11816);
or U12246 (N_12246,N_11859,N_11529);
and U12247 (N_12247,N_11193,N_10593);
nor U12248 (N_12248,N_10870,N_10841);
nand U12249 (N_12249,N_11810,N_11981);
or U12250 (N_12250,N_11754,N_11234);
nand U12251 (N_12251,N_10866,N_11059);
and U12252 (N_12252,N_10817,N_10814);
nor U12253 (N_12253,N_11076,N_11994);
xnor U12254 (N_12254,N_11413,N_11487);
or U12255 (N_12255,N_11159,N_11857);
or U12256 (N_12256,N_11775,N_10777);
xnor U12257 (N_12257,N_11927,N_10993);
nor U12258 (N_12258,N_11152,N_11439);
nor U12259 (N_12259,N_10770,N_10657);
or U12260 (N_12260,N_11044,N_11616);
nor U12261 (N_12261,N_11676,N_11273);
and U12262 (N_12262,N_11032,N_11277);
and U12263 (N_12263,N_11484,N_11985);
or U12264 (N_12264,N_11382,N_11948);
xor U12265 (N_12265,N_11752,N_11706);
or U12266 (N_12266,N_11693,N_11354);
and U12267 (N_12267,N_10527,N_10834);
or U12268 (N_12268,N_11200,N_11060);
and U12269 (N_12269,N_11545,N_11720);
or U12270 (N_12270,N_11839,N_10796);
nor U12271 (N_12271,N_11470,N_10826);
nand U12272 (N_12272,N_11805,N_11673);
xor U12273 (N_12273,N_10991,N_10806);
and U12274 (N_12274,N_10663,N_10910);
nand U12275 (N_12275,N_10744,N_10844);
or U12276 (N_12276,N_10539,N_11964);
xor U12277 (N_12277,N_11764,N_11992);
or U12278 (N_12278,N_11922,N_11814);
nor U12279 (N_12279,N_11282,N_10900);
xnor U12280 (N_12280,N_10523,N_10942);
xnor U12281 (N_12281,N_11309,N_11782);
and U12282 (N_12282,N_11511,N_10816);
nand U12283 (N_12283,N_11655,N_10570);
and U12284 (N_12284,N_11588,N_11518);
and U12285 (N_12285,N_11486,N_11206);
and U12286 (N_12286,N_11081,N_11409);
nand U12287 (N_12287,N_10528,N_10719);
nand U12288 (N_12288,N_11878,N_11558);
nand U12289 (N_12289,N_10655,N_11456);
xnor U12290 (N_12290,N_10636,N_11364);
and U12291 (N_12291,N_10863,N_11077);
and U12292 (N_12292,N_11398,N_10672);
nor U12293 (N_12293,N_10797,N_11246);
or U12294 (N_12294,N_11260,N_10682);
xnor U12295 (N_12295,N_10925,N_11855);
nand U12296 (N_12296,N_11120,N_10710);
or U12297 (N_12297,N_10781,N_10631);
xnor U12298 (N_12298,N_11983,N_11251);
or U12299 (N_12299,N_10613,N_11573);
or U12300 (N_12300,N_11660,N_10728);
xor U12301 (N_12301,N_10653,N_10941);
or U12302 (N_12302,N_11320,N_10592);
or U12303 (N_12303,N_10801,N_11851);
and U12304 (N_12304,N_11495,N_11729);
or U12305 (N_12305,N_11649,N_11777);
nor U12306 (N_12306,N_11126,N_11385);
and U12307 (N_12307,N_11958,N_11712);
or U12308 (N_12308,N_11182,N_11164);
xor U12309 (N_12309,N_11479,N_11407);
or U12310 (N_12310,N_11471,N_11381);
nand U12311 (N_12311,N_11007,N_11889);
or U12312 (N_12312,N_11885,N_11211);
and U12313 (N_12313,N_10525,N_11682);
xnor U12314 (N_12314,N_10859,N_11228);
nor U12315 (N_12315,N_11826,N_10765);
and U12316 (N_12316,N_11448,N_10774);
xnor U12317 (N_12317,N_10706,N_10955);
or U12318 (N_12318,N_11003,N_11057);
and U12319 (N_12319,N_10998,N_11405);
or U12320 (N_12320,N_11429,N_11629);
nor U12321 (N_12321,N_11383,N_10577);
nand U12322 (N_12322,N_11533,N_11109);
or U12323 (N_12323,N_10707,N_11960);
nand U12324 (N_12324,N_10952,N_11766);
xnor U12325 (N_12325,N_11372,N_10574);
and U12326 (N_12326,N_10673,N_11072);
xor U12327 (N_12327,N_11041,N_11204);
and U12328 (N_12328,N_11216,N_11863);
nor U12329 (N_12329,N_11537,N_10708);
or U12330 (N_12330,N_11648,N_10558);
xor U12331 (N_12331,N_11135,N_11280);
nand U12332 (N_12332,N_11401,N_11142);
or U12333 (N_12333,N_11895,N_11626);
nor U12334 (N_12334,N_11101,N_10837);
nor U12335 (N_12335,N_11733,N_11037);
xor U12336 (N_12336,N_11388,N_11546);
nor U12337 (N_12337,N_11928,N_11311);
xnor U12338 (N_12338,N_11399,N_11393);
and U12339 (N_12339,N_11351,N_10646);
and U12340 (N_12340,N_11040,N_11048);
and U12341 (N_12341,N_11473,N_10830);
and U12342 (N_12342,N_10599,N_10959);
xnor U12343 (N_12343,N_11286,N_11739);
and U12344 (N_12344,N_10988,N_11102);
xor U12345 (N_12345,N_11829,N_11387);
or U12346 (N_12346,N_10662,N_10919);
xor U12347 (N_12347,N_11887,N_10681);
or U12348 (N_12348,N_10701,N_10897);
nand U12349 (N_12349,N_10596,N_11674);
nand U12350 (N_12350,N_11988,N_10896);
xnor U12351 (N_12351,N_11725,N_11176);
and U12352 (N_12352,N_11136,N_10903);
xor U12353 (N_12353,N_11873,N_10754);
or U12354 (N_12354,N_11463,N_11404);
nand U12355 (N_12355,N_10552,N_11256);
xnor U12356 (N_12356,N_11549,N_11104);
nand U12357 (N_12357,N_11410,N_11593);
nand U12358 (N_12358,N_11756,N_11601);
nand U12359 (N_12359,N_11380,N_11867);
and U12360 (N_12360,N_10614,N_11502);
and U12361 (N_12361,N_11095,N_11902);
or U12362 (N_12362,N_10799,N_11550);
and U12363 (N_12363,N_11892,N_10555);
xnor U12364 (N_12364,N_10563,N_11893);
nand U12365 (N_12365,N_11941,N_10534);
and U12366 (N_12366,N_10930,N_11338);
nand U12367 (N_12367,N_10543,N_11052);
or U12368 (N_12368,N_10666,N_10659);
nand U12369 (N_12369,N_11205,N_11699);
and U12370 (N_12370,N_10937,N_11374);
nor U12371 (N_12371,N_10583,N_10909);
and U12372 (N_12372,N_11220,N_11089);
and U12373 (N_12373,N_11790,N_11905);
and U12374 (N_12374,N_11870,N_11971);
and U12375 (N_12375,N_10975,N_11798);
and U12376 (N_12376,N_11002,N_11708);
xor U12377 (N_12377,N_11209,N_10712);
nand U12378 (N_12378,N_11262,N_11812);
or U12379 (N_12379,N_11815,N_11963);
and U12380 (N_12380,N_10690,N_10782);
and U12381 (N_12381,N_11178,N_11792);
and U12382 (N_12382,N_11128,N_11494);
and U12383 (N_12383,N_10584,N_10836);
nand U12384 (N_12384,N_11313,N_10705);
xor U12385 (N_12385,N_11801,N_11075);
nor U12386 (N_12386,N_10787,N_11214);
and U12387 (N_12387,N_11916,N_10763);
nand U12388 (N_12388,N_11820,N_10618);
and U12389 (N_12389,N_10939,N_11303);
nand U12390 (N_12390,N_10761,N_10626);
xor U12391 (N_12391,N_11087,N_11105);
and U12392 (N_12392,N_10795,N_11086);
nor U12393 (N_12393,N_11619,N_11990);
nor U12394 (N_12394,N_11359,N_10633);
xnor U12395 (N_12395,N_11844,N_11575);
nand U12396 (N_12396,N_10773,N_11295);
or U12397 (N_12397,N_11476,N_11302);
nor U12398 (N_12398,N_11431,N_11637);
xnor U12399 (N_12399,N_11346,N_11270);
nand U12400 (N_12400,N_11541,N_11663);
nor U12401 (N_12401,N_10743,N_10727);
nor U12402 (N_12402,N_11531,N_10839);
nor U12403 (N_12403,N_10679,N_10518);
and U12404 (N_12404,N_10911,N_11478);
or U12405 (N_12405,N_10883,N_10760);
nor U12406 (N_12406,N_11450,N_10958);
nor U12407 (N_12407,N_10881,N_10905);
or U12408 (N_12408,N_11866,N_11083);
and U12409 (N_12409,N_11630,N_11447);
nor U12410 (N_12410,N_11788,N_11736);
nor U12411 (N_12411,N_11749,N_11403);
or U12412 (N_12412,N_10603,N_11612);
xnor U12413 (N_12413,N_11207,N_10597);
and U12414 (N_12414,N_10778,N_10746);
and U12415 (N_12415,N_11691,N_11012);
nand U12416 (N_12416,N_11850,N_11975);
nor U12417 (N_12417,N_11719,N_10625);
or U12418 (N_12418,N_11589,N_11175);
or U12419 (N_12419,N_10575,N_11090);
nor U12420 (N_12420,N_10802,N_11779);
nand U12421 (N_12421,N_11036,N_10893);
nand U12422 (N_12422,N_11112,N_10940);
nor U12423 (N_12423,N_11098,N_11778);
or U12424 (N_12424,N_11572,N_11858);
xor U12425 (N_12425,N_10590,N_11496);
nor U12426 (N_12426,N_10964,N_11853);
nand U12427 (N_12427,N_11623,N_10894);
nand U12428 (N_12428,N_11308,N_11116);
nor U12429 (N_12429,N_11763,N_11580);
nand U12430 (N_12430,N_10587,N_11307);
nand U12431 (N_12431,N_11901,N_11701);
or U12432 (N_12432,N_11349,N_10627);
xnor U12433 (N_12433,N_10954,N_11758);
xor U12434 (N_12434,N_10858,N_11053);
nor U12435 (N_12435,N_10589,N_11684);
nand U12436 (N_12436,N_10609,N_11442);
xor U12437 (N_12437,N_11773,N_11488);
xnor U12438 (N_12438,N_11898,N_10996);
or U12439 (N_12439,N_11344,N_11108);
xnor U12440 (N_12440,N_10871,N_11208);
nor U12441 (N_12441,N_11137,N_11015);
and U12442 (N_12442,N_11783,N_11830);
and U12443 (N_12443,N_11279,N_11697);
or U12444 (N_12444,N_10642,N_10530);
nand U12445 (N_12445,N_11947,N_11900);
nand U12446 (N_12446,N_11050,N_11757);
nor U12447 (N_12447,N_11606,N_11432);
and U12448 (N_12448,N_11139,N_10564);
nor U12449 (N_12449,N_11196,N_10768);
nor U12450 (N_12450,N_10689,N_11026);
xor U12451 (N_12451,N_11883,N_10753);
nor U12452 (N_12452,N_11329,N_11565);
and U12453 (N_12453,N_11014,N_10884);
nor U12454 (N_12454,N_11551,N_11970);
nor U12455 (N_12455,N_11955,N_11968);
nand U12456 (N_12456,N_10536,N_11995);
or U12457 (N_12457,N_11571,N_10585);
xor U12458 (N_12458,N_11064,N_11678);
nand U12459 (N_12459,N_10526,N_11240);
xor U12460 (N_12460,N_10579,N_11872);
or U12461 (N_12461,N_11653,N_11819);
or U12462 (N_12462,N_11809,N_10598);
or U12463 (N_12463,N_10967,N_11876);
nor U12464 (N_12464,N_11687,N_11942);
and U12465 (N_12465,N_10809,N_11296);
nand U12466 (N_12466,N_11989,N_11446);
nand U12467 (N_12467,N_11652,N_10723);
nand U12468 (N_12468,N_11031,N_11538);
nor U12469 (N_12469,N_10661,N_11528);
and U12470 (N_12470,N_11634,N_11977);
and U12471 (N_12471,N_10522,N_10828);
nor U12472 (N_12472,N_10845,N_11005);
nor U12473 (N_12473,N_11564,N_10704);
nor U12474 (N_12474,N_10800,N_11615);
nand U12475 (N_12475,N_11510,N_11950);
or U12476 (N_12476,N_11509,N_11400);
nand U12477 (N_12477,N_11497,N_10904);
and U12478 (N_12478,N_10922,N_10788);
nand U12479 (N_12479,N_11341,N_10885);
or U12480 (N_12480,N_11464,N_11453);
nand U12481 (N_12481,N_11848,N_11939);
nor U12482 (N_12482,N_11219,N_11919);
or U12483 (N_12483,N_11926,N_11321);
nand U12484 (N_12484,N_11542,N_11066);
xnor U12485 (N_12485,N_10572,N_10732);
xor U12486 (N_12486,N_11595,N_10976);
and U12487 (N_12487,N_11765,N_11638);
nor U12488 (N_12488,N_11907,N_11357);
nand U12489 (N_12489,N_10578,N_10700);
or U12490 (N_12490,N_11651,N_10935);
nand U12491 (N_12491,N_10927,N_11865);
or U12492 (N_12492,N_11582,N_11795);
xor U12493 (N_12493,N_11959,N_11556);
nor U12494 (N_12494,N_10960,N_11068);
and U12495 (N_12495,N_11468,N_11576);
nor U12496 (N_12496,N_10519,N_11728);
and U12497 (N_12497,N_10718,N_11585);
xor U12498 (N_12498,N_10970,N_10546);
nor U12499 (N_12499,N_11378,N_11625);
nand U12500 (N_12500,N_10860,N_11523);
xnor U12501 (N_12501,N_10901,N_11755);
or U12502 (N_12502,N_10692,N_10879);
nand U12503 (N_12503,N_10623,N_11143);
nor U12504 (N_12504,N_11972,N_10680);
nand U12505 (N_12505,N_10945,N_11093);
nand U12506 (N_12506,N_11908,N_11459);
nor U12507 (N_12507,N_11416,N_10822);
nor U12508 (N_12508,N_11345,N_10915);
nand U12509 (N_12509,N_10544,N_11656);
nor U12510 (N_12510,N_11864,N_11923);
nor U12511 (N_12511,N_11394,N_10949);
and U12512 (N_12512,N_11023,N_10550);
nand U12513 (N_12513,N_11285,N_11886);
nor U12514 (N_12514,N_11946,N_11647);
or U12515 (N_12515,N_11422,N_10855);
xnor U12516 (N_12516,N_10926,N_11018);
or U12517 (N_12517,N_10974,N_10667);
nand U12518 (N_12518,N_10882,N_10540);
or U12519 (N_12519,N_11369,N_10750);
nand U12520 (N_12520,N_11030,N_10693);
and U12521 (N_12521,N_11325,N_10600);
xnor U12522 (N_12522,N_11298,N_10634);
nand U12523 (N_12523,N_11904,N_11505);
nor U12524 (N_12524,N_10548,N_11896);
or U12525 (N_12525,N_11517,N_11227);
or U12526 (N_12526,N_10533,N_11917);
and U12527 (N_12527,N_11744,N_11482);
nor U12528 (N_12528,N_11823,N_11115);
nor U12529 (N_12529,N_11365,N_11633);
and U12530 (N_12530,N_10638,N_10873);
xor U12531 (N_12531,N_11943,N_11074);
nor U12532 (N_12532,N_10696,N_10509);
xor U12533 (N_12533,N_11133,N_11596);
nor U12534 (N_12534,N_11111,N_10843);
or U12535 (N_12535,N_11418,N_11278);
or U12536 (N_12536,N_11940,N_10971);
and U12537 (N_12537,N_11231,N_10854);
nand U12538 (N_12538,N_10868,N_10624);
and U12539 (N_12539,N_11426,N_10721);
and U12540 (N_12540,N_11474,N_10898);
nand U12541 (N_12541,N_10514,N_11522);
nor U12542 (N_12542,N_10720,N_11055);
nand U12543 (N_12543,N_11679,N_11704);
nor U12544 (N_12544,N_11071,N_11838);
or U12545 (N_12545,N_11698,N_11428);
xor U12546 (N_12546,N_11840,N_10582);
nand U12547 (N_12547,N_11337,N_10813);
nand U12548 (N_12548,N_11114,N_11578);
xor U12549 (N_12549,N_10686,N_11610);
nand U12550 (N_12550,N_11283,N_10513);
and U12551 (N_12551,N_11425,N_11085);
xor U12552 (N_12552,N_10654,N_10891);
xor U12553 (N_12553,N_11444,N_11353);
and U12554 (N_12554,N_10607,N_11342);
xor U12555 (N_12555,N_11915,N_10650);
nand U12556 (N_12556,N_11607,N_11748);
xor U12557 (N_12557,N_10517,N_11745);
nor U12558 (N_12558,N_11520,N_10601);
xnor U12559 (N_12559,N_10848,N_11033);
or U12560 (N_12560,N_11532,N_11371);
nand U12561 (N_12561,N_11125,N_10622);
xnor U12562 (N_12562,N_11006,N_10775);
xnor U12563 (N_12563,N_10946,N_10508);
xnor U12564 (N_12564,N_11455,N_11149);
or U12565 (N_12565,N_11566,N_11709);
nor U12566 (N_12566,N_11029,N_11110);
xnor U12567 (N_12567,N_11368,N_10931);
nand U12568 (N_12568,N_11480,N_11156);
nor U12569 (N_12569,N_11301,N_10670);
or U12570 (N_12570,N_11644,N_10846);
nor U12571 (N_12571,N_11367,N_11079);
or U12572 (N_12572,N_11562,N_11979);
nand U12573 (N_12573,N_11025,N_10923);
xnor U12574 (N_12574,N_11157,N_11785);
or U12575 (N_12575,N_10504,N_11224);
nand U12576 (N_12576,N_11909,N_11386);
xnor U12577 (N_12577,N_11569,N_11288);
nor U12578 (N_12578,N_10793,N_11925);
or U12579 (N_12579,N_11343,N_11186);
and U12580 (N_12580,N_11507,N_10957);
or U12581 (N_12581,N_10635,N_10805);
or U12582 (N_12582,N_11746,N_11718);
nand U12583 (N_12583,N_11265,N_10951);
nand U12584 (N_12584,N_10921,N_11614);
nor U12585 (N_12585,N_10505,N_11363);
xnor U12586 (N_12586,N_11899,N_10559);
nor U12587 (N_12587,N_10515,N_10565);
and U12588 (N_12588,N_10872,N_10762);
and U12589 (N_12589,N_11618,N_11170);
or U12590 (N_12590,N_11953,N_11065);
or U12591 (N_12591,N_10842,N_11483);
nand U12592 (N_12592,N_11461,N_11771);
xnor U12593 (N_12593,N_11049,N_11747);
and U12594 (N_12594,N_10929,N_11611);
nand U12595 (N_12595,N_11242,N_10714);
nor U12596 (N_12596,N_10520,N_10640);
nor U12597 (N_12597,N_11526,N_11512);
xnor U12598 (N_12598,N_10864,N_10554);
xor U12599 (N_12599,N_11658,N_11272);
nand U12600 (N_12600,N_11675,N_10803);
nor U12601 (N_12601,N_11384,N_10724);
nor U12602 (N_12602,N_11831,N_10857);
and U12603 (N_12603,N_11862,N_11806);
and U12604 (N_12604,N_11519,N_11808);
and U12605 (N_12605,N_11046,N_11058);
and U12606 (N_12606,N_10551,N_10950);
or U12607 (N_12607,N_10524,N_11661);
xor U12608 (N_12608,N_11910,N_10877);
xor U12609 (N_12609,N_10616,N_11348);
or U12610 (N_12610,N_11167,N_11022);
xnor U12611 (N_12611,N_11978,N_11841);
and U12612 (N_12612,N_11688,N_11761);
nor U12613 (N_12613,N_11177,N_11056);
or U12614 (N_12614,N_11489,N_10962);
nor U12615 (N_12615,N_11735,N_10573);
xnor U12616 (N_12616,N_11800,N_11158);
xnor U12617 (N_12617,N_10725,N_11190);
or U12618 (N_12618,N_10694,N_11632);
nor U12619 (N_12619,N_10611,N_11891);
nand U12620 (N_12620,N_11957,N_11004);
nand U12621 (N_12621,N_11402,N_11084);
nor U12622 (N_12622,N_11825,N_10567);
or U12623 (N_12623,N_10553,N_11500);
nor U12624 (N_12624,N_11132,N_10953);
nand U12625 (N_12625,N_11138,N_10606);
xnor U12626 (N_12626,N_10833,N_11221);
xnor U12627 (N_12627,N_11229,N_11659);
xor U12628 (N_12628,N_11621,N_11375);
nor U12629 (N_12629,N_11118,N_11171);
or U12630 (N_12630,N_11333,N_10880);
or U12631 (N_12631,N_11373,N_11297);
nand U12632 (N_12632,N_11292,N_11443);
nor U12633 (N_12633,N_10938,N_11336);
or U12634 (N_12634,N_11738,N_11834);
nand U12635 (N_12635,N_10771,N_11768);
or U12636 (N_12636,N_10688,N_11913);
or U12637 (N_12637,N_11119,N_11980);
nand U12638 (N_12638,N_10928,N_11743);
nor U12639 (N_12639,N_11347,N_11646);
and U12640 (N_12640,N_11472,N_11524);
xnor U12641 (N_12641,N_10943,N_11189);
nand U12642 (N_12642,N_11694,N_11011);
nand U12643 (N_12643,N_11350,N_11169);
nand U12644 (N_12644,N_11689,N_11918);
or U12645 (N_12645,N_11424,N_10751);
nand U12646 (N_12646,N_11767,N_11776);
and U12647 (N_12647,N_11753,N_11695);
nand U12648 (N_12648,N_11266,N_10798);
and U12649 (N_12649,N_10984,N_11881);
nor U12650 (N_12650,N_11837,N_11935);
or U12651 (N_12651,N_10594,N_11730);
and U12652 (N_12652,N_10906,N_11467);
nand U12653 (N_12653,N_11237,N_11263);
nand U12654 (N_12654,N_11920,N_11445);
or U12655 (N_12655,N_11868,N_11966);
nor U12656 (N_12656,N_11686,N_11936);
nand U12657 (N_12657,N_10722,N_11670);
or U12658 (N_12658,N_11683,N_11217);
xnor U12659 (N_12659,N_11181,N_11174);
and U12660 (N_12660,N_11434,N_11481);
nand U12661 (N_12661,N_11680,N_11880);
nand U12662 (N_12662,N_11039,N_10538);
nor U12663 (N_12663,N_10850,N_11530);
nor U12664 (N_12664,N_11144,N_11498);
nand U12665 (N_12665,N_10581,N_11427);
xnor U12666 (N_12666,N_11258,N_11836);
or U12667 (N_12667,N_11106,N_11961);
or U12668 (N_12668,N_11010,N_10887);
and U12669 (N_12669,N_11860,N_11700);
and U12670 (N_12670,N_10779,N_11276);
and U12671 (N_12671,N_11993,N_10933);
nor U12672 (N_12672,N_11604,N_11931);
or U12673 (N_12673,N_11107,N_11436);
and U12674 (N_12674,N_11440,N_10982);
and U12675 (N_12675,N_11460,N_11875);
or U12676 (N_12676,N_10914,N_10888);
and U12677 (N_12677,N_10749,N_10820);
nor U12678 (N_12678,N_11952,N_11390);
and U12679 (N_12679,N_10632,N_11962);
nand U12680 (N_12680,N_11949,N_10978);
nor U12681 (N_12681,N_11239,N_11594);
or U12682 (N_12682,N_10818,N_11188);
nor U12683 (N_12683,N_10852,N_10677);
nor U12684 (N_12684,N_11201,N_11099);
xor U12685 (N_12685,N_10902,N_11796);
nand U12686 (N_12686,N_11092,N_11274);
xor U12687 (N_12687,N_11454,N_10516);
nand U12688 (N_12688,N_11070,N_10913);
and U12689 (N_12689,N_10669,N_10968);
nand U12690 (N_12690,N_10997,N_11635);
xnor U12691 (N_12691,N_11561,N_11259);
xnor U12692 (N_12692,N_11877,N_10747);
and U12693 (N_12693,N_10675,N_11713);
and U12694 (N_12694,N_11869,N_10697);
nand U12695 (N_12695,N_10981,N_10979);
xor U12696 (N_12696,N_10823,N_10726);
nor U12697 (N_12697,N_10752,N_11247);
or U12698 (N_12698,N_10656,N_11290);
nor U12699 (N_12699,N_11540,N_10502);
or U12700 (N_12700,N_11244,N_11852);
or U12701 (N_12701,N_11724,N_11599);
or U12702 (N_12702,N_10963,N_11944);
and U12703 (N_12703,N_11121,N_11871);
or U12704 (N_12704,N_11956,N_11914);
and U12705 (N_12705,N_11078,N_11710);
nor U12706 (N_12706,N_11548,N_11620);
and U12707 (N_12707,N_11412,N_11772);
nor U12708 (N_12708,N_10772,N_11141);
or U12709 (N_12709,N_11254,N_11539);
nor U12710 (N_12710,N_10562,N_11584);
nor U12711 (N_12711,N_10856,N_11250);
xor U12712 (N_12712,N_11998,N_11912);
nand U12713 (N_12713,N_10995,N_11327);
nand U12714 (N_12714,N_10956,N_10532);
xnor U12715 (N_12715,N_10886,N_11069);
nand U12716 (N_12716,N_11641,N_11430);
xnor U12717 (N_12717,N_11165,N_10907);
nand U12718 (N_12718,N_11232,N_10874);
nor U12719 (N_12719,N_11299,N_11665);
nor U12720 (N_12720,N_11361,N_10755);
and U12721 (N_12721,N_11191,N_10895);
xor U12722 (N_12722,N_11466,N_10745);
nor U12723 (N_12723,N_11627,N_11903);
or U12724 (N_12724,N_11377,N_11017);
or U12725 (N_12725,N_10812,N_11515);
and U12726 (N_12726,N_11124,N_10838);
nand U12727 (N_12727,N_11696,N_11937);
nor U12728 (N_12728,N_11587,N_11934);
nor U12729 (N_12729,N_10867,N_11236);
and U12730 (N_12730,N_11845,N_10557);
nand U12731 (N_12731,N_11631,N_11516);
xnor U12732 (N_12732,N_10985,N_11088);
xnor U12733 (N_12733,N_11969,N_10702);
and U12734 (N_12734,N_11210,N_11316);
nor U12735 (N_12735,N_11458,N_10994);
xnor U12736 (N_12736,N_10716,N_11705);
nor U12737 (N_12737,N_11043,N_11168);
and U12738 (N_12738,N_10862,N_11760);
nand U12739 (N_12739,N_11155,N_11951);
nor U12740 (N_12740,N_11230,N_10678);
nor U12741 (N_12741,N_10821,N_11843);
and U12742 (N_12742,N_11692,N_11310);
or U12743 (N_12743,N_11726,N_10620);
nand U12744 (N_12744,N_11932,N_10748);
or U12745 (N_12745,N_11322,N_11235);
nand U12746 (N_12746,N_11742,N_11624);
and U12747 (N_12747,N_11331,N_11020);
and U12748 (N_12748,N_10691,N_11574);
xnor U12749 (N_12749,N_10641,N_11243);
xnor U12750 (N_12750,N_10858,N_11318);
or U12751 (N_12751,N_10892,N_11798);
or U12752 (N_12752,N_11403,N_11652);
and U12753 (N_12753,N_11124,N_11033);
nor U12754 (N_12754,N_10993,N_11021);
or U12755 (N_12755,N_10782,N_11730);
or U12756 (N_12756,N_10990,N_11428);
nor U12757 (N_12757,N_11258,N_11541);
or U12758 (N_12758,N_11945,N_10507);
and U12759 (N_12759,N_10973,N_10622);
xnor U12760 (N_12760,N_11006,N_11047);
xnor U12761 (N_12761,N_11437,N_10731);
nor U12762 (N_12762,N_11938,N_11189);
or U12763 (N_12763,N_10928,N_10804);
xnor U12764 (N_12764,N_11346,N_11617);
or U12765 (N_12765,N_10943,N_10926);
nor U12766 (N_12766,N_11596,N_11643);
and U12767 (N_12767,N_11438,N_11441);
or U12768 (N_12768,N_11811,N_11153);
nor U12769 (N_12769,N_11413,N_11058);
nand U12770 (N_12770,N_11142,N_11079);
and U12771 (N_12771,N_11937,N_11291);
nand U12772 (N_12772,N_11877,N_11370);
nor U12773 (N_12773,N_11850,N_10788);
xor U12774 (N_12774,N_11507,N_11974);
and U12775 (N_12775,N_11467,N_11856);
nand U12776 (N_12776,N_11403,N_11160);
nor U12777 (N_12777,N_11605,N_10715);
or U12778 (N_12778,N_11983,N_11704);
xor U12779 (N_12779,N_10799,N_11275);
or U12780 (N_12780,N_11006,N_10677);
or U12781 (N_12781,N_11555,N_11064);
nor U12782 (N_12782,N_11016,N_11976);
nor U12783 (N_12783,N_11719,N_10911);
xor U12784 (N_12784,N_11047,N_10826);
nand U12785 (N_12785,N_10956,N_10545);
nand U12786 (N_12786,N_11940,N_11400);
nand U12787 (N_12787,N_11316,N_11877);
and U12788 (N_12788,N_11326,N_11977);
or U12789 (N_12789,N_10799,N_10622);
and U12790 (N_12790,N_10650,N_11406);
nand U12791 (N_12791,N_10744,N_10971);
nor U12792 (N_12792,N_10548,N_11355);
and U12793 (N_12793,N_10782,N_10691);
or U12794 (N_12794,N_10678,N_10549);
xor U12795 (N_12795,N_10798,N_11487);
or U12796 (N_12796,N_11061,N_11330);
nor U12797 (N_12797,N_11531,N_11749);
nand U12798 (N_12798,N_11779,N_10789);
xor U12799 (N_12799,N_11584,N_11375);
nand U12800 (N_12800,N_11286,N_11647);
nor U12801 (N_12801,N_11205,N_10838);
nor U12802 (N_12802,N_11223,N_10504);
or U12803 (N_12803,N_11820,N_11398);
or U12804 (N_12804,N_11510,N_11532);
nor U12805 (N_12805,N_10916,N_11573);
and U12806 (N_12806,N_10719,N_11281);
and U12807 (N_12807,N_11655,N_11238);
nand U12808 (N_12808,N_11488,N_11640);
or U12809 (N_12809,N_11102,N_11058);
or U12810 (N_12810,N_10837,N_11439);
xor U12811 (N_12811,N_10658,N_11445);
or U12812 (N_12812,N_11787,N_11899);
and U12813 (N_12813,N_11441,N_11780);
nor U12814 (N_12814,N_11365,N_10609);
or U12815 (N_12815,N_11704,N_11769);
or U12816 (N_12816,N_11026,N_11175);
nor U12817 (N_12817,N_11865,N_11782);
nor U12818 (N_12818,N_11358,N_11299);
or U12819 (N_12819,N_11180,N_11603);
xnor U12820 (N_12820,N_11382,N_10863);
xor U12821 (N_12821,N_11462,N_10981);
xor U12822 (N_12822,N_11452,N_11825);
or U12823 (N_12823,N_10861,N_10683);
and U12824 (N_12824,N_11281,N_10762);
nor U12825 (N_12825,N_11255,N_11682);
nor U12826 (N_12826,N_10861,N_11746);
and U12827 (N_12827,N_11414,N_11649);
nor U12828 (N_12828,N_11761,N_10573);
nor U12829 (N_12829,N_10974,N_11843);
or U12830 (N_12830,N_11185,N_11149);
nor U12831 (N_12831,N_10623,N_10797);
and U12832 (N_12832,N_10726,N_11294);
nand U12833 (N_12833,N_11229,N_11228);
nor U12834 (N_12834,N_11731,N_11459);
and U12835 (N_12835,N_11405,N_11487);
xor U12836 (N_12836,N_11224,N_11080);
or U12837 (N_12837,N_10780,N_10903);
nand U12838 (N_12838,N_11251,N_10938);
or U12839 (N_12839,N_11288,N_11172);
or U12840 (N_12840,N_11624,N_10637);
nor U12841 (N_12841,N_11206,N_11422);
nand U12842 (N_12842,N_10966,N_11629);
or U12843 (N_12843,N_11109,N_11668);
nand U12844 (N_12844,N_10653,N_11576);
nor U12845 (N_12845,N_10688,N_10535);
xor U12846 (N_12846,N_11404,N_11586);
xnor U12847 (N_12847,N_10600,N_11529);
nand U12848 (N_12848,N_11380,N_11878);
or U12849 (N_12849,N_11289,N_11456);
xnor U12850 (N_12850,N_11952,N_11609);
nand U12851 (N_12851,N_11421,N_11701);
xnor U12852 (N_12852,N_11550,N_11479);
and U12853 (N_12853,N_11667,N_10550);
nand U12854 (N_12854,N_11095,N_11456);
xnor U12855 (N_12855,N_10619,N_11368);
xnor U12856 (N_12856,N_11304,N_11464);
or U12857 (N_12857,N_11904,N_11815);
nor U12858 (N_12858,N_11531,N_10933);
xnor U12859 (N_12859,N_11883,N_11432);
nor U12860 (N_12860,N_11728,N_10944);
or U12861 (N_12861,N_11817,N_11353);
and U12862 (N_12862,N_11209,N_11457);
xnor U12863 (N_12863,N_11155,N_11704);
nor U12864 (N_12864,N_10850,N_11422);
nor U12865 (N_12865,N_10533,N_11537);
xor U12866 (N_12866,N_11940,N_10680);
xor U12867 (N_12867,N_10934,N_10720);
or U12868 (N_12868,N_11246,N_11023);
and U12869 (N_12869,N_11475,N_11979);
and U12870 (N_12870,N_11978,N_11918);
or U12871 (N_12871,N_10940,N_11789);
or U12872 (N_12872,N_10892,N_11595);
nor U12873 (N_12873,N_11085,N_10581);
xor U12874 (N_12874,N_11844,N_11646);
and U12875 (N_12875,N_10918,N_11396);
and U12876 (N_12876,N_11792,N_11500);
and U12877 (N_12877,N_11039,N_10769);
xnor U12878 (N_12878,N_10500,N_11980);
or U12879 (N_12879,N_11927,N_11680);
xor U12880 (N_12880,N_11903,N_11886);
nor U12881 (N_12881,N_11498,N_11146);
and U12882 (N_12882,N_10552,N_10996);
nand U12883 (N_12883,N_11439,N_10910);
nor U12884 (N_12884,N_10636,N_11881);
xnor U12885 (N_12885,N_11965,N_11249);
nor U12886 (N_12886,N_11893,N_10804);
and U12887 (N_12887,N_11567,N_11151);
or U12888 (N_12888,N_10776,N_11024);
or U12889 (N_12889,N_11832,N_11597);
or U12890 (N_12890,N_11630,N_11734);
xnor U12891 (N_12891,N_10672,N_10526);
or U12892 (N_12892,N_11927,N_11019);
xnor U12893 (N_12893,N_11445,N_10559);
nor U12894 (N_12894,N_11507,N_11595);
and U12895 (N_12895,N_10888,N_10538);
xor U12896 (N_12896,N_11249,N_11739);
or U12897 (N_12897,N_11409,N_10974);
xnor U12898 (N_12898,N_10503,N_11185);
and U12899 (N_12899,N_11559,N_11473);
xor U12900 (N_12900,N_11500,N_10951);
nor U12901 (N_12901,N_10699,N_11367);
nand U12902 (N_12902,N_11496,N_10910);
xor U12903 (N_12903,N_11533,N_10594);
and U12904 (N_12904,N_11059,N_11282);
nor U12905 (N_12905,N_11192,N_10545);
nor U12906 (N_12906,N_11256,N_11555);
or U12907 (N_12907,N_11304,N_10797);
or U12908 (N_12908,N_11825,N_11375);
nand U12909 (N_12909,N_10990,N_10820);
nand U12910 (N_12910,N_11175,N_10813);
nand U12911 (N_12911,N_10524,N_11416);
or U12912 (N_12912,N_11485,N_11974);
nor U12913 (N_12913,N_11425,N_10849);
or U12914 (N_12914,N_10920,N_11628);
or U12915 (N_12915,N_11757,N_11111);
or U12916 (N_12916,N_10503,N_11350);
and U12917 (N_12917,N_11243,N_10643);
nor U12918 (N_12918,N_10557,N_11230);
nor U12919 (N_12919,N_11052,N_11227);
xnor U12920 (N_12920,N_11774,N_10859);
nand U12921 (N_12921,N_10705,N_10821);
or U12922 (N_12922,N_11129,N_11320);
nor U12923 (N_12923,N_11268,N_10743);
xor U12924 (N_12924,N_11605,N_11221);
nor U12925 (N_12925,N_11168,N_10817);
nor U12926 (N_12926,N_11371,N_11435);
xor U12927 (N_12927,N_11134,N_11955);
xnor U12928 (N_12928,N_10839,N_11304);
xnor U12929 (N_12929,N_10600,N_10711);
nand U12930 (N_12930,N_10594,N_10512);
or U12931 (N_12931,N_11903,N_11391);
nor U12932 (N_12932,N_11183,N_11134);
nor U12933 (N_12933,N_11092,N_10693);
xnor U12934 (N_12934,N_10920,N_11360);
xor U12935 (N_12935,N_11128,N_11182);
or U12936 (N_12936,N_10958,N_11318);
and U12937 (N_12937,N_11067,N_11962);
xor U12938 (N_12938,N_10742,N_10980);
nand U12939 (N_12939,N_11040,N_10887);
nor U12940 (N_12940,N_11194,N_10521);
nor U12941 (N_12941,N_10918,N_10942);
and U12942 (N_12942,N_11965,N_11714);
or U12943 (N_12943,N_11032,N_11875);
nor U12944 (N_12944,N_11006,N_11642);
xnor U12945 (N_12945,N_10634,N_10636);
nand U12946 (N_12946,N_10925,N_11931);
nand U12947 (N_12947,N_10849,N_11103);
nor U12948 (N_12948,N_10849,N_11347);
xor U12949 (N_12949,N_11324,N_11561);
nand U12950 (N_12950,N_11983,N_10779);
nor U12951 (N_12951,N_11136,N_10847);
xor U12952 (N_12952,N_10919,N_11947);
or U12953 (N_12953,N_11586,N_10673);
nand U12954 (N_12954,N_11796,N_11159);
xor U12955 (N_12955,N_10966,N_10863);
or U12956 (N_12956,N_10982,N_11171);
nand U12957 (N_12957,N_11797,N_11856);
xnor U12958 (N_12958,N_11178,N_11341);
or U12959 (N_12959,N_10729,N_11523);
and U12960 (N_12960,N_10854,N_11895);
or U12961 (N_12961,N_10635,N_10659);
nor U12962 (N_12962,N_11006,N_10740);
nand U12963 (N_12963,N_11130,N_11018);
nand U12964 (N_12964,N_10981,N_11171);
nand U12965 (N_12965,N_10594,N_10588);
xor U12966 (N_12966,N_10743,N_11881);
xnor U12967 (N_12967,N_10715,N_11942);
and U12968 (N_12968,N_11316,N_10827);
nor U12969 (N_12969,N_10519,N_11833);
xor U12970 (N_12970,N_11863,N_11396);
xnor U12971 (N_12971,N_11767,N_10571);
and U12972 (N_12972,N_11369,N_11933);
or U12973 (N_12973,N_11055,N_11386);
nand U12974 (N_12974,N_11132,N_11049);
nor U12975 (N_12975,N_11467,N_11405);
nor U12976 (N_12976,N_10963,N_10695);
and U12977 (N_12977,N_11962,N_10847);
or U12978 (N_12978,N_11065,N_11288);
and U12979 (N_12979,N_11544,N_10514);
nand U12980 (N_12980,N_10577,N_10910);
xor U12981 (N_12981,N_11731,N_11363);
xor U12982 (N_12982,N_11827,N_11941);
nor U12983 (N_12983,N_10843,N_11715);
nand U12984 (N_12984,N_10771,N_11368);
xnor U12985 (N_12985,N_11408,N_11235);
nand U12986 (N_12986,N_11233,N_11651);
or U12987 (N_12987,N_11790,N_11359);
xnor U12988 (N_12988,N_11906,N_11339);
nand U12989 (N_12989,N_11501,N_11866);
nor U12990 (N_12990,N_11708,N_11930);
or U12991 (N_12991,N_11793,N_11133);
nand U12992 (N_12992,N_11277,N_11333);
or U12993 (N_12993,N_11793,N_11016);
xnor U12994 (N_12994,N_11815,N_11596);
nand U12995 (N_12995,N_11054,N_11871);
and U12996 (N_12996,N_10607,N_10883);
nor U12997 (N_12997,N_11247,N_10736);
nand U12998 (N_12998,N_11407,N_11484);
and U12999 (N_12999,N_11137,N_10897);
nand U13000 (N_13000,N_10979,N_11608);
nor U13001 (N_13001,N_11110,N_11237);
and U13002 (N_13002,N_10971,N_10791);
or U13003 (N_13003,N_10621,N_11599);
xor U13004 (N_13004,N_10852,N_10639);
nor U13005 (N_13005,N_11605,N_11188);
nor U13006 (N_13006,N_11595,N_11536);
nand U13007 (N_13007,N_11243,N_11146);
nand U13008 (N_13008,N_10874,N_11217);
and U13009 (N_13009,N_10620,N_10562);
nor U13010 (N_13010,N_11590,N_11545);
nor U13011 (N_13011,N_10966,N_10689);
nand U13012 (N_13012,N_11254,N_11997);
nand U13013 (N_13013,N_11069,N_11276);
xor U13014 (N_13014,N_11322,N_11663);
nand U13015 (N_13015,N_11068,N_11042);
xor U13016 (N_13016,N_11945,N_10567);
and U13017 (N_13017,N_11906,N_11182);
xor U13018 (N_13018,N_11970,N_10773);
and U13019 (N_13019,N_11722,N_11038);
nor U13020 (N_13020,N_10692,N_10946);
or U13021 (N_13021,N_10718,N_10627);
xor U13022 (N_13022,N_11290,N_10524);
nor U13023 (N_13023,N_11601,N_11649);
xor U13024 (N_13024,N_10670,N_11740);
xnor U13025 (N_13025,N_10539,N_10681);
nand U13026 (N_13026,N_11607,N_11656);
xor U13027 (N_13027,N_11590,N_10680);
and U13028 (N_13028,N_10766,N_11086);
and U13029 (N_13029,N_11357,N_11337);
and U13030 (N_13030,N_11409,N_11471);
nor U13031 (N_13031,N_11712,N_11114);
xnor U13032 (N_13032,N_11962,N_10563);
nor U13033 (N_13033,N_11515,N_11137);
or U13034 (N_13034,N_11269,N_11323);
and U13035 (N_13035,N_10809,N_11139);
nor U13036 (N_13036,N_10602,N_11517);
nor U13037 (N_13037,N_11870,N_10958);
nor U13038 (N_13038,N_10755,N_11683);
or U13039 (N_13039,N_10940,N_10989);
nor U13040 (N_13040,N_11280,N_11214);
nor U13041 (N_13041,N_10996,N_11991);
nand U13042 (N_13042,N_10534,N_10900);
nand U13043 (N_13043,N_11339,N_10678);
xor U13044 (N_13044,N_11802,N_10757);
nor U13045 (N_13045,N_11877,N_11023);
xor U13046 (N_13046,N_10598,N_11599);
or U13047 (N_13047,N_11810,N_11783);
nor U13048 (N_13048,N_10955,N_11459);
nor U13049 (N_13049,N_10671,N_11428);
xnor U13050 (N_13050,N_11542,N_10535);
nand U13051 (N_13051,N_11407,N_11570);
xor U13052 (N_13052,N_11431,N_11057);
xnor U13053 (N_13053,N_11660,N_11386);
nor U13054 (N_13054,N_11058,N_10687);
xnor U13055 (N_13055,N_10814,N_10736);
or U13056 (N_13056,N_11531,N_10776);
xnor U13057 (N_13057,N_11999,N_11765);
nand U13058 (N_13058,N_11121,N_11594);
nor U13059 (N_13059,N_11084,N_10938);
xor U13060 (N_13060,N_10719,N_10595);
nor U13061 (N_13061,N_10891,N_10668);
nand U13062 (N_13062,N_10977,N_11821);
xor U13063 (N_13063,N_11321,N_11120);
xor U13064 (N_13064,N_10790,N_10724);
and U13065 (N_13065,N_11065,N_11003);
nor U13066 (N_13066,N_11391,N_10679);
and U13067 (N_13067,N_10783,N_11109);
and U13068 (N_13068,N_10665,N_11058);
nand U13069 (N_13069,N_11924,N_11263);
and U13070 (N_13070,N_11858,N_11298);
and U13071 (N_13071,N_11771,N_11504);
nor U13072 (N_13072,N_11474,N_10985);
or U13073 (N_13073,N_11936,N_11352);
nand U13074 (N_13074,N_11941,N_11095);
and U13075 (N_13075,N_11225,N_10816);
nand U13076 (N_13076,N_11762,N_11847);
or U13077 (N_13077,N_10565,N_11756);
or U13078 (N_13078,N_11027,N_10912);
and U13079 (N_13079,N_10789,N_11995);
and U13080 (N_13080,N_11149,N_11575);
nand U13081 (N_13081,N_11903,N_10506);
or U13082 (N_13082,N_11052,N_10591);
or U13083 (N_13083,N_11908,N_11500);
nor U13084 (N_13084,N_11457,N_11822);
and U13085 (N_13085,N_11074,N_11484);
and U13086 (N_13086,N_11631,N_10709);
nand U13087 (N_13087,N_11428,N_11020);
xnor U13088 (N_13088,N_11333,N_10750);
or U13089 (N_13089,N_11819,N_10856);
nor U13090 (N_13090,N_10691,N_10952);
nor U13091 (N_13091,N_11110,N_10744);
and U13092 (N_13092,N_11708,N_11601);
nor U13093 (N_13093,N_11518,N_11252);
and U13094 (N_13094,N_10724,N_11489);
or U13095 (N_13095,N_11909,N_10771);
and U13096 (N_13096,N_10883,N_11967);
nand U13097 (N_13097,N_11764,N_11278);
or U13098 (N_13098,N_10581,N_11870);
and U13099 (N_13099,N_11275,N_11784);
nor U13100 (N_13100,N_11508,N_10541);
xnor U13101 (N_13101,N_11062,N_10981);
xor U13102 (N_13102,N_10983,N_10659);
nand U13103 (N_13103,N_11692,N_10779);
or U13104 (N_13104,N_10811,N_11847);
nand U13105 (N_13105,N_11575,N_10576);
nor U13106 (N_13106,N_10955,N_11918);
nand U13107 (N_13107,N_11519,N_11391);
nor U13108 (N_13108,N_10843,N_11900);
or U13109 (N_13109,N_11422,N_11268);
nand U13110 (N_13110,N_10845,N_10507);
nor U13111 (N_13111,N_10937,N_10986);
nand U13112 (N_13112,N_11634,N_11132);
nor U13113 (N_13113,N_10631,N_11547);
and U13114 (N_13114,N_10517,N_11478);
and U13115 (N_13115,N_11136,N_10747);
nand U13116 (N_13116,N_11612,N_11568);
xor U13117 (N_13117,N_11235,N_11742);
nand U13118 (N_13118,N_10864,N_11794);
xor U13119 (N_13119,N_10962,N_10918);
nand U13120 (N_13120,N_11181,N_10962);
and U13121 (N_13121,N_11026,N_10921);
and U13122 (N_13122,N_10574,N_11398);
or U13123 (N_13123,N_10602,N_11430);
or U13124 (N_13124,N_11846,N_11911);
or U13125 (N_13125,N_11473,N_11226);
nor U13126 (N_13126,N_11417,N_11514);
or U13127 (N_13127,N_10587,N_11822);
or U13128 (N_13128,N_10989,N_11215);
and U13129 (N_13129,N_11836,N_11231);
nand U13130 (N_13130,N_10547,N_10738);
and U13131 (N_13131,N_11563,N_11486);
nor U13132 (N_13132,N_10913,N_10989);
nor U13133 (N_13133,N_10715,N_11407);
xor U13134 (N_13134,N_11426,N_11138);
and U13135 (N_13135,N_11128,N_10534);
xor U13136 (N_13136,N_10597,N_11062);
or U13137 (N_13137,N_11298,N_11512);
nor U13138 (N_13138,N_11410,N_10532);
and U13139 (N_13139,N_11292,N_11723);
and U13140 (N_13140,N_11096,N_11634);
xnor U13141 (N_13141,N_11559,N_11741);
or U13142 (N_13142,N_10519,N_11711);
xor U13143 (N_13143,N_11689,N_10596);
or U13144 (N_13144,N_11575,N_11530);
xnor U13145 (N_13145,N_11069,N_11725);
and U13146 (N_13146,N_10648,N_11251);
and U13147 (N_13147,N_10553,N_11701);
or U13148 (N_13148,N_10653,N_11402);
nand U13149 (N_13149,N_11484,N_10660);
nor U13150 (N_13150,N_11689,N_10711);
nand U13151 (N_13151,N_10655,N_10579);
xor U13152 (N_13152,N_11149,N_11616);
and U13153 (N_13153,N_11488,N_10977);
or U13154 (N_13154,N_10686,N_10830);
and U13155 (N_13155,N_11882,N_11670);
xnor U13156 (N_13156,N_11870,N_10721);
or U13157 (N_13157,N_10707,N_10937);
nand U13158 (N_13158,N_11151,N_11111);
nand U13159 (N_13159,N_11573,N_11537);
and U13160 (N_13160,N_11733,N_11433);
nor U13161 (N_13161,N_11188,N_11346);
nor U13162 (N_13162,N_11617,N_11153);
and U13163 (N_13163,N_11085,N_11048);
nand U13164 (N_13164,N_11010,N_11697);
and U13165 (N_13165,N_11848,N_10983);
and U13166 (N_13166,N_10838,N_11808);
or U13167 (N_13167,N_11082,N_11058);
xnor U13168 (N_13168,N_10723,N_11183);
xor U13169 (N_13169,N_11837,N_11559);
and U13170 (N_13170,N_11598,N_11346);
or U13171 (N_13171,N_11039,N_11855);
nor U13172 (N_13172,N_11660,N_11556);
or U13173 (N_13173,N_10952,N_11015);
xor U13174 (N_13174,N_11689,N_10621);
nand U13175 (N_13175,N_11084,N_11286);
or U13176 (N_13176,N_10902,N_11183);
xor U13177 (N_13177,N_10832,N_11876);
and U13178 (N_13178,N_11208,N_11942);
xor U13179 (N_13179,N_11391,N_10771);
nand U13180 (N_13180,N_11110,N_11364);
nor U13181 (N_13181,N_10666,N_11813);
or U13182 (N_13182,N_11587,N_11544);
and U13183 (N_13183,N_11684,N_10633);
xnor U13184 (N_13184,N_11065,N_11645);
and U13185 (N_13185,N_10751,N_11245);
xnor U13186 (N_13186,N_11835,N_11130);
and U13187 (N_13187,N_11874,N_11550);
and U13188 (N_13188,N_10644,N_10910);
nor U13189 (N_13189,N_11718,N_11276);
xnor U13190 (N_13190,N_10515,N_10675);
and U13191 (N_13191,N_11349,N_10683);
xnor U13192 (N_13192,N_11661,N_10896);
and U13193 (N_13193,N_10787,N_10586);
nor U13194 (N_13194,N_11869,N_11276);
and U13195 (N_13195,N_10997,N_11445);
nor U13196 (N_13196,N_11575,N_11714);
nor U13197 (N_13197,N_11159,N_10662);
nor U13198 (N_13198,N_11912,N_11131);
nand U13199 (N_13199,N_11112,N_11011);
xor U13200 (N_13200,N_11508,N_11832);
or U13201 (N_13201,N_11750,N_10503);
xnor U13202 (N_13202,N_10691,N_10878);
nand U13203 (N_13203,N_11596,N_11823);
and U13204 (N_13204,N_11853,N_10716);
xnor U13205 (N_13205,N_11289,N_10853);
or U13206 (N_13206,N_11849,N_11157);
xor U13207 (N_13207,N_10616,N_11209);
nand U13208 (N_13208,N_11360,N_10596);
and U13209 (N_13209,N_10757,N_10768);
xor U13210 (N_13210,N_10607,N_11051);
or U13211 (N_13211,N_11058,N_11422);
xor U13212 (N_13212,N_10532,N_10765);
or U13213 (N_13213,N_11270,N_10649);
or U13214 (N_13214,N_11090,N_10780);
or U13215 (N_13215,N_11569,N_10766);
xnor U13216 (N_13216,N_11149,N_11016);
xor U13217 (N_13217,N_11846,N_11208);
nand U13218 (N_13218,N_11065,N_11619);
nand U13219 (N_13219,N_10927,N_10771);
and U13220 (N_13220,N_10547,N_11597);
nor U13221 (N_13221,N_10557,N_11873);
and U13222 (N_13222,N_11723,N_11118);
and U13223 (N_13223,N_11593,N_10988);
nor U13224 (N_13224,N_11419,N_11585);
xnor U13225 (N_13225,N_10581,N_10970);
nand U13226 (N_13226,N_10688,N_11719);
and U13227 (N_13227,N_11662,N_11129);
nand U13228 (N_13228,N_11489,N_11445);
nor U13229 (N_13229,N_10559,N_10955);
and U13230 (N_13230,N_11185,N_10920);
and U13231 (N_13231,N_10523,N_11977);
nor U13232 (N_13232,N_10707,N_11423);
xnor U13233 (N_13233,N_11196,N_11091);
nor U13234 (N_13234,N_11966,N_11202);
nor U13235 (N_13235,N_10801,N_10755);
or U13236 (N_13236,N_11682,N_11846);
xnor U13237 (N_13237,N_10953,N_11316);
or U13238 (N_13238,N_11240,N_10705);
nor U13239 (N_13239,N_10551,N_11839);
and U13240 (N_13240,N_10829,N_11496);
xor U13241 (N_13241,N_11887,N_10674);
or U13242 (N_13242,N_11862,N_11308);
or U13243 (N_13243,N_11993,N_10780);
nand U13244 (N_13244,N_10722,N_11174);
or U13245 (N_13245,N_10980,N_11569);
or U13246 (N_13246,N_10576,N_10807);
or U13247 (N_13247,N_11595,N_11654);
and U13248 (N_13248,N_11554,N_10569);
nand U13249 (N_13249,N_11192,N_11252);
and U13250 (N_13250,N_11012,N_11889);
and U13251 (N_13251,N_10514,N_10602);
xnor U13252 (N_13252,N_10863,N_10912);
xnor U13253 (N_13253,N_11884,N_11080);
or U13254 (N_13254,N_10574,N_11259);
nor U13255 (N_13255,N_11280,N_10677);
and U13256 (N_13256,N_10807,N_11725);
and U13257 (N_13257,N_11679,N_11733);
and U13258 (N_13258,N_11039,N_11398);
nand U13259 (N_13259,N_11228,N_11393);
or U13260 (N_13260,N_10906,N_10946);
or U13261 (N_13261,N_11853,N_11589);
and U13262 (N_13262,N_11597,N_10602);
nor U13263 (N_13263,N_10788,N_11380);
or U13264 (N_13264,N_10803,N_10854);
or U13265 (N_13265,N_10733,N_10511);
nor U13266 (N_13266,N_11808,N_11642);
nand U13267 (N_13267,N_10580,N_11362);
xor U13268 (N_13268,N_11442,N_11447);
nand U13269 (N_13269,N_11679,N_11418);
nand U13270 (N_13270,N_10812,N_11252);
xor U13271 (N_13271,N_11108,N_11889);
and U13272 (N_13272,N_11529,N_10996);
xor U13273 (N_13273,N_11878,N_11822);
and U13274 (N_13274,N_11043,N_11259);
nand U13275 (N_13275,N_10863,N_11128);
nor U13276 (N_13276,N_11158,N_11481);
nand U13277 (N_13277,N_11358,N_10601);
nor U13278 (N_13278,N_11366,N_11944);
xor U13279 (N_13279,N_11789,N_11610);
and U13280 (N_13280,N_11400,N_11718);
and U13281 (N_13281,N_11930,N_11177);
nor U13282 (N_13282,N_11271,N_10667);
xnor U13283 (N_13283,N_10763,N_10732);
or U13284 (N_13284,N_10749,N_10772);
xor U13285 (N_13285,N_11376,N_10619);
nand U13286 (N_13286,N_11237,N_11349);
and U13287 (N_13287,N_11977,N_11511);
xnor U13288 (N_13288,N_10608,N_11212);
nand U13289 (N_13289,N_11864,N_11445);
xnor U13290 (N_13290,N_11527,N_10647);
xnor U13291 (N_13291,N_10879,N_10529);
nand U13292 (N_13292,N_11405,N_10648);
nand U13293 (N_13293,N_11564,N_11361);
xnor U13294 (N_13294,N_10798,N_11409);
xor U13295 (N_13295,N_10754,N_11915);
and U13296 (N_13296,N_11479,N_11557);
xor U13297 (N_13297,N_11362,N_10810);
and U13298 (N_13298,N_10831,N_11432);
xor U13299 (N_13299,N_10711,N_11869);
or U13300 (N_13300,N_10857,N_11672);
nor U13301 (N_13301,N_11233,N_10597);
xnor U13302 (N_13302,N_10973,N_10746);
nand U13303 (N_13303,N_10984,N_11558);
or U13304 (N_13304,N_10952,N_11318);
xor U13305 (N_13305,N_11347,N_11203);
xnor U13306 (N_13306,N_11936,N_10943);
and U13307 (N_13307,N_11560,N_11084);
nand U13308 (N_13308,N_11322,N_11853);
nand U13309 (N_13309,N_11217,N_11916);
or U13310 (N_13310,N_11695,N_11604);
and U13311 (N_13311,N_10984,N_10514);
and U13312 (N_13312,N_11953,N_11254);
or U13313 (N_13313,N_11776,N_10831);
or U13314 (N_13314,N_11571,N_10638);
nor U13315 (N_13315,N_10892,N_10967);
and U13316 (N_13316,N_11402,N_11729);
or U13317 (N_13317,N_10825,N_11200);
xor U13318 (N_13318,N_11295,N_11254);
xor U13319 (N_13319,N_11827,N_10992);
nor U13320 (N_13320,N_10532,N_11610);
or U13321 (N_13321,N_11416,N_11223);
and U13322 (N_13322,N_11150,N_10544);
and U13323 (N_13323,N_11182,N_10551);
nand U13324 (N_13324,N_10715,N_11667);
and U13325 (N_13325,N_10670,N_11195);
or U13326 (N_13326,N_11546,N_11885);
xnor U13327 (N_13327,N_11259,N_10648);
or U13328 (N_13328,N_11257,N_11826);
xnor U13329 (N_13329,N_10896,N_11201);
nor U13330 (N_13330,N_11156,N_10763);
and U13331 (N_13331,N_10953,N_11929);
or U13332 (N_13332,N_11597,N_11877);
nor U13333 (N_13333,N_11029,N_11891);
and U13334 (N_13334,N_10935,N_11786);
nor U13335 (N_13335,N_11730,N_10947);
xor U13336 (N_13336,N_11813,N_10572);
nor U13337 (N_13337,N_10702,N_11442);
nand U13338 (N_13338,N_10747,N_11071);
xnor U13339 (N_13339,N_11656,N_11933);
or U13340 (N_13340,N_11405,N_10614);
and U13341 (N_13341,N_10550,N_11679);
and U13342 (N_13342,N_10782,N_11589);
nand U13343 (N_13343,N_10707,N_10887);
and U13344 (N_13344,N_11918,N_11485);
nand U13345 (N_13345,N_11458,N_11802);
nand U13346 (N_13346,N_11204,N_11632);
and U13347 (N_13347,N_10817,N_10913);
nor U13348 (N_13348,N_11494,N_11914);
nor U13349 (N_13349,N_11297,N_10586);
xnor U13350 (N_13350,N_11768,N_11001);
and U13351 (N_13351,N_11168,N_11737);
xor U13352 (N_13352,N_10629,N_10946);
and U13353 (N_13353,N_11268,N_11277);
and U13354 (N_13354,N_11564,N_11129);
nand U13355 (N_13355,N_11902,N_11081);
xor U13356 (N_13356,N_10606,N_11511);
nand U13357 (N_13357,N_11463,N_10564);
xor U13358 (N_13358,N_11184,N_10535);
xnor U13359 (N_13359,N_11498,N_11002);
xor U13360 (N_13360,N_11663,N_11040);
xnor U13361 (N_13361,N_10803,N_11634);
nor U13362 (N_13362,N_11476,N_11472);
xor U13363 (N_13363,N_11491,N_10569);
xor U13364 (N_13364,N_10975,N_11327);
xor U13365 (N_13365,N_11146,N_11427);
nand U13366 (N_13366,N_11521,N_10944);
and U13367 (N_13367,N_11001,N_11806);
or U13368 (N_13368,N_10935,N_10527);
xor U13369 (N_13369,N_10520,N_10689);
xnor U13370 (N_13370,N_11366,N_11866);
and U13371 (N_13371,N_11139,N_11754);
xor U13372 (N_13372,N_10560,N_11997);
nor U13373 (N_13373,N_11295,N_11764);
nor U13374 (N_13374,N_10792,N_11675);
nor U13375 (N_13375,N_11983,N_11363);
or U13376 (N_13376,N_10508,N_11740);
and U13377 (N_13377,N_11126,N_11764);
or U13378 (N_13378,N_11408,N_10863);
xor U13379 (N_13379,N_11535,N_11332);
and U13380 (N_13380,N_10681,N_10537);
and U13381 (N_13381,N_11432,N_10550);
nand U13382 (N_13382,N_11775,N_11168);
nor U13383 (N_13383,N_10746,N_11905);
or U13384 (N_13384,N_10723,N_11197);
nor U13385 (N_13385,N_11206,N_11550);
nand U13386 (N_13386,N_11267,N_11455);
or U13387 (N_13387,N_10715,N_10590);
nor U13388 (N_13388,N_10976,N_11390);
xnor U13389 (N_13389,N_10577,N_11820);
nor U13390 (N_13390,N_11019,N_11021);
or U13391 (N_13391,N_11398,N_10710);
nor U13392 (N_13392,N_11307,N_10898);
or U13393 (N_13393,N_10635,N_10540);
xor U13394 (N_13394,N_11421,N_11571);
xnor U13395 (N_13395,N_11112,N_11453);
nor U13396 (N_13396,N_10741,N_10848);
and U13397 (N_13397,N_11235,N_11422);
nand U13398 (N_13398,N_11576,N_10710);
or U13399 (N_13399,N_10536,N_10636);
xor U13400 (N_13400,N_11510,N_11257);
nor U13401 (N_13401,N_10691,N_11825);
xor U13402 (N_13402,N_10701,N_10756);
nand U13403 (N_13403,N_11430,N_10854);
and U13404 (N_13404,N_10775,N_11204);
nor U13405 (N_13405,N_10942,N_11710);
nor U13406 (N_13406,N_11867,N_11448);
or U13407 (N_13407,N_10813,N_11118);
nand U13408 (N_13408,N_10521,N_11757);
nand U13409 (N_13409,N_11809,N_11448);
and U13410 (N_13410,N_11465,N_11501);
xnor U13411 (N_13411,N_10511,N_11208);
and U13412 (N_13412,N_11711,N_11121);
and U13413 (N_13413,N_11207,N_10702);
nor U13414 (N_13414,N_10761,N_10852);
and U13415 (N_13415,N_10607,N_11741);
xor U13416 (N_13416,N_11852,N_11172);
xor U13417 (N_13417,N_10576,N_11877);
or U13418 (N_13418,N_11480,N_11947);
nand U13419 (N_13419,N_11687,N_11783);
and U13420 (N_13420,N_11264,N_11722);
and U13421 (N_13421,N_11740,N_10796);
xnor U13422 (N_13422,N_11337,N_11918);
or U13423 (N_13423,N_10533,N_10970);
xnor U13424 (N_13424,N_10504,N_10800);
or U13425 (N_13425,N_11276,N_10998);
or U13426 (N_13426,N_11652,N_10564);
xnor U13427 (N_13427,N_11136,N_11680);
nand U13428 (N_13428,N_10881,N_11923);
nand U13429 (N_13429,N_11636,N_11218);
and U13430 (N_13430,N_11408,N_11565);
nor U13431 (N_13431,N_10658,N_11801);
xor U13432 (N_13432,N_11924,N_10982);
nor U13433 (N_13433,N_11558,N_11599);
nand U13434 (N_13434,N_11341,N_10547);
nand U13435 (N_13435,N_11576,N_11760);
nand U13436 (N_13436,N_10967,N_11423);
nand U13437 (N_13437,N_10713,N_11213);
or U13438 (N_13438,N_10885,N_11420);
nor U13439 (N_13439,N_11024,N_11276);
nor U13440 (N_13440,N_11345,N_10660);
nand U13441 (N_13441,N_11558,N_11992);
or U13442 (N_13442,N_11980,N_11204);
nor U13443 (N_13443,N_10522,N_11978);
nor U13444 (N_13444,N_11467,N_10903);
nand U13445 (N_13445,N_11352,N_11549);
nand U13446 (N_13446,N_11997,N_11866);
and U13447 (N_13447,N_11605,N_11855);
or U13448 (N_13448,N_11100,N_11404);
or U13449 (N_13449,N_11266,N_11118);
and U13450 (N_13450,N_11235,N_11450);
or U13451 (N_13451,N_11072,N_11617);
or U13452 (N_13452,N_11581,N_11940);
xor U13453 (N_13453,N_11281,N_11087);
or U13454 (N_13454,N_11445,N_10763);
and U13455 (N_13455,N_10822,N_11015);
nor U13456 (N_13456,N_11188,N_10729);
or U13457 (N_13457,N_10797,N_10759);
nor U13458 (N_13458,N_11906,N_11092);
or U13459 (N_13459,N_11670,N_10622);
xnor U13460 (N_13460,N_10789,N_10522);
and U13461 (N_13461,N_10801,N_11818);
and U13462 (N_13462,N_11225,N_11595);
and U13463 (N_13463,N_11402,N_10800);
and U13464 (N_13464,N_11788,N_10684);
and U13465 (N_13465,N_11874,N_10660);
nand U13466 (N_13466,N_10552,N_10564);
nand U13467 (N_13467,N_10835,N_10679);
nor U13468 (N_13468,N_11612,N_11482);
and U13469 (N_13469,N_10906,N_11790);
xnor U13470 (N_13470,N_10700,N_11476);
xnor U13471 (N_13471,N_11043,N_10623);
and U13472 (N_13472,N_10908,N_11180);
xnor U13473 (N_13473,N_11171,N_11161);
nor U13474 (N_13474,N_11205,N_11867);
xnor U13475 (N_13475,N_11990,N_11565);
nor U13476 (N_13476,N_10899,N_11041);
nand U13477 (N_13477,N_10883,N_11792);
and U13478 (N_13478,N_11883,N_11370);
xnor U13479 (N_13479,N_11460,N_11985);
or U13480 (N_13480,N_11099,N_10509);
nor U13481 (N_13481,N_10588,N_10615);
xor U13482 (N_13482,N_11729,N_11707);
and U13483 (N_13483,N_10675,N_11305);
nand U13484 (N_13484,N_11019,N_11872);
nor U13485 (N_13485,N_11574,N_11780);
or U13486 (N_13486,N_11767,N_10620);
xnor U13487 (N_13487,N_11061,N_11305);
and U13488 (N_13488,N_11193,N_11844);
xnor U13489 (N_13489,N_10577,N_10985);
nand U13490 (N_13490,N_11090,N_11532);
nand U13491 (N_13491,N_10689,N_11010);
nor U13492 (N_13492,N_11319,N_11884);
and U13493 (N_13493,N_11970,N_10991);
or U13494 (N_13494,N_11181,N_10505);
and U13495 (N_13495,N_11253,N_11178);
nor U13496 (N_13496,N_10567,N_10611);
and U13497 (N_13497,N_11975,N_11523);
or U13498 (N_13498,N_11496,N_11649);
xnor U13499 (N_13499,N_11277,N_11047);
nor U13500 (N_13500,N_12957,N_12796);
nand U13501 (N_13501,N_12429,N_12004);
and U13502 (N_13502,N_12071,N_12400);
and U13503 (N_13503,N_12402,N_12376);
or U13504 (N_13504,N_12977,N_12146);
nand U13505 (N_13505,N_12663,N_12061);
xnor U13506 (N_13506,N_13036,N_12544);
and U13507 (N_13507,N_13458,N_12394);
nand U13508 (N_13508,N_13177,N_13027);
or U13509 (N_13509,N_13439,N_13258);
nand U13510 (N_13510,N_13499,N_12831);
or U13511 (N_13511,N_12870,N_12139);
or U13512 (N_13512,N_13208,N_12412);
and U13513 (N_13513,N_13248,N_12221);
and U13514 (N_13514,N_12133,N_12558);
nor U13515 (N_13515,N_12587,N_12756);
xnor U13516 (N_13516,N_12742,N_12958);
xor U13517 (N_13517,N_12506,N_13081);
nor U13518 (N_13518,N_13107,N_12880);
nand U13519 (N_13519,N_13199,N_12056);
nor U13520 (N_13520,N_12464,N_12074);
nand U13521 (N_13521,N_13174,N_12382);
and U13522 (N_13522,N_12784,N_12678);
xnor U13523 (N_13523,N_12175,N_12185);
nand U13524 (N_13524,N_13162,N_13183);
and U13525 (N_13525,N_13334,N_12967);
nor U13526 (N_13526,N_13069,N_12703);
and U13527 (N_13527,N_12640,N_12332);
and U13528 (N_13528,N_12241,N_12651);
or U13529 (N_13529,N_13126,N_12953);
xor U13530 (N_13530,N_12954,N_12355);
or U13531 (N_13531,N_12040,N_13382);
or U13532 (N_13532,N_12539,N_12344);
or U13533 (N_13533,N_12530,N_12369);
nand U13534 (N_13534,N_12961,N_12931);
and U13535 (N_13535,N_12285,N_12368);
nor U13536 (N_13536,N_13379,N_13485);
and U13537 (N_13537,N_12391,N_12610);
nor U13538 (N_13538,N_12296,N_13342);
and U13539 (N_13539,N_12821,N_12264);
and U13540 (N_13540,N_13414,N_12916);
or U13541 (N_13541,N_12066,N_13431);
and U13542 (N_13542,N_13156,N_12016);
and U13543 (N_13543,N_13244,N_13321);
or U13544 (N_13544,N_12365,N_12103);
and U13545 (N_13545,N_12037,N_12352);
or U13546 (N_13546,N_12110,N_12462);
or U13547 (N_13547,N_12787,N_13063);
and U13548 (N_13548,N_12050,N_13223);
xor U13549 (N_13549,N_13429,N_12235);
nor U13550 (N_13550,N_13186,N_13021);
or U13551 (N_13551,N_12727,N_12287);
and U13552 (N_13552,N_13221,N_12380);
nor U13553 (N_13553,N_12490,N_12208);
xor U13554 (N_13554,N_13415,N_12997);
xor U13555 (N_13555,N_13189,N_13234);
nor U13556 (N_13556,N_12865,N_13122);
xor U13557 (N_13557,N_13127,N_12613);
and U13558 (N_13558,N_13262,N_12205);
xnor U13559 (N_13559,N_12731,N_12011);
and U13560 (N_13560,N_12006,N_13071);
nand U13561 (N_13561,N_12135,N_12327);
xor U13562 (N_13562,N_13222,N_12533);
nor U13563 (N_13563,N_13190,N_12969);
or U13564 (N_13564,N_12128,N_12802);
and U13565 (N_13565,N_12392,N_12333);
and U13566 (N_13566,N_12407,N_13481);
xor U13567 (N_13567,N_13293,N_12662);
or U13568 (N_13568,N_12196,N_12091);
xor U13569 (N_13569,N_13358,N_12622);
xnor U13570 (N_13570,N_13020,N_12884);
nand U13571 (N_13571,N_12574,N_12976);
or U13572 (N_13572,N_13087,N_12633);
nor U13573 (N_13573,N_12614,N_13067);
xor U13574 (N_13574,N_13076,N_13062);
xor U13575 (N_13575,N_12039,N_12902);
nand U13576 (N_13576,N_12240,N_12960);
or U13577 (N_13577,N_12728,N_12024);
xor U13578 (N_13578,N_13343,N_12090);
xnor U13579 (N_13579,N_13460,N_12409);
nand U13580 (N_13580,N_13236,N_12147);
or U13581 (N_13581,N_12955,N_13375);
or U13582 (N_13582,N_13135,N_12681);
xor U13583 (N_13583,N_13496,N_12435);
or U13584 (N_13584,N_12766,N_12864);
nand U13585 (N_13585,N_13272,N_12151);
nor U13586 (N_13586,N_12304,N_12867);
nor U13587 (N_13587,N_12187,N_13312);
or U13588 (N_13588,N_12142,N_12647);
or U13589 (N_13589,N_13057,N_13104);
or U13590 (N_13590,N_12912,N_13164);
nor U13591 (N_13591,N_13163,N_12941);
or U13592 (N_13592,N_12478,N_12340);
nor U13593 (N_13593,N_12803,N_12087);
and U13594 (N_13594,N_12713,N_13048);
nor U13595 (N_13595,N_12830,N_12975);
xnor U13596 (N_13596,N_13360,N_13184);
or U13597 (N_13597,N_12973,N_12511);
or U13598 (N_13598,N_13191,N_13402);
xnor U13599 (N_13599,N_12566,N_12044);
xor U13600 (N_13600,N_12120,N_12419);
and U13601 (N_13601,N_12126,N_13399);
xor U13602 (N_13602,N_12234,N_12937);
or U13603 (N_13603,N_12768,N_13207);
or U13604 (N_13604,N_12172,N_12670);
xnor U13605 (N_13605,N_12148,N_12914);
nand U13606 (N_13606,N_13477,N_13227);
nand U13607 (N_13607,N_13351,N_12053);
xor U13608 (N_13608,N_12454,N_12008);
or U13609 (N_13609,N_13058,N_12682);
nand U13610 (N_13610,N_12986,N_12620);
and U13611 (N_13611,N_13396,N_13483);
xor U13612 (N_13612,N_13366,N_13279);
or U13613 (N_13613,N_13388,N_12984);
xor U13614 (N_13614,N_12470,N_12580);
nor U13615 (N_13615,N_13344,N_12092);
nand U13616 (N_13616,N_12212,N_13490);
xnor U13617 (N_13617,N_13290,N_13153);
or U13618 (N_13618,N_13369,N_12904);
nor U13619 (N_13619,N_12452,N_12604);
or U13620 (N_13620,N_13406,N_12833);
nor U13621 (N_13621,N_13088,N_12512);
xnor U13622 (N_13622,N_12232,N_12656);
and U13623 (N_13623,N_12164,N_13436);
nand U13624 (N_13624,N_12301,N_13480);
nor U13625 (N_13625,N_12204,N_12117);
and U13626 (N_13626,N_12358,N_13040);
nor U13627 (N_13627,N_13214,N_12137);
nand U13628 (N_13628,N_12105,N_13023);
xor U13629 (N_13629,N_13079,N_12216);
nand U13630 (N_13630,N_12259,N_13130);
or U13631 (N_13631,N_12313,N_12206);
and U13632 (N_13632,N_12900,N_12882);
nand U13633 (N_13633,N_12222,N_12348);
nor U13634 (N_13634,N_12752,N_12238);
nor U13635 (N_13635,N_12167,N_13319);
nor U13636 (N_13636,N_12998,N_13187);
and U13637 (N_13637,N_12992,N_12810);
xor U13638 (N_13638,N_13120,N_13446);
nor U13639 (N_13639,N_12709,N_13347);
xor U13640 (N_13640,N_13111,N_13251);
xnor U13641 (N_13641,N_13075,N_12174);
or U13642 (N_13642,N_12494,N_12085);
nand U13643 (N_13643,N_13484,N_12180);
xnor U13644 (N_13644,N_13387,N_12903);
and U13645 (N_13645,N_12173,N_12388);
nor U13646 (N_13646,N_13148,N_13030);
nor U13647 (N_13647,N_12568,N_12252);
nor U13648 (N_13648,N_12453,N_12168);
nor U13649 (N_13649,N_12588,N_12943);
nor U13650 (N_13650,N_12189,N_13110);
nand U13651 (N_13651,N_12847,N_12022);
and U13652 (N_13652,N_13210,N_12769);
xor U13653 (N_13653,N_12193,N_12537);
xnor U13654 (N_13654,N_12809,N_13171);
or U13655 (N_13655,N_12243,N_12503);
and U13656 (N_13656,N_13447,N_12486);
and U13657 (N_13657,N_12635,N_12165);
nand U13658 (N_13658,N_12226,N_12638);
nand U13659 (N_13659,N_12846,N_13442);
and U13660 (N_13660,N_12561,N_12569);
and U13661 (N_13661,N_13026,N_12772);
or U13662 (N_13662,N_12051,N_12307);
nor U13663 (N_13663,N_13105,N_13314);
or U13664 (N_13664,N_13006,N_12456);
nor U13665 (N_13665,N_12650,N_12602);
xnor U13666 (N_13666,N_12124,N_13381);
and U13667 (N_13667,N_13451,N_12716);
or U13668 (N_13668,N_12156,N_12263);
or U13669 (N_13669,N_12149,N_13359);
and U13670 (N_13670,N_12928,N_12401);
xor U13671 (N_13671,N_12526,N_13330);
xor U13672 (N_13672,N_12999,N_13232);
and U13673 (N_13673,N_12162,N_12542);
and U13674 (N_13674,N_12201,N_13149);
xor U13675 (N_13675,N_13405,N_12956);
and U13676 (N_13676,N_13365,N_12339);
and U13677 (N_13677,N_12191,N_12551);
nand U13678 (N_13678,N_12045,N_12458);
xnor U13679 (N_13679,N_12776,N_13488);
nand U13680 (N_13680,N_13361,N_13091);
or U13681 (N_13681,N_12671,N_12009);
and U13682 (N_13682,N_12321,N_12646);
xor U13683 (N_13683,N_12711,N_12145);
or U13684 (N_13684,N_12118,N_12981);
and U13685 (N_13685,N_12033,N_13452);
nand U13686 (N_13686,N_13425,N_12632);
xor U13687 (N_13687,N_12080,N_12411);
or U13688 (N_13688,N_13012,N_12098);
nand U13689 (N_13689,N_12477,N_12781);
nor U13690 (N_13690,N_12326,N_12143);
nand U13691 (N_13691,N_12379,N_13167);
nor U13692 (N_13692,N_12323,N_13136);
or U13693 (N_13693,N_13470,N_13059);
or U13694 (N_13694,N_12715,N_13464);
xnor U13695 (N_13695,N_12788,N_12480);
nor U13696 (N_13696,N_12269,N_12338);
and U13697 (N_13697,N_12030,N_13169);
nor U13698 (N_13698,N_12334,N_12576);
nor U13699 (N_13699,N_12179,N_12873);
and U13700 (N_13700,N_12808,N_12832);
and U13701 (N_13701,N_12759,N_12209);
xnor U13702 (N_13702,N_13150,N_13422);
and U13703 (N_13703,N_12459,N_12354);
xor U13704 (N_13704,N_12468,N_13082);
nand U13705 (N_13705,N_13175,N_13313);
and U13706 (N_13706,N_13157,N_12306);
xnor U13707 (N_13707,N_12405,N_12994);
xnor U13708 (N_13708,N_12214,N_12607);
or U13709 (N_13709,N_12217,N_13435);
xor U13710 (N_13710,N_12929,N_12723);
xor U13711 (N_13711,N_13173,N_12237);
or U13712 (N_13712,N_13098,N_12911);
xnor U13713 (N_13713,N_13260,N_12730);
or U13714 (N_13714,N_12778,N_12572);
or U13715 (N_13715,N_13336,N_12856);
xor U13716 (N_13716,N_12014,N_12457);
nor U13717 (N_13717,N_12230,N_12186);
or U13718 (N_13718,N_13476,N_12372);
xnor U13719 (N_13719,N_13391,N_13471);
or U13720 (N_13720,N_13498,N_12414);
xor U13721 (N_13721,N_12177,N_12442);
xor U13722 (N_13722,N_12311,N_12905);
nand U13723 (N_13723,N_13225,N_13116);
nand U13724 (N_13724,N_12978,N_12679);
nand U13725 (N_13725,N_12988,N_12774);
nor U13726 (N_13726,N_13095,N_12095);
and U13727 (N_13727,N_12019,N_12842);
or U13728 (N_13728,N_12758,N_13393);
or U13729 (N_13729,N_12780,N_12626);
or U13730 (N_13730,N_12700,N_12293);
nor U13731 (N_13731,N_13441,N_13317);
xor U13732 (N_13732,N_12699,N_13300);
or U13733 (N_13733,N_13253,N_12195);
nor U13734 (N_13734,N_13377,N_12159);
and U13735 (N_13735,N_12826,N_12753);
nand U13736 (N_13736,N_12007,N_12823);
or U13737 (N_13737,N_12274,N_12498);
and U13738 (N_13738,N_13028,N_12406);
and U13739 (N_13739,N_13025,N_13117);
nand U13740 (N_13740,N_12199,N_13403);
nand U13741 (N_13741,N_12879,N_12356);
nor U13742 (N_13742,N_12298,N_13219);
nor U13743 (N_13743,N_12962,N_12347);
nand U13744 (N_13744,N_12852,N_13383);
nand U13745 (N_13745,N_13230,N_12863);
nand U13746 (N_13746,N_12874,N_13401);
nor U13747 (N_13747,N_12262,N_12026);
xor U13748 (N_13748,N_12472,N_12712);
nand U13749 (N_13749,N_12155,N_12972);
or U13750 (N_13750,N_12416,N_12592);
nor U13751 (N_13751,N_12277,N_12343);
or U13752 (N_13752,N_13487,N_13151);
nor U13753 (N_13753,N_13310,N_12265);
or U13754 (N_13754,N_13348,N_12415);
xnor U13755 (N_13755,N_13473,N_12469);
and U13756 (N_13756,N_13008,N_12611);
or U13757 (N_13757,N_13440,N_12390);
nand U13758 (N_13758,N_12331,N_12249);
or U13759 (N_13759,N_12898,N_12946);
nand U13760 (N_13760,N_12673,N_12518);
nor U13761 (N_13761,N_13266,N_13448);
nor U13762 (N_13762,N_12479,N_12844);
nand U13763 (N_13763,N_13017,N_13165);
and U13764 (N_13764,N_13109,N_12325);
nand U13765 (N_13765,N_12005,N_12420);
and U13766 (N_13766,N_12920,N_12102);
or U13767 (N_13767,N_12578,N_12585);
nand U13768 (N_13768,N_12440,N_12163);
or U13769 (N_13769,N_12996,N_13013);
nand U13770 (N_13770,N_12936,N_12793);
or U13771 (N_13771,N_12507,N_13242);
nand U13772 (N_13772,N_12562,N_12595);
and U13773 (N_13773,N_12746,N_13255);
and U13774 (N_13774,N_13418,N_12658);
xnor U13775 (N_13775,N_13323,N_13289);
nor U13776 (N_13776,N_12483,N_13101);
and U13777 (N_13777,N_12229,N_12897);
xnor U13778 (N_13778,N_12528,N_12068);
nand U13779 (N_13779,N_12674,N_12702);
nor U13780 (N_13780,N_12942,N_13096);
and U13781 (N_13781,N_12919,N_13287);
xor U13782 (N_13782,N_12115,N_12247);
nand U13783 (N_13783,N_12465,N_13283);
and U13784 (N_13784,N_12403,N_12218);
nor U13785 (N_13785,N_13426,N_13000);
or U13786 (N_13786,N_12560,N_13265);
or U13787 (N_13787,N_13074,N_12820);
nand U13788 (N_13788,N_12351,N_12603);
or U13789 (N_13789,N_12827,N_12375);
or U13790 (N_13790,N_12303,N_12563);
nand U13791 (N_13791,N_13103,N_13044);
xor U13792 (N_13792,N_13353,N_13131);
nor U13793 (N_13793,N_12686,N_12584);
nand U13794 (N_13794,N_12549,N_12853);
and U13795 (N_13795,N_12575,N_13029);
and U13796 (N_13796,N_13416,N_12282);
and U13797 (N_13797,N_12875,N_12838);
xor U13798 (N_13798,N_12959,N_12529);
and U13799 (N_13799,N_12361,N_12714);
xnor U13800 (N_13800,N_12540,N_13462);
or U13801 (N_13801,N_12745,N_13052);
nor U13802 (N_13802,N_12268,N_12850);
nand U13803 (N_13803,N_12088,N_12485);
xor U13804 (N_13804,N_13297,N_12767);
nor U13805 (N_13805,N_13205,N_13332);
or U13806 (N_13806,N_13072,N_12851);
or U13807 (N_13807,N_13202,N_12619);
xor U13808 (N_13808,N_13302,N_13064);
and U13809 (N_13809,N_12965,N_12600);
and U13810 (N_13810,N_13438,N_12161);
nand U13811 (N_13811,N_12048,N_12719);
or U13812 (N_13812,N_12925,N_12565);
or U13813 (N_13813,N_12461,N_12015);
and U13814 (N_13814,N_13015,N_12178);
xor U13815 (N_13815,N_12691,N_12181);
and U13816 (N_13816,N_12508,N_12707);
or U13817 (N_13817,N_12215,N_12545);
xor U13818 (N_13818,N_12983,N_13065);
nand U13819 (N_13819,N_12108,N_12680);
nand U13820 (N_13820,N_12862,N_12963);
nor U13821 (N_13821,N_13014,N_13491);
nand U13822 (N_13822,N_12913,N_13115);
nand U13823 (N_13823,N_12615,N_13235);
nand U13824 (N_13824,N_13329,N_12939);
nand U13825 (N_13825,N_13413,N_13271);
xnor U13826 (N_13826,N_12608,N_12665);
or U13827 (N_13827,N_12288,N_12096);
and U13828 (N_13828,N_12836,N_12849);
xnor U13829 (N_13829,N_13125,N_12207);
or U13830 (N_13830,N_12063,N_13123);
xor U13831 (N_13831,N_12297,N_12104);
or U13832 (N_13832,N_13245,N_12664);
xor U13833 (N_13833,N_12740,N_12153);
nand U13834 (N_13834,N_12738,N_12131);
nor U13835 (N_13835,N_13482,N_13408);
nor U13836 (N_13836,N_13384,N_12741);
and U13837 (N_13837,N_13182,N_13465);
xor U13838 (N_13838,N_13367,N_13051);
or U13839 (N_13839,N_12233,N_12430);
nor U13840 (N_13840,N_12743,N_12527);
xnor U13841 (N_13841,N_12581,N_12099);
xnor U13842 (N_13842,N_12437,N_12399);
nor U13843 (N_13843,N_13419,N_12076);
nor U13844 (N_13844,N_12038,N_13003);
nor U13845 (N_13845,N_13124,N_12696);
and U13846 (N_13846,N_13019,N_12636);
nand U13847 (N_13847,N_13154,N_12428);
and U13848 (N_13848,N_13363,N_13284);
nand U13849 (N_13849,N_12521,N_12938);
and U13850 (N_13850,N_12718,N_13159);
or U13851 (N_13851,N_12762,N_12089);
xnor U13852 (N_13852,N_12519,N_13263);
nand U13853 (N_13853,N_13032,N_13288);
or U13854 (N_13854,N_12497,N_13309);
nor U13855 (N_13855,N_12493,N_12598);
nor U13856 (N_13856,N_12672,N_13112);
nor U13857 (N_13857,N_12492,N_13392);
xnor U13858 (N_13858,N_12570,N_13385);
and U13859 (N_13859,N_13394,N_13331);
xnor U13860 (N_13860,N_12018,N_12446);
nand U13861 (N_13861,N_12289,N_12735);
nand U13862 (N_13862,N_13291,N_12449);
or U13863 (N_13863,N_12434,N_12641);
nand U13864 (N_13864,N_12889,N_12083);
and U13865 (N_13865,N_12861,N_13145);
nor U13866 (N_13866,N_12476,N_12227);
or U13867 (N_13867,N_13489,N_12097);
nor U13868 (N_13868,N_13276,N_12035);
xor U13869 (N_13869,N_12345,N_12475);
nor U13870 (N_13870,N_13195,N_13412);
and U13871 (N_13871,N_12722,N_13427);
xnor U13872 (N_13872,N_12773,N_12599);
and U13873 (N_13873,N_12499,N_12517);
nand U13874 (N_13874,N_13185,N_12425);
and U13875 (N_13875,N_12123,N_13209);
or U13876 (N_13876,N_13089,N_12654);
nand U13877 (N_13877,N_12628,N_13001);
nor U13878 (N_13878,N_13168,N_12360);
and U13879 (N_13879,N_13108,N_13322);
and U13880 (N_13880,N_12547,N_13224);
nand U13881 (N_13881,N_13172,N_12794);
nor U13882 (N_13882,N_12724,N_13410);
and U13883 (N_13883,N_13469,N_12257);
or U13884 (N_13884,N_12531,N_12447);
nor U13885 (N_13885,N_13400,N_12381);
xnor U13886 (N_13886,N_13229,N_12239);
nand U13887 (N_13887,N_12583,N_12789);
xnor U13888 (N_13888,N_12933,N_12797);
or U13889 (N_13889,N_12384,N_13049);
or U13890 (N_13890,N_12652,N_12374);
xor U13891 (N_13891,N_13445,N_12086);
xor U13892 (N_13892,N_12445,N_12495);
nand U13893 (N_13893,N_12822,N_12819);
xor U13894 (N_13894,N_12166,N_13339);
or U13895 (N_13895,N_13077,N_12272);
nor U13896 (N_13896,N_13100,N_12667);
nand U13897 (N_13897,N_13018,N_12894);
nand U13898 (N_13898,N_12582,N_12859);
nand U13899 (N_13899,N_13233,N_13129);
nand U13900 (N_13900,N_13390,N_12275);
or U13901 (N_13901,N_12049,N_12748);
xor U13902 (N_13902,N_12642,N_13340);
or U13903 (N_13903,N_12036,N_13311);
or U13904 (N_13904,N_12421,N_12127);
xor U13905 (N_13905,N_12386,N_12878);
or U13906 (N_13906,N_12278,N_12467);
nor U13907 (N_13907,N_12502,N_13237);
nand U13908 (N_13908,N_12899,N_12991);
nand U13909 (N_13909,N_13134,N_12330);
nand U13910 (N_13910,N_12021,N_13256);
xor U13911 (N_13911,N_12790,N_13022);
xnor U13912 (N_13912,N_13139,N_13078);
or U13913 (N_13913,N_13099,N_12487);
xnor U13914 (N_13914,N_12775,N_13254);
nand U13915 (N_13915,N_12194,N_13212);
nor U13916 (N_13916,N_13142,N_12591);
nand U13917 (N_13917,N_12786,N_13298);
or U13918 (N_13918,N_12052,N_12130);
nor U13919 (N_13919,N_12660,N_12291);
and U13920 (N_13920,N_12924,N_12012);
xnor U13921 (N_13921,N_12329,N_13411);
nand U13922 (N_13922,N_12107,N_12322);
or U13923 (N_13923,N_12951,N_12064);
or U13924 (N_13924,N_12328,N_12985);
or U13925 (N_13925,N_13243,N_12885);
and U13926 (N_13926,N_12246,N_13454);
xor U13927 (N_13927,N_13324,N_13246);
nor U13928 (N_13928,N_12000,N_12749);
and U13929 (N_13929,N_13166,N_12764);
xor U13930 (N_13930,N_12688,N_12605);
xor U13931 (N_13931,N_13395,N_12706);
nand U13932 (N_13932,N_12557,N_12612);
or U13933 (N_13933,N_12101,N_13325);
nor U13934 (N_13934,N_12947,N_13011);
nand U13935 (N_13935,N_13231,N_13080);
or U13936 (N_13936,N_12136,N_12645);
xor U13937 (N_13937,N_12886,N_13327);
nor U13938 (N_13938,N_12825,N_12708);
and U13939 (N_13939,N_12154,N_12644);
nor U13940 (N_13940,N_12169,N_12152);
xor U13941 (N_13941,N_12245,N_13444);
xnor U13942 (N_13942,N_13315,N_13409);
or U13943 (N_13943,N_12653,N_12661);
nor U13944 (N_13944,N_12944,N_13467);
nand U13945 (N_13945,N_12017,N_12378);
and U13946 (N_13946,N_13090,N_12948);
nor U13947 (N_13947,N_12593,N_12250);
nand U13948 (N_13948,N_12132,N_13270);
nor U13949 (N_13949,N_13362,N_13226);
nand U13950 (N_13950,N_12320,N_13005);
nor U13951 (N_13951,N_12757,N_13220);
xor U13952 (N_13952,N_12283,N_13137);
and U13953 (N_13953,N_12966,N_12763);
or U13954 (N_13954,N_13228,N_12210);
nand U13955 (N_13955,N_12513,N_12455);
xnor U13956 (N_13956,N_13114,N_12460);
nor U13957 (N_13957,N_12890,N_13193);
and U13958 (N_13958,N_13200,N_12798);
nand U13959 (N_13959,N_12029,N_12891);
nand U13960 (N_13960,N_13188,N_12617);
nand U13961 (N_13961,N_12100,N_12777);
and U13962 (N_13962,N_12812,N_12032);
and U13963 (N_13963,N_13397,N_12744);
nor U13964 (N_13964,N_12310,N_12034);
xnor U13965 (N_13965,N_13449,N_12385);
nand U13966 (N_13966,N_12559,N_12726);
xnor U13967 (N_13967,N_13495,N_12505);
and U13968 (N_13968,N_12424,N_12121);
or U13969 (N_13969,N_12639,N_13198);
xor U13970 (N_13970,N_12119,N_12413);
nor U13971 (N_13971,N_13341,N_12625);
xor U13972 (N_13972,N_13303,N_13016);
or U13973 (N_13973,N_12276,N_12341);
or U13974 (N_13974,N_12279,N_13128);
xor U13975 (N_13975,N_13038,N_12281);
or U13976 (N_13976,N_13034,N_12556);
nor U13977 (N_13977,N_12448,N_12292);
or U13978 (N_13978,N_12466,N_13463);
and U13979 (N_13979,N_12267,N_13264);
or U13980 (N_13980,N_12111,N_12990);
or U13981 (N_13981,N_12655,N_13380);
xnor U13982 (N_13982,N_12949,N_13474);
xnor U13983 (N_13983,N_13144,N_12041);
xor U13984 (N_13984,N_12266,N_12138);
nand U13985 (N_13985,N_12940,N_13143);
and U13986 (N_13986,N_12701,N_12536);
nor U13987 (N_13987,N_13170,N_12028);
nand U13988 (N_13988,N_12729,N_12950);
nand U13989 (N_13989,N_12077,N_13035);
xor U13990 (N_13990,N_13196,N_12396);
xor U13991 (N_13991,N_12171,N_12979);
xnor U13992 (N_13992,N_12150,N_12188);
and U13993 (N_13993,N_13466,N_12698);
nor U13994 (N_13994,N_12463,N_13268);
and U13995 (N_13995,N_13345,N_12002);
nor U13996 (N_13996,N_13478,N_12782);
nand U13997 (N_13997,N_12922,N_12971);
or U13998 (N_13998,N_13430,N_12754);
nor U13999 (N_13999,N_12106,N_12197);
nand U14000 (N_14000,N_12223,N_12860);
or U14001 (N_14001,N_12750,N_12273);
nor U14002 (N_14002,N_12324,N_12869);
xnor U14003 (N_14003,N_13453,N_12945);
and U14004 (N_14004,N_12302,N_13073);
nor U14005 (N_14005,N_12829,N_13056);
and U14006 (N_14006,N_13121,N_12824);
and U14007 (N_14007,N_12312,N_12710);
or U14008 (N_14008,N_13372,N_13320);
nor U14009 (N_14009,N_13178,N_12523);
and U14010 (N_14010,N_12771,N_12450);
nor U14011 (N_14011,N_12160,N_12815);
nor U14012 (N_14012,N_13141,N_13370);
xnor U14013 (N_14013,N_12065,N_13346);
nor U14014 (N_14014,N_12319,N_12251);
nor U14015 (N_14015,N_12573,N_12244);
nor U14016 (N_14016,N_12935,N_12550);
xnor U14017 (N_14017,N_12631,N_13031);
or U14018 (N_14018,N_12982,N_13285);
or U14019 (N_14019,N_12845,N_12546);
nor U14020 (N_14020,N_13434,N_12801);
and U14021 (N_14021,N_12255,N_13179);
and U14022 (N_14022,N_13060,N_13295);
nor U14023 (N_14023,N_13181,N_12634);
xor U14024 (N_14024,N_12923,N_12057);
xnor U14025 (N_14025,N_12284,N_12439);
or U14026 (N_14026,N_12915,N_13140);
nand U14027 (N_14027,N_13437,N_13216);
nand U14028 (N_14028,N_12818,N_12785);
nor U14029 (N_14029,N_12501,N_12687);
and U14030 (N_14030,N_12980,N_12734);
and U14031 (N_14031,N_12871,N_12256);
xnor U14032 (N_14032,N_12926,N_13450);
and U14033 (N_14033,N_13455,N_12995);
and U14034 (N_14034,N_12432,N_12514);
nand U14035 (N_14035,N_13269,N_13118);
and U14036 (N_14036,N_12286,N_12888);
nand U14037 (N_14037,N_12474,N_12917);
nand U14038 (N_14038,N_12444,N_12349);
nor U14039 (N_14039,N_13119,N_13252);
or U14040 (N_14040,N_12122,N_13138);
and U14041 (N_14041,N_12337,N_12489);
or U14042 (N_14042,N_12363,N_12657);
or U14043 (N_14043,N_12059,N_12770);
xnor U14044 (N_14044,N_13371,N_12877);
and U14045 (N_14045,N_13217,N_12834);
and U14046 (N_14046,N_12868,N_12705);
nor U14047 (N_14047,N_13368,N_12261);
nand U14048 (N_14048,N_12659,N_13155);
nand U14049 (N_14049,N_13146,N_12370);
nand U14050 (N_14050,N_12553,N_13386);
nor U14051 (N_14051,N_12042,N_12300);
xnor U14052 (N_14052,N_13066,N_12589);
nor U14053 (N_14053,N_13428,N_13278);
or U14054 (N_14054,N_13420,N_12073);
nor U14055 (N_14055,N_13161,N_12488);
and U14056 (N_14056,N_12564,N_13055);
nand U14057 (N_14057,N_13257,N_13356);
or U14058 (N_14058,N_12404,N_12848);
and U14059 (N_14059,N_12952,N_13147);
nor U14060 (N_14060,N_12484,N_12114);
nor U14061 (N_14061,N_12970,N_13204);
nand U14062 (N_14062,N_13357,N_12535);
nand U14063 (N_14063,N_13050,N_12228);
nand U14064 (N_14064,N_13176,N_13010);
or U14065 (N_14065,N_12677,N_12579);
and U14066 (N_14066,N_12318,N_12906);
and U14067 (N_14067,N_13249,N_12157);
xor U14068 (N_14068,N_12436,N_12316);
or U14069 (N_14069,N_12525,N_13355);
and U14070 (N_14070,N_13417,N_12141);
or U14071 (N_14071,N_12364,N_12075);
xor U14072 (N_14072,N_12047,N_12907);
and U14073 (N_14073,N_13404,N_12020);
and U14074 (N_14074,N_12586,N_12046);
xnor U14075 (N_14075,N_13113,N_12084);
nand U14076 (N_14076,N_13093,N_12013);
nor U14077 (N_14077,N_12854,N_12027);
and U14078 (N_14078,N_12236,N_13197);
nand U14079 (N_14079,N_13456,N_12471);
and U14080 (N_14080,N_13004,N_12067);
nor U14081 (N_14081,N_12079,N_12176);
nor U14082 (N_14082,N_13033,N_12609);
or U14083 (N_14083,N_12577,N_13497);
or U14084 (N_14084,N_13280,N_13338);
nor U14085 (N_14085,N_12695,N_12621);
and U14086 (N_14086,N_12335,N_12828);
nor U14087 (N_14087,N_13304,N_13286);
and U14088 (N_14088,N_12082,N_12383);
nand U14089 (N_14089,N_12253,N_12666);
nand U14090 (N_14090,N_12140,N_13424);
or U14091 (N_14091,N_12112,N_12520);
xor U14092 (N_14092,N_12733,N_12438);
or U14093 (N_14093,N_12817,N_12184);
xnor U14094 (N_14094,N_12792,N_12366);
nand U14095 (N_14095,N_12725,N_13261);
xor U14096 (N_14096,N_13250,N_12721);
or U14097 (N_14097,N_12134,N_12760);
nand U14098 (N_14098,N_13335,N_12552);
xor U14099 (N_14099,N_12807,N_12353);
nand U14100 (N_14100,N_12315,N_13492);
xor U14101 (N_14101,N_12901,N_12192);
nand U14102 (N_14102,N_12555,N_12417);
nor U14103 (N_14103,N_12630,N_12025);
nor U14104 (N_14104,N_13218,N_12078);
nand U14105 (N_14105,N_12685,N_13468);
nor U14106 (N_14106,N_12387,N_12183);
and U14107 (N_14107,N_12918,N_12813);
and U14108 (N_14108,N_12213,N_12491);
or U14109 (N_14109,N_12795,N_12554);
and U14110 (N_14110,N_12765,N_12129);
nand U14111 (N_14111,N_13158,N_12843);
nand U14112 (N_14112,N_12624,N_12800);
or U14113 (N_14113,N_12055,N_12254);
nand U14114 (N_14114,N_12500,N_12974);
nor U14115 (N_14115,N_12692,N_13267);
nor U14116 (N_14116,N_13349,N_12887);
nor U14117 (N_14117,N_13043,N_13299);
nor U14118 (N_14118,N_13432,N_13132);
or U14119 (N_14119,N_13152,N_12693);
and U14120 (N_14120,N_12910,N_12081);
xor U14121 (N_14121,N_12294,N_12840);
and U14122 (N_14122,N_13054,N_12431);
nand U14123 (N_14123,N_12805,N_12336);
nor U14124 (N_14124,N_13457,N_12377);
and U14125 (N_14125,N_13192,N_13086);
nor U14126 (N_14126,N_12516,N_13083);
xor U14127 (N_14127,N_12893,N_13337);
and U14128 (N_14128,N_12504,N_12422);
nand U14129 (N_14129,N_12876,N_12410);
nor U14130 (N_14130,N_13277,N_13486);
nand U14131 (N_14131,N_12606,N_12858);
or U14132 (N_14132,N_13407,N_12543);
xor U14133 (N_14133,N_12811,N_12932);
xor U14134 (N_14134,N_12094,N_13459);
nand U14135 (N_14135,N_12737,N_12541);
or U14136 (N_14136,N_13068,N_12314);
xor U14137 (N_14137,N_12220,N_12806);
xor U14138 (N_14138,N_12720,N_13041);
xnor U14139 (N_14139,N_12676,N_12704);
or U14140 (N_14140,N_12690,N_13106);
nor U14141 (N_14141,N_12072,N_12398);
nand U14142 (N_14142,N_12909,N_12855);
xnor U14143 (N_14143,N_12934,N_12144);
nor U14144 (N_14144,N_13133,N_12441);
and U14145 (N_14145,N_12054,N_13102);
or U14146 (N_14146,N_13273,N_13326);
nand U14147 (N_14147,N_12616,N_12623);
nand U14148 (N_14148,N_12567,N_13042);
and U14149 (N_14149,N_12571,N_12683);
or U14150 (N_14150,N_12755,N_12839);
nor U14151 (N_14151,N_12883,N_13007);
or U14152 (N_14152,N_12023,N_12697);
or U14153 (N_14153,N_13475,N_12203);
nor U14154 (N_14154,N_13316,N_13046);
nand U14155 (N_14155,N_12643,N_12993);
xnor U14156 (N_14156,N_13306,N_12443);
xor U14157 (N_14157,N_12231,N_12736);
and U14158 (N_14158,N_12732,N_12684);
nand U14159 (N_14159,N_12116,N_12694);
nor U14160 (N_14160,N_12481,N_12747);
nor U14161 (N_14161,N_12224,N_12473);
or U14162 (N_14162,N_12689,N_13494);
xnor U14163 (N_14163,N_13241,N_12482);
nor U14164 (N_14164,N_12423,N_13423);
nand U14165 (N_14165,N_13398,N_13364);
xnor U14166 (N_14166,N_12290,N_13239);
nand U14167 (N_14167,N_12675,N_12271);
and U14168 (N_14168,N_12751,N_13053);
or U14169 (N_14169,N_12804,N_12200);
or U14170 (N_14170,N_12739,N_12669);
and U14171 (N_14171,N_13247,N_12921);
and U14172 (N_14172,N_13307,N_12927);
and U14173 (N_14173,N_12389,N_12964);
nand U14174 (N_14174,N_13213,N_13292);
xnor U14175 (N_14175,N_12295,N_13037);
xor U14176 (N_14176,N_12373,N_12408);
xor U14177 (N_14177,N_12841,N_12534);
nor U14178 (N_14178,N_12892,N_13160);
or U14179 (N_14179,N_12857,N_12001);
and U14180 (N_14180,N_12305,N_13211);
or U14181 (N_14181,N_12367,N_12113);
xor U14182 (N_14182,N_13024,N_13308);
nor U14183 (N_14183,N_12371,N_13092);
nor U14184 (N_14184,N_13421,N_12280);
nor U14185 (N_14185,N_13296,N_12866);
nand U14186 (N_14186,N_13238,N_13240);
nand U14187 (N_14187,N_13328,N_12211);
or U14188 (N_14188,N_13045,N_13203);
nand U14189 (N_14189,N_12590,N_13206);
or U14190 (N_14190,N_13002,N_12601);
and U14191 (N_14191,N_12346,N_12835);
nand U14192 (N_14192,N_13097,N_12717);
and U14193 (N_14193,N_12668,N_12637);
xnor U14194 (N_14194,N_12597,N_12629);
nor U14195 (N_14195,N_13479,N_12426);
nand U14196 (N_14196,N_13374,N_12837);
nor U14197 (N_14197,N_12627,N_13350);
xnor U14198 (N_14198,N_12895,N_12393);
nand U14199 (N_14199,N_12814,N_12594);
xnor U14200 (N_14200,N_13094,N_12968);
or U14201 (N_14201,N_12791,N_13294);
nand U14202 (N_14202,N_12596,N_12308);
xor U14203 (N_14203,N_12060,N_12258);
nand U14204 (N_14204,N_13282,N_12270);
nand U14205 (N_14205,N_13039,N_12248);
and U14206 (N_14206,N_13070,N_12010);
xnor U14207 (N_14207,N_12109,N_12125);
nor U14208 (N_14208,N_13493,N_13259);
xor U14209 (N_14209,N_12170,N_13373);
nand U14210 (N_14210,N_12043,N_13201);
nand U14211 (N_14211,N_12058,N_12989);
xor U14212 (N_14212,N_12260,N_13047);
nor U14213 (N_14213,N_12350,N_12069);
xor U14214 (N_14214,N_12987,N_13472);
and U14215 (N_14215,N_12182,N_13194);
nor U14216 (N_14216,N_12357,N_12872);
and U14217 (N_14217,N_13376,N_12031);
or U14218 (N_14218,N_13318,N_12427);
nand U14219 (N_14219,N_12496,N_13301);
nor U14220 (N_14220,N_12783,N_12799);
and U14221 (N_14221,N_12816,N_13333);
or U14222 (N_14222,N_13215,N_13354);
or U14223 (N_14223,N_12433,N_12532);
and U14224 (N_14224,N_12761,N_12359);
nand U14225 (N_14225,N_12397,N_13378);
and U14226 (N_14226,N_12649,N_12538);
nand U14227 (N_14227,N_13084,N_12648);
nor U14228 (N_14228,N_13061,N_13274);
nor U14229 (N_14229,N_12930,N_13433);
and U14230 (N_14230,N_12908,N_13281);
and U14231 (N_14231,N_12342,N_13275);
xor U14232 (N_14232,N_12510,N_13009);
and U14233 (N_14233,N_12225,N_12509);
nand U14234 (N_14234,N_13443,N_12190);
nor U14235 (N_14235,N_12317,N_12618);
and U14236 (N_14236,N_12242,N_13352);
nand U14237 (N_14237,N_13389,N_12093);
xor U14238 (N_14238,N_12524,N_12395);
nand U14239 (N_14239,N_12062,N_12418);
nand U14240 (N_14240,N_12779,N_12309);
or U14241 (N_14241,N_12548,N_12202);
nor U14242 (N_14242,N_13180,N_12003);
nand U14243 (N_14243,N_12362,N_12219);
nor U14244 (N_14244,N_12158,N_12522);
nor U14245 (N_14245,N_12896,N_12515);
and U14246 (N_14246,N_12198,N_12881);
or U14247 (N_14247,N_13305,N_12070);
or U14248 (N_14248,N_13461,N_12451);
nand U14249 (N_14249,N_12299,N_13085);
and U14250 (N_14250,N_12761,N_13411);
nor U14251 (N_14251,N_13225,N_12277);
nor U14252 (N_14252,N_12718,N_12307);
xnor U14253 (N_14253,N_12777,N_12106);
and U14254 (N_14254,N_12123,N_13153);
or U14255 (N_14255,N_13426,N_12718);
nor U14256 (N_14256,N_12938,N_12066);
nand U14257 (N_14257,N_13133,N_12599);
nor U14258 (N_14258,N_13123,N_12319);
nor U14259 (N_14259,N_13018,N_13059);
or U14260 (N_14260,N_13305,N_13317);
or U14261 (N_14261,N_12994,N_13108);
nor U14262 (N_14262,N_13492,N_12693);
or U14263 (N_14263,N_13316,N_12320);
xor U14264 (N_14264,N_12034,N_12616);
xnor U14265 (N_14265,N_12219,N_12431);
nand U14266 (N_14266,N_13034,N_12102);
nand U14267 (N_14267,N_13126,N_13018);
xor U14268 (N_14268,N_13336,N_13457);
nand U14269 (N_14269,N_13272,N_13280);
nand U14270 (N_14270,N_12490,N_12832);
xor U14271 (N_14271,N_13306,N_13451);
and U14272 (N_14272,N_12096,N_12614);
xor U14273 (N_14273,N_13369,N_12144);
nor U14274 (N_14274,N_12819,N_13019);
and U14275 (N_14275,N_12717,N_12797);
xnor U14276 (N_14276,N_12374,N_13029);
nand U14277 (N_14277,N_13240,N_12410);
nand U14278 (N_14278,N_13122,N_12460);
nand U14279 (N_14279,N_13424,N_12127);
and U14280 (N_14280,N_12632,N_12332);
and U14281 (N_14281,N_13442,N_13047);
nand U14282 (N_14282,N_13203,N_12188);
xor U14283 (N_14283,N_12208,N_13054);
xnor U14284 (N_14284,N_12276,N_13137);
nor U14285 (N_14285,N_12089,N_12500);
and U14286 (N_14286,N_12801,N_13126);
nand U14287 (N_14287,N_12066,N_12996);
nand U14288 (N_14288,N_13129,N_12702);
nand U14289 (N_14289,N_13287,N_12043);
nor U14290 (N_14290,N_12195,N_13020);
nor U14291 (N_14291,N_13004,N_12682);
and U14292 (N_14292,N_13013,N_13385);
or U14293 (N_14293,N_12471,N_13040);
or U14294 (N_14294,N_13370,N_12844);
nand U14295 (N_14295,N_12872,N_12410);
nor U14296 (N_14296,N_12792,N_13095);
nor U14297 (N_14297,N_12327,N_13256);
and U14298 (N_14298,N_13446,N_12772);
xor U14299 (N_14299,N_12381,N_13064);
and U14300 (N_14300,N_12807,N_13272);
xor U14301 (N_14301,N_12852,N_13331);
xnor U14302 (N_14302,N_12107,N_13276);
nor U14303 (N_14303,N_12107,N_13493);
nor U14304 (N_14304,N_12299,N_12932);
and U14305 (N_14305,N_12737,N_12580);
or U14306 (N_14306,N_12457,N_12265);
xnor U14307 (N_14307,N_13033,N_13058);
nand U14308 (N_14308,N_13348,N_12183);
and U14309 (N_14309,N_13300,N_13424);
nand U14310 (N_14310,N_13352,N_12505);
or U14311 (N_14311,N_13101,N_12106);
xnor U14312 (N_14312,N_13273,N_12347);
nor U14313 (N_14313,N_13299,N_13100);
nor U14314 (N_14314,N_12768,N_13292);
nand U14315 (N_14315,N_13471,N_12441);
nor U14316 (N_14316,N_12322,N_13315);
nand U14317 (N_14317,N_12284,N_12543);
nand U14318 (N_14318,N_12980,N_12297);
nand U14319 (N_14319,N_13266,N_12384);
or U14320 (N_14320,N_13413,N_13398);
xnor U14321 (N_14321,N_12297,N_13099);
xor U14322 (N_14322,N_12042,N_12260);
xor U14323 (N_14323,N_12740,N_12421);
or U14324 (N_14324,N_13299,N_13133);
nand U14325 (N_14325,N_12625,N_12189);
nand U14326 (N_14326,N_12423,N_12540);
nor U14327 (N_14327,N_12811,N_12061);
and U14328 (N_14328,N_13065,N_12662);
or U14329 (N_14329,N_12377,N_12661);
xor U14330 (N_14330,N_13169,N_12245);
or U14331 (N_14331,N_12773,N_13098);
nor U14332 (N_14332,N_12249,N_12147);
nor U14333 (N_14333,N_13187,N_13462);
or U14334 (N_14334,N_12560,N_12107);
and U14335 (N_14335,N_12627,N_12626);
nor U14336 (N_14336,N_13498,N_12621);
xnor U14337 (N_14337,N_13336,N_12741);
and U14338 (N_14338,N_12126,N_13264);
nand U14339 (N_14339,N_12769,N_12977);
and U14340 (N_14340,N_12542,N_13062);
xor U14341 (N_14341,N_13479,N_12167);
or U14342 (N_14342,N_12446,N_12851);
or U14343 (N_14343,N_12316,N_12162);
xnor U14344 (N_14344,N_12493,N_12211);
and U14345 (N_14345,N_12353,N_13197);
and U14346 (N_14346,N_12031,N_12017);
nand U14347 (N_14347,N_13030,N_12706);
nand U14348 (N_14348,N_12271,N_13018);
nor U14349 (N_14349,N_12298,N_12141);
or U14350 (N_14350,N_13056,N_12280);
xor U14351 (N_14351,N_13483,N_12947);
xor U14352 (N_14352,N_12379,N_12326);
and U14353 (N_14353,N_13467,N_13189);
or U14354 (N_14354,N_12901,N_12686);
and U14355 (N_14355,N_12049,N_13372);
xor U14356 (N_14356,N_13240,N_12441);
nor U14357 (N_14357,N_12660,N_12784);
or U14358 (N_14358,N_12083,N_12180);
nor U14359 (N_14359,N_13340,N_12919);
or U14360 (N_14360,N_12761,N_12850);
xnor U14361 (N_14361,N_12035,N_12147);
and U14362 (N_14362,N_13026,N_12052);
nor U14363 (N_14363,N_13438,N_12585);
and U14364 (N_14364,N_12246,N_13474);
and U14365 (N_14365,N_13141,N_12552);
nor U14366 (N_14366,N_12623,N_13285);
nor U14367 (N_14367,N_13220,N_12024);
or U14368 (N_14368,N_12554,N_12598);
and U14369 (N_14369,N_13476,N_12048);
or U14370 (N_14370,N_12078,N_12247);
or U14371 (N_14371,N_12410,N_12562);
or U14372 (N_14372,N_12160,N_12537);
xor U14373 (N_14373,N_12400,N_12970);
or U14374 (N_14374,N_12100,N_12451);
nand U14375 (N_14375,N_12983,N_12250);
nor U14376 (N_14376,N_12602,N_12241);
nor U14377 (N_14377,N_12924,N_13238);
nor U14378 (N_14378,N_12762,N_13311);
or U14379 (N_14379,N_12590,N_12311);
nor U14380 (N_14380,N_12474,N_12654);
and U14381 (N_14381,N_13383,N_12382);
and U14382 (N_14382,N_13408,N_13325);
xor U14383 (N_14383,N_12520,N_12728);
xor U14384 (N_14384,N_12238,N_12966);
xor U14385 (N_14385,N_12878,N_12687);
and U14386 (N_14386,N_13429,N_13069);
or U14387 (N_14387,N_13360,N_12475);
nand U14388 (N_14388,N_12570,N_12758);
nand U14389 (N_14389,N_13032,N_13456);
nand U14390 (N_14390,N_13093,N_12518);
nor U14391 (N_14391,N_12503,N_12761);
nor U14392 (N_14392,N_13098,N_12316);
and U14393 (N_14393,N_12920,N_13149);
and U14394 (N_14394,N_13094,N_12312);
or U14395 (N_14395,N_12747,N_12584);
nor U14396 (N_14396,N_12841,N_12729);
nor U14397 (N_14397,N_12625,N_12380);
or U14398 (N_14398,N_13019,N_12831);
xnor U14399 (N_14399,N_13473,N_13105);
and U14400 (N_14400,N_12205,N_12456);
xnor U14401 (N_14401,N_13016,N_13042);
xor U14402 (N_14402,N_13482,N_13160);
and U14403 (N_14403,N_12822,N_12846);
and U14404 (N_14404,N_12741,N_13129);
nand U14405 (N_14405,N_13380,N_13260);
nor U14406 (N_14406,N_12741,N_12774);
nor U14407 (N_14407,N_13343,N_12651);
nand U14408 (N_14408,N_12966,N_13338);
nand U14409 (N_14409,N_12746,N_13364);
nor U14410 (N_14410,N_13288,N_12493);
nand U14411 (N_14411,N_12807,N_12172);
nor U14412 (N_14412,N_13006,N_13000);
and U14413 (N_14413,N_12195,N_13288);
nand U14414 (N_14414,N_12351,N_13157);
or U14415 (N_14415,N_13498,N_12009);
nand U14416 (N_14416,N_12298,N_13179);
or U14417 (N_14417,N_12686,N_12570);
nand U14418 (N_14418,N_13405,N_12706);
or U14419 (N_14419,N_12338,N_12616);
and U14420 (N_14420,N_12332,N_12160);
nand U14421 (N_14421,N_12776,N_13432);
nand U14422 (N_14422,N_13106,N_12925);
or U14423 (N_14423,N_12450,N_13106);
nand U14424 (N_14424,N_12294,N_13275);
and U14425 (N_14425,N_12678,N_12623);
and U14426 (N_14426,N_13045,N_12015);
nor U14427 (N_14427,N_13276,N_12400);
and U14428 (N_14428,N_13063,N_12046);
and U14429 (N_14429,N_12190,N_12924);
xor U14430 (N_14430,N_12817,N_13070);
and U14431 (N_14431,N_12669,N_13347);
and U14432 (N_14432,N_13239,N_12643);
or U14433 (N_14433,N_13163,N_12686);
xor U14434 (N_14434,N_13103,N_13071);
nor U14435 (N_14435,N_12646,N_13337);
and U14436 (N_14436,N_12668,N_13491);
or U14437 (N_14437,N_13309,N_12364);
xor U14438 (N_14438,N_12335,N_12537);
xor U14439 (N_14439,N_13330,N_12994);
and U14440 (N_14440,N_12053,N_12065);
nand U14441 (N_14441,N_12393,N_12135);
nor U14442 (N_14442,N_12269,N_13243);
xnor U14443 (N_14443,N_13108,N_12888);
nor U14444 (N_14444,N_12100,N_12763);
xor U14445 (N_14445,N_12331,N_12372);
or U14446 (N_14446,N_12752,N_12675);
and U14447 (N_14447,N_12152,N_12269);
nand U14448 (N_14448,N_12191,N_12465);
xor U14449 (N_14449,N_12796,N_13257);
nor U14450 (N_14450,N_12110,N_12035);
and U14451 (N_14451,N_12126,N_12436);
nand U14452 (N_14452,N_13242,N_12386);
and U14453 (N_14453,N_12808,N_12509);
nor U14454 (N_14454,N_13307,N_13250);
or U14455 (N_14455,N_12120,N_12453);
xor U14456 (N_14456,N_12557,N_12999);
and U14457 (N_14457,N_13295,N_12100);
and U14458 (N_14458,N_12456,N_13014);
nor U14459 (N_14459,N_13388,N_12505);
nand U14460 (N_14460,N_12733,N_12604);
nor U14461 (N_14461,N_13432,N_13074);
nand U14462 (N_14462,N_13429,N_12665);
and U14463 (N_14463,N_13337,N_13165);
xor U14464 (N_14464,N_12568,N_12276);
xor U14465 (N_14465,N_13317,N_12849);
or U14466 (N_14466,N_13222,N_13088);
or U14467 (N_14467,N_12710,N_12009);
nand U14468 (N_14468,N_13093,N_12679);
nor U14469 (N_14469,N_12288,N_12914);
nand U14470 (N_14470,N_13325,N_13076);
nor U14471 (N_14471,N_12156,N_13178);
nor U14472 (N_14472,N_13038,N_13174);
nand U14473 (N_14473,N_12911,N_12343);
nand U14474 (N_14474,N_13376,N_12363);
nor U14475 (N_14475,N_12147,N_12780);
or U14476 (N_14476,N_12710,N_12727);
nor U14477 (N_14477,N_12260,N_12230);
and U14478 (N_14478,N_13153,N_12811);
nor U14479 (N_14479,N_13395,N_12935);
xor U14480 (N_14480,N_12361,N_12970);
and U14481 (N_14481,N_12465,N_12329);
nand U14482 (N_14482,N_12695,N_13181);
nor U14483 (N_14483,N_12873,N_12885);
or U14484 (N_14484,N_12351,N_12359);
nand U14485 (N_14485,N_12809,N_13441);
or U14486 (N_14486,N_12163,N_12296);
or U14487 (N_14487,N_12755,N_13335);
nand U14488 (N_14488,N_12691,N_12985);
nor U14489 (N_14489,N_13117,N_12212);
nor U14490 (N_14490,N_13073,N_13200);
or U14491 (N_14491,N_13469,N_12125);
nand U14492 (N_14492,N_13391,N_12869);
nor U14493 (N_14493,N_12940,N_12452);
or U14494 (N_14494,N_12376,N_12616);
nor U14495 (N_14495,N_12878,N_13332);
nor U14496 (N_14496,N_12800,N_12664);
and U14497 (N_14497,N_12545,N_12539);
nor U14498 (N_14498,N_12052,N_12376);
xnor U14499 (N_14499,N_12470,N_13389);
or U14500 (N_14500,N_12701,N_12681);
xnor U14501 (N_14501,N_12338,N_12765);
or U14502 (N_14502,N_12413,N_12076);
and U14503 (N_14503,N_12791,N_12832);
nor U14504 (N_14504,N_12210,N_12375);
xor U14505 (N_14505,N_13138,N_13145);
nand U14506 (N_14506,N_12969,N_12056);
and U14507 (N_14507,N_12724,N_12389);
and U14508 (N_14508,N_12223,N_12988);
nand U14509 (N_14509,N_12966,N_12772);
nor U14510 (N_14510,N_13294,N_12085);
or U14511 (N_14511,N_13393,N_12488);
nand U14512 (N_14512,N_12518,N_12386);
xor U14513 (N_14513,N_12812,N_12436);
or U14514 (N_14514,N_12603,N_12225);
or U14515 (N_14515,N_12300,N_12752);
nor U14516 (N_14516,N_13088,N_13131);
xnor U14517 (N_14517,N_12212,N_12035);
xnor U14518 (N_14518,N_12048,N_13464);
or U14519 (N_14519,N_12931,N_12405);
or U14520 (N_14520,N_12571,N_12264);
and U14521 (N_14521,N_12176,N_13130);
and U14522 (N_14522,N_12086,N_12624);
and U14523 (N_14523,N_13309,N_13193);
nand U14524 (N_14524,N_12120,N_12377);
and U14525 (N_14525,N_12421,N_12795);
nor U14526 (N_14526,N_13344,N_13421);
or U14527 (N_14527,N_13211,N_13158);
xor U14528 (N_14528,N_12327,N_13047);
or U14529 (N_14529,N_12943,N_12889);
nand U14530 (N_14530,N_12045,N_13091);
and U14531 (N_14531,N_12519,N_12043);
xnor U14532 (N_14532,N_12671,N_13082);
xor U14533 (N_14533,N_12409,N_13241);
nand U14534 (N_14534,N_12916,N_13290);
nor U14535 (N_14535,N_12996,N_13239);
or U14536 (N_14536,N_12878,N_12216);
and U14537 (N_14537,N_12960,N_12432);
xor U14538 (N_14538,N_12867,N_12177);
xnor U14539 (N_14539,N_12665,N_12334);
or U14540 (N_14540,N_12692,N_13314);
xor U14541 (N_14541,N_12296,N_13480);
nand U14542 (N_14542,N_13429,N_12111);
and U14543 (N_14543,N_13419,N_12114);
and U14544 (N_14544,N_12305,N_12112);
xor U14545 (N_14545,N_13084,N_13230);
or U14546 (N_14546,N_13371,N_13325);
nor U14547 (N_14547,N_12049,N_12722);
xor U14548 (N_14548,N_12649,N_13122);
xnor U14549 (N_14549,N_12793,N_12192);
xnor U14550 (N_14550,N_12745,N_12105);
nand U14551 (N_14551,N_13397,N_12558);
nand U14552 (N_14552,N_12413,N_13007);
or U14553 (N_14553,N_13067,N_12102);
xnor U14554 (N_14554,N_13174,N_13367);
nor U14555 (N_14555,N_12366,N_12085);
or U14556 (N_14556,N_12801,N_12006);
or U14557 (N_14557,N_13334,N_12498);
xor U14558 (N_14558,N_13437,N_12088);
or U14559 (N_14559,N_12878,N_13380);
or U14560 (N_14560,N_13407,N_13015);
nor U14561 (N_14561,N_12713,N_12651);
xor U14562 (N_14562,N_13269,N_12765);
and U14563 (N_14563,N_12418,N_13447);
nand U14564 (N_14564,N_13361,N_12376);
xnor U14565 (N_14565,N_12607,N_12289);
nand U14566 (N_14566,N_12544,N_13144);
xor U14567 (N_14567,N_12727,N_13374);
or U14568 (N_14568,N_12782,N_12679);
nand U14569 (N_14569,N_12669,N_12363);
or U14570 (N_14570,N_12141,N_12304);
xor U14571 (N_14571,N_12042,N_13456);
and U14572 (N_14572,N_13401,N_13465);
and U14573 (N_14573,N_12600,N_12409);
and U14574 (N_14574,N_13370,N_13209);
xor U14575 (N_14575,N_12583,N_13011);
nor U14576 (N_14576,N_12643,N_12296);
xor U14577 (N_14577,N_12776,N_12684);
nor U14578 (N_14578,N_13013,N_13027);
or U14579 (N_14579,N_12787,N_13285);
nor U14580 (N_14580,N_12980,N_13078);
or U14581 (N_14581,N_12420,N_12376);
nand U14582 (N_14582,N_12963,N_12364);
nand U14583 (N_14583,N_13470,N_12942);
nand U14584 (N_14584,N_12725,N_13022);
and U14585 (N_14585,N_12126,N_12816);
xor U14586 (N_14586,N_12249,N_12833);
and U14587 (N_14587,N_13020,N_12751);
xnor U14588 (N_14588,N_12867,N_12741);
or U14589 (N_14589,N_12013,N_12083);
nand U14590 (N_14590,N_12549,N_12227);
and U14591 (N_14591,N_13391,N_12704);
xnor U14592 (N_14592,N_13445,N_13340);
nor U14593 (N_14593,N_12986,N_12946);
or U14594 (N_14594,N_12770,N_12847);
nor U14595 (N_14595,N_13430,N_12807);
xor U14596 (N_14596,N_13490,N_12661);
and U14597 (N_14597,N_13200,N_13096);
nand U14598 (N_14598,N_12456,N_13493);
nand U14599 (N_14599,N_12184,N_13053);
xnor U14600 (N_14600,N_13244,N_12583);
nand U14601 (N_14601,N_13300,N_12115);
or U14602 (N_14602,N_13253,N_12846);
xor U14603 (N_14603,N_13405,N_12686);
and U14604 (N_14604,N_12852,N_12578);
nor U14605 (N_14605,N_12554,N_12402);
and U14606 (N_14606,N_13324,N_12076);
or U14607 (N_14607,N_12143,N_12768);
or U14608 (N_14608,N_12223,N_13177);
nand U14609 (N_14609,N_13199,N_12238);
nor U14610 (N_14610,N_12313,N_12516);
xnor U14611 (N_14611,N_13240,N_12078);
xor U14612 (N_14612,N_12101,N_12461);
and U14613 (N_14613,N_12208,N_13056);
nor U14614 (N_14614,N_12097,N_12433);
nor U14615 (N_14615,N_13113,N_12190);
xor U14616 (N_14616,N_12972,N_12896);
and U14617 (N_14617,N_13119,N_13420);
nor U14618 (N_14618,N_12538,N_12568);
and U14619 (N_14619,N_13118,N_13206);
and U14620 (N_14620,N_12241,N_12668);
nor U14621 (N_14621,N_13128,N_13014);
nand U14622 (N_14622,N_13074,N_13301);
and U14623 (N_14623,N_13469,N_12060);
nor U14624 (N_14624,N_12085,N_12683);
and U14625 (N_14625,N_12878,N_12402);
and U14626 (N_14626,N_13261,N_12010);
xor U14627 (N_14627,N_12430,N_12505);
xnor U14628 (N_14628,N_12204,N_13156);
or U14629 (N_14629,N_13461,N_12964);
nor U14630 (N_14630,N_13052,N_12567);
or U14631 (N_14631,N_12625,N_12509);
or U14632 (N_14632,N_12316,N_12151);
xnor U14633 (N_14633,N_12570,N_12043);
nor U14634 (N_14634,N_12699,N_12594);
or U14635 (N_14635,N_12870,N_13465);
nor U14636 (N_14636,N_12378,N_13043);
xor U14637 (N_14637,N_13085,N_13447);
nor U14638 (N_14638,N_12087,N_12332);
or U14639 (N_14639,N_13209,N_12511);
and U14640 (N_14640,N_12317,N_12885);
and U14641 (N_14641,N_12339,N_12472);
nor U14642 (N_14642,N_13269,N_13194);
or U14643 (N_14643,N_12570,N_12915);
nor U14644 (N_14644,N_13411,N_12564);
and U14645 (N_14645,N_12421,N_13492);
and U14646 (N_14646,N_13057,N_12304);
nand U14647 (N_14647,N_12802,N_12626);
and U14648 (N_14648,N_13281,N_12681);
and U14649 (N_14649,N_13248,N_13361);
nor U14650 (N_14650,N_13262,N_12128);
or U14651 (N_14651,N_13256,N_12500);
or U14652 (N_14652,N_12203,N_12289);
nand U14653 (N_14653,N_12032,N_13377);
nand U14654 (N_14654,N_12659,N_12071);
or U14655 (N_14655,N_13141,N_13417);
and U14656 (N_14656,N_13414,N_12154);
and U14657 (N_14657,N_13397,N_13424);
and U14658 (N_14658,N_13480,N_13248);
or U14659 (N_14659,N_12743,N_13388);
nand U14660 (N_14660,N_12399,N_12530);
nor U14661 (N_14661,N_12449,N_12400);
nor U14662 (N_14662,N_13364,N_12598);
xnor U14663 (N_14663,N_12557,N_12672);
xor U14664 (N_14664,N_13419,N_13407);
or U14665 (N_14665,N_12983,N_12791);
and U14666 (N_14666,N_12735,N_12831);
or U14667 (N_14667,N_12349,N_12608);
or U14668 (N_14668,N_12101,N_12793);
xnor U14669 (N_14669,N_12389,N_12574);
or U14670 (N_14670,N_12259,N_12360);
or U14671 (N_14671,N_12808,N_12716);
nand U14672 (N_14672,N_12285,N_12144);
and U14673 (N_14673,N_12927,N_13073);
or U14674 (N_14674,N_12220,N_12235);
xor U14675 (N_14675,N_13187,N_12482);
xnor U14676 (N_14676,N_12288,N_12756);
nor U14677 (N_14677,N_13395,N_13341);
nor U14678 (N_14678,N_13199,N_12752);
xnor U14679 (N_14679,N_12717,N_13460);
and U14680 (N_14680,N_13074,N_12257);
xor U14681 (N_14681,N_12309,N_12767);
xor U14682 (N_14682,N_12862,N_12166);
and U14683 (N_14683,N_12673,N_12825);
or U14684 (N_14684,N_12348,N_13214);
nor U14685 (N_14685,N_12400,N_13038);
nor U14686 (N_14686,N_12197,N_13414);
and U14687 (N_14687,N_12939,N_13183);
or U14688 (N_14688,N_12158,N_12467);
xor U14689 (N_14689,N_13446,N_12190);
and U14690 (N_14690,N_13266,N_12645);
or U14691 (N_14691,N_12993,N_12240);
and U14692 (N_14692,N_13093,N_12675);
and U14693 (N_14693,N_12558,N_13456);
and U14694 (N_14694,N_13476,N_13294);
xnor U14695 (N_14695,N_12958,N_12114);
or U14696 (N_14696,N_12885,N_12283);
nor U14697 (N_14697,N_12704,N_12632);
and U14698 (N_14698,N_12095,N_12652);
or U14699 (N_14699,N_12298,N_12466);
and U14700 (N_14700,N_13034,N_12701);
nand U14701 (N_14701,N_12978,N_12137);
nand U14702 (N_14702,N_12974,N_13374);
xnor U14703 (N_14703,N_12379,N_12535);
or U14704 (N_14704,N_12047,N_13443);
nand U14705 (N_14705,N_13183,N_12236);
and U14706 (N_14706,N_12879,N_13201);
and U14707 (N_14707,N_12318,N_13040);
xnor U14708 (N_14708,N_12936,N_12969);
xor U14709 (N_14709,N_12931,N_12784);
and U14710 (N_14710,N_12683,N_12493);
nor U14711 (N_14711,N_12755,N_12622);
and U14712 (N_14712,N_12242,N_12137);
nand U14713 (N_14713,N_13243,N_12299);
and U14714 (N_14714,N_13040,N_13353);
or U14715 (N_14715,N_12471,N_12909);
xnor U14716 (N_14716,N_13081,N_12131);
nand U14717 (N_14717,N_12769,N_12686);
nand U14718 (N_14718,N_13220,N_12507);
xnor U14719 (N_14719,N_13039,N_13492);
xor U14720 (N_14720,N_13120,N_13167);
nor U14721 (N_14721,N_12012,N_12776);
and U14722 (N_14722,N_13459,N_12272);
or U14723 (N_14723,N_13123,N_13066);
or U14724 (N_14724,N_12396,N_12079);
nand U14725 (N_14725,N_13277,N_13099);
nand U14726 (N_14726,N_12289,N_12013);
xnor U14727 (N_14727,N_12306,N_12196);
or U14728 (N_14728,N_13188,N_12308);
and U14729 (N_14729,N_12598,N_12342);
nand U14730 (N_14730,N_12625,N_12121);
or U14731 (N_14731,N_12877,N_13210);
nand U14732 (N_14732,N_12608,N_12642);
xor U14733 (N_14733,N_12788,N_12531);
nor U14734 (N_14734,N_12113,N_13383);
nand U14735 (N_14735,N_12045,N_12964);
xor U14736 (N_14736,N_12829,N_12563);
nand U14737 (N_14737,N_12068,N_12168);
nand U14738 (N_14738,N_12112,N_12442);
nand U14739 (N_14739,N_13393,N_13296);
xnor U14740 (N_14740,N_13067,N_12228);
xnor U14741 (N_14741,N_13404,N_12664);
nand U14742 (N_14742,N_13445,N_12322);
or U14743 (N_14743,N_12361,N_12183);
or U14744 (N_14744,N_12801,N_13196);
and U14745 (N_14745,N_12445,N_13381);
and U14746 (N_14746,N_12869,N_12395);
nand U14747 (N_14747,N_13386,N_12683);
nand U14748 (N_14748,N_12069,N_13484);
nor U14749 (N_14749,N_12493,N_12194);
nor U14750 (N_14750,N_12812,N_12721);
and U14751 (N_14751,N_12574,N_12413);
nor U14752 (N_14752,N_13241,N_12133);
nor U14753 (N_14753,N_13154,N_13076);
and U14754 (N_14754,N_12323,N_12723);
nor U14755 (N_14755,N_13231,N_13222);
or U14756 (N_14756,N_12638,N_13363);
and U14757 (N_14757,N_12341,N_12711);
and U14758 (N_14758,N_12034,N_13399);
and U14759 (N_14759,N_13444,N_12897);
or U14760 (N_14760,N_13489,N_12044);
nand U14761 (N_14761,N_12526,N_13368);
nor U14762 (N_14762,N_12270,N_12097);
xnor U14763 (N_14763,N_13106,N_13095);
or U14764 (N_14764,N_13319,N_12360);
and U14765 (N_14765,N_13060,N_12297);
nand U14766 (N_14766,N_13364,N_12013);
nand U14767 (N_14767,N_12102,N_13007);
and U14768 (N_14768,N_12385,N_13383);
and U14769 (N_14769,N_12593,N_12812);
and U14770 (N_14770,N_13287,N_12089);
or U14771 (N_14771,N_12022,N_13395);
or U14772 (N_14772,N_12642,N_13326);
xor U14773 (N_14773,N_12672,N_13376);
xor U14774 (N_14774,N_13304,N_12195);
or U14775 (N_14775,N_13498,N_12803);
nand U14776 (N_14776,N_13433,N_12635);
and U14777 (N_14777,N_12131,N_12489);
and U14778 (N_14778,N_13297,N_12635);
and U14779 (N_14779,N_12215,N_12272);
and U14780 (N_14780,N_12925,N_12138);
or U14781 (N_14781,N_12474,N_12951);
nor U14782 (N_14782,N_13244,N_13395);
nand U14783 (N_14783,N_12903,N_12995);
nor U14784 (N_14784,N_12750,N_13288);
or U14785 (N_14785,N_12514,N_13305);
nand U14786 (N_14786,N_12224,N_12232);
nand U14787 (N_14787,N_13250,N_13483);
xnor U14788 (N_14788,N_12459,N_12269);
xnor U14789 (N_14789,N_12139,N_12117);
xor U14790 (N_14790,N_12842,N_12811);
nand U14791 (N_14791,N_13346,N_12840);
nor U14792 (N_14792,N_12369,N_12698);
or U14793 (N_14793,N_12288,N_13086);
nand U14794 (N_14794,N_12683,N_12101);
xor U14795 (N_14795,N_12611,N_12616);
xnor U14796 (N_14796,N_13433,N_12222);
nand U14797 (N_14797,N_12795,N_13167);
nor U14798 (N_14798,N_13267,N_12659);
nand U14799 (N_14799,N_12554,N_12933);
xnor U14800 (N_14800,N_12992,N_13279);
or U14801 (N_14801,N_12954,N_13365);
nand U14802 (N_14802,N_13131,N_12241);
and U14803 (N_14803,N_12217,N_12836);
and U14804 (N_14804,N_12993,N_12312);
or U14805 (N_14805,N_12597,N_13007);
xnor U14806 (N_14806,N_12737,N_13016);
nor U14807 (N_14807,N_12703,N_12937);
and U14808 (N_14808,N_13086,N_12821);
nor U14809 (N_14809,N_13124,N_12252);
and U14810 (N_14810,N_12848,N_12484);
nand U14811 (N_14811,N_13398,N_13289);
or U14812 (N_14812,N_13266,N_13223);
nor U14813 (N_14813,N_13427,N_13164);
xnor U14814 (N_14814,N_13263,N_12856);
nor U14815 (N_14815,N_12208,N_12925);
and U14816 (N_14816,N_12987,N_12189);
xnor U14817 (N_14817,N_13058,N_12350);
nor U14818 (N_14818,N_12321,N_12706);
nor U14819 (N_14819,N_12092,N_12023);
and U14820 (N_14820,N_13329,N_13105);
nor U14821 (N_14821,N_12359,N_13170);
nor U14822 (N_14822,N_12967,N_13141);
or U14823 (N_14823,N_12000,N_12420);
nor U14824 (N_14824,N_12332,N_12127);
xor U14825 (N_14825,N_13096,N_12609);
and U14826 (N_14826,N_12273,N_12144);
xnor U14827 (N_14827,N_12023,N_13391);
or U14828 (N_14828,N_12782,N_12179);
nand U14829 (N_14829,N_12547,N_13184);
or U14830 (N_14830,N_12383,N_12248);
nor U14831 (N_14831,N_12674,N_12982);
and U14832 (N_14832,N_12637,N_12109);
xor U14833 (N_14833,N_12281,N_13281);
nand U14834 (N_14834,N_13413,N_12500);
xnor U14835 (N_14835,N_12198,N_13354);
nor U14836 (N_14836,N_13238,N_12528);
nand U14837 (N_14837,N_12632,N_12362);
nand U14838 (N_14838,N_12566,N_12579);
nand U14839 (N_14839,N_13212,N_12334);
and U14840 (N_14840,N_12693,N_13289);
nand U14841 (N_14841,N_12040,N_13065);
or U14842 (N_14842,N_13435,N_12662);
and U14843 (N_14843,N_12899,N_13179);
nand U14844 (N_14844,N_13410,N_12919);
xnor U14845 (N_14845,N_12383,N_13287);
nand U14846 (N_14846,N_12638,N_12284);
and U14847 (N_14847,N_12724,N_12501);
xor U14848 (N_14848,N_13394,N_12850);
and U14849 (N_14849,N_12832,N_13108);
and U14850 (N_14850,N_12392,N_12563);
nand U14851 (N_14851,N_12738,N_12500);
nor U14852 (N_14852,N_13237,N_12447);
nand U14853 (N_14853,N_13431,N_12858);
xnor U14854 (N_14854,N_12470,N_12614);
nor U14855 (N_14855,N_12779,N_12340);
xnor U14856 (N_14856,N_12211,N_12230);
or U14857 (N_14857,N_12306,N_12460);
nand U14858 (N_14858,N_12435,N_12004);
nor U14859 (N_14859,N_12350,N_12125);
nor U14860 (N_14860,N_12174,N_12805);
and U14861 (N_14861,N_12830,N_12766);
xnor U14862 (N_14862,N_12825,N_13054);
and U14863 (N_14863,N_13320,N_12071);
xnor U14864 (N_14864,N_12602,N_13442);
nor U14865 (N_14865,N_12290,N_13206);
nor U14866 (N_14866,N_13097,N_12183);
nand U14867 (N_14867,N_13248,N_12161);
xnor U14868 (N_14868,N_13398,N_13236);
or U14869 (N_14869,N_12359,N_12613);
nand U14870 (N_14870,N_13470,N_12775);
xor U14871 (N_14871,N_12951,N_12822);
nand U14872 (N_14872,N_12314,N_12418);
nor U14873 (N_14873,N_12925,N_13116);
nor U14874 (N_14874,N_12110,N_13304);
nand U14875 (N_14875,N_12173,N_12756);
xnor U14876 (N_14876,N_12998,N_13427);
nor U14877 (N_14877,N_12418,N_12647);
xor U14878 (N_14878,N_12234,N_12506);
nor U14879 (N_14879,N_12378,N_12397);
nor U14880 (N_14880,N_12956,N_12364);
nand U14881 (N_14881,N_12397,N_12973);
or U14882 (N_14882,N_13455,N_12150);
nor U14883 (N_14883,N_12839,N_12802);
or U14884 (N_14884,N_12466,N_12976);
xnor U14885 (N_14885,N_12559,N_12415);
and U14886 (N_14886,N_12997,N_12543);
or U14887 (N_14887,N_13442,N_12104);
nor U14888 (N_14888,N_12096,N_12370);
nand U14889 (N_14889,N_13199,N_13300);
and U14890 (N_14890,N_13010,N_13021);
xnor U14891 (N_14891,N_12484,N_12931);
or U14892 (N_14892,N_12048,N_12137);
and U14893 (N_14893,N_12385,N_13294);
or U14894 (N_14894,N_12326,N_13187);
xnor U14895 (N_14895,N_12613,N_13398);
xnor U14896 (N_14896,N_12359,N_12824);
nand U14897 (N_14897,N_12272,N_13353);
nand U14898 (N_14898,N_13288,N_12894);
xnor U14899 (N_14899,N_12446,N_13471);
nor U14900 (N_14900,N_12205,N_12403);
xor U14901 (N_14901,N_12570,N_12243);
and U14902 (N_14902,N_12001,N_12101);
and U14903 (N_14903,N_12209,N_12210);
and U14904 (N_14904,N_12082,N_13260);
xor U14905 (N_14905,N_12904,N_12122);
xor U14906 (N_14906,N_12652,N_12310);
nand U14907 (N_14907,N_12666,N_13089);
nand U14908 (N_14908,N_13174,N_13110);
and U14909 (N_14909,N_13154,N_13228);
and U14910 (N_14910,N_12339,N_12059);
xnor U14911 (N_14911,N_12125,N_12113);
nor U14912 (N_14912,N_12701,N_13134);
and U14913 (N_14913,N_13437,N_12958);
nor U14914 (N_14914,N_13026,N_12494);
nand U14915 (N_14915,N_13054,N_12709);
or U14916 (N_14916,N_12582,N_12640);
nand U14917 (N_14917,N_12296,N_12974);
xor U14918 (N_14918,N_12535,N_13174);
nor U14919 (N_14919,N_12073,N_12166);
or U14920 (N_14920,N_12131,N_12135);
or U14921 (N_14921,N_13008,N_12061);
nor U14922 (N_14922,N_12058,N_12574);
or U14923 (N_14923,N_12295,N_12227);
xnor U14924 (N_14924,N_13215,N_13401);
or U14925 (N_14925,N_13092,N_12198);
nand U14926 (N_14926,N_13083,N_13368);
nor U14927 (N_14927,N_13273,N_13263);
nor U14928 (N_14928,N_12176,N_12834);
nor U14929 (N_14929,N_12979,N_13073);
or U14930 (N_14930,N_13490,N_13200);
and U14931 (N_14931,N_12054,N_12826);
nor U14932 (N_14932,N_12992,N_12651);
or U14933 (N_14933,N_12484,N_13417);
and U14934 (N_14934,N_12382,N_13076);
nand U14935 (N_14935,N_12952,N_13123);
and U14936 (N_14936,N_13499,N_12120);
xor U14937 (N_14937,N_13149,N_13407);
or U14938 (N_14938,N_13414,N_12947);
and U14939 (N_14939,N_13385,N_12940);
or U14940 (N_14940,N_12180,N_12986);
xnor U14941 (N_14941,N_13275,N_13418);
or U14942 (N_14942,N_12858,N_12640);
xnor U14943 (N_14943,N_13036,N_12089);
nand U14944 (N_14944,N_13134,N_12522);
nand U14945 (N_14945,N_12706,N_12612);
nor U14946 (N_14946,N_12000,N_12852);
and U14947 (N_14947,N_13221,N_12413);
xor U14948 (N_14948,N_12177,N_12897);
and U14949 (N_14949,N_13003,N_12554);
nand U14950 (N_14950,N_12851,N_12330);
or U14951 (N_14951,N_13310,N_12586);
nor U14952 (N_14952,N_13293,N_12370);
nand U14953 (N_14953,N_13175,N_12761);
nor U14954 (N_14954,N_12417,N_12538);
nand U14955 (N_14955,N_12831,N_13154);
xnor U14956 (N_14956,N_13448,N_13192);
xor U14957 (N_14957,N_13181,N_12655);
nand U14958 (N_14958,N_13378,N_13169);
nor U14959 (N_14959,N_12850,N_12441);
xor U14960 (N_14960,N_12897,N_12011);
nand U14961 (N_14961,N_12653,N_12780);
xnor U14962 (N_14962,N_12243,N_12019);
nand U14963 (N_14963,N_13005,N_12213);
or U14964 (N_14964,N_12010,N_13174);
and U14965 (N_14965,N_12083,N_12841);
nor U14966 (N_14966,N_12379,N_12478);
or U14967 (N_14967,N_13099,N_12079);
nand U14968 (N_14968,N_12243,N_12428);
and U14969 (N_14969,N_13269,N_13260);
nor U14970 (N_14970,N_13437,N_13243);
xnor U14971 (N_14971,N_12370,N_13153);
nor U14972 (N_14972,N_13400,N_12462);
nand U14973 (N_14973,N_12255,N_13277);
and U14974 (N_14974,N_12948,N_12860);
nand U14975 (N_14975,N_12718,N_13191);
nand U14976 (N_14976,N_12671,N_12347);
nand U14977 (N_14977,N_13200,N_12018);
xor U14978 (N_14978,N_12782,N_13291);
xnor U14979 (N_14979,N_13237,N_12269);
xnor U14980 (N_14980,N_13356,N_12373);
nand U14981 (N_14981,N_12868,N_13491);
nor U14982 (N_14982,N_12181,N_13183);
or U14983 (N_14983,N_12484,N_12886);
nor U14984 (N_14984,N_13273,N_13101);
nand U14985 (N_14985,N_12738,N_12940);
xor U14986 (N_14986,N_12595,N_12031);
and U14987 (N_14987,N_12015,N_13325);
nand U14988 (N_14988,N_13342,N_12219);
or U14989 (N_14989,N_12551,N_12537);
or U14990 (N_14990,N_12192,N_13364);
or U14991 (N_14991,N_12685,N_13283);
xor U14992 (N_14992,N_12293,N_12861);
nor U14993 (N_14993,N_12120,N_12338);
xnor U14994 (N_14994,N_13370,N_12285);
and U14995 (N_14995,N_12199,N_12453);
xor U14996 (N_14996,N_12456,N_12063);
nor U14997 (N_14997,N_12895,N_12509);
xnor U14998 (N_14998,N_12875,N_13364);
and U14999 (N_14999,N_12332,N_12107);
nand UO_0 (O_0,N_13698,N_14380);
and UO_1 (O_1,N_13814,N_13829);
and UO_2 (O_2,N_14469,N_14580);
nand UO_3 (O_3,N_14165,N_13892);
or UO_4 (O_4,N_13570,N_13601);
xor UO_5 (O_5,N_14574,N_13554);
and UO_6 (O_6,N_13887,N_14014);
or UO_7 (O_7,N_14339,N_13864);
xnor UO_8 (O_8,N_13974,N_14067);
nand UO_9 (O_9,N_14579,N_14711);
nand UO_10 (O_10,N_14447,N_14297);
nor UO_11 (O_11,N_14115,N_14201);
nand UO_12 (O_12,N_13672,N_13705);
nand UO_13 (O_13,N_13637,N_14345);
or UO_14 (O_14,N_14076,N_14240);
or UO_15 (O_15,N_14806,N_14865);
xor UO_16 (O_16,N_14528,N_14203);
or UO_17 (O_17,N_13866,N_14448);
nor UO_18 (O_18,N_14163,N_14891);
nor UO_19 (O_19,N_13583,N_14931);
nor UO_20 (O_20,N_14667,N_14735);
nor UO_21 (O_21,N_13796,N_14134);
nor UO_22 (O_22,N_14591,N_14706);
nor UO_23 (O_23,N_14133,N_14625);
and UO_24 (O_24,N_13692,N_14744);
nor UO_25 (O_25,N_14436,N_14830);
and UO_26 (O_26,N_14600,N_13549);
xor UO_27 (O_27,N_14928,N_14455);
and UO_28 (O_28,N_13807,N_14614);
nor UO_29 (O_29,N_14334,N_13643);
nor UO_30 (O_30,N_13815,N_14142);
or UO_31 (O_31,N_14803,N_14034);
nand UO_32 (O_32,N_14598,N_13857);
or UO_33 (O_33,N_14585,N_14100);
nor UO_34 (O_34,N_14826,N_14964);
or UO_35 (O_35,N_14534,N_13560);
xnor UO_36 (O_36,N_14210,N_13627);
xnor UO_37 (O_37,N_13721,N_14452);
xnor UO_38 (O_38,N_14799,N_14660);
xor UO_39 (O_39,N_13582,N_14227);
and UO_40 (O_40,N_14286,N_13526);
or UO_41 (O_41,N_13641,N_14899);
nor UO_42 (O_42,N_14065,N_13562);
nor UO_43 (O_43,N_13738,N_14661);
and UO_44 (O_44,N_14418,N_13747);
or UO_45 (O_45,N_14129,N_13851);
and UO_46 (O_46,N_14800,N_13666);
and UO_47 (O_47,N_13517,N_13848);
nand UO_48 (O_48,N_14536,N_13586);
nand UO_49 (O_49,N_14130,N_13856);
nor UO_50 (O_50,N_14486,N_14841);
nor UO_51 (O_51,N_13633,N_14679);
or UO_52 (O_52,N_14973,N_14649);
or UO_53 (O_53,N_13736,N_14620);
and UO_54 (O_54,N_14463,N_14650);
or UO_55 (O_55,N_13676,N_13605);
nand UO_56 (O_56,N_14836,N_13520);
nor UO_57 (O_57,N_14155,N_14874);
nand UO_58 (O_58,N_13654,N_13952);
xor UO_59 (O_59,N_13537,N_14063);
xor UO_60 (O_60,N_14814,N_14499);
nor UO_61 (O_61,N_14689,N_14219);
or UO_62 (O_62,N_13776,N_14125);
xnor UO_63 (O_63,N_13630,N_14853);
nand UO_64 (O_64,N_14244,N_14717);
nand UO_65 (O_65,N_14838,N_14762);
nor UO_66 (O_66,N_14484,N_14358);
nor UO_67 (O_67,N_13836,N_14843);
nor UO_68 (O_68,N_14618,N_14208);
nor UO_69 (O_69,N_13806,N_14186);
nor UO_70 (O_70,N_14225,N_14916);
and UO_71 (O_71,N_13896,N_14350);
xor UO_72 (O_72,N_13906,N_13763);
xnor UO_73 (O_73,N_14429,N_14777);
and UO_74 (O_74,N_14688,N_14426);
nand UO_75 (O_75,N_13865,N_13659);
or UO_76 (O_76,N_13548,N_14007);
or UO_77 (O_77,N_14589,N_13700);
or UO_78 (O_78,N_14521,N_13876);
or UO_79 (O_79,N_14386,N_14875);
or UO_80 (O_80,N_14375,N_14260);
xnor UO_81 (O_81,N_14236,N_14287);
xnor UO_82 (O_82,N_13935,N_14882);
nor UO_83 (O_83,N_13505,N_14432);
or UO_84 (O_84,N_14757,N_14329);
and UO_85 (O_85,N_14941,N_13936);
or UO_86 (O_86,N_13832,N_14220);
xor UO_87 (O_87,N_13702,N_13731);
and UO_88 (O_88,N_13536,N_13804);
or UO_89 (O_89,N_14046,N_14718);
and UO_90 (O_90,N_14617,N_13579);
xnor UO_91 (O_91,N_14795,N_14975);
and UO_92 (O_92,N_14283,N_14682);
and UO_93 (O_93,N_14226,N_14316);
and UO_94 (O_94,N_14561,N_13991);
nand UO_95 (O_95,N_14075,N_14867);
nor UO_96 (O_96,N_14372,N_13810);
nand UO_97 (O_97,N_14274,N_13675);
nand UO_98 (O_98,N_14554,N_14467);
nand UO_99 (O_99,N_14745,N_13594);
nor UO_100 (O_100,N_13874,N_13539);
nand UO_101 (O_101,N_14529,N_14383);
and UO_102 (O_102,N_14560,N_14877);
and UO_103 (O_103,N_13772,N_14263);
xnor UO_104 (O_104,N_14581,N_13743);
nor UO_105 (O_105,N_13577,N_13996);
and UO_106 (O_106,N_14824,N_14179);
nand UO_107 (O_107,N_14629,N_14030);
xnor UO_108 (O_108,N_13571,N_14572);
xnor UO_109 (O_109,N_14387,N_13541);
xor UO_110 (O_110,N_14000,N_13744);
nor UO_111 (O_111,N_13985,N_14754);
nand UO_112 (O_112,N_14045,N_13972);
nor UO_113 (O_113,N_14002,N_14073);
and UO_114 (O_114,N_14296,N_13703);
nand UO_115 (O_115,N_14478,N_14623);
nor UO_116 (O_116,N_13746,N_14793);
or UO_117 (O_117,N_14051,N_14072);
xor UO_118 (O_118,N_14936,N_14999);
nand UO_119 (O_119,N_14475,N_13715);
xor UO_120 (O_120,N_13839,N_14972);
xor UO_121 (O_121,N_14898,N_14815);
xor UO_122 (O_122,N_14098,N_14729);
xor UO_123 (O_123,N_14465,N_14720);
xor UO_124 (O_124,N_14050,N_14828);
nand UO_125 (O_125,N_13793,N_14987);
and UO_126 (O_126,N_14769,N_13532);
or UO_127 (O_127,N_14171,N_14214);
nand UO_128 (O_128,N_14593,N_13689);
nand UO_129 (O_129,N_14594,N_14366);
xnor UO_130 (O_130,N_13800,N_13679);
and UO_131 (O_131,N_14449,N_14077);
nor UO_132 (O_132,N_14110,N_14330);
and UO_133 (O_133,N_14866,N_14848);
and UO_134 (O_134,N_14004,N_13784);
or UO_135 (O_135,N_13949,N_13830);
and UO_136 (O_136,N_13841,N_14578);
xor UO_137 (O_137,N_14342,N_14481);
or UO_138 (O_138,N_14279,N_14114);
or UO_139 (O_139,N_14253,N_13955);
or UO_140 (O_140,N_14121,N_14553);
and UO_141 (O_141,N_14859,N_14218);
and UO_142 (O_142,N_14736,N_14373);
nor UO_143 (O_143,N_13727,N_13948);
nand UO_144 (O_144,N_14801,N_14099);
or UO_145 (O_145,N_14568,N_14992);
or UO_146 (O_146,N_13982,N_14362);
nand UO_147 (O_147,N_14507,N_14792);
nor UO_148 (O_148,N_14854,N_14923);
xnor UO_149 (O_149,N_13669,N_14710);
nand UO_150 (O_150,N_13947,N_14335);
and UO_151 (O_151,N_14023,N_13895);
xor UO_152 (O_152,N_13998,N_13501);
and UO_153 (O_153,N_13651,N_14080);
xnor UO_154 (O_154,N_13535,N_14681);
and UO_155 (O_155,N_14333,N_14108);
nand UO_156 (O_156,N_14331,N_13681);
nand UO_157 (O_157,N_14611,N_14892);
and UO_158 (O_158,N_14963,N_13889);
nand UO_159 (O_159,N_14543,N_14889);
xor UO_160 (O_160,N_14040,N_14157);
nand UO_161 (O_161,N_14758,N_14621);
nand UO_162 (O_162,N_14054,N_14038);
nand UO_163 (O_163,N_13894,N_14317);
xnor UO_164 (O_164,N_13886,N_14785);
nor UO_165 (O_165,N_13922,N_13656);
xnor UO_166 (O_166,N_14596,N_13735);
nor UO_167 (O_167,N_13683,N_14135);
nand UO_168 (O_168,N_14950,N_13811);
or UO_169 (O_169,N_13591,N_14784);
nand UO_170 (O_170,N_13785,N_14370);
and UO_171 (O_171,N_13777,N_13901);
nand UO_172 (O_172,N_14247,N_13623);
or UO_173 (O_173,N_13649,N_13657);
nand UO_174 (O_174,N_14187,N_13572);
nand UO_175 (O_175,N_13515,N_14140);
nand UO_176 (O_176,N_14281,N_14737);
nand UO_177 (O_177,N_13607,N_13580);
or UO_178 (O_178,N_14196,N_13644);
and UO_179 (O_179,N_14860,N_14085);
nor UO_180 (O_180,N_14492,N_14403);
nand UO_181 (O_181,N_14061,N_13919);
and UO_182 (O_182,N_14913,N_13559);
xor UO_183 (O_183,N_14783,N_14172);
nand UO_184 (O_184,N_14986,N_14044);
nor UO_185 (O_185,N_13879,N_13965);
nor UO_186 (O_186,N_14779,N_14609);
or UO_187 (O_187,N_14068,N_14359);
and UO_188 (O_188,N_14693,N_14789);
nor UO_189 (O_189,N_13592,N_14907);
and UO_190 (O_190,N_14107,N_14053);
or UO_191 (O_191,N_13826,N_14739);
or UO_192 (O_192,N_13913,N_14103);
xnor UO_193 (O_193,N_13691,N_13693);
xor UO_194 (O_194,N_14645,N_14940);
or UO_195 (O_195,N_14074,N_14340);
nand UO_196 (O_196,N_14636,N_14816);
and UO_197 (O_197,N_14648,N_14303);
xor UO_198 (O_198,N_13749,N_13805);
and UO_199 (O_199,N_14658,N_13714);
or UO_200 (O_200,N_13771,N_14791);
or UO_201 (O_201,N_13640,N_14532);
nor UO_202 (O_202,N_14419,N_14926);
nor UO_203 (O_203,N_14835,N_14774);
nand UO_204 (O_204,N_14357,N_14035);
nor UO_205 (O_205,N_14879,N_14632);
or UO_206 (O_206,N_14722,N_14150);
xor UO_207 (O_207,N_14153,N_14293);
xor UO_208 (O_208,N_13604,N_14746);
xnor UO_209 (O_209,N_13635,N_13665);
xnor UO_210 (O_210,N_14016,N_13927);
nand UO_211 (O_211,N_13525,N_13709);
nor UO_212 (O_212,N_14673,N_13696);
nor UO_213 (O_213,N_14610,N_13512);
and UO_214 (O_214,N_14542,N_14396);
xnor UO_215 (O_215,N_14470,N_13500);
nor UO_216 (O_216,N_14540,N_14850);
nor UO_217 (O_217,N_14057,N_14683);
nor UO_218 (O_218,N_13625,N_14275);
and UO_219 (O_219,N_14969,N_13650);
nand UO_220 (O_220,N_14787,N_13843);
xnor UO_221 (O_221,N_14217,N_14491);
nand UO_222 (O_222,N_13611,N_14863);
nor UO_223 (O_223,N_14434,N_14912);
and UO_224 (O_224,N_13544,N_14302);
or UO_225 (O_225,N_14984,N_14195);
nor UO_226 (O_226,N_14438,N_13711);
and UO_227 (O_227,N_13523,N_14713);
nand UO_228 (O_228,N_13853,N_14490);
or UO_229 (O_229,N_14404,N_14437);
xnor UO_230 (O_230,N_14606,N_13567);
xor UO_231 (O_231,N_14310,N_14919);
nor UO_232 (O_232,N_13509,N_13957);
nor UO_233 (O_233,N_13897,N_14117);
and UO_234 (O_234,N_13827,N_14991);
xnor UO_235 (O_235,N_14237,N_14116);
or UO_236 (O_236,N_14932,N_13566);
or UO_237 (O_237,N_14805,N_14476);
or UO_238 (O_238,N_13860,N_14304);
or UO_239 (O_239,N_14748,N_14104);
nand UO_240 (O_240,N_14687,N_14551);
nand UO_241 (O_241,N_14678,N_14101);
nor UO_242 (O_242,N_13992,N_14336);
nor UO_243 (O_243,N_14152,N_13802);
nand UO_244 (O_244,N_14262,N_13950);
and UO_245 (O_245,N_14890,N_13699);
nor UO_246 (O_246,N_14485,N_14137);
nand UO_247 (O_247,N_14430,N_14385);
xnor UO_248 (O_248,N_14307,N_13729);
nor UO_249 (O_249,N_13930,N_14974);
xor UO_250 (O_250,N_14708,N_13734);
or UO_251 (O_251,N_14457,N_14368);
nand UO_252 (O_252,N_13921,N_14680);
nand UO_253 (O_253,N_14313,N_14977);
nor UO_254 (O_254,N_13733,N_14665);
or UO_255 (O_255,N_13759,N_14181);
or UO_256 (O_256,N_14136,N_14138);
xor UO_257 (O_257,N_14164,N_14894);
or UO_258 (O_258,N_13503,N_14381);
xor UO_259 (O_259,N_13756,N_14451);
nor UO_260 (O_260,N_14628,N_14184);
nand UO_261 (O_261,N_14753,N_13621);
and UO_262 (O_262,N_14078,N_14031);
or UO_263 (O_263,N_14692,N_13531);
or UO_264 (O_264,N_14059,N_14527);
and UO_265 (O_265,N_14128,N_14505);
or UO_266 (O_266,N_13911,N_14906);
or UO_267 (O_267,N_14238,N_14514);
nand UO_268 (O_268,N_14288,N_13979);
nor UO_269 (O_269,N_13717,N_14592);
nand UO_270 (O_270,N_14763,N_14962);
nand UO_271 (O_271,N_14233,N_13719);
xnor UO_272 (O_272,N_13694,N_14024);
and UO_273 (O_273,N_14361,N_13540);
nor UO_274 (O_274,N_14020,N_13534);
nand UO_275 (O_275,N_13612,N_14167);
or UO_276 (O_276,N_14901,N_14555);
or UO_277 (O_277,N_13620,N_13929);
nand UO_278 (O_278,N_14111,N_14160);
or UO_279 (O_279,N_14563,N_14959);
and UO_280 (O_280,N_13993,N_13510);
nand UO_281 (O_281,N_13902,N_14669);
xor UO_282 (O_282,N_13631,N_14670);
or UO_283 (O_283,N_13511,N_14444);
nor UO_284 (O_284,N_14539,N_14526);
nand UO_285 (O_285,N_13903,N_14011);
xor UO_286 (O_286,N_14338,N_14326);
nor UO_287 (O_287,N_14041,N_14935);
or UO_288 (O_288,N_14768,N_14633);
xor UO_289 (O_289,N_14407,N_14740);
and UO_290 (O_290,N_14946,N_14119);
xor UO_291 (O_291,N_14885,N_13602);
xor UO_292 (O_292,N_14272,N_14096);
xor UO_293 (O_293,N_14849,N_14559);
xnor UO_294 (O_294,N_13909,N_14276);
and UO_295 (O_295,N_14668,N_13755);
and UO_296 (O_296,N_14637,N_13575);
nor UO_297 (O_297,N_14249,N_14215);
xor UO_298 (O_298,N_14696,N_14066);
nor UO_299 (O_299,N_14425,N_13639);
nor UO_300 (O_300,N_13712,N_14869);
and UO_301 (O_301,N_14684,N_14749);
or UO_302 (O_302,N_14643,N_13870);
xor UO_303 (O_303,N_13761,N_14765);
and UO_304 (O_304,N_13568,N_13661);
nand UO_305 (O_305,N_14771,N_13923);
xor UO_306 (O_306,N_14832,N_14821);
xnor UO_307 (O_307,N_13783,N_14520);
nor UO_308 (O_308,N_14945,N_14388);
or UO_309 (O_309,N_14151,N_14017);
nand UO_310 (O_310,N_14966,N_13975);
nand UO_311 (O_311,N_13619,N_13924);
or UO_312 (O_312,N_13545,N_14691);
nand UO_313 (O_313,N_13859,N_14466);
xnor UO_314 (O_314,N_13742,N_14515);
nand UO_315 (O_315,N_13688,N_14410);
nor UO_316 (O_316,N_14881,N_13646);
and UO_317 (O_317,N_14599,N_13518);
and UO_318 (O_318,N_13762,N_13662);
nand UO_319 (O_319,N_14012,N_13524);
or UO_320 (O_320,N_13697,N_13752);
or UO_321 (O_321,N_14095,N_14988);
or UO_322 (O_322,N_14391,N_14558);
nor UO_323 (O_323,N_13613,N_13645);
nand UO_324 (O_324,N_14369,N_14106);
or UO_325 (O_325,N_14209,N_14423);
nand UO_326 (O_326,N_14174,N_14062);
or UO_327 (O_327,N_14378,N_14995);
or UO_328 (O_328,N_13881,N_14587);
nand UO_329 (O_329,N_13615,N_13838);
xnor UO_330 (O_330,N_14207,N_13969);
nand UO_331 (O_331,N_14944,N_13674);
nor UO_332 (O_332,N_14318,N_13953);
or UO_333 (O_333,N_14725,N_14773);
nand UO_334 (O_334,N_14188,N_14595);
nor UO_335 (O_335,N_14639,N_14290);
xor UO_336 (O_336,N_14797,N_14379);
nand UO_337 (O_337,N_14270,N_14531);
nand UO_338 (O_338,N_14462,N_13724);
xnor UO_339 (O_339,N_14042,N_13816);
xor UO_340 (O_340,N_13614,N_13822);
nor UO_341 (O_341,N_14474,N_13946);
and UO_342 (O_342,N_14615,N_14958);
nand UO_343 (O_343,N_13622,N_14189);
xnor UO_344 (O_344,N_14728,N_14489);
xnor UO_345 (O_345,N_14093,N_14346);
or UO_346 (O_346,N_14003,N_13642);
nor UO_347 (O_347,N_13732,N_14231);
xor UO_348 (O_348,N_14126,N_14788);
and UO_349 (O_349,N_14158,N_14390);
nor UO_350 (O_350,N_14605,N_14212);
nor UO_351 (O_351,N_13934,N_14228);
xnor UO_352 (O_352,N_14056,N_14384);
and UO_353 (O_353,N_13823,N_14493);
or UO_354 (O_354,N_13561,N_14433);
nand UO_355 (O_355,N_13847,N_14084);
xnor UO_356 (O_356,N_13671,N_14471);
xor UO_357 (O_357,N_13799,N_14659);
xnor UO_358 (O_358,N_14353,N_14770);
nor UO_359 (O_359,N_14674,N_14312);
and UO_360 (O_360,N_13942,N_14925);
nor UO_361 (O_361,N_14976,N_13907);
nor UO_362 (O_362,N_13720,N_14967);
or UO_363 (O_363,N_14970,N_14397);
xor UO_364 (O_364,N_14817,N_14804);
nor UO_365 (O_365,N_14915,N_14535);
xor UO_366 (O_366,N_14392,N_14845);
nor UO_367 (O_367,N_14701,N_13716);
nor UO_368 (O_368,N_13920,N_13775);
xor UO_369 (O_369,N_14435,N_13758);
nand UO_370 (O_370,N_14036,N_14834);
and UO_371 (O_371,N_14147,N_14734);
nand UO_372 (O_372,N_14624,N_13900);
nand UO_373 (O_373,N_14344,N_13835);
and UO_374 (O_374,N_13600,N_13877);
xnor UO_375 (O_375,N_14025,N_13854);
nand UO_376 (O_376,N_14494,N_13730);
xnor UO_377 (O_377,N_14979,N_14778);
and UO_378 (O_378,N_14355,N_14176);
and UO_379 (O_379,N_13837,N_13686);
nand UO_380 (O_380,N_13739,N_14756);
and UO_381 (O_381,N_14052,N_14464);
nand UO_382 (O_382,N_14809,N_13967);
xnor UO_383 (O_383,N_13628,N_14571);
xnor UO_384 (O_384,N_14306,N_14268);
or UO_385 (O_385,N_14064,N_13863);
nor UO_386 (O_386,N_13677,N_14569);
nand UO_387 (O_387,N_13753,N_14252);
and UO_388 (O_388,N_14168,N_13995);
xor UO_389 (O_389,N_14477,N_14092);
nand UO_390 (O_390,N_14978,N_14401);
nand UO_391 (O_391,N_13812,N_13825);
nand UO_392 (O_392,N_13905,N_13610);
nand UO_393 (O_393,N_13981,N_14256);
nand UO_394 (O_394,N_14439,N_14193);
and UO_395 (O_395,N_14980,N_14199);
xor UO_396 (O_396,N_14254,N_13648);
nor UO_397 (O_397,N_14652,N_13754);
nand UO_398 (O_398,N_14402,N_14232);
or UO_399 (O_399,N_14173,N_14332);
or UO_400 (O_400,N_14417,N_14582);
or UO_401 (O_401,N_14127,N_14170);
nor UO_402 (O_402,N_13558,N_13585);
or UO_403 (O_403,N_14182,N_13740);
or UO_404 (O_404,N_13831,N_14314);
xnor UO_405 (O_405,N_13587,N_14008);
nand UO_406 (O_406,N_14604,N_14896);
nand UO_407 (O_407,N_13868,N_14458);
or UO_408 (O_408,N_13668,N_14700);
or UO_409 (O_409,N_14741,N_13867);
xnor UO_410 (O_410,N_14685,N_14951);
xor UO_411 (O_411,N_14200,N_14445);
and UO_412 (O_412,N_13533,N_14886);
or UO_413 (O_413,N_14523,N_13928);
xor UO_414 (O_414,N_13757,N_13767);
and UO_415 (O_415,N_14183,N_14010);
xor UO_416 (O_416,N_13550,N_14938);
and UO_417 (O_417,N_14141,N_13728);
nor UO_418 (O_418,N_13556,N_13774);
nor UO_419 (O_419,N_14686,N_13552);
and UO_420 (O_420,N_14006,N_13855);
and UO_421 (O_421,N_13765,N_14122);
and UO_422 (O_422,N_13680,N_14185);
nor UO_423 (O_423,N_13846,N_14197);
nor UO_424 (O_424,N_14862,N_14724);
and UO_425 (O_425,N_13987,N_13940);
nor UO_426 (O_426,N_13655,N_13820);
and UO_427 (O_427,N_14933,N_14942);
nor UO_428 (O_428,N_13880,N_14698);
nand UO_429 (O_429,N_13597,N_13933);
xor UO_430 (O_430,N_13595,N_14562);
nor UO_431 (O_431,N_14246,N_13722);
or UO_432 (O_432,N_14619,N_13663);
and UO_433 (O_433,N_14440,N_13875);
nor UO_434 (O_434,N_14833,N_13673);
xor UO_435 (O_435,N_13917,N_14413);
or UO_436 (O_436,N_13926,N_13617);
or UO_437 (O_437,N_14144,N_14608);
and UO_438 (O_438,N_14510,N_13899);
nand UO_439 (O_439,N_14731,N_13773);
and UO_440 (O_440,N_14230,N_14666);
nor UO_441 (O_441,N_13660,N_13817);
nor UO_442 (O_442,N_13707,N_14261);
and UO_443 (O_443,N_13710,N_14905);
or UO_444 (O_444,N_13861,N_14767);
xnor UO_445 (O_445,N_13989,N_13690);
or UO_446 (O_446,N_14612,N_13576);
nand UO_447 (O_447,N_13821,N_14794);
xnor UO_448 (O_448,N_14638,N_13939);
and UO_449 (O_449,N_14613,N_13593);
nor UO_450 (O_450,N_14903,N_14377);
nor UO_451 (O_451,N_13977,N_14202);
or UO_452 (O_452,N_14504,N_14308);
xor UO_453 (O_453,N_14271,N_14205);
or UO_454 (O_454,N_14395,N_14884);
nand UO_455 (O_455,N_14947,N_14411);
and UO_456 (O_456,N_14294,N_14154);
or UO_457 (O_457,N_13961,N_14132);
nor UO_458 (O_458,N_13932,N_14319);
or UO_459 (O_459,N_14421,N_13898);
and UO_460 (O_460,N_13547,N_14577);
xor UO_461 (O_461,N_13893,N_13522);
nand UO_462 (O_462,N_14782,N_14583);
and UO_463 (O_463,N_14323,N_14211);
and UO_464 (O_464,N_14878,N_14516);
xor UO_465 (O_465,N_14204,N_14295);
nor UO_466 (O_466,N_13647,N_14408);
or UO_467 (O_467,N_14086,N_13589);
and UO_468 (O_468,N_14921,N_14997);
and UO_469 (O_469,N_13748,N_14723);
xor UO_470 (O_470,N_14761,N_13883);
nand UO_471 (O_471,N_14989,N_14161);
or UO_472 (O_472,N_13653,N_13751);
xor UO_473 (O_473,N_14868,N_13956);
or UO_474 (O_474,N_13988,N_13912);
nor UO_475 (O_475,N_14699,N_13787);
and UO_476 (O_476,N_13596,N_13609);
nand UO_477 (O_477,N_13781,N_13543);
and UO_478 (O_478,N_13513,N_13701);
xnor UO_479 (O_479,N_14888,N_13789);
nor UO_480 (O_480,N_14055,N_13599);
nor UO_481 (O_481,N_13782,N_14811);
nor UO_482 (O_482,N_13845,N_14641);
nand UO_483 (O_483,N_14269,N_13869);
and UO_484 (O_484,N_13632,N_14714);
xnor UO_485 (O_485,N_14409,N_14088);
nand UO_486 (O_486,N_14503,N_14647);
and UO_487 (O_487,N_14677,N_13573);
xnor UO_488 (O_488,N_13658,N_14533);
nand UO_489 (O_489,N_14149,N_14416);
xnor UO_490 (O_490,N_14983,N_13584);
xor UO_491 (O_491,N_14043,N_14917);
nor UO_492 (O_492,N_14028,N_14022);
nor UO_493 (O_493,N_13968,N_14541);
nor UO_494 (O_494,N_14565,N_14083);
or UO_495 (O_495,N_13685,N_14364);
nand UO_496 (O_496,N_14655,N_13801);
and UO_497 (O_497,N_13983,N_14180);
and UO_498 (O_498,N_14376,N_14742);
or UO_499 (O_499,N_14810,N_14575);
xor UO_500 (O_500,N_14703,N_14190);
xnor UO_501 (O_501,N_14786,N_13999);
or UO_502 (O_502,N_14690,N_14780);
or UO_503 (O_503,N_14248,N_13652);
or UO_504 (O_504,N_14968,N_14732);
and UO_505 (O_505,N_14143,N_14552);
nand UO_506 (O_506,N_14846,N_14823);
nor UO_507 (O_507,N_13706,N_14813);
nand UO_508 (O_508,N_14299,N_14192);
or UO_509 (O_509,N_14234,N_14965);
or UO_510 (O_510,N_14148,N_14831);
and UO_511 (O_511,N_14672,N_14118);
and UO_512 (O_512,N_14341,N_13840);
nor UO_513 (O_513,N_14264,N_14229);
xor UO_514 (O_514,N_14420,N_13794);
nor UO_515 (O_515,N_14405,N_13629);
nor UO_516 (O_516,N_14663,N_14861);
and UO_517 (O_517,N_13986,N_13862);
or UO_518 (O_518,N_14829,N_14631);
and UO_519 (O_519,N_14827,N_13590);
or UO_520 (O_520,N_13764,N_14524);
nor UO_521 (O_521,N_14626,N_13971);
or UO_522 (O_522,N_14070,N_13973);
xor UO_523 (O_523,N_14267,N_14960);
or UO_524 (O_524,N_13873,N_14911);
nand UO_525 (O_525,N_14343,N_13916);
and UO_526 (O_526,N_13626,N_13606);
and UO_527 (O_527,N_14442,N_13670);
and UO_528 (O_528,N_14424,N_13780);
and UO_529 (O_529,N_14443,N_13557);
or UO_530 (O_530,N_14738,N_14955);
nor UO_531 (O_531,N_14544,N_14566);
xnor UO_532 (O_532,N_14537,N_14300);
nor UO_533 (O_533,N_14081,N_14258);
nor UO_534 (O_534,N_14897,N_14996);
nor UO_535 (O_535,N_13521,N_14627);
xnor UO_536 (O_536,N_14454,N_14428);
nand UO_537 (O_537,N_14949,N_14904);
and UO_538 (O_538,N_13964,N_14880);
xnor UO_539 (O_539,N_14759,N_13528);
nand UO_540 (O_540,N_14990,N_13616);
nor UO_541 (O_541,N_14519,N_14656);
nor UO_542 (O_542,N_14727,N_14671);
or UO_543 (O_543,N_13833,N_13850);
xnor UO_544 (O_544,N_14398,N_14037);
and UO_545 (O_545,N_14048,N_14576);
nand UO_546 (O_546,N_13667,N_13786);
nor UO_547 (O_547,N_14082,N_14363);
and UO_548 (O_548,N_14914,N_14764);
nand UO_549 (O_549,N_14642,N_14277);
or UO_550 (O_550,N_14517,N_13608);
or UO_551 (O_551,N_14726,N_14131);
nor UO_552 (O_552,N_14802,N_14909);
nand UO_553 (O_553,N_14545,N_14298);
nor UO_554 (O_554,N_13852,N_14751);
or UO_555 (O_555,N_14029,N_14586);
nor UO_556 (O_556,N_14772,N_13664);
or UO_557 (O_557,N_13943,N_14971);
and UO_558 (O_558,N_14399,N_14001);
and UO_559 (O_559,N_13984,N_14382);
nor UO_560 (O_560,N_14501,N_13925);
or UO_561 (O_561,N_14400,N_14223);
nand UO_562 (O_562,N_14159,N_14590);
and UO_563 (O_563,N_13564,N_14844);
or UO_564 (O_564,N_14374,N_13792);
nor UO_565 (O_565,N_14864,N_14169);
or UO_566 (O_566,N_14498,N_14351);
xnor UO_567 (O_567,N_14743,N_14887);
and UO_568 (O_568,N_14090,N_14356);
or UO_569 (O_569,N_13872,N_14512);
nand UO_570 (O_570,N_13791,N_14630);
nor UO_571 (O_571,N_13624,N_13885);
nand UO_572 (O_572,N_14216,N_14895);
and UO_573 (O_573,N_14352,N_13638);
nand UO_574 (O_574,N_14654,N_14089);
or UO_575 (O_575,N_13910,N_14360);
or UO_576 (O_576,N_13904,N_14750);
and UO_577 (O_577,N_13636,N_14285);
and UO_578 (O_578,N_14145,N_14124);
or UO_579 (O_579,N_14239,N_14243);
nor UO_580 (O_580,N_14930,N_13976);
or UO_581 (O_581,N_14640,N_14259);
nor UO_582 (O_582,N_13790,N_14354);
or UO_583 (O_583,N_14453,N_14939);
and UO_584 (O_584,N_14305,N_14224);
nand UO_585 (O_585,N_14123,N_14311);
xnor UO_586 (O_586,N_13813,N_13918);
nand UO_587 (O_587,N_14922,N_14837);
and UO_588 (O_588,N_13871,N_13938);
and UO_589 (O_589,N_14422,N_13529);
or UO_590 (O_590,N_13527,N_14328);
xnor UO_591 (O_591,N_14109,N_14394);
nand UO_592 (O_592,N_14675,N_13718);
and UO_593 (O_593,N_14557,N_14695);
nor UO_594 (O_594,N_13788,N_14245);
xor UO_595 (O_595,N_14456,N_14255);
nor UO_596 (O_596,N_14005,N_14807);
and UO_597 (O_597,N_14320,N_14495);
xnor UO_598 (O_598,N_14026,N_14957);
or UO_599 (O_599,N_14257,N_14146);
nor UO_600 (O_600,N_13737,N_14156);
or UO_601 (O_601,N_13941,N_14796);
or UO_602 (O_602,N_14511,N_14918);
and UO_603 (O_603,N_14694,N_14483);
and UO_604 (O_604,N_13588,N_14924);
and UO_605 (O_605,N_13516,N_13844);
nor UO_606 (O_606,N_14564,N_13507);
nand UO_607 (O_607,N_14525,N_14616);
or UO_608 (O_608,N_14284,N_14715);
nor UO_609 (O_609,N_13704,N_14752);
xnor UO_610 (O_610,N_14733,N_14112);
nor UO_611 (O_611,N_13891,N_13908);
and UO_612 (O_612,N_14927,N_14981);
and UO_613 (O_613,N_14712,N_14550);
nor UO_614 (O_614,N_14349,N_13687);
and UO_615 (O_615,N_14488,N_13884);
nor UO_616 (O_616,N_14337,N_14446);
nor UO_617 (O_617,N_14513,N_14191);
xor UO_618 (O_618,N_13682,N_14097);
or UO_619 (O_619,N_13770,N_14325);
xor UO_620 (O_620,N_13723,N_14993);
xor UO_621 (O_621,N_14943,N_14876);
xnor UO_622 (O_622,N_13779,N_13769);
nand UO_623 (O_623,N_13824,N_14952);
nor UO_624 (O_624,N_14820,N_14166);
nand UO_625 (O_625,N_14530,N_14635);
nand UO_626 (O_626,N_14570,N_14327);
or UO_627 (O_627,N_13504,N_14177);
and UO_628 (O_628,N_14178,N_14058);
and UO_629 (O_629,N_14021,N_14087);
nor UO_630 (O_630,N_13538,N_13768);
xnor UO_631 (O_631,N_13809,N_14509);
nor UO_632 (O_632,N_14646,N_13551);
nor UO_633 (O_633,N_14573,N_14548);
nor UO_634 (O_634,N_13798,N_14321);
xor UO_635 (O_635,N_14644,N_14468);
or UO_636 (O_636,N_13506,N_14603);
or UO_637 (O_637,N_14790,N_14954);
xor UO_638 (O_638,N_14102,N_14755);
and UO_639 (O_639,N_14760,N_13542);
or UO_640 (O_640,N_14709,N_14047);
and UO_641 (O_641,N_13819,N_14393);
or UO_642 (O_642,N_14664,N_13708);
or UO_643 (O_643,N_14389,N_13890);
xor UO_644 (O_644,N_14910,N_13980);
nor UO_645 (O_645,N_13958,N_14412);
and UO_646 (O_646,N_13514,N_13978);
xor UO_647 (O_647,N_14033,N_14985);
nand UO_648 (O_648,N_14009,N_14702);
nand UO_649 (O_649,N_14348,N_14441);
or UO_650 (O_650,N_14460,N_14496);
nand UO_651 (O_651,N_14929,N_13882);
and UO_652 (O_652,N_14347,N_13828);
and UO_653 (O_653,N_14459,N_13678);
and UO_654 (O_654,N_14819,N_14676);
nor UO_655 (O_655,N_13963,N_14602);
xnor UO_656 (O_656,N_13954,N_13578);
or UO_657 (O_657,N_14856,N_14497);
xnor UO_658 (O_658,N_14105,N_14538);
xnor UO_659 (O_659,N_13618,N_14235);
xnor UO_660 (O_660,N_14839,N_13603);
nand UO_661 (O_661,N_14473,N_13915);
and UO_662 (O_662,N_13842,N_14273);
xnor UO_663 (O_663,N_14301,N_14776);
or UO_664 (O_664,N_14719,N_14588);
xnor UO_665 (O_665,N_13750,N_14781);
xor UO_666 (O_666,N_14908,N_14071);
nand UO_667 (O_667,N_14406,N_14704);
and UO_668 (O_668,N_13745,N_13766);
nand UO_669 (O_669,N_13563,N_13970);
and UO_670 (O_670,N_14842,N_14634);
or UO_671 (O_671,N_14291,N_13888);
nand UO_672 (O_672,N_14998,N_14840);
or UO_673 (O_673,N_14251,N_13778);
nor UO_674 (O_674,N_13997,N_14292);
or UO_675 (O_675,N_13818,N_14902);
nor UO_676 (O_676,N_14747,N_14653);
and UO_677 (O_677,N_13725,N_14289);
nand UO_678 (O_678,N_14721,N_13914);
nand UO_679 (O_679,N_13713,N_13760);
xnor UO_680 (O_680,N_14818,N_14920);
xor UO_681 (O_681,N_13569,N_14651);
nand UO_682 (O_682,N_14213,N_14198);
or UO_683 (O_683,N_14522,N_14500);
and UO_684 (O_684,N_14415,N_14015);
nand UO_685 (O_685,N_14730,N_14309);
xnor UO_686 (O_686,N_14855,N_14250);
or UO_687 (O_687,N_14994,N_14697);
or UO_688 (O_688,N_14427,N_14487);
and UO_689 (O_689,N_14018,N_14852);
and UO_690 (O_690,N_13944,N_13808);
nand UO_691 (O_691,N_14120,N_14982);
nand UO_692 (O_692,N_14506,N_14556);
nand UO_693 (O_693,N_14798,N_13945);
nand UO_694 (O_694,N_13581,N_14547);
or UO_695 (O_695,N_14162,N_13951);
xor UO_696 (O_696,N_14549,N_13741);
nor UO_697 (O_697,N_14194,N_14242);
nor UO_698 (O_698,N_13598,N_14241);
xor UO_699 (O_699,N_14847,N_13553);
nor UO_700 (O_700,N_14662,N_14079);
nor UO_701 (O_701,N_13530,N_13695);
nand UO_702 (O_702,N_14893,N_13555);
nor UO_703 (O_703,N_13849,N_14934);
xnor UO_704 (O_704,N_14060,N_14707);
xor UO_705 (O_705,N_14324,N_14113);
nand UO_706 (O_706,N_14775,N_13878);
or UO_707 (O_707,N_14039,N_14716);
or UO_708 (O_708,N_14461,N_14479);
nor UO_709 (O_709,N_14206,N_13960);
xor UO_710 (O_710,N_13508,N_14872);
nor UO_711 (O_711,N_13797,N_14013);
and UO_712 (O_712,N_13931,N_14883);
or UO_713 (O_713,N_14139,N_14870);
and UO_714 (O_714,N_14937,N_14825);
and UO_715 (O_715,N_13803,N_14518);
nand UO_716 (O_716,N_14948,N_14069);
nor UO_717 (O_717,N_14450,N_13634);
or UO_718 (O_718,N_14280,N_13962);
or UO_719 (O_719,N_14705,N_14873);
nand UO_720 (O_720,N_14900,N_13966);
nor UO_721 (O_721,N_14032,N_13546);
nor UO_722 (O_722,N_13959,N_14091);
or UO_723 (O_723,N_14622,N_14480);
nor UO_724 (O_724,N_14812,N_14584);
nor UO_725 (O_725,N_13795,N_14502);
and UO_726 (O_726,N_14175,N_14266);
nand UO_727 (O_727,N_14278,N_14019);
xor UO_728 (O_728,N_13937,N_14822);
nand UO_729 (O_729,N_13565,N_14961);
nand UO_730 (O_730,N_13726,N_13834);
nor UO_731 (O_731,N_14221,N_14607);
nand UO_732 (O_732,N_14265,N_14851);
nand UO_733 (O_733,N_13994,N_14431);
or UO_734 (O_734,N_14049,N_14808);
or UO_735 (O_735,N_14472,N_14315);
and UO_736 (O_736,N_13502,N_14508);
or UO_737 (O_737,N_14766,N_14597);
and UO_738 (O_738,N_14857,N_14858);
and UO_739 (O_739,N_14482,N_13519);
and UO_740 (O_740,N_14657,N_14322);
xnor UO_741 (O_741,N_14365,N_14546);
nor UO_742 (O_742,N_14567,N_13574);
and UO_743 (O_743,N_14282,N_14027);
or UO_744 (O_744,N_13990,N_14601);
and UO_745 (O_745,N_14871,N_14956);
and UO_746 (O_746,N_13858,N_14367);
nand UO_747 (O_747,N_14953,N_14094);
and UO_748 (O_748,N_13684,N_14222);
nor UO_749 (O_749,N_14371,N_14414);
nor UO_750 (O_750,N_14253,N_13959);
and UO_751 (O_751,N_14840,N_14541);
or UO_752 (O_752,N_14671,N_13807);
xor UO_753 (O_753,N_14156,N_13515);
xor UO_754 (O_754,N_13952,N_13619);
nand UO_755 (O_755,N_13657,N_14976);
and UO_756 (O_756,N_14687,N_14240);
and UO_757 (O_757,N_13915,N_14935);
xnor UO_758 (O_758,N_13743,N_14658);
and UO_759 (O_759,N_14436,N_13897);
xnor UO_760 (O_760,N_14800,N_14558);
nor UO_761 (O_761,N_14707,N_14243);
xnor UO_762 (O_762,N_13586,N_13555);
nor UO_763 (O_763,N_14784,N_13592);
and UO_764 (O_764,N_14977,N_13514);
and UO_765 (O_765,N_14280,N_14419);
and UO_766 (O_766,N_13917,N_14894);
xnor UO_767 (O_767,N_14177,N_14364);
nand UO_768 (O_768,N_14835,N_13878);
or UO_769 (O_769,N_13553,N_14514);
xor UO_770 (O_770,N_14882,N_14593);
and UO_771 (O_771,N_13639,N_14042);
nand UO_772 (O_772,N_13928,N_14643);
nor UO_773 (O_773,N_14066,N_13578);
nor UO_774 (O_774,N_14907,N_14110);
nand UO_775 (O_775,N_13632,N_14101);
xnor UO_776 (O_776,N_14264,N_13516);
nand UO_777 (O_777,N_14883,N_13933);
or UO_778 (O_778,N_14288,N_14038);
xor UO_779 (O_779,N_14890,N_14334);
and UO_780 (O_780,N_14318,N_14014);
nor UO_781 (O_781,N_13766,N_13793);
nor UO_782 (O_782,N_13715,N_13972);
nor UO_783 (O_783,N_14415,N_14503);
nand UO_784 (O_784,N_14912,N_14242);
and UO_785 (O_785,N_14997,N_13621);
or UO_786 (O_786,N_13559,N_14660);
nor UO_787 (O_787,N_14403,N_14572);
and UO_788 (O_788,N_14150,N_14539);
nand UO_789 (O_789,N_14471,N_13908);
or UO_790 (O_790,N_14619,N_13688);
xor UO_791 (O_791,N_13985,N_14343);
xnor UO_792 (O_792,N_14794,N_14986);
nor UO_793 (O_793,N_13825,N_14114);
nand UO_794 (O_794,N_14081,N_14098);
nand UO_795 (O_795,N_13837,N_13669);
nand UO_796 (O_796,N_14437,N_13580);
nor UO_797 (O_797,N_14019,N_13865);
xnor UO_798 (O_798,N_14583,N_13943);
nand UO_799 (O_799,N_14500,N_13987);
nand UO_800 (O_800,N_14115,N_13799);
xor UO_801 (O_801,N_14072,N_14905);
xnor UO_802 (O_802,N_14541,N_14822);
nand UO_803 (O_803,N_13975,N_14219);
nand UO_804 (O_804,N_14389,N_14670);
or UO_805 (O_805,N_14435,N_13593);
or UO_806 (O_806,N_14155,N_14117);
nor UO_807 (O_807,N_13657,N_14144);
xor UO_808 (O_808,N_13675,N_13832);
nor UO_809 (O_809,N_14831,N_14980);
xnor UO_810 (O_810,N_14724,N_14237);
and UO_811 (O_811,N_14055,N_14529);
nor UO_812 (O_812,N_14910,N_14479);
xor UO_813 (O_813,N_13881,N_14218);
or UO_814 (O_814,N_14868,N_14881);
or UO_815 (O_815,N_13645,N_13524);
nor UO_816 (O_816,N_13747,N_14993);
nand UO_817 (O_817,N_14004,N_13820);
or UO_818 (O_818,N_14371,N_13743);
xnor UO_819 (O_819,N_14445,N_14212);
or UO_820 (O_820,N_14819,N_14417);
xor UO_821 (O_821,N_14702,N_13892);
nor UO_822 (O_822,N_14198,N_14961);
xnor UO_823 (O_823,N_13893,N_13962);
nand UO_824 (O_824,N_14275,N_14636);
nor UO_825 (O_825,N_14535,N_14026);
or UO_826 (O_826,N_14827,N_14697);
or UO_827 (O_827,N_14465,N_13703);
nand UO_828 (O_828,N_13566,N_14728);
or UO_829 (O_829,N_14947,N_14873);
nor UO_830 (O_830,N_14665,N_14478);
nand UO_831 (O_831,N_13852,N_14966);
and UO_832 (O_832,N_14532,N_13679);
or UO_833 (O_833,N_13711,N_14299);
or UO_834 (O_834,N_13535,N_13672);
xor UO_835 (O_835,N_14411,N_14899);
xor UO_836 (O_836,N_13715,N_14169);
nand UO_837 (O_837,N_13513,N_14463);
xnor UO_838 (O_838,N_14645,N_14152);
nor UO_839 (O_839,N_14942,N_14934);
or UO_840 (O_840,N_13912,N_14367);
or UO_841 (O_841,N_13584,N_14962);
xor UO_842 (O_842,N_14659,N_14947);
and UO_843 (O_843,N_14964,N_14686);
xnor UO_844 (O_844,N_13779,N_13757);
nand UO_845 (O_845,N_13515,N_13594);
xor UO_846 (O_846,N_14603,N_14289);
nor UO_847 (O_847,N_13838,N_14283);
nand UO_848 (O_848,N_14729,N_14625);
xnor UO_849 (O_849,N_13904,N_13768);
or UO_850 (O_850,N_14095,N_14255);
xor UO_851 (O_851,N_14176,N_13983);
xnor UO_852 (O_852,N_14225,N_14640);
or UO_853 (O_853,N_13872,N_14144);
nor UO_854 (O_854,N_14440,N_13667);
xnor UO_855 (O_855,N_14926,N_13694);
xnor UO_856 (O_856,N_14127,N_13918);
or UO_857 (O_857,N_14409,N_14531);
xnor UO_858 (O_858,N_14749,N_14511);
xor UO_859 (O_859,N_14044,N_13766);
xor UO_860 (O_860,N_14837,N_14486);
and UO_861 (O_861,N_14670,N_14263);
nor UO_862 (O_862,N_13637,N_14699);
nor UO_863 (O_863,N_14313,N_14075);
nor UO_864 (O_864,N_14763,N_14465);
xnor UO_865 (O_865,N_13781,N_13532);
or UO_866 (O_866,N_14702,N_14763);
xnor UO_867 (O_867,N_14588,N_14095);
nand UO_868 (O_868,N_14004,N_14008);
or UO_869 (O_869,N_13519,N_13637);
xnor UO_870 (O_870,N_13820,N_14870);
nor UO_871 (O_871,N_14054,N_14442);
nor UO_872 (O_872,N_14316,N_13554);
or UO_873 (O_873,N_14704,N_14893);
nor UO_874 (O_874,N_14867,N_13943);
xnor UO_875 (O_875,N_14333,N_14054);
and UO_876 (O_876,N_14590,N_14591);
and UO_877 (O_877,N_14496,N_13682);
nor UO_878 (O_878,N_14176,N_13510);
nand UO_879 (O_879,N_13528,N_14703);
and UO_880 (O_880,N_14637,N_14607);
and UO_881 (O_881,N_14399,N_14850);
and UO_882 (O_882,N_14451,N_14697);
nand UO_883 (O_883,N_14114,N_13590);
nand UO_884 (O_884,N_13814,N_14341);
and UO_885 (O_885,N_14590,N_14053);
and UO_886 (O_886,N_13660,N_13856);
or UO_887 (O_887,N_14211,N_13737);
nor UO_888 (O_888,N_14935,N_13500);
or UO_889 (O_889,N_14115,N_13904);
xnor UO_890 (O_890,N_13767,N_14733);
xnor UO_891 (O_891,N_14794,N_13988);
nor UO_892 (O_892,N_13754,N_14981);
or UO_893 (O_893,N_14323,N_14739);
nand UO_894 (O_894,N_13970,N_14477);
and UO_895 (O_895,N_13885,N_14686);
or UO_896 (O_896,N_14157,N_14989);
nand UO_897 (O_897,N_13958,N_14336);
nor UO_898 (O_898,N_14060,N_14829);
nor UO_899 (O_899,N_13836,N_14171);
or UO_900 (O_900,N_13556,N_13562);
nand UO_901 (O_901,N_13928,N_14551);
and UO_902 (O_902,N_13937,N_13952);
nor UO_903 (O_903,N_14770,N_14585);
nor UO_904 (O_904,N_13850,N_14322);
and UO_905 (O_905,N_14062,N_14999);
nor UO_906 (O_906,N_13830,N_13833);
nand UO_907 (O_907,N_13962,N_14951);
or UO_908 (O_908,N_13897,N_13669);
and UO_909 (O_909,N_13622,N_14223);
and UO_910 (O_910,N_14313,N_14842);
nand UO_911 (O_911,N_14117,N_14229);
and UO_912 (O_912,N_14151,N_14491);
nand UO_913 (O_913,N_14059,N_14698);
or UO_914 (O_914,N_14856,N_14899);
and UO_915 (O_915,N_13725,N_14525);
nand UO_916 (O_916,N_14508,N_14429);
nor UO_917 (O_917,N_14162,N_14429);
nor UO_918 (O_918,N_14558,N_13686);
and UO_919 (O_919,N_13626,N_14513);
nand UO_920 (O_920,N_13583,N_14323);
nand UO_921 (O_921,N_14575,N_14678);
or UO_922 (O_922,N_14678,N_14665);
or UO_923 (O_923,N_14030,N_13647);
nand UO_924 (O_924,N_14671,N_14077);
and UO_925 (O_925,N_14610,N_14095);
and UO_926 (O_926,N_14305,N_13828);
and UO_927 (O_927,N_13986,N_14765);
nor UO_928 (O_928,N_13874,N_13762);
and UO_929 (O_929,N_13983,N_14622);
xnor UO_930 (O_930,N_14942,N_14958);
nand UO_931 (O_931,N_14444,N_13912);
xnor UO_932 (O_932,N_13931,N_14343);
nor UO_933 (O_933,N_13529,N_13609);
and UO_934 (O_934,N_14974,N_14399);
and UO_935 (O_935,N_13903,N_14163);
or UO_936 (O_936,N_14902,N_14485);
xor UO_937 (O_937,N_14275,N_14402);
and UO_938 (O_938,N_14430,N_14227);
nor UO_939 (O_939,N_13695,N_14102);
nor UO_940 (O_940,N_14091,N_14108);
nor UO_941 (O_941,N_14636,N_14601);
xnor UO_942 (O_942,N_13989,N_13825);
and UO_943 (O_943,N_14503,N_14485);
and UO_944 (O_944,N_13617,N_14511);
nor UO_945 (O_945,N_14456,N_13789);
nor UO_946 (O_946,N_14381,N_14526);
or UO_947 (O_947,N_14010,N_14315);
xnor UO_948 (O_948,N_14638,N_13886);
nor UO_949 (O_949,N_13521,N_14425);
or UO_950 (O_950,N_14770,N_14932);
xor UO_951 (O_951,N_14732,N_14600);
or UO_952 (O_952,N_13536,N_13580);
xnor UO_953 (O_953,N_13823,N_13548);
or UO_954 (O_954,N_13525,N_14897);
nand UO_955 (O_955,N_14882,N_14451);
nand UO_956 (O_956,N_13597,N_14707);
and UO_957 (O_957,N_14403,N_13679);
and UO_958 (O_958,N_14676,N_14865);
and UO_959 (O_959,N_13855,N_13586);
nand UO_960 (O_960,N_14264,N_14190);
xor UO_961 (O_961,N_14410,N_14023);
nand UO_962 (O_962,N_14639,N_13971);
and UO_963 (O_963,N_14267,N_14926);
xor UO_964 (O_964,N_13501,N_13969);
and UO_965 (O_965,N_14856,N_14425);
nand UO_966 (O_966,N_14981,N_13590);
or UO_967 (O_967,N_14789,N_14089);
xor UO_968 (O_968,N_14502,N_13667);
xor UO_969 (O_969,N_14267,N_14096);
or UO_970 (O_970,N_14788,N_14872);
or UO_971 (O_971,N_14667,N_13877);
and UO_972 (O_972,N_14054,N_14306);
and UO_973 (O_973,N_13605,N_14506);
nor UO_974 (O_974,N_14053,N_14470);
nor UO_975 (O_975,N_14849,N_14293);
and UO_976 (O_976,N_14454,N_14943);
and UO_977 (O_977,N_13990,N_13759);
nand UO_978 (O_978,N_14492,N_14420);
nand UO_979 (O_979,N_14725,N_14197);
xnor UO_980 (O_980,N_14353,N_14833);
xor UO_981 (O_981,N_13794,N_14435);
or UO_982 (O_982,N_13831,N_13819);
and UO_983 (O_983,N_14285,N_14055);
nand UO_984 (O_984,N_14410,N_14595);
nand UO_985 (O_985,N_14981,N_13700);
nand UO_986 (O_986,N_14501,N_14924);
nand UO_987 (O_987,N_14209,N_14790);
nand UO_988 (O_988,N_14229,N_14948);
nor UO_989 (O_989,N_13848,N_14958);
nor UO_990 (O_990,N_14926,N_14502);
and UO_991 (O_991,N_13930,N_14711);
nor UO_992 (O_992,N_14327,N_14549);
or UO_993 (O_993,N_14868,N_13953);
nor UO_994 (O_994,N_14950,N_14545);
nand UO_995 (O_995,N_14728,N_13513);
nand UO_996 (O_996,N_14291,N_14116);
nor UO_997 (O_997,N_14116,N_14293);
xnor UO_998 (O_998,N_13523,N_13971);
and UO_999 (O_999,N_13803,N_13852);
and UO_1000 (O_1000,N_13782,N_14922);
nor UO_1001 (O_1001,N_14795,N_13982);
xor UO_1002 (O_1002,N_14734,N_13585);
or UO_1003 (O_1003,N_14878,N_13564);
nor UO_1004 (O_1004,N_14943,N_13665);
xor UO_1005 (O_1005,N_14697,N_14592);
or UO_1006 (O_1006,N_14898,N_14320);
nor UO_1007 (O_1007,N_14856,N_13994);
xnor UO_1008 (O_1008,N_14670,N_13588);
or UO_1009 (O_1009,N_14105,N_13656);
nand UO_1010 (O_1010,N_14743,N_14818);
xnor UO_1011 (O_1011,N_14487,N_14380);
nor UO_1012 (O_1012,N_14123,N_13862);
and UO_1013 (O_1013,N_14021,N_14447);
xnor UO_1014 (O_1014,N_14117,N_13546);
or UO_1015 (O_1015,N_13657,N_13695);
or UO_1016 (O_1016,N_13867,N_14000);
or UO_1017 (O_1017,N_13999,N_13710);
nor UO_1018 (O_1018,N_14026,N_14832);
nand UO_1019 (O_1019,N_14537,N_13866);
nor UO_1020 (O_1020,N_14526,N_14241);
xnor UO_1021 (O_1021,N_13996,N_14746);
nand UO_1022 (O_1022,N_13792,N_13778);
nand UO_1023 (O_1023,N_14161,N_14421);
xnor UO_1024 (O_1024,N_13729,N_14535);
xnor UO_1025 (O_1025,N_14934,N_14663);
nor UO_1026 (O_1026,N_13955,N_14743);
and UO_1027 (O_1027,N_14240,N_14545);
or UO_1028 (O_1028,N_13662,N_14322);
and UO_1029 (O_1029,N_14153,N_13655);
nand UO_1030 (O_1030,N_14473,N_13858);
and UO_1031 (O_1031,N_13935,N_14675);
nor UO_1032 (O_1032,N_14882,N_13959);
nor UO_1033 (O_1033,N_14858,N_14094);
nor UO_1034 (O_1034,N_13885,N_13535);
or UO_1035 (O_1035,N_13775,N_14422);
or UO_1036 (O_1036,N_14831,N_13599);
nor UO_1037 (O_1037,N_14342,N_13823);
and UO_1038 (O_1038,N_13529,N_14745);
nand UO_1039 (O_1039,N_13761,N_14579);
nor UO_1040 (O_1040,N_13759,N_14710);
xor UO_1041 (O_1041,N_14277,N_13813);
xnor UO_1042 (O_1042,N_14429,N_14164);
nor UO_1043 (O_1043,N_13770,N_13560);
xor UO_1044 (O_1044,N_14583,N_14501);
xnor UO_1045 (O_1045,N_14825,N_13667);
nand UO_1046 (O_1046,N_14584,N_14084);
or UO_1047 (O_1047,N_14648,N_13778);
nand UO_1048 (O_1048,N_14559,N_14210);
and UO_1049 (O_1049,N_14707,N_14650);
xor UO_1050 (O_1050,N_13708,N_14999);
or UO_1051 (O_1051,N_13595,N_13659);
nand UO_1052 (O_1052,N_14977,N_14264);
nor UO_1053 (O_1053,N_13791,N_14945);
xor UO_1054 (O_1054,N_13652,N_14660);
nor UO_1055 (O_1055,N_13768,N_13912);
nor UO_1056 (O_1056,N_13766,N_14917);
and UO_1057 (O_1057,N_13995,N_13759);
nand UO_1058 (O_1058,N_14442,N_13776);
nand UO_1059 (O_1059,N_13922,N_13526);
nand UO_1060 (O_1060,N_14432,N_13512);
xor UO_1061 (O_1061,N_14571,N_14243);
nand UO_1062 (O_1062,N_13942,N_14946);
nor UO_1063 (O_1063,N_13578,N_14646);
xor UO_1064 (O_1064,N_14119,N_14402);
nor UO_1065 (O_1065,N_14546,N_14770);
nand UO_1066 (O_1066,N_14548,N_14645);
and UO_1067 (O_1067,N_14944,N_13967);
xnor UO_1068 (O_1068,N_14017,N_14300);
nor UO_1069 (O_1069,N_14622,N_14824);
nand UO_1070 (O_1070,N_14574,N_14878);
or UO_1071 (O_1071,N_13597,N_14414);
nand UO_1072 (O_1072,N_14361,N_13987);
xor UO_1073 (O_1073,N_14349,N_14724);
nand UO_1074 (O_1074,N_14985,N_13687);
nor UO_1075 (O_1075,N_14079,N_14536);
nor UO_1076 (O_1076,N_13904,N_13912);
nand UO_1077 (O_1077,N_14350,N_14862);
nor UO_1078 (O_1078,N_13591,N_14104);
and UO_1079 (O_1079,N_14032,N_13627);
xnor UO_1080 (O_1080,N_13909,N_14543);
xor UO_1081 (O_1081,N_14215,N_14927);
xnor UO_1082 (O_1082,N_14055,N_14869);
nor UO_1083 (O_1083,N_14615,N_13906);
nor UO_1084 (O_1084,N_13697,N_14320);
or UO_1085 (O_1085,N_14611,N_13836);
nand UO_1086 (O_1086,N_14293,N_14901);
xnor UO_1087 (O_1087,N_14737,N_14744);
or UO_1088 (O_1088,N_14948,N_13738);
or UO_1089 (O_1089,N_14817,N_14333);
and UO_1090 (O_1090,N_14443,N_13765);
and UO_1091 (O_1091,N_13838,N_13646);
and UO_1092 (O_1092,N_13871,N_14349);
xor UO_1093 (O_1093,N_13532,N_14328);
nor UO_1094 (O_1094,N_14624,N_13994);
or UO_1095 (O_1095,N_13632,N_14331);
xor UO_1096 (O_1096,N_13981,N_13609);
and UO_1097 (O_1097,N_14928,N_13881);
and UO_1098 (O_1098,N_13944,N_14147);
or UO_1099 (O_1099,N_14179,N_14597);
and UO_1100 (O_1100,N_14597,N_13505);
nor UO_1101 (O_1101,N_14925,N_14195);
nand UO_1102 (O_1102,N_14116,N_14251);
nor UO_1103 (O_1103,N_14820,N_13801);
and UO_1104 (O_1104,N_14115,N_14917);
nor UO_1105 (O_1105,N_13802,N_14054);
nor UO_1106 (O_1106,N_13948,N_14718);
nor UO_1107 (O_1107,N_14871,N_14252);
xnor UO_1108 (O_1108,N_14784,N_13942);
xor UO_1109 (O_1109,N_14693,N_13800);
or UO_1110 (O_1110,N_14452,N_14683);
nand UO_1111 (O_1111,N_13643,N_14596);
and UO_1112 (O_1112,N_14779,N_13609);
nand UO_1113 (O_1113,N_13840,N_14791);
and UO_1114 (O_1114,N_14621,N_13606);
or UO_1115 (O_1115,N_13843,N_14177);
nand UO_1116 (O_1116,N_13542,N_13607);
or UO_1117 (O_1117,N_13549,N_14769);
or UO_1118 (O_1118,N_13808,N_13795);
xnor UO_1119 (O_1119,N_13867,N_14518);
xor UO_1120 (O_1120,N_14005,N_14373);
nand UO_1121 (O_1121,N_14517,N_13754);
or UO_1122 (O_1122,N_13545,N_14489);
or UO_1123 (O_1123,N_14644,N_14447);
nand UO_1124 (O_1124,N_13912,N_14020);
xnor UO_1125 (O_1125,N_14850,N_13574);
or UO_1126 (O_1126,N_14033,N_14454);
xnor UO_1127 (O_1127,N_14840,N_14456);
nor UO_1128 (O_1128,N_14674,N_14497);
xnor UO_1129 (O_1129,N_13770,N_14138);
xor UO_1130 (O_1130,N_14644,N_14155);
xnor UO_1131 (O_1131,N_14877,N_13876);
nand UO_1132 (O_1132,N_14350,N_13705);
nor UO_1133 (O_1133,N_14156,N_14247);
xnor UO_1134 (O_1134,N_14503,N_14701);
nand UO_1135 (O_1135,N_13976,N_13595);
xor UO_1136 (O_1136,N_14567,N_14218);
and UO_1137 (O_1137,N_14100,N_14462);
nand UO_1138 (O_1138,N_13938,N_14018);
nand UO_1139 (O_1139,N_13984,N_14755);
nand UO_1140 (O_1140,N_13564,N_14486);
nand UO_1141 (O_1141,N_14105,N_13667);
or UO_1142 (O_1142,N_14807,N_14295);
nand UO_1143 (O_1143,N_14643,N_14366);
nor UO_1144 (O_1144,N_13758,N_13917);
and UO_1145 (O_1145,N_14556,N_14654);
nor UO_1146 (O_1146,N_14028,N_13835);
nand UO_1147 (O_1147,N_14036,N_14362);
xnor UO_1148 (O_1148,N_14344,N_13973);
and UO_1149 (O_1149,N_13859,N_14569);
or UO_1150 (O_1150,N_14894,N_13720);
nor UO_1151 (O_1151,N_14297,N_14676);
nand UO_1152 (O_1152,N_13580,N_14784);
nor UO_1153 (O_1153,N_14236,N_13756);
nor UO_1154 (O_1154,N_13569,N_13881);
or UO_1155 (O_1155,N_14799,N_13505);
nand UO_1156 (O_1156,N_14092,N_14583);
xnor UO_1157 (O_1157,N_13746,N_14593);
xnor UO_1158 (O_1158,N_14813,N_14209);
or UO_1159 (O_1159,N_14524,N_14984);
xnor UO_1160 (O_1160,N_14762,N_13571);
or UO_1161 (O_1161,N_13574,N_13957);
or UO_1162 (O_1162,N_13611,N_14634);
xnor UO_1163 (O_1163,N_14393,N_13905);
and UO_1164 (O_1164,N_14611,N_14771);
or UO_1165 (O_1165,N_14049,N_14154);
and UO_1166 (O_1166,N_14681,N_14744);
nor UO_1167 (O_1167,N_14329,N_13586);
nor UO_1168 (O_1168,N_13841,N_14721);
xnor UO_1169 (O_1169,N_14540,N_14610);
and UO_1170 (O_1170,N_14176,N_13947);
and UO_1171 (O_1171,N_13911,N_13509);
xnor UO_1172 (O_1172,N_14628,N_14636);
or UO_1173 (O_1173,N_14940,N_14394);
nor UO_1174 (O_1174,N_13659,N_14206);
xor UO_1175 (O_1175,N_13670,N_14730);
or UO_1176 (O_1176,N_14991,N_13602);
or UO_1177 (O_1177,N_14806,N_14724);
nor UO_1178 (O_1178,N_14729,N_13829);
xnor UO_1179 (O_1179,N_13859,N_14878);
or UO_1180 (O_1180,N_13636,N_14877);
xnor UO_1181 (O_1181,N_13668,N_14461);
nor UO_1182 (O_1182,N_13564,N_14511);
or UO_1183 (O_1183,N_13757,N_14563);
and UO_1184 (O_1184,N_14515,N_14090);
or UO_1185 (O_1185,N_14989,N_14387);
or UO_1186 (O_1186,N_13869,N_14574);
and UO_1187 (O_1187,N_14413,N_14546);
xor UO_1188 (O_1188,N_13876,N_14619);
xnor UO_1189 (O_1189,N_14839,N_14214);
nor UO_1190 (O_1190,N_14785,N_14001);
nor UO_1191 (O_1191,N_13789,N_14482);
nor UO_1192 (O_1192,N_13888,N_13657);
nor UO_1193 (O_1193,N_14342,N_14598);
xnor UO_1194 (O_1194,N_14623,N_13942);
and UO_1195 (O_1195,N_13516,N_13791);
nand UO_1196 (O_1196,N_14043,N_14681);
nand UO_1197 (O_1197,N_14443,N_14185);
nand UO_1198 (O_1198,N_14770,N_14922);
nor UO_1199 (O_1199,N_14733,N_13891);
and UO_1200 (O_1200,N_13991,N_14284);
or UO_1201 (O_1201,N_13879,N_14067);
or UO_1202 (O_1202,N_13571,N_14456);
nand UO_1203 (O_1203,N_14805,N_14060);
or UO_1204 (O_1204,N_13736,N_14318);
and UO_1205 (O_1205,N_14348,N_14279);
xor UO_1206 (O_1206,N_13546,N_14972);
and UO_1207 (O_1207,N_14402,N_14087);
nor UO_1208 (O_1208,N_13764,N_13801);
xor UO_1209 (O_1209,N_14580,N_14080);
nand UO_1210 (O_1210,N_14218,N_14489);
nor UO_1211 (O_1211,N_14694,N_14774);
or UO_1212 (O_1212,N_13855,N_14043);
nand UO_1213 (O_1213,N_14997,N_13694);
and UO_1214 (O_1214,N_14056,N_13855);
or UO_1215 (O_1215,N_13730,N_14156);
or UO_1216 (O_1216,N_13589,N_14972);
nand UO_1217 (O_1217,N_14355,N_13706);
and UO_1218 (O_1218,N_14204,N_14190);
nand UO_1219 (O_1219,N_14665,N_14013);
xnor UO_1220 (O_1220,N_14628,N_14614);
or UO_1221 (O_1221,N_14871,N_14142);
nand UO_1222 (O_1222,N_14631,N_14065);
nand UO_1223 (O_1223,N_14952,N_14650);
and UO_1224 (O_1224,N_13986,N_14210);
and UO_1225 (O_1225,N_13815,N_14056);
and UO_1226 (O_1226,N_13639,N_14621);
or UO_1227 (O_1227,N_13918,N_14266);
nor UO_1228 (O_1228,N_13536,N_14541);
nand UO_1229 (O_1229,N_14219,N_14592);
nand UO_1230 (O_1230,N_13908,N_13768);
nand UO_1231 (O_1231,N_14819,N_14525);
nor UO_1232 (O_1232,N_14994,N_14361);
nor UO_1233 (O_1233,N_14788,N_13716);
or UO_1234 (O_1234,N_14341,N_14050);
nor UO_1235 (O_1235,N_13978,N_14435);
or UO_1236 (O_1236,N_14037,N_14177);
nor UO_1237 (O_1237,N_14242,N_14187);
xor UO_1238 (O_1238,N_14814,N_14723);
and UO_1239 (O_1239,N_14863,N_13633);
xor UO_1240 (O_1240,N_14321,N_14954);
xor UO_1241 (O_1241,N_14165,N_13763);
nand UO_1242 (O_1242,N_14641,N_14234);
or UO_1243 (O_1243,N_14564,N_14733);
nand UO_1244 (O_1244,N_14136,N_14301);
or UO_1245 (O_1245,N_14101,N_14624);
nand UO_1246 (O_1246,N_13599,N_14033);
xor UO_1247 (O_1247,N_14157,N_13970);
or UO_1248 (O_1248,N_14172,N_14005);
nor UO_1249 (O_1249,N_14476,N_14943);
or UO_1250 (O_1250,N_14355,N_14791);
nand UO_1251 (O_1251,N_14456,N_14926);
nand UO_1252 (O_1252,N_13737,N_13755);
xnor UO_1253 (O_1253,N_13747,N_14068);
or UO_1254 (O_1254,N_13771,N_14057);
nand UO_1255 (O_1255,N_14000,N_14862);
nand UO_1256 (O_1256,N_14603,N_14556);
xor UO_1257 (O_1257,N_13532,N_13581);
nor UO_1258 (O_1258,N_13691,N_14794);
xor UO_1259 (O_1259,N_14659,N_14443);
nor UO_1260 (O_1260,N_14090,N_14743);
or UO_1261 (O_1261,N_14330,N_14346);
and UO_1262 (O_1262,N_13830,N_13861);
nor UO_1263 (O_1263,N_14930,N_14835);
or UO_1264 (O_1264,N_14621,N_13537);
and UO_1265 (O_1265,N_14899,N_13649);
nor UO_1266 (O_1266,N_14897,N_13818);
nand UO_1267 (O_1267,N_14523,N_14645);
or UO_1268 (O_1268,N_14995,N_13869);
and UO_1269 (O_1269,N_14656,N_13643);
nor UO_1270 (O_1270,N_13711,N_13585);
nor UO_1271 (O_1271,N_14456,N_13750);
or UO_1272 (O_1272,N_13775,N_14135);
xor UO_1273 (O_1273,N_13852,N_14065);
nor UO_1274 (O_1274,N_14240,N_14671);
nand UO_1275 (O_1275,N_14541,N_14147);
xnor UO_1276 (O_1276,N_14338,N_13712);
and UO_1277 (O_1277,N_14395,N_14962);
nand UO_1278 (O_1278,N_14314,N_14892);
nand UO_1279 (O_1279,N_14617,N_14975);
or UO_1280 (O_1280,N_13671,N_14572);
and UO_1281 (O_1281,N_14419,N_14374);
xnor UO_1282 (O_1282,N_14144,N_13809);
and UO_1283 (O_1283,N_13981,N_13514);
nand UO_1284 (O_1284,N_14542,N_14693);
nand UO_1285 (O_1285,N_13727,N_14342);
or UO_1286 (O_1286,N_13594,N_14680);
nor UO_1287 (O_1287,N_13873,N_13712);
or UO_1288 (O_1288,N_13694,N_13608);
and UO_1289 (O_1289,N_13774,N_14997);
nand UO_1290 (O_1290,N_14033,N_13907);
and UO_1291 (O_1291,N_14621,N_14225);
nand UO_1292 (O_1292,N_13798,N_14215);
and UO_1293 (O_1293,N_13917,N_13572);
xor UO_1294 (O_1294,N_13761,N_14336);
or UO_1295 (O_1295,N_14579,N_13539);
nand UO_1296 (O_1296,N_14018,N_13517);
and UO_1297 (O_1297,N_13749,N_13822);
nand UO_1298 (O_1298,N_13978,N_13899);
nor UO_1299 (O_1299,N_13714,N_14577);
nand UO_1300 (O_1300,N_14600,N_13937);
xnor UO_1301 (O_1301,N_14606,N_14500);
xor UO_1302 (O_1302,N_13520,N_14987);
or UO_1303 (O_1303,N_14236,N_13910);
or UO_1304 (O_1304,N_14472,N_14823);
xor UO_1305 (O_1305,N_14991,N_14983);
nand UO_1306 (O_1306,N_14897,N_14078);
nor UO_1307 (O_1307,N_14452,N_14672);
nor UO_1308 (O_1308,N_14096,N_13526);
xnor UO_1309 (O_1309,N_13811,N_14100);
nor UO_1310 (O_1310,N_14466,N_14166);
nand UO_1311 (O_1311,N_14678,N_13860);
xnor UO_1312 (O_1312,N_14011,N_13581);
and UO_1313 (O_1313,N_14687,N_13697);
xnor UO_1314 (O_1314,N_13536,N_13821);
xnor UO_1315 (O_1315,N_14426,N_14052);
and UO_1316 (O_1316,N_14714,N_14162);
or UO_1317 (O_1317,N_13829,N_14413);
nor UO_1318 (O_1318,N_14262,N_14452);
nor UO_1319 (O_1319,N_13705,N_14672);
nor UO_1320 (O_1320,N_13560,N_13733);
xnor UO_1321 (O_1321,N_14941,N_14885);
or UO_1322 (O_1322,N_14634,N_13627);
and UO_1323 (O_1323,N_14763,N_14065);
nor UO_1324 (O_1324,N_14591,N_13803);
nand UO_1325 (O_1325,N_13549,N_14750);
and UO_1326 (O_1326,N_14062,N_13913);
nand UO_1327 (O_1327,N_14951,N_14816);
or UO_1328 (O_1328,N_14647,N_14531);
nand UO_1329 (O_1329,N_14984,N_14694);
nand UO_1330 (O_1330,N_13522,N_14786);
or UO_1331 (O_1331,N_14654,N_13597);
nor UO_1332 (O_1332,N_14849,N_14494);
nand UO_1333 (O_1333,N_14195,N_13508);
or UO_1334 (O_1334,N_14830,N_14048);
and UO_1335 (O_1335,N_13813,N_13671);
xor UO_1336 (O_1336,N_13883,N_13814);
or UO_1337 (O_1337,N_14764,N_14997);
or UO_1338 (O_1338,N_14934,N_14888);
nor UO_1339 (O_1339,N_14457,N_13572);
and UO_1340 (O_1340,N_14067,N_14911);
and UO_1341 (O_1341,N_14372,N_14620);
or UO_1342 (O_1342,N_13869,N_14707);
nand UO_1343 (O_1343,N_14916,N_14776);
nand UO_1344 (O_1344,N_14996,N_14154);
nand UO_1345 (O_1345,N_13512,N_13623);
or UO_1346 (O_1346,N_13507,N_13767);
and UO_1347 (O_1347,N_13629,N_14984);
xnor UO_1348 (O_1348,N_14339,N_14251);
and UO_1349 (O_1349,N_13808,N_14890);
xnor UO_1350 (O_1350,N_14882,N_14311);
and UO_1351 (O_1351,N_14277,N_14874);
and UO_1352 (O_1352,N_14131,N_13528);
and UO_1353 (O_1353,N_13687,N_13506);
nor UO_1354 (O_1354,N_14234,N_13834);
nand UO_1355 (O_1355,N_14107,N_14831);
or UO_1356 (O_1356,N_14839,N_13698);
nand UO_1357 (O_1357,N_14480,N_13885);
or UO_1358 (O_1358,N_13923,N_14818);
nand UO_1359 (O_1359,N_13596,N_13537);
xnor UO_1360 (O_1360,N_14884,N_14045);
xnor UO_1361 (O_1361,N_13529,N_14080);
and UO_1362 (O_1362,N_13732,N_13823);
or UO_1363 (O_1363,N_14506,N_14929);
or UO_1364 (O_1364,N_13935,N_14674);
and UO_1365 (O_1365,N_14825,N_13549);
nand UO_1366 (O_1366,N_14969,N_13667);
and UO_1367 (O_1367,N_13666,N_13549);
or UO_1368 (O_1368,N_14388,N_13797);
or UO_1369 (O_1369,N_13694,N_14900);
or UO_1370 (O_1370,N_14898,N_13533);
and UO_1371 (O_1371,N_14945,N_14574);
or UO_1372 (O_1372,N_14232,N_13840);
nand UO_1373 (O_1373,N_13830,N_14094);
nor UO_1374 (O_1374,N_13914,N_13621);
and UO_1375 (O_1375,N_14515,N_14784);
or UO_1376 (O_1376,N_14851,N_14255);
nor UO_1377 (O_1377,N_14766,N_14477);
nor UO_1378 (O_1378,N_14808,N_14553);
nand UO_1379 (O_1379,N_14499,N_14320);
and UO_1380 (O_1380,N_14177,N_14470);
xor UO_1381 (O_1381,N_14021,N_14361);
xor UO_1382 (O_1382,N_14849,N_14146);
nor UO_1383 (O_1383,N_14358,N_14598);
xor UO_1384 (O_1384,N_14606,N_14282);
nand UO_1385 (O_1385,N_14460,N_14402);
and UO_1386 (O_1386,N_14831,N_14797);
and UO_1387 (O_1387,N_14608,N_14030);
or UO_1388 (O_1388,N_14791,N_13732);
nand UO_1389 (O_1389,N_14245,N_13773);
xor UO_1390 (O_1390,N_14946,N_14428);
nor UO_1391 (O_1391,N_14311,N_14667);
nand UO_1392 (O_1392,N_14500,N_13609);
or UO_1393 (O_1393,N_14300,N_13513);
or UO_1394 (O_1394,N_14790,N_14712);
nand UO_1395 (O_1395,N_14302,N_13515);
nor UO_1396 (O_1396,N_14275,N_13973);
xor UO_1397 (O_1397,N_13831,N_14758);
xor UO_1398 (O_1398,N_13627,N_14143);
nor UO_1399 (O_1399,N_14463,N_14789);
xor UO_1400 (O_1400,N_14208,N_14677);
and UO_1401 (O_1401,N_13861,N_14514);
xor UO_1402 (O_1402,N_14224,N_14687);
xor UO_1403 (O_1403,N_14603,N_13882);
or UO_1404 (O_1404,N_14873,N_14024);
nand UO_1405 (O_1405,N_14716,N_13694);
and UO_1406 (O_1406,N_13965,N_14685);
nor UO_1407 (O_1407,N_13844,N_14899);
nand UO_1408 (O_1408,N_14625,N_13668);
or UO_1409 (O_1409,N_13727,N_14880);
and UO_1410 (O_1410,N_13603,N_14450);
nor UO_1411 (O_1411,N_14414,N_14843);
nor UO_1412 (O_1412,N_14766,N_13738);
and UO_1413 (O_1413,N_13651,N_14249);
xor UO_1414 (O_1414,N_14222,N_14940);
nand UO_1415 (O_1415,N_14281,N_13629);
xnor UO_1416 (O_1416,N_14099,N_13955);
nor UO_1417 (O_1417,N_14771,N_14702);
nor UO_1418 (O_1418,N_13699,N_14044);
nor UO_1419 (O_1419,N_13704,N_14122);
or UO_1420 (O_1420,N_14497,N_14484);
and UO_1421 (O_1421,N_14003,N_14781);
or UO_1422 (O_1422,N_14321,N_14164);
nand UO_1423 (O_1423,N_14385,N_14693);
nor UO_1424 (O_1424,N_14208,N_14626);
nor UO_1425 (O_1425,N_13677,N_14073);
or UO_1426 (O_1426,N_14594,N_14056);
or UO_1427 (O_1427,N_14488,N_13666);
and UO_1428 (O_1428,N_14061,N_13806);
or UO_1429 (O_1429,N_14570,N_13800);
xor UO_1430 (O_1430,N_14118,N_14958);
xnor UO_1431 (O_1431,N_14275,N_14005);
xnor UO_1432 (O_1432,N_14098,N_13807);
or UO_1433 (O_1433,N_13895,N_13727);
nor UO_1434 (O_1434,N_14186,N_13534);
and UO_1435 (O_1435,N_14524,N_14187);
and UO_1436 (O_1436,N_14417,N_13601);
nand UO_1437 (O_1437,N_14110,N_13964);
nand UO_1438 (O_1438,N_13876,N_13557);
and UO_1439 (O_1439,N_14896,N_13675);
or UO_1440 (O_1440,N_14256,N_13653);
or UO_1441 (O_1441,N_14942,N_13629);
and UO_1442 (O_1442,N_13958,N_13951);
xor UO_1443 (O_1443,N_13521,N_13584);
nor UO_1444 (O_1444,N_14133,N_13777);
or UO_1445 (O_1445,N_14761,N_14596);
nor UO_1446 (O_1446,N_13873,N_14286);
or UO_1447 (O_1447,N_14705,N_14011);
or UO_1448 (O_1448,N_14759,N_14276);
xor UO_1449 (O_1449,N_14997,N_14748);
and UO_1450 (O_1450,N_14551,N_13513);
or UO_1451 (O_1451,N_14401,N_14265);
nand UO_1452 (O_1452,N_13737,N_13561);
and UO_1453 (O_1453,N_14057,N_14735);
xnor UO_1454 (O_1454,N_14519,N_14716);
or UO_1455 (O_1455,N_13847,N_13548);
and UO_1456 (O_1456,N_14514,N_14450);
xor UO_1457 (O_1457,N_14528,N_14418);
nand UO_1458 (O_1458,N_14397,N_13902);
xnor UO_1459 (O_1459,N_14597,N_14265);
nand UO_1460 (O_1460,N_14214,N_14907);
xnor UO_1461 (O_1461,N_14479,N_14851);
nand UO_1462 (O_1462,N_13824,N_14955);
xnor UO_1463 (O_1463,N_13580,N_14922);
or UO_1464 (O_1464,N_13967,N_14205);
or UO_1465 (O_1465,N_14886,N_14163);
xor UO_1466 (O_1466,N_13575,N_13596);
and UO_1467 (O_1467,N_13778,N_14356);
nor UO_1468 (O_1468,N_14960,N_14082);
xnor UO_1469 (O_1469,N_14879,N_14821);
xnor UO_1470 (O_1470,N_14418,N_14775);
or UO_1471 (O_1471,N_13624,N_14692);
nand UO_1472 (O_1472,N_14447,N_13570);
xnor UO_1473 (O_1473,N_14034,N_14484);
xnor UO_1474 (O_1474,N_13552,N_13617);
or UO_1475 (O_1475,N_13711,N_14325);
or UO_1476 (O_1476,N_13619,N_13755);
or UO_1477 (O_1477,N_14331,N_14299);
xor UO_1478 (O_1478,N_14144,N_14016);
xor UO_1479 (O_1479,N_14890,N_13646);
nor UO_1480 (O_1480,N_14624,N_14846);
nand UO_1481 (O_1481,N_13723,N_14540);
and UO_1482 (O_1482,N_13694,N_13943);
nor UO_1483 (O_1483,N_14047,N_13675);
nand UO_1484 (O_1484,N_13765,N_14475);
nor UO_1485 (O_1485,N_14680,N_14179);
nand UO_1486 (O_1486,N_13756,N_13577);
nor UO_1487 (O_1487,N_13834,N_14091);
or UO_1488 (O_1488,N_14835,N_14335);
nor UO_1489 (O_1489,N_14419,N_14362);
xor UO_1490 (O_1490,N_13811,N_13534);
nor UO_1491 (O_1491,N_13833,N_14714);
and UO_1492 (O_1492,N_14872,N_13852);
or UO_1493 (O_1493,N_14299,N_14022);
nor UO_1494 (O_1494,N_14813,N_14236);
xnor UO_1495 (O_1495,N_14712,N_14138);
and UO_1496 (O_1496,N_14280,N_14303);
or UO_1497 (O_1497,N_13660,N_14820);
or UO_1498 (O_1498,N_14506,N_14291);
and UO_1499 (O_1499,N_14350,N_14167);
xor UO_1500 (O_1500,N_13528,N_13924);
xnor UO_1501 (O_1501,N_14045,N_13506);
or UO_1502 (O_1502,N_13551,N_13579);
and UO_1503 (O_1503,N_13762,N_14417);
nand UO_1504 (O_1504,N_14465,N_14439);
nand UO_1505 (O_1505,N_14290,N_14095);
and UO_1506 (O_1506,N_13523,N_14326);
and UO_1507 (O_1507,N_14687,N_14593);
nor UO_1508 (O_1508,N_14357,N_13799);
nor UO_1509 (O_1509,N_14244,N_14311);
nand UO_1510 (O_1510,N_14534,N_14493);
and UO_1511 (O_1511,N_14988,N_14151);
nand UO_1512 (O_1512,N_14622,N_14212);
xnor UO_1513 (O_1513,N_14408,N_13627);
nor UO_1514 (O_1514,N_14333,N_14521);
nor UO_1515 (O_1515,N_14291,N_13718);
nand UO_1516 (O_1516,N_14034,N_14809);
nand UO_1517 (O_1517,N_14780,N_13685);
xnor UO_1518 (O_1518,N_13690,N_14788);
nand UO_1519 (O_1519,N_14770,N_13954);
and UO_1520 (O_1520,N_13877,N_13970);
nand UO_1521 (O_1521,N_14982,N_13939);
or UO_1522 (O_1522,N_14652,N_13699);
nand UO_1523 (O_1523,N_13995,N_14356);
nand UO_1524 (O_1524,N_14215,N_14708);
or UO_1525 (O_1525,N_13579,N_14261);
xnor UO_1526 (O_1526,N_13994,N_13707);
and UO_1527 (O_1527,N_13957,N_13950);
nand UO_1528 (O_1528,N_13822,N_14675);
nor UO_1529 (O_1529,N_13803,N_14879);
nor UO_1530 (O_1530,N_13537,N_14681);
or UO_1531 (O_1531,N_14745,N_14820);
xor UO_1532 (O_1532,N_14818,N_14340);
or UO_1533 (O_1533,N_14299,N_14269);
xor UO_1534 (O_1534,N_14560,N_14158);
nor UO_1535 (O_1535,N_14827,N_14884);
nor UO_1536 (O_1536,N_13985,N_14404);
nand UO_1537 (O_1537,N_14785,N_14406);
nor UO_1538 (O_1538,N_13638,N_14005);
nand UO_1539 (O_1539,N_13626,N_14041);
nor UO_1540 (O_1540,N_13684,N_13897);
nor UO_1541 (O_1541,N_14958,N_13811);
xor UO_1542 (O_1542,N_14176,N_13583);
or UO_1543 (O_1543,N_13589,N_13765);
xnor UO_1544 (O_1544,N_14124,N_13731);
nor UO_1545 (O_1545,N_13708,N_14250);
xnor UO_1546 (O_1546,N_13890,N_13906);
or UO_1547 (O_1547,N_13764,N_13536);
and UO_1548 (O_1548,N_13752,N_13541);
xor UO_1549 (O_1549,N_14996,N_14821);
and UO_1550 (O_1550,N_13687,N_14759);
or UO_1551 (O_1551,N_13729,N_13555);
or UO_1552 (O_1552,N_13962,N_14089);
xor UO_1553 (O_1553,N_13931,N_14798);
nor UO_1554 (O_1554,N_14248,N_14735);
and UO_1555 (O_1555,N_13827,N_14959);
or UO_1556 (O_1556,N_14106,N_14038);
or UO_1557 (O_1557,N_14367,N_14687);
nand UO_1558 (O_1558,N_13941,N_14259);
nand UO_1559 (O_1559,N_14383,N_14648);
nand UO_1560 (O_1560,N_13554,N_14022);
nand UO_1561 (O_1561,N_14810,N_13738);
or UO_1562 (O_1562,N_14545,N_14631);
xnor UO_1563 (O_1563,N_13921,N_13525);
nor UO_1564 (O_1564,N_14891,N_13772);
and UO_1565 (O_1565,N_14915,N_14224);
nand UO_1566 (O_1566,N_14313,N_14558);
nor UO_1567 (O_1567,N_14538,N_14158);
nand UO_1568 (O_1568,N_13774,N_14263);
nand UO_1569 (O_1569,N_14990,N_13870);
nand UO_1570 (O_1570,N_14616,N_13882);
and UO_1571 (O_1571,N_14949,N_14596);
and UO_1572 (O_1572,N_14756,N_14696);
xor UO_1573 (O_1573,N_14338,N_13723);
nand UO_1574 (O_1574,N_14276,N_14111);
nand UO_1575 (O_1575,N_14797,N_14321);
and UO_1576 (O_1576,N_13681,N_14168);
nand UO_1577 (O_1577,N_14189,N_14194);
and UO_1578 (O_1578,N_13658,N_14054);
nand UO_1579 (O_1579,N_13644,N_14861);
xor UO_1580 (O_1580,N_14885,N_13897);
nor UO_1581 (O_1581,N_14077,N_14522);
nand UO_1582 (O_1582,N_14403,N_14611);
xor UO_1583 (O_1583,N_13977,N_14800);
or UO_1584 (O_1584,N_14534,N_13514);
and UO_1585 (O_1585,N_14337,N_13945);
or UO_1586 (O_1586,N_14056,N_14456);
nor UO_1587 (O_1587,N_14826,N_14982);
nand UO_1588 (O_1588,N_14630,N_14925);
xnor UO_1589 (O_1589,N_14341,N_14009);
and UO_1590 (O_1590,N_14748,N_13791);
and UO_1591 (O_1591,N_13553,N_14204);
and UO_1592 (O_1592,N_14208,N_14470);
nor UO_1593 (O_1593,N_13973,N_13921);
nand UO_1594 (O_1594,N_14862,N_14053);
xnor UO_1595 (O_1595,N_14241,N_14120);
and UO_1596 (O_1596,N_14470,N_13988);
and UO_1597 (O_1597,N_13891,N_14921);
nor UO_1598 (O_1598,N_13977,N_14608);
and UO_1599 (O_1599,N_13675,N_14179);
or UO_1600 (O_1600,N_14184,N_14812);
and UO_1601 (O_1601,N_14102,N_13977);
nor UO_1602 (O_1602,N_14180,N_14475);
and UO_1603 (O_1603,N_13830,N_14121);
nor UO_1604 (O_1604,N_14795,N_14866);
nand UO_1605 (O_1605,N_13805,N_14842);
nand UO_1606 (O_1606,N_14467,N_14567);
or UO_1607 (O_1607,N_14583,N_14931);
nor UO_1608 (O_1608,N_14263,N_14716);
xnor UO_1609 (O_1609,N_13636,N_14092);
nand UO_1610 (O_1610,N_13897,N_14147);
nand UO_1611 (O_1611,N_14507,N_14902);
nor UO_1612 (O_1612,N_14327,N_14633);
nand UO_1613 (O_1613,N_14504,N_13763);
and UO_1614 (O_1614,N_14424,N_13694);
nand UO_1615 (O_1615,N_14019,N_13911);
nor UO_1616 (O_1616,N_13901,N_13542);
nor UO_1617 (O_1617,N_13574,N_13533);
nor UO_1618 (O_1618,N_14617,N_14501);
nor UO_1619 (O_1619,N_14144,N_14067);
or UO_1620 (O_1620,N_13543,N_14615);
nor UO_1621 (O_1621,N_13723,N_14890);
and UO_1622 (O_1622,N_13686,N_14265);
nand UO_1623 (O_1623,N_14874,N_14810);
nand UO_1624 (O_1624,N_14978,N_13891);
and UO_1625 (O_1625,N_14658,N_13861);
nor UO_1626 (O_1626,N_14193,N_14110);
or UO_1627 (O_1627,N_14843,N_14842);
and UO_1628 (O_1628,N_14181,N_14580);
or UO_1629 (O_1629,N_14513,N_13917);
or UO_1630 (O_1630,N_14879,N_14424);
xnor UO_1631 (O_1631,N_13656,N_14988);
and UO_1632 (O_1632,N_14270,N_14380);
and UO_1633 (O_1633,N_13509,N_13866);
or UO_1634 (O_1634,N_13736,N_14670);
and UO_1635 (O_1635,N_14889,N_13554);
nor UO_1636 (O_1636,N_13992,N_13585);
xor UO_1637 (O_1637,N_14267,N_13621);
xor UO_1638 (O_1638,N_13962,N_14133);
or UO_1639 (O_1639,N_14902,N_14256);
nand UO_1640 (O_1640,N_13605,N_14050);
nor UO_1641 (O_1641,N_13534,N_14754);
nand UO_1642 (O_1642,N_14148,N_14996);
nor UO_1643 (O_1643,N_14283,N_14188);
nor UO_1644 (O_1644,N_14072,N_14275);
nor UO_1645 (O_1645,N_14006,N_14846);
nor UO_1646 (O_1646,N_13801,N_13805);
nor UO_1647 (O_1647,N_13888,N_14242);
and UO_1648 (O_1648,N_14452,N_13684);
or UO_1649 (O_1649,N_14744,N_14675);
and UO_1650 (O_1650,N_14616,N_14649);
nand UO_1651 (O_1651,N_13638,N_14391);
nand UO_1652 (O_1652,N_14813,N_14345);
or UO_1653 (O_1653,N_14122,N_14712);
or UO_1654 (O_1654,N_14200,N_14039);
or UO_1655 (O_1655,N_14875,N_13700);
nor UO_1656 (O_1656,N_13982,N_13743);
xor UO_1657 (O_1657,N_14312,N_14685);
nor UO_1658 (O_1658,N_13900,N_14256);
nor UO_1659 (O_1659,N_13721,N_13612);
nand UO_1660 (O_1660,N_13774,N_13621);
or UO_1661 (O_1661,N_14482,N_13834);
or UO_1662 (O_1662,N_13799,N_14897);
xor UO_1663 (O_1663,N_13734,N_14736);
xor UO_1664 (O_1664,N_14881,N_13698);
nor UO_1665 (O_1665,N_14230,N_13568);
or UO_1666 (O_1666,N_13653,N_14435);
nor UO_1667 (O_1667,N_14473,N_13605);
nand UO_1668 (O_1668,N_14050,N_14879);
or UO_1669 (O_1669,N_14498,N_13691);
or UO_1670 (O_1670,N_14091,N_14979);
nand UO_1671 (O_1671,N_13517,N_14167);
xnor UO_1672 (O_1672,N_14330,N_13879);
nor UO_1673 (O_1673,N_13862,N_13978);
or UO_1674 (O_1674,N_14989,N_14307);
nor UO_1675 (O_1675,N_14338,N_14471);
xnor UO_1676 (O_1676,N_14323,N_14879);
nor UO_1677 (O_1677,N_14587,N_13871);
and UO_1678 (O_1678,N_14271,N_14788);
xnor UO_1679 (O_1679,N_14781,N_14576);
xnor UO_1680 (O_1680,N_14736,N_13918);
xnor UO_1681 (O_1681,N_14761,N_13968);
nand UO_1682 (O_1682,N_14664,N_14212);
nor UO_1683 (O_1683,N_14012,N_14500);
nor UO_1684 (O_1684,N_13784,N_13834);
nor UO_1685 (O_1685,N_14223,N_13578);
and UO_1686 (O_1686,N_14007,N_14674);
nor UO_1687 (O_1687,N_14610,N_14963);
and UO_1688 (O_1688,N_14040,N_14395);
xnor UO_1689 (O_1689,N_14127,N_13953);
and UO_1690 (O_1690,N_14685,N_14222);
nor UO_1691 (O_1691,N_14170,N_13907);
or UO_1692 (O_1692,N_14207,N_14398);
or UO_1693 (O_1693,N_13583,N_13634);
and UO_1694 (O_1694,N_14333,N_14614);
nand UO_1695 (O_1695,N_14214,N_13651);
nand UO_1696 (O_1696,N_14197,N_14401);
xor UO_1697 (O_1697,N_14025,N_14989);
xnor UO_1698 (O_1698,N_14024,N_14237);
nor UO_1699 (O_1699,N_14470,N_14313);
nor UO_1700 (O_1700,N_14504,N_13656);
xnor UO_1701 (O_1701,N_14825,N_13993);
xor UO_1702 (O_1702,N_14890,N_14798);
xor UO_1703 (O_1703,N_13520,N_13539);
xnor UO_1704 (O_1704,N_14792,N_13594);
and UO_1705 (O_1705,N_13921,N_14642);
xor UO_1706 (O_1706,N_14448,N_14605);
and UO_1707 (O_1707,N_14288,N_14821);
xor UO_1708 (O_1708,N_13599,N_14285);
or UO_1709 (O_1709,N_13961,N_14743);
xnor UO_1710 (O_1710,N_13992,N_14697);
nand UO_1711 (O_1711,N_13774,N_13672);
and UO_1712 (O_1712,N_13905,N_14841);
xnor UO_1713 (O_1713,N_14447,N_13760);
nor UO_1714 (O_1714,N_14234,N_13619);
and UO_1715 (O_1715,N_13590,N_14208);
nand UO_1716 (O_1716,N_13874,N_14630);
nor UO_1717 (O_1717,N_14334,N_13628);
xnor UO_1718 (O_1718,N_14775,N_14913);
xnor UO_1719 (O_1719,N_14240,N_13806);
or UO_1720 (O_1720,N_13733,N_13677);
or UO_1721 (O_1721,N_14936,N_14961);
nor UO_1722 (O_1722,N_14218,N_14291);
and UO_1723 (O_1723,N_13663,N_14846);
and UO_1724 (O_1724,N_13598,N_14620);
or UO_1725 (O_1725,N_13976,N_14103);
xnor UO_1726 (O_1726,N_14375,N_14325);
or UO_1727 (O_1727,N_13912,N_14962);
nor UO_1728 (O_1728,N_14638,N_13811);
xor UO_1729 (O_1729,N_14870,N_14569);
and UO_1730 (O_1730,N_13554,N_13576);
or UO_1731 (O_1731,N_14829,N_14069);
or UO_1732 (O_1732,N_14290,N_13952);
nand UO_1733 (O_1733,N_14443,N_14826);
nand UO_1734 (O_1734,N_14929,N_14426);
and UO_1735 (O_1735,N_14636,N_13758);
or UO_1736 (O_1736,N_13665,N_13602);
and UO_1737 (O_1737,N_14109,N_14241);
or UO_1738 (O_1738,N_14578,N_14217);
and UO_1739 (O_1739,N_13747,N_14164);
and UO_1740 (O_1740,N_14007,N_14394);
and UO_1741 (O_1741,N_14024,N_14634);
or UO_1742 (O_1742,N_13968,N_14587);
xnor UO_1743 (O_1743,N_14864,N_14891);
or UO_1744 (O_1744,N_13701,N_14629);
xnor UO_1745 (O_1745,N_14939,N_14961);
nand UO_1746 (O_1746,N_13648,N_14479);
and UO_1747 (O_1747,N_14523,N_13906);
nor UO_1748 (O_1748,N_14098,N_13756);
and UO_1749 (O_1749,N_14698,N_14193);
xor UO_1750 (O_1750,N_14675,N_14289);
xnor UO_1751 (O_1751,N_13743,N_14304);
or UO_1752 (O_1752,N_14070,N_13534);
and UO_1753 (O_1753,N_14453,N_13867);
nand UO_1754 (O_1754,N_13720,N_13816);
xor UO_1755 (O_1755,N_13872,N_13913);
or UO_1756 (O_1756,N_14973,N_14295);
nand UO_1757 (O_1757,N_13724,N_14033);
xnor UO_1758 (O_1758,N_14220,N_13758);
nand UO_1759 (O_1759,N_14537,N_13869);
nor UO_1760 (O_1760,N_14500,N_14104);
or UO_1761 (O_1761,N_14721,N_14450);
nand UO_1762 (O_1762,N_13909,N_14090);
nor UO_1763 (O_1763,N_14271,N_13549);
nand UO_1764 (O_1764,N_14933,N_14236);
nor UO_1765 (O_1765,N_14764,N_14010);
or UO_1766 (O_1766,N_14507,N_14600);
or UO_1767 (O_1767,N_13560,N_13516);
nor UO_1768 (O_1768,N_14044,N_13737);
or UO_1769 (O_1769,N_13969,N_13884);
or UO_1770 (O_1770,N_14335,N_13708);
nand UO_1771 (O_1771,N_14743,N_13623);
nand UO_1772 (O_1772,N_13523,N_14064);
nor UO_1773 (O_1773,N_14905,N_13693);
xnor UO_1774 (O_1774,N_14073,N_14567);
nand UO_1775 (O_1775,N_14087,N_14934);
xnor UO_1776 (O_1776,N_13551,N_13650);
nand UO_1777 (O_1777,N_14050,N_13989);
nor UO_1778 (O_1778,N_14930,N_14321);
nand UO_1779 (O_1779,N_14279,N_14716);
nor UO_1780 (O_1780,N_13988,N_14043);
nor UO_1781 (O_1781,N_14802,N_14094);
nand UO_1782 (O_1782,N_14895,N_13606);
and UO_1783 (O_1783,N_13646,N_14591);
or UO_1784 (O_1784,N_14349,N_14256);
nor UO_1785 (O_1785,N_13964,N_13924);
or UO_1786 (O_1786,N_14178,N_14727);
or UO_1787 (O_1787,N_14064,N_14597);
nand UO_1788 (O_1788,N_13964,N_14637);
xor UO_1789 (O_1789,N_14808,N_14648);
xor UO_1790 (O_1790,N_14503,N_14837);
xnor UO_1791 (O_1791,N_13866,N_13959);
nor UO_1792 (O_1792,N_14626,N_14512);
xor UO_1793 (O_1793,N_14592,N_14125);
xnor UO_1794 (O_1794,N_14215,N_14767);
or UO_1795 (O_1795,N_14214,N_14393);
nand UO_1796 (O_1796,N_14662,N_14099);
and UO_1797 (O_1797,N_13731,N_14405);
nand UO_1798 (O_1798,N_14867,N_14740);
xnor UO_1799 (O_1799,N_13735,N_13533);
nand UO_1800 (O_1800,N_13538,N_14372);
nand UO_1801 (O_1801,N_14221,N_13500);
nor UO_1802 (O_1802,N_14130,N_14181);
nor UO_1803 (O_1803,N_14294,N_13945);
nor UO_1804 (O_1804,N_14480,N_14228);
and UO_1805 (O_1805,N_14384,N_14987);
and UO_1806 (O_1806,N_13993,N_13686);
nor UO_1807 (O_1807,N_13535,N_13736);
and UO_1808 (O_1808,N_14551,N_13958);
nand UO_1809 (O_1809,N_14617,N_13545);
nand UO_1810 (O_1810,N_13914,N_14324);
nand UO_1811 (O_1811,N_14871,N_13703);
and UO_1812 (O_1812,N_13662,N_13770);
nand UO_1813 (O_1813,N_14431,N_13850);
or UO_1814 (O_1814,N_14366,N_13721);
xnor UO_1815 (O_1815,N_14651,N_14786);
nor UO_1816 (O_1816,N_14922,N_14887);
nor UO_1817 (O_1817,N_13681,N_14877);
xnor UO_1818 (O_1818,N_14480,N_14920);
nor UO_1819 (O_1819,N_14170,N_13714);
xor UO_1820 (O_1820,N_14913,N_13799);
xnor UO_1821 (O_1821,N_14878,N_14218);
xnor UO_1822 (O_1822,N_13547,N_14568);
xor UO_1823 (O_1823,N_14356,N_13822);
xnor UO_1824 (O_1824,N_14276,N_14972);
nand UO_1825 (O_1825,N_14204,N_14127);
xnor UO_1826 (O_1826,N_13942,N_13699);
and UO_1827 (O_1827,N_13517,N_14446);
nand UO_1828 (O_1828,N_14217,N_13629);
or UO_1829 (O_1829,N_13726,N_13902);
xnor UO_1830 (O_1830,N_14562,N_14095);
nand UO_1831 (O_1831,N_13779,N_13959);
xnor UO_1832 (O_1832,N_14937,N_13887);
xor UO_1833 (O_1833,N_13639,N_14708);
nand UO_1834 (O_1834,N_14854,N_14502);
nand UO_1835 (O_1835,N_14923,N_14013);
or UO_1836 (O_1836,N_14699,N_14741);
xnor UO_1837 (O_1837,N_14812,N_13648);
or UO_1838 (O_1838,N_13892,N_13510);
xor UO_1839 (O_1839,N_14730,N_13504);
xnor UO_1840 (O_1840,N_13549,N_14403);
nor UO_1841 (O_1841,N_14685,N_14809);
nor UO_1842 (O_1842,N_13645,N_13868);
nand UO_1843 (O_1843,N_14584,N_13816);
and UO_1844 (O_1844,N_13761,N_14055);
or UO_1845 (O_1845,N_13849,N_14594);
nand UO_1846 (O_1846,N_14401,N_14939);
nor UO_1847 (O_1847,N_13661,N_14938);
nand UO_1848 (O_1848,N_13851,N_14724);
or UO_1849 (O_1849,N_14968,N_14587);
xnor UO_1850 (O_1850,N_14703,N_14214);
or UO_1851 (O_1851,N_14517,N_13948);
xor UO_1852 (O_1852,N_13640,N_14504);
xnor UO_1853 (O_1853,N_13788,N_14972);
nor UO_1854 (O_1854,N_14631,N_13541);
nand UO_1855 (O_1855,N_14134,N_13756);
or UO_1856 (O_1856,N_13500,N_14300);
xor UO_1857 (O_1857,N_14330,N_14474);
or UO_1858 (O_1858,N_14887,N_14929);
nor UO_1859 (O_1859,N_14658,N_14851);
xor UO_1860 (O_1860,N_13638,N_14578);
and UO_1861 (O_1861,N_14016,N_14004);
xor UO_1862 (O_1862,N_14553,N_14933);
nor UO_1863 (O_1863,N_14691,N_13854);
nand UO_1864 (O_1864,N_14733,N_13556);
and UO_1865 (O_1865,N_13872,N_14889);
xnor UO_1866 (O_1866,N_14517,N_14098);
and UO_1867 (O_1867,N_13673,N_14718);
or UO_1868 (O_1868,N_14815,N_13685);
or UO_1869 (O_1869,N_14341,N_14822);
and UO_1870 (O_1870,N_13962,N_13756);
nand UO_1871 (O_1871,N_14474,N_13874);
and UO_1872 (O_1872,N_14879,N_14517);
nand UO_1873 (O_1873,N_14979,N_13937);
or UO_1874 (O_1874,N_13554,N_14449);
xnor UO_1875 (O_1875,N_13754,N_13564);
nand UO_1876 (O_1876,N_14315,N_13622);
nand UO_1877 (O_1877,N_13711,N_14177);
nor UO_1878 (O_1878,N_14571,N_13716);
and UO_1879 (O_1879,N_14380,N_14485);
or UO_1880 (O_1880,N_14581,N_14602);
nor UO_1881 (O_1881,N_13721,N_14256);
and UO_1882 (O_1882,N_14001,N_14654);
xnor UO_1883 (O_1883,N_13884,N_14249);
nand UO_1884 (O_1884,N_14099,N_13731);
nor UO_1885 (O_1885,N_14628,N_14861);
or UO_1886 (O_1886,N_14119,N_13565);
nor UO_1887 (O_1887,N_13858,N_13881);
nor UO_1888 (O_1888,N_14151,N_14749);
nand UO_1889 (O_1889,N_14585,N_14134);
xnor UO_1890 (O_1890,N_14129,N_14999);
xnor UO_1891 (O_1891,N_13943,N_13586);
xor UO_1892 (O_1892,N_14813,N_14265);
and UO_1893 (O_1893,N_14425,N_13790);
or UO_1894 (O_1894,N_14120,N_13849);
nor UO_1895 (O_1895,N_14157,N_13676);
nand UO_1896 (O_1896,N_13840,N_14281);
nand UO_1897 (O_1897,N_14321,N_13804);
xor UO_1898 (O_1898,N_13555,N_14013);
or UO_1899 (O_1899,N_14446,N_14380);
or UO_1900 (O_1900,N_14319,N_13873);
and UO_1901 (O_1901,N_14700,N_13938);
nor UO_1902 (O_1902,N_14893,N_13759);
nor UO_1903 (O_1903,N_13647,N_14866);
nor UO_1904 (O_1904,N_14118,N_13857);
xnor UO_1905 (O_1905,N_14813,N_14454);
or UO_1906 (O_1906,N_14406,N_13869);
xor UO_1907 (O_1907,N_14635,N_14208);
and UO_1908 (O_1908,N_14280,N_14177);
nor UO_1909 (O_1909,N_14634,N_13750);
and UO_1910 (O_1910,N_14062,N_13897);
xnor UO_1911 (O_1911,N_14479,N_13963);
or UO_1912 (O_1912,N_14909,N_14972);
and UO_1913 (O_1913,N_13800,N_14800);
nor UO_1914 (O_1914,N_13505,N_14993);
and UO_1915 (O_1915,N_14603,N_14101);
nor UO_1916 (O_1916,N_14337,N_13602);
nor UO_1917 (O_1917,N_13953,N_14314);
nor UO_1918 (O_1918,N_14339,N_14779);
xnor UO_1919 (O_1919,N_14453,N_14296);
and UO_1920 (O_1920,N_14206,N_14441);
or UO_1921 (O_1921,N_14490,N_14948);
or UO_1922 (O_1922,N_14021,N_14035);
or UO_1923 (O_1923,N_13591,N_14112);
nor UO_1924 (O_1924,N_13989,N_13688);
nor UO_1925 (O_1925,N_14492,N_14776);
nor UO_1926 (O_1926,N_14109,N_14373);
xor UO_1927 (O_1927,N_14661,N_13502);
nand UO_1928 (O_1928,N_14687,N_14010);
or UO_1929 (O_1929,N_14165,N_14639);
nand UO_1930 (O_1930,N_13689,N_14102);
or UO_1931 (O_1931,N_14969,N_13961);
nand UO_1932 (O_1932,N_14610,N_14946);
nor UO_1933 (O_1933,N_13805,N_14020);
and UO_1934 (O_1934,N_13909,N_14652);
and UO_1935 (O_1935,N_13535,N_14356);
or UO_1936 (O_1936,N_14270,N_13785);
xnor UO_1937 (O_1937,N_14030,N_14544);
nor UO_1938 (O_1938,N_14522,N_14205);
and UO_1939 (O_1939,N_14559,N_14255);
xor UO_1940 (O_1940,N_14795,N_14225);
and UO_1941 (O_1941,N_14152,N_14479);
xnor UO_1942 (O_1942,N_13752,N_14779);
nor UO_1943 (O_1943,N_13770,N_14581);
nand UO_1944 (O_1944,N_14008,N_14932);
xnor UO_1945 (O_1945,N_14485,N_14933);
nor UO_1946 (O_1946,N_14689,N_13866);
nor UO_1947 (O_1947,N_14766,N_14128);
or UO_1948 (O_1948,N_13784,N_14028);
nor UO_1949 (O_1949,N_14594,N_14501);
xnor UO_1950 (O_1950,N_13603,N_13752);
nand UO_1951 (O_1951,N_14421,N_14396);
nand UO_1952 (O_1952,N_14452,N_14775);
and UO_1953 (O_1953,N_14102,N_14833);
or UO_1954 (O_1954,N_13823,N_14483);
and UO_1955 (O_1955,N_14366,N_14812);
and UO_1956 (O_1956,N_13559,N_13853);
nor UO_1957 (O_1957,N_14710,N_14922);
nor UO_1958 (O_1958,N_14074,N_14977);
and UO_1959 (O_1959,N_13571,N_14342);
xor UO_1960 (O_1960,N_14541,N_14582);
nor UO_1961 (O_1961,N_14738,N_14632);
nor UO_1962 (O_1962,N_13501,N_13890);
nand UO_1963 (O_1963,N_13857,N_14770);
xor UO_1964 (O_1964,N_14011,N_14599);
or UO_1965 (O_1965,N_14686,N_13904);
or UO_1966 (O_1966,N_14830,N_13654);
or UO_1967 (O_1967,N_13919,N_14796);
nor UO_1968 (O_1968,N_13949,N_14001);
xor UO_1969 (O_1969,N_14280,N_14345);
nor UO_1970 (O_1970,N_14366,N_13648);
nor UO_1971 (O_1971,N_13540,N_14179);
nor UO_1972 (O_1972,N_14810,N_13786);
and UO_1973 (O_1973,N_13663,N_14759);
or UO_1974 (O_1974,N_14497,N_14421);
and UO_1975 (O_1975,N_14929,N_14324);
nand UO_1976 (O_1976,N_14435,N_14967);
or UO_1977 (O_1977,N_14177,N_13588);
nand UO_1978 (O_1978,N_14390,N_14204);
and UO_1979 (O_1979,N_14683,N_14488);
xor UO_1980 (O_1980,N_14741,N_14498);
nand UO_1981 (O_1981,N_14366,N_14162);
or UO_1982 (O_1982,N_13500,N_13905);
and UO_1983 (O_1983,N_14502,N_14377);
or UO_1984 (O_1984,N_14729,N_13694);
nor UO_1985 (O_1985,N_13970,N_14386);
xnor UO_1986 (O_1986,N_14331,N_13605);
xnor UO_1987 (O_1987,N_14162,N_13956);
nand UO_1988 (O_1988,N_13911,N_14684);
nor UO_1989 (O_1989,N_14289,N_13873);
or UO_1990 (O_1990,N_14035,N_14435);
xnor UO_1991 (O_1991,N_14609,N_14281);
xnor UO_1992 (O_1992,N_13642,N_13711);
and UO_1993 (O_1993,N_14922,N_13898);
and UO_1994 (O_1994,N_14917,N_14095);
and UO_1995 (O_1995,N_14272,N_14019);
and UO_1996 (O_1996,N_14211,N_13582);
or UO_1997 (O_1997,N_14061,N_13674);
nand UO_1998 (O_1998,N_13660,N_14143);
nor UO_1999 (O_1999,N_14913,N_14029);
endmodule