module basic_1000_10000_1500_10_levels_2xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_384,In_216);
and U1 (N_1,In_786,In_112);
nor U2 (N_2,In_813,In_388);
and U3 (N_3,In_962,In_445);
or U4 (N_4,In_219,In_98);
and U5 (N_5,In_363,In_976);
and U6 (N_6,In_983,In_979);
nor U7 (N_7,In_119,In_614);
nand U8 (N_8,In_929,In_196);
and U9 (N_9,In_140,In_186);
and U10 (N_10,In_887,In_184);
or U11 (N_11,In_59,In_755);
and U12 (N_12,In_980,In_779);
or U13 (N_13,In_453,In_471);
or U14 (N_14,In_440,In_348);
and U15 (N_15,In_68,In_482);
or U16 (N_16,In_278,In_139);
and U17 (N_17,In_798,In_920);
and U18 (N_18,In_439,In_560);
and U19 (N_19,In_431,In_276);
or U20 (N_20,In_829,In_86);
nor U21 (N_21,In_896,In_650);
nor U22 (N_22,In_517,In_352);
xnor U23 (N_23,In_11,In_7);
or U24 (N_24,In_447,In_579);
and U25 (N_25,In_691,In_961);
nor U26 (N_26,In_587,In_902);
and U27 (N_27,In_940,In_475);
nor U28 (N_28,In_401,In_291);
nand U29 (N_29,In_75,In_48);
or U30 (N_30,In_154,In_690);
or U31 (N_31,In_429,In_378);
and U32 (N_32,In_875,In_558);
and U33 (N_33,In_211,In_677);
nor U34 (N_34,In_524,In_738);
nand U35 (N_35,In_808,In_342);
or U36 (N_36,In_965,In_823);
nand U37 (N_37,In_726,In_545);
or U38 (N_38,In_703,In_927);
nand U39 (N_39,In_52,In_575);
nand U40 (N_40,In_424,In_547);
or U41 (N_41,In_187,In_623);
nor U42 (N_42,In_529,In_830);
and U43 (N_43,In_303,In_485);
nor U44 (N_44,In_245,In_478);
nand U45 (N_45,In_47,In_644);
xor U46 (N_46,In_737,In_207);
and U47 (N_47,In_130,In_676);
or U48 (N_48,In_132,In_73);
nand U49 (N_49,In_850,In_831);
or U50 (N_50,In_402,In_859);
or U51 (N_51,In_700,In_995);
or U52 (N_52,In_491,In_170);
and U53 (N_53,In_665,In_598);
or U54 (N_54,In_915,In_495);
nand U55 (N_55,In_936,In_244);
or U56 (N_56,In_425,In_323);
or U57 (N_57,In_203,In_717);
nor U58 (N_58,In_627,In_556);
nor U59 (N_59,In_56,In_241);
and U60 (N_60,In_339,In_963);
or U61 (N_61,In_29,In_230);
and U62 (N_62,In_981,In_660);
nand U63 (N_63,In_883,In_543);
nor U64 (N_64,In_499,In_415);
nand U65 (N_65,In_654,In_254);
nor U66 (N_66,In_778,In_437);
or U67 (N_67,In_996,In_133);
and U68 (N_68,In_810,In_948);
and U69 (N_69,In_100,In_262);
and U70 (N_70,In_149,In_533);
nand U71 (N_71,In_32,In_316);
nand U72 (N_72,In_854,In_643);
and U73 (N_73,In_422,In_457);
nor U74 (N_74,In_452,In_742);
nor U75 (N_75,In_341,In_209);
nand U76 (N_76,In_76,In_777);
nor U77 (N_77,In_521,In_874);
nand U78 (N_78,In_226,In_34);
nand U79 (N_79,In_672,In_725);
or U80 (N_80,In_403,In_821);
nand U81 (N_81,In_550,In_651);
nand U82 (N_82,In_53,In_85);
or U83 (N_83,In_351,In_731);
or U84 (N_84,In_639,In_173);
nand U85 (N_85,In_855,In_836);
nor U86 (N_86,In_732,In_398);
or U87 (N_87,In_774,In_256);
and U88 (N_88,In_669,In_884);
nor U89 (N_89,In_120,In_467);
and U90 (N_90,In_880,In_835);
nor U91 (N_91,In_990,In_271);
and U92 (N_92,In_364,In_325);
or U93 (N_93,In_506,In_583);
nor U94 (N_94,In_395,In_773);
nor U95 (N_95,In_251,In_122);
or U96 (N_96,In_159,In_194);
nor U97 (N_97,In_542,In_421);
nand U98 (N_98,In_15,In_18);
or U99 (N_99,In_621,In_839);
and U100 (N_100,In_765,In_304);
nand U101 (N_101,In_716,In_527);
nor U102 (N_102,In_416,In_818);
or U103 (N_103,In_531,In_90);
nor U104 (N_104,In_695,In_247);
nor U105 (N_105,In_966,In_852);
nand U106 (N_106,In_292,In_815);
nor U107 (N_107,In_36,In_740);
or U108 (N_108,In_268,In_572);
or U109 (N_109,In_432,In_985);
nand U110 (N_110,In_620,In_897);
or U111 (N_111,In_608,In_78);
nor U112 (N_112,In_868,In_195);
and U113 (N_113,In_81,In_862);
nor U114 (N_114,In_169,In_313);
and U115 (N_115,In_782,In_6);
nor U116 (N_116,In_356,In_640);
nor U117 (N_117,In_763,In_306);
nor U118 (N_118,In_466,In_309);
nand U119 (N_119,In_381,In_320);
nand U120 (N_120,In_204,In_589);
nor U121 (N_121,In_557,In_576);
and U122 (N_122,In_391,In_92);
nand U123 (N_123,In_396,In_511);
nand U124 (N_124,In_879,In_997);
nor U125 (N_125,In_191,In_900);
nand U126 (N_126,In_565,In_793);
or U127 (N_127,In_799,In_780);
nor U128 (N_128,In_71,In_332);
or U129 (N_129,In_246,In_270);
nand U130 (N_130,In_790,In_175);
and U131 (N_131,In_947,In_824);
or U132 (N_132,In_4,In_967);
or U133 (N_133,In_188,In_597);
or U134 (N_134,In_974,In_519);
or U135 (N_135,In_603,In_260);
nor U136 (N_136,In_580,In_141);
and U137 (N_137,In_117,In_619);
nor U138 (N_138,In_370,In_911);
nor U139 (N_139,In_328,In_959);
nand U140 (N_140,In_462,In_872);
nor U141 (N_141,In_968,In_711);
nor U142 (N_142,In_893,In_93);
or U143 (N_143,In_470,In_702);
or U144 (N_144,In_393,In_661);
and U145 (N_145,In_420,In_759);
nor U146 (N_146,In_588,In_157);
nor U147 (N_147,In_944,In_26);
nor U148 (N_148,In_680,In_493);
and U149 (N_149,In_77,In_39);
nor U150 (N_150,In_827,In_108);
and U151 (N_151,In_97,In_455);
and U152 (N_152,In_789,In_595);
and U153 (N_153,In_227,In_986);
nor U154 (N_154,In_888,In_656);
and U155 (N_155,In_657,In_744);
nand U156 (N_156,In_435,In_111);
and U157 (N_157,In_544,In_9);
nand U158 (N_158,In_358,In_655);
nand U159 (N_159,In_300,In_606);
nor U160 (N_160,In_616,In_752);
nor U161 (N_161,In_630,In_183);
nor U162 (N_162,In_571,In_528);
or U163 (N_163,In_999,In_177);
nand U164 (N_164,In_973,In_2);
nor U165 (N_165,In_72,In_379);
and U166 (N_166,In_809,In_367);
or U167 (N_167,In_89,In_269);
nor U168 (N_168,In_324,In_197);
nand U169 (N_169,In_266,In_678);
or U170 (N_170,In_486,In_327);
or U171 (N_171,In_553,In_123);
and U172 (N_172,In_301,In_891);
and U173 (N_173,In_689,In_95);
or U174 (N_174,In_819,In_163);
and U175 (N_175,In_618,In_280);
nor U176 (N_176,In_182,In_24);
nand U177 (N_177,In_581,In_231);
nand U178 (N_178,In_613,In_50);
nor U179 (N_179,In_66,In_954);
or U180 (N_180,In_131,In_795);
nor U181 (N_181,In_205,In_242);
or U182 (N_182,In_258,In_769);
and U183 (N_183,In_624,In_237);
xnor U184 (N_184,In_135,In_642);
or U185 (N_185,In_265,In_629);
and U186 (N_186,In_277,In_261);
and U187 (N_187,In_514,In_788);
and U188 (N_188,In_0,In_42);
and U189 (N_189,In_259,In_10);
nor U190 (N_190,In_382,In_480);
or U191 (N_191,In_797,In_666);
or U192 (N_192,In_894,In_38);
nor U193 (N_193,In_935,In_670);
and U194 (N_194,In_941,In_710);
nor U195 (N_195,In_632,In_586);
or U196 (N_196,In_377,In_17);
nor U197 (N_197,In_413,In_733);
nand U198 (N_198,In_611,In_713);
nor U199 (N_199,In_361,In_791);
nor U200 (N_200,In_189,In_870);
xnor U201 (N_201,In_57,In_847);
nor U202 (N_202,In_950,In_848);
nor U203 (N_203,In_257,In_501);
or U204 (N_204,In_709,In_563);
nand U205 (N_205,In_373,In_27);
nand U206 (N_206,In_648,In_473);
xnor U207 (N_207,In_520,In_522);
nand U208 (N_208,In_932,In_489);
and U209 (N_209,In_80,In_193);
nor U210 (N_210,In_876,In_87);
nor U211 (N_211,In_409,In_505);
and U212 (N_212,In_23,In_882);
and U213 (N_213,In_321,In_807);
nand U214 (N_214,In_688,In_28);
and U215 (N_215,In_659,In_83);
and U216 (N_216,In_767,In_114);
and U217 (N_217,In_390,In_155);
or U218 (N_218,In_172,In_362);
and U219 (N_219,In_804,In_792);
nand U220 (N_220,In_610,In_296);
nand U221 (N_221,In_698,In_199);
or U222 (N_222,In_989,In_994);
and U223 (N_223,In_366,In_863);
or U224 (N_224,In_430,In_267);
nor U225 (N_225,In_147,In_113);
nand U226 (N_226,In_949,In_25);
nor U227 (N_227,In_443,In_224);
xnor U228 (N_228,In_392,In_434);
nand U229 (N_229,In_910,In_41);
nor U230 (N_230,In_164,In_336);
nor U231 (N_231,In_118,In_760);
nand U232 (N_232,In_568,In_771);
and U233 (N_233,In_58,In_903);
and U234 (N_234,In_410,In_222);
or U235 (N_235,In_512,In_518);
nand U236 (N_236,In_213,In_889);
or U237 (N_237,In_161,In_107);
nor U238 (N_238,In_368,In_743);
and U239 (N_239,In_972,In_969);
nor U240 (N_240,In_405,In_555);
and U241 (N_241,In_160,In_3);
or U242 (N_242,In_308,In_638);
and U243 (N_243,In_404,In_153);
and U244 (N_244,In_922,In_525);
and U245 (N_245,In_833,In_615);
nor U246 (N_246,In_333,In_919);
nor U247 (N_247,In_585,In_634);
nor U248 (N_248,In_134,In_238);
and U249 (N_249,In_145,In_886);
nand U250 (N_250,In_757,In_201);
nor U251 (N_251,In_747,In_722);
nor U252 (N_252,In_718,In_838);
and U253 (N_253,In_837,In_803);
nand U254 (N_254,In_549,In_626);
nand U255 (N_255,In_465,In_817);
nor U256 (N_256,In_275,In_329);
and U257 (N_257,In_14,In_653);
nor U258 (N_258,In_820,In_538);
nor U259 (N_259,In_551,In_449);
and U260 (N_260,In_720,In_347);
and U261 (N_261,In_335,In_696);
nor U262 (N_262,In_484,In_451);
and U263 (N_263,In_930,In_785);
nand U264 (N_264,In_925,In_192);
or U265 (N_265,In_843,In_735);
nor U266 (N_266,In_554,In_287);
nor U267 (N_267,In_281,In_592);
or U268 (N_268,In_487,In_234);
nand U269 (N_269,In_548,In_91);
or U270 (N_270,In_856,In_124);
nand U271 (N_271,In_857,In_539);
nand U272 (N_272,In_593,In_16);
nand U273 (N_273,In_507,In_878);
or U274 (N_274,In_776,In_450);
nand U275 (N_275,In_63,In_552);
nand U276 (N_276,In_464,In_494);
nand U277 (N_277,In_236,In_781);
or U278 (N_278,In_784,In_129);
nor U279 (N_279,In_998,In_322);
and U280 (N_280,In_562,In_476);
or U281 (N_281,In_21,In_165);
or U282 (N_282,In_283,In_754);
and U283 (N_283,In_683,In_783);
nor U284 (N_284,In_217,In_513);
or U285 (N_285,In_284,In_775);
or U286 (N_286,In_143,In_383);
or U287 (N_287,In_993,In_750);
or U288 (N_288,In_753,In_858);
nand U289 (N_289,In_933,In_208);
or U290 (N_290,In_516,In_946);
or U291 (N_291,In_806,In_293);
nand U292 (N_292,In_70,In_628);
or U293 (N_293,In_210,In_496);
and U294 (N_294,In_45,In_302);
or U295 (N_295,In_274,In_12);
nand U296 (N_296,In_667,In_715);
nand U297 (N_297,In_956,In_248);
nand U298 (N_298,In_570,In_55);
or U299 (N_299,In_729,In_745);
and U300 (N_300,In_637,In_851);
and U301 (N_301,In_357,In_37);
nor U302 (N_302,In_125,In_811);
nand U303 (N_303,In_805,In_61);
and U304 (N_304,In_239,In_479);
nand U305 (N_305,In_477,In_960);
nand U306 (N_306,In_906,In_96);
nand U307 (N_307,In_330,In_582);
or U308 (N_308,In_504,In_739);
nor U309 (N_309,In_685,In_901);
and U310 (N_310,In_79,In_290);
nor U311 (N_311,In_43,In_371);
nor U312 (N_312,In_841,In_353);
or U313 (N_313,In_179,In_701);
or U314 (N_314,In_346,In_181);
or U315 (N_315,In_905,In_913);
or U316 (N_316,In_397,In_109);
nor U317 (N_317,In_842,In_127);
or U318 (N_318,In_67,In_982);
or U319 (N_319,In_115,In_853);
and U320 (N_320,In_223,In_699);
or U321 (N_321,In_594,In_250);
nor U322 (N_322,In_584,In_899);
or U323 (N_323,In_386,In_546);
and U324 (N_324,In_567,In_908);
and U325 (N_325,In_106,In_446);
xor U326 (N_326,In_310,In_212);
or U327 (N_327,In_746,In_380);
nor U328 (N_328,In_564,In_158);
or U329 (N_329,In_49,In_350);
nor U330 (N_330,In_51,In_975);
and U331 (N_331,In_220,In_800);
or U332 (N_332,In_943,In_895);
or U333 (N_333,In_168,In_607);
nand U334 (N_334,In_456,In_64);
nand U335 (N_335,In_62,In_65);
nand U336 (N_336,In_142,In_633);
nand U337 (N_337,In_958,In_426);
and U338 (N_338,In_240,In_376);
and U339 (N_339,In_54,In_225);
and U340 (N_340,In_536,In_751);
or U341 (N_341,In_375,In_869);
and U342 (N_342,In_991,In_162);
and U343 (N_343,In_60,In_705);
and U344 (N_344,In_218,In_574);
xor U345 (N_345,In_772,In_178);
and U346 (N_346,In_916,In_82);
or U347 (N_347,In_591,In_299);
nand U348 (N_348,In_652,In_305);
nor U349 (N_349,In_679,In_126);
nand U350 (N_350,In_812,In_235);
or U351 (N_351,In_232,In_768);
nor U352 (N_352,In_939,In_461);
nor U353 (N_353,In_200,In_964);
and U354 (N_354,In_474,In_714);
and U355 (N_355,In_706,In_334);
nor U356 (N_356,In_697,In_796);
and U357 (N_357,In_249,In_861);
nor U358 (N_358,In_904,In_828);
nand U359 (N_359,In_566,In_442);
nand U360 (N_360,In_414,In_617);
and U361 (N_361,In_692,In_344);
or U362 (N_362,In_596,In_873);
nand U363 (N_363,In_631,In_885);
nor U364 (N_364,In_734,In_138);
nor U365 (N_365,In_448,In_770);
or U366 (N_366,In_612,In_826);
nor U367 (N_367,In_472,In_730);
nand U368 (N_368,In_417,In_801);
nand U369 (N_369,In_992,In_712);
and U370 (N_370,In_693,In_559);
nand U371 (N_371,In_340,In_40);
or U372 (N_372,In_490,In_736);
nor U373 (N_373,In_326,In_840);
nand U374 (N_374,In_288,In_116);
and U375 (N_375,In_105,In_233);
or U376 (N_376,In_69,In_272);
and U377 (N_377,In_816,In_311);
and U378 (N_378,In_454,In_337);
and U379 (N_379,In_762,In_314);
and U380 (N_380,In_822,In_469);
and U381 (N_381,In_399,In_599);
nor U382 (N_382,In_682,In_412);
nor U383 (N_383,In_206,In_372);
nand U384 (N_384,In_909,In_881);
nand U385 (N_385,In_924,In_704);
and U386 (N_386,In_898,In_331);
or U387 (N_387,In_934,In_914);
or U388 (N_388,In_46,In_957);
and U389 (N_389,In_917,In_988);
xor U390 (N_390,In_307,In_243);
and U391 (N_391,In_190,In_128);
nor U392 (N_392,In_317,In_625);
and U393 (N_393,In_294,In_526);
or U394 (N_394,In_406,In_719);
and U395 (N_395,In_360,In_864);
xnor U396 (N_396,In_646,In_955);
nand U397 (N_397,In_389,In_318);
and U398 (N_398,In_13,In_601);
or U399 (N_399,In_561,In_166);
and U400 (N_400,In_675,In_31);
or U401 (N_401,In_577,In_94);
or U402 (N_402,In_255,In_681);
nand U403 (N_403,In_540,In_912);
and U404 (N_404,In_860,In_541);
nand U405 (N_405,In_844,In_723);
and U406 (N_406,In_724,In_156);
or U407 (N_407,In_359,In_867);
nor U408 (N_408,In_508,In_264);
nor U409 (N_409,In_228,In_374);
or U410 (N_410,In_263,In_515);
nor U411 (N_411,In_534,In_411);
nor U412 (N_412,In_99,In_460);
nor U413 (N_413,In_537,In_33);
or U414 (N_414,In_152,In_459);
nand U415 (N_415,In_952,In_741);
or U416 (N_416,In_252,In_987);
nor U417 (N_417,In_794,In_662);
and U418 (N_418,In_766,In_673);
nor U419 (N_419,In_418,In_756);
nor U420 (N_420,In_185,In_892);
or U421 (N_421,In_215,In_102);
nand U422 (N_422,In_761,In_458);
nor U423 (N_423,In_167,In_953);
nor U424 (N_424,In_708,In_214);
nand U425 (N_425,In_877,In_136);
nand U426 (N_426,In_385,In_202);
or U427 (N_427,In_144,In_748);
xor U428 (N_428,In_503,In_951);
or U429 (N_429,In_918,In_419);
nand U430 (N_430,In_428,In_174);
and U431 (N_431,In_88,In_289);
and U432 (N_432,In_942,In_338);
and U433 (N_433,In_221,In_137);
and U434 (N_434,In_635,In_871);
and U435 (N_435,In_408,In_970);
nor U436 (N_436,In_35,In_834);
or U437 (N_437,In_315,In_279);
nand U438 (N_438,In_436,In_604);
or U439 (N_439,In_500,In_727);
nand U440 (N_440,In_394,In_121);
and U441 (N_441,In_441,In_647);
nor U442 (N_442,In_369,In_707);
or U443 (N_443,In_721,In_602);
or U444 (N_444,In_645,In_104);
or U445 (N_445,In_802,In_764);
nand U446 (N_446,In_229,In_671);
and U447 (N_447,In_907,In_433);
nor U448 (N_448,In_664,In_787);
nor U449 (N_449,In_605,In_674);
nand U450 (N_450,In_971,In_663);
or U451 (N_451,In_573,In_814);
and U452 (N_452,In_407,In_928);
and U453 (N_453,In_728,In_641);
nand U454 (N_454,In_365,In_686);
nor U455 (N_455,In_319,In_444);
nand U456 (N_456,In_483,In_285);
or U457 (N_457,In_658,In_845);
nand U458 (N_458,In_355,In_502);
nand U459 (N_459,In_253,In_866);
xor U460 (N_460,In_44,In_150);
and U461 (N_461,In_535,In_622);
or U462 (N_462,In_481,In_832);
nor U463 (N_463,In_20,In_569);
nor U464 (N_464,In_668,In_74);
nand U465 (N_465,In_497,In_926);
or U466 (N_466,In_694,In_921);
or U467 (N_467,In_492,In_427);
and U468 (N_468,In_890,In_488);
and U469 (N_469,In_937,In_176);
and U470 (N_470,In_5,In_298);
or U471 (N_471,In_354,In_345);
nor U472 (N_472,In_343,In_423);
nor U473 (N_473,In_295,In_825);
nand U474 (N_474,In_101,In_600);
and U475 (N_475,In_19,In_636);
nand U476 (N_476,In_1,In_180);
or U477 (N_477,In_312,In_687);
or U478 (N_478,In_923,In_578);
nor U479 (N_479,In_977,In_684);
nor U480 (N_480,In_498,In_286);
nand U481 (N_481,In_30,In_273);
and U482 (N_482,In_171,In_400);
or U483 (N_483,In_931,In_297);
nand U484 (N_484,In_387,In_349);
nand U485 (N_485,In_945,In_282);
and U486 (N_486,In_8,In_749);
and U487 (N_487,In_110,In_530);
nor U488 (N_488,In_849,In_84);
nand U489 (N_489,In_148,In_865);
and U490 (N_490,In_438,In_758);
or U491 (N_491,In_984,In_532);
nor U492 (N_492,In_649,In_510);
nand U493 (N_493,In_938,In_523);
or U494 (N_494,In_978,In_198);
nand U495 (N_495,In_590,In_468);
or U496 (N_496,In_151,In_103);
and U497 (N_497,In_463,In_509);
and U498 (N_498,In_146,In_846);
nand U499 (N_499,In_609,In_22);
nor U500 (N_500,In_164,In_498);
nand U501 (N_501,In_101,In_888);
nand U502 (N_502,In_376,In_288);
and U503 (N_503,In_671,In_472);
or U504 (N_504,In_201,In_615);
nor U505 (N_505,In_509,In_444);
or U506 (N_506,In_359,In_956);
or U507 (N_507,In_245,In_827);
nand U508 (N_508,In_479,In_735);
or U509 (N_509,In_439,In_698);
and U510 (N_510,In_756,In_917);
and U511 (N_511,In_327,In_289);
nand U512 (N_512,In_735,In_631);
nor U513 (N_513,In_883,In_228);
nand U514 (N_514,In_142,In_219);
or U515 (N_515,In_816,In_271);
and U516 (N_516,In_945,In_936);
nand U517 (N_517,In_357,In_318);
nand U518 (N_518,In_60,In_758);
or U519 (N_519,In_21,In_324);
and U520 (N_520,In_45,In_365);
nor U521 (N_521,In_848,In_61);
and U522 (N_522,In_374,In_387);
or U523 (N_523,In_631,In_195);
and U524 (N_524,In_615,In_296);
and U525 (N_525,In_769,In_729);
and U526 (N_526,In_917,In_455);
and U527 (N_527,In_709,In_490);
and U528 (N_528,In_217,In_290);
nor U529 (N_529,In_816,In_174);
and U530 (N_530,In_496,In_790);
and U531 (N_531,In_33,In_261);
and U532 (N_532,In_271,In_426);
and U533 (N_533,In_322,In_897);
nor U534 (N_534,In_840,In_304);
nor U535 (N_535,In_246,In_312);
or U536 (N_536,In_155,In_340);
nor U537 (N_537,In_20,In_71);
and U538 (N_538,In_110,In_121);
and U539 (N_539,In_406,In_747);
and U540 (N_540,In_810,In_645);
nor U541 (N_541,In_382,In_259);
or U542 (N_542,In_881,In_767);
nor U543 (N_543,In_464,In_684);
or U544 (N_544,In_273,In_1);
nand U545 (N_545,In_379,In_794);
nor U546 (N_546,In_469,In_47);
nand U547 (N_547,In_645,In_409);
and U548 (N_548,In_373,In_31);
nor U549 (N_549,In_782,In_592);
nor U550 (N_550,In_974,In_743);
nor U551 (N_551,In_255,In_412);
or U552 (N_552,In_652,In_386);
or U553 (N_553,In_90,In_503);
and U554 (N_554,In_405,In_307);
nor U555 (N_555,In_188,In_462);
nand U556 (N_556,In_729,In_456);
or U557 (N_557,In_784,In_971);
nor U558 (N_558,In_547,In_717);
and U559 (N_559,In_65,In_139);
or U560 (N_560,In_413,In_578);
and U561 (N_561,In_887,In_244);
nor U562 (N_562,In_800,In_932);
and U563 (N_563,In_85,In_342);
nand U564 (N_564,In_495,In_892);
nand U565 (N_565,In_338,In_61);
and U566 (N_566,In_344,In_775);
xor U567 (N_567,In_985,In_167);
nor U568 (N_568,In_668,In_279);
nand U569 (N_569,In_419,In_677);
or U570 (N_570,In_522,In_611);
or U571 (N_571,In_956,In_299);
nand U572 (N_572,In_84,In_339);
or U573 (N_573,In_712,In_924);
and U574 (N_574,In_947,In_187);
nand U575 (N_575,In_433,In_91);
and U576 (N_576,In_182,In_115);
xnor U577 (N_577,In_493,In_163);
or U578 (N_578,In_5,In_477);
nand U579 (N_579,In_215,In_58);
nor U580 (N_580,In_187,In_520);
nand U581 (N_581,In_86,In_958);
nand U582 (N_582,In_425,In_828);
nand U583 (N_583,In_80,In_300);
nor U584 (N_584,In_631,In_521);
and U585 (N_585,In_667,In_889);
nand U586 (N_586,In_69,In_263);
or U587 (N_587,In_106,In_114);
and U588 (N_588,In_186,In_229);
nor U589 (N_589,In_341,In_931);
or U590 (N_590,In_165,In_55);
or U591 (N_591,In_122,In_321);
or U592 (N_592,In_530,In_611);
xor U593 (N_593,In_108,In_575);
nor U594 (N_594,In_708,In_459);
nor U595 (N_595,In_603,In_191);
xnor U596 (N_596,In_915,In_979);
or U597 (N_597,In_812,In_125);
and U598 (N_598,In_369,In_47);
nor U599 (N_599,In_799,In_903);
or U600 (N_600,In_474,In_622);
and U601 (N_601,In_75,In_61);
nand U602 (N_602,In_224,In_449);
and U603 (N_603,In_261,In_137);
or U604 (N_604,In_382,In_812);
and U605 (N_605,In_350,In_628);
nor U606 (N_606,In_661,In_712);
or U607 (N_607,In_188,In_750);
nand U608 (N_608,In_113,In_687);
and U609 (N_609,In_503,In_187);
nand U610 (N_610,In_873,In_430);
nand U611 (N_611,In_722,In_3);
or U612 (N_612,In_112,In_878);
or U613 (N_613,In_692,In_59);
and U614 (N_614,In_434,In_598);
nor U615 (N_615,In_178,In_503);
nor U616 (N_616,In_114,In_262);
nor U617 (N_617,In_436,In_840);
or U618 (N_618,In_525,In_488);
nand U619 (N_619,In_474,In_1);
nand U620 (N_620,In_522,In_995);
and U621 (N_621,In_9,In_515);
nor U622 (N_622,In_834,In_718);
nand U623 (N_623,In_284,In_471);
and U624 (N_624,In_379,In_332);
nand U625 (N_625,In_331,In_712);
and U626 (N_626,In_13,In_403);
nor U627 (N_627,In_431,In_278);
and U628 (N_628,In_156,In_135);
or U629 (N_629,In_63,In_998);
and U630 (N_630,In_124,In_462);
and U631 (N_631,In_924,In_881);
or U632 (N_632,In_503,In_435);
nand U633 (N_633,In_420,In_663);
nand U634 (N_634,In_144,In_490);
and U635 (N_635,In_551,In_819);
and U636 (N_636,In_331,In_276);
and U637 (N_637,In_60,In_8);
nor U638 (N_638,In_713,In_499);
and U639 (N_639,In_507,In_244);
or U640 (N_640,In_104,In_316);
and U641 (N_641,In_137,In_782);
nor U642 (N_642,In_587,In_781);
nor U643 (N_643,In_292,In_183);
and U644 (N_644,In_672,In_295);
nand U645 (N_645,In_345,In_41);
or U646 (N_646,In_518,In_324);
nor U647 (N_647,In_271,In_81);
nor U648 (N_648,In_874,In_861);
nand U649 (N_649,In_661,In_203);
or U650 (N_650,In_155,In_752);
nand U651 (N_651,In_935,In_352);
nor U652 (N_652,In_362,In_978);
nor U653 (N_653,In_931,In_510);
or U654 (N_654,In_576,In_693);
or U655 (N_655,In_814,In_156);
nor U656 (N_656,In_656,In_8);
nand U657 (N_657,In_155,In_293);
nor U658 (N_658,In_317,In_404);
nor U659 (N_659,In_490,In_823);
or U660 (N_660,In_188,In_160);
nor U661 (N_661,In_37,In_865);
xnor U662 (N_662,In_628,In_176);
nor U663 (N_663,In_364,In_851);
nand U664 (N_664,In_991,In_697);
nand U665 (N_665,In_768,In_486);
nor U666 (N_666,In_525,In_504);
nand U667 (N_667,In_779,In_379);
nand U668 (N_668,In_7,In_220);
nand U669 (N_669,In_625,In_109);
and U670 (N_670,In_494,In_88);
and U671 (N_671,In_371,In_940);
nor U672 (N_672,In_528,In_308);
or U673 (N_673,In_995,In_655);
or U674 (N_674,In_612,In_744);
and U675 (N_675,In_910,In_650);
and U676 (N_676,In_873,In_301);
or U677 (N_677,In_605,In_858);
nor U678 (N_678,In_933,In_186);
nand U679 (N_679,In_117,In_980);
and U680 (N_680,In_229,In_673);
xor U681 (N_681,In_391,In_118);
or U682 (N_682,In_558,In_958);
or U683 (N_683,In_101,In_103);
and U684 (N_684,In_236,In_191);
nor U685 (N_685,In_294,In_398);
nor U686 (N_686,In_292,In_27);
nand U687 (N_687,In_837,In_562);
and U688 (N_688,In_194,In_930);
and U689 (N_689,In_920,In_440);
or U690 (N_690,In_726,In_765);
and U691 (N_691,In_277,In_662);
nand U692 (N_692,In_296,In_946);
or U693 (N_693,In_224,In_944);
nor U694 (N_694,In_828,In_674);
nand U695 (N_695,In_646,In_103);
nand U696 (N_696,In_126,In_943);
nand U697 (N_697,In_79,In_154);
and U698 (N_698,In_520,In_139);
nor U699 (N_699,In_60,In_874);
nand U700 (N_700,In_870,In_165);
and U701 (N_701,In_441,In_989);
or U702 (N_702,In_804,In_288);
or U703 (N_703,In_249,In_868);
nor U704 (N_704,In_115,In_294);
and U705 (N_705,In_527,In_567);
or U706 (N_706,In_899,In_875);
nor U707 (N_707,In_327,In_393);
and U708 (N_708,In_807,In_256);
nor U709 (N_709,In_522,In_555);
and U710 (N_710,In_114,In_999);
xnor U711 (N_711,In_961,In_549);
or U712 (N_712,In_654,In_392);
and U713 (N_713,In_20,In_127);
nand U714 (N_714,In_165,In_364);
nor U715 (N_715,In_866,In_156);
nand U716 (N_716,In_734,In_643);
and U717 (N_717,In_88,In_964);
or U718 (N_718,In_331,In_165);
and U719 (N_719,In_339,In_499);
nand U720 (N_720,In_97,In_122);
and U721 (N_721,In_268,In_921);
nand U722 (N_722,In_175,In_850);
or U723 (N_723,In_310,In_250);
nor U724 (N_724,In_993,In_23);
xor U725 (N_725,In_426,In_569);
and U726 (N_726,In_844,In_953);
and U727 (N_727,In_685,In_462);
nor U728 (N_728,In_721,In_620);
nor U729 (N_729,In_556,In_490);
xnor U730 (N_730,In_962,In_768);
or U731 (N_731,In_585,In_124);
nand U732 (N_732,In_931,In_431);
or U733 (N_733,In_796,In_0);
or U734 (N_734,In_283,In_474);
nand U735 (N_735,In_843,In_967);
nor U736 (N_736,In_916,In_692);
nor U737 (N_737,In_16,In_118);
and U738 (N_738,In_150,In_838);
nor U739 (N_739,In_867,In_473);
and U740 (N_740,In_59,In_366);
xnor U741 (N_741,In_64,In_992);
or U742 (N_742,In_965,In_695);
and U743 (N_743,In_419,In_147);
nand U744 (N_744,In_374,In_978);
nor U745 (N_745,In_685,In_354);
nand U746 (N_746,In_565,In_68);
or U747 (N_747,In_948,In_321);
nand U748 (N_748,In_73,In_675);
and U749 (N_749,In_703,In_978);
nor U750 (N_750,In_51,In_101);
and U751 (N_751,In_50,In_888);
nand U752 (N_752,In_840,In_889);
nor U753 (N_753,In_868,In_778);
and U754 (N_754,In_456,In_996);
or U755 (N_755,In_325,In_297);
nor U756 (N_756,In_884,In_483);
or U757 (N_757,In_81,In_328);
or U758 (N_758,In_878,In_796);
nor U759 (N_759,In_673,In_981);
and U760 (N_760,In_254,In_371);
and U761 (N_761,In_114,In_201);
or U762 (N_762,In_372,In_219);
and U763 (N_763,In_75,In_419);
nor U764 (N_764,In_274,In_83);
nor U765 (N_765,In_706,In_221);
and U766 (N_766,In_571,In_744);
nor U767 (N_767,In_283,In_779);
nor U768 (N_768,In_432,In_28);
nand U769 (N_769,In_939,In_490);
nand U770 (N_770,In_789,In_320);
or U771 (N_771,In_160,In_299);
nor U772 (N_772,In_16,In_53);
and U773 (N_773,In_856,In_847);
nand U774 (N_774,In_648,In_36);
or U775 (N_775,In_544,In_228);
nor U776 (N_776,In_941,In_593);
nor U777 (N_777,In_122,In_998);
nand U778 (N_778,In_951,In_263);
and U779 (N_779,In_222,In_806);
or U780 (N_780,In_899,In_139);
nor U781 (N_781,In_250,In_718);
or U782 (N_782,In_870,In_758);
nor U783 (N_783,In_288,In_458);
nor U784 (N_784,In_170,In_430);
and U785 (N_785,In_945,In_497);
or U786 (N_786,In_933,In_947);
nor U787 (N_787,In_545,In_205);
nor U788 (N_788,In_582,In_937);
or U789 (N_789,In_108,In_816);
nor U790 (N_790,In_778,In_252);
or U791 (N_791,In_581,In_709);
nand U792 (N_792,In_466,In_6);
nand U793 (N_793,In_225,In_214);
and U794 (N_794,In_48,In_830);
and U795 (N_795,In_377,In_6);
and U796 (N_796,In_711,In_950);
nor U797 (N_797,In_469,In_904);
and U798 (N_798,In_999,In_104);
or U799 (N_799,In_538,In_978);
and U800 (N_800,In_143,In_79);
and U801 (N_801,In_140,In_941);
nor U802 (N_802,In_213,In_973);
nand U803 (N_803,In_782,In_825);
and U804 (N_804,In_28,In_88);
nor U805 (N_805,In_771,In_6);
xnor U806 (N_806,In_161,In_236);
and U807 (N_807,In_400,In_449);
or U808 (N_808,In_142,In_291);
or U809 (N_809,In_834,In_864);
nand U810 (N_810,In_727,In_509);
or U811 (N_811,In_569,In_440);
nor U812 (N_812,In_616,In_533);
and U813 (N_813,In_775,In_945);
nor U814 (N_814,In_224,In_910);
nor U815 (N_815,In_200,In_11);
or U816 (N_816,In_457,In_443);
or U817 (N_817,In_192,In_880);
nor U818 (N_818,In_924,In_148);
nand U819 (N_819,In_998,In_493);
nand U820 (N_820,In_950,In_822);
and U821 (N_821,In_682,In_102);
nor U822 (N_822,In_187,In_251);
nor U823 (N_823,In_915,In_290);
and U824 (N_824,In_606,In_407);
nor U825 (N_825,In_209,In_528);
nand U826 (N_826,In_401,In_585);
and U827 (N_827,In_523,In_919);
nor U828 (N_828,In_621,In_129);
and U829 (N_829,In_47,In_675);
nand U830 (N_830,In_579,In_104);
and U831 (N_831,In_384,In_424);
or U832 (N_832,In_851,In_667);
nor U833 (N_833,In_947,In_166);
and U834 (N_834,In_230,In_103);
nor U835 (N_835,In_917,In_353);
nor U836 (N_836,In_461,In_740);
nor U837 (N_837,In_708,In_571);
nand U838 (N_838,In_671,In_425);
and U839 (N_839,In_987,In_630);
or U840 (N_840,In_255,In_348);
nor U841 (N_841,In_121,In_946);
nor U842 (N_842,In_499,In_840);
or U843 (N_843,In_124,In_1);
or U844 (N_844,In_669,In_339);
and U845 (N_845,In_152,In_268);
and U846 (N_846,In_337,In_380);
nand U847 (N_847,In_223,In_467);
nand U848 (N_848,In_395,In_851);
nand U849 (N_849,In_428,In_312);
nor U850 (N_850,In_511,In_810);
nor U851 (N_851,In_199,In_471);
or U852 (N_852,In_694,In_88);
nor U853 (N_853,In_972,In_298);
and U854 (N_854,In_599,In_764);
and U855 (N_855,In_735,In_635);
xnor U856 (N_856,In_724,In_959);
and U857 (N_857,In_963,In_633);
nor U858 (N_858,In_935,In_6);
or U859 (N_859,In_855,In_547);
nor U860 (N_860,In_504,In_729);
and U861 (N_861,In_152,In_428);
nor U862 (N_862,In_406,In_762);
nor U863 (N_863,In_874,In_927);
nand U864 (N_864,In_336,In_688);
nand U865 (N_865,In_561,In_137);
nor U866 (N_866,In_854,In_996);
nand U867 (N_867,In_316,In_444);
nor U868 (N_868,In_155,In_351);
and U869 (N_869,In_891,In_303);
and U870 (N_870,In_528,In_121);
or U871 (N_871,In_769,In_186);
nand U872 (N_872,In_587,In_822);
nand U873 (N_873,In_250,In_735);
nand U874 (N_874,In_250,In_175);
and U875 (N_875,In_157,In_449);
and U876 (N_876,In_429,In_956);
and U877 (N_877,In_325,In_802);
nand U878 (N_878,In_366,In_821);
nand U879 (N_879,In_182,In_532);
nand U880 (N_880,In_930,In_637);
nor U881 (N_881,In_896,In_945);
and U882 (N_882,In_719,In_414);
nor U883 (N_883,In_927,In_489);
or U884 (N_884,In_414,In_473);
nand U885 (N_885,In_721,In_764);
and U886 (N_886,In_266,In_226);
and U887 (N_887,In_73,In_488);
and U888 (N_888,In_673,In_167);
and U889 (N_889,In_861,In_368);
and U890 (N_890,In_884,In_239);
nand U891 (N_891,In_981,In_696);
nor U892 (N_892,In_944,In_23);
or U893 (N_893,In_972,In_581);
or U894 (N_894,In_715,In_672);
nor U895 (N_895,In_433,In_702);
nand U896 (N_896,In_814,In_333);
or U897 (N_897,In_796,In_905);
nand U898 (N_898,In_562,In_295);
nor U899 (N_899,In_291,In_641);
nor U900 (N_900,In_210,In_290);
nor U901 (N_901,In_758,In_987);
nor U902 (N_902,In_619,In_627);
nor U903 (N_903,In_674,In_831);
and U904 (N_904,In_259,In_784);
nor U905 (N_905,In_492,In_59);
nand U906 (N_906,In_513,In_343);
and U907 (N_907,In_926,In_965);
or U908 (N_908,In_681,In_167);
and U909 (N_909,In_522,In_766);
or U910 (N_910,In_303,In_168);
or U911 (N_911,In_857,In_498);
or U912 (N_912,In_696,In_849);
or U913 (N_913,In_666,In_946);
nand U914 (N_914,In_627,In_580);
or U915 (N_915,In_51,In_588);
nor U916 (N_916,In_150,In_217);
nand U917 (N_917,In_108,In_145);
nand U918 (N_918,In_173,In_778);
nor U919 (N_919,In_110,In_995);
nor U920 (N_920,In_178,In_672);
nand U921 (N_921,In_552,In_97);
nand U922 (N_922,In_582,In_942);
nor U923 (N_923,In_606,In_507);
nand U924 (N_924,In_341,In_686);
and U925 (N_925,In_37,In_268);
nand U926 (N_926,In_295,In_986);
nor U927 (N_927,In_877,In_191);
nor U928 (N_928,In_41,In_212);
nand U929 (N_929,In_36,In_873);
nand U930 (N_930,In_597,In_906);
and U931 (N_931,In_52,In_428);
nand U932 (N_932,In_690,In_788);
nor U933 (N_933,In_673,In_613);
or U934 (N_934,In_654,In_842);
or U935 (N_935,In_376,In_834);
or U936 (N_936,In_137,In_35);
nand U937 (N_937,In_93,In_624);
nor U938 (N_938,In_101,In_643);
and U939 (N_939,In_983,In_326);
or U940 (N_940,In_475,In_920);
xor U941 (N_941,In_13,In_320);
and U942 (N_942,In_519,In_678);
or U943 (N_943,In_352,In_570);
nor U944 (N_944,In_215,In_210);
nand U945 (N_945,In_766,In_353);
or U946 (N_946,In_627,In_599);
or U947 (N_947,In_933,In_30);
nor U948 (N_948,In_14,In_658);
nand U949 (N_949,In_426,In_56);
and U950 (N_950,In_219,In_377);
nand U951 (N_951,In_470,In_584);
or U952 (N_952,In_348,In_862);
or U953 (N_953,In_818,In_313);
nand U954 (N_954,In_167,In_175);
and U955 (N_955,In_970,In_454);
nand U956 (N_956,In_430,In_198);
and U957 (N_957,In_750,In_583);
nor U958 (N_958,In_198,In_603);
or U959 (N_959,In_650,In_911);
and U960 (N_960,In_266,In_93);
nor U961 (N_961,In_710,In_357);
nor U962 (N_962,In_606,In_580);
and U963 (N_963,In_422,In_445);
or U964 (N_964,In_155,In_737);
or U965 (N_965,In_422,In_935);
xnor U966 (N_966,In_515,In_495);
or U967 (N_967,In_307,In_577);
and U968 (N_968,In_648,In_408);
nor U969 (N_969,In_537,In_713);
or U970 (N_970,In_668,In_230);
nor U971 (N_971,In_772,In_931);
nor U972 (N_972,In_847,In_184);
or U973 (N_973,In_265,In_318);
nor U974 (N_974,In_268,In_129);
and U975 (N_975,In_867,In_931);
nor U976 (N_976,In_22,In_827);
or U977 (N_977,In_567,In_993);
or U978 (N_978,In_829,In_520);
nand U979 (N_979,In_914,In_39);
nor U980 (N_980,In_62,In_975);
or U981 (N_981,In_528,In_110);
nand U982 (N_982,In_7,In_572);
or U983 (N_983,In_433,In_653);
xor U984 (N_984,In_259,In_707);
nand U985 (N_985,In_976,In_29);
or U986 (N_986,In_962,In_863);
or U987 (N_987,In_678,In_670);
or U988 (N_988,In_837,In_724);
nor U989 (N_989,In_944,In_260);
and U990 (N_990,In_172,In_716);
xor U991 (N_991,In_6,In_882);
nor U992 (N_992,In_196,In_782);
nand U993 (N_993,In_690,In_393);
nor U994 (N_994,In_113,In_635);
or U995 (N_995,In_510,In_911);
and U996 (N_996,In_577,In_492);
nand U997 (N_997,In_670,In_189);
or U998 (N_998,In_710,In_24);
and U999 (N_999,In_305,In_651);
and U1000 (N_1000,N_287,N_387);
and U1001 (N_1001,N_180,N_777);
or U1002 (N_1002,N_259,N_700);
nor U1003 (N_1003,N_714,N_799);
and U1004 (N_1004,N_890,N_741);
nand U1005 (N_1005,N_83,N_970);
xor U1006 (N_1006,N_440,N_504);
and U1007 (N_1007,N_571,N_577);
and U1008 (N_1008,N_573,N_731);
nand U1009 (N_1009,N_385,N_167);
nand U1010 (N_1010,N_567,N_583);
and U1011 (N_1011,N_106,N_818);
and U1012 (N_1012,N_436,N_552);
nor U1013 (N_1013,N_726,N_177);
and U1014 (N_1014,N_626,N_304);
and U1015 (N_1015,N_527,N_399);
or U1016 (N_1016,N_319,N_644);
or U1017 (N_1017,N_640,N_401);
or U1018 (N_1018,N_851,N_457);
and U1019 (N_1019,N_913,N_963);
and U1020 (N_1020,N_172,N_797);
nor U1021 (N_1021,N_703,N_856);
or U1022 (N_1022,N_207,N_85);
nand U1023 (N_1023,N_189,N_569);
or U1024 (N_1024,N_697,N_730);
nor U1025 (N_1025,N_672,N_443);
or U1026 (N_1026,N_173,N_761);
nand U1027 (N_1027,N_953,N_84);
and U1028 (N_1028,N_434,N_215);
nor U1029 (N_1029,N_798,N_742);
nor U1030 (N_1030,N_525,N_727);
and U1031 (N_1031,N_439,N_29);
nor U1032 (N_1032,N_629,N_193);
or U1033 (N_1033,N_128,N_4);
nand U1034 (N_1034,N_598,N_398);
nor U1035 (N_1035,N_364,N_986);
nand U1036 (N_1036,N_283,N_668);
nand U1037 (N_1037,N_1,N_546);
xor U1038 (N_1038,N_45,N_297);
nor U1039 (N_1039,N_968,N_565);
and U1040 (N_1040,N_479,N_253);
nand U1041 (N_1041,N_605,N_365);
and U1042 (N_1042,N_371,N_453);
and U1043 (N_1043,N_660,N_770);
nand U1044 (N_1044,N_678,N_693);
or U1045 (N_1045,N_757,N_514);
or U1046 (N_1046,N_216,N_493);
or U1047 (N_1047,N_184,N_465);
and U1048 (N_1048,N_871,N_853);
nand U1049 (N_1049,N_114,N_395);
nand U1050 (N_1050,N_421,N_280);
and U1051 (N_1051,N_539,N_636);
or U1052 (N_1052,N_46,N_758);
and U1053 (N_1053,N_33,N_271);
or U1054 (N_1054,N_307,N_987);
or U1055 (N_1055,N_885,N_790);
nand U1056 (N_1056,N_725,N_136);
and U1057 (N_1057,N_554,N_494);
nand U1058 (N_1058,N_904,N_745);
or U1059 (N_1059,N_22,N_467);
nor U1060 (N_1060,N_409,N_833);
nand U1061 (N_1061,N_375,N_268);
and U1062 (N_1062,N_445,N_610);
nor U1063 (N_1063,N_767,N_562);
nand U1064 (N_1064,N_591,N_596);
xnor U1065 (N_1065,N_729,N_988);
and U1066 (N_1066,N_736,N_786);
or U1067 (N_1067,N_495,N_828);
and U1068 (N_1068,N_850,N_911);
nand U1069 (N_1069,N_463,N_775);
or U1070 (N_1070,N_196,N_219);
and U1071 (N_1071,N_373,N_405);
and U1072 (N_1072,N_928,N_93);
nor U1073 (N_1073,N_276,N_649);
or U1074 (N_1074,N_55,N_146);
nand U1075 (N_1075,N_151,N_901);
and U1076 (N_1076,N_972,N_766);
nand U1077 (N_1077,N_597,N_400);
and U1078 (N_1078,N_460,N_675);
nor U1079 (N_1079,N_31,N_165);
and U1080 (N_1080,N_367,N_892);
or U1081 (N_1081,N_903,N_582);
nor U1082 (N_1082,N_506,N_242);
and U1083 (N_1083,N_384,N_864);
nand U1084 (N_1084,N_108,N_210);
nand U1085 (N_1085,N_9,N_168);
nor U1086 (N_1086,N_221,N_360);
and U1087 (N_1087,N_921,N_812);
nand U1088 (N_1088,N_570,N_192);
or U1089 (N_1089,N_320,N_902);
and U1090 (N_1090,N_559,N_334);
nand U1091 (N_1091,N_336,N_578);
and U1092 (N_1092,N_388,N_366);
or U1093 (N_1093,N_540,N_809);
and U1094 (N_1094,N_279,N_915);
or U1095 (N_1095,N_608,N_769);
or U1096 (N_1096,N_722,N_148);
or U1097 (N_1097,N_2,N_286);
and U1098 (N_1098,N_438,N_485);
nor U1099 (N_1099,N_471,N_718);
or U1100 (N_1100,N_249,N_752);
or U1101 (N_1101,N_446,N_225);
nor U1102 (N_1102,N_819,N_138);
or U1103 (N_1103,N_418,N_352);
nor U1104 (N_1104,N_99,N_262);
and U1105 (N_1105,N_665,N_81);
and U1106 (N_1106,N_18,N_557);
xor U1107 (N_1107,N_916,N_228);
nor U1108 (N_1108,N_109,N_754);
and U1109 (N_1109,N_964,N_590);
and U1110 (N_1110,N_692,N_542);
or U1111 (N_1111,N_397,N_171);
nor U1112 (N_1112,N_240,N_734);
nor U1113 (N_1113,N_218,N_865);
and U1114 (N_1114,N_867,N_309);
and U1115 (N_1115,N_501,N_245);
nor U1116 (N_1116,N_5,N_427);
nand U1117 (N_1117,N_633,N_651);
or U1118 (N_1118,N_459,N_498);
nor U1119 (N_1119,N_881,N_480);
or U1120 (N_1120,N_611,N_404);
nor U1121 (N_1121,N_430,N_639);
or U1122 (N_1122,N_222,N_181);
and U1123 (N_1123,N_76,N_344);
or U1124 (N_1124,N_251,N_133);
or U1125 (N_1125,N_637,N_305);
xor U1126 (N_1126,N_792,N_879);
or U1127 (N_1127,N_878,N_90);
or U1128 (N_1128,N_842,N_95);
nand U1129 (N_1129,N_607,N_604);
nor U1130 (N_1130,N_803,N_947);
and U1131 (N_1131,N_965,N_310);
or U1132 (N_1132,N_325,N_298);
nand U1133 (N_1133,N_513,N_236);
or U1134 (N_1134,N_969,N_346);
and U1135 (N_1135,N_713,N_232);
nand U1136 (N_1136,N_635,N_201);
and U1137 (N_1137,N_424,N_743);
xor U1138 (N_1138,N_21,N_709);
nor U1139 (N_1139,N_353,N_120);
xor U1140 (N_1140,N_224,N_780);
nor U1141 (N_1141,N_813,N_117);
or U1142 (N_1142,N_744,N_950);
or U1143 (N_1143,N_343,N_348);
or U1144 (N_1144,N_284,N_464);
and U1145 (N_1145,N_671,N_720);
nor U1146 (N_1146,N_689,N_175);
or U1147 (N_1147,N_588,N_470);
nor U1148 (N_1148,N_795,N_526);
nor U1149 (N_1149,N_303,N_265);
nor U1150 (N_1150,N_428,N_302);
or U1151 (N_1151,N_42,N_179);
nor U1152 (N_1152,N_994,N_938);
and U1153 (N_1153,N_814,N_250);
nand U1154 (N_1154,N_535,N_980);
nor U1155 (N_1155,N_264,N_458);
nor U1156 (N_1156,N_880,N_740);
nand U1157 (N_1157,N_282,N_386);
nor U1158 (N_1158,N_505,N_581);
nor U1159 (N_1159,N_489,N_716);
xnor U1160 (N_1160,N_866,N_929);
nand U1161 (N_1161,N_43,N_337);
nor U1162 (N_1162,N_951,N_198);
or U1163 (N_1163,N_886,N_960);
nor U1164 (N_1164,N_503,N_350);
nor U1165 (N_1165,N_884,N_162);
or U1166 (N_1166,N_946,N_324);
and U1167 (N_1167,N_723,N_79);
or U1168 (N_1168,N_912,N_132);
nor U1169 (N_1169,N_876,N_482);
and U1170 (N_1170,N_149,N_357);
and U1171 (N_1171,N_593,N_241);
nand U1172 (N_1172,N_936,N_807);
nand U1173 (N_1173,N_724,N_783);
or U1174 (N_1174,N_231,N_696);
or U1175 (N_1175,N_256,N_155);
or U1176 (N_1176,N_707,N_558);
or U1177 (N_1177,N_389,N_316);
nor U1178 (N_1178,N_206,N_717);
or U1179 (N_1179,N_899,N_333);
nor U1180 (N_1180,N_134,N_574);
nand U1181 (N_1181,N_930,N_285);
nand U1182 (N_1182,N_174,N_39);
xor U1183 (N_1183,N_733,N_516);
or U1184 (N_1184,N_288,N_624);
or U1185 (N_1185,N_308,N_243);
or U1186 (N_1186,N_112,N_918);
nand U1187 (N_1187,N_983,N_555);
nand U1188 (N_1188,N_977,N_143);
nand U1189 (N_1189,N_273,N_802);
or U1190 (N_1190,N_50,N_576);
nor U1191 (N_1191,N_966,N_263);
nand U1192 (N_1192,N_234,N_419);
and U1193 (N_1193,N_200,N_104);
nand U1194 (N_1194,N_688,N_153);
and U1195 (N_1195,N_474,N_380);
and U1196 (N_1196,N_774,N_657);
or U1197 (N_1197,N_289,N_202);
or U1198 (N_1198,N_254,N_603);
or U1199 (N_1199,N_47,N_278);
xnor U1200 (N_1200,N_322,N_701);
nand U1201 (N_1201,N_166,N_759);
nand U1202 (N_1202,N_676,N_164);
and U1203 (N_1203,N_237,N_594);
nor U1204 (N_1204,N_585,N_580);
nand U1205 (N_1205,N_975,N_119);
nand U1206 (N_1206,N_383,N_49);
nor U1207 (N_1207,N_779,N_848);
nor U1208 (N_1208,N_19,N_57);
nand U1209 (N_1209,N_118,N_432);
nand U1210 (N_1210,N_919,N_486);
and U1211 (N_1211,N_822,N_313);
nor U1212 (N_1212,N_628,N_186);
nand U1213 (N_1213,N_417,N_52);
and U1214 (N_1214,N_997,N_408);
nand U1215 (N_1215,N_32,N_188);
nor U1216 (N_1216,N_238,N_961);
and U1217 (N_1217,N_497,N_949);
and U1218 (N_1218,N_13,N_3);
nor U1219 (N_1219,N_548,N_306);
nand U1220 (N_1220,N_553,N_156);
or U1221 (N_1221,N_187,N_959);
nand U1222 (N_1222,N_579,N_979);
nand U1223 (N_1223,N_650,N_61);
nor U1224 (N_1224,N_272,N_859);
and U1225 (N_1225,N_209,N_97);
or U1226 (N_1226,N_447,N_315);
xnor U1227 (N_1227,N_327,N_411);
or U1228 (N_1228,N_584,N_329);
nand U1229 (N_1229,N_53,N_995);
and U1230 (N_1230,N_875,N_528);
and U1231 (N_1231,N_220,N_169);
xor U1232 (N_1232,N_862,N_756);
nor U1233 (N_1233,N_163,N_361);
nand U1234 (N_1234,N_711,N_840);
nand U1235 (N_1235,N_437,N_37);
nand U1236 (N_1236,N_735,N_382);
or U1237 (N_1237,N_974,N_719);
or U1238 (N_1238,N_512,N_917);
or U1239 (N_1239,N_990,N_816);
nor U1240 (N_1240,N_423,N_147);
and U1241 (N_1241,N_834,N_748);
nor U1242 (N_1242,N_281,N_10);
and U1243 (N_1243,N_69,N_998);
nand U1244 (N_1244,N_907,N_652);
nand U1245 (N_1245,N_762,N_461);
nand U1246 (N_1246,N_127,N_900);
nor U1247 (N_1247,N_511,N_967);
nand U1248 (N_1248,N_372,N_673);
nor U1249 (N_1249,N_451,N_402);
or U1250 (N_1250,N_686,N_616);
nand U1251 (N_1251,N_931,N_868);
nand U1252 (N_1252,N_507,N_870);
nand U1253 (N_1253,N_606,N_541);
nor U1254 (N_1254,N_347,N_142);
nand U1255 (N_1255,N_369,N_80);
and U1256 (N_1256,N_623,N_768);
nand U1257 (N_1257,N_462,N_801);
or U1258 (N_1258,N_826,N_64);
or U1259 (N_1259,N_70,N_806);
nand U1260 (N_1260,N_92,N_292);
and U1261 (N_1261,N_277,N_137);
nand U1262 (N_1262,N_522,N_749);
nand U1263 (N_1263,N_269,N_661);
nor U1264 (N_1264,N_945,N_721);
nor U1265 (N_1265,N_784,N_121);
and U1266 (N_1266,N_510,N_294);
and U1267 (N_1267,N_993,N_519);
or U1268 (N_1268,N_564,N_690);
or U1269 (N_1269,N_508,N_587);
and U1270 (N_1270,N_659,N_65);
or U1271 (N_1271,N_26,N_328);
and U1272 (N_1272,N_331,N_176);
and U1273 (N_1273,N_183,N_499);
nand U1274 (N_1274,N_17,N_103);
nor U1275 (N_1275,N_299,N_185);
or U1276 (N_1276,N_252,N_877);
nor U1277 (N_1277,N_248,N_989);
xnor U1278 (N_1278,N_483,N_811);
or U1279 (N_1279,N_547,N_191);
nand U1280 (N_1280,N_356,N_999);
xor U1281 (N_1281,N_330,N_976);
and U1282 (N_1282,N_832,N_627);
or U1283 (N_1283,N_694,N_561);
nand U1284 (N_1284,N_394,N_379);
nand U1285 (N_1285,N_481,N_894);
and U1286 (N_1286,N_664,N_791);
nand U1287 (N_1287,N_469,N_182);
nand U1288 (N_1288,N_227,N_614);
nor U1289 (N_1289,N_72,N_837);
or U1290 (N_1290,N_684,N_750);
nand U1291 (N_1291,N_407,N_682);
or U1292 (N_1292,N_125,N_962);
and U1293 (N_1293,N_595,N_543);
nor U1294 (N_1294,N_533,N_293);
and U1295 (N_1295,N_170,N_641);
and U1296 (N_1296,N_58,N_520);
or U1297 (N_1297,N_488,N_345);
nand U1298 (N_1298,N_632,N_144);
and U1299 (N_1299,N_537,N_645);
and U1300 (N_1300,N_178,N_824);
and U1301 (N_1301,N_266,N_15);
or U1302 (N_1302,N_845,N_392);
and U1303 (N_1303,N_896,N_708);
and U1304 (N_1304,N_122,N_702);
and U1305 (N_1305,N_270,N_23);
nor U1306 (N_1306,N_924,N_35);
nor U1307 (N_1307,N_145,N_521);
nand U1308 (N_1308,N_781,N_937);
or U1309 (N_1309,N_27,N_821);
or U1310 (N_1310,N_891,N_883);
or U1311 (N_1311,N_914,N_638);
xnor U1312 (N_1312,N_468,N_620);
and U1313 (N_1313,N_41,N_442);
or U1314 (N_1314,N_981,N_698);
nor U1315 (N_1315,N_73,N_844);
nand U1316 (N_1316,N_422,N_575);
nor U1317 (N_1317,N_88,N_509);
and U1318 (N_1318,N_275,N_825);
and U1319 (N_1319,N_332,N_764);
nand U1320 (N_1320,N_454,N_518);
nor U1321 (N_1321,N_363,N_102);
and U1322 (N_1322,N_107,N_666);
nor U1323 (N_1323,N_190,N_955);
and U1324 (N_1324,N_158,N_496);
nand U1325 (N_1325,N_663,N_110);
or U1326 (N_1326,N_669,N_935);
nand U1327 (N_1327,N_341,N_323);
and U1328 (N_1328,N_476,N_592);
nor U1329 (N_1329,N_601,N_490);
nor U1330 (N_1330,N_441,N_551);
nand U1331 (N_1331,N_869,N_233);
or U1332 (N_1332,N_290,N_550);
and U1333 (N_1333,N_484,N_160);
and U1334 (N_1334,N_805,N_8);
or U1335 (N_1335,N_7,N_971);
or U1336 (N_1336,N_34,N_523);
nand U1337 (N_1337,N_159,N_808);
nor U1338 (N_1338,N_948,N_782);
nor U1339 (N_1339,N_391,N_670);
or U1340 (N_1340,N_785,N_625);
or U1341 (N_1341,N_213,N_91);
nand U1342 (N_1342,N_204,N_631);
nor U1343 (N_1343,N_530,N_849);
nand U1344 (N_1344,N_123,N_789);
and U1345 (N_1345,N_452,N_67);
nand U1346 (N_1346,N_679,N_939);
nor U1347 (N_1347,N_455,N_691);
nand U1348 (N_1348,N_429,N_773);
nand U1349 (N_1349,N_491,N_658);
and U1350 (N_1350,N_25,N_830);
xor U1351 (N_1351,N_677,N_942);
nor U1352 (N_1352,N_882,N_410);
or U1353 (N_1353,N_823,N_111);
and U1354 (N_1354,N_954,N_140);
or U1355 (N_1355,N_941,N_295);
nor U1356 (N_1356,N_154,N_314);
and U1357 (N_1357,N_362,N_642);
nand U1358 (N_1358,N_260,N_854);
or U1359 (N_1359,N_68,N_87);
or U1360 (N_1360,N_760,N_135);
and U1361 (N_1361,N_487,N_77);
nand U1362 (N_1362,N_472,N_318);
nor U1363 (N_1363,N_524,N_377);
and U1364 (N_1364,N_827,N_599);
and U1365 (N_1365,N_130,N_843);
nand U1366 (N_1366,N_621,N_98);
nand U1367 (N_1367,N_74,N_370);
and U1368 (N_1368,N_934,N_704);
and U1369 (N_1369,N_38,N_75);
and U1370 (N_1370,N_846,N_435);
nor U1371 (N_1371,N_923,N_630);
or U1372 (N_1372,N_985,N_208);
nor U1373 (N_1373,N_230,N_852);
or U1374 (N_1374,N_796,N_771);
xor U1375 (N_1375,N_211,N_710);
xor U1376 (N_1376,N_433,N_359);
nor U1377 (N_1377,N_393,N_214);
xnor U1378 (N_1378,N_246,N_197);
and U1379 (N_1379,N_887,N_728);
and U1380 (N_1380,N_312,N_247);
and U1381 (N_1381,N_71,N_705);
nor U1382 (N_1382,N_653,N_732);
and U1383 (N_1383,N_517,N_226);
nand U1384 (N_1384,N_534,N_431);
nand U1385 (N_1385,N_609,N_897);
or U1386 (N_1386,N_810,N_932);
or U1387 (N_1387,N_448,N_858);
and U1388 (N_1388,N_6,N_836);
nand U1389 (N_1389,N_763,N_847);
and U1390 (N_1390,N_681,N_612);
nand U1391 (N_1391,N_909,N_311);
or U1392 (N_1392,N_838,N_706);
or U1393 (N_1393,N_116,N_943);
and U1394 (N_1394,N_655,N_349);
nand U1395 (N_1395,N_376,N_910);
nor U1396 (N_1396,N_776,N_820);
nand U1397 (N_1397,N_96,N_863);
and U1398 (N_1398,N_82,N_478);
nor U1399 (N_1399,N_841,N_300);
nor U1400 (N_1400,N_56,N_667);
and U1401 (N_1401,N_321,N_893);
nand U1402 (N_1402,N_406,N_898);
nand U1403 (N_1403,N_0,N_340);
nor U1404 (N_1404,N_687,N_502);
and U1405 (N_1405,N_203,N_466);
nor U1406 (N_1406,N_531,N_982);
and U1407 (N_1407,N_683,N_63);
nor U1408 (N_1408,N_753,N_905);
and U1409 (N_1409,N_475,N_857);
nor U1410 (N_1410,N_992,N_60);
nand U1411 (N_1411,N_538,N_778);
and U1412 (N_1412,N_794,N_861);
nor U1413 (N_1413,N_831,N_456);
and U1414 (N_1414,N_355,N_100);
or U1415 (N_1415,N_933,N_205);
nand U1416 (N_1416,N_926,N_622);
nand U1417 (N_1417,N_925,N_450);
or U1418 (N_1418,N_66,N_24);
or U1419 (N_1419,N_712,N_229);
nor U1420 (N_1420,N_991,N_381);
or U1421 (N_1421,N_416,N_566);
nor U1422 (N_1422,N_788,N_16);
nand U1423 (N_1423,N_257,N_342);
xor U1424 (N_1424,N_646,N_973);
nor U1425 (N_1425,N_855,N_244);
or U1426 (N_1426,N_139,N_656);
and U1427 (N_1427,N_996,N_414);
and U1428 (N_1428,N_536,N_217);
nor U1429 (N_1429,N_426,N_415);
nand U1430 (N_1430,N_354,N_545);
or U1431 (N_1431,N_194,N_473);
or U1432 (N_1432,N_568,N_378);
nor U1433 (N_1433,N_772,N_685);
or U1434 (N_1434,N_793,N_739);
or U1435 (N_1435,N_787,N_358);
or U1436 (N_1436,N_927,N_680);
and U1437 (N_1437,N_89,N_14);
nand U1438 (N_1438,N_390,N_30);
nand U1439 (N_1439,N_940,N_413);
or U1440 (N_1440,N_560,N_105);
and U1441 (N_1441,N_695,N_78);
nor U1442 (N_1442,N_888,N_800);
nor U1443 (N_1443,N_860,N_738);
or U1444 (N_1444,N_634,N_563);
nand U1445 (N_1445,N_267,N_239);
nand U1446 (N_1446,N_500,N_150);
nand U1447 (N_1447,N_477,N_157);
nand U1448 (N_1448,N_296,N_124);
or U1449 (N_1449,N_544,N_746);
or U1450 (N_1450,N_54,N_195);
nor U1451 (N_1451,N_28,N_872);
or U1452 (N_1452,N_255,N_444);
or U1453 (N_1453,N_326,N_396);
nor U1454 (N_1454,N_532,N_335);
nor U1455 (N_1455,N_958,N_36);
nand U1456 (N_1456,N_12,N_835);
or U1457 (N_1457,N_374,N_600);
and U1458 (N_1458,N_908,N_152);
or U1459 (N_1459,N_952,N_161);
or U1460 (N_1460,N_619,N_40);
or U1461 (N_1461,N_86,N_339);
nor U1462 (N_1462,N_129,N_654);
or U1463 (N_1463,N_920,N_984);
or U1464 (N_1464,N_44,N_368);
nand U1465 (N_1465,N_301,N_11);
nor U1466 (N_1466,N_131,N_20);
or U1467 (N_1467,N_449,N_412);
and U1468 (N_1468,N_922,N_556);
or U1469 (N_1469,N_291,N_957);
or U1470 (N_1470,N_829,N_747);
nand U1471 (N_1471,N_515,N_648);
nor U1472 (N_1472,N_839,N_674);
nor U1473 (N_1473,N_895,N_715);
and U1474 (N_1474,N_425,N_62);
nor U1475 (N_1475,N_765,N_699);
nand U1476 (N_1476,N_572,N_873);
nand U1477 (N_1477,N_126,N_258);
or U1478 (N_1478,N_643,N_492);
nor U1479 (N_1479,N_115,N_817);
nor U1480 (N_1480,N_212,N_906);
or U1481 (N_1481,N_351,N_223);
nand U1482 (N_1482,N_94,N_549);
nand U1483 (N_1483,N_751,N_261);
and U1484 (N_1484,N_274,N_59);
nor U1485 (N_1485,N_48,N_617);
and U1486 (N_1486,N_529,N_317);
nand U1487 (N_1487,N_51,N_978);
or U1488 (N_1488,N_944,N_113);
or U1489 (N_1489,N_403,N_338);
nand U1490 (N_1490,N_647,N_589);
nor U1491 (N_1491,N_755,N_420);
and U1492 (N_1492,N_874,N_615);
xor U1493 (N_1493,N_199,N_602);
xnor U1494 (N_1494,N_804,N_737);
and U1495 (N_1495,N_235,N_889);
or U1496 (N_1496,N_618,N_101);
xnor U1497 (N_1497,N_586,N_613);
nand U1498 (N_1498,N_662,N_956);
and U1499 (N_1499,N_815,N_141);
and U1500 (N_1500,N_219,N_523);
or U1501 (N_1501,N_731,N_425);
nor U1502 (N_1502,N_540,N_414);
nand U1503 (N_1503,N_987,N_608);
nor U1504 (N_1504,N_390,N_256);
nand U1505 (N_1505,N_960,N_76);
nor U1506 (N_1506,N_742,N_94);
or U1507 (N_1507,N_34,N_710);
nor U1508 (N_1508,N_881,N_150);
and U1509 (N_1509,N_969,N_794);
nand U1510 (N_1510,N_994,N_513);
and U1511 (N_1511,N_611,N_171);
and U1512 (N_1512,N_926,N_899);
and U1513 (N_1513,N_564,N_892);
and U1514 (N_1514,N_234,N_157);
nand U1515 (N_1515,N_391,N_365);
nor U1516 (N_1516,N_421,N_859);
nand U1517 (N_1517,N_760,N_632);
nand U1518 (N_1518,N_796,N_96);
and U1519 (N_1519,N_98,N_321);
and U1520 (N_1520,N_701,N_235);
or U1521 (N_1521,N_971,N_878);
nand U1522 (N_1522,N_655,N_579);
nor U1523 (N_1523,N_795,N_816);
and U1524 (N_1524,N_719,N_563);
and U1525 (N_1525,N_356,N_134);
and U1526 (N_1526,N_549,N_961);
and U1527 (N_1527,N_101,N_368);
nand U1528 (N_1528,N_731,N_270);
and U1529 (N_1529,N_881,N_272);
or U1530 (N_1530,N_597,N_564);
xor U1531 (N_1531,N_13,N_99);
nor U1532 (N_1532,N_4,N_833);
nand U1533 (N_1533,N_305,N_48);
and U1534 (N_1534,N_778,N_505);
nand U1535 (N_1535,N_976,N_279);
nand U1536 (N_1536,N_981,N_928);
or U1537 (N_1537,N_926,N_445);
nand U1538 (N_1538,N_332,N_309);
and U1539 (N_1539,N_161,N_659);
nand U1540 (N_1540,N_733,N_308);
or U1541 (N_1541,N_58,N_118);
nand U1542 (N_1542,N_371,N_836);
and U1543 (N_1543,N_489,N_9);
nand U1544 (N_1544,N_403,N_100);
nor U1545 (N_1545,N_783,N_388);
nand U1546 (N_1546,N_622,N_786);
nand U1547 (N_1547,N_658,N_497);
or U1548 (N_1548,N_621,N_615);
and U1549 (N_1549,N_209,N_894);
nand U1550 (N_1550,N_627,N_226);
nand U1551 (N_1551,N_28,N_324);
or U1552 (N_1552,N_989,N_769);
and U1553 (N_1553,N_511,N_786);
or U1554 (N_1554,N_727,N_776);
or U1555 (N_1555,N_633,N_75);
or U1556 (N_1556,N_28,N_649);
nand U1557 (N_1557,N_841,N_409);
xor U1558 (N_1558,N_64,N_206);
or U1559 (N_1559,N_84,N_716);
or U1560 (N_1560,N_482,N_329);
nand U1561 (N_1561,N_193,N_258);
or U1562 (N_1562,N_460,N_366);
nor U1563 (N_1563,N_669,N_712);
nor U1564 (N_1564,N_710,N_97);
nor U1565 (N_1565,N_708,N_116);
or U1566 (N_1566,N_216,N_33);
or U1567 (N_1567,N_506,N_151);
and U1568 (N_1568,N_655,N_907);
nand U1569 (N_1569,N_648,N_78);
nor U1570 (N_1570,N_626,N_871);
nand U1571 (N_1571,N_60,N_816);
and U1572 (N_1572,N_47,N_579);
and U1573 (N_1573,N_620,N_263);
or U1574 (N_1574,N_434,N_226);
nor U1575 (N_1575,N_279,N_680);
nand U1576 (N_1576,N_849,N_263);
nor U1577 (N_1577,N_363,N_399);
nor U1578 (N_1578,N_45,N_945);
nor U1579 (N_1579,N_798,N_315);
or U1580 (N_1580,N_590,N_528);
and U1581 (N_1581,N_967,N_33);
and U1582 (N_1582,N_85,N_74);
nand U1583 (N_1583,N_620,N_676);
and U1584 (N_1584,N_733,N_242);
and U1585 (N_1585,N_27,N_684);
or U1586 (N_1586,N_623,N_713);
nand U1587 (N_1587,N_657,N_421);
nand U1588 (N_1588,N_170,N_406);
nand U1589 (N_1589,N_629,N_649);
and U1590 (N_1590,N_196,N_17);
nand U1591 (N_1591,N_637,N_403);
nand U1592 (N_1592,N_445,N_653);
or U1593 (N_1593,N_745,N_971);
nor U1594 (N_1594,N_428,N_985);
nor U1595 (N_1595,N_983,N_546);
nor U1596 (N_1596,N_692,N_947);
or U1597 (N_1597,N_281,N_826);
nor U1598 (N_1598,N_854,N_998);
nand U1599 (N_1599,N_802,N_402);
or U1600 (N_1600,N_56,N_130);
nor U1601 (N_1601,N_553,N_858);
or U1602 (N_1602,N_413,N_92);
nand U1603 (N_1603,N_131,N_676);
and U1604 (N_1604,N_334,N_930);
and U1605 (N_1605,N_526,N_251);
xnor U1606 (N_1606,N_527,N_259);
nand U1607 (N_1607,N_694,N_53);
nor U1608 (N_1608,N_812,N_601);
and U1609 (N_1609,N_636,N_967);
and U1610 (N_1610,N_699,N_623);
or U1611 (N_1611,N_342,N_661);
and U1612 (N_1612,N_643,N_756);
nand U1613 (N_1613,N_124,N_677);
nand U1614 (N_1614,N_764,N_423);
or U1615 (N_1615,N_704,N_656);
or U1616 (N_1616,N_697,N_703);
and U1617 (N_1617,N_987,N_821);
nand U1618 (N_1618,N_950,N_834);
or U1619 (N_1619,N_684,N_483);
nand U1620 (N_1620,N_710,N_815);
or U1621 (N_1621,N_754,N_250);
nand U1622 (N_1622,N_278,N_791);
nand U1623 (N_1623,N_904,N_690);
nand U1624 (N_1624,N_399,N_518);
or U1625 (N_1625,N_613,N_821);
nor U1626 (N_1626,N_915,N_205);
and U1627 (N_1627,N_776,N_713);
nand U1628 (N_1628,N_641,N_166);
and U1629 (N_1629,N_515,N_904);
nor U1630 (N_1630,N_827,N_450);
nand U1631 (N_1631,N_120,N_726);
nand U1632 (N_1632,N_759,N_915);
nand U1633 (N_1633,N_636,N_902);
and U1634 (N_1634,N_393,N_987);
xor U1635 (N_1635,N_92,N_988);
or U1636 (N_1636,N_495,N_704);
or U1637 (N_1637,N_979,N_209);
or U1638 (N_1638,N_716,N_633);
and U1639 (N_1639,N_47,N_789);
nand U1640 (N_1640,N_695,N_683);
or U1641 (N_1641,N_92,N_458);
nand U1642 (N_1642,N_8,N_849);
or U1643 (N_1643,N_844,N_501);
nor U1644 (N_1644,N_778,N_736);
nand U1645 (N_1645,N_507,N_430);
and U1646 (N_1646,N_940,N_275);
or U1647 (N_1647,N_651,N_561);
and U1648 (N_1648,N_80,N_840);
or U1649 (N_1649,N_315,N_490);
nor U1650 (N_1650,N_356,N_631);
nand U1651 (N_1651,N_10,N_48);
or U1652 (N_1652,N_235,N_308);
and U1653 (N_1653,N_958,N_808);
nand U1654 (N_1654,N_651,N_36);
or U1655 (N_1655,N_232,N_348);
nand U1656 (N_1656,N_836,N_933);
or U1657 (N_1657,N_244,N_219);
nand U1658 (N_1658,N_31,N_538);
or U1659 (N_1659,N_816,N_469);
nor U1660 (N_1660,N_59,N_566);
and U1661 (N_1661,N_21,N_81);
nand U1662 (N_1662,N_383,N_108);
nand U1663 (N_1663,N_374,N_847);
nand U1664 (N_1664,N_702,N_332);
nand U1665 (N_1665,N_64,N_70);
and U1666 (N_1666,N_684,N_693);
or U1667 (N_1667,N_785,N_880);
nand U1668 (N_1668,N_510,N_461);
or U1669 (N_1669,N_991,N_714);
nand U1670 (N_1670,N_937,N_896);
nand U1671 (N_1671,N_619,N_200);
and U1672 (N_1672,N_390,N_535);
nor U1673 (N_1673,N_322,N_98);
xnor U1674 (N_1674,N_471,N_72);
nand U1675 (N_1675,N_45,N_121);
and U1676 (N_1676,N_776,N_899);
nor U1677 (N_1677,N_598,N_972);
or U1678 (N_1678,N_283,N_399);
or U1679 (N_1679,N_349,N_33);
nor U1680 (N_1680,N_73,N_955);
nand U1681 (N_1681,N_488,N_39);
nor U1682 (N_1682,N_66,N_566);
and U1683 (N_1683,N_775,N_120);
nor U1684 (N_1684,N_485,N_357);
nor U1685 (N_1685,N_579,N_720);
nor U1686 (N_1686,N_268,N_614);
nand U1687 (N_1687,N_883,N_375);
and U1688 (N_1688,N_245,N_614);
nand U1689 (N_1689,N_985,N_169);
nand U1690 (N_1690,N_614,N_25);
nand U1691 (N_1691,N_881,N_238);
and U1692 (N_1692,N_839,N_423);
nor U1693 (N_1693,N_831,N_398);
or U1694 (N_1694,N_386,N_597);
nor U1695 (N_1695,N_377,N_974);
and U1696 (N_1696,N_320,N_29);
nor U1697 (N_1697,N_767,N_343);
or U1698 (N_1698,N_251,N_846);
or U1699 (N_1699,N_225,N_173);
or U1700 (N_1700,N_322,N_714);
or U1701 (N_1701,N_452,N_526);
nand U1702 (N_1702,N_14,N_956);
nor U1703 (N_1703,N_355,N_697);
nor U1704 (N_1704,N_149,N_782);
or U1705 (N_1705,N_57,N_686);
and U1706 (N_1706,N_716,N_809);
or U1707 (N_1707,N_19,N_617);
and U1708 (N_1708,N_3,N_694);
and U1709 (N_1709,N_54,N_867);
and U1710 (N_1710,N_923,N_965);
nand U1711 (N_1711,N_325,N_942);
nand U1712 (N_1712,N_861,N_269);
and U1713 (N_1713,N_374,N_617);
nand U1714 (N_1714,N_223,N_398);
nand U1715 (N_1715,N_382,N_328);
nand U1716 (N_1716,N_626,N_343);
and U1717 (N_1717,N_383,N_999);
or U1718 (N_1718,N_116,N_215);
or U1719 (N_1719,N_752,N_145);
or U1720 (N_1720,N_48,N_74);
nor U1721 (N_1721,N_751,N_496);
nor U1722 (N_1722,N_533,N_647);
and U1723 (N_1723,N_692,N_262);
or U1724 (N_1724,N_659,N_951);
nor U1725 (N_1725,N_643,N_34);
nand U1726 (N_1726,N_581,N_197);
nand U1727 (N_1727,N_789,N_669);
nand U1728 (N_1728,N_567,N_488);
and U1729 (N_1729,N_92,N_51);
or U1730 (N_1730,N_798,N_880);
and U1731 (N_1731,N_741,N_198);
and U1732 (N_1732,N_499,N_535);
nand U1733 (N_1733,N_59,N_821);
or U1734 (N_1734,N_939,N_954);
nor U1735 (N_1735,N_232,N_165);
nand U1736 (N_1736,N_387,N_830);
or U1737 (N_1737,N_389,N_99);
nand U1738 (N_1738,N_318,N_328);
and U1739 (N_1739,N_46,N_996);
or U1740 (N_1740,N_48,N_729);
or U1741 (N_1741,N_391,N_705);
and U1742 (N_1742,N_683,N_181);
or U1743 (N_1743,N_138,N_316);
or U1744 (N_1744,N_667,N_195);
nor U1745 (N_1745,N_688,N_104);
nand U1746 (N_1746,N_533,N_601);
nand U1747 (N_1747,N_942,N_37);
nand U1748 (N_1748,N_932,N_777);
or U1749 (N_1749,N_424,N_713);
or U1750 (N_1750,N_632,N_800);
nand U1751 (N_1751,N_630,N_67);
and U1752 (N_1752,N_557,N_987);
or U1753 (N_1753,N_188,N_257);
or U1754 (N_1754,N_565,N_961);
or U1755 (N_1755,N_33,N_991);
nor U1756 (N_1756,N_250,N_283);
nand U1757 (N_1757,N_55,N_552);
nor U1758 (N_1758,N_808,N_292);
nand U1759 (N_1759,N_32,N_723);
nand U1760 (N_1760,N_25,N_592);
nand U1761 (N_1761,N_755,N_411);
or U1762 (N_1762,N_76,N_394);
nand U1763 (N_1763,N_926,N_7);
nand U1764 (N_1764,N_709,N_367);
nand U1765 (N_1765,N_726,N_235);
nor U1766 (N_1766,N_797,N_165);
or U1767 (N_1767,N_960,N_899);
and U1768 (N_1768,N_821,N_714);
nand U1769 (N_1769,N_44,N_131);
and U1770 (N_1770,N_699,N_327);
or U1771 (N_1771,N_844,N_169);
nor U1772 (N_1772,N_573,N_142);
nand U1773 (N_1773,N_889,N_15);
nor U1774 (N_1774,N_651,N_256);
xnor U1775 (N_1775,N_847,N_10);
nand U1776 (N_1776,N_939,N_934);
and U1777 (N_1777,N_213,N_118);
nand U1778 (N_1778,N_113,N_147);
nor U1779 (N_1779,N_353,N_634);
nor U1780 (N_1780,N_651,N_465);
nand U1781 (N_1781,N_584,N_725);
nand U1782 (N_1782,N_636,N_371);
and U1783 (N_1783,N_704,N_725);
and U1784 (N_1784,N_536,N_248);
and U1785 (N_1785,N_974,N_534);
nand U1786 (N_1786,N_274,N_289);
and U1787 (N_1787,N_186,N_78);
and U1788 (N_1788,N_905,N_917);
nor U1789 (N_1789,N_950,N_383);
and U1790 (N_1790,N_5,N_869);
nand U1791 (N_1791,N_235,N_206);
nor U1792 (N_1792,N_253,N_747);
and U1793 (N_1793,N_261,N_213);
nand U1794 (N_1794,N_436,N_280);
or U1795 (N_1795,N_964,N_94);
nor U1796 (N_1796,N_673,N_422);
and U1797 (N_1797,N_229,N_672);
or U1798 (N_1798,N_872,N_319);
xnor U1799 (N_1799,N_635,N_464);
nor U1800 (N_1800,N_375,N_664);
nand U1801 (N_1801,N_829,N_126);
and U1802 (N_1802,N_884,N_668);
and U1803 (N_1803,N_713,N_974);
nand U1804 (N_1804,N_966,N_460);
nor U1805 (N_1805,N_452,N_439);
nand U1806 (N_1806,N_452,N_398);
and U1807 (N_1807,N_723,N_794);
nand U1808 (N_1808,N_602,N_211);
or U1809 (N_1809,N_140,N_719);
nand U1810 (N_1810,N_326,N_673);
and U1811 (N_1811,N_498,N_837);
nor U1812 (N_1812,N_240,N_714);
and U1813 (N_1813,N_316,N_253);
and U1814 (N_1814,N_653,N_329);
or U1815 (N_1815,N_511,N_795);
and U1816 (N_1816,N_990,N_265);
nor U1817 (N_1817,N_528,N_715);
nor U1818 (N_1818,N_868,N_493);
or U1819 (N_1819,N_262,N_163);
nor U1820 (N_1820,N_613,N_250);
and U1821 (N_1821,N_286,N_56);
and U1822 (N_1822,N_898,N_673);
nand U1823 (N_1823,N_676,N_151);
nand U1824 (N_1824,N_324,N_701);
nor U1825 (N_1825,N_332,N_839);
nor U1826 (N_1826,N_128,N_413);
nor U1827 (N_1827,N_193,N_822);
nor U1828 (N_1828,N_990,N_118);
and U1829 (N_1829,N_162,N_430);
and U1830 (N_1830,N_255,N_276);
nand U1831 (N_1831,N_134,N_656);
nor U1832 (N_1832,N_872,N_967);
or U1833 (N_1833,N_891,N_497);
and U1834 (N_1834,N_676,N_67);
and U1835 (N_1835,N_622,N_486);
nor U1836 (N_1836,N_648,N_983);
nor U1837 (N_1837,N_263,N_531);
or U1838 (N_1838,N_843,N_565);
and U1839 (N_1839,N_465,N_604);
nor U1840 (N_1840,N_973,N_83);
and U1841 (N_1841,N_894,N_314);
or U1842 (N_1842,N_635,N_625);
nor U1843 (N_1843,N_498,N_0);
nand U1844 (N_1844,N_483,N_687);
and U1845 (N_1845,N_849,N_867);
nor U1846 (N_1846,N_767,N_30);
nand U1847 (N_1847,N_48,N_324);
or U1848 (N_1848,N_918,N_340);
nor U1849 (N_1849,N_626,N_346);
nand U1850 (N_1850,N_762,N_727);
and U1851 (N_1851,N_316,N_566);
or U1852 (N_1852,N_828,N_930);
nor U1853 (N_1853,N_765,N_758);
nor U1854 (N_1854,N_653,N_110);
and U1855 (N_1855,N_738,N_975);
or U1856 (N_1856,N_161,N_376);
and U1857 (N_1857,N_823,N_609);
nand U1858 (N_1858,N_72,N_538);
nor U1859 (N_1859,N_528,N_271);
nor U1860 (N_1860,N_356,N_733);
and U1861 (N_1861,N_349,N_684);
and U1862 (N_1862,N_439,N_250);
and U1863 (N_1863,N_554,N_110);
or U1864 (N_1864,N_153,N_870);
and U1865 (N_1865,N_952,N_775);
or U1866 (N_1866,N_960,N_89);
xor U1867 (N_1867,N_923,N_503);
nand U1868 (N_1868,N_968,N_138);
nand U1869 (N_1869,N_556,N_101);
nor U1870 (N_1870,N_596,N_387);
and U1871 (N_1871,N_860,N_74);
nor U1872 (N_1872,N_619,N_695);
and U1873 (N_1873,N_631,N_492);
or U1874 (N_1874,N_760,N_909);
and U1875 (N_1875,N_23,N_489);
nand U1876 (N_1876,N_617,N_763);
and U1877 (N_1877,N_516,N_90);
and U1878 (N_1878,N_881,N_752);
or U1879 (N_1879,N_938,N_46);
and U1880 (N_1880,N_351,N_139);
and U1881 (N_1881,N_165,N_351);
or U1882 (N_1882,N_887,N_148);
nand U1883 (N_1883,N_154,N_395);
nand U1884 (N_1884,N_893,N_503);
or U1885 (N_1885,N_383,N_179);
or U1886 (N_1886,N_229,N_978);
nor U1887 (N_1887,N_419,N_668);
nor U1888 (N_1888,N_579,N_562);
nor U1889 (N_1889,N_321,N_70);
and U1890 (N_1890,N_612,N_650);
nor U1891 (N_1891,N_972,N_744);
nand U1892 (N_1892,N_772,N_824);
nand U1893 (N_1893,N_890,N_606);
xnor U1894 (N_1894,N_679,N_36);
nor U1895 (N_1895,N_55,N_298);
or U1896 (N_1896,N_914,N_682);
nor U1897 (N_1897,N_58,N_830);
nand U1898 (N_1898,N_622,N_372);
and U1899 (N_1899,N_22,N_487);
and U1900 (N_1900,N_423,N_197);
nor U1901 (N_1901,N_288,N_26);
and U1902 (N_1902,N_535,N_717);
or U1903 (N_1903,N_739,N_781);
nor U1904 (N_1904,N_601,N_933);
nor U1905 (N_1905,N_452,N_166);
or U1906 (N_1906,N_2,N_307);
nor U1907 (N_1907,N_286,N_582);
or U1908 (N_1908,N_536,N_552);
xor U1909 (N_1909,N_652,N_664);
or U1910 (N_1910,N_347,N_573);
nor U1911 (N_1911,N_670,N_586);
and U1912 (N_1912,N_127,N_864);
nand U1913 (N_1913,N_978,N_75);
or U1914 (N_1914,N_556,N_767);
and U1915 (N_1915,N_244,N_208);
nand U1916 (N_1916,N_555,N_457);
nand U1917 (N_1917,N_347,N_203);
and U1918 (N_1918,N_537,N_588);
nor U1919 (N_1919,N_215,N_135);
nor U1920 (N_1920,N_130,N_298);
nand U1921 (N_1921,N_450,N_956);
and U1922 (N_1922,N_435,N_906);
and U1923 (N_1923,N_213,N_135);
and U1924 (N_1924,N_995,N_377);
and U1925 (N_1925,N_133,N_758);
or U1926 (N_1926,N_252,N_797);
or U1927 (N_1927,N_762,N_172);
and U1928 (N_1928,N_914,N_887);
or U1929 (N_1929,N_863,N_564);
or U1930 (N_1930,N_635,N_795);
nand U1931 (N_1931,N_464,N_815);
or U1932 (N_1932,N_47,N_600);
nor U1933 (N_1933,N_257,N_287);
or U1934 (N_1934,N_953,N_376);
nand U1935 (N_1935,N_328,N_733);
or U1936 (N_1936,N_63,N_837);
and U1937 (N_1937,N_927,N_97);
or U1938 (N_1938,N_355,N_887);
and U1939 (N_1939,N_517,N_36);
nor U1940 (N_1940,N_59,N_591);
nor U1941 (N_1941,N_872,N_293);
or U1942 (N_1942,N_376,N_832);
nand U1943 (N_1943,N_353,N_551);
and U1944 (N_1944,N_928,N_536);
nor U1945 (N_1945,N_399,N_145);
nand U1946 (N_1946,N_458,N_735);
nand U1947 (N_1947,N_54,N_960);
nor U1948 (N_1948,N_536,N_235);
nand U1949 (N_1949,N_363,N_703);
nand U1950 (N_1950,N_851,N_497);
nand U1951 (N_1951,N_163,N_497);
nand U1952 (N_1952,N_848,N_245);
and U1953 (N_1953,N_461,N_422);
and U1954 (N_1954,N_54,N_139);
and U1955 (N_1955,N_820,N_984);
or U1956 (N_1956,N_351,N_462);
nor U1957 (N_1957,N_558,N_409);
and U1958 (N_1958,N_196,N_739);
and U1959 (N_1959,N_110,N_101);
and U1960 (N_1960,N_944,N_20);
nand U1961 (N_1961,N_657,N_828);
nand U1962 (N_1962,N_462,N_974);
and U1963 (N_1963,N_979,N_103);
or U1964 (N_1964,N_627,N_747);
and U1965 (N_1965,N_461,N_220);
or U1966 (N_1966,N_438,N_271);
or U1967 (N_1967,N_855,N_4);
nand U1968 (N_1968,N_323,N_951);
nand U1969 (N_1969,N_749,N_249);
and U1970 (N_1970,N_566,N_967);
nand U1971 (N_1971,N_921,N_673);
nor U1972 (N_1972,N_950,N_83);
or U1973 (N_1973,N_679,N_24);
or U1974 (N_1974,N_805,N_845);
nand U1975 (N_1975,N_817,N_995);
nor U1976 (N_1976,N_901,N_453);
and U1977 (N_1977,N_467,N_706);
nor U1978 (N_1978,N_581,N_647);
and U1979 (N_1979,N_852,N_23);
and U1980 (N_1980,N_516,N_75);
or U1981 (N_1981,N_391,N_407);
nand U1982 (N_1982,N_974,N_932);
or U1983 (N_1983,N_789,N_846);
or U1984 (N_1984,N_46,N_475);
nor U1985 (N_1985,N_916,N_865);
nand U1986 (N_1986,N_702,N_330);
nor U1987 (N_1987,N_991,N_526);
nand U1988 (N_1988,N_867,N_283);
or U1989 (N_1989,N_84,N_934);
nor U1990 (N_1990,N_527,N_387);
and U1991 (N_1991,N_443,N_466);
nor U1992 (N_1992,N_430,N_98);
and U1993 (N_1993,N_15,N_306);
or U1994 (N_1994,N_143,N_717);
nor U1995 (N_1995,N_312,N_940);
nand U1996 (N_1996,N_392,N_597);
nand U1997 (N_1997,N_43,N_496);
or U1998 (N_1998,N_663,N_497);
and U1999 (N_1999,N_995,N_721);
or U2000 (N_2000,N_1330,N_1618);
nor U2001 (N_2001,N_1572,N_1884);
xnor U2002 (N_2002,N_1526,N_1363);
and U2003 (N_2003,N_1491,N_1786);
nor U2004 (N_2004,N_1167,N_1084);
and U2005 (N_2005,N_1683,N_1818);
or U2006 (N_2006,N_1647,N_1894);
and U2007 (N_2007,N_1944,N_1510);
nor U2008 (N_2008,N_1761,N_1632);
xor U2009 (N_2009,N_1591,N_1223);
and U2010 (N_2010,N_1551,N_1154);
nor U2011 (N_2011,N_1738,N_1441);
nand U2012 (N_2012,N_1583,N_1875);
and U2013 (N_2013,N_1061,N_1197);
and U2014 (N_2014,N_1085,N_1984);
or U2015 (N_2015,N_1582,N_1982);
or U2016 (N_2016,N_1043,N_1711);
and U2017 (N_2017,N_1566,N_1764);
nor U2018 (N_2018,N_1854,N_1871);
and U2019 (N_2019,N_1055,N_1671);
or U2020 (N_2020,N_1012,N_1290);
and U2021 (N_2021,N_1292,N_1958);
and U2022 (N_2022,N_1258,N_1262);
nand U2023 (N_2023,N_1817,N_1476);
and U2024 (N_2024,N_1345,N_1421);
and U2025 (N_2025,N_1568,N_1864);
or U2026 (N_2026,N_1843,N_1614);
or U2027 (N_2027,N_1321,N_1237);
and U2028 (N_2028,N_1598,N_1781);
nor U2029 (N_2029,N_1298,N_1631);
nand U2030 (N_2030,N_1256,N_1992);
or U2031 (N_2031,N_1521,N_1682);
or U2032 (N_2032,N_1747,N_1800);
and U2033 (N_2033,N_1619,N_1293);
nor U2034 (N_2034,N_1855,N_1266);
or U2035 (N_2035,N_1165,N_1436);
and U2036 (N_2036,N_1932,N_1807);
and U2037 (N_2037,N_1606,N_1597);
or U2038 (N_2038,N_1703,N_1594);
nand U2039 (N_2039,N_1219,N_1644);
or U2040 (N_2040,N_1229,N_1208);
nor U2041 (N_2041,N_1525,N_1959);
or U2042 (N_2042,N_1556,N_1672);
nand U2043 (N_2043,N_1286,N_1744);
or U2044 (N_2044,N_1546,N_1075);
nand U2045 (N_2045,N_1387,N_1138);
nand U2046 (N_2046,N_1700,N_1479);
nand U2047 (N_2047,N_1039,N_1748);
nand U2048 (N_2048,N_1078,N_1726);
nor U2049 (N_2049,N_1485,N_1600);
nor U2050 (N_2050,N_1089,N_1163);
nand U2051 (N_2051,N_1770,N_1202);
xnor U2052 (N_2052,N_1396,N_1009);
or U2053 (N_2053,N_1327,N_1230);
nand U2054 (N_2054,N_1889,N_1112);
and U2055 (N_2055,N_1377,N_1863);
and U2056 (N_2056,N_1390,N_1979);
nand U2057 (N_2057,N_1697,N_1642);
or U2058 (N_2058,N_1414,N_1814);
and U2059 (N_2059,N_1067,N_1501);
or U2060 (N_2060,N_1406,N_1140);
nor U2061 (N_2061,N_1692,N_1657);
nor U2062 (N_2062,N_1563,N_1333);
or U2063 (N_2063,N_1402,N_1175);
or U2064 (N_2064,N_1472,N_1561);
or U2065 (N_2065,N_1985,N_1769);
or U2066 (N_2066,N_1896,N_1852);
nand U2067 (N_2067,N_1799,N_1082);
nor U2068 (N_2068,N_1560,N_1385);
or U2069 (N_2069,N_1162,N_1830);
nand U2070 (N_2070,N_1821,N_1735);
or U2071 (N_2071,N_1339,N_1802);
nand U2072 (N_2072,N_1059,N_1617);
nand U2073 (N_2073,N_1113,N_1437);
nor U2074 (N_2074,N_1119,N_1869);
or U2075 (N_2075,N_1831,N_1122);
nor U2076 (N_2076,N_1433,N_1260);
and U2077 (N_2077,N_1776,N_1705);
and U2078 (N_2078,N_1498,N_1372);
and U2079 (N_2079,N_1530,N_1307);
or U2080 (N_2080,N_1135,N_1584);
nor U2081 (N_2081,N_1648,N_1495);
nand U2082 (N_2082,N_1411,N_1684);
and U2083 (N_2083,N_1531,N_1562);
nand U2084 (N_2084,N_1173,N_1544);
and U2085 (N_2085,N_1473,N_1709);
or U2086 (N_2086,N_1021,N_1366);
or U2087 (N_2087,N_1997,N_1289);
or U2088 (N_2088,N_1767,N_1487);
nor U2089 (N_2089,N_1971,N_1376);
or U2090 (N_2090,N_1282,N_1742);
or U2091 (N_2091,N_1034,N_1909);
and U2092 (N_2092,N_1936,N_1028);
and U2093 (N_2093,N_1987,N_1212);
nor U2094 (N_2094,N_1353,N_1659);
or U2095 (N_2095,N_1465,N_1835);
nor U2096 (N_2096,N_1636,N_1284);
or U2097 (N_2097,N_1225,N_1215);
or U2098 (N_2098,N_1295,N_1183);
and U2099 (N_2099,N_1677,N_1155);
and U2100 (N_2100,N_1630,N_1558);
nor U2101 (N_2101,N_1731,N_1823);
nand U2102 (N_2102,N_1877,N_1840);
or U2103 (N_2103,N_1706,N_1620);
nand U2104 (N_2104,N_1027,N_1952);
nor U2105 (N_2105,N_1277,N_1837);
and U2106 (N_2106,N_1470,N_1270);
or U2107 (N_2107,N_1693,N_1740);
or U2108 (N_2108,N_1719,N_1131);
nor U2109 (N_2109,N_1115,N_1464);
nor U2110 (N_2110,N_1751,N_1056);
or U2111 (N_2111,N_1188,N_1991);
and U2112 (N_2112,N_1458,N_1246);
nor U2113 (N_2113,N_1279,N_1535);
nor U2114 (N_2114,N_1036,N_1542);
nand U2115 (N_2115,N_1453,N_1809);
and U2116 (N_2116,N_1904,N_1204);
nor U2117 (N_2117,N_1862,N_1086);
or U2118 (N_2118,N_1650,N_1434);
and U2119 (N_2119,N_1592,N_1319);
nor U2120 (N_2120,N_1189,N_1910);
nand U2121 (N_2121,N_1722,N_1841);
nand U2122 (N_2122,N_1996,N_1502);
nand U2123 (N_2123,N_1026,N_1793);
and U2124 (N_2124,N_1420,N_1364);
nand U2125 (N_2125,N_1765,N_1373);
and U2126 (N_2126,N_1815,N_1870);
nand U2127 (N_2127,N_1859,N_1294);
nand U2128 (N_2128,N_1497,N_1152);
nand U2129 (N_2129,N_1834,N_1418);
nor U2130 (N_2130,N_1348,N_1271);
and U2131 (N_2131,N_1861,N_1973);
and U2132 (N_2132,N_1788,N_1475);
nand U2133 (N_2133,N_1346,N_1024);
nor U2134 (N_2134,N_1371,N_1181);
nor U2135 (N_2135,N_1161,N_1916);
nand U2136 (N_2136,N_1132,N_1342);
nor U2137 (N_2137,N_1231,N_1431);
nor U2138 (N_2138,N_1578,N_1391);
nor U2139 (N_2139,N_1574,N_1825);
xnor U2140 (N_2140,N_1045,N_1389);
nand U2141 (N_2141,N_1914,N_1314);
or U2142 (N_2142,N_1281,N_1969);
nand U2143 (N_2143,N_1448,N_1020);
and U2144 (N_2144,N_1964,N_1865);
and U2145 (N_2145,N_1579,N_1961);
nor U2146 (N_2146,N_1176,N_1370);
nor U2147 (N_2147,N_1536,N_1882);
nor U2148 (N_2148,N_1790,N_1570);
or U2149 (N_2149,N_1892,N_1276);
nor U2150 (N_2150,N_1867,N_1095);
nand U2151 (N_2151,N_1068,N_1357);
nor U2152 (N_2152,N_1496,N_1939);
and U2153 (N_2153,N_1557,N_1733);
and U2154 (N_2154,N_1477,N_1957);
nand U2155 (N_2155,N_1766,N_1949);
and U2156 (N_2156,N_1750,N_1419);
xor U2157 (N_2157,N_1812,N_1567);
and U2158 (N_2158,N_1729,N_1233);
and U2159 (N_2159,N_1104,N_1743);
or U2160 (N_2160,N_1447,N_1927);
nand U2161 (N_2161,N_1918,N_1349);
or U2162 (N_2162,N_1395,N_1160);
and U2163 (N_2163,N_1407,N_1891);
nor U2164 (N_2164,N_1273,N_1232);
nor U2165 (N_2165,N_1948,N_1552);
nand U2166 (N_2166,N_1305,N_1621);
xnor U2167 (N_2167,N_1199,N_1783);
xor U2168 (N_2168,N_1652,N_1950);
nor U2169 (N_2169,N_1780,N_1895);
and U2170 (N_2170,N_1879,N_1885);
or U2171 (N_2171,N_1569,N_1446);
nor U2172 (N_2172,N_1032,N_1111);
xnor U2173 (N_2173,N_1150,N_1674);
and U2174 (N_2174,N_1325,N_1080);
nand U2175 (N_2175,N_1207,N_1773);
nor U2176 (N_2176,N_1604,N_1253);
and U2177 (N_2177,N_1749,N_1300);
nand U2178 (N_2178,N_1678,N_1608);
or U2179 (N_2179,N_1438,N_1216);
nor U2180 (N_2180,N_1670,N_1611);
and U2181 (N_2181,N_1509,N_1966);
nor U2182 (N_2182,N_1141,N_1541);
and U2183 (N_2183,N_1179,N_1934);
nor U2184 (N_2184,N_1585,N_1940);
and U2185 (N_2185,N_1782,N_1655);
and U2186 (N_2186,N_1635,N_1710);
nor U2187 (N_2187,N_1388,N_1715);
nor U2188 (N_2188,N_1013,N_1172);
and U2189 (N_2189,N_1022,N_1239);
and U2190 (N_2190,N_1323,N_1873);
and U2191 (N_2191,N_1913,N_1928);
nand U2192 (N_2192,N_1259,N_1439);
and U2193 (N_2193,N_1845,N_1504);
and U2194 (N_2194,N_1739,N_1299);
nor U2195 (N_2195,N_1519,N_1356);
nor U2196 (N_2196,N_1527,N_1899);
and U2197 (N_2197,N_1986,N_1951);
and U2198 (N_2198,N_1397,N_1915);
nor U2199 (N_2199,N_1716,N_1368);
nand U2200 (N_2200,N_1425,N_1275);
nor U2201 (N_2201,N_1053,N_1079);
and U2202 (N_2202,N_1014,N_1577);
or U2203 (N_2203,N_1432,N_1900);
xnor U2204 (N_2204,N_1144,N_1538);
and U2205 (N_2205,N_1129,N_1060);
or U2206 (N_2206,N_1901,N_1886);
nand U2207 (N_2207,N_1178,N_1746);
nor U2208 (N_2208,N_1675,N_1593);
nand U2209 (N_2209,N_1745,N_1412);
nor U2210 (N_2210,N_1603,N_1435);
nor U2211 (N_2211,N_1763,N_1283);
nand U2212 (N_2212,N_1306,N_1123);
nand U2213 (N_2213,N_1947,N_1444);
and U2214 (N_2214,N_1004,N_1555);
nand U2215 (N_2215,N_1313,N_1251);
nand U2216 (N_2216,N_1303,N_1250);
nand U2217 (N_2217,N_1590,N_1203);
or U2218 (N_2218,N_1627,N_1072);
nand U2219 (N_2219,N_1147,N_1404);
nand U2220 (N_2220,N_1532,N_1827);
or U2221 (N_2221,N_1860,N_1789);
xnor U2222 (N_2222,N_1310,N_1774);
and U2223 (N_2223,N_1066,N_1797);
nand U2224 (N_2224,N_1628,N_1226);
nor U2225 (N_2225,N_1117,N_1813);
nand U2226 (N_2226,N_1816,N_1828);
nor U2227 (N_2227,N_1576,N_1999);
nand U2228 (N_2228,N_1088,N_1515);
nand U2229 (N_2229,N_1461,N_1938);
nand U2230 (N_2230,N_1320,N_1553);
and U2231 (N_2231,N_1101,N_1685);
and U2232 (N_2232,N_1044,N_1097);
nor U2233 (N_2233,N_1612,N_1006);
and U2234 (N_2234,N_1480,N_1268);
nand U2235 (N_2235,N_1015,N_1272);
nor U2236 (N_2236,N_1960,N_1702);
and U2237 (N_2237,N_1919,N_1931);
nor U2238 (N_2238,N_1695,N_1634);
nor U2239 (N_2239,N_1484,N_1309);
nand U2240 (N_2240,N_1826,N_1010);
and U2241 (N_2241,N_1824,N_1287);
nor U2242 (N_2242,N_1070,N_1549);
or U2243 (N_2243,N_1409,N_1609);
or U2244 (N_2244,N_1090,N_1267);
or U2245 (N_2245,N_1925,N_1661);
or U2246 (N_2246,N_1482,N_1633);
or U2247 (N_2247,N_1350,N_1369);
and U2248 (N_2248,N_1533,N_1545);
or U2249 (N_2249,N_1898,N_1847);
nor U2250 (N_2250,N_1164,N_1317);
nand U2251 (N_2251,N_1408,N_1174);
nor U2252 (N_2252,N_1029,N_1694);
or U2253 (N_2253,N_1137,N_1980);
nand U2254 (N_2254,N_1429,N_1220);
or U2255 (N_2255,N_1354,N_1008);
nor U2256 (N_2256,N_1466,N_1049);
xnor U2257 (N_2257,N_1128,N_1981);
nor U2258 (N_2258,N_1255,N_1322);
and U2259 (N_2259,N_1427,N_1696);
and U2260 (N_2260,N_1838,N_1708);
nand U2261 (N_2261,N_1778,N_1588);
and U2262 (N_2262,N_1933,N_1505);
nand U2263 (N_2263,N_1822,N_1937);
nand U2264 (N_2264,N_1868,N_1146);
nor U2265 (N_2265,N_1265,N_1063);
nor U2266 (N_2266,N_1062,N_1798);
or U2267 (N_2267,N_1639,N_1094);
or U2268 (N_2268,N_1426,N_1905);
or U2269 (N_2269,N_1157,N_1967);
nand U2270 (N_2270,N_1721,N_1848);
and U2271 (N_2271,N_1196,N_1185);
or U2272 (N_2272,N_1153,N_1662);
nand U2273 (N_2273,N_1849,N_1151);
xnor U2274 (N_2274,N_1550,N_1236);
and U2275 (N_2275,N_1503,N_1732);
nor U2276 (N_2276,N_1471,N_1478);
and U2277 (N_2277,N_1454,N_1511);
nand U2278 (N_2278,N_1098,N_1423);
and U2279 (N_2279,N_1280,N_1442);
nand U2280 (N_2280,N_1954,N_1872);
nand U2281 (N_2281,N_1416,N_1539);
nand U2282 (N_2282,N_1341,N_1819);
or U2283 (N_2283,N_1083,N_1945);
nor U2284 (N_2284,N_1752,N_1336);
nand U2285 (N_2285,N_1888,N_1707);
and U2286 (N_2286,N_1074,N_1589);
nor U2287 (N_2287,N_1263,N_1058);
nand U2288 (N_2288,N_1194,N_1398);
nand U2289 (N_2289,N_1463,N_1110);
and U2290 (N_2290,N_1712,N_1076);
and U2291 (N_2291,N_1126,N_1071);
nor U2292 (N_2292,N_1332,N_1520);
nand U2293 (N_2293,N_1205,N_1718);
nand U2294 (N_2294,N_1874,N_1069);
nor U2295 (N_2295,N_1785,N_1836);
xnor U2296 (N_2296,N_1170,N_1252);
or U2297 (N_2297,N_1244,N_1638);
or U2298 (N_2298,N_1688,N_1492);
nand U2299 (N_2299,N_1955,N_1379);
or U2300 (N_2300,N_1134,N_1775);
or U2301 (N_2301,N_1610,N_1018);
nand U2302 (N_2302,N_1177,N_1459);
nand U2303 (N_2303,N_1974,N_1308);
nor U2304 (N_2304,N_1073,N_1846);
and U2305 (N_2305,N_1548,N_1092);
or U2306 (N_2306,N_1665,N_1613);
and U2307 (N_2307,N_1316,N_1842);
and U2308 (N_2308,N_1963,N_1374);
and U2309 (N_2309,N_1663,N_1238);
xor U2310 (N_2310,N_1030,N_1607);
nor U2311 (N_2311,N_1881,N_1400);
nor U2312 (N_2312,N_1640,N_1221);
and U2313 (N_2313,N_1003,N_1329);
xor U2314 (N_2314,N_1360,N_1965);
and U2315 (N_2315,N_1096,N_1344);
and U2316 (N_2316,N_1359,N_1756);
nor U2317 (N_2317,N_1362,N_1288);
or U2318 (N_2318,N_1235,N_1523);
nor U2319 (N_2319,N_1201,N_1048);
nor U2320 (N_2320,N_1540,N_1615);
nor U2321 (N_2321,N_1646,N_1093);
nor U2322 (N_2322,N_1334,N_1133);
or U2323 (N_2323,N_1832,N_1565);
or U2324 (N_2324,N_1143,N_1499);
and U2325 (N_2325,N_1649,N_1488);
nand U2326 (N_2326,N_1581,N_1956);
nor U2327 (N_2327,N_1656,N_1392);
nand U2328 (N_2328,N_1077,N_1573);
or U2329 (N_2329,N_1210,N_1033);
or U2330 (N_2330,N_1187,N_1587);
or U2331 (N_2331,N_1990,N_1804);
or U2332 (N_2332,N_1720,N_1717);
nand U2333 (N_2333,N_1050,N_1792);
nor U2334 (N_2334,N_1978,N_1193);
nor U2335 (N_2335,N_1559,N_1537);
nor U2336 (N_2336,N_1213,N_1120);
nor U2337 (N_2337,N_1035,N_1124);
nand U2338 (N_2338,N_1791,N_1462);
and U2339 (N_2339,N_1669,N_1424);
nor U2340 (N_2340,N_1468,N_1757);
or U2341 (N_2341,N_1031,N_1218);
or U2342 (N_2342,N_1993,N_1002);
nand U2343 (N_2343,N_1257,N_1728);
and U2344 (N_2344,N_1217,N_1803);
and U2345 (N_2345,N_1626,N_1241);
nor U2346 (N_2346,N_1857,N_1820);
nand U2347 (N_2347,N_1844,N_1771);
nor U2348 (N_2348,N_1211,N_1347);
and U2349 (N_2349,N_1629,N_1358);
nand U2350 (N_2350,N_1460,N_1736);
nand U2351 (N_2351,N_1668,N_1243);
and U2352 (N_2352,N_1651,N_1943);
or U2353 (N_2353,N_1930,N_1254);
xor U2354 (N_2354,N_1428,N_1839);
or U2355 (N_2355,N_1352,N_1806);
or U2356 (N_2356,N_1942,N_1302);
and U2357 (N_2357,N_1099,N_1109);
nand U2358 (N_2358,N_1195,N_1890);
nor U2359 (N_2359,N_1810,N_1198);
nand U2360 (N_2360,N_1601,N_1517);
nand U2361 (N_2361,N_1393,N_1328);
or U2362 (N_2362,N_1946,N_1474);
and U2363 (N_2363,N_1929,N_1417);
or U2364 (N_2364,N_1616,N_1041);
nand U2365 (N_2365,N_1228,N_1312);
and U2366 (N_2366,N_1000,N_1676);
and U2367 (N_2367,N_1318,N_1121);
nor U2368 (N_2368,N_1064,N_1403);
or U2369 (N_2369,N_1486,N_1159);
or U2370 (N_2370,N_1249,N_1725);
and U2371 (N_2371,N_1191,N_1297);
xnor U2372 (N_2372,N_1456,N_1394);
and U2373 (N_2373,N_1142,N_1779);
or U2374 (N_2374,N_1580,N_1169);
nor U2375 (N_2375,N_1730,N_1483);
and U2376 (N_2376,N_1017,N_1528);
and U2377 (N_2377,N_1941,N_1087);
and U2378 (N_2378,N_1443,N_1543);
or U2379 (N_2379,N_1125,N_1880);
or U2380 (N_2380,N_1508,N_1759);
and U2381 (N_2381,N_1851,N_1554);
nor U2382 (N_2382,N_1924,N_1200);
and U2383 (N_2383,N_1186,N_1304);
nor U2384 (N_2384,N_1724,N_1047);
or U2385 (N_2385,N_1575,N_1701);
and U2386 (N_2386,N_1489,N_1382);
or U2387 (N_2387,N_1968,N_1641);
nor U2388 (N_2388,N_1415,N_1274);
or U2389 (N_2389,N_1547,N_1469);
and U2390 (N_2390,N_1777,N_1833);
and U2391 (N_2391,N_1762,N_1737);
or U2392 (N_2392,N_1261,N_1184);
nor U2393 (N_2393,N_1787,N_1315);
nor U2394 (N_2394,N_1908,N_1296);
nor U2395 (N_2395,N_1052,N_1689);
or U2396 (N_2396,N_1324,N_1768);
nor U2397 (N_2397,N_1139,N_1935);
nor U2398 (N_2398,N_1168,N_1240);
or U2399 (N_2399,N_1953,N_1977);
nor U2400 (N_2400,N_1516,N_1989);
nand U2401 (N_2401,N_1326,N_1493);
and U2402 (N_2402,N_1445,N_1923);
nand U2403 (N_2403,N_1269,N_1224);
and U2404 (N_2404,N_1921,N_1887);
nor U2405 (N_2405,N_1522,N_1680);
nand U2406 (N_2406,N_1007,N_1534);
nor U2407 (N_2407,N_1926,N_1666);
and U2408 (N_2408,N_1422,N_1754);
nand U2409 (N_2409,N_1383,N_1698);
or U2410 (N_2410,N_1658,N_1149);
nor U2411 (N_2411,N_1405,N_1451);
or U2412 (N_2412,N_1214,N_1970);
nand U2413 (N_2413,N_1381,N_1166);
and U2414 (N_2414,N_1449,N_1040);
nor U2415 (N_2415,N_1513,N_1512);
nor U2416 (N_2416,N_1107,N_1679);
nand U2417 (N_2417,N_1625,N_1467);
nand U2418 (N_2418,N_1912,N_1983);
nor U2419 (N_2419,N_1922,N_1903);
and U2420 (N_2420,N_1876,N_1758);
nor U2421 (N_2421,N_1660,N_1452);
and U2422 (N_2422,N_1065,N_1386);
and U2423 (N_2423,N_1667,N_1005);
or U2424 (N_2424,N_1723,N_1524);
or U2425 (N_2425,N_1681,N_1054);
nand U2426 (N_2426,N_1158,N_1340);
nand U2427 (N_2427,N_1595,N_1507);
nor U2428 (N_2428,N_1038,N_1037);
xnor U2429 (N_2429,N_1623,N_1001);
nor U2430 (N_2430,N_1853,N_1046);
nor U2431 (N_2431,N_1481,N_1180);
nor U2432 (N_2432,N_1118,N_1727);
nand U2433 (N_2433,N_1850,N_1430);
and U2434 (N_2434,N_1878,N_1490);
and U2435 (N_2435,N_1278,N_1440);
and U2436 (N_2436,N_1384,N_1103);
and U2437 (N_2437,N_1622,N_1375);
nor U2438 (N_2438,N_1972,N_1116);
or U2439 (N_2439,N_1410,N_1713);
or U2440 (N_2440,N_1331,N_1906);
nor U2441 (N_2441,N_1367,N_1753);
nand U2442 (N_2442,N_1907,N_1130);
nor U2443 (N_2443,N_1156,N_1190);
nor U2444 (N_2444,N_1975,N_1399);
nor U2445 (N_2445,N_1518,N_1602);
or U2446 (N_2446,N_1760,N_1920);
and U2447 (N_2447,N_1605,N_1995);
and U2448 (N_2448,N_1011,N_1599);
nor U2449 (N_2449,N_1637,N_1866);
and U2450 (N_2450,N_1883,N_1686);
nor U2451 (N_2451,N_1976,N_1691);
and U2452 (N_2452,N_1148,N_1227);
and U2453 (N_2453,N_1338,N_1361);
nor U2454 (N_2454,N_1091,N_1343);
and U2455 (N_2455,N_1355,N_1192);
xor U2456 (N_2456,N_1019,N_1291);
and U2457 (N_2457,N_1285,N_1801);
nand U2458 (N_2458,N_1699,N_1596);
or U2459 (N_2459,N_1413,N_1401);
or U2460 (N_2460,N_1988,N_1714);
and U2461 (N_2461,N_1784,N_1264);
nor U2462 (N_2462,N_1335,N_1127);
nand U2463 (N_2463,N_1145,N_1893);
nand U2464 (N_2464,N_1506,N_1811);
and U2465 (N_2465,N_1455,N_1102);
and U2466 (N_2466,N_1016,N_1247);
and U2467 (N_2467,N_1171,N_1025);
and U2468 (N_2468,N_1829,N_1182);
nor U2469 (N_2469,N_1653,N_1337);
nor U2470 (N_2470,N_1023,N_1380);
nand U2471 (N_2471,N_1687,N_1529);
nor U2472 (N_2472,N_1772,N_1741);
nor U2473 (N_2473,N_1624,N_1917);
nand U2474 (N_2474,N_1245,N_1645);
or U2475 (N_2475,N_1643,N_1242);
or U2476 (N_2476,N_1500,N_1108);
and U2477 (N_2477,N_1042,N_1378);
nand U2478 (N_2478,N_1564,N_1494);
nor U2479 (N_2479,N_1571,N_1673);
nand U2480 (N_2480,N_1805,N_1902);
or U2481 (N_2481,N_1234,N_1734);
nor U2482 (N_2482,N_1209,N_1586);
or U2483 (N_2483,N_1897,N_1051);
nor U2484 (N_2484,N_1808,N_1690);
nor U2485 (N_2485,N_1057,N_1994);
and U2486 (N_2486,N_1794,N_1100);
nand U2487 (N_2487,N_1206,N_1795);
or U2488 (N_2488,N_1106,N_1248);
nor U2489 (N_2489,N_1114,N_1514);
nand U2490 (N_2490,N_1654,N_1105);
or U2491 (N_2491,N_1457,N_1856);
or U2492 (N_2492,N_1911,N_1311);
and U2493 (N_2493,N_1450,N_1301);
nand U2494 (N_2494,N_1365,N_1858);
xor U2495 (N_2495,N_1796,N_1962);
nand U2496 (N_2496,N_1755,N_1081);
or U2497 (N_2497,N_1351,N_1222);
or U2498 (N_2498,N_1136,N_1664);
and U2499 (N_2499,N_1704,N_1998);
nand U2500 (N_2500,N_1405,N_1431);
and U2501 (N_2501,N_1357,N_1823);
and U2502 (N_2502,N_1719,N_1483);
nor U2503 (N_2503,N_1052,N_1605);
nand U2504 (N_2504,N_1718,N_1783);
or U2505 (N_2505,N_1121,N_1389);
nand U2506 (N_2506,N_1051,N_1652);
nor U2507 (N_2507,N_1708,N_1783);
nand U2508 (N_2508,N_1938,N_1829);
nor U2509 (N_2509,N_1599,N_1062);
or U2510 (N_2510,N_1900,N_1801);
or U2511 (N_2511,N_1213,N_1045);
xor U2512 (N_2512,N_1231,N_1334);
or U2513 (N_2513,N_1799,N_1200);
nor U2514 (N_2514,N_1956,N_1048);
nor U2515 (N_2515,N_1175,N_1428);
and U2516 (N_2516,N_1408,N_1504);
xor U2517 (N_2517,N_1632,N_1268);
and U2518 (N_2518,N_1956,N_1744);
nand U2519 (N_2519,N_1339,N_1040);
or U2520 (N_2520,N_1609,N_1433);
or U2521 (N_2521,N_1826,N_1604);
nor U2522 (N_2522,N_1416,N_1214);
and U2523 (N_2523,N_1718,N_1994);
nand U2524 (N_2524,N_1026,N_1799);
nor U2525 (N_2525,N_1097,N_1639);
and U2526 (N_2526,N_1360,N_1296);
nand U2527 (N_2527,N_1365,N_1131);
and U2528 (N_2528,N_1802,N_1370);
nor U2529 (N_2529,N_1533,N_1543);
nor U2530 (N_2530,N_1630,N_1034);
nor U2531 (N_2531,N_1555,N_1672);
nor U2532 (N_2532,N_1352,N_1920);
xnor U2533 (N_2533,N_1463,N_1456);
nor U2534 (N_2534,N_1627,N_1402);
nor U2535 (N_2535,N_1612,N_1417);
nand U2536 (N_2536,N_1268,N_1458);
or U2537 (N_2537,N_1683,N_1987);
and U2538 (N_2538,N_1818,N_1975);
nand U2539 (N_2539,N_1614,N_1357);
and U2540 (N_2540,N_1353,N_1405);
or U2541 (N_2541,N_1150,N_1241);
xnor U2542 (N_2542,N_1269,N_1596);
nand U2543 (N_2543,N_1627,N_1348);
and U2544 (N_2544,N_1906,N_1076);
and U2545 (N_2545,N_1564,N_1181);
nand U2546 (N_2546,N_1204,N_1145);
nand U2547 (N_2547,N_1141,N_1334);
and U2548 (N_2548,N_1215,N_1341);
nand U2549 (N_2549,N_1732,N_1375);
nand U2550 (N_2550,N_1896,N_1541);
nor U2551 (N_2551,N_1701,N_1295);
nand U2552 (N_2552,N_1057,N_1713);
and U2553 (N_2553,N_1738,N_1092);
nor U2554 (N_2554,N_1837,N_1510);
nand U2555 (N_2555,N_1136,N_1859);
xor U2556 (N_2556,N_1776,N_1083);
nand U2557 (N_2557,N_1513,N_1900);
or U2558 (N_2558,N_1362,N_1309);
nor U2559 (N_2559,N_1721,N_1447);
nand U2560 (N_2560,N_1576,N_1594);
nor U2561 (N_2561,N_1444,N_1265);
and U2562 (N_2562,N_1547,N_1975);
or U2563 (N_2563,N_1408,N_1168);
nand U2564 (N_2564,N_1985,N_1403);
and U2565 (N_2565,N_1414,N_1203);
or U2566 (N_2566,N_1999,N_1577);
nand U2567 (N_2567,N_1432,N_1328);
and U2568 (N_2568,N_1627,N_1634);
nand U2569 (N_2569,N_1804,N_1249);
and U2570 (N_2570,N_1064,N_1039);
and U2571 (N_2571,N_1158,N_1153);
and U2572 (N_2572,N_1962,N_1344);
nor U2573 (N_2573,N_1915,N_1681);
nand U2574 (N_2574,N_1170,N_1742);
nor U2575 (N_2575,N_1481,N_1939);
and U2576 (N_2576,N_1212,N_1465);
or U2577 (N_2577,N_1828,N_1647);
or U2578 (N_2578,N_1037,N_1559);
and U2579 (N_2579,N_1118,N_1580);
nand U2580 (N_2580,N_1287,N_1544);
nand U2581 (N_2581,N_1791,N_1899);
and U2582 (N_2582,N_1241,N_1484);
and U2583 (N_2583,N_1520,N_1408);
or U2584 (N_2584,N_1494,N_1895);
or U2585 (N_2585,N_1678,N_1299);
nor U2586 (N_2586,N_1135,N_1958);
and U2587 (N_2587,N_1878,N_1863);
nand U2588 (N_2588,N_1360,N_1990);
nand U2589 (N_2589,N_1526,N_1955);
xor U2590 (N_2590,N_1050,N_1824);
nor U2591 (N_2591,N_1286,N_1974);
or U2592 (N_2592,N_1005,N_1359);
nor U2593 (N_2593,N_1892,N_1889);
and U2594 (N_2594,N_1205,N_1584);
or U2595 (N_2595,N_1235,N_1106);
nor U2596 (N_2596,N_1427,N_1270);
or U2597 (N_2597,N_1110,N_1304);
nor U2598 (N_2598,N_1786,N_1111);
nor U2599 (N_2599,N_1361,N_1207);
and U2600 (N_2600,N_1790,N_1595);
nand U2601 (N_2601,N_1848,N_1892);
nor U2602 (N_2602,N_1528,N_1113);
or U2603 (N_2603,N_1994,N_1367);
nor U2604 (N_2604,N_1784,N_1367);
nand U2605 (N_2605,N_1393,N_1760);
xnor U2606 (N_2606,N_1369,N_1214);
nand U2607 (N_2607,N_1271,N_1153);
nor U2608 (N_2608,N_1201,N_1989);
nand U2609 (N_2609,N_1674,N_1124);
nand U2610 (N_2610,N_1577,N_1147);
nand U2611 (N_2611,N_1973,N_1466);
nor U2612 (N_2612,N_1497,N_1902);
nor U2613 (N_2613,N_1716,N_1815);
nor U2614 (N_2614,N_1247,N_1678);
and U2615 (N_2615,N_1429,N_1608);
nor U2616 (N_2616,N_1827,N_1055);
nor U2617 (N_2617,N_1349,N_1739);
or U2618 (N_2618,N_1208,N_1581);
or U2619 (N_2619,N_1514,N_1253);
nor U2620 (N_2620,N_1295,N_1906);
nand U2621 (N_2621,N_1332,N_1453);
and U2622 (N_2622,N_1677,N_1449);
and U2623 (N_2623,N_1824,N_1650);
and U2624 (N_2624,N_1894,N_1902);
and U2625 (N_2625,N_1999,N_1842);
nor U2626 (N_2626,N_1418,N_1588);
or U2627 (N_2627,N_1284,N_1140);
and U2628 (N_2628,N_1207,N_1861);
or U2629 (N_2629,N_1538,N_1127);
nand U2630 (N_2630,N_1833,N_1711);
or U2631 (N_2631,N_1241,N_1413);
xnor U2632 (N_2632,N_1832,N_1210);
and U2633 (N_2633,N_1332,N_1800);
nand U2634 (N_2634,N_1484,N_1915);
nand U2635 (N_2635,N_1095,N_1781);
and U2636 (N_2636,N_1801,N_1845);
nand U2637 (N_2637,N_1964,N_1697);
or U2638 (N_2638,N_1461,N_1593);
or U2639 (N_2639,N_1454,N_1267);
nand U2640 (N_2640,N_1350,N_1829);
nand U2641 (N_2641,N_1616,N_1804);
or U2642 (N_2642,N_1839,N_1667);
and U2643 (N_2643,N_1442,N_1131);
or U2644 (N_2644,N_1008,N_1538);
nand U2645 (N_2645,N_1648,N_1316);
nand U2646 (N_2646,N_1822,N_1350);
nor U2647 (N_2647,N_1629,N_1575);
and U2648 (N_2648,N_1388,N_1744);
nor U2649 (N_2649,N_1011,N_1334);
or U2650 (N_2650,N_1513,N_1713);
nand U2651 (N_2651,N_1388,N_1488);
xor U2652 (N_2652,N_1175,N_1157);
or U2653 (N_2653,N_1226,N_1467);
nor U2654 (N_2654,N_1588,N_1402);
nand U2655 (N_2655,N_1481,N_1462);
or U2656 (N_2656,N_1224,N_1707);
or U2657 (N_2657,N_1795,N_1359);
nor U2658 (N_2658,N_1565,N_1116);
nand U2659 (N_2659,N_1103,N_1956);
nand U2660 (N_2660,N_1285,N_1126);
nand U2661 (N_2661,N_1732,N_1323);
nand U2662 (N_2662,N_1325,N_1706);
nand U2663 (N_2663,N_1103,N_1415);
nand U2664 (N_2664,N_1552,N_1965);
and U2665 (N_2665,N_1411,N_1056);
or U2666 (N_2666,N_1881,N_1414);
and U2667 (N_2667,N_1615,N_1209);
nor U2668 (N_2668,N_1714,N_1920);
nand U2669 (N_2669,N_1904,N_1399);
and U2670 (N_2670,N_1976,N_1042);
nor U2671 (N_2671,N_1846,N_1598);
xor U2672 (N_2672,N_1371,N_1767);
nand U2673 (N_2673,N_1514,N_1356);
or U2674 (N_2674,N_1481,N_1669);
nor U2675 (N_2675,N_1925,N_1405);
nor U2676 (N_2676,N_1281,N_1280);
xor U2677 (N_2677,N_1290,N_1339);
or U2678 (N_2678,N_1981,N_1717);
and U2679 (N_2679,N_1899,N_1660);
xnor U2680 (N_2680,N_1053,N_1509);
and U2681 (N_2681,N_1036,N_1710);
nand U2682 (N_2682,N_1282,N_1524);
nor U2683 (N_2683,N_1013,N_1274);
nor U2684 (N_2684,N_1439,N_1436);
or U2685 (N_2685,N_1657,N_1303);
and U2686 (N_2686,N_1922,N_1810);
nand U2687 (N_2687,N_1134,N_1575);
xnor U2688 (N_2688,N_1867,N_1724);
nand U2689 (N_2689,N_1441,N_1862);
nand U2690 (N_2690,N_1329,N_1521);
or U2691 (N_2691,N_1789,N_1132);
nand U2692 (N_2692,N_1636,N_1821);
nor U2693 (N_2693,N_1221,N_1845);
and U2694 (N_2694,N_1357,N_1193);
or U2695 (N_2695,N_1747,N_1329);
or U2696 (N_2696,N_1695,N_1534);
and U2697 (N_2697,N_1863,N_1418);
or U2698 (N_2698,N_1145,N_1461);
and U2699 (N_2699,N_1380,N_1584);
nand U2700 (N_2700,N_1313,N_1451);
nor U2701 (N_2701,N_1627,N_1502);
nor U2702 (N_2702,N_1747,N_1120);
and U2703 (N_2703,N_1153,N_1736);
or U2704 (N_2704,N_1107,N_1474);
and U2705 (N_2705,N_1534,N_1666);
and U2706 (N_2706,N_1622,N_1925);
nand U2707 (N_2707,N_1753,N_1597);
or U2708 (N_2708,N_1349,N_1446);
and U2709 (N_2709,N_1468,N_1177);
nand U2710 (N_2710,N_1500,N_1283);
nor U2711 (N_2711,N_1691,N_1818);
and U2712 (N_2712,N_1718,N_1124);
nand U2713 (N_2713,N_1072,N_1301);
and U2714 (N_2714,N_1080,N_1176);
and U2715 (N_2715,N_1554,N_1070);
and U2716 (N_2716,N_1426,N_1041);
nand U2717 (N_2717,N_1193,N_1133);
and U2718 (N_2718,N_1905,N_1679);
and U2719 (N_2719,N_1373,N_1567);
or U2720 (N_2720,N_1217,N_1605);
or U2721 (N_2721,N_1593,N_1606);
nor U2722 (N_2722,N_1196,N_1482);
xor U2723 (N_2723,N_1615,N_1842);
or U2724 (N_2724,N_1694,N_1493);
nand U2725 (N_2725,N_1975,N_1746);
and U2726 (N_2726,N_1939,N_1334);
nand U2727 (N_2727,N_1819,N_1184);
and U2728 (N_2728,N_1328,N_1978);
or U2729 (N_2729,N_1821,N_1556);
nor U2730 (N_2730,N_1254,N_1028);
and U2731 (N_2731,N_1827,N_1348);
nand U2732 (N_2732,N_1481,N_1553);
and U2733 (N_2733,N_1538,N_1850);
and U2734 (N_2734,N_1595,N_1913);
nand U2735 (N_2735,N_1698,N_1986);
or U2736 (N_2736,N_1667,N_1694);
nor U2737 (N_2737,N_1053,N_1985);
or U2738 (N_2738,N_1629,N_1588);
and U2739 (N_2739,N_1602,N_1358);
nand U2740 (N_2740,N_1493,N_1150);
nand U2741 (N_2741,N_1331,N_1948);
and U2742 (N_2742,N_1719,N_1717);
or U2743 (N_2743,N_1772,N_1747);
nand U2744 (N_2744,N_1982,N_1925);
nand U2745 (N_2745,N_1996,N_1555);
and U2746 (N_2746,N_1154,N_1570);
and U2747 (N_2747,N_1599,N_1660);
nor U2748 (N_2748,N_1276,N_1262);
nand U2749 (N_2749,N_1532,N_1964);
and U2750 (N_2750,N_1982,N_1851);
or U2751 (N_2751,N_1471,N_1224);
and U2752 (N_2752,N_1198,N_1160);
and U2753 (N_2753,N_1519,N_1005);
and U2754 (N_2754,N_1505,N_1659);
or U2755 (N_2755,N_1358,N_1960);
or U2756 (N_2756,N_1653,N_1192);
nand U2757 (N_2757,N_1753,N_1154);
nand U2758 (N_2758,N_1775,N_1076);
and U2759 (N_2759,N_1358,N_1522);
and U2760 (N_2760,N_1696,N_1712);
or U2761 (N_2761,N_1066,N_1097);
nor U2762 (N_2762,N_1072,N_1350);
nor U2763 (N_2763,N_1822,N_1249);
nand U2764 (N_2764,N_1798,N_1349);
and U2765 (N_2765,N_1851,N_1394);
nand U2766 (N_2766,N_1157,N_1028);
nand U2767 (N_2767,N_1589,N_1457);
nor U2768 (N_2768,N_1204,N_1962);
nor U2769 (N_2769,N_1345,N_1650);
nor U2770 (N_2770,N_1804,N_1948);
nand U2771 (N_2771,N_1059,N_1357);
nand U2772 (N_2772,N_1608,N_1098);
nand U2773 (N_2773,N_1757,N_1662);
nand U2774 (N_2774,N_1336,N_1356);
or U2775 (N_2775,N_1732,N_1438);
or U2776 (N_2776,N_1528,N_1521);
or U2777 (N_2777,N_1074,N_1551);
and U2778 (N_2778,N_1905,N_1714);
and U2779 (N_2779,N_1205,N_1138);
nor U2780 (N_2780,N_1896,N_1904);
and U2781 (N_2781,N_1189,N_1383);
and U2782 (N_2782,N_1829,N_1488);
and U2783 (N_2783,N_1576,N_1746);
or U2784 (N_2784,N_1198,N_1517);
and U2785 (N_2785,N_1153,N_1224);
nand U2786 (N_2786,N_1782,N_1050);
nand U2787 (N_2787,N_1494,N_1864);
and U2788 (N_2788,N_1075,N_1097);
nor U2789 (N_2789,N_1372,N_1749);
nor U2790 (N_2790,N_1991,N_1454);
or U2791 (N_2791,N_1594,N_1235);
and U2792 (N_2792,N_1188,N_1737);
nor U2793 (N_2793,N_1827,N_1466);
and U2794 (N_2794,N_1777,N_1556);
and U2795 (N_2795,N_1597,N_1438);
and U2796 (N_2796,N_1262,N_1705);
or U2797 (N_2797,N_1312,N_1099);
and U2798 (N_2798,N_1018,N_1384);
nand U2799 (N_2799,N_1706,N_1957);
nor U2800 (N_2800,N_1945,N_1236);
nand U2801 (N_2801,N_1086,N_1614);
and U2802 (N_2802,N_1268,N_1337);
nor U2803 (N_2803,N_1394,N_1503);
nor U2804 (N_2804,N_1087,N_1617);
or U2805 (N_2805,N_1187,N_1508);
nand U2806 (N_2806,N_1048,N_1970);
or U2807 (N_2807,N_1617,N_1986);
xor U2808 (N_2808,N_1867,N_1236);
nor U2809 (N_2809,N_1724,N_1410);
or U2810 (N_2810,N_1023,N_1584);
or U2811 (N_2811,N_1931,N_1161);
and U2812 (N_2812,N_1131,N_1952);
and U2813 (N_2813,N_1184,N_1341);
nor U2814 (N_2814,N_1374,N_1713);
nor U2815 (N_2815,N_1575,N_1310);
nor U2816 (N_2816,N_1908,N_1533);
nor U2817 (N_2817,N_1409,N_1371);
or U2818 (N_2818,N_1463,N_1827);
nand U2819 (N_2819,N_1788,N_1573);
and U2820 (N_2820,N_1783,N_1434);
nor U2821 (N_2821,N_1649,N_1734);
nand U2822 (N_2822,N_1304,N_1208);
nor U2823 (N_2823,N_1781,N_1387);
and U2824 (N_2824,N_1405,N_1340);
and U2825 (N_2825,N_1501,N_1114);
nand U2826 (N_2826,N_1195,N_1199);
nand U2827 (N_2827,N_1888,N_1120);
or U2828 (N_2828,N_1057,N_1193);
nand U2829 (N_2829,N_1733,N_1767);
nand U2830 (N_2830,N_1100,N_1961);
or U2831 (N_2831,N_1495,N_1625);
nor U2832 (N_2832,N_1639,N_1523);
nand U2833 (N_2833,N_1951,N_1375);
nor U2834 (N_2834,N_1406,N_1270);
or U2835 (N_2835,N_1680,N_1263);
and U2836 (N_2836,N_1786,N_1213);
and U2837 (N_2837,N_1891,N_1120);
and U2838 (N_2838,N_1862,N_1758);
or U2839 (N_2839,N_1329,N_1242);
nand U2840 (N_2840,N_1165,N_1274);
or U2841 (N_2841,N_1101,N_1126);
or U2842 (N_2842,N_1384,N_1495);
nand U2843 (N_2843,N_1962,N_1494);
nand U2844 (N_2844,N_1720,N_1906);
nor U2845 (N_2845,N_1111,N_1797);
or U2846 (N_2846,N_1376,N_1261);
or U2847 (N_2847,N_1617,N_1407);
and U2848 (N_2848,N_1714,N_1144);
nor U2849 (N_2849,N_1581,N_1914);
nand U2850 (N_2850,N_1807,N_1227);
nand U2851 (N_2851,N_1346,N_1255);
nor U2852 (N_2852,N_1148,N_1952);
or U2853 (N_2853,N_1478,N_1043);
nor U2854 (N_2854,N_1246,N_1394);
nor U2855 (N_2855,N_1413,N_1453);
xor U2856 (N_2856,N_1266,N_1813);
xor U2857 (N_2857,N_1683,N_1834);
or U2858 (N_2858,N_1344,N_1146);
nor U2859 (N_2859,N_1778,N_1079);
and U2860 (N_2860,N_1012,N_1270);
or U2861 (N_2861,N_1420,N_1295);
or U2862 (N_2862,N_1290,N_1765);
nor U2863 (N_2863,N_1053,N_1934);
or U2864 (N_2864,N_1539,N_1139);
and U2865 (N_2865,N_1357,N_1445);
and U2866 (N_2866,N_1554,N_1128);
and U2867 (N_2867,N_1379,N_1332);
and U2868 (N_2868,N_1676,N_1249);
and U2869 (N_2869,N_1148,N_1030);
nand U2870 (N_2870,N_1339,N_1835);
or U2871 (N_2871,N_1430,N_1272);
nand U2872 (N_2872,N_1979,N_1710);
nor U2873 (N_2873,N_1913,N_1812);
or U2874 (N_2874,N_1297,N_1835);
and U2875 (N_2875,N_1764,N_1640);
or U2876 (N_2876,N_1631,N_1329);
nor U2877 (N_2877,N_1544,N_1586);
and U2878 (N_2878,N_1807,N_1781);
nand U2879 (N_2879,N_1887,N_1955);
or U2880 (N_2880,N_1746,N_1289);
and U2881 (N_2881,N_1522,N_1162);
or U2882 (N_2882,N_1482,N_1327);
nor U2883 (N_2883,N_1741,N_1907);
or U2884 (N_2884,N_1832,N_1181);
nor U2885 (N_2885,N_1845,N_1278);
nand U2886 (N_2886,N_1555,N_1738);
and U2887 (N_2887,N_1390,N_1616);
nand U2888 (N_2888,N_1821,N_1597);
nor U2889 (N_2889,N_1763,N_1058);
nor U2890 (N_2890,N_1015,N_1253);
nand U2891 (N_2891,N_1573,N_1544);
and U2892 (N_2892,N_1980,N_1412);
nor U2893 (N_2893,N_1675,N_1632);
nand U2894 (N_2894,N_1248,N_1013);
nor U2895 (N_2895,N_1352,N_1967);
and U2896 (N_2896,N_1479,N_1995);
or U2897 (N_2897,N_1614,N_1367);
nor U2898 (N_2898,N_1180,N_1768);
nor U2899 (N_2899,N_1683,N_1313);
and U2900 (N_2900,N_1183,N_1684);
or U2901 (N_2901,N_1752,N_1825);
and U2902 (N_2902,N_1534,N_1382);
nor U2903 (N_2903,N_1551,N_1140);
or U2904 (N_2904,N_1917,N_1940);
and U2905 (N_2905,N_1464,N_1211);
nand U2906 (N_2906,N_1954,N_1254);
and U2907 (N_2907,N_1273,N_1246);
and U2908 (N_2908,N_1013,N_1149);
nor U2909 (N_2909,N_1168,N_1721);
nand U2910 (N_2910,N_1266,N_1217);
or U2911 (N_2911,N_1453,N_1550);
nor U2912 (N_2912,N_1308,N_1117);
or U2913 (N_2913,N_1973,N_1998);
and U2914 (N_2914,N_1824,N_1661);
and U2915 (N_2915,N_1146,N_1255);
and U2916 (N_2916,N_1098,N_1764);
xor U2917 (N_2917,N_1608,N_1871);
nand U2918 (N_2918,N_1448,N_1327);
nor U2919 (N_2919,N_1890,N_1132);
and U2920 (N_2920,N_1987,N_1868);
xnor U2921 (N_2921,N_1183,N_1846);
or U2922 (N_2922,N_1649,N_1169);
or U2923 (N_2923,N_1794,N_1635);
and U2924 (N_2924,N_1303,N_1680);
nand U2925 (N_2925,N_1030,N_1577);
and U2926 (N_2926,N_1454,N_1038);
or U2927 (N_2927,N_1648,N_1657);
nand U2928 (N_2928,N_1333,N_1668);
and U2929 (N_2929,N_1888,N_1931);
and U2930 (N_2930,N_1502,N_1944);
or U2931 (N_2931,N_1979,N_1251);
nand U2932 (N_2932,N_1566,N_1142);
nand U2933 (N_2933,N_1845,N_1670);
nor U2934 (N_2934,N_1702,N_1396);
nor U2935 (N_2935,N_1051,N_1991);
or U2936 (N_2936,N_1012,N_1421);
nand U2937 (N_2937,N_1350,N_1809);
and U2938 (N_2938,N_1792,N_1488);
nand U2939 (N_2939,N_1984,N_1431);
nor U2940 (N_2940,N_1163,N_1507);
nor U2941 (N_2941,N_1451,N_1011);
xnor U2942 (N_2942,N_1538,N_1765);
or U2943 (N_2943,N_1543,N_1181);
nor U2944 (N_2944,N_1868,N_1718);
nor U2945 (N_2945,N_1103,N_1816);
or U2946 (N_2946,N_1857,N_1503);
nor U2947 (N_2947,N_1105,N_1531);
or U2948 (N_2948,N_1122,N_1666);
and U2949 (N_2949,N_1874,N_1593);
nor U2950 (N_2950,N_1792,N_1336);
nand U2951 (N_2951,N_1606,N_1098);
nand U2952 (N_2952,N_1727,N_1973);
nand U2953 (N_2953,N_1045,N_1986);
or U2954 (N_2954,N_1742,N_1373);
nor U2955 (N_2955,N_1516,N_1583);
and U2956 (N_2956,N_1732,N_1925);
or U2957 (N_2957,N_1608,N_1126);
nand U2958 (N_2958,N_1714,N_1743);
and U2959 (N_2959,N_1702,N_1018);
and U2960 (N_2960,N_1467,N_1550);
or U2961 (N_2961,N_1149,N_1728);
nand U2962 (N_2962,N_1753,N_1773);
nor U2963 (N_2963,N_1669,N_1594);
and U2964 (N_2964,N_1806,N_1593);
and U2965 (N_2965,N_1264,N_1080);
and U2966 (N_2966,N_1124,N_1701);
or U2967 (N_2967,N_1790,N_1844);
nand U2968 (N_2968,N_1125,N_1361);
nor U2969 (N_2969,N_1942,N_1726);
nand U2970 (N_2970,N_1809,N_1371);
or U2971 (N_2971,N_1641,N_1477);
and U2972 (N_2972,N_1677,N_1236);
nor U2973 (N_2973,N_1867,N_1347);
nand U2974 (N_2974,N_1409,N_1901);
or U2975 (N_2975,N_1196,N_1253);
or U2976 (N_2976,N_1059,N_1510);
nor U2977 (N_2977,N_1986,N_1571);
nand U2978 (N_2978,N_1795,N_1717);
nor U2979 (N_2979,N_1508,N_1072);
nor U2980 (N_2980,N_1366,N_1005);
or U2981 (N_2981,N_1246,N_1656);
nor U2982 (N_2982,N_1489,N_1115);
nand U2983 (N_2983,N_1667,N_1755);
nor U2984 (N_2984,N_1430,N_1233);
and U2985 (N_2985,N_1505,N_1166);
or U2986 (N_2986,N_1965,N_1767);
nor U2987 (N_2987,N_1595,N_1030);
and U2988 (N_2988,N_1471,N_1929);
and U2989 (N_2989,N_1093,N_1838);
nor U2990 (N_2990,N_1639,N_1486);
or U2991 (N_2991,N_1088,N_1596);
or U2992 (N_2992,N_1196,N_1592);
nor U2993 (N_2993,N_1416,N_1220);
or U2994 (N_2994,N_1772,N_1307);
and U2995 (N_2995,N_1630,N_1456);
nand U2996 (N_2996,N_1023,N_1591);
or U2997 (N_2997,N_1082,N_1383);
and U2998 (N_2998,N_1420,N_1218);
or U2999 (N_2999,N_1242,N_1123);
nor U3000 (N_3000,N_2919,N_2343);
nor U3001 (N_3001,N_2554,N_2645);
and U3002 (N_3002,N_2702,N_2301);
nand U3003 (N_3003,N_2143,N_2329);
or U3004 (N_3004,N_2663,N_2442);
or U3005 (N_3005,N_2743,N_2277);
or U3006 (N_3006,N_2328,N_2956);
or U3007 (N_3007,N_2394,N_2647);
xor U3008 (N_3008,N_2062,N_2559);
and U3009 (N_3009,N_2855,N_2545);
nor U3010 (N_3010,N_2347,N_2157);
nor U3011 (N_3011,N_2473,N_2522);
nand U3012 (N_3012,N_2930,N_2144);
or U3013 (N_3013,N_2226,N_2345);
and U3014 (N_3014,N_2011,N_2198);
or U3015 (N_3015,N_2918,N_2570);
or U3016 (N_3016,N_2177,N_2646);
nor U3017 (N_3017,N_2699,N_2741);
and U3018 (N_3018,N_2366,N_2727);
nand U3019 (N_3019,N_2139,N_2450);
nor U3020 (N_3020,N_2117,N_2175);
nand U3021 (N_3021,N_2709,N_2395);
and U3022 (N_3022,N_2502,N_2245);
and U3023 (N_3023,N_2374,N_2035);
or U3024 (N_3024,N_2736,N_2611);
and U3025 (N_3025,N_2221,N_2170);
and U3026 (N_3026,N_2004,N_2029);
or U3027 (N_3027,N_2661,N_2444);
and U3028 (N_3028,N_2520,N_2514);
and U3029 (N_3029,N_2840,N_2882);
and U3030 (N_3030,N_2729,N_2862);
nand U3031 (N_3031,N_2106,N_2335);
nor U3032 (N_3032,N_2490,N_2353);
or U3033 (N_3033,N_2375,N_2952);
or U3034 (N_3034,N_2735,N_2419);
or U3035 (N_3035,N_2251,N_2385);
nand U3036 (N_3036,N_2298,N_2643);
nand U3037 (N_3037,N_2656,N_2551);
and U3038 (N_3038,N_2701,N_2449);
or U3039 (N_3039,N_2093,N_2481);
nand U3040 (N_3040,N_2732,N_2489);
and U3041 (N_3041,N_2432,N_2584);
and U3042 (N_3042,N_2210,N_2516);
or U3043 (N_3043,N_2608,N_2090);
nand U3044 (N_3044,N_2580,N_2047);
or U3045 (N_3045,N_2512,N_2379);
nor U3046 (N_3046,N_2823,N_2621);
and U3047 (N_3047,N_2873,N_2409);
nor U3048 (N_3048,N_2503,N_2601);
nand U3049 (N_3049,N_2839,N_2708);
nor U3050 (N_3050,N_2892,N_2475);
nor U3051 (N_3051,N_2519,N_2109);
and U3052 (N_3052,N_2931,N_2224);
and U3053 (N_3053,N_2542,N_2212);
or U3054 (N_3054,N_2453,N_2941);
and U3055 (N_3055,N_2742,N_2429);
nor U3056 (N_3056,N_2174,N_2695);
or U3057 (N_3057,N_2365,N_2228);
or U3058 (N_3058,N_2668,N_2414);
nand U3059 (N_3059,N_2402,N_2209);
and U3060 (N_3060,N_2197,N_2739);
and U3061 (N_3061,N_2960,N_2575);
nor U3062 (N_3062,N_2521,N_2119);
nor U3063 (N_3063,N_2002,N_2319);
and U3064 (N_3064,N_2880,N_2543);
nor U3065 (N_3065,N_2199,N_2779);
and U3066 (N_3066,N_2459,N_2641);
nor U3067 (N_3067,N_2162,N_2843);
and U3068 (N_3068,N_2994,N_2132);
and U3069 (N_3069,N_2965,N_2988);
or U3070 (N_3070,N_2883,N_2805);
or U3071 (N_3071,N_2412,N_2057);
nor U3072 (N_3072,N_2692,N_2636);
and U3073 (N_3073,N_2902,N_2286);
nand U3074 (N_3074,N_2788,N_2091);
nor U3075 (N_3075,N_2875,N_2336);
nor U3076 (N_3076,N_2416,N_2628);
nor U3077 (N_3077,N_2768,N_2907);
xor U3078 (N_3078,N_2420,N_2947);
nor U3079 (N_3079,N_2461,N_2786);
nand U3080 (N_3080,N_2678,N_2178);
and U3081 (N_3081,N_2484,N_2480);
or U3082 (N_3082,N_2242,N_2711);
nor U3083 (N_3083,N_2059,N_2186);
nor U3084 (N_3084,N_2651,N_2760);
nand U3085 (N_3085,N_2857,N_2725);
or U3086 (N_3086,N_2547,N_2368);
and U3087 (N_3087,N_2165,N_2748);
nor U3088 (N_3088,N_2120,N_2184);
nor U3089 (N_3089,N_2208,N_2518);
or U3090 (N_3090,N_2408,N_2285);
and U3091 (N_3091,N_2269,N_2346);
and U3092 (N_3092,N_2391,N_2278);
nand U3093 (N_3093,N_2785,N_2439);
nand U3094 (N_3094,N_2899,N_2326);
nand U3095 (N_3095,N_2150,N_2372);
or U3096 (N_3096,N_2548,N_2146);
nor U3097 (N_3097,N_2778,N_2496);
or U3098 (N_3098,N_2094,N_2889);
and U3099 (N_3099,N_2258,N_2822);
nor U3100 (N_3100,N_2361,N_2576);
or U3101 (N_3101,N_2142,N_2888);
nor U3102 (N_3102,N_2625,N_2176);
nand U3103 (N_3103,N_2722,N_2406);
and U3104 (N_3104,N_2044,N_2827);
nand U3105 (N_3105,N_2976,N_2891);
nor U3106 (N_3106,N_2943,N_2253);
or U3107 (N_3107,N_2008,N_2179);
nand U3108 (N_3108,N_2780,N_2043);
or U3109 (N_3109,N_2151,N_2819);
or U3110 (N_3110,N_2923,N_2334);
or U3111 (N_3111,N_2966,N_2793);
nand U3112 (N_3112,N_2130,N_2492);
nand U3113 (N_3113,N_2493,N_2967);
nor U3114 (N_3114,N_2055,N_2306);
nand U3115 (N_3115,N_2034,N_2979);
nand U3116 (N_3116,N_2160,N_2108);
or U3117 (N_3117,N_2844,N_2893);
or U3118 (N_3118,N_2980,N_2627);
nor U3119 (N_3119,N_2852,N_2288);
or U3120 (N_3120,N_2498,N_2389);
nand U3121 (N_3121,N_2540,N_2193);
nor U3122 (N_3122,N_2992,N_2972);
xor U3123 (N_3123,N_2549,N_2356);
nor U3124 (N_3124,N_2808,N_2148);
nor U3125 (N_3125,N_2039,N_2073);
and U3126 (N_3126,N_2957,N_2386);
or U3127 (N_3127,N_2504,N_2655);
nand U3128 (N_3128,N_2716,N_2024);
nor U3129 (N_3129,N_2604,N_2973);
nand U3130 (N_3130,N_2217,N_2917);
nand U3131 (N_3131,N_2050,N_2858);
and U3132 (N_3132,N_2854,N_2940);
or U3133 (N_3133,N_2403,N_2810);
or U3134 (N_3134,N_2938,N_2700);
nand U3135 (N_3135,N_2082,N_2796);
nor U3136 (N_3136,N_2758,N_2293);
nor U3137 (N_3137,N_2488,N_2592);
or U3138 (N_3138,N_2950,N_2266);
or U3139 (N_3139,N_2616,N_2623);
or U3140 (N_3140,N_2167,N_2820);
xor U3141 (N_3141,N_2946,N_2595);
nand U3142 (N_3142,N_2618,N_2640);
and U3143 (N_3143,N_2795,N_2136);
nor U3144 (N_3144,N_2593,N_2089);
nor U3145 (N_3145,N_2927,N_2614);
nor U3146 (N_3146,N_2737,N_2624);
nor U3147 (N_3147,N_2693,N_2418);
nor U3148 (N_3148,N_2898,N_2951);
nor U3149 (N_3149,N_2381,N_2715);
and U3150 (N_3150,N_2192,N_2964);
nand U3151 (N_3151,N_2141,N_2207);
or U3152 (N_3152,N_2527,N_2783);
nand U3153 (N_3153,N_2734,N_2316);
nand U3154 (N_3154,N_2685,N_2289);
nand U3155 (N_3155,N_2399,N_2222);
and U3156 (N_3156,N_2667,N_2849);
nor U3157 (N_3157,N_2817,N_2171);
and U3158 (N_3158,N_2046,N_2485);
nand U3159 (N_3159,N_2443,N_2309);
nor U3160 (N_3160,N_2659,N_2775);
nand U3161 (N_3161,N_2102,N_2415);
or U3162 (N_3162,N_2276,N_2860);
or U3163 (N_3163,N_2264,N_2010);
nor U3164 (N_3164,N_2291,N_2045);
nand U3165 (N_3165,N_2052,N_2427);
or U3166 (N_3166,N_2961,N_2187);
or U3167 (N_3167,N_2836,N_2241);
nand U3168 (N_3168,N_2870,N_2128);
nand U3169 (N_3169,N_2523,N_2405);
or U3170 (N_3170,N_2067,N_2376);
and U3171 (N_3171,N_2612,N_2189);
or U3172 (N_3172,N_2206,N_2639);
and U3173 (N_3173,N_2792,N_2666);
or U3174 (N_3174,N_2074,N_2662);
nand U3175 (N_3175,N_2006,N_2016);
or U3176 (N_3176,N_2607,N_2033);
or U3177 (N_3177,N_2782,N_2948);
nor U3178 (N_3178,N_2642,N_2755);
or U3179 (N_3179,N_2040,N_2740);
or U3180 (N_3180,N_2027,N_2384);
or U3181 (N_3181,N_2267,N_2332);
nor U3182 (N_3182,N_2677,N_2292);
or U3183 (N_3183,N_2798,N_2300);
xnor U3184 (N_3184,N_2903,N_2746);
xor U3185 (N_3185,N_2750,N_2993);
nand U3186 (N_3186,N_2697,N_2201);
nand U3187 (N_3187,N_2581,N_2265);
or U3188 (N_3188,N_2850,N_2652);
and U3189 (N_3189,N_2881,N_2477);
nand U3190 (N_3190,N_2660,N_2211);
nor U3191 (N_3191,N_2771,N_2280);
and U3192 (N_3192,N_2598,N_2654);
and U3193 (N_3193,N_2859,N_2632);
nor U3194 (N_3194,N_2003,N_2272);
and U3195 (N_3195,N_2116,N_2606);
nor U3196 (N_3196,N_2088,N_2400);
nor U3197 (N_3197,N_2552,N_2856);
and U3198 (N_3198,N_2437,N_2599);
or U3199 (N_3199,N_2445,N_2229);
or U3200 (N_3200,N_2537,N_2924);
and U3201 (N_3201,N_2683,N_2048);
nand U3202 (N_3202,N_2322,N_2686);
or U3203 (N_3203,N_2303,N_2674);
or U3204 (N_3204,N_2248,N_2842);
and U3205 (N_3205,N_2219,N_2704);
and U3206 (N_3206,N_2182,N_2049);
and U3207 (N_3207,N_2355,N_2991);
nand U3208 (N_3208,N_2825,N_2564);
and U3209 (N_3209,N_2246,N_2271);
and U3210 (N_3210,N_2113,N_2600);
and U3211 (N_3211,N_2491,N_2104);
nor U3212 (N_3212,N_2086,N_2235);
and U3213 (N_3213,N_2738,N_2001);
and U3214 (N_3214,N_2215,N_2020);
and U3215 (N_3215,N_2511,N_2318);
and U3216 (N_3216,N_2287,N_2107);
nor U3217 (N_3217,N_2804,N_2434);
or U3218 (N_3218,N_2273,N_2297);
and U3219 (N_3219,N_2833,N_2007);
nand U3220 (N_3220,N_2370,N_2083);
nor U3221 (N_3221,N_2214,N_2078);
nor U3222 (N_3222,N_2313,N_2868);
nand U3223 (N_3223,N_2626,N_2500);
or U3224 (N_3224,N_2865,N_2900);
and U3225 (N_3225,N_2784,N_2841);
nand U3226 (N_3226,N_2005,N_2482);
nor U3227 (N_3227,N_2634,N_2451);
and U3228 (N_3228,N_2230,N_2396);
nor U3229 (N_3229,N_2351,N_2851);
or U3230 (N_3230,N_2455,N_2095);
or U3231 (N_3231,N_2791,N_2350);
or U3232 (N_3232,N_2181,N_2495);
or U3233 (N_3233,N_2337,N_2173);
nand U3234 (N_3234,N_2259,N_2213);
and U3235 (N_3235,N_2470,N_2390);
nor U3236 (N_3236,N_2041,N_2986);
and U3237 (N_3237,N_2497,N_2731);
nor U3238 (N_3238,N_2526,N_2871);
nor U3239 (N_3239,N_2975,N_2204);
nor U3240 (N_3240,N_2435,N_2325);
nor U3241 (N_3241,N_2247,N_2814);
or U3242 (N_3242,N_2260,N_2354);
and U3243 (N_3243,N_2072,N_2362);
nor U3244 (N_3244,N_2312,N_2762);
nor U3245 (N_3245,N_2373,N_2115);
nand U3246 (N_3246,N_2720,N_2910);
or U3247 (N_3247,N_2932,N_2111);
or U3248 (N_3248,N_2431,N_2818);
nand U3249 (N_3249,N_2582,N_2687);
nor U3250 (N_3250,N_2462,N_2051);
and U3251 (N_3251,N_2525,N_2989);
or U3252 (N_3252,N_2487,N_2797);
or U3253 (N_3253,N_2556,N_2558);
nand U3254 (N_3254,N_2320,N_2773);
and U3255 (N_3255,N_2826,N_2331);
and U3256 (N_3256,N_2590,N_2605);
and U3257 (N_3257,N_2237,N_2220);
or U3258 (N_3258,N_2571,N_2154);
and U3259 (N_3259,N_2799,N_2188);
nand U3260 (N_3260,N_2617,N_2721);
nand U3261 (N_3261,N_2974,N_2939);
or U3262 (N_3262,N_2030,N_2425);
and U3263 (N_3263,N_2152,N_2065);
nand U3264 (N_3264,N_2829,N_2447);
nor U3265 (N_3265,N_2769,N_2284);
or U3266 (N_3266,N_2494,N_2996);
nor U3267 (N_3267,N_2270,N_2806);
nand U3268 (N_3268,N_2311,N_2125);
nand U3269 (N_3269,N_2648,N_2638);
nand U3270 (N_3270,N_2249,N_2848);
xor U3271 (N_3271,N_2096,N_2377);
or U3272 (N_3272,N_2834,N_2568);
nand U3273 (N_3273,N_2421,N_2454);
nand U3274 (N_3274,N_2506,N_2861);
xnor U3275 (N_3275,N_2921,N_2131);
nand U3276 (N_3276,N_2256,N_2250);
or U3277 (N_3277,N_2075,N_2025);
nand U3278 (N_3278,N_2529,N_2159);
and U3279 (N_3279,N_2909,N_2133);
and U3280 (N_3280,N_2507,N_2069);
nor U3281 (N_3281,N_2100,N_2982);
nor U3282 (N_3282,N_2790,N_2995);
and U3283 (N_3283,N_2935,N_2613);
nor U3284 (N_3284,N_2101,N_2754);
nand U3285 (N_3285,N_2751,N_2619);
and U3286 (N_3286,N_2528,N_2572);
nor U3287 (N_3287,N_2710,N_2036);
xnor U3288 (N_3288,N_2591,N_2717);
and U3289 (N_3289,N_2424,N_2916);
nand U3290 (N_3290,N_2673,N_2949);
and U3291 (N_3291,N_2501,N_2018);
nor U3292 (N_3292,N_2103,N_2315);
and U3293 (N_3293,N_2781,N_2080);
nor U3294 (N_3294,N_2837,N_2679);
or U3295 (N_3295,N_2539,N_2895);
and U3296 (N_3296,N_2962,N_2846);
nand U3297 (N_3297,N_2513,N_2596);
nand U3298 (N_3298,N_2535,N_2650);
or U3299 (N_3299,N_2594,N_2168);
nor U3300 (N_3300,N_2944,N_2299);
or U3301 (N_3301,N_2026,N_2963);
and U3302 (N_3302,N_2032,N_2438);
nor U3303 (N_3303,N_2359,N_2068);
nor U3304 (N_3304,N_2812,N_2426);
nor U3305 (N_3305,N_2227,N_2060);
and U3306 (N_3306,N_2759,N_2983);
and U3307 (N_3307,N_2901,N_2533);
nand U3308 (N_3308,N_2615,N_2585);
and U3309 (N_3309,N_2317,N_2969);
and U3310 (N_3310,N_2124,N_2586);
or U3311 (N_3311,N_2195,N_2824);
or U3312 (N_3312,N_2998,N_2555);
nand U3313 (N_3313,N_2885,N_2936);
nor U3314 (N_3314,N_2014,N_2565);
and U3315 (N_3315,N_2787,N_2452);
xor U3316 (N_3316,N_2573,N_2371);
or U3317 (N_3317,N_2509,N_2015);
or U3318 (N_3318,N_2971,N_2534);
or U3319 (N_3319,N_2216,N_2469);
nor U3320 (N_3320,N_2190,N_2231);
and U3321 (N_3321,N_2985,N_2122);
nand U3322 (N_3322,N_2838,N_2794);
nor U3323 (N_3323,N_2821,N_2436);
nand U3324 (N_3324,N_2672,N_2084);
nand U3325 (N_3325,N_2397,N_2314);
nand U3326 (N_3326,N_2205,N_2012);
nor U3327 (N_3327,N_2483,N_2149);
or U3328 (N_3328,N_2684,N_2079);
xnor U3329 (N_3329,N_2349,N_2433);
nor U3330 (N_3330,N_2990,N_2121);
nand U3331 (N_3331,N_2338,N_2257);
nand U3332 (N_3332,N_2290,N_2166);
nand U3333 (N_3333,N_2164,N_2926);
and U3334 (N_3334,N_2281,N_2383);
nor U3335 (N_3335,N_2728,N_2457);
nand U3336 (N_3336,N_2567,N_2587);
nor U3337 (N_3337,N_2904,N_2676);
and U3338 (N_3338,N_2610,N_2087);
nand U3339 (N_3339,N_2054,N_2766);
and U3340 (N_3340,N_2038,N_2378);
nand U3341 (N_3341,N_2458,N_2183);
and U3342 (N_3342,N_2310,N_2874);
and U3343 (N_3343,N_2000,N_2404);
or U3344 (N_3344,N_2369,N_2745);
or U3345 (N_3345,N_2879,N_2479);
nand U3346 (N_3346,N_2037,N_2382);
or U3347 (N_3347,N_2296,N_2588);
nand U3348 (N_3348,N_2254,N_2560);
or U3349 (N_3349,N_2392,N_2225);
and U3350 (N_3350,N_2063,N_2476);
nor U3351 (N_3351,N_2876,N_2689);
nand U3352 (N_3352,N_2756,N_2753);
nand U3353 (N_3353,N_2637,N_2255);
nand U3354 (N_3354,N_2077,N_2589);
and U3355 (N_3355,N_2200,N_2330);
or U3356 (N_3356,N_2423,N_2380);
nor U3357 (N_3357,N_2017,N_2723);
or U3358 (N_3358,N_2076,N_2097);
nand U3359 (N_3359,N_2955,N_2446);
and U3360 (N_3360,N_2933,N_2456);
or U3361 (N_3361,N_2691,N_2070);
or U3362 (N_3362,N_2911,N_2172);
nand U3363 (N_3363,N_2263,N_2920);
and U3364 (N_3364,N_2978,N_2765);
or U3365 (N_3365,N_2156,N_2649);
nand U3366 (N_3366,N_2776,N_2906);
nand U3367 (N_3367,N_2577,N_2872);
nor U3368 (N_3368,N_2180,N_2218);
nor U3369 (N_3369,N_2908,N_2092);
nand U3370 (N_3370,N_2105,N_2009);
and U3371 (N_3371,N_2147,N_2719);
or U3372 (N_3372,N_2407,N_2398);
and U3373 (N_3373,N_2863,N_2835);
or U3374 (N_3374,N_2321,N_2413);
and U3375 (N_3375,N_2367,N_2232);
or U3376 (N_3376,N_2510,N_2997);
and U3377 (N_3377,N_2544,N_2448);
nand U3378 (N_3378,N_2622,N_2644);
nand U3379 (N_3379,N_2896,N_2274);
or U3380 (N_3380,N_2262,N_2357);
or U3381 (N_3381,N_2811,N_2233);
or U3382 (N_3382,N_2411,N_2307);
and U3383 (N_3383,N_2730,N_2884);
xnor U3384 (N_3384,N_2864,N_2890);
and U3385 (N_3385,N_2013,N_2724);
nand U3386 (N_3386,N_2401,N_2134);
or U3387 (N_3387,N_2191,N_2464);
nor U3388 (N_3388,N_2410,N_2937);
nand U3389 (N_3389,N_2468,N_2913);
and U3390 (N_3390,N_2244,N_2688);
and U3391 (N_3391,N_2803,N_2866);
or U3392 (N_3392,N_2333,N_2364);
or U3393 (N_3393,N_2635,N_2118);
and U3394 (N_3394,N_2304,N_2505);
nor U3395 (N_3395,N_2532,N_2718);
nor U3396 (N_3396,N_2474,N_2238);
xnor U3397 (N_3397,N_2603,N_2912);
nor U3398 (N_3398,N_2553,N_2252);
and U3399 (N_3399,N_2878,N_2675);
and U3400 (N_3400,N_2914,N_2602);
nand U3401 (N_3401,N_2441,N_2158);
nand U3402 (N_3402,N_2282,N_2669);
nor U3403 (N_3403,N_2744,N_2275);
nor U3404 (N_3404,N_2153,N_2126);
nor U3405 (N_3405,N_2774,N_2085);
nor U3406 (N_3406,N_2800,N_2777);
nand U3407 (N_3407,N_2664,N_2524);
nand U3408 (N_3408,N_2772,N_2886);
and U3409 (N_3409,N_2752,N_2887);
nand U3410 (N_3410,N_2440,N_2620);
and U3411 (N_3411,N_2223,N_2053);
nand U3412 (N_3412,N_2705,N_2633);
nor U3413 (N_3413,N_2813,N_2422);
nor U3414 (N_3414,N_2802,N_2682);
or U3415 (N_3415,N_2023,N_2071);
nand U3416 (N_3416,N_2987,N_2929);
nor U3417 (N_3417,N_2531,N_2767);
nor U3418 (N_3418,N_2417,N_2294);
xor U3419 (N_3419,N_2653,N_2546);
or U3420 (N_3420,N_2344,N_2467);
and U3421 (N_3421,N_2706,N_2770);
or U3422 (N_3422,N_2393,N_2066);
or U3423 (N_3423,N_2845,N_2127);
and U3424 (N_3424,N_2163,N_2970);
or U3425 (N_3425,N_2726,N_2815);
or U3426 (N_3426,N_2135,N_2342);
nand U3427 (N_3427,N_2169,N_2999);
or U3428 (N_3428,N_2234,N_2463);
and U3429 (N_3429,N_2324,N_2283);
nor U3430 (N_3430,N_2968,N_2832);
nor U3431 (N_3431,N_2789,N_2945);
nor U3432 (N_3432,N_2138,N_2302);
nor U3433 (N_3433,N_2098,N_2236);
and U3434 (N_3434,N_2240,N_2478);
nand U3435 (N_3435,N_2022,N_2530);
nand U3436 (N_3436,N_2566,N_2112);
and U3437 (N_3437,N_2203,N_2562);
and U3438 (N_3438,N_2763,N_2757);
and U3439 (N_3439,N_2471,N_2696);
and U3440 (N_3440,N_2578,N_2323);
nor U3441 (N_3441,N_2694,N_2583);
or U3442 (N_3442,N_2922,N_2243);
and U3443 (N_3443,N_2630,N_2749);
nor U3444 (N_3444,N_2714,N_2561);
and U3445 (N_3445,N_2680,N_2959);
nand U3446 (N_3446,N_2194,N_2671);
nand U3447 (N_3447,N_2761,N_2472);
nand U3448 (N_3448,N_2031,N_2161);
and U3449 (N_3449,N_2764,N_2925);
nand U3450 (N_3450,N_2690,N_2609);
nand U3451 (N_3451,N_2123,N_2137);
and U3452 (N_3452,N_2064,N_2387);
or U3453 (N_3453,N_2028,N_2809);
and U3454 (N_3454,N_2466,N_2140);
and U3455 (N_3455,N_2733,N_2061);
nor U3456 (N_3456,N_2631,N_2550);
or U3457 (N_3457,N_2340,N_2894);
xnor U3458 (N_3458,N_2541,N_2579);
nor U3459 (N_3459,N_2905,N_2114);
nor U3460 (N_3460,N_2295,N_2499);
and U3461 (N_3461,N_2099,N_2430);
nand U3462 (N_3462,N_2597,N_2129);
or U3463 (N_3463,N_2363,N_2268);
xnor U3464 (N_3464,N_2185,N_2019);
nor U3465 (N_3465,N_2847,N_2897);
and U3466 (N_3466,N_2508,N_2830);
xnor U3467 (N_3467,N_2428,N_2110);
nand U3468 (N_3468,N_2352,N_2915);
nor U3469 (N_3469,N_2348,N_2981);
or U3470 (N_3470,N_2308,N_2747);
nand U3471 (N_3471,N_2958,N_2703);
nor U3472 (N_3472,N_2388,N_2536);
nand U3473 (N_3473,N_2977,N_2341);
nand U3474 (N_3474,N_2202,N_2707);
nor U3475 (N_3475,N_2953,N_2867);
nor U3476 (N_3476,N_2681,N_2465);
nor U3477 (N_3477,N_2665,N_2081);
and U3478 (N_3478,N_2574,N_2327);
nor U3479 (N_3479,N_2056,N_2486);
and U3480 (N_3480,N_2305,N_2934);
nand U3481 (N_3481,N_2698,N_2538);
or U3482 (N_3482,N_2629,N_2954);
or U3483 (N_3483,N_2928,N_2515);
or U3484 (N_3484,N_2155,N_2657);
nor U3485 (N_3485,N_2360,N_2239);
or U3486 (N_3486,N_2196,N_2339);
xor U3487 (N_3487,N_2816,N_2807);
and U3488 (N_3488,N_2670,N_2828);
and U3489 (N_3489,N_2563,N_2279);
and U3490 (N_3490,N_2557,N_2801);
and U3491 (N_3491,N_2358,N_2021);
nand U3492 (N_3492,N_2569,N_2712);
or U3493 (N_3493,N_2042,N_2831);
or U3494 (N_3494,N_2942,N_2713);
and U3495 (N_3495,N_2058,N_2877);
or U3496 (N_3496,N_2658,N_2984);
nand U3497 (N_3497,N_2517,N_2853);
or U3498 (N_3498,N_2145,N_2460);
nor U3499 (N_3499,N_2869,N_2261);
or U3500 (N_3500,N_2287,N_2364);
nand U3501 (N_3501,N_2759,N_2082);
and U3502 (N_3502,N_2136,N_2466);
nor U3503 (N_3503,N_2547,N_2255);
nand U3504 (N_3504,N_2934,N_2826);
nor U3505 (N_3505,N_2000,N_2632);
or U3506 (N_3506,N_2322,N_2008);
and U3507 (N_3507,N_2630,N_2867);
or U3508 (N_3508,N_2529,N_2728);
nor U3509 (N_3509,N_2984,N_2657);
or U3510 (N_3510,N_2071,N_2954);
or U3511 (N_3511,N_2357,N_2186);
nand U3512 (N_3512,N_2009,N_2997);
and U3513 (N_3513,N_2499,N_2837);
nand U3514 (N_3514,N_2043,N_2325);
nand U3515 (N_3515,N_2665,N_2080);
nand U3516 (N_3516,N_2400,N_2431);
and U3517 (N_3517,N_2400,N_2822);
and U3518 (N_3518,N_2226,N_2224);
and U3519 (N_3519,N_2203,N_2261);
nand U3520 (N_3520,N_2204,N_2661);
or U3521 (N_3521,N_2627,N_2073);
or U3522 (N_3522,N_2340,N_2508);
or U3523 (N_3523,N_2326,N_2962);
nand U3524 (N_3524,N_2346,N_2624);
nor U3525 (N_3525,N_2792,N_2618);
nand U3526 (N_3526,N_2381,N_2440);
or U3527 (N_3527,N_2006,N_2412);
nand U3528 (N_3528,N_2110,N_2931);
nor U3529 (N_3529,N_2876,N_2605);
or U3530 (N_3530,N_2838,N_2216);
and U3531 (N_3531,N_2641,N_2546);
nor U3532 (N_3532,N_2051,N_2163);
nor U3533 (N_3533,N_2979,N_2652);
nor U3534 (N_3534,N_2598,N_2132);
nand U3535 (N_3535,N_2789,N_2888);
and U3536 (N_3536,N_2603,N_2004);
or U3537 (N_3537,N_2360,N_2293);
nor U3538 (N_3538,N_2378,N_2463);
and U3539 (N_3539,N_2317,N_2613);
xor U3540 (N_3540,N_2313,N_2133);
or U3541 (N_3541,N_2765,N_2604);
nor U3542 (N_3542,N_2115,N_2829);
and U3543 (N_3543,N_2877,N_2204);
nand U3544 (N_3544,N_2795,N_2416);
nand U3545 (N_3545,N_2959,N_2804);
nor U3546 (N_3546,N_2104,N_2679);
nor U3547 (N_3547,N_2461,N_2029);
and U3548 (N_3548,N_2038,N_2423);
nor U3549 (N_3549,N_2196,N_2315);
nand U3550 (N_3550,N_2882,N_2828);
and U3551 (N_3551,N_2508,N_2933);
and U3552 (N_3552,N_2304,N_2466);
or U3553 (N_3553,N_2269,N_2694);
nor U3554 (N_3554,N_2978,N_2356);
or U3555 (N_3555,N_2180,N_2032);
or U3556 (N_3556,N_2382,N_2112);
xnor U3557 (N_3557,N_2684,N_2726);
nor U3558 (N_3558,N_2700,N_2563);
nand U3559 (N_3559,N_2161,N_2440);
and U3560 (N_3560,N_2233,N_2659);
nor U3561 (N_3561,N_2086,N_2742);
nor U3562 (N_3562,N_2398,N_2912);
nand U3563 (N_3563,N_2953,N_2353);
nand U3564 (N_3564,N_2136,N_2979);
or U3565 (N_3565,N_2183,N_2210);
xor U3566 (N_3566,N_2098,N_2493);
nand U3567 (N_3567,N_2926,N_2056);
nand U3568 (N_3568,N_2351,N_2373);
or U3569 (N_3569,N_2952,N_2079);
or U3570 (N_3570,N_2014,N_2111);
or U3571 (N_3571,N_2724,N_2014);
or U3572 (N_3572,N_2433,N_2029);
and U3573 (N_3573,N_2755,N_2816);
nand U3574 (N_3574,N_2824,N_2325);
and U3575 (N_3575,N_2017,N_2171);
and U3576 (N_3576,N_2608,N_2019);
nor U3577 (N_3577,N_2498,N_2475);
nand U3578 (N_3578,N_2278,N_2488);
and U3579 (N_3579,N_2341,N_2576);
nand U3580 (N_3580,N_2892,N_2529);
nor U3581 (N_3581,N_2539,N_2015);
or U3582 (N_3582,N_2272,N_2760);
or U3583 (N_3583,N_2265,N_2447);
xor U3584 (N_3584,N_2173,N_2691);
nand U3585 (N_3585,N_2082,N_2514);
or U3586 (N_3586,N_2644,N_2685);
nand U3587 (N_3587,N_2800,N_2114);
or U3588 (N_3588,N_2527,N_2688);
nand U3589 (N_3589,N_2466,N_2229);
and U3590 (N_3590,N_2663,N_2345);
and U3591 (N_3591,N_2172,N_2088);
and U3592 (N_3592,N_2639,N_2426);
and U3593 (N_3593,N_2680,N_2053);
or U3594 (N_3594,N_2270,N_2193);
nand U3595 (N_3595,N_2165,N_2303);
nand U3596 (N_3596,N_2899,N_2599);
nor U3597 (N_3597,N_2720,N_2838);
nor U3598 (N_3598,N_2983,N_2161);
and U3599 (N_3599,N_2218,N_2346);
nor U3600 (N_3600,N_2959,N_2306);
nand U3601 (N_3601,N_2443,N_2088);
nand U3602 (N_3602,N_2255,N_2551);
and U3603 (N_3603,N_2593,N_2704);
nand U3604 (N_3604,N_2850,N_2634);
nor U3605 (N_3605,N_2371,N_2656);
and U3606 (N_3606,N_2667,N_2869);
nand U3607 (N_3607,N_2959,N_2146);
xor U3608 (N_3608,N_2167,N_2912);
nor U3609 (N_3609,N_2857,N_2513);
nand U3610 (N_3610,N_2468,N_2342);
nor U3611 (N_3611,N_2741,N_2489);
nor U3612 (N_3612,N_2665,N_2323);
xnor U3613 (N_3613,N_2755,N_2351);
nor U3614 (N_3614,N_2608,N_2818);
or U3615 (N_3615,N_2174,N_2477);
or U3616 (N_3616,N_2809,N_2102);
nor U3617 (N_3617,N_2225,N_2712);
nor U3618 (N_3618,N_2602,N_2678);
and U3619 (N_3619,N_2653,N_2427);
nor U3620 (N_3620,N_2897,N_2812);
nor U3621 (N_3621,N_2089,N_2082);
nor U3622 (N_3622,N_2777,N_2749);
or U3623 (N_3623,N_2712,N_2588);
nor U3624 (N_3624,N_2593,N_2737);
nor U3625 (N_3625,N_2966,N_2017);
nand U3626 (N_3626,N_2844,N_2254);
nor U3627 (N_3627,N_2229,N_2453);
or U3628 (N_3628,N_2314,N_2851);
nand U3629 (N_3629,N_2945,N_2874);
or U3630 (N_3630,N_2252,N_2574);
or U3631 (N_3631,N_2553,N_2519);
and U3632 (N_3632,N_2282,N_2965);
or U3633 (N_3633,N_2728,N_2804);
nor U3634 (N_3634,N_2000,N_2861);
nand U3635 (N_3635,N_2295,N_2029);
or U3636 (N_3636,N_2053,N_2211);
xnor U3637 (N_3637,N_2787,N_2146);
xnor U3638 (N_3638,N_2307,N_2289);
and U3639 (N_3639,N_2132,N_2742);
nor U3640 (N_3640,N_2058,N_2573);
or U3641 (N_3641,N_2808,N_2523);
nor U3642 (N_3642,N_2071,N_2155);
or U3643 (N_3643,N_2079,N_2398);
or U3644 (N_3644,N_2366,N_2144);
or U3645 (N_3645,N_2793,N_2233);
nor U3646 (N_3646,N_2762,N_2033);
nor U3647 (N_3647,N_2180,N_2274);
or U3648 (N_3648,N_2900,N_2442);
or U3649 (N_3649,N_2449,N_2650);
nand U3650 (N_3650,N_2423,N_2463);
or U3651 (N_3651,N_2208,N_2644);
nor U3652 (N_3652,N_2959,N_2125);
nand U3653 (N_3653,N_2796,N_2117);
nand U3654 (N_3654,N_2874,N_2498);
nand U3655 (N_3655,N_2201,N_2242);
and U3656 (N_3656,N_2956,N_2160);
xnor U3657 (N_3657,N_2507,N_2541);
and U3658 (N_3658,N_2419,N_2543);
or U3659 (N_3659,N_2829,N_2075);
or U3660 (N_3660,N_2131,N_2666);
or U3661 (N_3661,N_2724,N_2099);
and U3662 (N_3662,N_2325,N_2066);
nor U3663 (N_3663,N_2155,N_2838);
nand U3664 (N_3664,N_2752,N_2322);
nand U3665 (N_3665,N_2355,N_2585);
and U3666 (N_3666,N_2589,N_2716);
and U3667 (N_3667,N_2109,N_2113);
nand U3668 (N_3668,N_2855,N_2991);
nand U3669 (N_3669,N_2022,N_2556);
nor U3670 (N_3670,N_2272,N_2411);
or U3671 (N_3671,N_2540,N_2131);
nand U3672 (N_3672,N_2259,N_2748);
and U3673 (N_3673,N_2200,N_2325);
or U3674 (N_3674,N_2991,N_2394);
nand U3675 (N_3675,N_2614,N_2803);
nor U3676 (N_3676,N_2307,N_2724);
nand U3677 (N_3677,N_2030,N_2158);
nor U3678 (N_3678,N_2455,N_2776);
and U3679 (N_3679,N_2464,N_2229);
nand U3680 (N_3680,N_2849,N_2975);
xnor U3681 (N_3681,N_2334,N_2839);
nand U3682 (N_3682,N_2233,N_2116);
and U3683 (N_3683,N_2980,N_2586);
or U3684 (N_3684,N_2622,N_2970);
or U3685 (N_3685,N_2863,N_2008);
xnor U3686 (N_3686,N_2201,N_2232);
or U3687 (N_3687,N_2405,N_2903);
or U3688 (N_3688,N_2739,N_2467);
or U3689 (N_3689,N_2192,N_2398);
nor U3690 (N_3690,N_2232,N_2732);
xnor U3691 (N_3691,N_2017,N_2676);
or U3692 (N_3692,N_2024,N_2377);
and U3693 (N_3693,N_2659,N_2514);
nand U3694 (N_3694,N_2105,N_2409);
or U3695 (N_3695,N_2061,N_2238);
nor U3696 (N_3696,N_2690,N_2541);
and U3697 (N_3697,N_2970,N_2812);
nor U3698 (N_3698,N_2962,N_2789);
or U3699 (N_3699,N_2794,N_2550);
nand U3700 (N_3700,N_2530,N_2993);
or U3701 (N_3701,N_2121,N_2213);
or U3702 (N_3702,N_2232,N_2832);
and U3703 (N_3703,N_2630,N_2573);
nand U3704 (N_3704,N_2767,N_2134);
or U3705 (N_3705,N_2986,N_2749);
or U3706 (N_3706,N_2801,N_2245);
and U3707 (N_3707,N_2781,N_2471);
nand U3708 (N_3708,N_2096,N_2015);
and U3709 (N_3709,N_2595,N_2494);
and U3710 (N_3710,N_2450,N_2575);
nand U3711 (N_3711,N_2342,N_2544);
nor U3712 (N_3712,N_2939,N_2374);
nand U3713 (N_3713,N_2869,N_2423);
and U3714 (N_3714,N_2129,N_2702);
nand U3715 (N_3715,N_2545,N_2553);
nor U3716 (N_3716,N_2851,N_2226);
or U3717 (N_3717,N_2496,N_2999);
and U3718 (N_3718,N_2339,N_2079);
and U3719 (N_3719,N_2024,N_2758);
and U3720 (N_3720,N_2309,N_2212);
xor U3721 (N_3721,N_2149,N_2589);
nor U3722 (N_3722,N_2488,N_2232);
or U3723 (N_3723,N_2586,N_2758);
nand U3724 (N_3724,N_2286,N_2553);
or U3725 (N_3725,N_2956,N_2571);
or U3726 (N_3726,N_2775,N_2943);
or U3727 (N_3727,N_2471,N_2098);
or U3728 (N_3728,N_2552,N_2866);
nand U3729 (N_3729,N_2390,N_2475);
or U3730 (N_3730,N_2521,N_2004);
or U3731 (N_3731,N_2290,N_2688);
nor U3732 (N_3732,N_2217,N_2287);
nor U3733 (N_3733,N_2073,N_2305);
or U3734 (N_3734,N_2369,N_2956);
or U3735 (N_3735,N_2009,N_2996);
nand U3736 (N_3736,N_2390,N_2435);
and U3737 (N_3737,N_2194,N_2192);
or U3738 (N_3738,N_2708,N_2442);
nand U3739 (N_3739,N_2741,N_2943);
nor U3740 (N_3740,N_2730,N_2052);
nand U3741 (N_3741,N_2106,N_2172);
nor U3742 (N_3742,N_2417,N_2714);
nor U3743 (N_3743,N_2800,N_2129);
and U3744 (N_3744,N_2754,N_2984);
and U3745 (N_3745,N_2799,N_2729);
nor U3746 (N_3746,N_2541,N_2758);
or U3747 (N_3747,N_2355,N_2870);
or U3748 (N_3748,N_2617,N_2730);
or U3749 (N_3749,N_2805,N_2558);
nor U3750 (N_3750,N_2774,N_2597);
or U3751 (N_3751,N_2489,N_2440);
nor U3752 (N_3752,N_2551,N_2337);
and U3753 (N_3753,N_2102,N_2410);
nor U3754 (N_3754,N_2049,N_2812);
or U3755 (N_3755,N_2794,N_2704);
and U3756 (N_3756,N_2258,N_2892);
nor U3757 (N_3757,N_2003,N_2847);
and U3758 (N_3758,N_2857,N_2482);
or U3759 (N_3759,N_2959,N_2759);
nor U3760 (N_3760,N_2144,N_2200);
nor U3761 (N_3761,N_2847,N_2569);
or U3762 (N_3762,N_2670,N_2372);
nor U3763 (N_3763,N_2936,N_2725);
and U3764 (N_3764,N_2027,N_2879);
and U3765 (N_3765,N_2886,N_2487);
nand U3766 (N_3766,N_2619,N_2639);
or U3767 (N_3767,N_2258,N_2887);
or U3768 (N_3768,N_2747,N_2860);
and U3769 (N_3769,N_2302,N_2732);
or U3770 (N_3770,N_2820,N_2754);
nand U3771 (N_3771,N_2689,N_2387);
nor U3772 (N_3772,N_2482,N_2096);
nand U3773 (N_3773,N_2163,N_2624);
and U3774 (N_3774,N_2921,N_2811);
nand U3775 (N_3775,N_2744,N_2075);
and U3776 (N_3776,N_2803,N_2887);
nor U3777 (N_3777,N_2356,N_2878);
nor U3778 (N_3778,N_2336,N_2873);
nand U3779 (N_3779,N_2477,N_2595);
nand U3780 (N_3780,N_2703,N_2846);
or U3781 (N_3781,N_2498,N_2986);
nand U3782 (N_3782,N_2411,N_2752);
nor U3783 (N_3783,N_2040,N_2498);
xnor U3784 (N_3784,N_2349,N_2341);
nor U3785 (N_3785,N_2560,N_2240);
or U3786 (N_3786,N_2964,N_2329);
and U3787 (N_3787,N_2590,N_2373);
or U3788 (N_3788,N_2809,N_2478);
and U3789 (N_3789,N_2786,N_2421);
nor U3790 (N_3790,N_2977,N_2892);
or U3791 (N_3791,N_2292,N_2609);
nor U3792 (N_3792,N_2667,N_2277);
and U3793 (N_3793,N_2401,N_2951);
nand U3794 (N_3794,N_2681,N_2992);
and U3795 (N_3795,N_2467,N_2173);
and U3796 (N_3796,N_2902,N_2552);
or U3797 (N_3797,N_2249,N_2049);
nor U3798 (N_3798,N_2222,N_2194);
nor U3799 (N_3799,N_2946,N_2119);
nand U3800 (N_3800,N_2250,N_2811);
nor U3801 (N_3801,N_2150,N_2892);
nor U3802 (N_3802,N_2008,N_2518);
xnor U3803 (N_3803,N_2823,N_2447);
nor U3804 (N_3804,N_2034,N_2221);
or U3805 (N_3805,N_2907,N_2767);
or U3806 (N_3806,N_2085,N_2696);
nand U3807 (N_3807,N_2666,N_2314);
and U3808 (N_3808,N_2091,N_2930);
and U3809 (N_3809,N_2271,N_2480);
xnor U3810 (N_3810,N_2514,N_2655);
nand U3811 (N_3811,N_2147,N_2476);
or U3812 (N_3812,N_2115,N_2283);
nor U3813 (N_3813,N_2760,N_2972);
nor U3814 (N_3814,N_2353,N_2527);
nand U3815 (N_3815,N_2926,N_2490);
nor U3816 (N_3816,N_2427,N_2928);
xnor U3817 (N_3817,N_2388,N_2696);
nor U3818 (N_3818,N_2442,N_2727);
and U3819 (N_3819,N_2035,N_2918);
or U3820 (N_3820,N_2077,N_2640);
nand U3821 (N_3821,N_2750,N_2648);
nand U3822 (N_3822,N_2134,N_2939);
or U3823 (N_3823,N_2203,N_2486);
or U3824 (N_3824,N_2901,N_2964);
or U3825 (N_3825,N_2050,N_2965);
nor U3826 (N_3826,N_2787,N_2786);
nand U3827 (N_3827,N_2610,N_2792);
and U3828 (N_3828,N_2596,N_2824);
nor U3829 (N_3829,N_2021,N_2361);
and U3830 (N_3830,N_2077,N_2245);
and U3831 (N_3831,N_2868,N_2878);
or U3832 (N_3832,N_2042,N_2270);
nand U3833 (N_3833,N_2410,N_2942);
nand U3834 (N_3834,N_2468,N_2207);
nor U3835 (N_3835,N_2906,N_2162);
and U3836 (N_3836,N_2591,N_2030);
and U3837 (N_3837,N_2898,N_2503);
nor U3838 (N_3838,N_2741,N_2004);
nor U3839 (N_3839,N_2579,N_2190);
or U3840 (N_3840,N_2789,N_2902);
nand U3841 (N_3841,N_2178,N_2421);
nor U3842 (N_3842,N_2992,N_2564);
nand U3843 (N_3843,N_2553,N_2785);
nand U3844 (N_3844,N_2667,N_2351);
nand U3845 (N_3845,N_2484,N_2165);
and U3846 (N_3846,N_2598,N_2518);
and U3847 (N_3847,N_2185,N_2717);
nand U3848 (N_3848,N_2080,N_2658);
nor U3849 (N_3849,N_2960,N_2551);
nor U3850 (N_3850,N_2805,N_2404);
or U3851 (N_3851,N_2003,N_2357);
nor U3852 (N_3852,N_2944,N_2272);
nor U3853 (N_3853,N_2153,N_2852);
nor U3854 (N_3854,N_2394,N_2542);
nand U3855 (N_3855,N_2815,N_2215);
nor U3856 (N_3856,N_2851,N_2122);
or U3857 (N_3857,N_2566,N_2821);
nand U3858 (N_3858,N_2151,N_2175);
nor U3859 (N_3859,N_2622,N_2955);
nand U3860 (N_3860,N_2948,N_2151);
or U3861 (N_3861,N_2542,N_2184);
nand U3862 (N_3862,N_2290,N_2271);
or U3863 (N_3863,N_2653,N_2445);
nand U3864 (N_3864,N_2848,N_2412);
and U3865 (N_3865,N_2397,N_2248);
nand U3866 (N_3866,N_2383,N_2340);
and U3867 (N_3867,N_2857,N_2500);
nand U3868 (N_3868,N_2427,N_2895);
and U3869 (N_3869,N_2927,N_2708);
nor U3870 (N_3870,N_2478,N_2707);
nand U3871 (N_3871,N_2545,N_2964);
nor U3872 (N_3872,N_2461,N_2114);
nand U3873 (N_3873,N_2871,N_2411);
nor U3874 (N_3874,N_2686,N_2163);
nand U3875 (N_3875,N_2695,N_2725);
nand U3876 (N_3876,N_2476,N_2302);
and U3877 (N_3877,N_2317,N_2107);
nand U3878 (N_3878,N_2349,N_2954);
and U3879 (N_3879,N_2856,N_2855);
nor U3880 (N_3880,N_2289,N_2351);
nand U3881 (N_3881,N_2720,N_2775);
nand U3882 (N_3882,N_2778,N_2865);
or U3883 (N_3883,N_2126,N_2546);
nand U3884 (N_3884,N_2349,N_2374);
nor U3885 (N_3885,N_2071,N_2224);
and U3886 (N_3886,N_2406,N_2633);
or U3887 (N_3887,N_2271,N_2536);
nor U3888 (N_3888,N_2067,N_2944);
nor U3889 (N_3889,N_2717,N_2429);
or U3890 (N_3890,N_2399,N_2306);
nor U3891 (N_3891,N_2333,N_2541);
nand U3892 (N_3892,N_2083,N_2303);
and U3893 (N_3893,N_2127,N_2791);
nand U3894 (N_3894,N_2072,N_2977);
or U3895 (N_3895,N_2472,N_2699);
and U3896 (N_3896,N_2323,N_2683);
nor U3897 (N_3897,N_2836,N_2625);
nor U3898 (N_3898,N_2718,N_2120);
and U3899 (N_3899,N_2477,N_2193);
or U3900 (N_3900,N_2716,N_2905);
nor U3901 (N_3901,N_2542,N_2685);
nor U3902 (N_3902,N_2341,N_2605);
or U3903 (N_3903,N_2155,N_2762);
nand U3904 (N_3904,N_2181,N_2644);
and U3905 (N_3905,N_2955,N_2467);
nand U3906 (N_3906,N_2457,N_2507);
or U3907 (N_3907,N_2293,N_2446);
nand U3908 (N_3908,N_2475,N_2586);
and U3909 (N_3909,N_2396,N_2783);
xnor U3910 (N_3910,N_2986,N_2647);
nor U3911 (N_3911,N_2414,N_2039);
or U3912 (N_3912,N_2039,N_2773);
nor U3913 (N_3913,N_2332,N_2830);
or U3914 (N_3914,N_2348,N_2954);
and U3915 (N_3915,N_2022,N_2041);
nor U3916 (N_3916,N_2557,N_2894);
and U3917 (N_3917,N_2634,N_2191);
or U3918 (N_3918,N_2458,N_2541);
and U3919 (N_3919,N_2938,N_2489);
nor U3920 (N_3920,N_2331,N_2876);
nand U3921 (N_3921,N_2882,N_2447);
nor U3922 (N_3922,N_2199,N_2750);
nor U3923 (N_3923,N_2896,N_2328);
and U3924 (N_3924,N_2177,N_2723);
and U3925 (N_3925,N_2577,N_2983);
or U3926 (N_3926,N_2804,N_2280);
or U3927 (N_3927,N_2160,N_2506);
and U3928 (N_3928,N_2078,N_2141);
or U3929 (N_3929,N_2031,N_2797);
nor U3930 (N_3930,N_2458,N_2358);
and U3931 (N_3931,N_2744,N_2146);
and U3932 (N_3932,N_2030,N_2756);
and U3933 (N_3933,N_2085,N_2421);
or U3934 (N_3934,N_2952,N_2062);
or U3935 (N_3935,N_2599,N_2010);
and U3936 (N_3936,N_2630,N_2168);
nand U3937 (N_3937,N_2272,N_2697);
or U3938 (N_3938,N_2271,N_2498);
or U3939 (N_3939,N_2776,N_2183);
nand U3940 (N_3940,N_2316,N_2004);
and U3941 (N_3941,N_2978,N_2726);
and U3942 (N_3942,N_2629,N_2205);
or U3943 (N_3943,N_2699,N_2414);
and U3944 (N_3944,N_2341,N_2493);
or U3945 (N_3945,N_2684,N_2407);
and U3946 (N_3946,N_2496,N_2167);
or U3947 (N_3947,N_2963,N_2423);
nor U3948 (N_3948,N_2565,N_2016);
nor U3949 (N_3949,N_2140,N_2553);
or U3950 (N_3950,N_2173,N_2393);
or U3951 (N_3951,N_2333,N_2264);
nand U3952 (N_3952,N_2521,N_2363);
or U3953 (N_3953,N_2576,N_2156);
and U3954 (N_3954,N_2811,N_2693);
nor U3955 (N_3955,N_2155,N_2857);
or U3956 (N_3956,N_2838,N_2548);
or U3957 (N_3957,N_2557,N_2481);
nor U3958 (N_3958,N_2710,N_2600);
and U3959 (N_3959,N_2036,N_2088);
nand U3960 (N_3960,N_2523,N_2084);
or U3961 (N_3961,N_2007,N_2045);
and U3962 (N_3962,N_2433,N_2472);
or U3963 (N_3963,N_2576,N_2182);
nor U3964 (N_3964,N_2642,N_2180);
nand U3965 (N_3965,N_2027,N_2442);
or U3966 (N_3966,N_2003,N_2910);
and U3967 (N_3967,N_2426,N_2469);
or U3968 (N_3968,N_2583,N_2024);
nand U3969 (N_3969,N_2516,N_2534);
and U3970 (N_3970,N_2028,N_2811);
and U3971 (N_3971,N_2111,N_2260);
nand U3972 (N_3972,N_2453,N_2314);
and U3973 (N_3973,N_2927,N_2575);
or U3974 (N_3974,N_2195,N_2293);
nor U3975 (N_3975,N_2657,N_2682);
or U3976 (N_3976,N_2692,N_2942);
and U3977 (N_3977,N_2296,N_2495);
or U3978 (N_3978,N_2369,N_2303);
nor U3979 (N_3979,N_2006,N_2202);
nor U3980 (N_3980,N_2990,N_2707);
and U3981 (N_3981,N_2277,N_2151);
or U3982 (N_3982,N_2186,N_2866);
nor U3983 (N_3983,N_2275,N_2551);
and U3984 (N_3984,N_2505,N_2271);
and U3985 (N_3985,N_2304,N_2323);
nand U3986 (N_3986,N_2799,N_2109);
and U3987 (N_3987,N_2712,N_2881);
or U3988 (N_3988,N_2353,N_2025);
nand U3989 (N_3989,N_2885,N_2040);
nor U3990 (N_3990,N_2754,N_2903);
or U3991 (N_3991,N_2479,N_2011);
or U3992 (N_3992,N_2165,N_2602);
nand U3993 (N_3993,N_2139,N_2821);
or U3994 (N_3994,N_2858,N_2928);
nor U3995 (N_3995,N_2049,N_2443);
and U3996 (N_3996,N_2990,N_2384);
and U3997 (N_3997,N_2170,N_2952);
or U3998 (N_3998,N_2658,N_2937);
nand U3999 (N_3999,N_2163,N_2701);
nand U4000 (N_4000,N_3901,N_3629);
and U4001 (N_4001,N_3972,N_3923);
and U4002 (N_4002,N_3360,N_3110);
and U4003 (N_4003,N_3606,N_3068);
or U4004 (N_4004,N_3796,N_3251);
nor U4005 (N_4005,N_3113,N_3354);
nand U4006 (N_4006,N_3968,N_3844);
or U4007 (N_4007,N_3105,N_3032);
and U4008 (N_4008,N_3045,N_3866);
nor U4009 (N_4009,N_3975,N_3569);
nand U4010 (N_4010,N_3521,N_3567);
nor U4011 (N_4011,N_3978,N_3457);
and U4012 (N_4012,N_3682,N_3698);
and U4013 (N_4013,N_3845,N_3990);
nor U4014 (N_4014,N_3580,N_3283);
or U4015 (N_4015,N_3986,N_3545);
nor U4016 (N_4016,N_3822,N_3176);
and U4017 (N_4017,N_3753,N_3481);
and U4018 (N_4018,N_3670,N_3500);
and U4019 (N_4019,N_3074,N_3393);
or U4020 (N_4020,N_3755,N_3915);
nand U4021 (N_4021,N_3769,N_3138);
nor U4022 (N_4022,N_3296,N_3692);
and U4023 (N_4023,N_3136,N_3135);
and U4024 (N_4024,N_3498,N_3970);
and U4025 (N_4025,N_3873,N_3720);
and U4026 (N_4026,N_3163,N_3938);
or U4027 (N_4027,N_3904,N_3798);
nand U4028 (N_4028,N_3564,N_3727);
nand U4029 (N_4029,N_3106,N_3111);
and U4030 (N_4030,N_3322,N_3468);
or U4031 (N_4031,N_3932,N_3061);
and U4032 (N_4032,N_3784,N_3856);
nand U4033 (N_4033,N_3751,N_3674);
nor U4034 (N_4034,N_3718,N_3108);
and U4035 (N_4035,N_3897,N_3701);
nand U4036 (N_4036,N_3519,N_3369);
or U4037 (N_4037,N_3517,N_3615);
or U4038 (N_4038,N_3367,N_3792);
nand U4039 (N_4039,N_3793,N_3477);
and U4040 (N_4040,N_3593,N_3276);
nor U4041 (N_4041,N_3834,N_3683);
nand U4042 (N_4042,N_3955,N_3420);
nand U4043 (N_4043,N_3390,N_3401);
or U4044 (N_4044,N_3294,N_3435);
or U4045 (N_4045,N_3456,N_3903);
nor U4046 (N_4046,N_3402,N_3353);
and U4047 (N_4047,N_3054,N_3047);
nand U4048 (N_4048,N_3738,N_3756);
and U4049 (N_4049,N_3374,N_3744);
and U4050 (N_4050,N_3981,N_3359);
nor U4051 (N_4051,N_3413,N_3766);
or U4052 (N_4052,N_3969,N_3589);
xor U4053 (N_4053,N_3836,N_3781);
or U4054 (N_4054,N_3672,N_3247);
nand U4055 (N_4055,N_3802,N_3826);
and U4056 (N_4056,N_3710,N_3576);
and U4057 (N_4057,N_3308,N_3385);
and U4058 (N_4058,N_3151,N_3691);
nand U4059 (N_4059,N_3289,N_3243);
or U4060 (N_4060,N_3381,N_3510);
and U4061 (N_4061,N_3333,N_3134);
nand U4062 (N_4062,N_3819,N_3741);
or U4063 (N_4063,N_3869,N_3592);
nor U4064 (N_4064,N_3697,N_3795);
nor U4065 (N_4065,N_3411,N_3088);
or U4066 (N_4066,N_3528,N_3488);
nor U4067 (N_4067,N_3315,N_3408);
nor U4068 (N_4068,N_3542,N_3320);
nor U4069 (N_4069,N_3258,N_3570);
or U4070 (N_4070,N_3987,N_3616);
nand U4071 (N_4071,N_3638,N_3448);
nor U4072 (N_4072,N_3817,N_3870);
and U4073 (N_4073,N_3996,N_3187);
nand U4074 (N_4074,N_3452,N_3478);
nand U4075 (N_4075,N_3582,N_3806);
and U4076 (N_4076,N_3234,N_3807);
nor U4077 (N_4077,N_3335,N_3921);
nor U4078 (N_4078,N_3330,N_3036);
and U4079 (N_4079,N_3416,N_3573);
or U4080 (N_4080,N_3131,N_3679);
and U4081 (N_4081,N_3703,N_3167);
or U4082 (N_4082,N_3022,N_3365);
or U4083 (N_4083,N_3208,N_3862);
and U4084 (N_4084,N_3801,N_3958);
or U4085 (N_4085,N_3148,N_3891);
and U4086 (N_4086,N_3377,N_3746);
nor U4087 (N_4087,N_3336,N_3998);
xnor U4088 (N_4088,N_3613,N_3070);
or U4089 (N_4089,N_3577,N_3889);
and U4090 (N_4090,N_3091,N_3715);
nor U4091 (N_4091,N_3306,N_3145);
or U4092 (N_4092,N_3585,N_3757);
and U4093 (N_4093,N_3497,N_3042);
and U4094 (N_4094,N_3493,N_3415);
nor U4095 (N_4095,N_3546,N_3052);
or U4096 (N_4096,N_3489,N_3737);
and U4097 (N_4097,N_3527,N_3681);
or U4098 (N_4098,N_3641,N_3455);
and U4099 (N_4099,N_3121,N_3168);
or U4100 (N_4100,N_3021,N_3763);
and U4101 (N_4101,N_3877,N_3395);
nand U4102 (N_4102,N_3098,N_3890);
and U4103 (N_4103,N_3103,N_3093);
nor U4104 (N_4104,N_3449,N_3874);
and U4105 (N_4105,N_3038,N_3094);
or U4106 (N_4106,N_3946,N_3706);
nor U4107 (N_4107,N_3699,N_3494);
nor U4108 (N_4108,N_3730,N_3438);
nor U4109 (N_4109,N_3409,N_3848);
or U4110 (N_4110,N_3568,N_3442);
nand U4111 (N_4111,N_3140,N_3952);
and U4112 (N_4112,N_3941,N_3599);
or U4113 (N_4113,N_3429,N_3329);
nand U4114 (N_4114,N_3099,N_3123);
nand U4115 (N_4115,N_3624,N_3398);
nand U4116 (N_4116,N_3547,N_3198);
xnor U4117 (N_4117,N_3112,N_3752);
xor U4118 (N_4118,N_3403,N_3461);
nand U4119 (N_4119,N_3153,N_3551);
or U4120 (N_4120,N_3314,N_3013);
and U4121 (N_4121,N_3612,N_3159);
or U4122 (N_4122,N_3900,N_3799);
nand U4123 (N_4123,N_3383,N_3646);
and U4124 (N_4124,N_3973,N_3954);
nor U4125 (N_4125,N_3120,N_3876);
and U4126 (N_4126,N_3345,N_3885);
xor U4127 (N_4127,N_3609,N_3273);
xnor U4128 (N_4128,N_3685,N_3522);
nand U4129 (N_4129,N_3237,N_3157);
nor U4130 (N_4130,N_3161,N_3927);
or U4131 (N_4131,N_3963,N_3808);
nand U4132 (N_4132,N_3195,N_3643);
nand U4133 (N_4133,N_3141,N_3201);
nor U4134 (N_4134,N_3989,N_3884);
nor U4135 (N_4135,N_3150,N_3464);
and U4136 (N_4136,N_3666,N_3266);
and U4137 (N_4137,N_3003,N_3469);
nor U4138 (N_4138,N_3172,N_3248);
nand U4139 (N_4139,N_3083,N_3236);
xnor U4140 (N_4140,N_3827,N_3950);
or U4141 (N_4141,N_3858,N_3122);
and U4142 (N_4142,N_3199,N_3659);
and U4143 (N_4143,N_3011,N_3774);
nor U4144 (N_4144,N_3561,N_3653);
nand U4145 (N_4145,N_3541,N_3770);
and U4146 (N_4146,N_3081,N_3964);
or U4147 (N_4147,N_3439,N_3450);
or U4148 (N_4148,N_3611,N_3747);
and U4149 (N_4149,N_3942,N_3531);
nor U4150 (N_4150,N_3832,N_3344);
nor U4151 (N_4151,N_3290,N_3212);
or U4152 (N_4152,N_3888,N_3459);
or U4153 (N_4153,N_3282,N_3017);
nor U4154 (N_4154,N_3860,N_3684);
and U4155 (N_4155,N_3244,N_3279);
or U4156 (N_4156,N_3667,N_3712);
and U4157 (N_4157,N_3125,N_3914);
or U4158 (N_4158,N_3265,N_3355);
nor U4159 (N_4159,N_3905,N_3332);
nor U4160 (N_4160,N_3171,N_3264);
and U4161 (N_4161,N_3441,N_3132);
and U4162 (N_4162,N_3233,N_3060);
and U4163 (N_4163,N_3484,N_3767);
and U4164 (N_4164,N_3286,N_3959);
xor U4165 (N_4165,N_3924,N_3312);
nand U4166 (N_4166,N_3508,N_3118);
nor U4167 (N_4167,N_3217,N_3940);
nor U4168 (N_4168,N_3626,N_3086);
and U4169 (N_4169,N_3104,N_3254);
nand U4170 (N_4170,N_3392,N_3949);
nor U4171 (N_4171,N_3039,N_3048);
nor U4172 (N_4172,N_3040,N_3533);
nor U4173 (N_4173,N_3584,N_3049);
nor U4174 (N_4174,N_3544,N_3700);
and U4175 (N_4175,N_3421,N_3944);
or U4176 (N_4176,N_3278,N_3370);
and U4177 (N_4177,N_3215,N_3075);
and U4178 (N_4178,N_3100,N_3102);
and U4179 (N_4179,N_3407,N_3334);
or U4180 (N_4180,N_3852,N_3230);
nand U4181 (N_4181,N_3337,N_3078);
and U4182 (N_4182,N_3902,N_3444);
or U4183 (N_4183,N_3768,N_3661);
nand U4184 (N_4184,N_3688,N_3879);
nand U4185 (N_4185,N_3809,N_3499);
and U4186 (N_4186,N_3341,N_3053);
nor U4187 (N_4187,N_3027,N_3779);
nor U4188 (N_4188,N_3956,N_3200);
or U4189 (N_4189,N_3675,N_3384);
nor U4190 (N_4190,N_3908,N_3622);
and U4191 (N_4191,N_3197,N_3705);
nor U4192 (N_4192,N_3175,N_3490);
nand U4193 (N_4193,N_3304,N_3742);
and U4194 (N_4194,N_3831,N_3257);
xor U4195 (N_4195,N_3635,N_3250);
or U4196 (N_4196,N_3919,N_3910);
and U4197 (N_4197,N_3361,N_3620);
and U4198 (N_4198,N_3191,N_3300);
xor U4199 (N_4199,N_3658,N_3604);
or U4200 (N_4200,N_3400,N_3911);
and U4201 (N_4201,N_3818,N_3758);
or U4202 (N_4202,N_3850,N_3841);
nand U4203 (N_4203,N_3591,N_3028);
nor U4204 (N_4204,N_3026,N_3227);
or U4205 (N_4205,N_3595,N_3479);
nor U4206 (N_4206,N_3553,N_3980);
and U4207 (N_4207,N_3581,N_3431);
nor U4208 (N_4208,N_3324,N_3565);
nor U4209 (N_4209,N_3596,N_3548);
nand U4210 (N_4210,N_3926,N_3824);
and U4211 (N_4211,N_3302,N_3443);
nor U4212 (N_4212,N_3472,N_3023);
or U4213 (N_4213,N_3694,N_3607);
and U4214 (N_4214,N_3260,N_3405);
nor U4215 (N_4215,N_3109,N_3614);
or U4216 (N_4216,N_3480,N_3645);
nand U4217 (N_4217,N_3292,N_3843);
nor U4218 (N_4218,N_3909,N_3853);
nor U4219 (N_4219,N_3886,N_3967);
nor U4220 (N_4220,N_3433,N_3186);
nor U4221 (N_4221,N_3647,N_3644);
nand U4222 (N_4222,N_3539,N_3155);
or U4223 (N_4223,N_3739,N_3864);
or U4224 (N_4224,N_3363,N_3725);
nand U4225 (N_4225,N_3487,N_3812);
and U4226 (N_4226,N_3673,N_3029);
nor U4227 (N_4227,N_3339,N_3437);
nand U4228 (N_4228,N_3868,N_3055);
and U4229 (N_4229,N_3702,N_3291);
nand U4230 (N_4230,N_3242,N_3623);
nor U4231 (N_4231,N_3976,N_3496);
or U4232 (N_4232,N_3253,N_3765);
and U4233 (N_4233,N_3618,N_3693);
or U4234 (N_4234,N_3997,N_3880);
nand U4235 (N_4235,N_3636,N_3628);
nor U4236 (N_4236,N_3837,N_3209);
and U4237 (N_4237,N_3371,N_3759);
nand U4238 (N_4238,N_3362,N_3096);
or U4239 (N_4239,N_3979,N_3351);
nand U4240 (N_4240,N_3259,N_3139);
and U4241 (N_4241,N_3610,N_3313);
nor U4242 (N_4242,N_3662,N_3695);
nor U4243 (N_4243,N_3358,N_3617);
or U4244 (N_4244,N_3419,N_3085);
and U4245 (N_4245,N_3722,N_3648);
and U4246 (N_4246,N_3147,N_3734);
nor U4247 (N_4247,N_3503,N_3925);
nand U4248 (N_4248,N_3960,N_3937);
and U4249 (N_4249,N_3930,N_3660);
nor U4250 (N_4250,N_3557,N_3426);
nor U4251 (N_4251,N_3872,N_3238);
or U4252 (N_4252,N_3019,N_3931);
or U4253 (N_4253,N_3422,N_3424);
nor U4254 (N_4254,N_3458,N_3632);
nor U4255 (N_4255,N_3000,N_3775);
nor U4256 (N_4256,N_3318,N_3284);
xor U4257 (N_4257,N_3562,N_3537);
nand U4258 (N_4258,N_3387,N_3597);
nand U4259 (N_4259,N_3764,N_3847);
or U4260 (N_4260,N_3263,N_3368);
nor U4261 (N_4261,N_3785,N_3310);
and U4262 (N_4262,N_3550,N_3740);
or U4263 (N_4263,N_3031,N_3811);
nor U4264 (N_4264,N_3440,N_3823);
nand U4265 (N_4265,N_3579,N_3182);
nand U4266 (N_4266,N_3446,N_3948);
nor U4267 (N_4267,N_3035,N_3771);
and U4268 (N_4268,N_3729,N_3530);
and U4269 (N_4269,N_3605,N_3558);
or U4270 (N_4270,N_3838,N_3721);
xor U4271 (N_4271,N_3087,N_3736);
nor U4272 (N_4272,N_3297,N_3945);
or U4273 (N_4273,N_3574,N_3192);
or U4274 (N_4274,N_3575,N_3277);
nand U4275 (N_4275,N_3507,N_3486);
or U4276 (N_4276,N_3214,N_3231);
or U4277 (N_4277,N_3995,N_3092);
xnor U4278 (N_4278,N_3194,N_3057);
and U4279 (N_4279,N_3012,N_3878);
nand U4280 (N_4280,N_3229,N_3349);
nand U4281 (N_4281,N_3514,N_3689);
or U4282 (N_4282,N_3654,N_3893);
or U4283 (N_4283,N_3492,N_3495);
nand U4284 (N_4284,N_3177,N_3883);
nor U4285 (N_4285,N_3301,N_3482);
or U4286 (N_4286,N_3239,N_3603);
nor U4287 (N_4287,N_3228,N_3154);
or U4288 (N_4288,N_3529,N_3166);
and U4289 (N_4289,N_3509,N_3114);
and U4290 (N_4290,N_3745,N_3571);
nand U4291 (N_4291,N_3786,N_3828);
or U4292 (N_4292,N_3261,N_3916);
and U4293 (N_4293,N_3906,N_3887);
and U4294 (N_4294,N_3476,N_3224);
nand U4295 (N_4295,N_3203,N_3071);
and U4296 (N_4296,N_3327,N_3241);
or U4297 (N_4297,N_3193,N_3379);
nor U4298 (N_4298,N_3156,N_3311);
and U4299 (N_4299,N_3185,N_3144);
nor U4300 (N_4300,N_3412,N_3555);
and U4301 (N_4301,N_3563,N_3044);
nand U4302 (N_4302,N_3274,N_3732);
nand U4303 (N_4303,N_3414,N_3994);
or U4304 (N_4304,N_3714,N_3307);
or U4305 (N_4305,N_3829,N_3350);
or U4306 (N_4306,N_3762,N_3898);
nor U4307 (N_4307,N_3119,N_3189);
or U4308 (N_4308,N_3303,N_3338);
and U4309 (N_4309,N_3268,N_3041);
nand U4310 (N_4310,N_3859,N_3833);
and U4311 (N_4311,N_3184,N_3787);
nand U4312 (N_4312,N_3825,N_3309);
or U4313 (N_4313,N_3221,N_3583);
nor U4314 (N_4314,N_3116,N_3525);
and U4315 (N_4315,N_3957,N_3892);
and U4316 (N_4316,N_3608,N_3735);
or U4317 (N_4317,N_3418,N_3373);
and U4318 (N_4318,N_3552,N_3559);
nand U4319 (N_4319,N_3578,N_3406);
or U4320 (N_4320,N_3849,N_3634);
or U4321 (N_4321,N_3272,N_3206);
or U4322 (N_4322,N_3881,N_3470);
nor U4323 (N_4323,N_3164,N_3137);
nand U4324 (N_4324,N_3066,N_3475);
nor U4325 (N_4325,N_3502,N_3707);
and U4326 (N_4326,N_3839,N_3204);
nor U4327 (N_4327,N_3375,N_3077);
nand U4328 (N_4328,N_3394,N_3115);
and U4329 (N_4329,N_3471,N_3984);
and U4330 (N_4330,N_3804,N_3665);
nor U4331 (N_4331,N_3343,N_3999);
and U4332 (N_4332,N_3162,N_3907);
nand U4333 (N_4333,N_3299,N_3222);
or U4334 (N_4334,N_3271,N_3328);
nor U4335 (N_4335,N_3962,N_3025);
nor U4336 (N_4336,N_3621,N_3983);
or U4337 (N_4337,N_3467,N_3794);
and U4338 (N_4338,N_3971,N_3797);
nand U4339 (N_4339,N_3535,N_3965);
and U4340 (N_4340,N_3639,N_3778);
nor U4341 (N_4341,N_3425,N_3226);
nand U4342 (N_4342,N_3427,N_3046);
or U4343 (N_4343,N_3002,N_3953);
nand U4344 (N_4344,N_3505,N_3196);
and U4345 (N_4345,N_3451,N_3010);
and U4346 (N_4346,N_3678,N_3586);
or U4347 (N_4347,N_3602,N_3388);
nor U4348 (N_4348,N_3939,N_3922);
or U4349 (N_4349,N_3249,N_3174);
nor U4350 (N_4350,N_3269,N_3202);
nand U4351 (N_4351,N_3669,N_3149);
nor U4352 (N_4352,N_3788,N_3076);
and U4353 (N_4353,N_3245,N_3783);
nor U4354 (N_4354,N_3178,N_3319);
nor U4355 (N_4355,N_3287,N_3773);
and U4356 (N_4356,N_3594,N_3225);
or U4357 (N_4357,N_3107,N_3777);
nand U4358 (N_4358,N_3170,N_3504);
and U4359 (N_4359,N_3072,N_3985);
and U4360 (N_4360,N_3380,N_3912);
xor U4361 (N_4361,N_3992,N_3625);
and U4362 (N_4362,N_3899,N_3356);
nand U4363 (N_4363,N_3453,N_3855);
nor U4364 (N_4364,N_3124,N_3724);
and U4365 (N_4365,N_3791,N_3513);
nor U4366 (N_4366,N_3761,N_3275);
nand U4367 (N_4367,N_3929,N_3235);
nand U4368 (N_4368,N_3428,N_3895);
nand U4369 (N_4369,N_3947,N_3396);
nand U4370 (N_4370,N_3445,N_3749);
nand U4371 (N_4371,N_3117,N_3127);
or U4372 (N_4372,N_3821,N_3656);
nor U4373 (N_4373,N_3520,N_3090);
nand U4374 (N_4374,N_3460,N_3340);
or U4375 (N_4375,N_3917,N_3524);
nand U4376 (N_4376,N_3378,N_3295);
or U4377 (N_4377,N_3423,N_3095);
or U4378 (N_4378,N_3627,N_3084);
nand U4379 (N_4379,N_3069,N_3058);
nor U4380 (N_4380,N_3007,N_3814);
and U4381 (N_4381,N_3005,N_3820);
nand U4382 (N_4382,N_3491,N_3160);
and U4383 (N_4383,N_3101,N_3650);
nand U4384 (N_4384,N_3943,N_3326);
and U4385 (N_4385,N_3642,N_3130);
nand U4386 (N_4386,N_3894,N_3432);
and U4387 (N_4387,N_3165,N_3861);
nand U4388 (N_4388,N_3065,N_3073);
nand U4389 (N_4389,N_3213,N_3466);
xnor U4390 (N_4390,N_3686,N_3668);
or U4391 (N_4391,N_3006,N_3079);
nor U4392 (N_4392,N_3754,N_3216);
nand U4393 (N_4393,N_3713,N_3974);
nor U4394 (N_4394,N_3928,N_3372);
nand U4395 (N_4395,N_3267,N_3549);
or U4396 (N_4396,N_3346,N_3382);
and U4397 (N_4397,N_3803,N_3146);
nand U4398 (N_4398,N_3810,N_3731);
nand U4399 (N_4399,N_3474,N_3342);
nand U4400 (N_4400,N_3205,N_3728);
and U4401 (N_4401,N_3410,N_3704);
xnor U4402 (N_4402,N_3142,N_3252);
nand U4403 (N_4403,N_3554,N_3780);
and U4404 (N_4404,N_3158,N_3321);
nand U4405 (N_4405,N_3056,N_3867);
nand U4406 (N_4406,N_3188,N_3434);
and U4407 (N_4407,N_3436,N_3128);
nor U4408 (N_4408,N_3256,N_3080);
nand U4409 (N_4409,N_3133,N_3364);
nand U4410 (N_4410,N_3951,N_3050);
and U4411 (N_4411,N_3063,N_3454);
or U4412 (N_4412,N_3143,N_3001);
and U4413 (N_4413,N_3210,N_3920);
nand U4414 (N_4414,N_3566,N_3357);
and U4415 (N_4415,N_3572,N_3220);
nor U4416 (N_4416,N_3316,N_3966);
nor U4417 (N_4417,N_3556,N_3536);
nand U4418 (N_4418,N_3386,N_3207);
and U4419 (N_4419,N_3211,N_3232);
nor U4420 (N_4420,N_3936,N_3181);
and U4421 (N_4421,N_3726,N_3750);
nor U4422 (N_4422,N_3863,N_3716);
nor U4423 (N_4423,N_3082,N_3179);
and U4424 (N_4424,N_3598,N_3851);
and U4425 (N_4425,N_3991,N_3298);
and U4426 (N_4426,N_3352,N_3501);
and U4427 (N_4427,N_3523,N_3323);
or U4428 (N_4428,N_3218,N_3588);
and U4429 (N_4429,N_3652,N_3180);
xnor U4430 (N_4430,N_3526,N_3748);
nor U4431 (N_4431,N_3590,N_3875);
and U4432 (N_4432,N_3717,N_3516);
nand U4433 (N_4433,N_3782,N_3173);
or U4434 (N_4434,N_3865,N_3913);
or U4435 (N_4435,N_3776,N_3034);
nor U4436 (N_4436,N_3018,N_3015);
nand U4437 (N_4437,N_3815,N_3033);
xnor U4438 (N_4438,N_3262,N_3677);
and U4439 (N_4439,N_3089,N_3240);
and U4440 (N_4440,N_3934,N_3534);
or U4441 (N_4441,N_3657,N_3982);
and U4442 (N_4442,N_3655,N_3835);
nor U4443 (N_4443,N_3830,N_3465);
and U4444 (N_4444,N_3709,N_3399);
nand U4445 (N_4445,N_3511,N_3126);
nor U4446 (N_4446,N_3169,N_3671);
and U4447 (N_4447,N_3760,N_3772);
xor U4448 (N_4448,N_3462,N_3918);
nand U4449 (N_4449,N_3067,N_3030);
nor U4450 (N_4450,N_3430,N_3348);
nor U4451 (N_4451,N_3518,N_3037);
nand U4452 (N_4452,N_3532,N_3014);
and U4453 (N_4453,N_3325,N_3649);
nand U4454 (N_4454,N_3871,N_3246);
nand U4455 (N_4455,N_3854,N_3270);
and U4456 (N_4456,N_3129,N_3619);
nor U4457 (N_4457,N_3483,N_3664);
nor U4458 (N_4458,N_3933,N_3506);
or U4459 (N_4459,N_3059,N_3285);
nor U4460 (N_4460,N_3538,N_3813);
or U4461 (N_4461,N_3255,N_3447);
xor U4462 (N_4462,N_3687,N_3417);
and U4463 (N_4463,N_3711,N_3663);
xor U4464 (N_4464,N_3281,N_3977);
or U4465 (N_4465,N_3543,N_3800);
nor U4466 (N_4466,N_3600,N_3840);
xnor U4467 (N_4467,N_3631,N_3391);
or U4468 (N_4468,N_3016,N_3293);
xor U4469 (N_4469,N_3882,N_3690);
nand U4470 (N_4470,N_3183,N_3024);
nand U4471 (N_4471,N_3004,N_3305);
or U4472 (N_4472,N_3789,N_3988);
nand U4473 (N_4473,N_3723,N_3708);
xnor U4474 (N_4474,N_3935,N_3601);
nand U4475 (N_4475,N_3331,N_3009);
nor U4476 (N_4476,N_3317,N_3630);
xor U4477 (N_4477,N_3397,N_3680);
or U4478 (N_4478,N_3463,N_3280);
or U4479 (N_4479,N_3540,N_3719);
and U4480 (N_4480,N_3376,N_3473);
or U4481 (N_4481,N_3790,N_3051);
nor U4482 (N_4482,N_3020,N_3857);
and U4483 (N_4483,N_3223,N_3515);
or U4484 (N_4484,N_3676,N_3062);
nor U4485 (N_4485,N_3560,N_3733);
nand U4486 (N_4486,N_3190,N_3640);
or U4487 (N_4487,N_3961,N_3097);
nand U4488 (N_4488,N_3389,N_3366);
nor U4489 (N_4489,N_3637,N_3485);
nand U4490 (N_4490,N_3743,N_3043);
nor U4491 (N_4491,N_3993,N_3696);
or U4492 (N_4492,N_3512,N_3896);
or U4493 (N_4493,N_3008,N_3633);
nand U4494 (N_4494,N_3842,N_3651);
nor U4495 (N_4495,N_3805,N_3152);
and U4496 (N_4496,N_3846,N_3587);
nor U4497 (N_4497,N_3219,N_3064);
and U4498 (N_4498,N_3347,N_3288);
nor U4499 (N_4499,N_3404,N_3816);
and U4500 (N_4500,N_3493,N_3903);
and U4501 (N_4501,N_3523,N_3476);
nand U4502 (N_4502,N_3600,N_3736);
nand U4503 (N_4503,N_3314,N_3832);
nand U4504 (N_4504,N_3227,N_3553);
and U4505 (N_4505,N_3733,N_3476);
nand U4506 (N_4506,N_3984,N_3978);
or U4507 (N_4507,N_3705,N_3921);
or U4508 (N_4508,N_3552,N_3505);
xnor U4509 (N_4509,N_3379,N_3525);
and U4510 (N_4510,N_3807,N_3020);
nor U4511 (N_4511,N_3210,N_3162);
nor U4512 (N_4512,N_3294,N_3765);
nand U4513 (N_4513,N_3467,N_3904);
and U4514 (N_4514,N_3149,N_3908);
and U4515 (N_4515,N_3462,N_3015);
or U4516 (N_4516,N_3050,N_3467);
nand U4517 (N_4517,N_3825,N_3667);
nor U4518 (N_4518,N_3131,N_3259);
nand U4519 (N_4519,N_3170,N_3930);
nand U4520 (N_4520,N_3236,N_3456);
nor U4521 (N_4521,N_3330,N_3332);
or U4522 (N_4522,N_3608,N_3554);
xnor U4523 (N_4523,N_3640,N_3262);
nand U4524 (N_4524,N_3918,N_3788);
or U4525 (N_4525,N_3026,N_3557);
and U4526 (N_4526,N_3156,N_3099);
nand U4527 (N_4527,N_3244,N_3822);
or U4528 (N_4528,N_3262,N_3844);
or U4529 (N_4529,N_3681,N_3399);
or U4530 (N_4530,N_3815,N_3864);
nand U4531 (N_4531,N_3211,N_3369);
nand U4532 (N_4532,N_3781,N_3503);
nand U4533 (N_4533,N_3389,N_3655);
nor U4534 (N_4534,N_3397,N_3629);
nand U4535 (N_4535,N_3495,N_3774);
or U4536 (N_4536,N_3968,N_3658);
and U4537 (N_4537,N_3682,N_3446);
or U4538 (N_4538,N_3386,N_3157);
or U4539 (N_4539,N_3217,N_3393);
nor U4540 (N_4540,N_3362,N_3953);
or U4541 (N_4541,N_3285,N_3684);
or U4542 (N_4542,N_3730,N_3617);
or U4543 (N_4543,N_3951,N_3129);
nand U4544 (N_4544,N_3122,N_3732);
xnor U4545 (N_4545,N_3877,N_3114);
xnor U4546 (N_4546,N_3463,N_3593);
or U4547 (N_4547,N_3115,N_3112);
and U4548 (N_4548,N_3783,N_3273);
nor U4549 (N_4549,N_3990,N_3701);
or U4550 (N_4550,N_3074,N_3717);
nand U4551 (N_4551,N_3496,N_3012);
nor U4552 (N_4552,N_3024,N_3934);
and U4553 (N_4553,N_3025,N_3872);
nand U4554 (N_4554,N_3047,N_3529);
nand U4555 (N_4555,N_3147,N_3962);
and U4556 (N_4556,N_3491,N_3013);
nand U4557 (N_4557,N_3410,N_3085);
or U4558 (N_4558,N_3709,N_3927);
xnor U4559 (N_4559,N_3069,N_3286);
or U4560 (N_4560,N_3274,N_3183);
or U4561 (N_4561,N_3514,N_3616);
nand U4562 (N_4562,N_3730,N_3502);
and U4563 (N_4563,N_3487,N_3230);
nor U4564 (N_4564,N_3043,N_3132);
and U4565 (N_4565,N_3966,N_3291);
and U4566 (N_4566,N_3945,N_3015);
and U4567 (N_4567,N_3924,N_3076);
nor U4568 (N_4568,N_3539,N_3846);
nand U4569 (N_4569,N_3836,N_3164);
nand U4570 (N_4570,N_3577,N_3107);
nand U4571 (N_4571,N_3273,N_3884);
nand U4572 (N_4572,N_3614,N_3968);
or U4573 (N_4573,N_3752,N_3929);
nand U4574 (N_4574,N_3564,N_3439);
and U4575 (N_4575,N_3936,N_3982);
nand U4576 (N_4576,N_3536,N_3844);
or U4577 (N_4577,N_3756,N_3031);
or U4578 (N_4578,N_3631,N_3523);
nor U4579 (N_4579,N_3206,N_3580);
nor U4580 (N_4580,N_3479,N_3011);
nand U4581 (N_4581,N_3649,N_3148);
nand U4582 (N_4582,N_3841,N_3995);
and U4583 (N_4583,N_3509,N_3125);
or U4584 (N_4584,N_3581,N_3425);
and U4585 (N_4585,N_3370,N_3004);
or U4586 (N_4586,N_3373,N_3269);
nand U4587 (N_4587,N_3607,N_3750);
and U4588 (N_4588,N_3101,N_3187);
or U4589 (N_4589,N_3648,N_3052);
or U4590 (N_4590,N_3696,N_3683);
and U4591 (N_4591,N_3708,N_3942);
or U4592 (N_4592,N_3669,N_3880);
and U4593 (N_4593,N_3367,N_3817);
nor U4594 (N_4594,N_3613,N_3862);
nand U4595 (N_4595,N_3473,N_3909);
and U4596 (N_4596,N_3336,N_3600);
xnor U4597 (N_4597,N_3900,N_3590);
nor U4598 (N_4598,N_3449,N_3750);
and U4599 (N_4599,N_3470,N_3093);
nand U4600 (N_4600,N_3092,N_3303);
or U4601 (N_4601,N_3452,N_3544);
and U4602 (N_4602,N_3352,N_3379);
and U4603 (N_4603,N_3492,N_3791);
and U4604 (N_4604,N_3619,N_3437);
nor U4605 (N_4605,N_3560,N_3008);
nand U4606 (N_4606,N_3147,N_3463);
nor U4607 (N_4607,N_3935,N_3365);
nor U4608 (N_4608,N_3662,N_3777);
and U4609 (N_4609,N_3855,N_3738);
nand U4610 (N_4610,N_3956,N_3401);
or U4611 (N_4611,N_3573,N_3935);
nor U4612 (N_4612,N_3464,N_3535);
nor U4613 (N_4613,N_3001,N_3519);
or U4614 (N_4614,N_3384,N_3702);
or U4615 (N_4615,N_3288,N_3757);
or U4616 (N_4616,N_3184,N_3680);
and U4617 (N_4617,N_3438,N_3736);
or U4618 (N_4618,N_3408,N_3055);
nor U4619 (N_4619,N_3901,N_3336);
nand U4620 (N_4620,N_3680,N_3603);
and U4621 (N_4621,N_3242,N_3267);
or U4622 (N_4622,N_3598,N_3323);
and U4623 (N_4623,N_3273,N_3500);
or U4624 (N_4624,N_3428,N_3495);
or U4625 (N_4625,N_3948,N_3356);
nand U4626 (N_4626,N_3561,N_3771);
xnor U4627 (N_4627,N_3924,N_3130);
or U4628 (N_4628,N_3544,N_3054);
nor U4629 (N_4629,N_3552,N_3107);
and U4630 (N_4630,N_3700,N_3314);
nor U4631 (N_4631,N_3848,N_3118);
or U4632 (N_4632,N_3661,N_3104);
nand U4633 (N_4633,N_3693,N_3830);
nand U4634 (N_4634,N_3117,N_3756);
nor U4635 (N_4635,N_3877,N_3917);
and U4636 (N_4636,N_3544,N_3567);
and U4637 (N_4637,N_3699,N_3031);
or U4638 (N_4638,N_3214,N_3850);
and U4639 (N_4639,N_3294,N_3061);
nor U4640 (N_4640,N_3974,N_3102);
or U4641 (N_4641,N_3891,N_3144);
and U4642 (N_4642,N_3254,N_3206);
xnor U4643 (N_4643,N_3632,N_3952);
or U4644 (N_4644,N_3250,N_3140);
or U4645 (N_4645,N_3196,N_3923);
nand U4646 (N_4646,N_3527,N_3644);
or U4647 (N_4647,N_3542,N_3444);
or U4648 (N_4648,N_3936,N_3742);
nand U4649 (N_4649,N_3873,N_3001);
nand U4650 (N_4650,N_3343,N_3992);
and U4651 (N_4651,N_3091,N_3787);
and U4652 (N_4652,N_3830,N_3366);
nor U4653 (N_4653,N_3681,N_3165);
and U4654 (N_4654,N_3574,N_3289);
and U4655 (N_4655,N_3440,N_3389);
or U4656 (N_4656,N_3677,N_3480);
or U4657 (N_4657,N_3542,N_3877);
or U4658 (N_4658,N_3613,N_3361);
and U4659 (N_4659,N_3085,N_3201);
or U4660 (N_4660,N_3221,N_3272);
nor U4661 (N_4661,N_3640,N_3566);
or U4662 (N_4662,N_3429,N_3498);
nand U4663 (N_4663,N_3278,N_3528);
and U4664 (N_4664,N_3214,N_3564);
or U4665 (N_4665,N_3580,N_3899);
nand U4666 (N_4666,N_3982,N_3459);
nand U4667 (N_4667,N_3940,N_3377);
nor U4668 (N_4668,N_3597,N_3418);
or U4669 (N_4669,N_3093,N_3790);
nor U4670 (N_4670,N_3523,N_3218);
nand U4671 (N_4671,N_3069,N_3089);
nor U4672 (N_4672,N_3335,N_3696);
or U4673 (N_4673,N_3632,N_3496);
nor U4674 (N_4674,N_3027,N_3769);
or U4675 (N_4675,N_3253,N_3032);
nor U4676 (N_4676,N_3636,N_3676);
nand U4677 (N_4677,N_3666,N_3148);
or U4678 (N_4678,N_3997,N_3686);
nor U4679 (N_4679,N_3904,N_3882);
nor U4680 (N_4680,N_3630,N_3588);
or U4681 (N_4681,N_3382,N_3860);
or U4682 (N_4682,N_3520,N_3361);
or U4683 (N_4683,N_3713,N_3190);
or U4684 (N_4684,N_3684,N_3275);
and U4685 (N_4685,N_3043,N_3481);
or U4686 (N_4686,N_3313,N_3669);
nand U4687 (N_4687,N_3946,N_3375);
and U4688 (N_4688,N_3310,N_3440);
and U4689 (N_4689,N_3046,N_3734);
and U4690 (N_4690,N_3195,N_3660);
nor U4691 (N_4691,N_3426,N_3001);
nor U4692 (N_4692,N_3524,N_3018);
nor U4693 (N_4693,N_3979,N_3324);
nand U4694 (N_4694,N_3983,N_3297);
nor U4695 (N_4695,N_3017,N_3502);
nor U4696 (N_4696,N_3997,N_3328);
or U4697 (N_4697,N_3054,N_3540);
nor U4698 (N_4698,N_3295,N_3290);
nor U4699 (N_4699,N_3183,N_3688);
nand U4700 (N_4700,N_3690,N_3542);
and U4701 (N_4701,N_3325,N_3809);
nor U4702 (N_4702,N_3489,N_3366);
nand U4703 (N_4703,N_3319,N_3988);
nor U4704 (N_4704,N_3866,N_3073);
or U4705 (N_4705,N_3955,N_3392);
nand U4706 (N_4706,N_3846,N_3319);
nor U4707 (N_4707,N_3616,N_3019);
nor U4708 (N_4708,N_3134,N_3818);
or U4709 (N_4709,N_3504,N_3007);
or U4710 (N_4710,N_3495,N_3535);
nor U4711 (N_4711,N_3760,N_3069);
or U4712 (N_4712,N_3150,N_3142);
nand U4713 (N_4713,N_3025,N_3068);
nor U4714 (N_4714,N_3481,N_3064);
nor U4715 (N_4715,N_3957,N_3363);
and U4716 (N_4716,N_3459,N_3947);
nand U4717 (N_4717,N_3250,N_3383);
nor U4718 (N_4718,N_3597,N_3267);
and U4719 (N_4719,N_3889,N_3127);
or U4720 (N_4720,N_3865,N_3208);
nor U4721 (N_4721,N_3061,N_3908);
or U4722 (N_4722,N_3514,N_3016);
nand U4723 (N_4723,N_3593,N_3652);
nor U4724 (N_4724,N_3806,N_3314);
and U4725 (N_4725,N_3002,N_3005);
xnor U4726 (N_4726,N_3920,N_3432);
nand U4727 (N_4727,N_3688,N_3293);
or U4728 (N_4728,N_3705,N_3562);
or U4729 (N_4729,N_3265,N_3918);
nor U4730 (N_4730,N_3846,N_3595);
and U4731 (N_4731,N_3249,N_3850);
and U4732 (N_4732,N_3558,N_3903);
nor U4733 (N_4733,N_3401,N_3850);
nor U4734 (N_4734,N_3298,N_3803);
and U4735 (N_4735,N_3510,N_3728);
and U4736 (N_4736,N_3483,N_3157);
nor U4737 (N_4737,N_3521,N_3400);
nor U4738 (N_4738,N_3799,N_3742);
nand U4739 (N_4739,N_3158,N_3950);
or U4740 (N_4740,N_3429,N_3741);
and U4741 (N_4741,N_3417,N_3408);
or U4742 (N_4742,N_3910,N_3849);
and U4743 (N_4743,N_3921,N_3812);
or U4744 (N_4744,N_3985,N_3835);
nor U4745 (N_4745,N_3324,N_3546);
and U4746 (N_4746,N_3559,N_3150);
nand U4747 (N_4747,N_3121,N_3280);
and U4748 (N_4748,N_3712,N_3641);
nand U4749 (N_4749,N_3286,N_3820);
nor U4750 (N_4750,N_3876,N_3341);
or U4751 (N_4751,N_3508,N_3142);
or U4752 (N_4752,N_3874,N_3718);
nor U4753 (N_4753,N_3653,N_3774);
or U4754 (N_4754,N_3651,N_3042);
or U4755 (N_4755,N_3578,N_3412);
or U4756 (N_4756,N_3304,N_3188);
nor U4757 (N_4757,N_3803,N_3139);
or U4758 (N_4758,N_3935,N_3120);
and U4759 (N_4759,N_3519,N_3759);
nand U4760 (N_4760,N_3219,N_3184);
nand U4761 (N_4761,N_3119,N_3736);
nor U4762 (N_4762,N_3495,N_3481);
or U4763 (N_4763,N_3633,N_3452);
nor U4764 (N_4764,N_3018,N_3739);
and U4765 (N_4765,N_3451,N_3202);
and U4766 (N_4766,N_3156,N_3788);
xor U4767 (N_4767,N_3126,N_3083);
or U4768 (N_4768,N_3936,N_3988);
or U4769 (N_4769,N_3091,N_3705);
nand U4770 (N_4770,N_3976,N_3499);
and U4771 (N_4771,N_3396,N_3065);
or U4772 (N_4772,N_3994,N_3413);
nor U4773 (N_4773,N_3641,N_3815);
and U4774 (N_4774,N_3829,N_3288);
and U4775 (N_4775,N_3375,N_3941);
nor U4776 (N_4776,N_3960,N_3229);
and U4777 (N_4777,N_3694,N_3534);
and U4778 (N_4778,N_3097,N_3910);
nand U4779 (N_4779,N_3832,N_3270);
nor U4780 (N_4780,N_3538,N_3936);
nand U4781 (N_4781,N_3070,N_3675);
nor U4782 (N_4782,N_3318,N_3762);
or U4783 (N_4783,N_3802,N_3775);
or U4784 (N_4784,N_3903,N_3132);
nor U4785 (N_4785,N_3448,N_3513);
nor U4786 (N_4786,N_3880,N_3624);
nand U4787 (N_4787,N_3735,N_3985);
nand U4788 (N_4788,N_3506,N_3418);
nand U4789 (N_4789,N_3114,N_3481);
and U4790 (N_4790,N_3043,N_3341);
nor U4791 (N_4791,N_3395,N_3239);
and U4792 (N_4792,N_3165,N_3238);
or U4793 (N_4793,N_3159,N_3749);
nand U4794 (N_4794,N_3099,N_3961);
nor U4795 (N_4795,N_3479,N_3452);
or U4796 (N_4796,N_3153,N_3990);
nor U4797 (N_4797,N_3191,N_3459);
and U4798 (N_4798,N_3748,N_3692);
and U4799 (N_4799,N_3841,N_3507);
or U4800 (N_4800,N_3221,N_3373);
nand U4801 (N_4801,N_3216,N_3319);
and U4802 (N_4802,N_3003,N_3309);
nand U4803 (N_4803,N_3391,N_3179);
nor U4804 (N_4804,N_3776,N_3382);
or U4805 (N_4805,N_3465,N_3882);
nand U4806 (N_4806,N_3154,N_3226);
and U4807 (N_4807,N_3405,N_3258);
and U4808 (N_4808,N_3245,N_3886);
or U4809 (N_4809,N_3388,N_3065);
nand U4810 (N_4810,N_3347,N_3340);
and U4811 (N_4811,N_3710,N_3122);
or U4812 (N_4812,N_3417,N_3741);
nor U4813 (N_4813,N_3167,N_3499);
and U4814 (N_4814,N_3218,N_3221);
or U4815 (N_4815,N_3594,N_3018);
or U4816 (N_4816,N_3916,N_3010);
nor U4817 (N_4817,N_3722,N_3085);
nand U4818 (N_4818,N_3713,N_3465);
or U4819 (N_4819,N_3324,N_3770);
and U4820 (N_4820,N_3793,N_3263);
or U4821 (N_4821,N_3507,N_3314);
nor U4822 (N_4822,N_3475,N_3630);
nand U4823 (N_4823,N_3784,N_3470);
or U4824 (N_4824,N_3676,N_3398);
nor U4825 (N_4825,N_3036,N_3798);
nand U4826 (N_4826,N_3917,N_3028);
nand U4827 (N_4827,N_3312,N_3352);
nor U4828 (N_4828,N_3721,N_3474);
or U4829 (N_4829,N_3688,N_3938);
and U4830 (N_4830,N_3290,N_3659);
or U4831 (N_4831,N_3784,N_3799);
nand U4832 (N_4832,N_3005,N_3498);
nand U4833 (N_4833,N_3479,N_3321);
or U4834 (N_4834,N_3838,N_3875);
or U4835 (N_4835,N_3119,N_3609);
nor U4836 (N_4836,N_3986,N_3281);
and U4837 (N_4837,N_3326,N_3327);
or U4838 (N_4838,N_3227,N_3533);
and U4839 (N_4839,N_3481,N_3040);
nor U4840 (N_4840,N_3292,N_3072);
nand U4841 (N_4841,N_3311,N_3146);
nand U4842 (N_4842,N_3321,N_3419);
nand U4843 (N_4843,N_3163,N_3617);
nor U4844 (N_4844,N_3148,N_3870);
or U4845 (N_4845,N_3352,N_3456);
nor U4846 (N_4846,N_3104,N_3913);
nor U4847 (N_4847,N_3657,N_3403);
and U4848 (N_4848,N_3574,N_3989);
and U4849 (N_4849,N_3192,N_3103);
or U4850 (N_4850,N_3638,N_3663);
or U4851 (N_4851,N_3699,N_3905);
and U4852 (N_4852,N_3615,N_3225);
and U4853 (N_4853,N_3742,N_3267);
and U4854 (N_4854,N_3952,N_3093);
nor U4855 (N_4855,N_3048,N_3902);
or U4856 (N_4856,N_3751,N_3632);
or U4857 (N_4857,N_3401,N_3921);
nand U4858 (N_4858,N_3796,N_3789);
or U4859 (N_4859,N_3268,N_3081);
and U4860 (N_4860,N_3704,N_3810);
nand U4861 (N_4861,N_3834,N_3428);
and U4862 (N_4862,N_3650,N_3376);
and U4863 (N_4863,N_3882,N_3860);
nor U4864 (N_4864,N_3154,N_3358);
or U4865 (N_4865,N_3262,N_3318);
and U4866 (N_4866,N_3671,N_3199);
nand U4867 (N_4867,N_3905,N_3760);
nor U4868 (N_4868,N_3546,N_3665);
nor U4869 (N_4869,N_3573,N_3644);
nand U4870 (N_4870,N_3403,N_3306);
or U4871 (N_4871,N_3785,N_3079);
and U4872 (N_4872,N_3546,N_3399);
or U4873 (N_4873,N_3758,N_3591);
xnor U4874 (N_4874,N_3638,N_3775);
or U4875 (N_4875,N_3335,N_3030);
nor U4876 (N_4876,N_3288,N_3224);
nor U4877 (N_4877,N_3455,N_3365);
and U4878 (N_4878,N_3880,N_3031);
nand U4879 (N_4879,N_3620,N_3356);
nand U4880 (N_4880,N_3039,N_3502);
nor U4881 (N_4881,N_3530,N_3518);
and U4882 (N_4882,N_3050,N_3904);
or U4883 (N_4883,N_3685,N_3709);
nand U4884 (N_4884,N_3236,N_3878);
and U4885 (N_4885,N_3867,N_3265);
and U4886 (N_4886,N_3901,N_3265);
and U4887 (N_4887,N_3704,N_3734);
or U4888 (N_4888,N_3748,N_3238);
and U4889 (N_4889,N_3187,N_3862);
and U4890 (N_4890,N_3600,N_3944);
nor U4891 (N_4891,N_3662,N_3087);
nand U4892 (N_4892,N_3399,N_3968);
nand U4893 (N_4893,N_3496,N_3916);
nand U4894 (N_4894,N_3014,N_3483);
nand U4895 (N_4895,N_3540,N_3355);
xnor U4896 (N_4896,N_3849,N_3785);
nor U4897 (N_4897,N_3582,N_3759);
or U4898 (N_4898,N_3144,N_3257);
nor U4899 (N_4899,N_3829,N_3022);
or U4900 (N_4900,N_3385,N_3005);
or U4901 (N_4901,N_3861,N_3947);
nand U4902 (N_4902,N_3658,N_3622);
and U4903 (N_4903,N_3982,N_3120);
or U4904 (N_4904,N_3456,N_3939);
xnor U4905 (N_4905,N_3468,N_3715);
nand U4906 (N_4906,N_3569,N_3087);
and U4907 (N_4907,N_3884,N_3359);
or U4908 (N_4908,N_3093,N_3784);
nand U4909 (N_4909,N_3939,N_3113);
or U4910 (N_4910,N_3812,N_3742);
or U4911 (N_4911,N_3706,N_3593);
nand U4912 (N_4912,N_3225,N_3605);
or U4913 (N_4913,N_3557,N_3413);
nand U4914 (N_4914,N_3790,N_3425);
and U4915 (N_4915,N_3370,N_3455);
nand U4916 (N_4916,N_3217,N_3759);
and U4917 (N_4917,N_3496,N_3643);
or U4918 (N_4918,N_3963,N_3379);
nor U4919 (N_4919,N_3849,N_3851);
nor U4920 (N_4920,N_3485,N_3051);
nor U4921 (N_4921,N_3926,N_3031);
nor U4922 (N_4922,N_3059,N_3490);
xor U4923 (N_4923,N_3887,N_3060);
nor U4924 (N_4924,N_3929,N_3294);
and U4925 (N_4925,N_3683,N_3702);
nand U4926 (N_4926,N_3956,N_3356);
and U4927 (N_4927,N_3006,N_3360);
and U4928 (N_4928,N_3423,N_3370);
or U4929 (N_4929,N_3368,N_3269);
nor U4930 (N_4930,N_3611,N_3155);
and U4931 (N_4931,N_3317,N_3247);
or U4932 (N_4932,N_3724,N_3852);
or U4933 (N_4933,N_3228,N_3766);
nand U4934 (N_4934,N_3598,N_3939);
and U4935 (N_4935,N_3427,N_3931);
nor U4936 (N_4936,N_3096,N_3921);
nor U4937 (N_4937,N_3495,N_3797);
and U4938 (N_4938,N_3039,N_3513);
nor U4939 (N_4939,N_3368,N_3516);
nand U4940 (N_4940,N_3976,N_3221);
nor U4941 (N_4941,N_3710,N_3949);
nand U4942 (N_4942,N_3672,N_3976);
nor U4943 (N_4943,N_3932,N_3977);
or U4944 (N_4944,N_3378,N_3873);
or U4945 (N_4945,N_3343,N_3173);
or U4946 (N_4946,N_3271,N_3373);
and U4947 (N_4947,N_3500,N_3796);
nand U4948 (N_4948,N_3314,N_3297);
nor U4949 (N_4949,N_3513,N_3223);
nor U4950 (N_4950,N_3624,N_3053);
nor U4951 (N_4951,N_3817,N_3515);
and U4952 (N_4952,N_3505,N_3604);
and U4953 (N_4953,N_3694,N_3938);
or U4954 (N_4954,N_3356,N_3768);
or U4955 (N_4955,N_3492,N_3201);
nand U4956 (N_4956,N_3920,N_3670);
or U4957 (N_4957,N_3539,N_3867);
or U4958 (N_4958,N_3959,N_3483);
nor U4959 (N_4959,N_3308,N_3091);
nand U4960 (N_4960,N_3922,N_3256);
nor U4961 (N_4961,N_3444,N_3762);
nand U4962 (N_4962,N_3463,N_3867);
nor U4963 (N_4963,N_3427,N_3542);
and U4964 (N_4964,N_3367,N_3283);
nor U4965 (N_4965,N_3715,N_3900);
or U4966 (N_4966,N_3706,N_3883);
and U4967 (N_4967,N_3758,N_3085);
nor U4968 (N_4968,N_3267,N_3457);
and U4969 (N_4969,N_3507,N_3668);
and U4970 (N_4970,N_3388,N_3347);
nor U4971 (N_4971,N_3918,N_3706);
and U4972 (N_4972,N_3013,N_3749);
and U4973 (N_4973,N_3571,N_3874);
nor U4974 (N_4974,N_3237,N_3935);
and U4975 (N_4975,N_3925,N_3965);
nand U4976 (N_4976,N_3939,N_3269);
nor U4977 (N_4977,N_3551,N_3917);
or U4978 (N_4978,N_3305,N_3273);
or U4979 (N_4979,N_3326,N_3384);
nand U4980 (N_4980,N_3597,N_3864);
nor U4981 (N_4981,N_3217,N_3383);
nor U4982 (N_4982,N_3226,N_3070);
nand U4983 (N_4983,N_3028,N_3947);
and U4984 (N_4984,N_3640,N_3132);
or U4985 (N_4985,N_3827,N_3973);
nand U4986 (N_4986,N_3093,N_3257);
and U4987 (N_4987,N_3782,N_3499);
and U4988 (N_4988,N_3961,N_3537);
nor U4989 (N_4989,N_3045,N_3082);
and U4990 (N_4990,N_3293,N_3812);
nand U4991 (N_4991,N_3043,N_3463);
or U4992 (N_4992,N_3129,N_3494);
and U4993 (N_4993,N_3150,N_3963);
and U4994 (N_4994,N_3346,N_3018);
or U4995 (N_4995,N_3254,N_3722);
and U4996 (N_4996,N_3755,N_3178);
or U4997 (N_4997,N_3233,N_3150);
or U4998 (N_4998,N_3718,N_3263);
nand U4999 (N_4999,N_3156,N_3589);
nand U5000 (N_5000,N_4780,N_4709);
and U5001 (N_5001,N_4050,N_4524);
xor U5002 (N_5002,N_4778,N_4249);
nand U5003 (N_5003,N_4988,N_4942);
nand U5004 (N_5004,N_4868,N_4782);
nand U5005 (N_5005,N_4769,N_4454);
nor U5006 (N_5006,N_4033,N_4626);
or U5007 (N_5007,N_4911,N_4895);
and U5008 (N_5008,N_4802,N_4196);
nand U5009 (N_5009,N_4761,N_4822);
nand U5010 (N_5010,N_4189,N_4439);
and U5011 (N_5011,N_4979,N_4512);
and U5012 (N_5012,N_4443,N_4351);
or U5013 (N_5013,N_4920,N_4426);
nand U5014 (N_5014,N_4501,N_4046);
xor U5015 (N_5015,N_4362,N_4131);
nor U5016 (N_5016,N_4392,N_4264);
nor U5017 (N_5017,N_4531,N_4469);
nor U5018 (N_5018,N_4041,N_4358);
or U5019 (N_5019,N_4089,N_4651);
nand U5020 (N_5020,N_4913,N_4420);
and U5021 (N_5021,N_4019,N_4954);
nand U5022 (N_5022,N_4768,N_4779);
or U5023 (N_5023,N_4659,N_4929);
nand U5024 (N_5024,N_4687,N_4560);
or U5025 (N_5025,N_4835,N_4969);
nor U5026 (N_5026,N_4744,N_4243);
and U5027 (N_5027,N_4676,N_4239);
nand U5028 (N_5028,N_4902,N_4923);
nand U5029 (N_5029,N_4149,N_4349);
and U5030 (N_5030,N_4061,N_4649);
nor U5031 (N_5031,N_4409,N_4506);
xor U5032 (N_5032,N_4135,N_4887);
or U5033 (N_5033,N_4881,N_4217);
or U5034 (N_5034,N_4719,N_4322);
or U5035 (N_5035,N_4573,N_4009);
nand U5036 (N_5036,N_4773,N_4260);
nand U5037 (N_5037,N_4021,N_4825);
nor U5038 (N_5038,N_4927,N_4488);
nand U5039 (N_5039,N_4419,N_4701);
nand U5040 (N_5040,N_4346,N_4974);
nor U5041 (N_5041,N_4291,N_4675);
or U5042 (N_5042,N_4532,N_4357);
nand U5043 (N_5043,N_4637,N_4574);
nand U5044 (N_5044,N_4998,N_4111);
nor U5045 (N_5045,N_4638,N_4229);
nor U5046 (N_5046,N_4630,N_4422);
and U5047 (N_5047,N_4334,N_4765);
and U5048 (N_5048,N_4302,N_4284);
nor U5049 (N_5049,N_4300,N_4254);
xor U5050 (N_5050,N_4916,N_4003);
nor U5051 (N_5051,N_4533,N_4490);
nand U5052 (N_5052,N_4672,N_4017);
or U5053 (N_5053,N_4953,N_4310);
nand U5054 (N_5054,N_4604,N_4746);
or U5055 (N_5055,N_4461,N_4048);
or U5056 (N_5056,N_4318,N_4722);
nand U5057 (N_5057,N_4278,N_4222);
nand U5058 (N_5058,N_4355,N_4184);
or U5059 (N_5059,N_4363,N_4801);
nor U5060 (N_5060,N_4192,N_4495);
or U5061 (N_5061,N_4014,N_4126);
and U5062 (N_5062,N_4353,N_4809);
nand U5063 (N_5063,N_4097,N_4319);
and U5064 (N_5064,N_4085,N_4516);
or U5065 (N_5065,N_4551,N_4095);
nand U5066 (N_5066,N_4082,N_4981);
or U5067 (N_5067,N_4669,N_4772);
and U5068 (N_5068,N_4452,N_4839);
nand U5069 (N_5069,N_4579,N_4416);
nand U5070 (N_5070,N_4288,N_4663);
nor U5071 (N_5071,N_4083,N_4108);
and U5072 (N_5072,N_4486,N_4550);
and U5073 (N_5073,N_4038,N_4614);
and U5074 (N_5074,N_4618,N_4889);
nand U5075 (N_5075,N_4647,N_4892);
nand U5076 (N_5076,N_4955,N_4536);
nand U5077 (N_5077,N_4143,N_4205);
and U5078 (N_5078,N_4695,N_4186);
and U5079 (N_5079,N_4323,N_4157);
and U5080 (N_5080,N_4390,N_4577);
and U5081 (N_5081,N_4811,N_4987);
nand U5082 (N_5082,N_4151,N_4689);
or U5083 (N_5083,N_4933,N_4924);
nor U5084 (N_5084,N_4241,N_4863);
nor U5085 (N_5085,N_4406,N_4044);
nor U5086 (N_5086,N_4795,N_4330);
nor U5087 (N_5087,N_4563,N_4633);
nand U5088 (N_5088,N_4738,N_4487);
or U5089 (N_5089,N_4166,N_4005);
nand U5090 (N_5090,N_4571,N_4505);
or U5091 (N_5091,N_4843,N_4263);
and U5092 (N_5092,N_4088,N_4712);
or U5093 (N_5093,N_4656,N_4567);
or U5094 (N_5094,N_4584,N_4645);
nand U5095 (N_5095,N_4666,N_4527);
and U5096 (N_5096,N_4716,N_4748);
nand U5097 (N_5097,N_4446,N_4627);
nand U5098 (N_5098,N_4803,N_4921);
xor U5099 (N_5099,N_4429,N_4326);
or U5100 (N_5100,N_4673,N_4432);
nor U5101 (N_5101,N_4824,N_4960);
nor U5102 (N_5102,N_4437,N_4128);
and U5103 (N_5103,N_4220,N_4417);
nor U5104 (N_5104,N_4029,N_4674);
or U5105 (N_5105,N_4086,N_4664);
and U5106 (N_5106,N_4093,N_4818);
nand U5107 (N_5107,N_4070,N_4671);
or U5108 (N_5108,N_4631,N_4256);
nand U5109 (N_5109,N_4472,N_4226);
nor U5110 (N_5110,N_4950,N_4413);
and U5111 (N_5111,N_4228,N_4043);
xnor U5112 (N_5112,N_4606,N_4332);
nor U5113 (N_5113,N_4344,N_4366);
and U5114 (N_5114,N_4207,N_4183);
and U5115 (N_5115,N_4667,N_4977);
or U5116 (N_5116,N_4290,N_4855);
nand U5117 (N_5117,N_4042,N_4542);
or U5118 (N_5118,N_4588,N_4138);
and U5119 (N_5119,N_4583,N_4371);
nand U5120 (N_5120,N_4150,N_4745);
xnor U5121 (N_5121,N_4838,N_4657);
or U5122 (N_5122,N_4990,N_4342);
nand U5123 (N_5123,N_4211,N_4703);
nor U5124 (N_5124,N_4098,N_4543);
nand U5125 (N_5125,N_4939,N_4653);
or U5126 (N_5126,N_4575,N_4327);
or U5127 (N_5127,N_4770,N_4849);
and U5128 (N_5128,N_4023,N_4844);
nor U5129 (N_5129,N_4841,N_4224);
or U5130 (N_5130,N_4137,N_4576);
nand U5131 (N_5131,N_4236,N_4870);
nor U5132 (N_5132,N_4293,N_4530);
nand U5133 (N_5133,N_4002,N_4741);
and U5134 (N_5134,N_4521,N_4539);
nor U5135 (N_5135,N_4265,N_4785);
nand U5136 (N_5136,N_4368,N_4589);
nand U5137 (N_5137,N_4733,N_4523);
and U5138 (N_5138,N_4548,N_4142);
or U5139 (N_5139,N_4750,N_4297);
nand U5140 (N_5140,N_4430,N_4641);
or U5141 (N_5141,N_4018,N_4391);
nor U5142 (N_5142,N_4154,N_4118);
and U5143 (N_5143,N_4752,N_4888);
nand U5144 (N_5144,N_4103,N_4175);
and U5145 (N_5145,N_4807,N_4587);
and U5146 (N_5146,N_4713,N_4360);
and U5147 (N_5147,N_4985,N_4001);
nand U5148 (N_5148,N_4743,N_4075);
nor U5149 (N_5149,N_4427,N_4514);
or U5150 (N_5150,N_4938,N_4590);
or U5151 (N_5151,N_4312,N_4145);
or U5152 (N_5152,N_4296,N_4854);
and U5153 (N_5153,N_4796,N_4279);
nand U5154 (N_5154,N_4528,N_4833);
and U5155 (N_5155,N_4845,N_4066);
or U5156 (N_5156,N_4295,N_4515);
nand U5157 (N_5157,N_4139,N_4130);
nor U5158 (N_5158,N_4156,N_4476);
and U5159 (N_5159,N_4110,N_4946);
nor U5160 (N_5160,N_4966,N_4678);
nor U5161 (N_5161,N_4181,N_4388);
nand U5162 (N_5162,N_4073,N_4337);
or U5163 (N_5163,N_4777,N_4707);
nand U5164 (N_5164,N_4629,N_4679);
or U5165 (N_5165,N_4037,N_4850);
and U5166 (N_5166,N_4068,N_4596);
and U5167 (N_5167,N_4307,N_4899);
nor U5168 (N_5168,N_4072,N_4943);
nor U5169 (N_5169,N_4176,N_4737);
nor U5170 (N_5170,N_4553,N_4306);
and U5171 (N_5171,N_4136,N_4159);
nor U5172 (N_5172,N_4727,N_4755);
or U5173 (N_5173,N_4791,N_4798);
and U5174 (N_5174,N_4564,N_4127);
and U5175 (N_5175,N_4754,N_4435);
or U5176 (N_5176,N_4853,N_4878);
and U5177 (N_5177,N_4901,N_4994);
nand U5178 (N_5178,N_4153,N_4930);
or U5179 (N_5179,N_4370,N_4753);
nand U5180 (N_5180,N_4786,N_4873);
and U5181 (N_5181,N_4794,N_4393);
or U5182 (N_5182,N_4039,N_4094);
nand U5183 (N_5183,N_4340,N_4812);
or U5184 (N_5184,N_4418,N_4065);
nand U5185 (N_5185,N_4174,N_4040);
and U5186 (N_5186,N_4456,N_4080);
nor U5187 (N_5187,N_4078,N_4747);
nor U5188 (N_5188,N_4926,N_4210);
nand U5189 (N_5189,N_4504,N_4815);
nor U5190 (N_5190,N_4261,N_4190);
and U5191 (N_5191,N_4721,N_4771);
or U5192 (N_5192,N_4117,N_4757);
nand U5193 (N_5193,N_4864,N_4968);
nor U5194 (N_5194,N_4762,N_4509);
nand U5195 (N_5195,N_4299,N_4125);
or U5196 (N_5196,N_4062,N_4272);
or U5197 (N_5197,N_4467,N_4394);
or U5198 (N_5198,N_4329,N_4036);
nor U5199 (N_5199,N_4244,N_4789);
nand U5200 (N_5200,N_4975,N_4114);
nor U5201 (N_5201,N_4891,N_4980);
nand U5202 (N_5202,N_4706,N_4012);
nand U5203 (N_5203,N_4423,N_4221);
or U5204 (N_5204,N_4644,N_4875);
and U5205 (N_5205,N_4623,N_4556);
nand U5206 (N_5206,N_4376,N_4354);
or U5207 (N_5207,N_4882,N_4661);
nand U5208 (N_5208,N_4378,N_4460);
and U5209 (N_5209,N_4711,N_4121);
and U5210 (N_5210,N_4739,N_4298);
nand U5211 (N_5211,N_4045,N_4397);
or U5212 (N_5212,N_4714,N_4544);
nand U5213 (N_5213,N_4011,N_4986);
or U5214 (N_5214,N_4652,N_4250);
or U5215 (N_5215,N_4113,N_4890);
and U5216 (N_5216,N_4705,N_4897);
nand U5217 (N_5217,N_4381,N_4999);
nand U5218 (N_5218,N_4235,N_4022);
nor U5219 (N_5219,N_4615,N_4101);
nand U5220 (N_5220,N_4962,N_4328);
nand U5221 (N_5221,N_4335,N_4790);
nand U5222 (N_5222,N_4425,N_4496);
or U5223 (N_5223,N_4559,N_4925);
nor U5224 (N_5224,N_4144,N_4814);
or U5225 (N_5225,N_4494,N_4348);
or U5226 (N_5226,N_4106,N_4102);
and U5227 (N_5227,N_4374,N_4997);
nand U5228 (N_5228,N_4379,N_4160);
or U5229 (N_5229,N_4280,N_4438);
nand U5230 (N_5230,N_4493,N_4594);
and U5231 (N_5231,N_4453,N_4421);
or U5232 (N_5232,N_4808,N_4350);
and U5233 (N_5233,N_4941,N_4252);
and U5234 (N_5234,N_4030,N_4026);
nor U5235 (N_5235,N_4459,N_4133);
nor U5236 (N_5236,N_4386,N_4313);
or U5237 (N_5237,N_4625,N_4917);
or U5238 (N_5238,N_4225,N_4991);
nor U5239 (N_5239,N_4598,N_4027);
or U5240 (N_5240,N_4134,N_4107);
nor U5241 (N_5241,N_4016,N_4325);
and U5242 (N_5242,N_4315,N_4451);
xnor U5243 (N_5243,N_4465,N_4591);
nor U5244 (N_5244,N_4056,N_4281);
or U5245 (N_5245,N_4170,N_4862);
and U5246 (N_5246,N_4908,N_4586);
nand U5247 (N_5247,N_4874,N_4468);
xor U5248 (N_5248,N_4540,N_4356);
and U5249 (N_5249,N_4555,N_4398);
nand U5250 (N_5250,N_4499,N_4407);
nand U5251 (N_5251,N_4665,N_4728);
and U5252 (N_5252,N_4508,N_4526);
nor U5253 (N_5253,N_4013,N_4823);
nand U5254 (N_5254,N_4502,N_4436);
nand U5255 (N_5255,N_4879,N_4377);
nor U5256 (N_5256,N_4147,N_4247);
nand U5257 (N_5257,N_4694,N_4231);
xnor U5258 (N_5258,N_4763,N_4783);
nand U5259 (N_5259,N_4820,N_4047);
and U5260 (N_5260,N_4698,N_4015);
or U5261 (N_5261,N_4266,N_4064);
nor U5262 (N_5262,N_4304,N_4333);
nor U5263 (N_5263,N_4457,N_4240);
xnor U5264 (N_5264,N_4865,N_4268);
and U5265 (N_5265,N_4475,N_4905);
or U5266 (N_5266,N_4466,N_4740);
nand U5267 (N_5267,N_4970,N_4336);
nor U5268 (N_5268,N_4074,N_4720);
and U5269 (N_5269,N_4058,N_4491);
or U5270 (N_5270,N_4119,N_4518);
nand U5271 (N_5271,N_4682,N_4431);
nand U5272 (N_5272,N_4028,N_4819);
and U5273 (N_5273,N_4402,N_4316);
nand U5274 (N_5274,N_4934,N_4828);
xnor U5275 (N_5275,N_4301,N_4681);
nand U5276 (N_5276,N_4936,N_4214);
nor U5277 (N_5277,N_4766,N_4867);
or U5278 (N_5278,N_4602,N_4163);
or U5279 (N_5279,N_4995,N_4520);
nor U5280 (N_5280,N_4758,N_4498);
nand U5281 (N_5281,N_4624,N_4906);
nor U5282 (N_5282,N_4294,N_4096);
or U5283 (N_5283,N_4219,N_4578);
and U5284 (N_5284,N_4052,N_4091);
and U5285 (N_5285,N_4636,N_4537);
or U5286 (N_5286,N_4580,N_4051);
nor U5287 (N_5287,N_4730,N_4872);
or U5288 (N_5288,N_4285,N_4158);
nor U5289 (N_5289,N_4399,N_4683);
or U5290 (N_5290,N_4725,N_4948);
nand U5291 (N_5291,N_4635,N_4433);
nor U5292 (N_5292,N_4230,N_4200);
and U5293 (N_5293,N_4617,N_4063);
nand U5294 (N_5294,N_4759,N_4479);
or U5295 (N_5295,N_4582,N_4640);
nand U5296 (N_5296,N_4947,N_4538);
nand U5297 (N_5297,N_4726,N_4704);
or U5298 (N_5298,N_4736,N_4919);
and U5299 (N_5299,N_4463,N_4481);
nor U5300 (N_5300,N_4203,N_4206);
or U5301 (N_5301,N_4100,N_4507);
and U5302 (N_5302,N_4610,N_4477);
or U5303 (N_5303,N_4834,N_4984);
nand U5304 (N_5304,N_4165,N_4444);
nand U5305 (N_5305,N_4049,N_4982);
nand U5306 (N_5306,N_4836,N_4710);
or U5307 (N_5307,N_4896,N_4218);
or U5308 (N_5308,N_4359,N_4367);
and U5309 (N_5309,N_4480,N_4961);
and U5310 (N_5310,N_4233,N_4621);
or U5311 (N_5311,N_4731,N_4776);
or U5312 (N_5312,N_4059,N_4613);
nand U5313 (N_5313,N_4851,N_4006);
or U5314 (N_5314,N_4688,N_4167);
and U5315 (N_5315,N_4213,N_4522);
or U5316 (N_5316,N_4568,N_4104);
and U5317 (N_5317,N_4020,N_4848);
xor U5318 (N_5318,N_4470,N_4842);
nand U5319 (N_5319,N_4648,N_4952);
nand U5320 (N_5320,N_4384,N_4311);
and U5321 (N_5321,N_4866,N_4338);
nand U5322 (N_5322,N_4308,N_4549);
nor U5323 (N_5323,N_4497,N_4248);
or U5324 (N_5324,N_4109,N_4566);
or U5325 (N_5325,N_4650,N_4403);
nor U5326 (N_5326,N_4025,N_4081);
nor U5327 (N_5327,N_4788,N_4963);
nand U5328 (N_5328,N_4662,N_4259);
nand U5329 (N_5329,N_4519,N_4034);
nand U5330 (N_5330,N_4199,N_4309);
or U5331 (N_5331,N_4529,N_4632);
nand U5332 (N_5332,N_4171,N_4369);
and U5333 (N_5333,N_4935,N_4320);
and U5334 (N_5334,N_4283,N_4169);
nand U5335 (N_5335,N_4116,N_4185);
or U5336 (N_5336,N_4352,N_4816);
and U5337 (N_5337,N_4639,N_4373);
nand U5338 (N_5338,N_4215,N_4900);
or U5339 (N_5339,N_4484,N_4668);
nor U5340 (N_5340,N_4305,N_4057);
nand U5341 (N_5341,N_4742,N_4907);
nand U5342 (N_5342,N_4365,N_4105);
nand U5343 (N_5343,N_4691,N_4408);
or U5344 (N_5344,N_4274,N_4751);
or U5345 (N_5345,N_4071,N_4992);
and U5346 (N_5346,N_4869,N_4122);
or U5347 (N_5347,N_4646,N_4194);
and U5348 (N_5348,N_4445,N_4172);
nand U5349 (N_5349,N_4428,N_4784);
xnor U5350 (N_5350,N_4546,N_4148);
nand U5351 (N_5351,N_4871,N_4565);
nand U5352 (N_5352,N_4204,N_4561);
nand U5353 (N_5353,N_4455,N_4547);
nor U5354 (N_5354,N_4655,N_4570);
or U5355 (N_5355,N_4774,N_4599);
and U5356 (N_5356,N_4702,N_4084);
nand U5357 (N_5357,N_4967,N_4182);
nor U5358 (N_5358,N_4880,N_4846);
or U5359 (N_5359,N_4931,N_4004);
nor U5360 (N_5360,N_4282,N_4152);
xnor U5361 (N_5361,N_4483,N_4735);
nand U5362 (N_5362,N_4690,N_4608);
or U5363 (N_5363,N_4609,N_4343);
or U5364 (N_5364,N_4956,N_4799);
and U5365 (N_5365,N_4164,N_4600);
and U5366 (N_5366,N_4054,N_4077);
or U5367 (N_5367,N_4861,N_4729);
or U5368 (N_5368,N_4092,N_4115);
nand U5369 (N_5369,N_4775,N_4922);
nor U5370 (N_5370,N_4797,N_4595);
nand U5371 (N_5371,N_4462,N_4654);
and U5372 (N_5372,N_4303,N_4603);
nand U5373 (N_5373,N_4400,N_4840);
and U5374 (N_5374,N_4383,N_4535);
or U5375 (N_5375,N_4976,N_4940);
nor U5376 (N_5376,N_4918,N_4253);
nor U5377 (N_5377,N_4271,N_4411);
nor U5378 (N_5378,N_4187,N_4670);
nand U5379 (N_5379,N_4723,N_4197);
and U5380 (N_5380,N_4267,N_4904);
nor U5381 (N_5381,N_4345,N_4611);
nor U5382 (N_5382,N_4964,N_4767);
and U5383 (N_5383,N_4972,N_4511);
nor U5384 (N_5384,N_4517,N_4804);
or U5385 (N_5385,N_4464,N_4162);
or U5386 (N_5386,N_4557,N_4837);
and U5387 (N_5387,N_4489,N_4658);
or U5388 (N_5388,N_4257,N_4831);
nand U5389 (N_5389,N_4697,N_4593);
or U5390 (N_5390,N_4852,N_4572);
and U5391 (N_5391,N_4717,N_4692);
or U5392 (N_5392,N_4718,N_4525);
xor U5393 (N_5393,N_4958,N_4513);
nor U5394 (N_5394,N_4592,N_4277);
and U5395 (N_5395,N_4680,N_4826);
or U5396 (N_5396,N_4321,N_4292);
and U5397 (N_5397,N_4860,N_4492);
nand U5398 (N_5398,N_4474,N_4545);
nor U5399 (N_5399,N_4700,N_4434);
nor U5400 (N_5400,N_4450,N_4605);
and U5401 (N_5401,N_4541,N_4937);
nor U5402 (N_5402,N_4732,N_4251);
and U5403 (N_5403,N_4708,N_4275);
or U5404 (N_5404,N_4877,N_4234);
nor U5405 (N_5405,N_4957,N_4202);
nor U5406 (N_5406,N_4188,N_4415);
nand U5407 (N_5407,N_4724,N_4031);
nor U5408 (N_5408,N_4010,N_4597);
and U5409 (N_5409,N_4120,N_4781);
and U5410 (N_5410,N_4983,N_4227);
nand U5411 (N_5411,N_4569,N_4060);
or U5412 (N_5412,N_4696,N_4485);
nor U5413 (N_5413,N_4686,N_4414);
or U5414 (N_5414,N_4500,N_4859);
nand U5415 (N_5415,N_4827,N_4339);
or U5416 (N_5416,N_4405,N_4684);
nand U5417 (N_5417,N_4699,N_4076);
nor U5418 (N_5418,N_4959,N_4317);
nor U5419 (N_5419,N_4255,N_4915);
nand U5420 (N_5420,N_4364,N_4734);
and U5421 (N_5421,N_4912,N_4032);
or U5422 (N_5422,N_4643,N_4884);
and U5423 (N_5423,N_4458,N_4314);
nand U5424 (N_5424,N_4375,N_4246);
nor U5425 (N_5425,N_4619,N_4404);
xnor U5426 (N_5426,N_4806,N_4178);
nand U5427 (N_5427,N_4140,N_4971);
or U5428 (N_5428,N_4155,N_4909);
or U5429 (N_5429,N_4829,N_4885);
nand U5430 (N_5430,N_4069,N_4287);
and U5431 (N_5431,N_4132,N_4989);
or U5432 (N_5432,N_4607,N_4024);
or U5433 (N_5433,N_4331,N_4223);
nor U5434 (N_5434,N_4847,N_4389);
nor U5435 (N_5435,N_4764,N_4787);
or U5436 (N_5436,N_4800,N_4198);
or U5437 (N_5437,N_4601,N_4914);
nand U5438 (N_5438,N_4793,N_4558);
nand U5439 (N_5439,N_4035,N_4622);
nand U5440 (N_5440,N_4996,N_4396);
and U5441 (N_5441,N_4146,N_4441);
nand U5442 (N_5442,N_4616,N_4099);
or U5443 (N_5443,N_4173,N_4289);
nor U5444 (N_5444,N_4554,N_4760);
nor U5445 (N_5445,N_4201,N_4876);
xnor U5446 (N_5446,N_4993,N_4324);
or U5447 (N_5447,N_4447,N_4628);
or U5448 (N_5448,N_4893,N_4269);
nand U5449 (N_5449,N_4478,N_4382);
or U5450 (N_5450,N_4112,N_4424);
or U5451 (N_5451,N_4124,N_4756);
and U5452 (N_5452,N_4749,N_4195);
nand U5453 (N_5453,N_4237,N_4471);
or U5454 (N_5454,N_4448,N_4715);
or U5455 (N_5455,N_4238,N_4642);
or U5456 (N_5456,N_4886,N_4007);
or U5457 (N_5457,N_4341,N_4067);
nor U5458 (N_5458,N_4090,N_4932);
and U5459 (N_5459,N_4191,N_4161);
nand U5460 (N_5460,N_4832,N_4562);
or U5461 (N_5461,N_4830,N_4581);
nand U5462 (N_5462,N_4440,N_4612);
nor U5463 (N_5463,N_4087,N_4928);
and U5464 (N_5464,N_4817,N_4180);
or U5465 (N_5465,N_4973,N_4473);
or U5466 (N_5466,N_4380,N_4693);
nor U5467 (N_5467,N_4401,N_4810);
and U5468 (N_5468,N_4945,N_4193);
and U5469 (N_5469,N_4805,N_4168);
or U5470 (N_5470,N_4552,N_4898);
nor U5471 (N_5471,N_4858,N_4055);
and U5472 (N_5472,N_4449,N_4442);
nor U5473 (N_5473,N_4209,N_4245);
and U5474 (N_5474,N_4258,N_4482);
or U5475 (N_5475,N_4179,N_4372);
nor U5476 (N_5476,N_4262,N_4008);
or U5477 (N_5477,N_4141,N_4242);
or U5478 (N_5478,N_4270,N_4903);
and U5479 (N_5479,N_4129,N_4177);
or U5480 (N_5480,N_4660,N_4232);
nor U5481 (N_5481,N_4620,N_4978);
and U5482 (N_5482,N_4079,N_4894);
nor U5483 (N_5483,N_4216,N_4412);
or U5484 (N_5484,N_4000,N_4910);
or U5485 (N_5485,N_4212,N_4385);
nor U5486 (N_5486,N_4634,N_4510);
nor U5487 (N_5487,N_4286,N_4387);
nand U5488 (N_5488,N_4347,N_4410);
or U5489 (N_5489,N_4856,N_4685);
nand U5490 (N_5490,N_4273,N_4949);
or U5491 (N_5491,N_4208,N_4944);
and U5492 (N_5492,N_4857,N_4677);
nand U5493 (N_5493,N_4821,N_4503);
nor U5494 (N_5494,N_4792,N_4585);
nor U5495 (N_5495,N_4395,N_4813);
nand U5496 (N_5496,N_4965,N_4053);
nor U5497 (N_5497,N_4123,N_4951);
nor U5498 (N_5498,N_4534,N_4276);
and U5499 (N_5499,N_4883,N_4361);
nand U5500 (N_5500,N_4947,N_4079);
and U5501 (N_5501,N_4116,N_4156);
and U5502 (N_5502,N_4752,N_4247);
and U5503 (N_5503,N_4832,N_4544);
nand U5504 (N_5504,N_4446,N_4335);
nand U5505 (N_5505,N_4692,N_4118);
and U5506 (N_5506,N_4503,N_4522);
nor U5507 (N_5507,N_4183,N_4767);
and U5508 (N_5508,N_4066,N_4317);
and U5509 (N_5509,N_4667,N_4682);
or U5510 (N_5510,N_4470,N_4688);
nand U5511 (N_5511,N_4789,N_4700);
and U5512 (N_5512,N_4994,N_4973);
or U5513 (N_5513,N_4275,N_4441);
nor U5514 (N_5514,N_4453,N_4130);
or U5515 (N_5515,N_4817,N_4179);
or U5516 (N_5516,N_4428,N_4225);
nor U5517 (N_5517,N_4265,N_4542);
or U5518 (N_5518,N_4108,N_4324);
nand U5519 (N_5519,N_4091,N_4928);
and U5520 (N_5520,N_4618,N_4229);
or U5521 (N_5521,N_4957,N_4699);
or U5522 (N_5522,N_4923,N_4619);
nand U5523 (N_5523,N_4232,N_4079);
and U5524 (N_5524,N_4138,N_4633);
nand U5525 (N_5525,N_4475,N_4855);
nand U5526 (N_5526,N_4859,N_4040);
nand U5527 (N_5527,N_4632,N_4920);
nor U5528 (N_5528,N_4783,N_4498);
xnor U5529 (N_5529,N_4806,N_4796);
nor U5530 (N_5530,N_4180,N_4905);
nor U5531 (N_5531,N_4873,N_4980);
xnor U5532 (N_5532,N_4347,N_4476);
and U5533 (N_5533,N_4013,N_4147);
or U5534 (N_5534,N_4168,N_4456);
and U5535 (N_5535,N_4833,N_4824);
nor U5536 (N_5536,N_4383,N_4564);
and U5537 (N_5537,N_4580,N_4120);
or U5538 (N_5538,N_4972,N_4929);
xor U5539 (N_5539,N_4521,N_4631);
or U5540 (N_5540,N_4989,N_4054);
nand U5541 (N_5541,N_4599,N_4466);
nor U5542 (N_5542,N_4953,N_4815);
xor U5543 (N_5543,N_4704,N_4149);
nor U5544 (N_5544,N_4238,N_4499);
and U5545 (N_5545,N_4831,N_4541);
nand U5546 (N_5546,N_4013,N_4979);
or U5547 (N_5547,N_4359,N_4252);
or U5548 (N_5548,N_4641,N_4363);
nand U5549 (N_5549,N_4583,N_4159);
or U5550 (N_5550,N_4127,N_4940);
or U5551 (N_5551,N_4052,N_4511);
and U5552 (N_5552,N_4020,N_4941);
xnor U5553 (N_5553,N_4086,N_4540);
and U5554 (N_5554,N_4948,N_4047);
nand U5555 (N_5555,N_4332,N_4882);
nor U5556 (N_5556,N_4806,N_4873);
xnor U5557 (N_5557,N_4008,N_4342);
or U5558 (N_5558,N_4019,N_4631);
nor U5559 (N_5559,N_4985,N_4837);
nor U5560 (N_5560,N_4186,N_4769);
nand U5561 (N_5561,N_4936,N_4013);
nand U5562 (N_5562,N_4903,N_4630);
or U5563 (N_5563,N_4013,N_4868);
nor U5564 (N_5564,N_4856,N_4720);
xnor U5565 (N_5565,N_4386,N_4037);
nor U5566 (N_5566,N_4107,N_4517);
nor U5567 (N_5567,N_4769,N_4020);
or U5568 (N_5568,N_4966,N_4617);
nor U5569 (N_5569,N_4764,N_4895);
or U5570 (N_5570,N_4852,N_4663);
and U5571 (N_5571,N_4525,N_4835);
and U5572 (N_5572,N_4328,N_4487);
or U5573 (N_5573,N_4122,N_4410);
xor U5574 (N_5574,N_4185,N_4428);
nand U5575 (N_5575,N_4985,N_4019);
or U5576 (N_5576,N_4319,N_4042);
nand U5577 (N_5577,N_4304,N_4514);
nor U5578 (N_5578,N_4422,N_4011);
nand U5579 (N_5579,N_4266,N_4953);
and U5580 (N_5580,N_4493,N_4836);
nor U5581 (N_5581,N_4966,N_4498);
nor U5582 (N_5582,N_4418,N_4520);
or U5583 (N_5583,N_4908,N_4723);
nand U5584 (N_5584,N_4771,N_4504);
and U5585 (N_5585,N_4118,N_4583);
nor U5586 (N_5586,N_4532,N_4902);
or U5587 (N_5587,N_4380,N_4299);
nand U5588 (N_5588,N_4099,N_4390);
and U5589 (N_5589,N_4786,N_4028);
nor U5590 (N_5590,N_4906,N_4301);
or U5591 (N_5591,N_4492,N_4982);
nand U5592 (N_5592,N_4775,N_4263);
or U5593 (N_5593,N_4226,N_4307);
or U5594 (N_5594,N_4009,N_4184);
nand U5595 (N_5595,N_4005,N_4940);
nor U5596 (N_5596,N_4382,N_4553);
or U5597 (N_5597,N_4941,N_4361);
nor U5598 (N_5598,N_4205,N_4853);
or U5599 (N_5599,N_4888,N_4761);
nand U5600 (N_5600,N_4063,N_4905);
nand U5601 (N_5601,N_4485,N_4591);
nor U5602 (N_5602,N_4928,N_4055);
nor U5603 (N_5603,N_4312,N_4279);
xor U5604 (N_5604,N_4383,N_4189);
and U5605 (N_5605,N_4899,N_4456);
or U5606 (N_5606,N_4162,N_4442);
or U5607 (N_5607,N_4820,N_4230);
and U5608 (N_5608,N_4268,N_4601);
nand U5609 (N_5609,N_4605,N_4372);
and U5610 (N_5610,N_4137,N_4518);
nand U5611 (N_5611,N_4548,N_4745);
nor U5612 (N_5612,N_4973,N_4800);
and U5613 (N_5613,N_4201,N_4326);
or U5614 (N_5614,N_4841,N_4176);
or U5615 (N_5615,N_4548,N_4733);
nor U5616 (N_5616,N_4303,N_4166);
or U5617 (N_5617,N_4699,N_4022);
or U5618 (N_5618,N_4508,N_4502);
nor U5619 (N_5619,N_4922,N_4020);
nand U5620 (N_5620,N_4968,N_4229);
and U5621 (N_5621,N_4805,N_4655);
nand U5622 (N_5622,N_4408,N_4327);
nor U5623 (N_5623,N_4470,N_4241);
xnor U5624 (N_5624,N_4025,N_4651);
and U5625 (N_5625,N_4456,N_4729);
nor U5626 (N_5626,N_4012,N_4450);
nor U5627 (N_5627,N_4327,N_4133);
or U5628 (N_5628,N_4544,N_4111);
nor U5629 (N_5629,N_4751,N_4551);
nor U5630 (N_5630,N_4214,N_4047);
or U5631 (N_5631,N_4554,N_4213);
or U5632 (N_5632,N_4436,N_4101);
or U5633 (N_5633,N_4680,N_4609);
and U5634 (N_5634,N_4228,N_4736);
or U5635 (N_5635,N_4208,N_4367);
and U5636 (N_5636,N_4572,N_4203);
or U5637 (N_5637,N_4855,N_4697);
nor U5638 (N_5638,N_4971,N_4490);
and U5639 (N_5639,N_4397,N_4522);
or U5640 (N_5640,N_4230,N_4895);
nor U5641 (N_5641,N_4827,N_4884);
nor U5642 (N_5642,N_4772,N_4082);
nor U5643 (N_5643,N_4741,N_4585);
nor U5644 (N_5644,N_4206,N_4196);
or U5645 (N_5645,N_4207,N_4876);
and U5646 (N_5646,N_4489,N_4249);
and U5647 (N_5647,N_4848,N_4190);
and U5648 (N_5648,N_4856,N_4443);
nor U5649 (N_5649,N_4402,N_4363);
and U5650 (N_5650,N_4284,N_4694);
or U5651 (N_5651,N_4439,N_4454);
xor U5652 (N_5652,N_4851,N_4173);
nor U5653 (N_5653,N_4691,N_4300);
and U5654 (N_5654,N_4067,N_4811);
nand U5655 (N_5655,N_4969,N_4679);
nor U5656 (N_5656,N_4125,N_4208);
nor U5657 (N_5657,N_4319,N_4480);
and U5658 (N_5658,N_4497,N_4474);
or U5659 (N_5659,N_4926,N_4326);
nand U5660 (N_5660,N_4856,N_4893);
nand U5661 (N_5661,N_4777,N_4889);
nand U5662 (N_5662,N_4017,N_4384);
and U5663 (N_5663,N_4270,N_4585);
nor U5664 (N_5664,N_4502,N_4950);
nand U5665 (N_5665,N_4721,N_4513);
nor U5666 (N_5666,N_4540,N_4932);
and U5667 (N_5667,N_4621,N_4948);
nand U5668 (N_5668,N_4915,N_4405);
and U5669 (N_5669,N_4764,N_4007);
nor U5670 (N_5670,N_4492,N_4517);
nor U5671 (N_5671,N_4481,N_4539);
and U5672 (N_5672,N_4981,N_4836);
or U5673 (N_5673,N_4617,N_4576);
or U5674 (N_5674,N_4041,N_4304);
nand U5675 (N_5675,N_4554,N_4621);
nand U5676 (N_5676,N_4234,N_4660);
nor U5677 (N_5677,N_4580,N_4506);
nand U5678 (N_5678,N_4143,N_4518);
nor U5679 (N_5679,N_4960,N_4505);
or U5680 (N_5680,N_4967,N_4830);
or U5681 (N_5681,N_4053,N_4517);
xor U5682 (N_5682,N_4438,N_4822);
nand U5683 (N_5683,N_4839,N_4665);
nand U5684 (N_5684,N_4153,N_4708);
or U5685 (N_5685,N_4908,N_4178);
nand U5686 (N_5686,N_4451,N_4185);
and U5687 (N_5687,N_4143,N_4497);
or U5688 (N_5688,N_4344,N_4969);
xnor U5689 (N_5689,N_4536,N_4121);
nor U5690 (N_5690,N_4316,N_4883);
nor U5691 (N_5691,N_4858,N_4199);
or U5692 (N_5692,N_4513,N_4285);
nor U5693 (N_5693,N_4668,N_4444);
and U5694 (N_5694,N_4188,N_4553);
or U5695 (N_5695,N_4785,N_4887);
nor U5696 (N_5696,N_4083,N_4031);
xnor U5697 (N_5697,N_4617,N_4918);
xor U5698 (N_5698,N_4915,N_4935);
nand U5699 (N_5699,N_4406,N_4245);
nor U5700 (N_5700,N_4123,N_4529);
or U5701 (N_5701,N_4106,N_4004);
nor U5702 (N_5702,N_4348,N_4691);
or U5703 (N_5703,N_4969,N_4173);
nor U5704 (N_5704,N_4711,N_4187);
nor U5705 (N_5705,N_4799,N_4483);
or U5706 (N_5706,N_4326,N_4231);
nand U5707 (N_5707,N_4510,N_4480);
and U5708 (N_5708,N_4204,N_4123);
or U5709 (N_5709,N_4384,N_4100);
xor U5710 (N_5710,N_4661,N_4118);
nand U5711 (N_5711,N_4832,N_4652);
or U5712 (N_5712,N_4945,N_4519);
nand U5713 (N_5713,N_4114,N_4365);
or U5714 (N_5714,N_4786,N_4544);
nor U5715 (N_5715,N_4651,N_4567);
nand U5716 (N_5716,N_4998,N_4910);
xor U5717 (N_5717,N_4843,N_4414);
or U5718 (N_5718,N_4820,N_4570);
nor U5719 (N_5719,N_4159,N_4078);
nand U5720 (N_5720,N_4994,N_4621);
or U5721 (N_5721,N_4597,N_4933);
nand U5722 (N_5722,N_4445,N_4536);
and U5723 (N_5723,N_4689,N_4912);
or U5724 (N_5724,N_4527,N_4472);
and U5725 (N_5725,N_4472,N_4089);
nor U5726 (N_5726,N_4787,N_4339);
nand U5727 (N_5727,N_4019,N_4962);
xnor U5728 (N_5728,N_4906,N_4382);
nand U5729 (N_5729,N_4974,N_4702);
nor U5730 (N_5730,N_4090,N_4991);
and U5731 (N_5731,N_4712,N_4846);
nor U5732 (N_5732,N_4673,N_4636);
and U5733 (N_5733,N_4732,N_4967);
nor U5734 (N_5734,N_4703,N_4872);
nor U5735 (N_5735,N_4672,N_4844);
nor U5736 (N_5736,N_4186,N_4914);
nor U5737 (N_5737,N_4782,N_4340);
nor U5738 (N_5738,N_4402,N_4674);
nand U5739 (N_5739,N_4381,N_4035);
nand U5740 (N_5740,N_4092,N_4743);
and U5741 (N_5741,N_4703,N_4491);
and U5742 (N_5742,N_4896,N_4409);
and U5743 (N_5743,N_4574,N_4005);
and U5744 (N_5744,N_4538,N_4252);
nor U5745 (N_5745,N_4258,N_4499);
nand U5746 (N_5746,N_4547,N_4156);
nor U5747 (N_5747,N_4167,N_4621);
nor U5748 (N_5748,N_4835,N_4860);
or U5749 (N_5749,N_4878,N_4386);
or U5750 (N_5750,N_4085,N_4008);
nand U5751 (N_5751,N_4590,N_4257);
nand U5752 (N_5752,N_4966,N_4141);
and U5753 (N_5753,N_4177,N_4111);
nor U5754 (N_5754,N_4962,N_4561);
nand U5755 (N_5755,N_4203,N_4343);
or U5756 (N_5756,N_4531,N_4004);
nand U5757 (N_5757,N_4446,N_4256);
and U5758 (N_5758,N_4968,N_4262);
nor U5759 (N_5759,N_4892,N_4248);
and U5760 (N_5760,N_4622,N_4940);
nand U5761 (N_5761,N_4800,N_4269);
and U5762 (N_5762,N_4291,N_4175);
nor U5763 (N_5763,N_4330,N_4002);
nand U5764 (N_5764,N_4809,N_4072);
or U5765 (N_5765,N_4408,N_4256);
xnor U5766 (N_5766,N_4131,N_4679);
nor U5767 (N_5767,N_4644,N_4401);
nand U5768 (N_5768,N_4173,N_4438);
nor U5769 (N_5769,N_4394,N_4622);
nand U5770 (N_5770,N_4179,N_4156);
or U5771 (N_5771,N_4083,N_4701);
xnor U5772 (N_5772,N_4805,N_4389);
nor U5773 (N_5773,N_4947,N_4468);
nor U5774 (N_5774,N_4849,N_4453);
or U5775 (N_5775,N_4751,N_4370);
nand U5776 (N_5776,N_4450,N_4791);
or U5777 (N_5777,N_4672,N_4771);
or U5778 (N_5778,N_4829,N_4956);
nor U5779 (N_5779,N_4654,N_4521);
nand U5780 (N_5780,N_4195,N_4164);
nand U5781 (N_5781,N_4352,N_4026);
or U5782 (N_5782,N_4099,N_4010);
and U5783 (N_5783,N_4916,N_4650);
or U5784 (N_5784,N_4122,N_4069);
nor U5785 (N_5785,N_4662,N_4903);
nor U5786 (N_5786,N_4056,N_4633);
nor U5787 (N_5787,N_4673,N_4104);
nand U5788 (N_5788,N_4173,N_4897);
or U5789 (N_5789,N_4826,N_4272);
or U5790 (N_5790,N_4510,N_4905);
or U5791 (N_5791,N_4864,N_4815);
nor U5792 (N_5792,N_4057,N_4428);
and U5793 (N_5793,N_4457,N_4922);
nor U5794 (N_5794,N_4183,N_4827);
nand U5795 (N_5795,N_4031,N_4388);
nand U5796 (N_5796,N_4490,N_4680);
nand U5797 (N_5797,N_4229,N_4394);
or U5798 (N_5798,N_4348,N_4873);
nor U5799 (N_5799,N_4867,N_4631);
and U5800 (N_5800,N_4691,N_4518);
or U5801 (N_5801,N_4088,N_4966);
nor U5802 (N_5802,N_4582,N_4940);
or U5803 (N_5803,N_4564,N_4587);
nand U5804 (N_5804,N_4192,N_4127);
nor U5805 (N_5805,N_4765,N_4494);
nor U5806 (N_5806,N_4387,N_4708);
and U5807 (N_5807,N_4689,N_4481);
nor U5808 (N_5808,N_4179,N_4734);
nand U5809 (N_5809,N_4833,N_4467);
nor U5810 (N_5810,N_4976,N_4660);
nor U5811 (N_5811,N_4487,N_4655);
or U5812 (N_5812,N_4818,N_4540);
nor U5813 (N_5813,N_4998,N_4802);
nor U5814 (N_5814,N_4068,N_4681);
nand U5815 (N_5815,N_4554,N_4396);
nand U5816 (N_5816,N_4470,N_4445);
nor U5817 (N_5817,N_4669,N_4470);
and U5818 (N_5818,N_4401,N_4005);
nor U5819 (N_5819,N_4164,N_4771);
or U5820 (N_5820,N_4359,N_4031);
and U5821 (N_5821,N_4485,N_4645);
xor U5822 (N_5822,N_4913,N_4994);
nand U5823 (N_5823,N_4944,N_4308);
nand U5824 (N_5824,N_4340,N_4384);
and U5825 (N_5825,N_4675,N_4406);
or U5826 (N_5826,N_4935,N_4618);
nand U5827 (N_5827,N_4989,N_4774);
nand U5828 (N_5828,N_4948,N_4830);
nand U5829 (N_5829,N_4450,N_4135);
and U5830 (N_5830,N_4569,N_4870);
nand U5831 (N_5831,N_4047,N_4521);
nand U5832 (N_5832,N_4683,N_4522);
or U5833 (N_5833,N_4478,N_4144);
or U5834 (N_5834,N_4353,N_4965);
and U5835 (N_5835,N_4584,N_4935);
or U5836 (N_5836,N_4140,N_4984);
and U5837 (N_5837,N_4778,N_4424);
nor U5838 (N_5838,N_4649,N_4968);
or U5839 (N_5839,N_4482,N_4930);
and U5840 (N_5840,N_4227,N_4592);
and U5841 (N_5841,N_4328,N_4151);
and U5842 (N_5842,N_4849,N_4276);
nor U5843 (N_5843,N_4958,N_4152);
nand U5844 (N_5844,N_4441,N_4677);
or U5845 (N_5845,N_4307,N_4562);
and U5846 (N_5846,N_4136,N_4412);
or U5847 (N_5847,N_4650,N_4647);
xnor U5848 (N_5848,N_4237,N_4475);
nor U5849 (N_5849,N_4137,N_4997);
or U5850 (N_5850,N_4948,N_4177);
nand U5851 (N_5851,N_4666,N_4565);
nor U5852 (N_5852,N_4029,N_4585);
nor U5853 (N_5853,N_4303,N_4586);
or U5854 (N_5854,N_4259,N_4168);
or U5855 (N_5855,N_4772,N_4596);
and U5856 (N_5856,N_4482,N_4048);
or U5857 (N_5857,N_4969,N_4307);
or U5858 (N_5858,N_4184,N_4962);
or U5859 (N_5859,N_4108,N_4371);
and U5860 (N_5860,N_4161,N_4769);
and U5861 (N_5861,N_4445,N_4848);
nand U5862 (N_5862,N_4822,N_4724);
nand U5863 (N_5863,N_4529,N_4121);
or U5864 (N_5864,N_4944,N_4572);
nor U5865 (N_5865,N_4266,N_4947);
or U5866 (N_5866,N_4328,N_4970);
and U5867 (N_5867,N_4359,N_4365);
nor U5868 (N_5868,N_4082,N_4417);
or U5869 (N_5869,N_4917,N_4657);
and U5870 (N_5870,N_4883,N_4143);
nand U5871 (N_5871,N_4462,N_4918);
and U5872 (N_5872,N_4319,N_4180);
and U5873 (N_5873,N_4495,N_4847);
nand U5874 (N_5874,N_4032,N_4977);
and U5875 (N_5875,N_4256,N_4513);
nand U5876 (N_5876,N_4903,N_4336);
and U5877 (N_5877,N_4872,N_4043);
nor U5878 (N_5878,N_4515,N_4572);
or U5879 (N_5879,N_4439,N_4386);
and U5880 (N_5880,N_4913,N_4935);
or U5881 (N_5881,N_4973,N_4055);
or U5882 (N_5882,N_4334,N_4508);
nand U5883 (N_5883,N_4730,N_4579);
nor U5884 (N_5884,N_4573,N_4753);
xor U5885 (N_5885,N_4972,N_4621);
and U5886 (N_5886,N_4351,N_4044);
nor U5887 (N_5887,N_4543,N_4340);
and U5888 (N_5888,N_4485,N_4269);
and U5889 (N_5889,N_4191,N_4538);
nor U5890 (N_5890,N_4587,N_4393);
and U5891 (N_5891,N_4745,N_4496);
or U5892 (N_5892,N_4851,N_4440);
and U5893 (N_5893,N_4004,N_4543);
nor U5894 (N_5894,N_4268,N_4959);
nand U5895 (N_5895,N_4765,N_4096);
and U5896 (N_5896,N_4034,N_4454);
and U5897 (N_5897,N_4153,N_4561);
nand U5898 (N_5898,N_4008,N_4111);
nand U5899 (N_5899,N_4432,N_4286);
or U5900 (N_5900,N_4252,N_4193);
or U5901 (N_5901,N_4121,N_4495);
or U5902 (N_5902,N_4621,N_4711);
nor U5903 (N_5903,N_4851,N_4976);
or U5904 (N_5904,N_4010,N_4888);
or U5905 (N_5905,N_4123,N_4117);
and U5906 (N_5906,N_4789,N_4730);
xor U5907 (N_5907,N_4274,N_4750);
and U5908 (N_5908,N_4004,N_4157);
nor U5909 (N_5909,N_4437,N_4169);
nand U5910 (N_5910,N_4963,N_4821);
nor U5911 (N_5911,N_4308,N_4267);
nand U5912 (N_5912,N_4332,N_4098);
nand U5913 (N_5913,N_4852,N_4918);
and U5914 (N_5914,N_4121,N_4818);
and U5915 (N_5915,N_4761,N_4821);
nor U5916 (N_5916,N_4396,N_4693);
nor U5917 (N_5917,N_4799,N_4781);
nand U5918 (N_5918,N_4379,N_4419);
nor U5919 (N_5919,N_4538,N_4279);
nor U5920 (N_5920,N_4621,N_4611);
or U5921 (N_5921,N_4703,N_4073);
or U5922 (N_5922,N_4219,N_4651);
or U5923 (N_5923,N_4755,N_4190);
nor U5924 (N_5924,N_4064,N_4208);
nor U5925 (N_5925,N_4598,N_4782);
or U5926 (N_5926,N_4454,N_4550);
nor U5927 (N_5927,N_4184,N_4795);
nand U5928 (N_5928,N_4535,N_4498);
nand U5929 (N_5929,N_4415,N_4755);
and U5930 (N_5930,N_4106,N_4138);
nor U5931 (N_5931,N_4829,N_4567);
nor U5932 (N_5932,N_4253,N_4789);
or U5933 (N_5933,N_4115,N_4392);
nor U5934 (N_5934,N_4611,N_4982);
and U5935 (N_5935,N_4370,N_4619);
and U5936 (N_5936,N_4742,N_4232);
and U5937 (N_5937,N_4363,N_4937);
nor U5938 (N_5938,N_4693,N_4478);
and U5939 (N_5939,N_4551,N_4352);
nor U5940 (N_5940,N_4762,N_4359);
nand U5941 (N_5941,N_4883,N_4334);
nand U5942 (N_5942,N_4903,N_4038);
or U5943 (N_5943,N_4177,N_4699);
nand U5944 (N_5944,N_4963,N_4630);
nor U5945 (N_5945,N_4569,N_4703);
and U5946 (N_5946,N_4341,N_4004);
nor U5947 (N_5947,N_4746,N_4030);
nor U5948 (N_5948,N_4791,N_4315);
nand U5949 (N_5949,N_4990,N_4780);
nor U5950 (N_5950,N_4653,N_4903);
nor U5951 (N_5951,N_4646,N_4428);
xnor U5952 (N_5952,N_4657,N_4888);
and U5953 (N_5953,N_4401,N_4108);
and U5954 (N_5954,N_4979,N_4254);
xor U5955 (N_5955,N_4328,N_4741);
and U5956 (N_5956,N_4932,N_4930);
nor U5957 (N_5957,N_4648,N_4369);
nand U5958 (N_5958,N_4505,N_4481);
nand U5959 (N_5959,N_4468,N_4554);
and U5960 (N_5960,N_4753,N_4457);
or U5961 (N_5961,N_4815,N_4083);
nand U5962 (N_5962,N_4673,N_4465);
nor U5963 (N_5963,N_4557,N_4826);
and U5964 (N_5964,N_4574,N_4347);
nand U5965 (N_5965,N_4009,N_4839);
or U5966 (N_5966,N_4955,N_4672);
and U5967 (N_5967,N_4903,N_4163);
or U5968 (N_5968,N_4382,N_4944);
nand U5969 (N_5969,N_4195,N_4248);
nand U5970 (N_5970,N_4005,N_4784);
or U5971 (N_5971,N_4499,N_4642);
or U5972 (N_5972,N_4846,N_4457);
nor U5973 (N_5973,N_4889,N_4087);
and U5974 (N_5974,N_4132,N_4327);
nor U5975 (N_5975,N_4502,N_4965);
or U5976 (N_5976,N_4388,N_4625);
or U5977 (N_5977,N_4425,N_4083);
and U5978 (N_5978,N_4288,N_4588);
or U5979 (N_5979,N_4175,N_4375);
nand U5980 (N_5980,N_4864,N_4609);
nand U5981 (N_5981,N_4963,N_4367);
nand U5982 (N_5982,N_4476,N_4049);
nor U5983 (N_5983,N_4934,N_4849);
or U5984 (N_5984,N_4421,N_4760);
xnor U5985 (N_5985,N_4768,N_4111);
and U5986 (N_5986,N_4738,N_4313);
nor U5987 (N_5987,N_4230,N_4199);
nand U5988 (N_5988,N_4213,N_4688);
nand U5989 (N_5989,N_4543,N_4842);
or U5990 (N_5990,N_4915,N_4397);
nand U5991 (N_5991,N_4368,N_4759);
nand U5992 (N_5992,N_4725,N_4061);
nand U5993 (N_5993,N_4872,N_4915);
nor U5994 (N_5994,N_4514,N_4069);
nand U5995 (N_5995,N_4985,N_4190);
nor U5996 (N_5996,N_4926,N_4492);
nand U5997 (N_5997,N_4098,N_4960);
nand U5998 (N_5998,N_4037,N_4385);
or U5999 (N_5999,N_4953,N_4738);
nand U6000 (N_6000,N_5848,N_5141);
and U6001 (N_6001,N_5833,N_5021);
nor U6002 (N_6002,N_5253,N_5987);
and U6003 (N_6003,N_5338,N_5049);
nor U6004 (N_6004,N_5305,N_5990);
or U6005 (N_6005,N_5301,N_5358);
nand U6006 (N_6006,N_5834,N_5551);
and U6007 (N_6007,N_5667,N_5095);
and U6008 (N_6008,N_5793,N_5383);
nor U6009 (N_6009,N_5539,N_5210);
nand U6010 (N_6010,N_5438,N_5757);
and U6011 (N_6011,N_5492,N_5318);
and U6012 (N_6012,N_5302,N_5405);
nand U6013 (N_6013,N_5138,N_5741);
and U6014 (N_6014,N_5533,N_5634);
or U6015 (N_6015,N_5411,N_5925);
or U6016 (N_6016,N_5408,N_5343);
nor U6017 (N_6017,N_5291,N_5867);
nand U6018 (N_6018,N_5683,N_5165);
and U6019 (N_6019,N_5929,N_5749);
nor U6020 (N_6020,N_5842,N_5797);
nor U6021 (N_6021,N_5384,N_5190);
nor U6022 (N_6022,N_5538,N_5317);
or U6023 (N_6023,N_5396,N_5732);
or U6024 (N_6024,N_5537,N_5666);
nand U6025 (N_6025,N_5006,N_5450);
and U6026 (N_6026,N_5824,N_5646);
nor U6027 (N_6027,N_5541,N_5944);
and U6028 (N_6028,N_5489,N_5314);
nand U6029 (N_6029,N_5671,N_5898);
nand U6030 (N_6030,N_5599,N_5163);
and U6031 (N_6031,N_5779,N_5642);
and U6032 (N_6032,N_5673,N_5407);
or U6033 (N_6033,N_5373,N_5258);
or U6034 (N_6034,N_5044,N_5563);
nor U6035 (N_6035,N_5289,N_5410);
nand U6036 (N_6036,N_5882,N_5730);
or U6037 (N_6037,N_5160,N_5084);
nor U6038 (N_6038,N_5062,N_5085);
or U6039 (N_6039,N_5886,N_5781);
nand U6040 (N_6040,N_5452,N_5211);
nand U6041 (N_6041,N_5355,N_5294);
nor U6042 (N_6042,N_5065,N_5575);
or U6043 (N_6043,N_5821,N_5958);
and U6044 (N_6044,N_5823,N_5512);
nor U6045 (N_6045,N_5056,N_5625);
nor U6046 (N_6046,N_5287,N_5529);
nor U6047 (N_6047,N_5904,N_5024);
or U6048 (N_6048,N_5152,N_5030);
nand U6049 (N_6049,N_5362,N_5515);
nand U6050 (N_6050,N_5376,N_5369);
or U6051 (N_6051,N_5572,N_5052);
and U6052 (N_6052,N_5354,N_5387);
xnor U6053 (N_6053,N_5285,N_5893);
or U6054 (N_6054,N_5943,N_5491);
or U6055 (N_6055,N_5744,N_5696);
nor U6056 (N_6056,N_5914,N_5991);
or U6057 (N_6057,N_5618,N_5184);
nor U6058 (N_6058,N_5207,N_5416);
nor U6059 (N_6059,N_5272,N_5193);
and U6060 (N_6060,N_5947,N_5262);
and U6061 (N_6061,N_5892,N_5585);
or U6062 (N_6062,N_5829,N_5574);
and U6063 (N_6063,N_5009,N_5584);
or U6064 (N_6064,N_5740,N_5462);
nor U6065 (N_6065,N_5609,N_5051);
nor U6066 (N_6066,N_5391,N_5276);
and U6067 (N_6067,N_5068,N_5337);
or U6068 (N_6068,N_5487,N_5280);
and U6069 (N_6069,N_5994,N_5425);
and U6070 (N_6070,N_5257,N_5299);
or U6071 (N_6071,N_5135,N_5791);
nand U6072 (N_6072,N_5669,N_5508);
nand U6073 (N_6073,N_5891,N_5389);
and U6074 (N_6074,N_5436,N_5706);
nor U6075 (N_6075,N_5493,N_5229);
or U6076 (N_6076,N_5869,N_5456);
and U6077 (N_6077,N_5132,N_5327);
xnor U6078 (N_6078,N_5308,N_5061);
nor U6079 (N_6079,N_5303,N_5951);
nor U6080 (N_6080,N_5116,N_5079);
or U6081 (N_6081,N_5169,N_5888);
nand U6082 (N_6082,N_5738,N_5709);
nand U6083 (N_6083,N_5345,N_5502);
or U6084 (N_6084,N_5249,N_5698);
and U6085 (N_6085,N_5478,N_5640);
nand U6086 (N_6086,N_5873,N_5617);
or U6087 (N_6087,N_5370,N_5969);
nor U6088 (N_6088,N_5259,N_5764);
nand U6089 (N_6089,N_5861,N_5759);
nor U6090 (N_6090,N_5128,N_5550);
nor U6091 (N_6091,N_5907,N_5518);
nand U6092 (N_6092,N_5035,N_5535);
or U6093 (N_6093,N_5279,N_5765);
or U6094 (N_6094,N_5310,N_5392);
and U6095 (N_6095,N_5610,N_5260);
nor U6096 (N_6096,N_5427,N_5737);
nand U6097 (N_6097,N_5374,N_5560);
nand U6098 (N_6098,N_5729,N_5763);
or U6099 (N_6099,N_5615,N_5507);
nand U6100 (N_6100,N_5244,N_5311);
and U6101 (N_6101,N_5500,N_5851);
or U6102 (N_6102,N_5554,N_5209);
and U6103 (N_6103,N_5909,N_5724);
and U6104 (N_6104,N_5269,N_5498);
xnor U6105 (N_6105,N_5880,N_5826);
nand U6106 (N_6106,N_5717,N_5570);
nor U6107 (N_6107,N_5034,N_5927);
and U6108 (N_6108,N_5840,N_5134);
or U6109 (N_6109,N_5736,N_5393);
nand U6110 (N_6110,N_5017,N_5961);
or U6111 (N_6111,N_5964,N_5041);
or U6112 (N_6112,N_5072,N_5720);
or U6113 (N_6113,N_5655,N_5334);
nand U6114 (N_6114,N_5549,N_5237);
nand U6115 (N_6115,N_5012,N_5164);
nor U6116 (N_6116,N_5651,N_5449);
nand U6117 (N_6117,N_5708,N_5526);
nor U6118 (N_6118,N_5999,N_5045);
nand U6119 (N_6119,N_5479,N_5379);
nor U6120 (N_6120,N_5812,N_5693);
and U6121 (N_6121,N_5963,N_5441);
and U6122 (N_6122,N_5212,N_5790);
nor U6123 (N_6123,N_5418,N_5948);
nand U6124 (N_6124,N_5633,N_5876);
and U6125 (N_6125,N_5081,N_5581);
nor U6126 (N_6126,N_5320,N_5566);
and U6127 (N_6127,N_5647,N_5710);
or U6128 (N_6128,N_5144,N_5265);
nor U6129 (N_6129,N_5366,N_5966);
and U6130 (N_6130,N_5010,N_5348);
nor U6131 (N_6131,N_5553,N_5819);
nand U6132 (N_6132,N_5868,N_5684);
nor U6133 (N_6133,N_5118,N_5274);
nand U6134 (N_6134,N_5723,N_5154);
nand U6135 (N_6135,N_5266,N_5580);
or U6136 (N_6136,N_5286,N_5126);
nor U6137 (N_6137,N_5573,N_5205);
nand U6138 (N_6138,N_5780,N_5748);
and U6139 (N_6139,N_5579,N_5546);
nand U6140 (N_6140,N_5182,N_5847);
nand U6141 (N_6141,N_5364,N_5103);
nor U6142 (N_6142,N_5620,N_5926);
or U6143 (N_6143,N_5101,N_5481);
nor U6144 (N_6144,N_5234,N_5372);
and U6145 (N_6145,N_5578,N_5149);
and U6146 (N_6146,N_5428,N_5545);
or U6147 (N_6147,N_5915,N_5071);
and U6148 (N_6148,N_5798,N_5517);
and U6149 (N_6149,N_5335,N_5505);
nand U6150 (N_6150,N_5476,N_5340);
and U6151 (N_6151,N_5363,N_5704);
nor U6152 (N_6152,N_5050,N_5202);
and U6153 (N_6153,N_5971,N_5858);
xnor U6154 (N_6154,N_5702,N_5268);
and U6155 (N_6155,N_5176,N_5668);
and U6156 (N_6156,N_5424,N_5046);
and U6157 (N_6157,N_5766,N_5214);
or U6158 (N_6158,N_5356,N_5241);
and U6159 (N_6159,N_5658,N_5697);
nand U6160 (N_6160,N_5716,N_5722);
nor U6161 (N_6161,N_5622,N_5175);
or U6162 (N_6162,N_5104,N_5739);
nand U6163 (N_6163,N_5296,N_5544);
nand U6164 (N_6164,N_5236,N_5040);
xnor U6165 (N_6165,N_5001,N_5036);
and U6166 (N_6166,N_5004,N_5980);
nor U6167 (N_6167,N_5231,N_5621);
nor U6168 (N_6168,N_5965,N_5552);
and U6169 (N_6169,N_5180,N_5931);
or U6170 (N_6170,N_5339,N_5271);
or U6171 (N_6171,N_5807,N_5174);
and U6172 (N_6172,N_5083,N_5460);
nand U6173 (N_6173,N_5381,N_5419);
or U6174 (N_6174,N_5769,N_5801);
and U6175 (N_6175,N_5974,N_5523);
and U6176 (N_6176,N_5557,N_5583);
or U6177 (N_6177,N_5592,N_5270);
nand U6178 (N_6178,N_5525,N_5319);
nand U6179 (N_6179,N_5057,N_5707);
nor U6180 (N_6180,N_5775,N_5839);
and U6181 (N_6181,N_5995,N_5119);
and U6182 (N_6182,N_5090,N_5559);
xor U6183 (N_6183,N_5813,N_5582);
nand U6184 (N_6184,N_5000,N_5605);
and U6185 (N_6185,N_5879,N_5347);
xnor U6186 (N_6186,N_5242,N_5604);
xor U6187 (N_6187,N_5199,N_5243);
nor U6188 (N_6188,N_5981,N_5235);
nand U6189 (N_6189,N_5501,N_5323);
or U6190 (N_6190,N_5624,N_5192);
and U6191 (N_6191,N_5412,N_5458);
xor U6192 (N_6192,N_5254,N_5705);
nand U6193 (N_6193,N_5540,N_5222);
or U6194 (N_6194,N_5043,N_5881);
nor U6195 (N_6195,N_5316,N_5569);
nor U6196 (N_6196,N_5718,N_5467);
nand U6197 (N_6197,N_5166,N_5466);
xnor U6198 (N_6198,N_5186,N_5196);
or U6199 (N_6199,N_5435,N_5714);
and U6200 (N_6200,N_5855,N_5039);
or U6201 (N_6201,N_5332,N_5735);
or U6202 (N_6202,N_5497,N_5437);
nand U6203 (N_6203,N_5465,N_5528);
xor U6204 (N_6204,N_5787,N_5018);
or U6205 (N_6205,N_5828,N_5913);
or U6206 (N_6206,N_5984,N_5679);
and U6207 (N_6207,N_5850,N_5681);
or U6208 (N_6208,N_5457,N_5070);
nor U6209 (N_6209,N_5283,N_5972);
nor U6210 (N_6210,N_5031,N_5108);
or U6211 (N_6211,N_5406,N_5692);
nor U6212 (N_6212,N_5946,N_5002);
or U6213 (N_6213,N_5923,N_5688);
nand U6214 (N_6214,N_5288,N_5504);
nor U6215 (N_6215,N_5066,N_5386);
or U6216 (N_6216,N_5495,N_5415);
nand U6217 (N_6217,N_5510,N_5985);
or U6218 (N_6218,N_5155,N_5921);
xor U6219 (N_6219,N_5019,N_5076);
or U6220 (N_6220,N_5020,N_5426);
nand U6221 (N_6221,N_5611,N_5371);
or U6222 (N_6222,N_5854,N_5808);
xnor U6223 (N_6223,N_5409,N_5659);
nand U6224 (N_6224,N_5281,N_5173);
nand U6225 (N_6225,N_5639,N_5261);
and U6226 (N_6226,N_5846,N_5794);
or U6227 (N_6227,N_5256,N_5792);
nand U6228 (N_6228,N_5635,N_5420);
nor U6229 (N_6229,N_5513,N_5967);
nand U6230 (N_6230,N_5007,N_5142);
or U6231 (N_6231,N_5413,N_5900);
nand U6232 (N_6232,N_5630,N_5774);
nand U6233 (N_6233,N_5799,N_5509);
nor U6234 (N_6234,N_5077,N_5607);
or U6235 (N_6235,N_5295,N_5430);
nand U6236 (N_6236,N_5565,N_5171);
or U6237 (N_6237,N_5827,N_5168);
or U6238 (N_6238,N_5555,N_5472);
nor U6239 (N_6239,N_5177,N_5013);
nor U6240 (N_6240,N_5567,N_5664);
and U6241 (N_6241,N_5970,N_5564);
nor U6242 (N_6242,N_5852,N_5751);
nand U6243 (N_6243,N_5400,N_5014);
or U6244 (N_6244,N_5473,N_5073);
and U6245 (N_6245,N_5357,N_5298);
nand U6246 (N_6246,N_5753,N_5742);
and U6247 (N_6247,N_5015,N_5960);
nand U6248 (N_6248,N_5940,N_5894);
or U6249 (N_6249,N_5631,N_5150);
nor U6250 (N_6250,N_5404,N_5147);
or U6251 (N_6251,N_5841,N_5315);
nor U6252 (N_6252,N_5112,N_5747);
and U6253 (N_6253,N_5005,N_5521);
nor U6254 (N_6254,N_5760,N_5455);
nand U6255 (N_6255,N_5871,N_5663);
or U6256 (N_6256,N_5482,N_5156);
nor U6257 (N_6257,N_5058,N_5962);
and U6258 (N_6258,N_5378,N_5571);
and U6259 (N_6259,N_5477,N_5527);
nor U6260 (N_6260,N_5843,N_5422);
or U6261 (N_6261,N_5350,N_5758);
or U6262 (N_6262,N_5761,N_5092);
or U6263 (N_6263,N_5752,N_5522);
and U6264 (N_6264,N_5161,N_5403);
or U6265 (N_6265,N_5952,N_5830);
nor U6266 (N_6266,N_5989,N_5776);
nand U6267 (N_6267,N_5726,N_5377);
nand U6268 (N_6268,N_5390,N_5206);
nand U6269 (N_6269,N_5835,N_5930);
or U6270 (N_6270,N_5292,N_5221);
nand U6271 (N_6271,N_5181,N_5531);
nand U6272 (N_6272,N_5795,N_5938);
and U6273 (N_6273,N_5945,N_5804);
and U6274 (N_6274,N_5360,N_5796);
nand U6275 (N_6275,N_5053,N_5815);
nor U6276 (N_6276,N_5576,N_5686);
nor U6277 (N_6277,N_5448,N_5048);
or U6278 (N_6278,N_5883,N_5973);
nand U6279 (N_6279,N_5468,N_5542);
nor U6280 (N_6280,N_5859,N_5198);
nor U6281 (N_6281,N_5649,N_5800);
and U6282 (N_6282,N_5113,N_5145);
or U6283 (N_6283,N_5297,N_5956);
nand U6284 (N_6284,N_5548,N_5516);
or U6285 (N_6285,N_5591,N_5897);
and U6286 (N_6286,N_5088,N_5245);
or U6287 (N_6287,N_5300,N_5628);
nand U6288 (N_6288,N_5695,N_5711);
nor U6289 (N_6289,N_5324,N_5399);
nand U6290 (N_6290,N_5148,N_5082);
nor U6291 (N_6291,N_5157,N_5650);
nor U6292 (N_6292,N_5240,N_5398);
nand U6293 (N_6293,N_5106,N_5028);
xnor U6294 (N_6294,N_5762,N_5195);
nand U6295 (N_6295,N_5225,N_5250);
or U6296 (N_6296,N_5342,N_5187);
and U6297 (N_6297,N_5837,N_5784);
or U6298 (N_6298,N_5115,N_5469);
xor U6299 (N_6299,N_5238,N_5033);
nand U6300 (N_6300,N_5100,N_5474);
nand U6301 (N_6301,N_5375,N_5179);
nor U6302 (N_6302,N_5352,N_5331);
nand U6303 (N_6303,N_5822,N_5414);
nand U6304 (N_6304,N_5330,N_5601);
or U6305 (N_6305,N_5853,N_5228);
and U6306 (N_6306,N_5110,N_5949);
and U6307 (N_6307,N_5080,N_5887);
nor U6308 (N_6308,N_5439,N_5086);
nor U6309 (N_6309,N_5998,N_5870);
nand U6310 (N_6310,N_5820,N_5463);
and U6311 (N_6311,N_5594,N_5992);
or U6312 (N_6312,N_5977,N_5768);
and U6313 (N_6313,N_5277,N_5032);
and U6314 (N_6314,N_5983,N_5503);
and U6315 (N_6315,N_5170,N_5197);
and U6316 (N_6316,N_5637,N_5789);
nand U6317 (N_6317,N_5562,N_5865);
xnor U6318 (N_6318,N_5255,N_5120);
xor U6319 (N_6319,N_5968,N_5614);
nand U6320 (N_6320,N_5444,N_5454);
xor U6321 (N_6321,N_5252,N_5219);
nor U6322 (N_6322,N_5590,N_5933);
nor U6323 (N_6323,N_5485,N_5442);
nand U6324 (N_6324,N_5661,N_5220);
and U6325 (N_6325,N_5899,N_5862);
nand U6326 (N_6326,N_5464,N_5770);
nand U6327 (N_6327,N_5682,N_5459);
nor U6328 (N_6328,N_5959,N_5874);
nor U6329 (N_6329,N_5860,N_5447);
and U6330 (N_6330,N_5644,N_5385);
and U6331 (N_6331,N_5975,N_5486);
and U6332 (N_6332,N_5519,N_5587);
and U6333 (N_6333,N_5825,N_5623);
nand U6334 (N_6334,N_5475,N_5434);
nand U6335 (N_6335,N_5836,N_5603);
or U6336 (N_6336,N_5122,N_5136);
nand U6337 (N_6337,N_5616,N_5896);
nand U6338 (N_6338,N_5885,N_5857);
or U6339 (N_6339,N_5499,N_5638);
nor U6340 (N_6340,N_5514,N_5188);
or U6341 (N_6341,N_5151,N_5670);
and U6342 (N_6342,N_5461,N_5232);
nor U6343 (N_6343,N_5304,N_5351);
and U6344 (N_6344,N_5189,N_5172);
or U6345 (N_6345,N_5431,N_5856);
or U6346 (N_6346,N_5451,N_5606);
nand U6347 (N_6347,N_5380,N_5123);
nor U6348 (N_6348,N_5676,N_5201);
nor U6349 (N_6349,N_5251,N_5936);
nor U6350 (N_6350,N_5941,N_5312);
and U6351 (N_6351,N_5532,N_5440);
or U6352 (N_6352,N_5719,N_5109);
nand U6353 (N_6353,N_5890,N_5809);
or U6354 (N_6354,N_5783,N_5786);
and U6355 (N_6355,N_5713,N_5785);
and U6356 (N_6356,N_5680,N_5916);
and U6357 (N_6357,N_5361,N_5677);
nor U6358 (N_6358,N_5613,N_5042);
and U6359 (N_6359,N_5596,N_5932);
or U6360 (N_6360,N_5908,N_5208);
nor U6361 (N_6361,N_5657,N_5388);
nand U6362 (N_6362,N_5600,N_5227);
nand U6363 (N_6363,N_5645,N_5832);
nand U6364 (N_6364,N_5026,N_5648);
nand U6365 (N_6365,N_5248,N_5233);
or U6366 (N_6366,N_5098,N_5107);
nand U6367 (N_6367,N_5217,N_5367);
and U6368 (N_6368,N_5619,N_5520);
nor U6369 (N_6369,N_5656,N_5275);
nand U6370 (N_6370,N_5875,N_5223);
nor U6371 (N_6371,N_5105,N_5102);
or U6372 (N_6372,N_5845,N_5950);
or U6373 (N_6373,N_5029,N_5060);
nor U6374 (N_6374,N_5325,N_5771);
nand U6375 (N_6375,N_5675,N_5247);
or U6376 (N_6376,N_5063,N_5097);
nor U6377 (N_6377,N_5685,N_5778);
or U6378 (N_6378,N_5586,N_5423);
and U6379 (N_6379,N_5877,N_5471);
nor U6380 (N_6380,N_5359,N_5889);
nand U6381 (N_6381,N_5701,N_5937);
and U6382 (N_6382,N_5712,N_5397);
nand U6383 (N_6383,N_5153,N_5745);
or U6384 (N_6384,N_5588,N_5446);
and U6385 (N_6385,N_5678,N_5731);
or U6386 (N_6386,N_5114,N_5577);
nor U6387 (N_6387,N_5593,N_5831);
nand U6388 (N_6388,N_5922,N_5878);
nor U6389 (N_6389,N_5755,N_5353);
nand U6390 (N_6390,N_5864,N_5777);
nand U6391 (N_6391,N_5912,N_5750);
and U6392 (N_6392,N_5928,N_5011);
and U6393 (N_6393,N_5127,N_5178);
nand U6394 (N_6394,N_5556,N_5125);
xnor U6395 (N_6395,N_5313,N_5986);
or U6396 (N_6396,N_5534,N_5849);
nor U6397 (N_6397,N_5918,N_5075);
nand U6398 (N_6398,N_5595,N_5365);
and U6399 (N_6399,N_5293,N_5121);
or U6400 (N_6400,N_5494,N_5906);
nor U6401 (N_6401,N_5782,N_5674);
and U6402 (N_6402,N_5612,N_5810);
nand U6403 (N_6403,N_5733,N_5417);
or U6404 (N_6404,N_5699,N_5204);
or U6405 (N_6405,N_5988,N_5054);
nand U6406 (N_6406,N_5935,N_5341);
nand U6407 (N_6407,N_5530,N_5903);
xnor U6408 (N_6408,N_5336,N_5982);
or U6409 (N_6409,N_5641,N_5662);
nand U6410 (N_6410,N_5200,N_5027);
nor U6411 (N_6411,N_5817,N_5598);
nand U6412 (N_6412,N_5401,N_5047);
nand U6413 (N_6413,N_5349,N_5602);
or U6414 (N_6414,N_5978,N_5558);
nand U6415 (N_6415,N_5382,N_5432);
nand U6416 (N_6416,N_5003,N_5660);
nor U6417 (N_6417,N_5939,N_5568);
or U6418 (N_6418,N_5993,N_5484);
or U6419 (N_6419,N_5158,N_5480);
nand U6420 (N_6420,N_5524,N_5278);
or U6421 (N_6421,N_5183,N_5997);
or U6422 (N_6422,N_5597,N_5743);
and U6423 (N_6423,N_5901,N_5213);
and U6424 (N_6424,N_5627,N_5905);
or U6425 (N_6425,N_5037,N_5394);
nand U6426 (N_6426,N_5734,N_5273);
nor U6427 (N_6427,N_5239,N_5282);
nand U6428 (N_6428,N_5767,N_5654);
nand U6429 (N_6429,N_5218,N_5547);
and U6430 (N_6430,N_5653,N_5055);
or U6431 (N_6431,N_5159,N_5395);
and U6432 (N_6432,N_5167,N_5344);
nand U6433 (N_6433,N_5911,N_5694);
and U6434 (N_6434,N_5087,N_5920);
or U6435 (N_6435,N_5124,N_5703);
xnor U6436 (N_6436,N_5091,N_5133);
nor U6437 (N_6437,N_5470,N_5069);
xor U6438 (N_6438,N_5067,N_5139);
nand U6439 (N_6439,N_5216,N_5093);
nand U6440 (N_6440,N_5895,N_5230);
or U6441 (N_6441,N_5094,N_5016);
nand U6442 (N_6442,N_5589,N_5818);
or U6443 (N_6443,N_5146,N_5117);
nor U6444 (N_6444,N_5421,N_5746);
nand U6445 (N_6445,N_5957,N_5140);
nand U6446 (N_6446,N_5402,N_5038);
nor U6447 (N_6447,N_5064,N_5805);
and U6448 (N_6448,N_5838,N_5643);
nand U6449 (N_6449,N_5309,N_5488);
nand U6450 (N_6450,N_5725,N_5727);
nand U6451 (N_6451,N_5321,N_5099);
nand U6452 (N_6452,N_5445,N_5672);
nand U6453 (N_6453,N_5059,N_5691);
nor U6454 (N_6454,N_5264,N_5756);
nand U6455 (N_6455,N_5561,N_5863);
nor U6456 (N_6456,N_5872,N_5074);
nor U6457 (N_6457,N_5246,N_5089);
nand U6458 (N_6458,N_5111,N_5215);
nand U6459 (N_6459,N_5806,N_5976);
nand U6460 (N_6460,N_5811,N_5025);
or U6461 (N_6461,N_5665,N_5129);
and U6462 (N_6462,N_5919,N_5307);
and U6463 (N_6463,N_5721,N_5917);
nand U6464 (N_6464,N_5803,N_5652);
and U6465 (N_6465,N_5866,N_5483);
nand U6466 (N_6466,N_5008,N_5511);
nand U6467 (N_6467,N_5715,N_5306);
or U6468 (N_6468,N_5078,N_5433);
nor U6469 (N_6469,N_5772,N_5226);
or U6470 (N_6470,N_5884,N_5629);
nand U6471 (N_6471,N_5954,N_5773);
nor U6472 (N_6472,N_5689,N_5934);
and U6473 (N_6473,N_5203,N_5955);
nor U6474 (N_6474,N_5536,N_5443);
and U6475 (N_6475,N_5162,N_5191);
and U6476 (N_6476,N_5143,N_5626);
and U6477 (N_6477,N_5632,N_5290);
xnor U6478 (N_6478,N_5329,N_5022);
nand U6479 (N_6479,N_5267,N_5346);
and U6480 (N_6480,N_5326,N_5754);
nand U6481 (N_6481,N_5902,N_5429);
nor U6482 (N_6482,N_5137,N_5690);
and U6483 (N_6483,N_5333,N_5608);
nor U6484 (N_6484,N_5368,N_5023);
or U6485 (N_6485,N_5636,N_5322);
nand U6486 (N_6486,N_5814,N_5700);
and U6487 (N_6487,N_5096,N_5953);
nand U6488 (N_6488,N_5788,N_5453);
nand U6489 (N_6489,N_5816,N_5910);
nor U6490 (N_6490,N_5284,N_5506);
or U6491 (N_6491,N_5543,N_5185);
nand U6492 (N_6492,N_5263,N_5924);
nor U6493 (N_6493,N_5328,N_5687);
or U6494 (N_6494,N_5728,N_5490);
or U6495 (N_6495,N_5496,N_5844);
xor U6496 (N_6496,N_5131,N_5979);
nor U6497 (N_6497,N_5130,N_5996);
xor U6498 (N_6498,N_5224,N_5802);
nor U6499 (N_6499,N_5194,N_5942);
or U6500 (N_6500,N_5470,N_5671);
nor U6501 (N_6501,N_5355,N_5024);
and U6502 (N_6502,N_5529,N_5054);
nor U6503 (N_6503,N_5404,N_5161);
nand U6504 (N_6504,N_5302,N_5746);
nand U6505 (N_6505,N_5344,N_5662);
and U6506 (N_6506,N_5341,N_5187);
xor U6507 (N_6507,N_5322,N_5022);
and U6508 (N_6508,N_5835,N_5613);
nor U6509 (N_6509,N_5649,N_5669);
nor U6510 (N_6510,N_5280,N_5023);
xor U6511 (N_6511,N_5805,N_5021);
and U6512 (N_6512,N_5997,N_5484);
and U6513 (N_6513,N_5858,N_5130);
or U6514 (N_6514,N_5299,N_5896);
nand U6515 (N_6515,N_5277,N_5403);
nor U6516 (N_6516,N_5768,N_5702);
nor U6517 (N_6517,N_5088,N_5596);
or U6518 (N_6518,N_5434,N_5953);
nor U6519 (N_6519,N_5915,N_5510);
xor U6520 (N_6520,N_5249,N_5080);
nand U6521 (N_6521,N_5421,N_5553);
or U6522 (N_6522,N_5085,N_5230);
or U6523 (N_6523,N_5813,N_5309);
nor U6524 (N_6524,N_5611,N_5431);
nand U6525 (N_6525,N_5724,N_5741);
nor U6526 (N_6526,N_5698,N_5222);
nor U6527 (N_6527,N_5651,N_5953);
or U6528 (N_6528,N_5927,N_5882);
and U6529 (N_6529,N_5518,N_5358);
and U6530 (N_6530,N_5099,N_5372);
and U6531 (N_6531,N_5689,N_5406);
nor U6532 (N_6532,N_5018,N_5336);
nor U6533 (N_6533,N_5069,N_5459);
or U6534 (N_6534,N_5343,N_5486);
and U6535 (N_6535,N_5027,N_5212);
nor U6536 (N_6536,N_5179,N_5308);
nor U6537 (N_6537,N_5828,N_5559);
or U6538 (N_6538,N_5898,N_5575);
xor U6539 (N_6539,N_5206,N_5840);
xor U6540 (N_6540,N_5061,N_5932);
nand U6541 (N_6541,N_5645,N_5556);
nor U6542 (N_6542,N_5774,N_5679);
nor U6543 (N_6543,N_5075,N_5206);
nand U6544 (N_6544,N_5404,N_5846);
nor U6545 (N_6545,N_5943,N_5347);
and U6546 (N_6546,N_5331,N_5815);
or U6547 (N_6547,N_5801,N_5408);
and U6548 (N_6548,N_5258,N_5175);
or U6549 (N_6549,N_5732,N_5828);
nand U6550 (N_6550,N_5935,N_5636);
nor U6551 (N_6551,N_5872,N_5459);
nor U6552 (N_6552,N_5937,N_5179);
nor U6553 (N_6553,N_5884,N_5944);
or U6554 (N_6554,N_5019,N_5955);
or U6555 (N_6555,N_5115,N_5486);
nand U6556 (N_6556,N_5722,N_5682);
and U6557 (N_6557,N_5665,N_5989);
nor U6558 (N_6558,N_5509,N_5253);
nor U6559 (N_6559,N_5980,N_5714);
and U6560 (N_6560,N_5740,N_5295);
nor U6561 (N_6561,N_5288,N_5294);
and U6562 (N_6562,N_5908,N_5295);
nand U6563 (N_6563,N_5759,N_5564);
xor U6564 (N_6564,N_5762,N_5642);
and U6565 (N_6565,N_5878,N_5968);
nor U6566 (N_6566,N_5825,N_5618);
and U6567 (N_6567,N_5982,N_5055);
and U6568 (N_6568,N_5616,N_5563);
nor U6569 (N_6569,N_5142,N_5689);
xnor U6570 (N_6570,N_5991,N_5216);
and U6571 (N_6571,N_5184,N_5373);
or U6572 (N_6572,N_5064,N_5463);
and U6573 (N_6573,N_5321,N_5938);
nand U6574 (N_6574,N_5315,N_5688);
nand U6575 (N_6575,N_5889,N_5987);
and U6576 (N_6576,N_5073,N_5933);
or U6577 (N_6577,N_5652,N_5867);
and U6578 (N_6578,N_5149,N_5139);
and U6579 (N_6579,N_5982,N_5881);
or U6580 (N_6580,N_5635,N_5845);
nand U6581 (N_6581,N_5783,N_5594);
nor U6582 (N_6582,N_5397,N_5249);
nor U6583 (N_6583,N_5331,N_5854);
nand U6584 (N_6584,N_5591,N_5101);
nand U6585 (N_6585,N_5987,N_5236);
or U6586 (N_6586,N_5134,N_5486);
nand U6587 (N_6587,N_5938,N_5579);
nor U6588 (N_6588,N_5104,N_5016);
or U6589 (N_6589,N_5808,N_5889);
or U6590 (N_6590,N_5014,N_5470);
and U6591 (N_6591,N_5092,N_5922);
nor U6592 (N_6592,N_5239,N_5948);
and U6593 (N_6593,N_5926,N_5100);
nand U6594 (N_6594,N_5757,N_5675);
xor U6595 (N_6595,N_5709,N_5312);
or U6596 (N_6596,N_5846,N_5996);
nand U6597 (N_6597,N_5735,N_5420);
or U6598 (N_6598,N_5358,N_5499);
nand U6599 (N_6599,N_5446,N_5823);
nor U6600 (N_6600,N_5898,N_5651);
and U6601 (N_6601,N_5854,N_5343);
or U6602 (N_6602,N_5620,N_5043);
xnor U6603 (N_6603,N_5877,N_5035);
or U6604 (N_6604,N_5785,N_5272);
nand U6605 (N_6605,N_5939,N_5406);
or U6606 (N_6606,N_5064,N_5902);
and U6607 (N_6607,N_5705,N_5274);
and U6608 (N_6608,N_5175,N_5319);
nand U6609 (N_6609,N_5063,N_5974);
and U6610 (N_6610,N_5223,N_5626);
nand U6611 (N_6611,N_5640,N_5150);
or U6612 (N_6612,N_5907,N_5066);
nor U6613 (N_6613,N_5189,N_5222);
nor U6614 (N_6614,N_5067,N_5200);
or U6615 (N_6615,N_5709,N_5340);
nor U6616 (N_6616,N_5904,N_5481);
and U6617 (N_6617,N_5725,N_5821);
nand U6618 (N_6618,N_5654,N_5389);
nor U6619 (N_6619,N_5117,N_5088);
and U6620 (N_6620,N_5710,N_5475);
and U6621 (N_6621,N_5279,N_5617);
nand U6622 (N_6622,N_5132,N_5492);
and U6623 (N_6623,N_5844,N_5219);
nand U6624 (N_6624,N_5683,N_5329);
nor U6625 (N_6625,N_5972,N_5534);
xnor U6626 (N_6626,N_5128,N_5034);
nand U6627 (N_6627,N_5350,N_5944);
or U6628 (N_6628,N_5368,N_5963);
or U6629 (N_6629,N_5819,N_5014);
and U6630 (N_6630,N_5240,N_5006);
and U6631 (N_6631,N_5124,N_5548);
nand U6632 (N_6632,N_5772,N_5249);
nor U6633 (N_6633,N_5681,N_5621);
and U6634 (N_6634,N_5908,N_5964);
nor U6635 (N_6635,N_5947,N_5249);
and U6636 (N_6636,N_5873,N_5326);
xor U6637 (N_6637,N_5805,N_5167);
nor U6638 (N_6638,N_5370,N_5567);
xnor U6639 (N_6639,N_5113,N_5052);
nand U6640 (N_6640,N_5103,N_5648);
or U6641 (N_6641,N_5203,N_5017);
and U6642 (N_6642,N_5518,N_5996);
nand U6643 (N_6643,N_5706,N_5423);
or U6644 (N_6644,N_5140,N_5432);
or U6645 (N_6645,N_5668,N_5842);
or U6646 (N_6646,N_5163,N_5251);
and U6647 (N_6647,N_5770,N_5111);
or U6648 (N_6648,N_5126,N_5884);
or U6649 (N_6649,N_5943,N_5307);
or U6650 (N_6650,N_5380,N_5343);
nand U6651 (N_6651,N_5099,N_5019);
or U6652 (N_6652,N_5153,N_5345);
or U6653 (N_6653,N_5528,N_5654);
xnor U6654 (N_6654,N_5439,N_5191);
or U6655 (N_6655,N_5423,N_5237);
xnor U6656 (N_6656,N_5917,N_5504);
xnor U6657 (N_6657,N_5798,N_5473);
nand U6658 (N_6658,N_5792,N_5970);
and U6659 (N_6659,N_5865,N_5329);
or U6660 (N_6660,N_5555,N_5711);
and U6661 (N_6661,N_5411,N_5801);
or U6662 (N_6662,N_5862,N_5584);
nand U6663 (N_6663,N_5295,N_5464);
or U6664 (N_6664,N_5128,N_5151);
or U6665 (N_6665,N_5929,N_5763);
or U6666 (N_6666,N_5412,N_5575);
or U6667 (N_6667,N_5214,N_5969);
nor U6668 (N_6668,N_5404,N_5416);
nor U6669 (N_6669,N_5270,N_5985);
nor U6670 (N_6670,N_5053,N_5816);
nand U6671 (N_6671,N_5294,N_5109);
or U6672 (N_6672,N_5703,N_5348);
and U6673 (N_6673,N_5913,N_5267);
and U6674 (N_6674,N_5011,N_5214);
nand U6675 (N_6675,N_5457,N_5891);
or U6676 (N_6676,N_5909,N_5238);
nand U6677 (N_6677,N_5171,N_5296);
nor U6678 (N_6678,N_5242,N_5559);
or U6679 (N_6679,N_5519,N_5914);
nor U6680 (N_6680,N_5624,N_5546);
nand U6681 (N_6681,N_5453,N_5032);
or U6682 (N_6682,N_5876,N_5999);
nor U6683 (N_6683,N_5815,N_5738);
and U6684 (N_6684,N_5110,N_5439);
nor U6685 (N_6685,N_5438,N_5844);
nor U6686 (N_6686,N_5425,N_5526);
nor U6687 (N_6687,N_5414,N_5834);
nand U6688 (N_6688,N_5449,N_5178);
nor U6689 (N_6689,N_5087,N_5164);
nand U6690 (N_6690,N_5337,N_5194);
nor U6691 (N_6691,N_5149,N_5635);
and U6692 (N_6692,N_5519,N_5032);
nor U6693 (N_6693,N_5997,N_5260);
and U6694 (N_6694,N_5908,N_5235);
nand U6695 (N_6695,N_5241,N_5799);
nor U6696 (N_6696,N_5204,N_5693);
nand U6697 (N_6697,N_5441,N_5283);
or U6698 (N_6698,N_5306,N_5599);
nand U6699 (N_6699,N_5210,N_5075);
nor U6700 (N_6700,N_5192,N_5775);
nand U6701 (N_6701,N_5808,N_5717);
nand U6702 (N_6702,N_5020,N_5840);
nor U6703 (N_6703,N_5142,N_5991);
and U6704 (N_6704,N_5687,N_5325);
and U6705 (N_6705,N_5625,N_5058);
or U6706 (N_6706,N_5199,N_5507);
or U6707 (N_6707,N_5649,N_5850);
nand U6708 (N_6708,N_5817,N_5878);
nand U6709 (N_6709,N_5116,N_5134);
nand U6710 (N_6710,N_5537,N_5255);
nand U6711 (N_6711,N_5014,N_5659);
xnor U6712 (N_6712,N_5975,N_5905);
or U6713 (N_6713,N_5706,N_5173);
and U6714 (N_6714,N_5026,N_5012);
nand U6715 (N_6715,N_5831,N_5295);
and U6716 (N_6716,N_5848,N_5010);
nand U6717 (N_6717,N_5961,N_5386);
and U6718 (N_6718,N_5915,N_5518);
nor U6719 (N_6719,N_5884,N_5280);
nor U6720 (N_6720,N_5270,N_5529);
or U6721 (N_6721,N_5881,N_5986);
nor U6722 (N_6722,N_5695,N_5489);
and U6723 (N_6723,N_5443,N_5722);
and U6724 (N_6724,N_5973,N_5751);
nand U6725 (N_6725,N_5151,N_5085);
nor U6726 (N_6726,N_5985,N_5128);
nor U6727 (N_6727,N_5345,N_5298);
and U6728 (N_6728,N_5253,N_5413);
and U6729 (N_6729,N_5413,N_5158);
xor U6730 (N_6730,N_5348,N_5910);
or U6731 (N_6731,N_5864,N_5345);
and U6732 (N_6732,N_5650,N_5733);
nor U6733 (N_6733,N_5875,N_5412);
nor U6734 (N_6734,N_5158,N_5947);
xor U6735 (N_6735,N_5042,N_5784);
and U6736 (N_6736,N_5595,N_5836);
or U6737 (N_6737,N_5186,N_5366);
and U6738 (N_6738,N_5965,N_5806);
and U6739 (N_6739,N_5153,N_5026);
nor U6740 (N_6740,N_5813,N_5160);
and U6741 (N_6741,N_5755,N_5756);
or U6742 (N_6742,N_5867,N_5088);
nor U6743 (N_6743,N_5484,N_5463);
and U6744 (N_6744,N_5435,N_5764);
or U6745 (N_6745,N_5924,N_5136);
nor U6746 (N_6746,N_5290,N_5723);
nor U6747 (N_6747,N_5121,N_5029);
and U6748 (N_6748,N_5343,N_5304);
nor U6749 (N_6749,N_5324,N_5906);
nand U6750 (N_6750,N_5178,N_5498);
nand U6751 (N_6751,N_5927,N_5140);
nor U6752 (N_6752,N_5712,N_5715);
nand U6753 (N_6753,N_5876,N_5296);
or U6754 (N_6754,N_5521,N_5792);
nor U6755 (N_6755,N_5144,N_5234);
or U6756 (N_6756,N_5840,N_5507);
and U6757 (N_6757,N_5301,N_5265);
xor U6758 (N_6758,N_5882,N_5803);
xor U6759 (N_6759,N_5021,N_5125);
or U6760 (N_6760,N_5260,N_5748);
and U6761 (N_6761,N_5061,N_5596);
and U6762 (N_6762,N_5037,N_5645);
nor U6763 (N_6763,N_5887,N_5399);
or U6764 (N_6764,N_5468,N_5241);
nand U6765 (N_6765,N_5425,N_5636);
nor U6766 (N_6766,N_5146,N_5443);
and U6767 (N_6767,N_5507,N_5012);
or U6768 (N_6768,N_5669,N_5284);
nor U6769 (N_6769,N_5733,N_5455);
nand U6770 (N_6770,N_5149,N_5171);
nand U6771 (N_6771,N_5034,N_5661);
nor U6772 (N_6772,N_5121,N_5814);
or U6773 (N_6773,N_5627,N_5648);
and U6774 (N_6774,N_5811,N_5238);
nand U6775 (N_6775,N_5266,N_5443);
or U6776 (N_6776,N_5677,N_5328);
nand U6777 (N_6777,N_5678,N_5490);
or U6778 (N_6778,N_5599,N_5631);
nand U6779 (N_6779,N_5388,N_5922);
nor U6780 (N_6780,N_5360,N_5378);
nor U6781 (N_6781,N_5915,N_5536);
and U6782 (N_6782,N_5230,N_5108);
and U6783 (N_6783,N_5493,N_5266);
nor U6784 (N_6784,N_5180,N_5991);
nor U6785 (N_6785,N_5678,N_5976);
nand U6786 (N_6786,N_5492,N_5180);
nor U6787 (N_6787,N_5556,N_5633);
nor U6788 (N_6788,N_5038,N_5291);
nor U6789 (N_6789,N_5174,N_5241);
and U6790 (N_6790,N_5430,N_5680);
and U6791 (N_6791,N_5234,N_5448);
nand U6792 (N_6792,N_5101,N_5361);
and U6793 (N_6793,N_5292,N_5987);
or U6794 (N_6794,N_5458,N_5075);
nor U6795 (N_6795,N_5551,N_5301);
or U6796 (N_6796,N_5340,N_5850);
nand U6797 (N_6797,N_5465,N_5368);
nand U6798 (N_6798,N_5594,N_5192);
or U6799 (N_6799,N_5159,N_5022);
nor U6800 (N_6800,N_5037,N_5287);
xor U6801 (N_6801,N_5867,N_5222);
nor U6802 (N_6802,N_5483,N_5399);
nor U6803 (N_6803,N_5370,N_5086);
nor U6804 (N_6804,N_5451,N_5817);
nor U6805 (N_6805,N_5720,N_5298);
nand U6806 (N_6806,N_5296,N_5365);
or U6807 (N_6807,N_5313,N_5519);
and U6808 (N_6808,N_5003,N_5797);
and U6809 (N_6809,N_5353,N_5006);
or U6810 (N_6810,N_5648,N_5706);
nand U6811 (N_6811,N_5067,N_5934);
and U6812 (N_6812,N_5935,N_5450);
nand U6813 (N_6813,N_5130,N_5762);
and U6814 (N_6814,N_5623,N_5665);
or U6815 (N_6815,N_5855,N_5236);
nand U6816 (N_6816,N_5042,N_5928);
and U6817 (N_6817,N_5903,N_5370);
nand U6818 (N_6818,N_5711,N_5903);
nor U6819 (N_6819,N_5541,N_5897);
or U6820 (N_6820,N_5851,N_5017);
nor U6821 (N_6821,N_5417,N_5437);
or U6822 (N_6822,N_5792,N_5225);
or U6823 (N_6823,N_5513,N_5990);
nand U6824 (N_6824,N_5317,N_5568);
nand U6825 (N_6825,N_5826,N_5871);
nand U6826 (N_6826,N_5863,N_5472);
and U6827 (N_6827,N_5243,N_5361);
or U6828 (N_6828,N_5472,N_5226);
nor U6829 (N_6829,N_5137,N_5822);
and U6830 (N_6830,N_5080,N_5070);
nor U6831 (N_6831,N_5306,N_5913);
nand U6832 (N_6832,N_5953,N_5545);
or U6833 (N_6833,N_5226,N_5738);
nand U6834 (N_6834,N_5554,N_5437);
or U6835 (N_6835,N_5962,N_5145);
nor U6836 (N_6836,N_5685,N_5787);
or U6837 (N_6837,N_5602,N_5823);
nor U6838 (N_6838,N_5806,N_5121);
nor U6839 (N_6839,N_5067,N_5540);
nor U6840 (N_6840,N_5035,N_5375);
nor U6841 (N_6841,N_5356,N_5713);
and U6842 (N_6842,N_5690,N_5232);
and U6843 (N_6843,N_5312,N_5732);
or U6844 (N_6844,N_5721,N_5577);
nand U6845 (N_6845,N_5750,N_5647);
or U6846 (N_6846,N_5483,N_5487);
or U6847 (N_6847,N_5712,N_5029);
or U6848 (N_6848,N_5475,N_5084);
nor U6849 (N_6849,N_5547,N_5708);
nor U6850 (N_6850,N_5361,N_5393);
nor U6851 (N_6851,N_5234,N_5830);
nor U6852 (N_6852,N_5462,N_5003);
or U6853 (N_6853,N_5305,N_5534);
and U6854 (N_6854,N_5097,N_5012);
or U6855 (N_6855,N_5303,N_5024);
nand U6856 (N_6856,N_5386,N_5949);
nand U6857 (N_6857,N_5413,N_5606);
and U6858 (N_6858,N_5059,N_5338);
nand U6859 (N_6859,N_5561,N_5577);
nor U6860 (N_6860,N_5824,N_5743);
nand U6861 (N_6861,N_5726,N_5508);
or U6862 (N_6862,N_5299,N_5889);
and U6863 (N_6863,N_5727,N_5526);
nand U6864 (N_6864,N_5030,N_5452);
or U6865 (N_6865,N_5359,N_5875);
and U6866 (N_6866,N_5063,N_5719);
nor U6867 (N_6867,N_5882,N_5633);
nor U6868 (N_6868,N_5853,N_5368);
nor U6869 (N_6869,N_5987,N_5183);
nor U6870 (N_6870,N_5392,N_5232);
and U6871 (N_6871,N_5514,N_5356);
nor U6872 (N_6872,N_5282,N_5215);
and U6873 (N_6873,N_5112,N_5061);
or U6874 (N_6874,N_5068,N_5361);
or U6875 (N_6875,N_5003,N_5638);
and U6876 (N_6876,N_5951,N_5533);
nand U6877 (N_6877,N_5954,N_5513);
nand U6878 (N_6878,N_5688,N_5173);
or U6879 (N_6879,N_5500,N_5382);
nor U6880 (N_6880,N_5156,N_5698);
nand U6881 (N_6881,N_5748,N_5469);
or U6882 (N_6882,N_5523,N_5893);
and U6883 (N_6883,N_5707,N_5922);
xnor U6884 (N_6884,N_5728,N_5112);
nand U6885 (N_6885,N_5433,N_5917);
nand U6886 (N_6886,N_5238,N_5202);
nand U6887 (N_6887,N_5385,N_5038);
and U6888 (N_6888,N_5747,N_5346);
nand U6889 (N_6889,N_5219,N_5990);
nand U6890 (N_6890,N_5161,N_5857);
nor U6891 (N_6891,N_5923,N_5846);
or U6892 (N_6892,N_5235,N_5387);
or U6893 (N_6893,N_5796,N_5916);
nand U6894 (N_6894,N_5967,N_5249);
nor U6895 (N_6895,N_5161,N_5298);
nor U6896 (N_6896,N_5126,N_5220);
nor U6897 (N_6897,N_5778,N_5355);
nand U6898 (N_6898,N_5325,N_5256);
and U6899 (N_6899,N_5817,N_5806);
nand U6900 (N_6900,N_5195,N_5300);
nor U6901 (N_6901,N_5442,N_5697);
or U6902 (N_6902,N_5216,N_5309);
and U6903 (N_6903,N_5307,N_5455);
nand U6904 (N_6904,N_5725,N_5578);
nand U6905 (N_6905,N_5516,N_5996);
or U6906 (N_6906,N_5434,N_5280);
or U6907 (N_6907,N_5999,N_5774);
and U6908 (N_6908,N_5452,N_5488);
xnor U6909 (N_6909,N_5734,N_5348);
nor U6910 (N_6910,N_5405,N_5639);
or U6911 (N_6911,N_5740,N_5621);
and U6912 (N_6912,N_5240,N_5331);
nand U6913 (N_6913,N_5999,N_5797);
and U6914 (N_6914,N_5780,N_5589);
or U6915 (N_6915,N_5998,N_5286);
or U6916 (N_6916,N_5603,N_5492);
and U6917 (N_6917,N_5632,N_5335);
nand U6918 (N_6918,N_5749,N_5501);
nand U6919 (N_6919,N_5837,N_5072);
or U6920 (N_6920,N_5031,N_5690);
and U6921 (N_6921,N_5001,N_5068);
and U6922 (N_6922,N_5055,N_5850);
or U6923 (N_6923,N_5082,N_5217);
nand U6924 (N_6924,N_5805,N_5037);
and U6925 (N_6925,N_5920,N_5658);
nand U6926 (N_6926,N_5135,N_5126);
nand U6927 (N_6927,N_5891,N_5241);
nor U6928 (N_6928,N_5990,N_5392);
nor U6929 (N_6929,N_5171,N_5497);
and U6930 (N_6930,N_5617,N_5517);
nand U6931 (N_6931,N_5778,N_5444);
and U6932 (N_6932,N_5571,N_5146);
nand U6933 (N_6933,N_5011,N_5019);
nand U6934 (N_6934,N_5490,N_5053);
nand U6935 (N_6935,N_5244,N_5184);
nor U6936 (N_6936,N_5524,N_5282);
or U6937 (N_6937,N_5438,N_5828);
nand U6938 (N_6938,N_5881,N_5534);
nand U6939 (N_6939,N_5466,N_5644);
nand U6940 (N_6940,N_5158,N_5018);
nand U6941 (N_6941,N_5226,N_5834);
nand U6942 (N_6942,N_5698,N_5270);
nand U6943 (N_6943,N_5103,N_5847);
nand U6944 (N_6944,N_5612,N_5279);
nand U6945 (N_6945,N_5898,N_5772);
nor U6946 (N_6946,N_5058,N_5490);
nor U6947 (N_6947,N_5129,N_5379);
nand U6948 (N_6948,N_5367,N_5101);
or U6949 (N_6949,N_5181,N_5534);
nand U6950 (N_6950,N_5599,N_5690);
or U6951 (N_6951,N_5849,N_5597);
and U6952 (N_6952,N_5195,N_5402);
or U6953 (N_6953,N_5604,N_5804);
and U6954 (N_6954,N_5914,N_5963);
and U6955 (N_6955,N_5110,N_5915);
nor U6956 (N_6956,N_5219,N_5788);
and U6957 (N_6957,N_5492,N_5672);
or U6958 (N_6958,N_5810,N_5554);
or U6959 (N_6959,N_5849,N_5851);
nor U6960 (N_6960,N_5295,N_5352);
nor U6961 (N_6961,N_5285,N_5110);
nor U6962 (N_6962,N_5711,N_5197);
and U6963 (N_6963,N_5997,N_5441);
nor U6964 (N_6964,N_5815,N_5783);
nor U6965 (N_6965,N_5825,N_5233);
nor U6966 (N_6966,N_5004,N_5532);
or U6967 (N_6967,N_5671,N_5572);
nor U6968 (N_6968,N_5745,N_5741);
or U6969 (N_6969,N_5810,N_5747);
nand U6970 (N_6970,N_5790,N_5876);
nor U6971 (N_6971,N_5884,N_5623);
or U6972 (N_6972,N_5149,N_5488);
or U6973 (N_6973,N_5832,N_5862);
nand U6974 (N_6974,N_5117,N_5462);
nand U6975 (N_6975,N_5644,N_5164);
nand U6976 (N_6976,N_5541,N_5497);
xnor U6977 (N_6977,N_5712,N_5613);
nand U6978 (N_6978,N_5716,N_5827);
and U6979 (N_6979,N_5367,N_5264);
and U6980 (N_6980,N_5689,N_5354);
and U6981 (N_6981,N_5252,N_5432);
or U6982 (N_6982,N_5876,N_5177);
nor U6983 (N_6983,N_5512,N_5859);
or U6984 (N_6984,N_5158,N_5422);
nor U6985 (N_6985,N_5465,N_5170);
or U6986 (N_6986,N_5110,N_5581);
nor U6987 (N_6987,N_5780,N_5250);
and U6988 (N_6988,N_5431,N_5652);
or U6989 (N_6989,N_5709,N_5765);
or U6990 (N_6990,N_5231,N_5839);
nand U6991 (N_6991,N_5699,N_5375);
and U6992 (N_6992,N_5092,N_5388);
or U6993 (N_6993,N_5990,N_5590);
or U6994 (N_6994,N_5362,N_5501);
and U6995 (N_6995,N_5111,N_5912);
or U6996 (N_6996,N_5286,N_5659);
nor U6997 (N_6997,N_5416,N_5127);
nor U6998 (N_6998,N_5940,N_5252);
nand U6999 (N_6999,N_5645,N_5099);
nor U7000 (N_7000,N_6763,N_6988);
and U7001 (N_7001,N_6286,N_6245);
and U7002 (N_7002,N_6063,N_6880);
and U7003 (N_7003,N_6761,N_6142);
nor U7004 (N_7004,N_6876,N_6923);
nor U7005 (N_7005,N_6412,N_6180);
and U7006 (N_7006,N_6048,N_6429);
and U7007 (N_7007,N_6592,N_6331);
and U7008 (N_7008,N_6096,N_6773);
xnor U7009 (N_7009,N_6453,N_6261);
nor U7010 (N_7010,N_6955,N_6571);
nand U7011 (N_7011,N_6706,N_6410);
or U7012 (N_7012,N_6863,N_6817);
or U7013 (N_7013,N_6242,N_6626);
nor U7014 (N_7014,N_6846,N_6864);
or U7015 (N_7015,N_6290,N_6100);
or U7016 (N_7016,N_6523,N_6591);
or U7017 (N_7017,N_6214,N_6499);
and U7018 (N_7018,N_6418,N_6255);
nor U7019 (N_7019,N_6752,N_6918);
nand U7020 (N_7020,N_6220,N_6833);
xor U7021 (N_7021,N_6073,N_6606);
and U7022 (N_7022,N_6145,N_6685);
and U7023 (N_7023,N_6692,N_6722);
and U7024 (N_7024,N_6912,N_6733);
nor U7025 (N_7025,N_6162,N_6550);
nor U7026 (N_7026,N_6960,N_6598);
nor U7027 (N_7027,N_6356,N_6901);
nand U7028 (N_7028,N_6350,N_6460);
and U7029 (N_7029,N_6679,N_6738);
nor U7030 (N_7030,N_6989,N_6485);
and U7031 (N_7031,N_6602,N_6470);
nor U7032 (N_7032,N_6294,N_6518);
and U7033 (N_7033,N_6888,N_6737);
nand U7034 (N_7034,N_6328,N_6446);
nand U7035 (N_7035,N_6316,N_6312);
nand U7036 (N_7036,N_6040,N_6428);
or U7037 (N_7037,N_6198,N_6249);
or U7038 (N_7038,N_6366,N_6292);
or U7039 (N_7039,N_6395,N_6781);
and U7040 (N_7040,N_6502,N_6925);
nor U7041 (N_7041,N_6820,N_6108);
and U7042 (N_7042,N_6965,N_6035);
and U7043 (N_7043,N_6235,N_6767);
or U7044 (N_7044,N_6546,N_6802);
or U7045 (N_7045,N_6522,N_6194);
xor U7046 (N_7046,N_6101,N_6950);
or U7047 (N_7047,N_6060,N_6528);
or U7048 (N_7048,N_6259,N_6174);
and U7049 (N_7049,N_6822,N_6654);
nand U7050 (N_7050,N_6870,N_6910);
xnor U7051 (N_7051,N_6014,N_6646);
or U7052 (N_7052,N_6344,N_6951);
nor U7053 (N_7053,N_6199,N_6478);
nor U7054 (N_7054,N_6757,N_6287);
or U7055 (N_7055,N_6323,N_6452);
nand U7056 (N_7056,N_6547,N_6457);
nand U7057 (N_7057,N_6922,N_6930);
xor U7058 (N_7058,N_6791,N_6387);
nand U7059 (N_7059,N_6443,N_6610);
nor U7060 (N_7060,N_6620,N_6031);
nand U7061 (N_7061,N_6732,N_6437);
or U7062 (N_7062,N_6488,N_6309);
and U7063 (N_7063,N_6714,N_6021);
nor U7064 (N_7064,N_6717,N_6230);
nor U7065 (N_7065,N_6956,N_6560);
or U7066 (N_7066,N_6049,N_6422);
or U7067 (N_7067,N_6771,N_6223);
and U7068 (N_7068,N_6143,N_6374);
and U7069 (N_7069,N_6854,N_6621);
xnor U7070 (N_7070,N_6891,N_6744);
and U7071 (N_7071,N_6052,N_6419);
nor U7072 (N_7072,N_6203,N_6532);
or U7073 (N_7073,N_6128,N_6713);
and U7074 (N_7074,N_6015,N_6920);
or U7075 (N_7075,N_6293,N_6949);
nand U7076 (N_7076,N_6298,N_6787);
and U7077 (N_7077,N_6970,N_6897);
or U7078 (N_7078,N_6932,N_6961);
nand U7079 (N_7079,N_6990,N_6420);
nand U7080 (N_7080,N_6458,N_6144);
and U7081 (N_7081,N_6633,N_6436);
nor U7082 (N_7082,N_6608,N_6510);
nand U7083 (N_7083,N_6678,N_6012);
nor U7084 (N_7084,N_6303,N_6262);
nor U7085 (N_7085,N_6613,N_6110);
nor U7086 (N_7086,N_6728,N_6637);
or U7087 (N_7087,N_6931,N_6671);
and U7088 (N_7088,N_6795,N_6697);
nand U7089 (N_7089,N_6612,N_6302);
nor U7090 (N_7090,N_6946,N_6189);
nand U7091 (N_7091,N_6657,N_6830);
nand U7092 (N_7092,N_6248,N_6469);
or U7093 (N_7093,N_6721,N_6967);
nor U7094 (N_7094,N_6396,N_6579);
nor U7095 (N_7095,N_6667,N_6941);
and U7096 (N_7096,N_6739,N_6136);
nor U7097 (N_7097,N_6423,N_6115);
or U7098 (N_7098,N_6152,N_6158);
or U7099 (N_7099,N_6253,N_6719);
nor U7100 (N_7100,N_6688,N_6583);
and U7101 (N_7101,N_6748,N_6824);
nand U7102 (N_7102,N_6167,N_6804);
or U7103 (N_7103,N_6025,N_6276);
or U7104 (N_7104,N_6069,N_6887);
nand U7105 (N_7105,N_6630,N_6674);
nand U7106 (N_7106,N_6132,N_6206);
nor U7107 (N_7107,N_6789,N_6424);
or U7108 (N_7108,N_6801,N_6906);
nand U7109 (N_7109,N_6680,N_6165);
nand U7110 (N_7110,N_6736,N_6670);
and U7111 (N_7111,N_6994,N_6260);
nand U7112 (N_7112,N_6991,N_6465);
nand U7113 (N_7113,N_6102,N_6289);
xor U7114 (N_7114,N_6215,N_6002);
or U7115 (N_7115,N_6619,N_6234);
and U7116 (N_7116,N_6740,N_6053);
nand U7117 (N_7117,N_6020,N_6751);
and U7118 (N_7118,N_6477,N_6001);
or U7119 (N_7119,N_6588,N_6272);
and U7120 (N_7120,N_6668,N_6122);
xor U7121 (N_7121,N_6898,N_6508);
nor U7122 (N_7122,N_6027,N_6661);
or U7123 (N_7123,N_6828,N_6557);
nand U7124 (N_7124,N_6936,N_6154);
or U7125 (N_7125,N_6568,N_6482);
or U7126 (N_7126,N_6300,N_6120);
nand U7127 (N_7127,N_6202,N_6024);
or U7128 (N_7128,N_6584,N_6987);
nor U7129 (N_7129,N_6064,N_6785);
nand U7130 (N_7130,N_6777,N_6345);
or U7131 (N_7131,N_6903,N_6107);
nand U7132 (N_7132,N_6228,N_6690);
nand U7133 (N_7133,N_6765,N_6219);
nor U7134 (N_7134,N_6834,N_6582);
and U7135 (N_7135,N_6836,N_6501);
nand U7136 (N_7136,N_6747,N_6386);
nor U7137 (N_7137,N_6275,N_6217);
nand U7138 (N_7138,N_6258,N_6483);
xor U7139 (N_7139,N_6576,N_6393);
or U7140 (N_7140,N_6239,N_6947);
and U7141 (N_7141,N_6377,N_6317);
or U7142 (N_7142,N_6796,N_6288);
nand U7143 (N_7143,N_6181,N_6456);
nor U7144 (N_7144,N_6831,N_6811);
nor U7145 (N_7145,N_6384,N_6790);
or U7146 (N_7146,N_6558,N_6365);
xnor U7147 (N_7147,N_6225,N_6676);
nand U7148 (N_7148,N_6699,N_6195);
and U7149 (N_7149,N_6130,N_6640);
nand U7150 (N_7150,N_6911,N_6720);
xor U7151 (N_7151,N_6066,N_6611);
or U7152 (N_7152,N_6326,N_6121);
nor U7153 (N_7153,N_6004,N_6388);
and U7154 (N_7154,N_6807,N_6071);
nor U7155 (N_7155,N_6319,N_6570);
or U7156 (N_7156,N_6475,N_6937);
nand U7157 (N_7157,N_6335,N_6271);
or U7158 (N_7158,N_6940,N_6373);
nand U7159 (N_7159,N_6171,N_6754);
nand U7160 (N_7160,N_6094,N_6934);
and U7161 (N_7161,N_6809,N_6995);
nand U7162 (N_7162,N_6586,N_6694);
nor U7163 (N_7163,N_6869,N_6042);
nor U7164 (N_7164,N_6871,N_6684);
or U7165 (N_7165,N_6018,N_6352);
nand U7166 (N_7166,N_6417,N_6322);
and U7167 (N_7167,N_6603,N_6561);
nor U7168 (N_7168,N_6095,N_6074);
and U7169 (N_7169,N_6472,N_6686);
or U7170 (N_7170,N_6524,N_6845);
or U7171 (N_7171,N_6186,N_6484);
or U7172 (N_7172,N_6803,N_6779);
nand U7173 (N_7173,N_6404,N_6370);
and U7174 (N_7174,N_6541,N_6486);
nand U7175 (N_7175,N_6459,N_6118);
nand U7176 (N_7176,N_6858,N_6046);
nand U7177 (N_7177,N_6638,N_6026);
and U7178 (N_7178,N_6147,N_6116);
nand U7179 (N_7179,N_6361,N_6081);
nand U7180 (N_7180,N_6173,N_6474);
nand U7181 (N_7181,N_6496,N_6425);
nor U7182 (N_7182,N_6650,N_6376);
or U7183 (N_7183,N_6859,N_6448);
nand U7184 (N_7184,N_6498,N_6764);
nand U7185 (N_7185,N_6881,N_6939);
nor U7186 (N_7186,N_6749,N_6003);
nor U7187 (N_7187,N_6562,N_6051);
and U7188 (N_7188,N_6529,N_6282);
xor U7189 (N_7189,N_6839,N_6433);
or U7190 (N_7190,N_6503,N_6634);
and U7191 (N_7191,N_6770,N_6653);
nor U7192 (N_7192,N_6466,N_6392);
or U7193 (N_7193,N_6601,N_6954);
or U7194 (N_7194,N_6971,N_6758);
nand U7195 (N_7195,N_6264,N_6759);
and U7196 (N_7196,N_6281,N_6175);
and U7197 (N_7197,N_6237,N_6111);
nand U7198 (N_7198,N_6236,N_6375);
and U7199 (N_7199,N_6315,N_6605);
and U7200 (N_7200,N_6379,N_6170);
nor U7201 (N_7201,N_6882,N_6179);
nor U7202 (N_7202,N_6567,N_6982);
nand U7203 (N_7203,N_6246,N_6251);
or U7204 (N_7204,N_6127,N_6389);
nand U7205 (N_7205,N_6663,N_6092);
and U7206 (N_7206,N_6347,N_6016);
or U7207 (N_7207,N_6059,N_6408);
nand U7208 (N_7208,N_6163,N_6900);
xor U7209 (N_7209,N_6964,N_6993);
nand U7210 (N_7210,N_6036,N_6378);
nor U7211 (N_7211,N_6124,N_6471);
nor U7212 (N_7212,N_6409,N_6691);
nand U7213 (N_7213,N_6886,N_6543);
nand U7214 (N_7214,N_6509,N_6193);
nand U7215 (N_7215,N_6278,N_6357);
or U7216 (N_7216,N_6464,N_6873);
nand U7217 (N_7217,N_6097,N_6868);
nor U7218 (N_7218,N_6844,N_6957);
nor U7219 (N_7219,N_6243,N_6599);
nor U7220 (N_7220,N_6829,N_6632);
nand U7221 (N_7221,N_6521,N_6683);
nand U7222 (N_7222,N_6105,N_6700);
nand U7223 (N_7223,N_6310,N_6734);
and U7224 (N_7224,N_6559,N_6304);
nor U7225 (N_7225,N_6526,N_6150);
or U7226 (N_7226,N_6673,N_6123);
nor U7227 (N_7227,N_6682,N_6256);
and U7228 (N_7228,N_6977,N_6702);
or U7229 (N_7229,N_6642,N_6782);
nand U7230 (N_7230,N_6889,N_6695);
or U7231 (N_7231,N_6197,N_6953);
and U7232 (N_7232,N_6712,N_6454);
xnor U7233 (N_7233,N_6119,N_6774);
nor U7234 (N_7234,N_6535,N_6390);
and U7235 (N_7235,N_6070,N_6826);
nor U7236 (N_7236,N_6212,N_6134);
nor U7237 (N_7237,N_6821,N_6400);
or U7238 (N_7238,N_6841,N_6735);
or U7239 (N_7239,N_6226,N_6628);
nand U7240 (N_7240,N_6146,N_6159);
nor U7241 (N_7241,N_6835,N_6011);
or U7242 (N_7242,N_6086,N_6346);
nor U7243 (N_7243,N_6468,N_6382);
and U7244 (N_7244,N_6072,N_6615);
nand U7245 (N_7245,N_6183,N_6296);
or U7246 (N_7246,N_6681,N_6114);
nor U7247 (N_7247,N_6495,N_6339);
or U7248 (N_7248,N_6704,N_6353);
or U7249 (N_7249,N_6609,N_6851);
nand U7250 (N_7250,N_6155,N_6233);
nor U7251 (N_7251,N_6455,N_6489);
nor U7252 (N_7252,N_6277,N_6336);
nor U7253 (N_7253,N_6385,N_6330);
or U7254 (N_7254,N_6872,N_6103);
nor U7255 (N_7255,N_6861,N_6444);
nand U7256 (N_7256,N_6525,N_6113);
nor U7257 (N_7257,N_6625,N_6693);
nand U7258 (N_7258,N_6211,N_6314);
xnor U7259 (N_7259,N_6698,N_6087);
or U7260 (N_7260,N_6311,N_6263);
and U7261 (N_7261,N_6088,N_6805);
nand U7262 (N_7262,N_6921,N_6877);
nand U7263 (N_7263,N_6125,N_6224);
and U7264 (N_7264,N_6677,N_6649);
nor U7265 (N_7265,N_6769,N_6825);
xnor U7266 (N_7266,N_6656,N_6966);
nor U7267 (N_7267,N_6729,N_6098);
and U7268 (N_7268,N_6574,N_6614);
nor U7269 (N_7269,N_6666,N_6527);
nand U7270 (N_7270,N_6129,N_6435);
nand U7271 (N_7271,N_6112,N_6209);
and U7272 (N_7272,N_6952,N_6624);
and U7273 (N_7273,N_6916,N_6847);
and U7274 (N_7274,N_6270,N_6082);
nand U7275 (N_7275,N_6157,N_6291);
and U7276 (N_7276,N_6449,N_6655);
nor U7277 (N_7277,N_6514,N_6711);
and U7278 (N_7278,N_6280,N_6553);
and U7279 (N_7279,N_6549,N_6265);
nor U7280 (N_7280,N_6492,N_6138);
or U7281 (N_7281,N_6305,N_6324);
xor U7282 (N_7282,N_6511,N_6430);
nand U7283 (N_7283,N_6061,N_6569);
nor U7284 (N_7284,N_6089,N_6504);
nand U7285 (N_7285,N_6427,N_6505);
and U7286 (N_7286,N_6581,N_6044);
and U7287 (N_7287,N_6359,N_6340);
or U7288 (N_7288,N_6268,N_6516);
or U7289 (N_7289,N_6369,N_6078);
nor U7290 (N_7290,N_6812,N_6057);
nor U7291 (N_7291,N_6329,N_6832);
nand U7292 (N_7292,N_6651,N_6038);
nor U7293 (N_7293,N_6766,N_6141);
or U7294 (N_7294,N_6421,N_6867);
nand U7295 (N_7295,N_6325,N_6857);
nor U7296 (N_7296,N_6659,N_6076);
or U7297 (N_7297,N_6639,N_6629);
nand U7298 (N_7298,N_6058,N_6414);
and U7299 (N_7299,N_6067,N_6772);
nand U7300 (N_7300,N_6973,N_6506);
or U7301 (N_7301,N_6945,N_6978);
and U7302 (N_7302,N_6896,N_6908);
or U7303 (N_7303,N_6267,N_6963);
and U7304 (N_7304,N_6017,N_6731);
nor U7305 (N_7305,N_6252,N_6367);
and U7306 (N_7306,N_6342,N_6274);
and U7307 (N_7307,N_6850,N_6065);
and U7308 (N_7308,N_6227,N_6572);
and U7309 (N_7309,N_6983,N_6109);
nor U7310 (N_7310,N_6718,N_6687);
or U7311 (N_7311,N_6878,N_6139);
nand U7312 (N_7312,N_6213,N_6318);
xnor U7313 (N_7313,N_6919,N_6462);
or U7314 (N_7314,N_6515,N_6976);
and U7315 (N_7315,N_6182,N_6823);
nor U7316 (N_7316,N_6244,N_6743);
and U7317 (N_7317,N_6348,N_6536);
nor U7318 (N_7318,N_6813,N_6783);
or U7319 (N_7319,N_6257,N_6725);
and U7320 (N_7320,N_6797,N_6085);
and U7321 (N_7321,N_6792,N_6411);
nor U7322 (N_7322,N_6343,N_6442);
or U7323 (N_7323,N_6091,N_6283);
and U7324 (N_7324,N_6075,N_6578);
and U7325 (N_7325,N_6381,N_6126);
nand U7326 (N_7326,N_6727,N_6848);
nand U7327 (N_7327,N_6726,N_6996);
nand U7328 (N_7328,N_6467,N_6840);
nor U7329 (N_7329,N_6914,N_6476);
and U7330 (N_7330,N_6391,N_6513);
xor U7331 (N_7331,N_6814,N_6500);
or U7332 (N_7332,N_6593,N_6556);
nor U7333 (N_7333,N_6705,N_6079);
nor U7334 (N_7334,N_6297,N_6520);
xnor U7335 (N_7335,N_6301,N_6043);
nand U7336 (N_7336,N_6883,N_6517);
nor U7337 (N_7337,N_6644,N_6313);
or U7338 (N_7338,N_6196,N_6636);
nor U7339 (N_7339,N_6191,N_6926);
or U7340 (N_7340,N_6816,N_6218);
and U7341 (N_7341,N_6487,N_6788);
or U7342 (N_7342,N_6247,N_6497);
xor U7343 (N_7343,N_6306,N_6852);
nand U7344 (N_7344,N_6407,N_6355);
or U7345 (N_7345,N_6929,N_6439);
or U7346 (N_7346,N_6210,N_6222);
or U7347 (N_7347,N_6153,N_6493);
nand U7348 (N_7348,N_6207,N_6715);
nand U7349 (N_7349,N_6415,N_6140);
nor U7350 (N_7350,N_6969,N_6786);
and U7351 (N_7351,N_6548,N_6627);
or U7352 (N_7352,N_6019,N_6710);
and U7353 (N_7353,N_6587,N_6007);
nor U7354 (N_7354,N_6169,N_6837);
nor U7355 (N_7355,N_6806,N_6716);
or U7356 (N_7356,N_6545,N_6450);
or U7357 (N_7357,N_6432,N_6622);
nand U7358 (N_7358,N_6295,N_6665);
and U7359 (N_7359,N_6037,N_6902);
and U7360 (N_7360,N_6984,N_6885);
nor U7361 (N_7361,N_6013,N_6133);
and U7362 (N_7362,N_6463,N_6148);
nor U7363 (N_7363,N_6756,N_6090);
or U7364 (N_7364,N_6707,N_6413);
and U7365 (N_7365,N_6172,N_6308);
and U7366 (N_7366,N_6907,N_6077);
and U7367 (N_7367,N_6349,N_6371);
and U7368 (N_7368,N_6724,N_6942);
nand U7369 (N_7369,N_6600,N_6190);
and U7370 (N_7370,N_6648,N_6358);
and U7371 (N_7371,N_6856,N_6538);
or U7372 (N_7372,N_6798,N_6968);
or U7373 (N_7373,N_6778,N_6943);
or U7374 (N_7374,N_6332,N_6607);
xor U7375 (N_7375,N_6068,N_6447);
nor U7376 (N_7376,N_6997,N_6838);
nand U7377 (N_7377,N_6539,N_6975);
nand U7378 (N_7378,N_6652,N_6009);
or U7379 (N_7379,N_6641,N_6405);
nor U7380 (N_7380,N_6917,N_6985);
nand U7381 (N_7381,N_6083,N_6451);
and U7382 (N_7382,N_6709,N_6808);
or U7383 (N_7383,N_6551,N_6029);
and U7384 (N_7384,N_6426,N_6321);
and U7385 (N_7385,N_6573,N_6564);
nor U7386 (N_7386,N_6662,N_6494);
nor U7387 (N_7387,N_6056,N_6168);
and U7388 (N_7388,N_6689,N_6842);
or U7389 (N_7389,N_6555,N_6696);
nor U7390 (N_7390,N_6238,N_6793);
or U7391 (N_7391,N_6552,N_6534);
or U7392 (N_7392,N_6701,N_6580);
or U7393 (N_7393,N_6855,N_6406);
and U7394 (N_7394,N_6892,N_6895);
or U7395 (N_7395,N_6819,N_6185);
nand U7396 (N_7396,N_6337,N_6364);
and U7397 (N_7397,N_6401,N_6047);
nor U7398 (N_7398,N_6320,N_6669);
nand U7399 (N_7399,N_6055,N_6924);
or U7400 (N_7400,N_6944,N_6512);
nor U7401 (N_7401,N_6742,N_6618);
nor U7402 (N_7402,N_6104,N_6338);
nand U7403 (N_7403,N_6480,N_6490);
nor U7404 (N_7404,N_6229,N_6032);
and U7405 (N_7405,N_6519,N_6273);
nand U7406 (N_7406,N_6928,N_6034);
nand U7407 (N_7407,N_6479,N_6200);
and U7408 (N_7408,N_6980,N_6981);
nand U7409 (N_7409,N_6799,N_6723);
and U7410 (N_7410,N_6491,N_6904);
or U7411 (N_7411,N_6383,N_6050);
nor U7412 (N_7412,N_6776,N_6341);
and U7413 (N_7413,N_6431,N_6445);
or U7414 (N_7414,N_6589,N_6979);
and U7415 (N_7415,N_6998,N_6062);
nand U7416 (N_7416,N_6327,N_6810);
nor U7417 (N_7417,N_6204,N_6554);
and U7418 (N_7418,N_6531,N_6645);
nand U7419 (N_7419,N_6865,N_6708);
and U7420 (N_7420,N_6815,N_6905);
nor U7421 (N_7421,N_6800,N_6672);
nor U7422 (N_7422,N_6750,N_6794);
nand U7423 (N_7423,N_6284,N_6232);
or U7424 (N_7424,N_6533,N_6354);
and U7425 (N_7425,N_6184,N_6137);
or U7426 (N_7426,N_6565,N_6166);
nand U7427 (N_7427,N_6664,N_6010);
nor U7428 (N_7428,N_6473,N_6240);
nand U7429 (N_7429,N_6658,N_6616);
nand U7430 (N_7430,N_6635,N_6334);
nor U7431 (N_7431,N_6893,N_6192);
nor U7432 (N_7432,N_6080,N_6333);
or U7433 (N_7433,N_6205,N_6879);
and U7434 (N_7434,N_6351,N_6481);
nand U7435 (N_7435,N_6590,N_6544);
or U7436 (N_7436,N_6755,N_6999);
and U7437 (N_7437,N_6285,N_6241);
or U7438 (N_7438,N_6507,N_6030);
or U7439 (N_7439,N_6647,N_6563);
nand U7440 (N_7440,N_6775,N_6595);
and U7441 (N_7441,N_6927,N_6675);
nand U7442 (N_7442,N_6986,N_6397);
and U7443 (N_7443,N_6875,N_6992);
and U7444 (N_7444,N_6000,N_6760);
and U7445 (N_7445,N_6022,N_6862);
or U7446 (N_7446,N_6041,N_6948);
nand U7447 (N_7447,N_6741,N_6023);
or U7448 (N_7448,N_6006,N_6201);
or U7449 (N_7449,N_6577,N_6660);
and U7450 (N_7450,N_6398,N_6177);
and U7451 (N_7451,N_6894,N_6540);
or U7452 (N_7452,N_6160,N_6178);
xor U7453 (N_7453,N_6005,N_6818);
nor U7454 (N_7454,N_6208,N_6368);
nor U7455 (N_7455,N_6753,N_6631);
or U7456 (N_7456,N_6935,N_6585);
nand U7457 (N_7457,N_6131,N_6380);
nand U7458 (N_7458,N_6441,N_6746);
xor U7459 (N_7459,N_6890,N_6542);
nor U7460 (N_7460,N_6394,N_6360);
or U7461 (N_7461,N_6221,N_6537);
and U7462 (N_7462,N_6958,N_6938);
nor U7463 (N_7463,N_6416,N_6363);
and U7464 (N_7464,N_6176,N_6597);
nand U7465 (N_7465,N_6530,N_6151);
or U7466 (N_7466,N_6106,N_6962);
or U7467 (N_7467,N_6250,N_6461);
xor U7468 (N_7468,N_6874,N_6399);
or U7469 (N_7469,N_6254,N_6594);
and U7470 (N_7470,N_6866,N_6054);
or U7471 (N_7471,N_6440,N_6566);
and U7472 (N_7472,N_6623,N_6161);
nand U7473 (N_7473,N_6617,N_6913);
or U7474 (N_7474,N_6972,N_6149);
or U7475 (N_7475,N_6372,N_6884);
or U7476 (N_7476,N_6084,N_6784);
and U7477 (N_7477,N_6434,N_6216);
and U7478 (N_7478,N_6307,N_6188);
and U7479 (N_7479,N_6156,N_6099);
nor U7480 (N_7480,N_6909,N_6231);
and U7481 (N_7481,N_6269,N_6762);
or U7482 (N_7482,N_6899,N_6008);
nor U7483 (N_7483,N_6299,N_6703);
nand U7484 (N_7484,N_6093,N_6915);
nand U7485 (N_7485,N_6575,N_6039);
nand U7486 (N_7486,N_6117,N_6849);
nand U7487 (N_7487,N_6279,N_6045);
or U7488 (N_7488,N_6028,N_6164);
or U7489 (N_7489,N_6959,N_6780);
nand U7490 (N_7490,N_6843,N_6827);
or U7491 (N_7491,N_6604,N_6403);
nor U7492 (N_7492,N_6135,N_6768);
and U7493 (N_7493,N_6974,N_6033);
nand U7494 (N_7494,N_6187,N_6745);
and U7495 (N_7495,N_6933,N_6853);
or U7496 (N_7496,N_6402,N_6266);
nand U7497 (N_7497,N_6438,N_6730);
or U7498 (N_7498,N_6596,N_6643);
xor U7499 (N_7499,N_6860,N_6362);
xor U7500 (N_7500,N_6968,N_6326);
nand U7501 (N_7501,N_6168,N_6289);
and U7502 (N_7502,N_6579,N_6809);
and U7503 (N_7503,N_6669,N_6909);
nor U7504 (N_7504,N_6451,N_6615);
nand U7505 (N_7505,N_6755,N_6239);
nor U7506 (N_7506,N_6895,N_6551);
nor U7507 (N_7507,N_6717,N_6186);
or U7508 (N_7508,N_6464,N_6581);
nor U7509 (N_7509,N_6994,N_6089);
or U7510 (N_7510,N_6377,N_6263);
and U7511 (N_7511,N_6231,N_6391);
nand U7512 (N_7512,N_6394,N_6282);
nor U7513 (N_7513,N_6363,N_6497);
nand U7514 (N_7514,N_6778,N_6432);
or U7515 (N_7515,N_6398,N_6846);
nor U7516 (N_7516,N_6854,N_6789);
and U7517 (N_7517,N_6583,N_6849);
and U7518 (N_7518,N_6353,N_6261);
nand U7519 (N_7519,N_6255,N_6832);
nand U7520 (N_7520,N_6225,N_6302);
nand U7521 (N_7521,N_6291,N_6743);
nor U7522 (N_7522,N_6721,N_6179);
nor U7523 (N_7523,N_6719,N_6964);
nor U7524 (N_7524,N_6852,N_6822);
nand U7525 (N_7525,N_6110,N_6306);
or U7526 (N_7526,N_6880,N_6945);
nor U7527 (N_7527,N_6764,N_6345);
or U7528 (N_7528,N_6172,N_6936);
nand U7529 (N_7529,N_6045,N_6100);
and U7530 (N_7530,N_6849,N_6872);
nand U7531 (N_7531,N_6471,N_6759);
or U7532 (N_7532,N_6926,N_6842);
and U7533 (N_7533,N_6927,N_6192);
or U7534 (N_7534,N_6386,N_6658);
nand U7535 (N_7535,N_6417,N_6986);
and U7536 (N_7536,N_6745,N_6413);
and U7537 (N_7537,N_6321,N_6130);
nand U7538 (N_7538,N_6719,N_6992);
or U7539 (N_7539,N_6612,N_6380);
nor U7540 (N_7540,N_6810,N_6445);
nor U7541 (N_7541,N_6818,N_6939);
nor U7542 (N_7542,N_6619,N_6252);
nor U7543 (N_7543,N_6474,N_6131);
nor U7544 (N_7544,N_6090,N_6519);
and U7545 (N_7545,N_6983,N_6191);
nor U7546 (N_7546,N_6148,N_6963);
or U7547 (N_7547,N_6437,N_6041);
nand U7548 (N_7548,N_6218,N_6934);
and U7549 (N_7549,N_6693,N_6651);
and U7550 (N_7550,N_6781,N_6635);
nor U7551 (N_7551,N_6039,N_6176);
and U7552 (N_7552,N_6334,N_6251);
and U7553 (N_7553,N_6175,N_6546);
and U7554 (N_7554,N_6393,N_6256);
or U7555 (N_7555,N_6444,N_6166);
nand U7556 (N_7556,N_6402,N_6700);
xor U7557 (N_7557,N_6484,N_6550);
nor U7558 (N_7558,N_6546,N_6950);
nor U7559 (N_7559,N_6499,N_6278);
nor U7560 (N_7560,N_6282,N_6831);
nand U7561 (N_7561,N_6235,N_6681);
and U7562 (N_7562,N_6363,N_6042);
nand U7563 (N_7563,N_6396,N_6059);
nand U7564 (N_7564,N_6967,N_6013);
nand U7565 (N_7565,N_6629,N_6561);
or U7566 (N_7566,N_6623,N_6867);
or U7567 (N_7567,N_6139,N_6577);
nand U7568 (N_7568,N_6402,N_6489);
nor U7569 (N_7569,N_6333,N_6691);
or U7570 (N_7570,N_6204,N_6292);
nor U7571 (N_7571,N_6214,N_6032);
or U7572 (N_7572,N_6120,N_6179);
nand U7573 (N_7573,N_6134,N_6168);
nand U7574 (N_7574,N_6612,N_6574);
nor U7575 (N_7575,N_6706,N_6969);
or U7576 (N_7576,N_6555,N_6475);
nor U7577 (N_7577,N_6662,N_6371);
or U7578 (N_7578,N_6635,N_6644);
xor U7579 (N_7579,N_6938,N_6864);
nor U7580 (N_7580,N_6390,N_6209);
xor U7581 (N_7581,N_6737,N_6899);
nand U7582 (N_7582,N_6444,N_6527);
or U7583 (N_7583,N_6462,N_6098);
and U7584 (N_7584,N_6399,N_6030);
and U7585 (N_7585,N_6506,N_6324);
or U7586 (N_7586,N_6619,N_6900);
nor U7587 (N_7587,N_6288,N_6859);
nand U7588 (N_7588,N_6349,N_6494);
nand U7589 (N_7589,N_6350,N_6921);
nor U7590 (N_7590,N_6414,N_6241);
and U7591 (N_7591,N_6553,N_6590);
or U7592 (N_7592,N_6363,N_6237);
nor U7593 (N_7593,N_6410,N_6161);
nor U7594 (N_7594,N_6557,N_6992);
and U7595 (N_7595,N_6520,N_6683);
and U7596 (N_7596,N_6784,N_6332);
or U7597 (N_7597,N_6253,N_6731);
nand U7598 (N_7598,N_6104,N_6869);
nor U7599 (N_7599,N_6322,N_6066);
or U7600 (N_7600,N_6792,N_6909);
and U7601 (N_7601,N_6487,N_6357);
nor U7602 (N_7602,N_6930,N_6614);
and U7603 (N_7603,N_6418,N_6434);
and U7604 (N_7604,N_6079,N_6192);
and U7605 (N_7605,N_6026,N_6814);
xnor U7606 (N_7606,N_6046,N_6972);
or U7607 (N_7607,N_6597,N_6331);
and U7608 (N_7608,N_6772,N_6586);
nor U7609 (N_7609,N_6949,N_6472);
nor U7610 (N_7610,N_6153,N_6998);
nand U7611 (N_7611,N_6993,N_6381);
nor U7612 (N_7612,N_6742,N_6812);
and U7613 (N_7613,N_6448,N_6863);
nand U7614 (N_7614,N_6540,N_6049);
or U7615 (N_7615,N_6882,N_6825);
nand U7616 (N_7616,N_6270,N_6062);
nor U7617 (N_7617,N_6289,N_6488);
nor U7618 (N_7618,N_6462,N_6642);
and U7619 (N_7619,N_6372,N_6354);
nand U7620 (N_7620,N_6720,N_6114);
or U7621 (N_7621,N_6249,N_6185);
nand U7622 (N_7622,N_6976,N_6585);
nor U7623 (N_7623,N_6060,N_6230);
xnor U7624 (N_7624,N_6363,N_6429);
xnor U7625 (N_7625,N_6385,N_6638);
and U7626 (N_7626,N_6495,N_6784);
or U7627 (N_7627,N_6454,N_6031);
and U7628 (N_7628,N_6185,N_6649);
nor U7629 (N_7629,N_6603,N_6291);
nor U7630 (N_7630,N_6096,N_6264);
and U7631 (N_7631,N_6914,N_6399);
nor U7632 (N_7632,N_6985,N_6384);
or U7633 (N_7633,N_6296,N_6294);
and U7634 (N_7634,N_6618,N_6928);
or U7635 (N_7635,N_6204,N_6651);
nand U7636 (N_7636,N_6880,N_6576);
nor U7637 (N_7637,N_6382,N_6496);
or U7638 (N_7638,N_6654,N_6397);
or U7639 (N_7639,N_6185,N_6449);
nand U7640 (N_7640,N_6920,N_6866);
or U7641 (N_7641,N_6269,N_6544);
nor U7642 (N_7642,N_6108,N_6037);
nand U7643 (N_7643,N_6162,N_6693);
or U7644 (N_7644,N_6028,N_6397);
nand U7645 (N_7645,N_6172,N_6822);
nand U7646 (N_7646,N_6105,N_6981);
or U7647 (N_7647,N_6687,N_6538);
nor U7648 (N_7648,N_6187,N_6488);
and U7649 (N_7649,N_6248,N_6422);
nor U7650 (N_7650,N_6756,N_6381);
and U7651 (N_7651,N_6072,N_6003);
or U7652 (N_7652,N_6859,N_6811);
xnor U7653 (N_7653,N_6559,N_6181);
and U7654 (N_7654,N_6415,N_6381);
and U7655 (N_7655,N_6904,N_6712);
and U7656 (N_7656,N_6914,N_6815);
and U7657 (N_7657,N_6158,N_6800);
and U7658 (N_7658,N_6930,N_6912);
and U7659 (N_7659,N_6907,N_6691);
nand U7660 (N_7660,N_6577,N_6905);
nor U7661 (N_7661,N_6679,N_6503);
or U7662 (N_7662,N_6473,N_6720);
nand U7663 (N_7663,N_6071,N_6942);
nand U7664 (N_7664,N_6965,N_6087);
or U7665 (N_7665,N_6922,N_6849);
nand U7666 (N_7666,N_6592,N_6435);
and U7667 (N_7667,N_6273,N_6713);
nor U7668 (N_7668,N_6940,N_6605);
nor U7669 (N_7669,N_6618,N_6453);
or U7670 (N_7670,N_6650,N_6194);
and U7671 (N_7671,N_6682,N_6502);
nand U7672 (N_7672,N_6393,N_6848);
nand U7673 (N_7673,N_6656,N_6653);
nor U7674 (N_7674,N_6084,N_6770);
or U7675 (N_7675,N_6460,N_6937);
and U7676 (N_7676,N_6547,N_6447);
or U7677 (N_7677,N_6119,N_6590);
nand U7678 (N_7678,N_6150,N_6364);
and U7679 (N_7679,N_6105,N_6529);
and U7680 (N_7680,N_6534,N_6103);
nand U7681 (N_7681,N_6463,N_6403);
nand U7682 (N_7682,N_6638,N_6157);
nor U7683 (N_7683,N_6701,N_6116);
nand U7684 (N_7684,N_6383,N_6409);
and U7685 (N_7685,N_6330,N_6668);
nand U7686 (N_7686,N_6943,N_6525);
nor U7687 (N_7687,N_6435,N_6070);
nand U7688 (N_7688,N_6910,N_6079);
and U7689 (N_7689,N_6188,N_6577);
nor U7690 (N_7690,N_6462,N_6046);
and U7691 (N_7691,N_6019,N_6847);
nor U7692 (N_7692,N_6076,N_6770);
and U7693 (N_7693,N_6270,N_6085);
nand U7694 (N_7694,N_6278,N_6008);
nor U7695 (N_7695,N_6154,N_6736);
or U7696 (N_7696,N_6967,N_6711);
nand U7697 (N_7697,N_6447,N_6643);
or U7698 (N_7698,N_6250,N_6357);
nand U7699 (N_7699,N_6498,N_6525);
nor U7700 (N_7700,N_6739,N_6439);
nor U7701 (N_7701,N_6238,N_6405);
nor U7702 (N_7702,N_6535,N_6787);
and U7703 (N_7703,N_6318,N_6447);
nand U7704 (N_7704,N_6512,N_6170);
nand U7705 (N_7705,N_6766,N_6268);
nor U7706 (N_7706,N_6466,N_6790);
or U7707 (N_7707,N_6100,N_6669);
and U7708 (N_7708,N_6638,N_6774);
nand U7709 (N_7709,N_6484,N_6413);
and U7710 (N_7710,N_6020,N_6758);
nand U7711 (N_7711,N_6119,N_6584);
or U7712 (N_7712,N_6630,N_6490);
nor U7713 (N_7713,N_6088,N_6662);
or U7714 (N_7714,N_6443,N_6240);
nor U7715 (N_7715,N_6358,N_6225);
and U7716 (N_7716,N_6836,N_6673);
nand U7717 (N_7717,N_6408,N_6062);
nor U7718 (N_7718,N_6311,N_6528);
and U7719 (N_7719,N_6327,N_6072);
or U7720 (N_7720,N_6179,N_6686);
nand U7721 (N_7721,N_6125,N_6174);
nand U7722 (N_7722,N_6402,N_6463);
or U7723 (N_7723,N_6562,N_6773);
nand U7724 (N_7724,N_6920,N_6413);
nand U7725 (N_7725,N_6303,N_6402);
or U7726 (N_7726,N_6055,N_6702);
and U7727 (N_7727,N_6556,N_6175);
or U7728 (N_7728,N_6836,N_6276);
or U7729 (N_7729,N_6578,N_6126);
and U7730 (N_7730,N_6698,N_6051);
and U7731 (N_7731,N_6052,N_6687);
nor U7732 (N_7732,N_6839,N_6121);
nor U7733 (N_7733,N_6704,N_6253);
and U7734 (N_7734,N_6451,N_6453);
nand U7735 (N_7735,N_6192,N_6046);
and U7736 (N_7736,N_6844,N_6520);
nor U7737 (N_7737,N_6236,N_6289);
or U7738 (N_7738,N_6861,N_6283);
nor U7739 (N_7739,N_6746,N_6548);
nand U7740 (N_7740,N_6238,N_6408);
and U7741 (N_7741,N_6955,N_6704);
or U7742 (N_7742,N_6993,N_6125);
nor U7743 (N_7743,N_6984,N_6985);
nand U7744 (N_7744,N_6883,N_6790);
and U7745 (N_7745,N_6038,N_6969);
and U7746 (N_7746,N_6648,N_6140);
nor U7747 (N_7747,N_6974,N_6092);
nand U7748 (N_7748,N_6666,N_6271);
nor U7749 (N_7749,N_6932,N_6070);
or U7750 (N_7750,N_6546,N_6380);
nand U7751 (N_7751,N_6111,N_6527);
or U7752 (N_7752,N_6022,N_6233);
or U7753 (N_7753,N_6297,N_6414);
nor U7754 (N_7754,N_6570,N_6217);
nand U7755 (N_7755,N_6650,N_6441);
and U7756 (N_7756,N_6841,N_6121);
nand U7757 (N_7757,N_6086,N_6907);
or U7758 (N_7758,N_6661,N_6625);
nor U7759 (N_7759,N_6798,N_6274);
and U7760 (N_7760,N_6146,N_6986);
nor U7761 (N_7761,N_6738,N_6394);
nor U7762 (N_7762,N_6928,N_6531);
or U7763 (N_7763,N_6231,N_6359);
nor U7764 (N_7764,N_6456,N_6122);
and U7765 (N_7765,N_6923,N_6626);
nand U7766 (N_7766,N_6507,N_6124);
nor U7767 (N_7767,N_6382,N_6504);
and U7768 (N_7768,N_6725,N_6505);
and U7769 (N_7769,N_6276,N_6658);
or U7770 (N_7770,N_6035,N_6774);
nor U7771 (N_7771,N_6125,N_6072);
nor U7772 (N_7772,N_6853,N_6263);
and U7773 (N_7773,N_6513,N_6101);
nor U7774 (N_7774,N_6644,N_6114);
and U7775 (N_7775,N_6159,N_6397);
nand U7776 (N_7776,N_6511,N_6697);
nand U7777 (N_7777,N_6649,N_6789);
and U7778 (N_7778,N_6902,N_6979);
nand U7779 (N_7779,N_6333,N_6744);
nor U7780 (N_7780,N_6654,N_6965);
xnor U7781 (N_7781,N_6721,N_6034);
and U7782 (N_7782,N_6575,N_6502);
nand U7783 (N_7783,N_6473,N_6241);
or U7784 (N_7784,N_6035,N_6467);
or U7785 (N_7785,N_6892,N_6710);
and U7786 (N_7786,N_6903,N_6502);
nand U7787 (N_7787,N_6805,N_6802);
and U7788 (N_7788,N_6332,N_6221);
nand U7789 (N_7789,N_6435,N_6340);
or U7790 (N_7790,N_6276,N_6133);
nor U7791 (N_7791,N_6504,N_6476);
nor U7792 (N_7792,N_6122,N_6533);
nor U7793 (N_7793,N_6878,N_6940);
nor U7794 (N_7794,N_6824,N_6327);
nor U7795 (N_7795,N_6408,N_6613);
or U7796 (N_7796,N_6479,N_6766);
nand U7797 (N_7797,N_6372,N_6240);
and U7798 (N_7798,N_6829,N_6801);
or U7799 (N_7799,N_6231,N_6456);
nor U7800 (N_7800,N_6804,N_6062);
or U7801 (N_7801,N_6914,N_6837);
or U7802 (N_7802,N_6548,N_6634);
nor U7803 (N_7803,N_6081,N_6107);
or U7804 (N_7804,N_6368,N_6988);
and U7805 (N_7805,N_6625,N_6882);
and U7806 (N_7806,N_6104,N_6245);
or U7807 (N_7807,N_6022,N_6972);
nor U7808 (N_7808,N_6691,N_6899);
nand U7809 (N_7809,N_6964,N_6091);
nor U7810 (N_7810,N_6379,N_6736);
or U7811 (N_7811,N_6638,N_6858);
and U7812 (N_7812,N_6889,N_6214);
and U7813 (N_7813,N_6907,N_6895);
xor U7814 (N_7814,N_6836,N_6724);
or U7815 (N_7815,N_6994,N_6911);
and U7816 (N_7816,N_6352,N_6058);
and U7817 (N_7817,N_6451,N_6082);
and U7818 (N_7818,N_6735,N_6567);
nor U7819 (N_7819,N_6459,N_6738);
and U7820 (N_7820,N_6001,N_6534);
nand U7821 (N_7821,N_6084,N_6284);
nor U7822 (N_7822,N_6248,N_6753);
nand U7823 (N_7823,N_6693,N_6727);
nor U7824 (N_7824,N_6508,N_6102);
nand U7825 (N_7825,N_6284,N_6462);
nor U7826 (N_7826,N_6642,N_6267);
nor U7827 (N_7827,N_6149,N_6102);
or U7828 (N_7828,N_6432,N_6474);
xnor U7829 (N_7829,N_6942,N_6525);
nor U7830 (N_7830,N_6625,N_6803);
nor U7831 (N_7831,N_6562,N_6948);
and U7832 (N_7832,N_6431,N_6950);
nand U7833 (N_7833,N_6870,N_6440);
and U7834 (N_7834,N_6314,N_6566);
nand U7835 (N_7835,N_6561,N_6019);
nand U7836 (N_7836,N_6284,N_6351);
nor U7837 (N_7837,N_6271,N_6619);
nand U7838 (N_7838,N_6191,N_6916);
and U7839 (N_7839,N_6931,N_6976);
or U7840 (N_7840,N_6755,N_6908);
nor U7841 (N_7841,N_6532,N_6836);
or U7842 (N_7842,N_6740,N_6781);
and U7843 (N_7843,N_6026,N_6686);
or U7844 (N_7844,N_6270,N_6974);
and U7845 (N_7845,N_6214,N_6251);
and U7846 (N_7846,N_6406,N_6093);
nand U7847 (N_7847,N_6598,N_6277);
nor U7848 (N_7848,N_6287,N_6330);
nor U7849 (N_7849,N_6533,N_6412);
nor U7850 (N_7850,N_6762,N_6568);
nand U7851 (N_7851,N_6365,N_6739);
nor U7852 (N_7852,N_6015,N_6168);
and U7853 (N_7853,N_6246,N_6987);
nor U7854 (N_7854,N_6096,N_6834);
or U7855 (N_7855,N_6383,N_6121);
nand U7856 (N_7856,N_6200,N_6730);
nand U7857 (N_7857,N_6290,N_6261);
nand U7858 (N_7858,N_6560,N_6819);
nor U7859 (N_7859,N_6108,N_6702);
or U7860 (N_7860,N_6614,N_6660);
xor U7861 (N_7861,N_6041,N_6040);
or U7862 (N_7862,N_6456,N_6391);
xor U7863 (N_7863,N_6674,N_6434);
nor U7864 (N_7864,N_6277,N_6611);
nor U7865 (N_7865,N_6696,N_6294);
and U7866 (N_7866,N_6919,N_6995);
or U7867 (N_7867,N_6153,N_6013);
nand U7868 (N_7868,N_6581,N_6403);
nand U7869 (N_7869,N_6013,N_6124);
and U7870 (N_7870,N_6807,N_6916);
and U7871 (N_7871,N_6956,N_6065);
nand U7872 (N_7872,N_6133,N_6203);
or U7873 (N_7873,N_6541,N_6147);
nand U7874 (N_7874,N_6360,N_6219);
nor U7875 (N_7875,N_6187,N_6211);
or U7876 (N_7876,N_6875,N_6486);
and U7877 (N_7877,N_6163,N_6354);
nand U7878 (N_7878,N_6950,N_6763);
or U7879 (N_7879,N_6148,N_6792);
or U7880 (N_7880,N_6866,N_6404);
nor U7881 (N_7881,N_6058,N_6849);
nor U7882 (N_7882,N_6030,N_6906);
nand U7883 (N_7883,N_6178,N_6347);
nor U7884 (N_7884,N_6077,N_6894);
and U7885 (N_7885,N_6874,N_6499);
nor U7886 (N_7886,N_6198,N_6125);
and U7887 (N_7887,N_6604,N_6692);
and U7888 (N_7888,N_6286,N_6102);
nand U7889 (N_7889,N_6993,N_6275);
or U7890 (N_7890,N_6523,N_6205);
nand U7891 (N_7891,N_6169,N_6087);
or U7892 (N_7892,N_6204,N_6142);
and U7893 (N_7893,N_6379,N_6555);
and U7894 (N_7894,N_6545,N_6721);
and U7895 (N_7895,N_6664,N_6956);
nor U7896 (N_7896,N_6476,N_6845);
nand U7897 (N_7897,N_6636,N_6697);
or U7898 (N_7898,N_6821,N_6272);
nor U7899 (N_7899,N_6713,N_6913);
nand U7900 (N_7900,N_6377,N_6282);
or U7901 (N_7901,N_6204,N_6960);
nand U7902 (N_7902,N_6840,N_6147);
nand U7903 (N_7903,N_6887,N_6991);
or U7904 (N_7904,N_6325,N_6930);
or U7905 (N_7905,N_6518,N_6028);
nor U7906 (N_7906,N_6930,N_6229);
or U7907 (N_7907,N_6588,N_6363);
xnor U7908 (N_7908,N_6634,N_6465);
or U7909 (N_7909,N_6076,N_6874);
nor U7910 (N_7910,N_6411,N_6778);
nor U7911 (N_7911,N_6312,N_6832);
nand U7912 (N_7912,N_6427,N_6682);
and U7913 (N_7913,N_6125,N_6294);
or U7914 (N_7914,N_6515,N_6088);
or U7915 (N_7915,N_6093,N_6309);
or U7916 (N_7916,N_6444,N_6715);
and U7917 (N_7917,N_6011,N_6916);
nand U7918 (N_7918,N_6829,N_6164);
or U7919 (N_7919,N_6029,N_6696);
nor U7920 (N_7920,N_6175,N_6414);
or U7921 (N_7921,N_6430,N_6787);
xnor U7922 (N_7922,N_6678,N_6126);
and U7923 (N_7923,N_6264,N_6177);
or U7924 (N_7924,N_6516,N_6022);
nor U7925 (N_7925,N_6501,N_6316);
nand U7926 (N_7926,N_6374,N_6314);
or U7927 (N_7927,N_6906,N_6680);
nand U7928 (N_7928,N_6326,N_6824);
and U7929 (N_7929,N_6504,N_6735);
and U7930 (N_7930,N_6255,N_6961);
or U7931 (N_7931,N_6598,N_6122);
nor U7932 (N_7932,N_6792,N_6225);
or U7933 (N_7933,N_6866,N_6867);
nor U7934 (N_7934,N_6858,N_6261);
nand U7935 (N_7935,N_6652,N_6843);
and U7936 (N_7936,N_6651,N_6609);
nor U7937 (N_7937,N_6517,N_6937);
or U7938 (N_7938,N_6805,N_6774);
nor U7939 (N_7939,N_6497,N_6494);
nor U7940 (N_7940,N_6105,N_6175);
and U7941 (N_7941,N_6465,N_6971);
and U7942 (N_7942,N_6547,N_6379);
nor U7943 (N_7943,N_6317,N_6800);
nor U7944 (N_7944,N_6475,N_6200);
or U7945 (N_7945,N_6314,N_6256);
and U7946 (N_7946,N_6693,N_6445);
or U7947 (N_7947,N_6538,N_6960);
and U7948 (N_7948,N_6704,N_6214);
and U7949 (N_7949,N_6435,N_6296);
and U7950 (N_7950,N_6663,N_6510);
nor U7951 (N_7951,N_6019,N_6551);
and U7952 (N_7952,N_6421,N_6658);
or U7953 (N_7953,N_6019,N_6022);
and U7954 (N_7954,N_6767,N_6800);
and U7955 (N_7955,N_6355,N_6527);
or U7956 (N_7956,N_6088,N_6887);
xnor U7957 (N_7957,N_6231,N_6341);
and U7958 (N_7958,N_6631,N_6060);
and U7959 (N_7959,N_6377,N_6053);
and U7960 (N_7960,N_6738,N_6215);
or U7961 (N_7961,N_6572,N_6701);
nand U7962 (N_7962,N_6125,N_6078);
and U7963 (N_7963,N_6481,N_6923);
nand U7964 (N_7964,N_6498,N_6797);
or U7965 (N_7965,N_6568,N_6810);
or U7966 (N_7966,N_6456,N_6702);
nor U7967 (N_7967,N_6330,N_6005);
nand U7968 (N_7968,N_6622,N_6773);
or U7969 (N_7969,N_6534,N_6080);
or U7970 (N_7970,N_6927,N_6894);
nor U7971 (N_7971,N_6451,N_6221);
or U7972 (N_7972,N_6208,N_6480);
and U7973 (N_7973,N_6027,N_6456);
nand U7974 (N_7974,N_6895,N_6714);
and U7975 (N_7975,N_6390,N_6072);
xor U7976 (N_7976,N_6647,N_6790);
or U7977 (N_7977,N_6324,N_6377);
nand U7978 (N_7978,N_6087,N_6236);
nand U7979 (N_7979,N_6885,N_6942);
nand U7980 (N_7980,N_6337,N_6267);
nor U7981 (N_7981,N_6568,N_6545);
nand U7982 (N_7982,N_6411,N_6988);
nor U7983 (N_7983,N_6564,N_6839);
nor U7984 (N_7984,N_6819,N_6081);
or U7985 (N_7985,N_6734,N_6882);
nor U7986 (N_7986,N_6608,N_6259);
or U7987 (N_7987,N_6123,N_6390);
nand U7988 (N_7988,N_6502,N_6435);
or U7989 (N_7989,N_6392,N_6376);
nand U7990 (N_7990,N_6594,N_6907);
nand U7991 (N_7991,N_6918,N_6407);
and U7992 (N_7992,N_6154,N_6565);
or U7993 (N_7993,N_6691,N_6605);
nand U7994 (N_7994,N_6508,N_6111);
or U7995 (N_7995,N_6008,N_6795);
nand U7996 (N_7996,N_6112,N_6939);
nor U7997 (N_7997,N_6676,N_6971);
nand U7998 (N_7998,N_6166,N_6526);
and U7999 (N_7999,N_6446,N_6255);
nand U8000 (N_8000,N_7269,N_7076);
nand U8001 (N_8001,N_7597,N_7032);
nor U8002 (N_8002,N_7748,N_7384);
or U8003 (N_8003,N_7713,N_7120);
and U8004 (N_8004,N_7729,N_7387);
nor U8005 (N_8005,N_7179,N_7295);
nand U8006 (N_8006,N_7945,N_7954);
nor U8007 (N_8007,N_7836,N_7990);
nor U8008 (N_8008,N_7425,N_7916);
and U8009 (N_8009,N_7920,N_7173);
nand U8010 (N_8010,N_7195,N_7490);
nor U8011 (N_8011,N_7083,N_7242);
nand U8012 (N_8012,N_7587,N_7725);
and U8013 (N_8013,N_7449,N_7999);
and U8014 (N_8014,N_7872,N_7839);
nor U8015 (N_8015,N_7797,N_7416);
and U8016 (N_8016,N_7311,N_7393);
and U8017 (N_8017,N_7708,N_7956);
or U8018 (N_8018,N_7306,N_7352);
nand U8019 (N_8019,N_7267,N_7706);
and U8020 (N_8020,N_7506,N_7875);
and U8021 (N_8021,N_7130,N_7517);
and U8022 (N_8022,N_7371,N_7879);
or U8023 (N_8023,N_7344,N_7996);
or U8024 (N_8024,N_7511,N_7833);
nand U8025 (N_8025,N_7027,N_7781);
and U8026 (N_8026,N_7564,N_7756);
or U8027 (N_8027,N_7318,N_7406);
and U8028 (N_8028,N_7635,N_7753);
nand U8029 (N_8029,N_7168,N_7657);
nor U8030 (N_8030,N_7923,N_7550);
and U8031 (N_8031,N_7855,N_7759);
or U8032 (N_8032,N_7377,N_7693);
nor U8033 (N_8033,N_7200,N_7362);
nor U8034 (N_8034,N_7335,N_7622);
xnor U8035 (N_8035,N_7626,N_7779);
nand U8036 (N_8036,N_7094,N_7343);
and U8037 (N_8037,N_7128,N_7261);
nor U8038 (N_8038,N_7003,N_7288);
and U8039 (N_8039,N_7176,N_7818);
or U8040 (N_8040,N_7798,N_7356);
and U8041 (N_8041,N_7840,N_7978);
nand U8042 (N_8042,N_7791,N_7562);
nor U8043 (N_8043,N_7915,N_7320);
nor U8044 (N_8044,N_7736,N_7323);
or U8045 (N_8045,N_7560,N_7628);
nand U8046 (N_8046,N_7636,N_7512);
nor U8047 (N_8047,N_7040,N_7240);
nand U8048 (N_8048,N_7935,N_7627);
and U8049 (N_8049,N_7378,N_7086);
nand U8050 (N_8050,N_7846,N_7165);
nor U8051 (N_8051,N_7834,N_7680);
or U8052 (N_8052,N_7334,N_7767);
nand U8053 (N_8053,N_7896,N_7648);
and U8054 (N_8054,N_7357,N_7676);
and U8055 (N_8055,N_7654,N_7848);
nor U8056 (N_8056,N_7073,N_7022);
or U8057 (N_8057,N_7931,N_7375);
or U8058 (N_8058,N_7556,N_7910);
nand U8059 (N_8059,N_7229,N_7289);
nor U8060 (N_8060,N_7755,N_7031);
or U8061 (N_8061,N_7230,N_7637);
nor U8062 (N_8062,N_7749,N_7919);
nor U8063 (N_8063,N_7614,N_7763);
and U8064 (N_8064,N_7710,N_7889);
and U8065 (N_8065,N_7442,N_7381);
or U8066 (N_8066,N_7502,N_7093);
nor U8067 (N_8067,N_7095,N_7743);
nand U8068 (N_8068,N_7629,N_7058);
nand U8069 (N_8069,N_7390,N_7816);
and U8070 (N_8070,N_7973,N_7015);
nor U8071 (N_8071,N_7801,N_7547);
and U8072 (N_8072,N_7067,N_7604);
nor U8073 (N_8073,N_7471,N_7479);
or U8074 (N_8074,N_7528,N_7602);
nand U8075 (N_8075,N_7035,N_7227);
nor U8076 (N_8076,N_7109,N_7641);
nand U8077 (N_8077,N_7431,N_7665);
and U8078 (N_8078,N_7762,N_7147);
nor U8079 (N_8079,N_7868,N_7582);
and U8080 (N_8080,N_7145,N_7522);
nor U8081 (N_8081,N_7722,N_7744);
and U8082 (N_8082,N_7829,N_7687);
nand U8083 (N_8083,N_7271,N_7215);
and U8084 (N_8084,N_7853,N_7322);
or U8085 (N_8085,N_7606,N_7050);
nor U8086 (N_8086,N_7433,N_7194);
and U8087 (N_8087,N_7129,N_7890);
nor U8088 (N_8088,N_7441,N_7161);
or U8089 (N_8089,N_7366,N_7893);
or U8090 (N_8090,N_7373,N_7102);
nand U8091 (N_8091,N_7470,N_7809);
and U8092 (N_8092,N_7402,N_7336);
and U8093 (N_8093,N_7877,N_7752);
nand U8094 (N_8094,N_7515,N_7726);
nand U8095 (N_8095,N_7354,N_7066);
nand U8096 (N_8096,N_7467,N_7717);
and U8097 (N_8097,N_7319,N_7014);
or U8098 (N_8098,N_7538,N_7851);
or U8099 (N_8099,N_7291,N_7447);
and U8100 (N_8100,N_7980,N_7424);
and U8101 (N_8101,N_7972,N_7939);
or U8102 (N_8102,N_7151,N_7598);
and U8103 (N_8103,N_7225,N_7118);
or U8104 (N_8104,N_7566,N_7312);
and U8105 (N_8105,N_7827,N_7503);
or U8106 (N_8106,N_7274,N_7302);
nor U8107 (N_8107,N_7739,N_7976);
nand U8108 (N_8108,N_7684,N_7310);
nand U8109 (N_8109,N_7347,N_7983);
and U8110 (N_8110,N_7329,N_7513);
nor U8111 (N_8111,N_7041,N_7080);
and U8112 (N_8112,N_7037,N_7616);
and U8113 (N_8113,N_7519,N_7249);
and U8114 (N_8114,N_7531,N_7601);
and U8115 (N_8115,N_7077,N_7275);
nand U8116 (N_8116,N_7212,N_7303);
and U8117 (N_8117,N_7305,N_7675);
or U8118 (N_8118,N_7325,N_7141);
nand U8119 (N_8119,N_7894,N_7158);
nand U8120 (N_8120,N_7439,N_7313);
nor U8121 (N_8121,N_7104,N_7701);
or U8122 (N_8122,N_7218,N_7279);
nand U8123 (N_8123,N_7097,N_7644);
or U8124 (N_8124,N_7340,N_7811);
or U8125 (N_8125,N_7342,N_7221);
or U8126 (N_8126,N_7255,N_7475);
nand U8127 (N_8127,N_7584,N_7409);
nand U8128 (N_8128,N_7984,N_7370);
nor U8129 (N_8129,N_7679,N_7139);
or U8130 (N_8130,N_7551,N_7777);
or U8131 (N_8131,N_7133,N_7651);
nor U8132 (N_8132,N_7741,N_7328);
nand U8133 (N_8133,N_7337,N_7078);
nand U8134 (N_8134,N_7673,N_7204);
or U8135 (N_8135,N_7874,N_7062);
nand U8136 (N_8136,N_7787,N_7349);
or U8137 (N_8137,N_7166,N_7188);
and U8138 (N_8138,N_7464,N_7012);
and U8139 (N_8139,N_7647,N_7358);
nand U8140 (N_8140,N_7826,N_7643);
nor U8141 (N_8141,N_7652,N_7908);
and U8142 (N_8142,N_7707,N_7505);
or U8143 (N_8143,N_7510,N_7430);
and U8144 (N_8144,N_7966,N_7372);
nor U8145 (N_8145,N_7880,N_7087);
xor U8146 (N_8146,N_7786,N_7599);
nor U8147 (N_8147,N_7485,N_7364);
nand U8148 (N_8148,N_7253,N_7290);
nor U8149 (N_8149,N_7557,N_7903);
nand U8150 (N_8150,N_7806,N_7454);
or U8151 (N_8151,N_7382,N_7633);
nand U8152 (N_8152,N_7114,N_7921);
or U8153 (N_8153,N_7583,N_7124);
nand U8154 (N_8154,N_7049,N_7157);
or U8155 (N_8155,N_7656,N_7742);
nand U8156 (N_8156,N_7055,N_7233);
or U8157 (N_8157,N_7611,N_7177);
nor U8158 (N_8158,N_7207,N_7285);
xor U8159 (N_8159,N_7388,N_7304);
or U8160 (N_8160,N_7594,N_7723);
nor U8161 (N_8161,N_7365,N_7103);
nor U8162 (N_8162,N_7167,N_7435);
and U8163 (N_8163,N_7383,N_7521);
nand U8164 (N_8164,N_7010,N_7169);
nand U8165 (N_8165,N_7420,N_7272);
and U8166 (N_8166,N_7771,N_7257);
nand U8167 (N_8167,N_7936,N_7061);
nor U8168 (N_8168,N_7397,N_7994);
nor U8169 (N_8169,N_7700,N_7712);
nand U8170 (N_8170,N_7250,N_7882);
or U8171 (N_8171,N_7974,N_7821);
nor U8172 (N_8172,N_7526,N_7533);
or U8173 (N_8173,N_7793,N_7761);
or U8174 (N_8174,N_7243,N_7842);
and U8175 (N_8175,N_7444,N_7478);
or U8176 (N_8176,N_7105,N_7278);
and U8177 (N_8177,N_7205,N_7688);
or U8178 (N_8178,N_7053,N_7123);
or U8179 (N_8179,N_7500,N_7986);
nand U8180 (N_8180,N_7831,N_7523);
and U8181 (N_8181,N_7704,N_7620);
or U8182 (N_8182,N_7719,N_7495);
and U8183 (N_8183,N_7121,N_7823);
and U8184 (N_8184,N_7541,N_7489);
or U8185 (N_8185,N_7149,N_7664);
nand U8186 (N_8186,N_7640,N_7537);
or U8187 (N_8187,N_7969,N_7029);
nor U8188 (N_8188,N_7197,N_7369);
and U8189 (N_8189,N_7333,N_7101);
nand U8190 (N_8190,N_7987,N_7548);
nand U8191 (N_8191,N_7281,N_7294);
nand U8192 (N_8192,N_7768,N_7934);
nor U8193 (N_8193,N_7993,N_7573);
nor U8194 (N_8194,N_7196,N_7895);
nand U8195 (N_8195,N_7011,N_7330);
or U8196 (N_8196,N_7082,N_7957);
nor U8197 (N_8197,N_7219,N_7808);
nor U8198 (N_8198,N_7810,N_7824);
nor U8199 (N_8199,N_7552,N_7125);
nand U8200 (N_8200,N_7509,N_7033);
and U8201 (N_8201,N_7572,N_7461);
or U8202 (N_8202,N_7985,N_7091);
nand U8203 (N_8203,N_7711,N_7621);
nor U8204 (N_8204,N_7396,N_7142);
and U8205 (N_8205,N_7198,N_7905);
xnor U8206 (N_8206,N_7738,N_7422);
or U8207 (N_8207,N_7849,N_7991);
nand U8208 (N_8208,N_7327,N_7235);
nand U8209 (N_8209,N_7886,N_7171);
or U8210 (N_8210,N_7930,N_7608);
nor U8211 (N_8211,N_7596,N_7293);
and U8212 (N_8212,N_7455,N_7134);
or U8213 (N_8213,N_7491,N_7828);
or U8214 (N_8214,N_7152,N_7263);
nand U8215 (N_8215,N_7429,N_7052);
nor U8216 (N_8216,N_7023,N_7353);
nor U8217 (N_8217,N_7870,N_7778);
nand U8218 (N_8218,N_7059,N_7765);
nand U8219 (N_8219,N_7926,N_7858);
and U8220 (N_8220,N_7803,N_7757);
and U8221 (N_8221,N_7692,N_7020);
and U8222 (N_8222,N_7578,N_7232);
nand U8223 (N_8223,N_7266,N_7309);
nor U8224 (N_8224,N_7544,N_7789);
nor U8225 (N_8225,N_7256,N_7702);
or U8226 (N_8226,N_7662,N_7264);
nand U8227 (N_8227,N_7308,N_7137);
xnor U8228 (N_8228,N_7792,N_7518);
and U8229 (N_8229,N_7554,N_7414);
nand U8230 (N_8230,N_7861,N_7773);
xnor U8231 (N_8231,N_7856,N_7838);
or U8232 (N_8232,N_7822,N_7452);
nand U8233 (N_8233,N_7610,N_7075);
nand U8234 (N_8234,N_7678,N_7048);
and U8235 (N_8235,N_7160,N_7262);
nand U8236 (N_8236,N_7018,N_7958);
nor U8237 (N_8237,N_7909,N_7203);
nand U8238 (N_8238,N_7057,N_7570);
or U8239 (N_8239,N_7697,N_7876);
xor U8240 (N_8240,N_7952,N_7835);
or U8241 (N_8241,N_7585,N_7951);
or U8242 (N_8242,N_7054,N_7539);
nand U8243 (N_8243,N_7655,N_7317);
and U8244 (N_8244,N_7047,N_7534);
or U8245 (N_8245,N_7480,N_7911);
or U8246 (N_8246,N_7477,N_7244);
and U8247 (N_8247,N_7407,N_7222);
nor U8248 (N_8248,N_7445,N_7888);
and U8249 (N_8249,N_7282,N_7072);
nor U8250 (N_8250,N_7758,N_7216);
and U8251 (N_8251,N_7639,N_7691);
and U8252 (N_8252,N_7411,N_7260);
and U8253 (N_8253,N_7026,N_7163);
nor U8254 (N_8254,N_7967,N_7507);
and U8255 (N_8255,N_7535,N_7780);
nand U8256 (N_8256,N_7747,N_7258);
nand U8257 (N_8257,N_7805,N_7988);
and U8258 (N_8258,N_7790,N_7590);
nor U8259 (N_8259,N_7600,N_7796);
or U8260 (N_8260,N_7389,N_7668);
nand U8261 (N_8261,N_7374,N_7110);
or U8262 (N_8262,N_7013,N_7817);
nor U8263 (N_8263,N_7284,N_7943);
and U8264 (N_8264,N_7937,N_7553);
nor U8265 (N_8265,N_7440,N_7714);
nor U8266 (N_8266,N_7208,N_7944);
nor U8267 (N_8267,N_7751,N_7841);
nor U8268 (N_8268,N_7079,N_7653);
nand U8269 (N_8269,N_7246,N_7496);
and U8270 (N_8270,N_7226,N_7997);
nor U8271 (N_8271,N_7887,N_7532);
or U8272 (N_8272,N_7332,N_7112);
and U8273 (N_8273,N_7060,N_7941);
and U8274 (N_8274,N_7427,N_7400);
nand U8275 (N_8275,N_7069,N_7938);
nand U8276 (N_8276,N_7613,N_7146);
or U8277 (N_8277,N_7144,N_7223);
nand U8278 (N_8278,N_7775,N_7116);
or U8279 (N_8279,N_7398,N_7056);
and U8280 (N_8280,N_7183,N_7820);
and U8281 (N_8281,N_7497,N_7184);
and U8282 (N_8282,N_7459,N_7307);
nand U8283 (N_8283,N_7525,N_7892);
or U8284 (N_8284,N_7850,N_7933);
nand U8285 (N_8285,N_7321,N_7899);
and U8286 (N_8286,N_7536,N_7395);
nor U8287 (N_8287,N_7437,N_7501);
or U8288 (N_8288,N_7001,N_7348);
nand U8289 (N_8289,N_7224,N_7603);
nand U8290 (N_8290,N_7254,N_7927);
nor U8291 (N_8291,N_7660,N_7737);
and U8292 (N_8292,N_7772,N_7760);
nand U8293 (N_8293,N_7642,N_7898);
nor U8294 (N_8294,N_7273,N_7063);
or U8295 (N_8295,N_7609,N_7351);
and U8296 (N_8296,N_7415,N_7034);
and U8297 (N_8297,N_7917,N_7466);
and U8298 (N_8298,N_7115,N_7297);
nor U8299 (N_8299,N_7669,N_7995);
nor U8300 (N_8300,N_7686,N_7667);
nand U8301 (N_8301,N_7481,N_7098);
nor U8302 (N_8302,N_7925,N_7568);
nor U8303 (N_8303,N_7953,N_7376);
and U8304 (N_8304,N_7326,N_7117);
nor U8305 (N_8305,N_7009,N_7493);
nor U8306 (N_8306,N_7918,N_7902);
and U8307 (N_8307,N_7617,N_7624);
nand U8308 (N_8308,N_7961,N_7426);
or U8309 (N_8309,N_7410,N_7385);
nor U8310 (N_8310,N_7843,N_7979);
nor U8311 (N_8311,N_7090,N_7579);
and U8312 (N_8312,N_7071,N_7645);
nand U8313 (N_8313,N_7576,N_7650);
and U8314 (N_8314,N_7785,N_7718);
nand U8315 (N_8315,N_7367,N_7689);
and U8316 (N_8316,N_7259,N_7542);
nor U8317 (N_8317,N_7000,N_7646);
or U8318 (N_8318,N_7499,N_7153);
or U8319 (N_8319,N_7912,N_7180);
xnor U8320 (N_8320,N_7068,N_7287);
nor U8321 (N_8321,N_7844,N_7251);
and U8322 (N_8322,N_7784,N_7913);
and U8323 (N_8323,N_7588,N_7355);
nand U8324 (N_8324,N_7039,N_7595);
or U8325 (N_8325,N_7030,N_7942);
nor U8326 (N_8326,N_7314,N_7571);
nand U8327 (N_8327,N_7800,N_7472);
and U8328 (N_8328,N_7100,N_7042);
nor U8329 (N_8329,N_7659,N_7649);
and U8330 (N_8330,N_7214,N_7156);
nand U8331 (N_8331,N_7473,N_7405);
or U8332 (N_8332,N_7631,N_7460);
or U8333 (N_8333,N_7486,N_7754);
or U8334 (N_8334,N_7770,N_7119);
nor U8335 (N_8335,N_7476,N_7730);
and U8336 (N_8336,N_7530,N_7735);
nor U8337 (N_8337,N_7563,N_7202);
and U8338 (N_8338,N_7940,N_7783);
nor U8339 (N_8339,N_7731,N_7099);
xor U8340 (N_8340,N_7514,N_7448);
nor U8341 (N_8341,N_7217,N_7181);
nand U8342 (N_8342,N_7960,N_7891);
and U8343 (N_8343,N_7113,N_7096);
or U8344 (N_8344,N_7782,N_7559);
nand U8345 (N_8345,N_7605,N_7270);
and U8346 (N_8346,N_7612,N_7740);
or U8347 (N_8347,N_7458,N_7607);
nor U8348 (N_8348,N_7932,N_7446);
or U8349 (N_8349,N_7699,N_7025);
or U8350 (N_8350,N_7038,N_7462);
nor U8351 (N_8351,N_7696,N_7432);
nor U8352 (N_8352,N_7106,N_7469);
nor U8353 (N_8353,N_7565,N_7252);
nor U8354 (N_8354,N_7339,N_7036);
or U8355 (N_8355,N_7807,N_7619);
and U8356 (N_8356,N_7236,N_7316);
nand U8357 (N_8357,N_7854,N_7592);
nor U8358 (N_8358,N_7482,N_7949);
or U8359 (N_8359,N_7296,N_7992);
nor U8360 (N_8360,N_7845,N_7331);
or U8361 (N_8361,N_7685,N_7185);
nand U8362 (N_8362,N_7589,N_7136);
or U8363 (N_8363,N_7248,N_7863);
nor U8364 (N_8364,N_7638,N_7301);
nor U8365 (N_8365,N_7391,N_7417);
nor U8366 (N_8366,N_7663,N_7092);
xor U8367 (N_8367,N_7081,N_7733);
and U8368 (N_8368,N_7088,N_7265);
nor U8369 (N_8369,N_7211,N_7690);
and U8370 (N_8370,N_7418,N_7581);
nor U8371 (N_8371,N_7543,N_7172);
or U8372 (N_8372,N_7138,N_7703);
nand U8373 (N_8373,N_7666,N_7392);
nand U8374 (N_8374,N_7971,N_7412);
nor U8375 (N_8375,N_7764,N_7237);
or U8376 (N_8376,N_7401,N_7928);
nor U8377 (N_8377,N_7324,N_7450);
or U8378 (N_8378,N_7508,N_7989);
or U8379 (N_8379,N_7127,N_7878);
and U8380 (N_8380,N_7819,N_7209);
nand U8381 (N_8381,N_7002,N_7210);
nand U8382 (N_8382,N_7540,N_7231);
nor U8383 (N_8383,N_7745,N_7558);
and U8384 (N_8384,N_7277,N_7494);
xnor U8385 (N_8385,N_7338,N_7982);
and U8386 (N_8386,N_7632,N_7955);
nor U8387 (N_8387,N_7457,N_7276);
xnor U8388 (N_8388,N_7948,N_7857);
nand U8389 (N_8389,N_7709,N_7070);
nor U8390 (N_8390,N_7677,N_7492);
or U8391 (N_8391,N_7871,N_7008);
or U8392 (N_8392,N_7866,N_7865);
nor U8393 (N_8393,N_7404,N_7924);
nand U8394 (N_8394,N_7716,N_7715);
nor U8395 (N_8395,N_7017,N_7591);
or U8396 (N_8396,N_7436,N_7970);
xor U8397 (N_8397,N_7463,N_7623);
nand U8398 (N_8398,N_7837,N_7734);
nor U8399 (N_8399,N_7150,N_7520);
and U8400 (N_8400,N_7132,N_7577);
and U8401 (N_8401,N_7245,N_7064);
nand U8402 (N_8402,N_7728,N_7089);
and U8403 (N_8403,N_7228,N_7883);
or U8404 (N_8404,N_7658,N_7812);
and U8405 (N_8405,N_7794,N_7549);
or U8406 (N_8406,N_7674,N_7695);
or U8407 (N_8407,N_7074,N_7746);
and U8408 (N_8408,N_7732,N_7998);
nand U8409 (N_8409,N_7201,N_7561);
and U8410 (N_8410,N_7286,N_7832);
or U8411 (N_8411,N_7964,N_7268);
nand U8412 (N_8412,N_7825,N_7683);
nor U8413 (N_8413,N_7044,N_7804);
or U8414 (N_8414,N_7051,N_7199);
or U8415 (N_8415,N_7394,N_7187);
or U8416 (N_8416,N_7618,N_7345);
and U8417 (N_8417,N_7705,N_7359);
or U8418 (N_8418,N_7859,N_7045);
nand U8419 (N_8419,N_7122,N_7456);
nand U8420 (N_8420,N_7421,N_7174);
nor U8421 (N_8421,N_7929,N_7164);
or U8422 (N_8422,N_7043,N_7852);
or U8423 (N_8423,N_7914,N_7085);
nor U8424 (N_8424,N_7155,N_7413);
nand U8425 (N_8425,N_7965,N_7191);
and U8426 (N_8426,N_7024,N_7682);
nor U8427 (N_8427,N_7885,N_7451);
nor U8428 (N_8428,N_7574,N_7815);
nand U8429 (N_8429,N_7484,N_7131);
nand U8430 (N_8430,N_7443,N_7907);
or U8431 (N_8431,N_7884,N_7922);
nor U8432 (N_8432,N_7504,N_7453);
and U8433 (N_8433,N_7795,N_7963);
xor U8434 (N_8434,N_7292,N_7488);
nor U8435 (N_8435,N_7419,N_7769);
xnor U8436 (N_8436,N_7386,N_7140);
or U8437 (N_8437,N_7004,N_7108);
nand U8438 (N_8438,N_7867,N_7586);
nand U8439 (N_8439,N_7159,N_7774);
and U8440 (N_8440,N_7428,N_7192);
nand U8441 (N_8441,N_7946,N_7901);
or U8442 (N_8442,N_7016,N_7234);
or U8443 (N_8443,N_7465,N_7698);
and U8444 (N_8444,N_7615,N_7238);
nand U8445 (N_8445,N_7799,N_7724);
and U8446 (N_8446,N_7981,N_7766);
and U8447 (N_8447,N_7111,N_7213);
nand U8448 (N_8448,N_7315,N_7175);
and U8449 (N_8449,N_7399,N_7904);
nand U8450 (N_8450,N_7487,N_7084);
xnor U8451 (N_8451,N_7360,N_7671);
or U8452 (N_8452,N_7408,N_7962);
and U8453 (N_8453,N_7634,N_7727);
and U8454 (N_8454,N_7283,N_7438);
or U8455 (N_8455,N_7830,N_7720);
or U8456 (N_8456,N_7661,N_7968);
nor U8457 (N_8457,N_7897,N_7247);
nand U8458 (N_8458,N_7046,N_7379);
and U8459 (N_8459,N_7468,N_7670);
and U8460 (N_8460,N_7529,N_7681);
or U8461 (N_8461,N_7788,N_7019);
nand U8462 (N_8462,N_7524,N_7575);
and U8463 (N_8463,N_7241,N_7006);
or U8464 (N_8464,N_7947,N_7546);
nand U8465 (N_8465,N_7350,N_7190);
nand U8466 (N_8466,N_7900,N_7299);
and U8467 (N_8467,N_7135,N_7721);
nand U8468 (N_8468,N_7813,N_7380);
and U8469 (N_8469,N_7672,N_7434);
xor U8470 (N_8470,N_7814,N_7423);
or U8471 (N_8471,N_7363,N_7143);
or U8472 (N_8472,N_7298,N_7107);
nand U8473 (N_8473,N_7483,N_7300);
nand U8474 (N_8474,N_7346,N_7178);
or U8475 (N_8475,N_7750,N_7906);
nor U8476 (N_8476,N_7869,N_7126);
or U8477 (N_8477,N_7516,N_7498);
or U8478 (N_8478,N_7341,N_7802);
nor U8479 (N_8479,N_7148,N_7555);
and U8480 (N_8480,N_7776,N_7593);
nor U8481 (N_8481,N_7860,N_7065);
nor U8482 (N_8482,N_7170,N_7545);
or U8483 (N_8483,N_7162,N_7527);
and U8484 (N_8484,N_7239,N_7580);
or U8485 (N_8485,N_7007,N_7630);
and U8486 (N_8486,N_7881,N_7182);
nor U8487 (N_8487,N_7028,N_7206);
nand U8488 (N_8488,N_7474,N_7368);
xor U8489 (N_8489,N_7189,N_7567);
nand U8490 (N_8490,N_7847,N_7864);
nor U8491 (N_8491,N_7959,N_7403);
nor U8492 (N_8492,N_7977,N_7280);
nor U8493 (N_8493,N_7975,N_7220);
and U8494 (N_8494,N_7950,N_7694);
nand U8495 (N_8495,N_7021,N_7005);
nand U8496 (N_8496,N_7625,N_7193);
or U8497 (N_8497,N_7361,N_7569);
nand U8498 (N_8498,N_7873,N_7154);
and U8499 (N_8499,N_7862,N_7186);
nor U8500 (N_8500,N_7117,N_7667);
nand U8501 (N_8501,N_7672,N_7952);
and U8502 (N_8502,N_7904,N_7996);
or U8503 (N_8503,N_7559,N_7726);
nor U8504 (N_8504,N_7896,N_7658);
nand U8505 (N_8505,N_7570,N_7856);
and U8506 (N_8506,N_7890,N_7342);
nand U8507 (N_8507,N_7322,N_7600);
nand U8508 (N_8508,N_7710,N_7286);
or U8509 (N_8509,N_7497,N_7043);
nor U8510 (N_8510,N_7754,N_7708);
or U8511 (N_8511,N_7278,N_7810);
nor U8512 (N_8512,N_7456,N_7772);
or U8513 (N_8513,N_7179,N_7998);
and U8514 (N_8514,N_7719,N_7859);
or U8515 (N_8515,N_7909,N_7308);
nor U8516 (N_8516,N_7296,N_7436);
or U8517 (N_8517,N_7084,N_7631);
nand U8518 (N_8518,N_7048,N_7007);
and U8519 (N_8519,N_7705,N_7037);
and U8520 (N_8520,N_7844,N_7041);
nand U8521 (N_8521,N_7948,N_7459);
nor U8522 (N_8522,N_7796,N_7588);
and U8523 (N_8523,N_7035,N_7177);
and U8524 (N_8524,N_7131,N_7825);
nor U8525 (N_8525,N_7941,N_7163);
nor U8526 (N_8526,N_7977,N_7655);
and U8527 (N_8527,N_7763,N_7196);
nor U8528 (N_8528,N_7803,N_7242);
and U8529 (N_8529,N_7503,N_7834);
or U8530 (N_8530,N_7193,N_7273);
or U8531 (N_8531,N_7622,N_7373);
nor U8532 (N_8532,N_7635,N_7738);
nand U8533 (N_8533,N_7659,N_7473);
or U8534 (N_8534,N_7281,N_7541);
and U8535 (N_8535,N_7673,N_7664);
and U8536 (N_8536,N_7213,N_7229);
or U8537 (N_8537,N_7775,N_7895);
nand U8538 (N_8538,N_7861,N_7456);
and U8539 (N_8539,N_7179,N_7423);
and U8540 (N_8540,N_7106,N_7844);
nand U8541 (N_8541,N_7131,N_7976);
nand U8542 (N_8542,N_7777,N_7497);
and U8543 (N_8543,N_7341,N_7711);
and U8544 (N_8544,N_7006,N_7854);
nand U8545 (N_8545,N_7756,N_7430);
nor U8546 (N_8546,N_7397,N_7973);
nand U8547 (N_8547,N_7583,N_7263);
nor U8548 (N_8548,N_7158,N_7051);
nand U8549 (N_8549,N_7587,N_7579);
and U8550 (N_8550,N_7304,N_7631);
and U8551 (N_8551,N_7606,N_7231);
nand U8552 (N_8552,N_7550,N_7916);
and U8553 (N_8553,N_7933,N_7107);
nand U8554 (N_8554,N_7696,N_7578);
or U8555 (N_8555,N_7997,N_7627);
or U8556 (N_8556,N_7938,N_7866);
nor U8557 (N_8557,N_7873,N_7674);
or U8558 (N_8558,N_7930,N_7887);
or U8559 (N_8559,N_7424,N_7777);
or U8560 (N_8560,N_7425,N_7872);
nor U8561 (N_8561,N_7329,N_7205);
nor U8562 (N_8562,N_7956,N_7093);
and U8563 (N_8563,N_7403,N_7291);
or U8564 (N_8564,N_7545,N_7878);
or U8565 (N_8565,N_7495,N_7984);
and U8566 (N_8566,N_7963,N_7567);
and U8567 (N_8567,N_7075,N_7698);
or U8568 (N_8568,N_7536,N_7967);
and U8569 (N_8569,N_7935,N_7260);
nor U8570 (N_8570,N_7458,N_7814);
nor U8571 (N_8571,N_7258,N_7787);
nand U8572 (N_8572,N_7037,N_7701);
nand U8573 (N_8573,N_7793,N_7716);
or U8574 (N_8574,N_7717,N_7530);
nand U8575 (N_8575,N_7318,N_7459);
or U8576 (N_8576,N_7687,N_7666);
nand U8577 (N_8577,N_7533,N_7687);
xor U8578 (N_8578,N_7502,N_7010);
nor U8579 (N_8579,N_7415,N_7914);
nor U8580 (N_8580,N_7266,N_7994);
and U8581 (N_8581,N_7001,N_7580);
nor U8582 (N_8582,N_7552,N_7372);
and U8583 (N_8583,N_7704,N_7659);
nor U8584 (N_8584,N_7163,N_7400);
nor U8585 (N_8585,N_7642,N_7401);
xor U8586 (N_8586,N_7846,N_7553);
and U8587 (N_8587,N_7514,N_7009);
or U8588 (N_8588,N_7306,N_7154);
nand U8589 (N_8589,N_7153,N_7515);
or U8590 (N_8590,N_7666,N_7866);
or U8591 (N_8591,N_7215,N_7672);
nor U8592 (N_8592,N_7345,N_7131);
nand U8593 (N_8593,N_7299,N_7351);
nand U8594 (N_8594,N_7887,N_7209);
nor U8595 (N_8595,N_7904,N_7461);
xor U8596 (N_8596,N_7627,N_7394);
nand U8597 (N_8597,N_7769,N_7739);
nand U8598 (N_8598,N_7716,N_7511);
nor U8599 (N_8599,N_7825,N_7185);
nor U8600 (N_8600,N_7530,N_7056);
nor U8601 (N_8601,N_7811,N_7696);
nor U8602 (N_8602,N_7101,N_7611);
and U8603 (N_8603,N_7720,N_7766);
nor U8604 (N_8604,N_7003,N_7782);
and U8605 (N_8605,N_7854,N_7876);
or U8606 (N_8606,N_7181,N_7777);
nand U8607 (N_8607,N_7922,N_7481);
and U8608 (N_8608,N_7805,N_7047);
and U8609 (N_8609,N_7882,N_7754);
or U8610 (N_8610,N_7901,N_7601);
nor U8611 (N_8611,N_7466,N_7170);
nor U8612 (N_8612,N_7826,N_7113);
nor U8613 (N_8613,N_7183,N_7198);
nand U8614 (N_8614,N_7186,N_7824);
nor U8615 (N_8615,N_7617,N_7174);
or U8616 (N_8616,N_7676,N_7261);
or U8617 (N_8617,N_7723,N_7973);
nor U8618 (N_8618,N_7571,N_7823);
nand U8619 (N_8619,N_7720,N_7150);
nand U8620 (N_8620,N_7974,N_7645);
nor U8621 (N_8621,N_7358,N_7623);
and U8622 (N_8622,N_7296,N_7974);
nand U8623 (N_8623,N_7276,N_7327);
or U8624 (N_8624,N_7836,N_7049);
nand U8625 (N_8625,N_7734,N_7752);
nor U8626 (N_8626,N_7131,N_7731);
nand U8627 (N_8627,N_7717,N_7900);
or U8628 (N_8628,N_7988,N_7885);
nor U8629 (N_8629,N_7037,N_7435);
nand U8630 (N_8630,N_7700,N_7959);
and U8631 (N_8631,N_7195,N_7283);
nand U8632 (N_8632,N_7379,N_7821);
nand U8633 (N_8633,N_7818,N_7606);
or U8634 (N_8634,N_7812,N_7758);
nand U8635 (N_8635,N_7013,N_7128);
and U8636 (N_8636,N_7532,N_7583);
nor U8637 (N_8637,N_7565,N_7842);
and U8638 (N_8638,N_7728,N_7634);
nor U8639 (N_8639,N_7613,N_7136);
or U8640 (N_8640,N_7640,N_7591);
or U8641 (N_8641,N_7762,N_7304);
and U8642 (N_8642,N_7884,N_7439);
and U8643 (N_8643,N_7190,N_7979);
or U8644 (N_8644,N_7753,N_7299);
nand U8645 (N_8645,N_7202,N_7999);
nor U8646 (N_8646,N_7226,N_7471);
or U8647 (N_8647,N_7629,N_7051);
and U8648 (N_8648,N_7304,N_7010);
nand U8649 (N_8649,N_7507,N_7947);
nor U8650 (N_8650,N_7865,N_7664);
and U8651 (N_8651,N_7430,N_7935);
and U8652 (N_8652,N_7738,N_7772);
or U8653 (N_8653,N_7491,N_7227);
nor U8654 (N_8654,N_7153,N_7801);
or U8655 (N_8655,N_7428,N_7032);
or U8656 (N_8656,N_7294,N_7012);
nand U8657 (N_8657,N_7401,N_7890);
and U8658 (N_8658,N_7222,N_7580);
and U8659 (N_8659,N_7024,N_7334);
and U8660 (N_8660,N_7960,N_7140);
or U8661 (N_8661,N_7996,N_7927);
and U8662 (N_8662,N_7651,N_7838);
or U8663 (N_8663,N_7919,N_7915);
or U8664 (N_8664,N_7734,N_7295);
or U8665 (N_8665,N_7925,N_7183);
nand U8666 (N_8666,N_7704,N_7463);
nor U8667 (N_8667,N_7373,N_7530);
or U8668 (N_8668,N_7664,N_7759);
nor U8669 (N_8669,N_7847,N_7853);
and U8670 (N_8670,N_7964,N_7230);
or U8671 (N_8671,N_7701,N_7429);
nand U8672 (N_8672,N_7193,N_7610);
and U8673 (N_8673,N_7543,N_7726);
nand U8674 (N_8674,N_7147,N_7376);
and U8675 (N_8675,N_7696,N_7838);
nor U8676 (N_8676,N_7446,N_7658);
or U8677 (N_8677,N_7253,N_7936);
xnor U8678 (N_8678,N_7130,N_7396);
or U8679 (N_8679,N_7232,N_7136);
nor U8680 (N_8680,N_7111,N_7110);
nor U8681 (N_8681,N_7587,N_7121);
nand U8682 (N_8682,N_7627,N_7327);
nor U8683 (N_8683,N_7376,N_7948);
and U8684 (N_8684,N_7412,N_7147);
nor U8685 (N_8685,N_7624,N_7031);
xnor U8686 (N_8686,N_7390,N_7171);
nand U8687 (N_8687,N_7532,N_7747);
or U8688 (N_8688,N_7902,N_7004);
nand U8689 (N_8689,N_7720,N_7467);
or U8690 (N_8690,N_7780,N_7634);
or U8691 (N_8691,N_7467,N_7123);
and U8692 (N_8692,N_7862,N_7184);
or U8693 (N_8693,N_7060,N_7112);
and U8694 (N_8694,N_7640,N_7610);
and U8695 (N_8695,N_7271,N_7392);
xor U8696 (N_8696,N_7245,N_7618);
or U8697 (N_8697,N_7054,N_7909);
nor U8698 (N_8698,N_7892,N_7798);
nor U8699 (N_8699,N_7917,N_7011);
nand U8700 (N_8700,N_7699,N_7787);
nor U8701 (N_8701,N_7135,N_7956);
xnor U8702 (N_8702,N_7723,N_7950);
nor U8703 (N_8703,N_7367,N_7138);
or U8704 (N_8704,N_7878,N_7222);
and U8705 (N_8705,N_7662,N_7096);
nand U8706 (N_8706,N_7518,N_7505);
xnor U8707 (N_8707,N_7917,N_7985);
nor U8708 (N_8708,N_7821,N_7983);
and U8709 (N_8709,N_7361,N_7896);
nor U8710 (N_8710,N_7635,N_7450);
and U8711 (N_8711,N_7741,N_7001);
or U8712 (N_8712,N_7180,N_7733);
or U8713 (N_8713,N_7602,N_7385);
nand U8714 (N_8714,N_7794,N_7504);
or U8715 (N_8715,N_7437,N_7439);
xor U8716 (N_8716,N_7691,N_7210);
or U8717 (N_8717,N_7138,N_7882);
or U8718 (N_8718,N_7775,N_7308);
nand U8719 (N_8719,N_7069,N_7685);
or U8720 (N_8720,N_7017,N_7618);
nand U8721 (N_8721,N_7147,N_7434);
and U8722 (N_8722,N_7129,N_7044);
and U8723 (N_8723,N_7465,N_7873);
nand U8724 (N_8724,N_7308,N_7147);
nor U8725 (N_8725,N_7494,N_7379);
or U8726 (N_8726,N_7654,N_7456);
or U8727 (N_8727,N_7255,N_7586);
and U8728 (N_8728,N_7083,N_7791);
and U8729 (N_8729,N_7808,N_7544);
nand U8730 (N_8730,N_7528,N_7304);
and U8731 (N_8731,N_7202,N_7415);
nor U8732 (N_8732,N_7929,N_7938);
or U8733 (N_8733,N_7740,N_7819);
nand U8734 (N_8734,N_7538,N_7605);
or U8735 (N_8735,N_7932,N_7674);
or U8736 (N_8736,N_7232,N_7997);
nand U8737 (N_8737,N_7372,N_7821);
nor U8738 (N_8738,N_7900,N_7770);
nor U8739 (N_8739,N_7123,N_7286);
or U8740 (N_8740,N_7668,N_7155);
or U8741 (N_8741,N_7579,N_7896);
or U8742 (N_8742,N_7532,N_7163);
nand U8743 (N_8743,N_7470,N_7484);
nor U8744 (N_8744,N_7826,N_7877);
nor U8745 (N_8745,N_7704,N_7173);
and U8746 (N_8746,N_7084,N_7329);
nand U8747 (N_8747,N_7901,N_7109);
and U8748 (N_8748,N_7938,N_7559);
or U8749 (N_8749,N_7163,N_7887);
or U8750 (N_8750,N_7449,N_7859);
nor U8751 (N_8751,N_7943,N_7618);
nand U8752 (N_8752,N_7922,N_7525);
and U8753 (N_8753,N_7539,N_7422);
and U8754 (N_8754,N_7596,N_7814);
nor U8755 (N_8755,N_7302,N_7538);
nand U8756 (N_8756,N_7003,N_7685);
nor U8757 (N_8757,N_7759,N_7162);
and U8758 (N_8758,N_7098,N_7461);
nand U8759 (N_8759,N_7049,N_7258);
or U8760 (N_8760,N_7785,N_7873);
or U8761 (N_8761,N_7167,N_7580);
or U8762 (N_8762,N_7234,N_7063);
and U8763 (N_8763,N_7843,N_7780);
nand U8764 (N_8764,N_7349,N_7665);
and U8765 (N_8765,N_7848,N_7990);
and U8766 (N_8766,N_7749,N_7145);
nand U8767 (N_8767,N_7596,N_7363);
nor U8768 (N_8768,N_7366,N_7211);
or U8769 (N_8769,N_7393,N_7550);
nand U8770 (N_8770,N_7458,N_7517);
nand U8771 (N_8771,N_7283,N_7583);
or U8772 (N_8772,N_7915,N_7714);
or U8773 (N_8773,N_7326,N_7181);
nand U8774 (N_8774,N_7516,N_7229);
or U8775 (N_8775,N_7784,N_7874);
nor U8776 (N_8776,N_7692,N_7961);
or U8777 (N_8777,N_7161,N_7875);
or U8778 (N_8778,N_7168,N_7669);
nand U8779 (N_8779,N_7275,N_7494);
and U8780 (N_8780,N_7217,N_7312);
nand U8781 (N_8781,N_7895,N_7684);
nand U8782 (N_8782,N_7281,N_7880);
and U8783 (N_8783,N_7034,N_7530);
or U8784 (N_8784,N_7112,N_7758);
or U8785 (N_8785,N_7405,N_7648);
and U8786 (N_8786,N_7177,N_7968);
nor U8787 (N_8787,N_7026,N_7082);
nand U8788 (N_8788,N_7925,N_7590);
or U8789 (N_8789,N_7502,N_7851);
and U8790 (N_8790,N_7558,N_7895);
nor U8791 (N_8791,N_7218,N_7729);
nor U8792 (N_8792,N_7083,N_7980);
nand U8793 (N_8793,N_7664,N_7288);
nand U8794 (N_8794,N_7085,N_7011);
nand U8795 (N_8795,N_7092,N_7983);
nor U8796 (N_8796,N_7844,N_7734);
or U8797 (N_8797,N_7975,N_7948);
xnor U8798 (N_8798,N_7991,N_7422);
xor U8799 (N_8799,N_7414,N_7476);
xnor U8800 (N_8800,N_7661,N_7808);
nand U8801 (N_8801,N_7036,N_7443);
xor U8802 (N_8802,N_7018,N_7415);
nand U8803 (N_8803,N_7431,N_7574);
or U8804 (N_8804,N_7038,N_7315);
nor U8805 (N_8805,N_7219,N_7377);
or U8806 (N_8806,N_7943,N_7364);
or U8807 (N_8807,N_7728,N_7545);
and U8808 (N_8808,N_7053,N_7727);
and U8809 (N_8809,N_7687,N_7595);
and U8810 (N_8810,N_7265,N_7232);
or U8811 (N_8811,N_7651,N_7861);
and U8812 (N_8812,N_7135,N_7366);
and U8813 (N_8813,N_7027,N_7296);
nor U8814 (N_8814,N_7359,N_7100);
or U8815 (N_8815,N_7282,N_7335);
and U8816 (N_8816,N_7782,N_7313);
and U8817 (N_8817,N_7488,N_7679);
nand U8818 (N_8818,N_7110,N_7853);
nor U8819 (N_8819,N_7840,N_7081);
or U8820 (N_8820,N_7949,N_7200);
or U8821 (N_8821,N_7429,N_7771);
nand U8822 (N_8822,N_7218,N_7151);
nor U8823 (N_8823,N_7256,N_7222);
or U8824 (N_8824,N_7766,N_7738);
nor U8825 (N_8825,N_7418,N_7409);
nor U8826 (N_8826,N_7369,N_7875);
and U8827 (N_8827,N_7425,N_7611);
nand U8828 (N_8828,N_7905,N_7144);
nand U8829 (N_8829,N_7436,N_7916);
nor U8830 (N_8830,N_7999,N_7105);
nand U8831 (N_8831,N_7358,N_7648);
nand U8832 (N_8832,N_7597,N_7257);
nor U8833 (N_8833,N_7295,N_7906);
nor U8834 (N_8834,N_7715,N_7969);
xnor U8835 (N_8835,N_7421,N_7853);
nand U8836 (N_8836,N_7663,N_7378);
nand U8837 (N_8837,N_7574,N_7135);
and U8838 (N_8838,N_7622,N_7266);
nand U8839 (N_8839,N_7314,N_7179);
or U8840 (N_8840,N_7670,N_7333);
nor U8841 (N_8841,N_7371,N_7565);
xnor U8842 (N_8842,N_7692,N_7205);
xor U8843 (N_8843,N_7042,N_7750);
nor U8844 (N_8844,N_7839,N_7162);
nor U8845 (N_8845,N_7012,N_7597);
nand U8846 (N_8846,N_7869,N_7611);
or U8847 (N_8847,N_7365,N_7769);
or U8848 (N_8848,N_7226,N_7258);
nor U8849 (N_8849,N_7940,N_7788);
nand U8850 (N_8850,N_7652,N_7565);
xor U8851 (N_8851,N_7780,N_7552);
nand U8852 (N_8852,N_7869,N_7298);
nand U8853 (N_8853,N_7680,N_7228);
nand U8854 (N_8854,N_7520,N_7219);
nor U8855 (N_8855,N_7619,N_7778);
nand U8856 (N_8856,N_7174,N_7509);
nand U8857 (N_8857,N_7652,N_7980);
or U8858 (N_8858,N_7836,N_7350);
or U8859 (N_8859,N_7071,N_7058);
or U8860 (N_8860,N_7560,N_7558);
nand U8861 (N_8861,N_7413,N_7365);
or U8862 (N_8862,N_7152,N_7339);
nor U8863 (N_8863,N_7989,N_7024);
or U8864 (N_8864,N_7977,N_7854);
and U8865 (N_8865,N_7121,N_7661);
and U8866 (N_8866,N_7506,N_7735);
nand U8867 (N_8867,N_7062,N_7515);
nor U8868 (N_8868,N_7362,N_7801);
nor U8869 (N_8869,N_7157,N_7262);
nand U8870 (N_8870,N_7843,N_7317);
and U8871 (N_8871,N_7845,N_7392);
nand U8872 (N_8872,N_7776,N_7242);
or U8873 (N_8873,N_7608,N_7140);
nor U8874 (N_8874,N_7619,N_7184);
nor U8875 (N_8875,N_7226,N_7137);
nand U8876 (N_8876,N_7657,N_7900);
or U8877 (N_8877,N_7886,N_7851);
and U8878 (N_8878,N_7434,N_7184);
and U8879 (N_8879,N_7961,N_7994);
nor U8880 (N_8880,N_7105,N_7275);
nand U8881 (N_8881,N_7545,N_7654);
nor U8882 (N_8882,N_7041,N_7584);
nand U8883 (N_8883,N_7063,N_7073);
or U8884 (N_8884,N_7242,N_7493);
and U8885 (N_8885,N_7113,N_7584);
nand U8886 (N_8886,N_7101,N_7222);
nand U8887 (N_8887,N_7781,N_7063);
or U8888 (N_8888,N_7901,N_7645);
nor U8889 (N_8889,N_7168,N_7760);
nor U8890 (N_8890,N_7311,N_7352);
nor U8891 (N_8891,N_7010,N_7847);
and U8892 (N_8892,N_7139,N_7934);
or U8893 (N_8893,N_7420,N_7569);
nor U8894 (N_8894,N_7174,N_7196);
nor U8895 (N_8895,N_7202,N_7359);
or U8896 (N_8896,N_7410,N_7447);
nor U8897 (N_8897,N_7592,N_7661);
nor U8898 (N_8898,N_7422,N_7853);
nor U8899 (N_8899,N_7296,N_7635);
nand U8900 (N_8900,N_7091,N_7377);
or U8901 (N_8901,N_7021,N_7814);
nor U8902 (N_8902,N_7990,N_7546);
or U8903 (N_8903,N_7358,N_7562);
nand U8904 (N_8904,N_7869,N_7007);
and U8905 (N_8905,N_7795,N_7085);
and U8906 (N_8906,N_7095,N_7911);
or U8907 (N_8907,N_7162,N_7211);
nor U8908 (N_8908,N_7082,N_7055);
nor U8909 (N_8909,N_7192,N_7900);
or U8910 (N_8910,N_7951,N_7737);
and U8911 (N_8911,N_7491,N_7521);
nor U8912 (N_8912,N_7079,N_7119);
nor U8913 (N_8913,N_7785,N_7104);
or U8914 (N_8914,N_7472,N_7206);
or U8915 (N_8915,N_7112,N_7212);
or U8916 (N_8916,N_7847,N_7988);
nand U8917 (N_8917,N_7282,N_7076);
nor U8918 (N_8918,N_7886,N_7920);
or U8919 (N_8919,N_7299,N_7962);
or U8920 (N_8920,N_7596,N_7700);
or U8921 (N_8921,N_7225,N_7231);
and U8922 (N_8922,N_7745,N_7309);
or U8923 (N_8923,N_7785,N_7944);
nor U8924 (N_8924,N_7165,N_7114);
nor U8925 (N_8925,N_7126,N_7248);
and U8926 (N_8926,N_7343,N_7643);
nand U8927 (N_8927,N_7722,N_7670);
or U8928 (N_8928,N_7104,N_7320);
nand U8929 (N_8929,N_7324,N_7035);
nor U8930 (N_8930,N_7044,N_7713);
and U8931 (N_8931,N_7834,N_7094);
nand U8932 (N_8932,N_7412,N_7132);
nand U8933 (N_8933,N_7286,N_7243);
and U8934 (N_8934,N_7159,N_7470);
and U8935 (N_8935,N_7767,N_7244);
nand U8936 (N_8936,N_7850,N_7993);
nand U8937 (N_8937,N_7237,N_7960);
nand U8938 (N_8938,N_7984,N_7884);
or U8939 (N_8939,N_7562,N_7812);
nand U8940 (N_8940,N_7726,N_7778);
nor U8941 (N_8941,N_7452,N_7999);
nor U8942 (N_8942,N_7523,N_7455);
and U8943 (N_8943,N_7748,N_7094);
or U8944 (N_8944,N_7897,N_7861);
nand U8945 (N_8945,N_7949,N_7456);
and U8946 (N_8946,N_7457,N_7161);
nand U8947 (N_8947,N_7307,N_7183);
and U8948 (N_8948,N_7888,N_7621);
nand U8949 (N_8949,N_7450,N_7347);
nor U8950 (N_8950,N_7302,N_7608);
nor U8951 (N_8951,N_7273,N_7616);
and U8952 (N_8952,N_7108,N_7315);
nand U8953 (N_8953,N_7299,N_7583);
or U8954 (N_8954,N_7296,N_7294);
and U8955 (N_8955,N_7379,N_7286);
nand U8956 (N_8956,N_7953,N_7306);
nand U8957 (N_8957,N_7606,N_7167);
xnor U8958 (N_8958,N_7626,N_7281);
nand U8959 (N_8959,N_7022,N_7693);
nand U8960 (N_8960,N_7498,N_7250);
nand U8961 (N_8961,N_7100,N_7781);
or U8962 (N_8962,N_7820,N_7388);
nand U8963 (N_8963,N_7012,N_7353);
nor U8964 (N_8964,N_7261,N_7271);
or U8965 (N_8965,N_7010,N_7680);
nor U8966 (N_8966,N_7994,N_7850);
nor U8967 (N_8967,N_7147,N_7691);
nand U8968 (N_8968,N_7875,N_7837);
xnor U8969 (N_8969,N_7182,N_7602);
nor U8970 (N_8970,N_7895,N_7027);
nor U8971 (N_8971,N_7880,N_7206);
and U8972 (N_8972,N_7984,N_7971);
and U8973 (N_8973,N_7014,N_7156);
nor U8974 (N_8974,N_7782,N_7684);
and U8975 (N_8975,N_7984,N_7827);
or U8976 (N_8976,N_7181,N_7556);
nand U8977 (N_8977,N_7174,N_7860);
or U8978 (N_8978,N_7715,N_7683);
nand U8979 (N_8979,N_7081,N_7743);
nand U8980 (N_8980,N_7808,N_7958);
nor U8981 (N_8981,N_7483,N_7124);
and U8982 (N_8982,N_7376,N_7847);
nand U8983 (N_8983,N_7033,N_7894);
nor U8984 (N_8984,N_7056,N_7320);
nand U8985 (N_8985,N_7252,N_7687);
or U8986 (N_8986,N_7690,N_7780);
or U8987 (N_8987,N_7130,N_7162);
nand U8988 (N_8988,N_7294,N_7882);
or U8989 (N_8989,N_7091,N_7360);
and U8990 (N_8990,N_7811,N_7047);
or U8991 (N_8991,N_7300,N_7440);
or U8992 (N_8992,N_7216,N_7094);
nand U8993 (N_8993,N_7731,N_7071);
nor U8994 (N_8994,N_7715,N_7124);
or U8995 (N_8995,N_7413,N_7885);
and U8996 (N_8996,N_7357,N_7513);
nand U8997 (N_8997,N_7699,N_7618);
nor U8998 (N_8998,N_7705,N_7122);
xnor U8999 (N_8999,N_7188,N_7393);
nand U9000 (N_9000,N_8038,N_8698);
and U9001 (N_9001,N_8601,N_8501);
nand U9002 (N_9002,N_8006,N_8670);
and U9003 (N_9003,N_8811,N_8378);
or U9004 (N_9004,N_8380,N_8312);
nand U9005 (N_9005,N_8548,N_8233);
nor U9006 (N_9006,N_8503,N_8214);
nand U9007 (N_9007,N_8858,N_8276);
nand U9008 (N_9008,N_8124,N_8030);
nand U9009 (N_9009,N_8460,N_8407);
and U9010 (N_9010,N_8779,N_8660);
and U9011 (N_9011,N_8777,N_8907);
nand U9012 (N_9012,N_8212,N_8827);
and U9013 (N_9013,N_8415,N_8425);
and U9014 (N_9014,N_8438,N_8235);
nor U9015 (N_9015,N_8324,N_8513);
xnor U9016 (N_9016,N_8010,N_8547);
nor U9017 (N_9017,N_8910,N_8571);
nand U9018 (N_9018,N_8563,N_8171);
or U9019 (N_9019,N_8556,N_8027);
nor U9020 (N_9020,N_8263,N_8577);
nand U9021 (N_9021,N_8645,N_8163);
or U9022 (N_9022,N_8238,N_8929);
and U9023 (N_9023,N_8874,N_8139);
nor U9024 (N_9024,N_8491,N_8453);
nor U9025 (N_9025,N_8274,N_8300);
and U9026 (N_9026,N_8031,N_8061);
nor U9027 (N_9027,N_8986,N_8681);
and U9028 (N_9028,N_8140,N_8213);
nor U9029 (N_9029,N_8266,N_8516);
and U9030 (N_9030,N_8689,N_8111);
nor U9031 (N_9031,N_8841,N_8450);
or U9032 (N_9032,N_8461,N_8419);
and U9033 (N_9033,N_8867,N_8344);
or U9034 (N_9034,N_8083,N_8889);
nand U9035 (N_9035,N_8114,N_8988);
or U9036 (N_9036,N_8695,N_8877);
or U9037 (N_9037,N_8246,N_8924);
or U9038 (N_9038,N_8925,N_8764);
nand U9039 (N_9039,N_8589,N_8794);
and U9040 (N_9040,N_8922,N_8394);
and U9041 (N_9041,N_8041,N_8222);
nor U9042 (N_9042,N_8781,N_8927);
or U9043 (N_9043,N_8624,N_8719);
nand U9044 (N_9044,N_8742,N_8999);
nand U9045 (N_9045,N_8744,N_8609);
and U9046 (N_9046,N_8280,N_8220);
nand U9047 (N_9047,N_8353,N_8991);
or U9048 (N_9048,N_8409,N_8562);
and U9049 (N_9049,N_8046,N_8495);
and U9050 (N_9050,N_8330,N_8357);
xnor U9051 (N_9051,N_8549,N_8025);
nand U9052 (N_9052,N_8241,N_8070);
nand U9053 (N_9053,N_8985,N_8473);
nand U9054 (N_9054,N_8928,N_8679);
nand U9055 (N_9055,N_8334,N_8199);
nor U9056 (N_9056,N_8420,N_8890);
nand U9057 (N_9057,N_8658,N_8383);
nand U9058 (N_9058,N_8250,N_8422);
nand U9059 (N_9059,N_8789,N_8955);
nor U9060 (N_9060,N_8743,N_8641);
nor U9061 (N_9061,N_8126,N_8160);
nand U9062 (N_9062,N_8313,N_8686);
and U9063 (N_9063,N_8035,N_8131);
nand U9064 (N_9064,N_8170,N_8154);
or U9065 (N_9065,N_8375,N_8847);
or U9066 (N_9066,N_8539,N_8612);
or U9067 (N_9067,N_8807,N_8203);
nor U9068 (N_9068,N_8016,N_8650);
nor U9069 (N_9069,N_8172,N_8391);
and U9070 (N_9070,N_8125,N_8531);
and U9071 (N_9071,N_8224,N_8443);
nand U9072 (N_9072,N_8965,N_8879);
and U9073 (N_9073,N_8333,N_8084);
or U9074 (N_9074,N_8173,N_8261);
nor U9075 (N_9075,N_8078,N_8859);
nor U9076 (N_9076,N_8273,N_8778);
nor U9077 (N_9077,N_8147,N_8341);
nand U9078 (N_9078,N_8487,N_8356);
nand U9079 (N_9079,N_8236,N_8270);
and U9080 (N_9080,N_8785,N_8672);
and U9081 (N_9081,N_8321,N_8098);
nor U9082 (N_9082,N_8286,N_8683);
nor U9083 (N_9083,N_8845,N_8463);
nor U9084 (N_9084,N_8348,N_8995);
nand U9085 (N_9085,N_8944,N_8979);
and U9086 (N_9086,N_8718,N_8795);
and U9087 (N_9087,N_8020,N_8036);
and U9088 (N_9088,N_8726,N_8336);
nor U9089 (N_9089,N_8846,N_8521);
nand U9090 (N_9090,N_8754,N_8287);
nand U9091 (N_9091,N_8446,N_8984);
and U9092 (N_9092,N_8860,N_8676);
nor U9093 (N_9093,N_8242,N_8533);
or U9094 (N_9094,N_8893,N_8509);
nand U9095 (N_9095,N_8145,N_8382);
nor U9096 (N_9096,N_8350,N_8730);
xnor U9097 (N_9097,N_8223,N_8723);
or U9098 (N_9098,N_8833,N_8081);
nor U9099 (N_9099,N_8554,N_8525);
nor U9100 (N_9100,N_8505,N_8322);
and U9101 (N_9101,N_8133,N_8099);
nand U9102 (N_9102,N_8392,N_8408);
or U9103 (N_9103,N_8054,N_8064);
nand U9104 (N_9104,N_8970,N_8788);
and U9105 (N_9105,N_8216,N_8143);
and U9106 (N_9106,N_8062,N_8331);
and U9107 (N_9107,N_8857,N_8468);
nand U9108 (N_9108,N_8417,N_8558);
nand U9109 (N_9109,N_8427,N_8507);
or U9110 (N_9110,N_8756,N_8192);
nand U9111 (N_9111,N_8663,N_8106);
nor U9112 (N_9112,N_8901,N_8015);
nand U9113 (N_9113,N_8080,N_8464);
nand U9114 (N_9114,N_8178,N_8195);
and U9115 (N_9115,N_8949,N_8042);
or U9116 (N_9116,N_8423,N_8814);
nand U9117 (N_9117,N_8724,N_8349);
or U9118 (N_9118,N_8024,N_8174);
or U9119 (N_9119,N_8390,N_8141);
and U9120 (N_9120,N_8694,N_8467);
and U9121 (N_9121,N_8760,N_8844);
and U9122 (N_9122,N_8977,N_8715);
nor U9123 (N_9123,N_8520,N_8699);
nand U9124 (N_9124,N_8614,N_8234);
nand U9125 (N_9125,N_8152,N_8532);
nor U9126 (N_9126,N_8588,N_8630);
nand U9127 (N_9127,N_8295,N_8921);
or U9128 (N_9128,N_8604,N_8388);
nand U9129 (N_9129,N_8570,N_8720);
and U9130 (N_9130,N_8668,N_8197);
or U9131 (N_9131,N_8477,N_8882);
nand U9132 (N_9132,N_8637,N_8886);
or U9133 (N_9133,N_8307,N_8484);
nor U9134 (N_9134,N_8960,N_8166);
nor U9135 (N_9135,N_8191,N_8018);
nand U9136 (N_9136,N_8937,N_8204);
or U9137 (N_9137,N_8871,N_8414);
or U9138 (N_9138,N_8586,N_8411);
nor U9139 (N_9139,N_8073,N_8297);
nor U9140 (N_9140,N_8705,N_8623);
nor U9141 (N_9141,N_8413,N_8369);
or U9142 (N_9142,N_8763,N_8475);
and U9143 (N_9143,N_8014,N_8958);
nor U9144 (N_9144,N_8625,N_8696);
nand U9145 (N_9145,N_8673,N_8605);
and U9146 (N_9146,N_8135,N_8856);
nor U9147 (N_9147,N_8915,N_8485);
nor U9148 (N_9148,N_8825,N_8264);
or U9149 (N_9149,N_8346,N_8308);
nor U9150 (N_9150,N_8112,N_8189);
and U9151 (N_9151,N_8034,N_8864);
or U9152 (N_9152,N_8952,N_8664);
or U9153 (N_9153,N_8768,N_8741);
and U9154 (N_9154,N_8838,N_8755);
or U9155 (N_9155,N_8550,N_8682);
nor U9156 (N_9156,N_8832,N_8530);
or U9157 (N_9157,N_8736,N_8130);
and U9158 (N_9158,N_8721,N_8524);
nor U9159 (N_9159,N_8607,N_8181);
and U9160 (N_9160,N_8410,N_8608);
nor U9161 (N_9161,N_8469,N_8745);
nand U9162 (N_9162,N_8567,N_8622);
nand U9163 (N_9163,N_8265,N_8587);
or U9164 (N_9164,N_8938,N_8662);
nand U9165 (N_9165,N_8474,N_8431);
or U9166 (N_9166,N_8087,N_8455);
and U9167 (N_9167,N_8366,N_8218);
nor U9168 (N_9168,N_8058,N_8956);
and U9169 (N_9169,N_8717,N_8905);
or U9170 (N_9170,N_8129,N_8167);
and U9171 (N_9171,N_8826,N_8542);
nand U9172 (N_9172,N_8319,N_8998);
nor U9173 (N_9173,N_8289,N_8972);
or U9174 (N_9174,N_8177,N_8506);
and U9175 (N_9175,N_8045,N_8941);
and U9176 (N_9176,N_8361,N_8365);
nand U9177 (N_9177,N_8499,N_8797);
or U9178 (N_9178,N_8186,N_8003);
nor U9179 (N_9179,N_8428,N_8594);
nor U9180 (N_9180,N_8296,N_8386);
xnor U9181 (N_9181,N_8316,N_8596);
and U9182 (N_9182,N_8101,N_8619);
nand U9183 (N_9183,N_8399,N_8783);
and U9184 (N_9184,N_8787,N_8028);
nand U9185 (N_9185,N_8254,N_8648);
and U9186 (N_9186,N_8272,N_8740);
and U9187 (N_9187,N_8066,N_8279);
nor U9188 (N_9188,N_8175,N_8592);
or U9189 (N_9189,N_8339,N_8470);
nor U9190 (N_9190,N_8931,N_8896);
and U9191 (N_9191,N_8733,N_8458);
or U9192 (N_9192,N_8561,N_8688);
nor U9193 (N_9193,N_8643,N_8968);
and U9194 (N_9194,N_8818,N_8828);
or U9195 (N_9195,N_8945,N_8578);
nor U9196 (N_9196,N_8712,N_8440);
and U9197 (N_9197,N_8540,N_8466);
nor U9198 (N_9198,N_8076,N_8703);
nand U9199 (N_9199,N_8009,N_8198);
and U9200 (N_9200,N_8278,N_8819);
or U9201 (N_9201,N_8259,N_8606);
and U9202 (N_9202,N_8320,N_8872);
or U9203 (N_9203,N_8044,N_8429);
nor U9204 (N_9204,N_8104,N_8151);
nand U9205 (N_9205,N_8528,N_8784);
nor U9206 (N_9206,N_8217,N_8775);
or U9207 (N_9207,N_8687,N_8884);
nand U9208 (N_9208,N_8978,N_8284);
or U9209 (N_9209,N_8400,N_8600);
nor U9210 (N_9210,N_8888,N_8653);
and U9211 (N_9211,N_8674,N_8919);
nand U9212 (N_9212,N_8823,N_8808);
and U9213 (N_9213,N_8100,N_8142);
and U9214 (N_9214,N_8959,N_8916);
or U9215 (N_9215,N_8817,N_8961);
nor U9216 (N_9216,N_8615,N_8761);
xnor U9217 (N_9217,N_8875,N_8725);
nand U9218 (N_9218,N_8515,N_8148);
nand U9219 (N_9219,N_8634,N_8940);
nand U9220 (N_9220,N_8822,N_8591);
or U9221 (N_9221,N_8019,N_8881);
or U9222 (N_9222,N_8997,N_8168);
nor U9223 (N_9223,N_8180,N_8776);
and U9224 (N_9224,N_8982,N_8337);
nor U9225 (N_9225,N_8667,N_8512);
nand U9226 (N_9226,N_8576,N_8702);
nand U9227 (N_9227,N_8281,N_8082);
or U9228 (N_9228,N_8950,N_8059);
nand U9229 (N_9229,N_8404,N_8226);
or U9230 (N_9230,N_8208,N_8060);
and U9231 (N_9231,N_8363,N_8465);
nand U9232 (N_9232,N_8457,N_8255);
nor U9233 (N_9233,N_8671,N_8117);
nand U9234 (N_9234,N_8086,N_8815);
and U9235 (N_9235,N_8435,N_8831);
nand U9236 (N_9236,N_8697,N_8240);
or U9237 (N_9237,N_8138,N_8498);
and U9238 (N_9238,N_8462,N_8853);
or U9239 (N_9239,N_8360,N_8275);
nand U9240 (N_9240,N_8948,N_8656);
or U9241 (N_9241,N_8782,N_8071);
or U9242 (N_9242,N_8870,N_8115);
and U9243 (N_9243,N_8969,N_8711);
nor U9244 (N_9244,N_8047,N_8362);
nor U9245 (N_9245,N_8966,N_8902);
nor U9246 (N_9246,N_8579,N_8793);
and U9247 (N_9247,N_8747,N_8483);
or U9248 (N_9248,N_8627,N_8529);
or U9249 (N_9249,N_8885,N_8231);
and U9250 (N_9250,N_8370,N_8454);
and U9251 (N_9251,N_8574,N_8210);
nand U9252 (N_9252,N_8200,N_8056);
nand U9253 (N_9253,N_8573,N_8633);
nor U9254 (N_9254,N_8611,N_8708);
or U9255 (N_9255,N_8824,N_8017);
nor U9256 (N_9256,N_8481,N_8786);
nand U9257 (N_9257,N_8479,N_8748);
or U9258 (N_9258,N_8480,N_8839);
nand U9259 (N_9259,N_8790,N_8401);
nor U9260 (N_9260,N_8471,N_8368);
and U9261 (N_9261,N_8892,N_8813);
nand U9262 (N_9262,N_8759,N_8862);
or U9263 (N_9263,N_8150,N_8700);
nor U9264 (N_9264,N_8749,N_8716);
nor U9265 (N_9265,N_8773,N_8335);
or U9266 (N_9266,N_8476,N_8644);
and U9267 (N_9267,N_8447,N_8780);
and U9268 (N_9268,N_8001,N_8290);
and U9269 (N_9269,N_8434,N_8387);
nand U9270 (N_9270,N_8555,N_8232);
or U9271 (N_9271,N_8936,N_8315);
and U9272 (N_9272,N_8632,N_8108);
or U9273 (N_9273,N_8738,N_8920);
and U9274 (N_9274,N_8109,N_8523);
nand U9275 (N_9275,N_8635,N_8305);
or U9276 (N_9276,N_8367,N_8957);
and U9277 (N_9277,N_8048,N_8156);
nor U9278 (N_9278,N_8918,N_8973);
nor U9279 (N_9279,N_8758,N_8753);
nand U9280 (N_9280,N_8183,N_8165);
nor U9281 (N_9281,N_8205,N_8136);
nand U9282 (N_9282,N_8294,N_8618);
nor U9283 (N_9283,N_8534,N_8565);
nand U9284 (N_9284,N_8908,N_8057);
nor U9285 (N_9285,N_8580,N_8221);
nor U9286 (N_9286,N_8526,N_8193);
nand U9287 (N_9287,N_8436,N_8626);
and U9288 (N_9288,N_8628,N_8169);
nand U9289 (N_9289,N_8842,N_8906);
nand U9290 (N_9290,N_8654,N_8092);
xor U9291 (N_9291,N_8327,N_8582);
nor U9292 (N_9292,N_8829,N_8868);
and U9293 (N_9293,N_8739,N_8439);
or U9294 (N_9294,N_8544,N_8089);
and U9295 (N_9295,N_8291,N_8381);
and U9296 (N_9296,N_8980,N_8848);
and U9297 (N_9297,N_8283,N_8012);
and U9298 (N_9298,N_8005,N_8405);
and U9299 (N_9299,N_8621,N_8248);
nand U9300 (N_9300,N_8207,N_8299);
nand U9301 (N_9301,N_8752,N_8954);
nor U9302 (N_9302,N_8993,N_8351);
nor U9303 (N_9303,N_8735,N_8772);
nand U9304 (N_9304,N_8202,N_8655);
and U9305 (N_9305,N_8063,N_8861);
nor U9306 (N_9306,N_8159,N_8900);
or U9307 (N_9307,N_8091,N_8511);
nor U9308 (N_9308,N_8430,N_8182);
nand U9309 (N_9309,N_8727,N_8282);
nor U9310 (N_9310,N_8432,N_8103);
nor U9311 (N_9311,N_8732,N_8052);
nand U9312 (N_9312,N_8271,N_8134);
or U9313 (N_9313,N_8347,N_8489);
or U9314 (N_9314,N_8209,N_8116);
nand U9315 (N_9315,N_8545,N_8564);
nor U9316 (N_9316,N_8765,N_8096);
or U9317 (N_9317,N_8358,N_8424);
nor U9318 (N_9318,N_8445,N_8118);
nand U9319 (N_9319,N_8854,N_8559);
xor U9320 (N_9320,N_8459,N_8904);
nor U9321 (N_9321,N_8963,N_8298);
nand U9322 (N_9322,N_8691,N_8593);
and U9323 (N_9323,N_8933,N_8267);
nor U9324 (N_9324,N_8917,N_8396);
nor U9325 (N_9325,N_8049,N_8494);
nor U9326 (N_9326,N_8799,N_8373);
nand U9327 (N_9327,N_8575,N_8206);
or U9328 (N_9328,N_8569,N_8566);
or U9329 (N_9329,N_8137,N_8535);
nor U9330 (N_9330,N_8376,N_8403);
nor U9331 (N_9331,N_8983,N_8887);
nand U9332 (N_9332,N_8119,N_8769);
and U9333 (N_9333,N_8004,N_8364);
nand U9334 (N_9334,N_8301,N_8728);
nand U9335 (N_9335,N_8433,N_8478);
nand U9336 (N_9336,N_8899,N_8328);
and U9337 (N_9337,N_8514,N_8994);
and U9338 (N_9338,N_8398,N_8646);
and U9339 (N_9339,N_8157,N_8597);
nor U9340 (N_9340,N_8876,N_8690);
nand U9341 (N_9341,N_8449,N_8040);
and U9342 (N_9342,N_8293,N_8803);
or U9343 (N_9343,N_8196,N_8603);
nor U9344 (N_9344,N_8680,N_8493);
and U9345 (N_9345,N_8029,N_8215);
and U9346 (N_9346,N_8402,N_8093);
nand U9347 (N_9347,N_8714,N_8964);
nor U9348 (N_9348,N_8770,N_8201);
nor U9349 (N_9349,N_8065,N_8069);
nor U9350 (N_9350,N_8572,N_8537);
and U9351 (N_9351,N_8821,N_8345);
nor U9352 (N_9352,N_8568,N_8602);
or U9353 (N_9353,N_8000,N_8317);
or U9354 (N_9354,N_8657,N_8472);
nand U9355 (N_9355,N_8406,N_8228);
nor U9356 (N_9356,N_8187,N_8026);
nor U9357 (N_9357,N_8522,N_8962);
or U9358 (N_9358,N_8384,N_8309);
nand U9359 (N_9359,N_8891,N_8923);
and U9360 (N_9360,N_8132,N_8704);
nand U9361 (N_9361,N_8379,N_8149);
or U9362 (N_9362,N_8258,N_8395);
nand U9363 (N_9363,N_8551,N_8385);
or U9364 (N_9364,N_8895,N_8932);
or U9365 (N_9365,N_8510,N_8975);
or U9366 (N_9366,N_8865,N_8880);
or U9367 (N_9367,N_8437,N_8153);
or U9368 (N_9368,N_8620,N_8541);
and U9369 (N_9369,N_8584,N_8072);
and U9370 (N_9370,N_8176,N_8912);
xor U9371 (N_9371,N_8179,N_8863);
xnor U9372 (N_9372,N_8022,N_8120);
nand U9373 (N_9373,N_8053,N_8194);
nor U9374 (N_9374,N_8237,N_8710);
nor U9375 (N_9375,N_8771,N_8037);
nand U9376 (N_9376,N_8251,N_8393);
nand U9377 (N_9377,N_8849,N_8837);
xor U9378 (N_9378,N_8617,N_8444);
nand U9379 (N_9379,N_8926,N_8946);
nor U9380 (N_9380,N_8951,N_8903);
nor U9381 (N_9381,N_8722,N_8989);
nor U9382 (N_9382,N_8277,N_8935);
or U9383 (N_9383,N_8750,N_8894);
and U9384 (N_9384,N_8225,N_8599);
nor U9385 (N_9385,N_8050,N_8067);
and U9386 (N_9386,N_8372,N_8023);
nor U9387 (N_9387,N_8798,N_8074);
nor U9388 (N_9388,N_8253,N_8441);
nor U9389 (N_9389,N_8371,N_8007);
and U9390 (N_9390,N_8943,N_8734);
nand U9391 (N_9391,N_8883,N_8377);
nand U9392 (N_9392,N_8075,N_8757);
nand U9393 (N_9393,N_8032,N_8247);
nand U9394 (N_9394,N_8342,N_8737);
or U9395 (N_9395,N_8397,N_8389);
and U9396 (N_9396,N_8102,N_8546);
or U9397 (N_9397,N_8557,N_8105);
or U9398 (N_9398,N_8302,N_8836);
or U9399 (N_9399,N_8068,N_8585);
or U9400 (N_9400,N_8911,N_8185);
and U9401 (N_9401,N_8939,N_8971);
or U9402 (N_9402,N_8002,N_8640);
nand U9403 (N_9403,N_8451,N_8517);
and U9404 (N_9404,N_8245,N_8416);
nor U9405 (N_9405,N_8636,N_8482);
or U9406 (N_9406,N_8590,N_8610);
nor U9407 (N_9407,N_8113,N_8990);
nand U9408 (N_9408,N_8260,N_8638);
or U9409 (N_9409,N_8269,N_8581);
and U9410 (N_9410,N_8190,N_8709);
or U9411 (N_9411,N_8033,N_8981);
nand U9412 (N_9412,N_8805,N_8292);
nor U9413 (N_9413,N_8996,N_8613);
or U9414 (N_9414,N_8162,N_8751);
nor U9415 (N_9415,N_8107,N_8852);
or U9416 (N_9416,N_8230,N_8536);
or U9417 (N_9417,N_8332,N_8707);
nand U9418 (N_9418,N_8873,N_8791);
nand U9419 (N_9419,N_8519,N_8122);
nor U9420 (N_9420,N_8155,N_8898);
nand U9421 (N_9421,N_8502,N_8097);
nand U9422 (N_9422,N_8810,N_8184);
and U9423 (N_9423,N_8835,N_8303);
xor U9424 (N_9424,N_8079,N_8318);
nand U9425 (N_9425,N_8110,N_8974);
nor U9426 (N_9426,N_8947,N_8088);
and U9427 (N_9427,N_8008,N_8121);
nor U9428 (N_9428,N_8128,N_8869);
nand U9429 (N_9429,N_8639,N_8085);
or U9430 (N_9430,N_8352,N_8488);
nor U9431 (N_9431,N_8412,N_8508);
nand U9432 (N_9432,N_8011,N_8843);
xor U9433 (N_9433,N_8518,N_8953);
nand U9434 (N_9434,N_8486,N_8942);
xnor U9435 (N_9435,N_8675,N_8649);
or U9436 (N_9436,N_8796,N_8161);
nor U9437 (N_9437,N_8355,N_8314);
nand U9438 (N_9438,N_8693,N_8834);
nand U9439 (N_9439,N_8325,N_8665);
or U9440 (N_9440,N_8806,N_8329);
nand U9441 (N_9441,N_8661,N_8914);
or U9442 (N_9442,N_8598,N_8731);
nor U9443 (N_9443,N_8774,N_8692);
and U9444 (N_9444,N_8629,N_8909);
and U9445 (N_9445,N_8252,N_8285);
nand U9446 (N_9446,N_8496,N_8310);
or U9447 (N_9447,N_8897,N_8164);
nor U9448 (N_9448,N_8338,N_8262);
nor U9449 (N_9449,N_8851,N_8144);
or U9450 (N_9450,N_8616,N_8840);
nand U9451 (N_9451,N_8802,N_8792);
nor U9452 (N_9452,N_8452,N_8538);
and U9453 (N_9453,N_8677,N_8326);
and U9454 (N_9454,N_8659,N_8583);
and U9455 (N_9455,N_8244,N_8543);
or U9456 (N_9456,N_8306,N_8878);
and U9457 (N_9457,N_8227,N_8448);
and U9458 (N_9458,N_8504,N_8219);
or U9459 (N_9459,N_8767,N_8374);
and U9460 (N_9460,N_8766,N_8340);
nand U9461 (N_9461,N_8684,N_8268);
or U9462 (N_9462,N_8497,N_8490);
nand U9463 (N_9463,N_8229,N_8553);
nand U9464 (N_9464,N_8354,N_8746);
nor U9465 (N_9465,N_8527,N_8256);
nand U9466 (N_9466,N_8850,N_8456);
and U9467 (N_9467,N_8642,N_8442);
nor U9468 (N_9468,N_8678,N_8651);
nand U9469 (N_9469,N_8685,N_8560);
and U9470 (N_9470,N_8158,N_8595);
and U9471 (N_9471,N_8976,N_8934);
nor U9472 (N_9472,N_8418,N_8090);
nand U9473 (N_9473,N_8647,N_8426);
nand U9474 (N_9474,N_8013,N_8866);
and U9475 (N_9475,N_8987,N_8830);
nand U9476 (N_9476,N_8077,N_8631);
nor U9477 (N_9477,N_8762,N_8288);
and U9478 (N_9478,N_8188,N_8500);
or U9479 (N_9479,N_8239,N_8855);
nand U9480 (N_9480,N_8304,N_8094);
and U9481 (N_9481,N_8801,N_8343);
or U9482 (N_9482,N_8812,N_8055);
or U9483 (N_9483,N_8243,N_8051);
nor U9484 (N_9484,N_8804,N_8913);
or U9485 (N_9485,N_8127,N_8311);
nor U9486 (N_9486,N_8492,N_8706);
or U9487 (N_9487,N_8123,N_8421);
nor U9488 (N_9488,N_8021,N_8701);
or U9489 (N_9489,N_8729,N_8211);
and U9490 (N_9490,N_8359,N_8669);
and U9491 (N_9491,N_8992,N_8820);
or U9492 (N_9492,N_8652,N_8323);
or U9493 (N_9493,N_8043,N_8713);
or U9494 (N_9494,N_8552,N_8039);
and U9495 (N_9495,N_8257,N_8666);
nor U9496 (N_9496,N_8249,N_8809);
or U9497 (N_9497,N_8095,N_8816);
and U9498 (N_9498,N_8930,N_8146);
nor U9499 (N_9499,N_8967,N_8800);
and U9500 (N_9500,N_8303,N_8527);
nor U9501 (N_9501,N_8790,N_8866);
xor U9502 (N_9502,N_8721,N_8681);
nand U9503 (N_9503,N_8922,N_8590);
and U9504 (N_9504,N_8732,N_8721);
and U9505 (N_9505,N_8440,N_8044);
nor U9506 (N_9506,N_8121,N_8896);
and U9507 (N_9507,N_8374,N_8725);
nand U9508 (N_9508,N_8684,N_8677);
nand U9509 (N_9509,N_8586,N_8023);
nand U9510 (N_9510,N_8387,N_8156);
and U9511 (N_9511,N_8907,N_8325);
and U9512 (N_9512,N_8356,N_8500);
nor U9513 (N_9513,N_8930,N_8009);
nor U9514 (N_9514,N_8888,N_8615);
nand U9515 (N_9515,N_8270,N_8520);
nor U9516 (N_9516,N_8753,N_8477);
nand U9517 (N_9517,N_8305,N_8838);
nand U9518 (N_9518,N_8228,N_8886);
and U9519 (N_9519,N_8373,N_8336);
nor U9520 (N_9520,N_8756,N_8541);
and U9521 (N_9521,N_8937,N_8248);
or U9522 (N_9522,N_8069,N_8482);
or U9523 (N_9523,N_8165,N_8779);
or U9524 (N_9524,N_8965,N_8057);
or U9525 (N_9525,N_8658,N_8282);
xor U9526 (N_9526,N_8818,N_8117);
xor U9527 (N_9527,N_8670,N_8652);
nor U9528 (N_9528,N_8323,N_8411);
nand U9529 (N_9529,N_8277,N_8880);
nand U9530 (N_9530,N_8997,N_8020);
or U9531 (N_9531,N_8182,N_8342);
or U9532 (N_9532,N_8312,N_8908);
nand U9533 (N_9533,N_8273,N_8220);
nor U9534 (N_9534,N_8904,N_8900);
nor U9535 (N_9535,N_8592,N_8844);
and U9536 (N_9536,N_8077,N_8987);
nor U9537 (N_9537,N_8678,N_8761);
nor U9538 (N_9538,N_8252,N_8590);
nand U9539 (N_9539,N_8977,N_8778);
nand U9540 (N_9540,N_8823,N_8508);
or U9541 (N_9541,N_8654,N_8727);
nor U9542 (N_9542,N_8184,N_8026);
and U9543 (N_9543,N_8506,N_8266);
and U9544 (N_9544,N_8791,N_8652);
nor U9545 (N_9545,N_8994,N_8613);
and U9546 (N_9546,N_8701,N_8227);
and U9547 (N_9547,N_8405,N_8532);
nand U9548 (N_9548,N_8430,N_8714);
and U9549 (N_9549,N_8116,N_8479);
nor U9550 (N_9550,N_8765,N_8342);
and U9551 (N_9551,N_8109,N_8876);
or U9552 (N_9552,N_8450,N_8105);
nand U9553 (N_9553,N_8154,N_8985);
or U9554 (N_9554,N_8902,N_8607);
nor U9555 (N_9555,N_8647,N_8592);
or U9556 (N_9556,N_8959,N_8827);
nand U9557 (N_9557,N_8270,N_8746);
or U9558 (N_9558,N_8396,N_8263);
nor U9559 (N_9559,N_8389,N_8244);
xor U9560 (N_9560,N_8679,N_8105);
or U9561 (N_9561,N_8920,N_8384);
or U9562 (N_9562,N_8813,N_8021);
or U9563 (N_9563,N_8314,N_8748);
nand U9564 (N_9564,N_8897,N_8936);
or U9565 (N_9565,N_8574,N_8546);
nor U9566 (N_9566,N_8582,N_8608);
or U9567 (N_9567,N_8235,N_8159);
nor U9568 (N_9568,N_8269,N_8458);
or U9569 (N_9569,N_8300,N_8252);
nor U9570 (N_9570,N_8221,N_8626);
xor U9571 (N_9571,N_8333,N_8655);
nand U9572 (N_9572,N_8523,N_8326);
and U9573 (N_9573,N_8122,N_8937);
and U9574 (N_9574,N_8965,N_8391);
nand U9575 (N_9575,N_8019,N_8409);
or U9576 (N_9576,N_8039,N_8860);
nand U9577 (N_9577,N_8485,N_8092);
nor U9578 (N_9578,N_8582,N_8687);
or U9579 (N_9579,N_8653,N_8542);
xnor U9580 (N_9580,N_8005,N_8598);
and U9581 (N_9581,N_8896,N_8052);
nor U9582 (N_9582,N_8418,N_8869);
nor U9583 (N_9583,N_8015,N_8079);
nor U9584 (N_9584,N_8960,N_8314);
or U9585 (N_9585,N_8277,N_8182);
and U9586 (N_9586,N_8300,N_8122);
nor U9587 (N_9587,N_8554,N_8450);
nor U9588 (N_9588,N_8269,N_8695);
and U9589 (N_9589,N_8590,N_8567);
and U9590 (N_9590,N_8947,N_8170);
or U9591 (N_9591,N_8047,N_8512);
and U9592 (N_9592,N_8122,N_8838);
nand U9593 (N_9593,N_8734,N_8759);
or U9594 (N_9594,N_8984,N_8987);
or U9595 (N_9595,N_8260,N_8307);
nand U9596 (N_9596,N_8496,N_8788);
nand U9597 (N_9597,N_8788,N_8538);
nand U9598 (N_9598,N_8269,N_8981);
nand U9599 (N_9599,N_8923,N_8174);
or U9600 (N_9600,N_8518,N_8590);
or U9601 (N_9601,N_8956,N_8076);
and U9602 (N_9602,N_8738,N_8122);
and U9603 (N_9603,N_8382,N_8211);
and U9604 (N_9604,N_8565,N_8908);
nor U9605 (N_9605,N_8963,N_8003);
xnor U9606 (N_9606,N_8034,N_8081);
and U9607 (N_9607,N_8933,N_8217);
or U9608 (N_9608,N_8790,N_8908);
nand U9609 (N_9609,N_8171,N_8319);
xnor U9610 (N_9610,N_8473,N_8417);
nor U9611 (N_9611,N_8039,N_8436);
xor U9612 (N_9612,N_8990,N_8251);
and U9613 (N_9613,N_8046,N_8007);
nor U9614 (N_9614,N_8406,N_8524);
or U9615 (N_9615,N_8125,N_8955);
and U9616 (N_9616,N_8956,N_8572);
xnor U9617 (N_9617,N_8762,N_8790);
or U9618 (N_9618,N_8344,N_8168);
or U9619 (N_9619,N_8526,N_8651);
nor U9620 (N_9620,N_8102,N_8152);
nor U9621 (N_9621,N_8829,N_8889);
nor U9622 (N_9622,N_8890,N_8521);
nor U9623 (N_9623,N_8849,N_8057);
nor U9624 (N_9624,N_8014,N_8306);
or U9625 (N_9625,N_8657,N_8290);
nand U9626 (N_9626,N_8388,N_8995);
and U9627 (N_9627,N_8186,N_8760);
nand U9628 (N_9628,N_8788,N_8424);
nand U9629 (N_9629,N_8122,N_8257);
nor U9630 (N_9630,N_8866,N_8217);
nor U9631 (N_9631,N_8246,N_8627);
and U9632 (N_9632,N_8028,N_8218);
or U9633 (N_9633,N_8651,N_8983);
nand U9634 (N_9634,N_8850,N_8467);
nor U9635 (N_9635,N_8770,N_8193);
nand U9636 (N_9636,N_8908,N_8905);
or U9637 (N_9637,N_8912,N_8201);
or U9638 (N_9638,N_8574,N_8628);
nor U9639 (N_9639,N_8733,N_8644);
nor U9640 (N_9640,N_8125,N_8868);
and U9641 (N_9641,N_8763,N_8061);
nor U9642 (N_9642,N_8211,N_8968);
or U9643 (N_9643,N_8810,N_8613);
and U9644 (N_9644,N_8920,N_8504);
nor U9645 (N_9645,N_8425,N_8911);
nor U9646 (N_9646,N_8333,N_8437);
and U9647 (N_9647,N_8721,N_8332);
nor U9648 (N_9648,N_8273,N_8102);
or U9649 (N_9649,N_8415,N_8991);
nor U9650 (N_9650,N_8031,N_8943);
and U9651 (N_9651,N_8405,N_8732);
and U9652 (N_9652,N_8321,N_8917);
nor U9653 (N_9653,N_8972,N_8773);
or U9654 (N_9654,N_8181,N_8582);
and U9655 (N_9655,N_8392,N_8401);
or U9656 (N_9656,N_8384,N_8083);
and U9657 (N_9657,N_8643,N_8832);
nor U9658 (N_9658,N_8000,N_8491);
nand U9659 (N_9659,N_8878,N_8105);
nor U9660 (N_9660,N_8337,N_8984);
and U9661 (N_9661,N_8483,N_8712);
or U9662 (N_9662,N_8033,N_8533);
nor U9663 (N_9663,N_8246,N_8130);
nor U9664 (N_9664,N_8285,N_8775);
xor U9665 (N_9665,N_8484,N_8971);
nor U9666 (N_9666,N_8509,N_8471);
or U9667 (N_9667,N_8458,N_8832);
nand U9668 (N_9668,N_8989,N_8999);
or U9669 (N_9669,N_8108,N_8702);
nand U9670 (N_9670,N_8422,N_8403);
and U9671 (N_9671,N_8067,N_8396);
nand U9672 (N_9672,N_8911,N_8099);
or U9673 (N_9673,N_8957,N_8169);
nor U9674 (N_9674,N_8663,N_8224);
and U9675 (N_9675,N_8758,N_8939);
and U9676 (N_9676,N_8814,N_8756);
nand U9677 (N_9677,N_8362,N_8032);
nand U9678 (N_9678,N_8412,N_8454);
nand U9679 (N_9679,N_8365,N_8933);
nor U9680 (N_9680,N_8048,N_8436);
nor U9681 (N_9681,N_8648,N_8762);
nand U9682 (N_9682,N_8047,N_8321);
nand U9683 (N_9683,N_8329,N_8829);
or U9684 (N_9684,N_8964,N_8933);
or U9685 (N_9685,N_8312,N_8587);
nand U9686 (N_9686,N_8576,N_8986);
or U9687 (N_9687,N_8500,N_8385);
or U9688 (N_9688,N_8209,N_8890);
nor U9689 (N_9689,N_8900,N_8084);
nor U9690 (N_9690,N_8352,N_8168);
nand U9691 (N_9691,N_8526,N_8990);
or U9692 (N_9692,N_8453,N_8300);
nor U9693 (N_9693,N_8999,N_8069);
or U9694 (N_9694,N_8517,N_8225);
nor U9695 (N_9695,N_8982,N_8184);
and U9696 (N_9696,N_8484,N_8788);
nor U9697 (N_9697,N_8794,N_8696);
xor U9698 (N_9698,N_8732,N_8226);
nand U9699 (N_9699,N_8847,N_8735);
nand U9700 (N_9700,N_8599,N_8110);
or U9701 (N_9701,N_8578,N_8890);
xnor U9702 (N_9702,N_8719,N_8303);
or U9703 (N_9703,N_8838,N_8334);
nand U9704 (N_9704,N_8984,N_8098);
nand U9705 (N_9705,N_8342,N_8484);
and U9706 (N_9706,N_8270,N_8030);
and U9707 (N_9707,N_8337,N_8863);
and U9708 (N_9708,N_8591,N_8043);
nor U9709 (N_9709,N_8100,N_8549);
or U9710 (N_9710,N_8948,N_8649);
and U9711 (N_9711,N_8685,N_8619);
nor U9712 (N_9712,N_8055,N_8227);
and U9713 (N_9713,N_8496,N_8016);
or U9714 (N_9714,N_8796,N_8083);
or U9715 (N_9715,N_8635,N_8787);
nor U9716 (N_9716,N_8605,N_8652);
and U9717 (N_9717,N_8955,N_8468);
and U9718 (N_9718,N_8071,N_8499);
nand U9719 (N_9719,N_8227,N_8277);
nand U9720 (N_9720,N_8605,N_8059);
nand U9721 (N_9721,N_8105,N_8665);
nand U9722 (N_9722,N_8408,N_8933);
and U9723 (N_9723,N_8893,N_8320);
or U9724 (N_9724,N_8465,N_8116);
or U9725 (N_9725,N_8305,N_8784);
nor U9726 (N_9726,N_8511,N_8554);
nand U9727 (N_9727,N_8969,N_8387);
and U9728 (N_9728,N_8490,N_8263);
xor U9729 (N_9729,N_8716,N_8426);
nor U9730 (N_9730,N_8623,N_8558);
and U9731 (N_9731,N_8851,N_8263);
nand U9732 (N_9732,N_8078,N_8103);
nor U9733 (N_9733,N_8441,N_8655);
nor U9734 (N_9734,N_8939,N_8075);
nor U9735 (N_9735,N_8913,N_8082);
xnor U9736 (N_9736,N_8695,N_8906);
xnor U9737 (N_9737,N_8267,N_8053);
or U9738 (N_9738,N_8137,N_8725);
and U9739 (N_9739,N_8443,N_8292);
and U9740 (N_9740,N_8819,N_8270);
nor U9741 (N_9741,N_8665,N_8193);
nand U9742 (N_9742,N_8466,N_8842);
or U9743 (N_9743,N_8454,N_8834);
nand U9744 (N_9744,N_8922,N_8434);
and U9745 (N_9745,N_8949,N_8206);
nand U9746 (N_9746,N_8022,N_8709);
nand U9747 (N_9747,N_8775,N_8596);
nor U9748 (N_9748,N_8049,N_8115);
and U9749 (N_9749,N_8375,N_8528);
and U9750 (N_9750,N_8097,N_8087);
nand U9751 (N_9751,N_8883,N_8066);
and U9752 (N_9752,N_8031,N_8141);
and U9753 (N_9753,N_8861,N_8709);
xnor U9754 (N_9754,N_8097,N_8944);
nor U9755 (N_9755,N_8180,N_8173);
nor U9756 (N_9756,N_8628,N_8561);
nand U9757 (N_9757,N_8458,N_8541);
nand U9758 (N_9758,N_8756,N_8789);
nand U9759 (N_9759,N_8057,N_8951);
and U9760 (N_9760,N_8813,N_8533);
or U9761 (N_9761,N_8746,N_8335);
nand U9762 (N_9762,N_8020,N_8006);
or U9763 (N_9763,N_8029,N_8363);
nand U9764 (N_9764,N_8560,N_8952);
and U9765 (N_9765,N_8449,N_8986);
or U9766 (N_9766,N_8481,N_8138);
and U9767 (N_9767,N_8918,N_8081);
nand U9768 (N_9768,N_8225,N_8248);
xor U9769 (N_9769,N_8278,N_8171);
and U9770 (N_9770,N_8741,N_8920);
and U9771 (N_9771,N_8775,N_8414);
nand U9772 (N_9772,N_8646,N_8959);
and U9773 (N_9773,N_8395,N_8256);
and U9774 (N_9774,N_8329,N_8328);
nor U9775 (N_9775,N_8705,N_8245);
nor U9776 (N_9776,N_8398,N_8200);
and U9777 (N_9777,N_8366,N_8247);
nand U9778 (N_9778,N_8842,N_8086);
nor U9779 (N_9779,N_8929,N_8954);
and U9780 (N_9780,N_8348,N_8616);
nor U9781 (N_9781,N_8867,N_8927);
and U9782 (N_9782,N_8542,N_8995);
nor U9783 (N_9783,N_8312,N_8150);
nand U9784 (N_9784,N_8318,N_8661);
or U9785 (N_9785,N_8453,N_8636);
nor U9786 (N_9786,N_8500,N_8993);
or U9787 (N_9787,N_8069,N_8429);
or U9788 (N_9788,N_8331,N_8294);
nor U9789 (N_9789,N_8215,N_8421);
and U9790 (N_9790,N_8026,N_8150);
or U9791 (N_9791,N_8590,N_8080);
nand U9792 (N_9792,N_8742,N_8243);
or U9793 (N_9793,N_8957,N_8808);
or U9794 (N_9794,N_8455,N_8205);
and U9795 (N_9795,N_8832,N_8406);
nor U9796 (N_9796,N_8611,N_8529);
nor U9797 (N_9797,N_8305,N_8874);
and U9798 (N_9798,N_8461,N_8831);
nand U9799 (N_9799,N_8925,N_8168);
nor U9800 (N_9800,N_8860,N_8017);
or U9801 (N_9801,N_8574,N_8244);
or U9802 (N_9802,N_8649,N_8137);
and U9803 (N_9803,N_8891,N_8888);
nand U9804 (N_9804,N_8530,N_8157);
nor U9805 (N_9805,N_8773,N_8256);
nand U9806 (N_9806,N_8090,N_8906);
or U9807 (N_9807,N_8446,N_8048);
or U9808 (N_9808,N_8270,N_8981);
nor U9809 (N_9809,N_8644,N_8153);
nor U9810 (N_9810,N_8663,N_8480);
or U9811 (N_9811,N_8782,N_8752);
nor U9812 (N_9812,N_8893,N_8108);
nor U9813 (N_9813,N_8074,N_8784);
or U9814 (N_9814,N_8924,N_8102);
and U9815 (N_9815,N_8370,N_8864);
or U9816 (N_9816,N_8894,N_8642);
nand U9817 (N_9817,N_8686,N_8142);
or U9818 (N_9818,N_8513,N_8768);
nor U9819 (N_9819,N_8289,N_8863);
nor U9820 (N_9820,N_8568,N_8880);
and U9821 (N_9821,N_8650,N_8965);
nor U9822 (N_9822,N_8327,N_8843);
nand U9823 (N_9823,N_8659,N_8461);
or U9824 (N_9824,N_8021,N_8315);
and U9825 (N_9825,N_8434,N_8382);
nor U9826 (N_9826,N_8593,N_8887);
and U9827 (N_9827,N_8250,N_8022);
or U9828 (N_9828,N_8276,N_8845);
nand U9829 (N_9829,N_8964,N_8230);
or U9830 (N_9830,N_8383,N_8711);
and U9831 (N_9831,N_8929,N_8875);
and U9832 (N_9832,N_8275,N_8641);
nor U9833 (N_9833,N_8197,N_8950);
or U9834 (N_9834,N_8320,N_8868);
nand U9835 (N_9835,N_8780,N_8076);
nor U9836 (N_9836,N_8966,N_8939);
nor U9837 (N_9837,N_8990,N_8211);
nor U9838 (N_9838,N_8055,N_8216);
and U9839 (N_9839,N_8048,N_8376);
and U9840 (N_9840,N_8539,N_8963);
nor U9841 (N_9841,N_8054,N_8238);
and U9842 (N_9842,N_8991,N_8786);
nor U9843 (N_9843,N_8435,N_8341);
or U9844 (N_9844,N_8498,N_8329);
or U9845 (N_9845,N_8788,N_8846);
and U9846 (N_9846,N_8628,N_8993);
nand U9847 (N_9847,N_8706,N_8996);
or U9848 (N_9848,N_8132,N_8757);
nand U9849 (N_9849,N_8696,N_8096);
or U9850 (N_9850,N_8767,N_8343);
nor U9851 (N_9851,N_8562,N_8456);
or U9852 (N_9852,N_8673,N_8345);
and U9853 (N_9853,N_8409,N_8899);
nand U9854 (N_9854,N_8890,N_8726);
nor U9855 (N_9855,N_8789,N_8763);
and U9856 (N_9856,N_8117,N_8938);
or U9857 (N_9857,N_8502,N_8886);
nor U9858 (N_9858,N_8961,N_8243);
nand U9859 (N_9859,N_8343,N_8722);
nor U9860 (N_9860,N_8238,N_8720);
and U9861 (N_9861,N_8847,N_8393);
nor U9862 (N_9862,N_8065,N_8612);
and U9863 (N_9863,N_8018,N_8064);
xnor U9864 (N_9864,N_8041,N_8090);
and U9865 (N_9865,N_8647,N_8401);
and U9866 (N_9866,N_8323,N_8005);
and U9867 (N_9867,N_8746,N_8850);
and U9868 (N_9868,N_8628,N_8370);
or U9869 (N_9869,N_8933,N_8168);
nand U9870 (N_9870,N_8724,N_8308);
and U9871 (N_9871,N_8320,N_8310);
nor U9872 (N_9872,N_8611,N_8725);
nor U9873 (N_9873,N_8858,N_8064);
and U9874 (N_9874,N_8750,N_8628);
and U9875 (N_9875,N_8368,N_8498);
and U9876 (N_9876,N_8575,N_8068);
nor U9877 (N_9877,N_8899,N_8218);
nand U9878 (N_9878,N_8634,N_8912);
and U9879 (N_9879,N_8122,N_8453);
and U9880 (N_9880,N_8535,N_8165);
nor U9881 (N_9881,N_8197,N_8199);
nor U9882 (N_9882,N_8765,N_8140);
nor U9883 (N_9883,N_8835,N_8317);
and U9884 (N_9884,N_8118,N_8622);
or U9885 (N_9885,N_8300,N_8802);
or U9886 (N_9886,N_8385,N_8246);
nor U9887 (N_9887,N_8585,N_8786);
or U9888 (N_9888,N_8966,N_8856);
or U9889 (N_9889,N_8461,N_8481);
and U9890 (N_9890,N_8880,N_8454);
or U9891 (N_9891,N_8753,N_8931);
nand U9892 (N_9892,N_8964,N_8664);
and U9893 (N_9893,N_8866,N_8360);
and U9894 (N_9894,N_8660,N_8740);
nand U9895 (N_9895,N_8503,N_8563);
nor U9896 (N_9896,N_8020,N_8275);
and U9897 (N_9897,N_8386,N_8642);
and U9898 (N_9898,N_8419,N_8874);
nor U9899 (N_9899,N_8238,N_8899);
nand U9900 (N_9900,N_8830,N_8094);
and U9901 (N_9901,N_8015,N_8493);
nand U9902 (N_9902,N_8398,N_8092);
and U9903 (N_9903,N_8588,N_8776);
or U9904 (N_9904,N_8279,N_8610);
nor U9905 (N_9905,N_8731,N_8289);
and U9906 (N_9906,N_8565,N_8285);
or U9907 (N_9907,N_8029,N_8384);
nand U9908 (N_9908,N_8028,N_8123);
and U9909 (N_9909,N_8501,N_8833);
nor U9910 (N_9910,N_8173,N_8592);
xor U9911 (N_9911,N_8670,N_8796);
or U9912 (N_9912,N_8757,N_8060);
nor U9913 (N_9913,N_8126,N_8082);
nand U9914 (N_9914,N_8539,N_8015);
or U9915 (N_9915,N_8599,N_8533);
and U9916 (N_9916,N_8939,N_8237);
xor U9917 (N_9917,N_8274,N_8351);
nand U9918 (N_9918,N_8646,N_8963);
and U9919 (N_9919,N_8488,N_8938);
and U9920 (N_9920,N_8495,N_8095);
or U9921 (N_9921,N_8756,N_8430);
nand U9922 (N_9922,N_8170,N_8189);
and U9923 (N_9923,N_8423,N_8903);
or U9924 (N_9924,N_8906,N_8244);
nor U9925 (N_9925,N_8103,N_8986);
nand U9926 (N_9926,N_8662,N_8546);
nor U9927 (N_9927,N_8452,N_8473);
nor U9928 (N_9928,N_8215,N_8647);
and U9929 (N_9929,N_8019,N_8393);
nand U9930 (N_9930,N_8935,N_8107);
nor U9931 (N_9931,N_8351,N_8032);
and U9932 (N_9932,N_8037,N_8766);
nor U9933 (N_9933,N_8251,N_8839);
nand U9934 (N_9934,N_8039,N_8168);
or U9935 (N_9935,N_8029,N_8327);
nand U9936 (N_9936,N_8847,N_8198);
nand U9937 (N_9937,N_8027,N_8695);
or U9938 (N_9938,N_8025,N_8712);
and U9939 (N_9939,N_8001,N_8492);
or U9940 (N_9940,N_8489,N_8468);
or U9941 (N_9941,N_8315,N_8111);
and U9942 (N_9942,N_8385,N_8187);
nand U9943 (N_9943,N_8275,N_8705);
nand U9944 (N_9944,N_8085,N_8067);
nor U9945 (N_9945,N_8854,N_8026);
and U9946 (N_9946,N_8391,N_8284);
and U9947 (N_9947,N_8280,N_8587);
and U9948 (N_9948,N_8288,N_8017);
nor U9949 (N_9949,N_8176,N_8534);
nand U9950 (N_9950,N_8676,N_8010);
or U9951 (N_9951,N_8336,N_8541);
or U9952 (N_9952,N_8287,N_8461);
or U9953 (N_9953,N_8066,N_8362);
nand U9954 (N_9954,N_8616,N_8274);
or U9955 (N_9955,N_8927,N_8154);
nor U9956 (N_9956,N_8235,N_8368);
nor U9957 (N_9957,N_8094,N_8516);
and U9958 (N_9958,N_8508,N_8530);
nand U9959 (N_9959,N_8203,N_8189);
and U9960 (N_9960,N_8495,N_8547);
and U9961 (N_9961,N_8011,N_8546);
or U9962 (N_9962,N_8341,N_8437);
nor U9963 (N_9963,N_8761,N_8619);
and U9964 (N_9964,N_8672,N_8740);
nor U9965 (N_9965,N_8949,N_8364);
and U9966 (N_9966,N_8368,N_8429);
nand U9967 (N_9967,N_8694,N_8487);
xnor U9968 (N_9968,N_8646,N_8895);
nand U9969 (N_9969,N_8076,N_8404);
or U9970 (N_9970,N_8250,N_8544);
and U9971 (N_9971,N_8025,N_8575);
nor U9972 (N_9972,N_8119,N_8764);
or U9973 (N_9973,N_8334,N_8926);
and U9974 (N_9974,N_8874,N_8780);
and U9975 (N_9975,N_8311,N_8648);
or U9976 (N_9976,N_8013,N_8722);
or U9977 (N_9977,N_8679,N_8068);
xor U9978 (N_9978,N_8392,N_8579);
nor U9979 (N_9979,N_8664,N_8333);
nand U9980 (N_9980,N_8417,N_8105);
and U9981 (N_9981,N_8658,N_8038);
nand U9982 (N_9982,N_8964,N_8415);
nor U9983 (N_9983,N_8696,N_8175);
nor U9984 (N_9984,N_8933,N_8210);
nand U9985 (N_9985,N_8263,N_8437);
and U9986 (N_9986,N_8076,N_8099);
and U9987 (N_9987,N_8466,N_8131);
or U9988 (N_9988,N_8362,N_8593);
nor U9989 (N_9989,N_8155,N_8773);
or U9990 (N_9990,N_8340,N_8229);
or U9991 (N_9991,N_8000,N_8480);
and U9992 (N_9992,N_8042,N_8134);
or U9993 (N_9993,N_8932,N_8962);
nor U9994 (N_9994,N_8888,N_8770);
nor U9995 (N_9995,N_8409,N_8679);
nand U9996 (N_9996,N_8985,N_8063);
nand U9997 (N_9997,N_8299,N_8288);
nand U9998 (N_9998,N_8234,N_8249);
and U9999 (N_9999,N_8135,N_8110);
nor UO_0 (O_0,N_9803,N_9569);
or UO_1 (O_1,N_9830,N_9339);
and UO_2 (O_2,N_9831,N_9291);
and UO_3 (O_3,N_9510,N_9144);
or UO_4 (O_4,N_9108,N_9813);
or UO_5 (O_5,N_9231,N_9160);
or UO_6 (O_6,N_9701,N_9725);
or UO_7 (O_7,N_9362,N_9804);
or UO_8 (O_8,N_9364,N_9507);
and UO_9 (O_9,N_9734,N_9678);
and UO_10 (O_10,N_9002,N_9748);
nand UO_11 (O_11,N_9642,N_9083);
and UO_12 (O_12,N_9590,N_9959);
nand UO_13 (O_13,N_9630,N_9110);
nand UO_14 (O_14,N_9694,N_9553);
and UO_15 (O_15,N_9352,N_9326);
nor UO_16 (O_16,N_9320,N_9226);
and UO_17 (O_17,N_9312,N_9723);
or UO_18 (O_18,N_9600,N_9764);
nor UO_19 (O_19,N_9202,N_9861);
or UO_20 (O_20,N_9969,N_9404);
or UO_21 (O_21,N_9473,N_9766);
or UO_22 (O_22,N_9490,N_9011);
or UO_23 (O_23,N_9058,N_9325);
nor UO_24 (O_24,N_9900,N_9797);
nand UO_25 (O_25,N_9172,N_9494);
and UO_26 (O_26,N_9495,N_9342);
or UO_27 (O_27,N_9169,N_9407);
and UO_28 (O_28,N_9760,N_9999);
or UO_29 (O_29,N_9469,N_9755);
and UO_30 (O_30,N_9781,N_9433);
or UO_31 (O_31,N_9982,N_9016);
nor UO_32 (O_32,N_9387,N_9513);
and UO_33 (O_33,N_9220,N_9731);
nand UO_34 (O_34,N_9155,N_9647);
and UO_35 (O_35,N_9257,N_9145);
nand UO_36 (O_36,N_9921,N_9782);
and UO_37 (O_37,N_9898,N_9233);
nand UO_38 (O_38,N_9613,N_9099);
or UO_39 (O_39,N_9120,N_9255);
or UO_40 (O_40,N_9902,N_9078);
nand UO_41 (O_41,N_9640,N_9281);
or UO_42 (O_42,N_9182,N_9164);
nand UO_43 (O_43,N_9081,N_9392);
xnor UO_44 (O_44,N_9505,N_9103);
or UO_45 (O_45,N_9137,N_9873);
nand UO_46 (O_46,N_9771,N_9024);
nor UO_47 (O_47,N_9915,N_9747);
nand UO_48 (O_48,N_9534,N_9034);
nand UO_49 (O_49,N_9390,N_9159);
nor UO_50 (O_50,N_9882,N_9268);
nand UO_51 (O_51,N_9406,N_9643);
and UO_52 (O_52,N_9295,N_9558);
and UO_53 (O_53,N_9128,N_9323);
and UO_54 (O_54,N_9129,N_9153);
and UO_55 (O_55,N_9179,N_9043);
nor UO_56 (O_56,N_9267,N_9874);
and UO_57 (O_57,N_9814,N_9181);
nor UO_58 (O_58,N_9920,N_9437);
nand UO_59 (O_59,N_9062,N_9464);
nand UO_60 (O_60,N_9310,N_9089);
or UO_61 (O_61,N_9798,N_9366);
nand UO_62 (O_62,N_9113,N_9971);
nand UO_63 (O_63,N_9676,N_9588);
or UO_64 (O_64,N_9041,N_9822);
xor UO_65 (O_65,N_9991,N_9355);
and UO_66 (O_66,N_9250,N_9708);
nor UO_67 (O_67,N_9865,N_9492);
nor UO_68 (O_68,N_9662,N_9562);
nor UO_69 (O_69,N_9005,N_9953);
and UO_70 (O_70,N_9358,N_9141);
nor UO_71 (O_71,N_9488,N_9270);
nor UO_72 (O_72,N_9401,N_9092);
or UO_73 (O_73,N_9879,N_9330);
and UO_74 (O_74,N_9857,N_9703);
and UO_75 (O_75,N_9225,N_9173);
nor UO_76 (O_76,N_9934,N_9810);
nor UO_77 (O_77,N_9974,N_9065);
nand UO_78 (O_78,N_9875,N_9780);
or UO_79 (O_79,N_9858,N_9462);
nand UO_80 (O_80,N_9637,N_9080);
and UO_81 (O_81,N_9891,N_9009);
nor UO_82 (O_82,N_9393,N_9408);
nor UO_83 (O_83,N_9795,N_9936);
nor UO_84 (O_84,N_9787,N_9540);
nor UO_85 (O_85,N_9333,N_9596);
nor UO_86 (O_86,N_9026,N_9014);
nor UO_87 (O_87,N_9612,N_9232);
nand UO_88 (O_88,N_9792,N_9204);
nor UO_89 (O_89,N_9163,N_9086);
nor UO_90 (O_90,N_9463,N_9881);
nor UO_91 (O_91,N_9894,N_9631);
or UO_92 (O_92,N_9811,N_9504);
or UO_93 (O_93,N_9743,N_9100);
nand UO_94 (O_94,N_9728,N_9947);
nor UO_95 (O_95,N_9605,N_9962);
and UO_96 (O_96,N_9668,N_9876);
and UO_97 (O_97,N_9691,N_9314);
nor UO_98 (O_98,N_9402,N_9863);
xor UO_99 (O_99,N_9796,N_9308);
nor UO_100 (O_100,N_9719,N_9574);
nor UO_101 (O_101,N_9253,N_9130);
nor UO_102 (O_102,N_9745,N_9298);
nor UO_103 (O_103,N_9721,N_9101);
or UO_104 (O_104,N_9430,N_9154);
or UO_105 (O_105,N_9967,N_9859);
or UO_106 (O_106,N_9617,N_9475);
nand UO_107 (O_107,N_9122,N_9059);
and UO_108 (O_108,N_9531,N_9357);
and UO_109 (O_109,N_9292,N_9116);
and UO_110 (O_110,N_9055,N_9950);
and UO_111 (O_111,N_9907,N_9580);
or UO_112 (O_112,N_9530,N_9335);
or UO_113 (O_113,N_9709,N_9935);
nand UO_114 (O_114,N_9658,N_9761);
nor UO_115 (O_115,N_9618,N_9966);
nor UO_116 (O_116,N_9987,N_9832);
xnor UO_117 (O_117,N_9178,N_9854);
nand UO_118 (O_118,N_9884,N_9177);
and UO_119 (O_119,N_9757,N_9560);
or UO_120 (O_120,N_9478,N_9542);
and UO_121 (O_121,N_9415,N_9697);
or UO_122 (O_122,N_9443,N_9954);
nand UO_123 (O_123,N_9050,N_9125);
and UO_124 (O_124,N_9603,N_9886);
and UO_125 (O_125,N_9968,N_9940);
or UO_126 (O_126,N_9910,N_9517);
and UO_127 (O_127,N_9418,N_9274);
nand UO_128 (O_128,N_9946,N_9664);
nor UO_129 (O_129,N_9399,N_9850);
or UO_130 (O_130,N_9245,N_9397);
nand UO_131 (O_131,N_9503,N_9369);
and UO_132 (O_132,N_9783,N_9692);
or UO_133 (O_133,N_9571,N_9821);
nand UO_134 (O_134,N_9230,N_9459);
nand UO_135 (O_135,N_9114,N_9975);
nor UO_136 (O_136,N_9944,N_9147);
nand UO_137 (O_137,N_9716,N_9301);
or UO_138 (O_138,N_9727,N_9575);
and UO_139 (O_139,N_9460,N_9284);
nor UO_140 (O_140,N_9029,N_9604);
xor UO_141 (O_141,N_9895,N_9527);
or UO_142 (O_142,N_9749,N_9076);
and UO_143 (O_143,N_9998,N_9012);
nor UO_144 (O_144,N_9309,N_9023);
nand UO_145 (O_145,N_9218,N_9396);
nand UO_146 (O_146,N_9579,N_9428);
nor UO_147 (O_147,N_9941,N_9567);
or UO_148 (O_148,N_9679,N_9649);
nor UO_149 (O_149,N_9511,N_9037);
and UO_150 (O_150,N_9269,N_9445);
or UO_151 (O_151,N_9119,N_9389);
nor UO_152 (O_152,N_9931,N_9045);
and UO_153 (O_153,N_9261,N_9289);
or UO_154 (O_154,N_9509,N_9138);
and UO_155 (O_155,N_9514,N_9619);
nor UO_156 (O_156,N_9240,N_9834);
and UO_157 (O_157,N_9949,N_9121);
or UO_158 (O_158,N_9887,N_9526);
nand UO_159 (O_159,N_9123,N_9450);
nand UO_160 (O_160,N_9072,N_9677);
nand UO_161 (O_161,N_9115,N_9290);
or UO_162 (O_162,N_9238,N_9102);
nor UO_163 (O_163,N_9484,N_9652);
nor UO_164 (O_164,N_9550,N_9572);
or UO_165 (O_165,N_9251,N_9582);
nor UO_166 (O_166,N_9805,N_9318);
nor UO_167 (O_167,N_9090,N_9063);
or UO_168 (O_168,N_9243,N_9278);
nor UO_169 (O_169,N_9151,N_9215);
or UO_170 (O_170,N_9897,N_9791);
and UO_171 (O_171,N_9801,N_9197);
nor UO_172 (O_172,N_9471,N_9223);
nand UO_173 (O_173,N_9586,N_9273);
nor UO_174 (O_174,N_9918,N_9939);
and UO_175 (O_175,N_9221,N_9316);
and UO_176 (O_176,N_9321,N_9127);
and UO_177 (O_177,N_9786,N_9768);
nand UO_178 (O_178,N_9200,N_9807);
and UO_179 (O_179,N_9093,N_9061);
and UO_180 (O_180,N_9790,N_9075);
or UO_181 (O_181,N_9539,N_9970);
nor UO_182 (O_182,N_9070,N_9555);
and UO_183 (O_183,N_9167,N_9046);
or UO_184 (O_184,N_9247,N_9265);
and UO_185 (O_185,N_9754,N_9957);
or UO_186 (O_186,N_9239,N_9585);
nor UO_187 (O_187,N_9903,N_9104);
or UO_188 (O_188,N_9106,N_9933);
nor UO_189 (O_189,N_9922,N_9565);
and UO_190 (O_190,N_9844,N_9979);
nand UO_191 (O_191,N_9248,N_9896);
nand UO_192 (O_192,N_9906,N_9729);
and UO_193 (O_193,N_9688,N_9563);
or UO_194 (O_194,N_9961,N_9327);
nor UO_195 (O_195,N_9964,N_9126);
xnor UO_196 (O_196,N_9136,N_9978);
or UO_197 (O_197,N_9280,N_9395);
nand UO_198 (O_198,N_9758,N_9942);
nor UO_199 (O_199,N_9071,N_9332);
and UO_200 (O_200,N_9623,N_9347);
nand UO_201 (O_201,N_9673,N_9271);
and UO_202 (O_202,N_9930,N_9343);
nand UO_203 (O_203,N_9235,N_9328);
nand UO_204 (O_204,N_9837,N_9912);
nand UO_205 (O_205,N_9105,N_9717);
nor UO_206 (O_206,N_9480,N_9763);
and UO_207 (O_207,N_9094,N_9213);
or UO_208 (O_208,N_9589,N_9435);
and UO_209 (O_209,N_9194,N_9502);
or UO_210 (O_210,N_9338,N_9685);
xor UO_211 (O_211,N_9913,N_9568);
or UO_212 (O_212,N_9520,N_9909);
or UO_213 (O_213,N_9756,N_9442);
nor UO_214 (O_214,N_9833,N_9241);
and UO_215 (O_215,N_9340,N_9955);
nor UO_216 (O_216,N_9234,N_9146);
and UO_217 (O_217,N_9789,N_9726);
and UO_218 (O_218,N_9373,N_9557);
nand UO_219 (O_219,N_9282,N_9952);
and UO_220 (O_220,N_9965,N_9324);
nor UO_221 (O_221,N_9730,N_9537);
and UO_222 (O_222,N_9995,N_9224);
and UO_223 (O_223,N_9482,N_9926);
or UO_224 (O_224,N_9047,N_9622);
or UO_225 (O_225,N_9535,N_9650);
nand UO_226 (O_226,N_9470,N_9044);
or UO_227 (O_227,N_9293,N_9827);
nand UO_228 (O_228,N_9776,N_9707);
nor UO_229 (O_229,N_9523,N_9824);
and UO_230 (O_230,N_9158,N_9772);
nor UO_231 (O_231,N_9350,N_9739);
nand UO_232 (O_232,N_9483,N_9107);
and UO_233 (O_233,N_9860,N_9162);
nor UO_234 (O_234,N_9455,N_9751);
and UO_235 (O_235,N_9413,N_9744);
nor UO_236 (O_236,N_9015,N_9544);
xnor UO_237 (O_237,N_9489,N_9032);
and UO_238 (O_238,N_9191,N_9476);
and UO_239 (O_239,N_9485,N_9746);
nand UO_240 (O_240,N_9778,N_9246);
nand UO_241 (O_241,N_9254,N_9963);
nor UO_242 (O_242,N_9187,N_9140);
nand UO_243 (O_243,N_9997,N_9356);
nor UO_244 (O_244,N_9020,N_9607);
nor UO_245 (O_245,N_9769,N_9938);
nand UO_246 (O_246,N_9199,N_9111);
nand UO_247 (O_247,N_9411,N_9227);
nor UO_248 (O_248,N_9210,N_9412);
or UO_249 (O_249,N_9663,N_9917);
and UO_250 (O_250,N_9381,N_9275);
nand UO_251 (O_251,N_9989,N_9515);
and UO_252 (O_252,N_9570,N_9219);
or UO_253 (O_253,N_9417,N_9904);
and UO_254 (O_254,N_9852,N_9519);
and UO_255 (O_255,N_9304,N_9767);
or UO_256 (O_256,N_9846,N_9712);
nand UO_257 (O_257,N_9626,N_9168);
xnor UO_258 (O_258,N_9862,N_9665);
nand UO_259 (O_259,N_9845,N_9561);
or UO_260 (O_260,N_9698,N_9436);
nor UO_261 (O_261,N_9983,N_9131);
and UO_262 (O_262,N_9752,N_9710);
nand UO_263 (O_263,N_9217,N_9262);
and UO_264 (O_264,N_9583,N_9578);
nor UO_265 (O_265,N_9943,N_9774);
and UO_266 (O_266,N_9236,N_9336);
nor UO_267 (O_267,N_9693,N_9735);
nand UO_268 (O_268,N_9960,N_9244);
and UO_269 (O_269,N_9499,N_9048);
xnor UO_270 (O_270,N_9378,N_9205);
and UO_271 (O_271,N_9715,N_9806);
and UO_272 (O_272,N_9890,N_9359);
or UO_273 (O_273,N_9036,N_9452);
nand UO_274 (O_274,N_9263,N_9670);
or UO_275 (O_275,N_9928,N_9867);
nor UO_276 (O_276,N_9564,N_9405);
nor UO_277 (O_277,N_9815,N_9165);
xor UO_278 (O_278,N_9932,N_9714);
and UO_279 (O_279,N_9671,N_9142);
nor UO_280 (O_280,N_9360,N_9004);
nor UO_281 (O_281,N_9628,N_9276);
or UO_282 (O_282,N_9028,N_9214);
or UO_283 (O_283,N_9195,N_9367);
or UO_284 (O_284,N_9283,N_9299);
nand UO_285 (O_285,N_9646,N_9741);
and UO_286 (O_286,N_9908,N_9419);
nor UO_287 (O_287,N_9272,N_9541);
nor UO_288 (O_288,N_9866,N_9054);
or UO_289 (O_289,N_9666,N_9794);
or UO_290 (O_290,N_9878,N_9883);
or UO_291 (O_291,N_9302,N_9064);
or UO_292 (O_292,N_9929,N_9980);
and UO_293 (O_293,N_9351,N_9809);
nor UO_294 (O_294,N_9724,N_9872);
nand UO_295 (O_295,N_9538,N_9258);
nand UO_296 (O_296,N_9681,N_9545);
or UO_297 (O_297,N_9069,N_9669);
nor UO_298 (O_298,N_9374,N_9958);
and UO_299 (O_299,N_9148,N_9098);
nor UO_300 (O_300,N_9458,N_9423);
nand UO_301 (O_301,N_9348,N_9410);
and UO_302 (O_302,N_9639,N_9134);
and UO_303 (O_303,N_9429,N_9638);
nand UO_304 (O_304,N_9259,N_9161);
nand UO_305 (O_305,N_9157,N_9775);
or UO_306 (O_306,N_9587,N_9923);
nand UO_307 (O_307,N_9117,N_9656);
nor UO_308 (O_308,N_9888,N_9184);
or UO_309 (O_309,N_9644,N_9152);
nor UO_310 (O_310,N_9512,N_9424);
nor UO_311 (O_311,N_9819,N_9740);
nor UO_312 (O_312,N_9493,N_9889);
nor UO_313 (O_313,N_9013,N_9864);
nand UO_314 (O_314,N_9203,N_9385);
and UO_315 (O_315,N_9529,N_9851);
and UO_316 (O_316,N_9421,N_9087);
or UO_317 (O_317,N_9633,N_9427);
xnor UO_318 (O_318,N_9547,N_9657);
and UO_319 (O_319,N_9474,N_9193);
nand UO_320 (O_320,N_9597,N_9174);
or UO_321 (O_321,N_9322,N_9277);
nor UO_322 (O_322,N_9695,N_9085);
nor UO_323 (O_323,N_9361,N_9892);
nor UO_324 (O_324,N_9409,N_9143);
and UO_325 (O_325,N_9847,N_9438);
nor UO_326 (O_326,N_9525,N_9440);
and UO_327 (O_327,N_9593,N_9479);
nand UO_328 (O_328,N_9853,N_9993);
nand UO_329 (O_329,N_9738,N_9190);
nor UO_330 (O_330,N_9311,N_9635);
or UO_331 (O_331,N_9003,N_9208);
nand UO_332 (O_332,N_9901,N_9508);
nand UO_333 (O_333,N_9305,N_9486);
nand UO_334 (O_334,N_9759,N_9687);
nand UO_335 (O_335,N_9856,N_9077);
nor UO_336 (O_336,N_9842,N_9264);
xor UO_337 (O_337,N_9848,N_9216);
nand UO_338 (O_338,N_9109,N_9300);
nand UO_339 (O_339,N_9288,N_9266);
nand UO_340 (O_340,N_9286,N_9849);
or UO_341 (O_341,N_9212,N_9285);
or UO_342 (O_342,N_9431,N_9648);
nand UO_343 (O_343,N_9711,N_9051);
or UO_344 (O_344,N_9880,N_9770);
and UO_345 (O_345,N_9592,N_9307);
nand UO_346 (O_346,N_9654,N_9672);
nand UO_347 (O_347,N_9765,N_9820);
or UO_348 (O_348,N_9802,N_9398);
and UO_349 (O_349,N_9491,N_9344);
nor UO_350 (O_350,N_9426,N_9006);
or UO_351 (O_351,N_9990,N_9602);
or UO_352 (O_352,N_9074,N_9737);
and UO_353 (O_353,N_9893,N_9546);
nor UO_354 (O_354,N_9988,N_9713);
nor UO_355 (O_355,N_9595,N_9391);
nor UO_356 (O_356,N_9451,N_9793);
nand UO_357 (O_357,N_9441,N_9388);
and UO_358 (O_358,N_9718,N_9185);
nor UO_359 (O_359,N_9675,N_9722);
or UO_360 (O_360,N_9186,N_9466);
and UO_361 (O_361,N_9838,N_9655);
or UO_362 (O_362,N_9835,N_9620);
nand UO_363 (O_363,N_9825,N_9616);
nor UO_364 (O_364,N_9461,N_9702);
or UO_365 (O_365,N_9196,N_9035);
or UO_366 (O_366,N_9610,N_9403);
and UO_367 (O_367,N_9641,N_9532);
or UO_368 (O_368,N_9319,N_9629);
or UO_369 (O_369,N_9924,N_9449);
xor UO_370 (O_370,N_9294,N_9249);
nand UO_371 (O_371,N_9189,N_9981);
or UO_372 (O_372,N_9624,N_9543);
nor UO_373 (O_373,N_9287,N_9383);
or UO_374 (O_374,N_9150,N_9201);
nand UO_375 (O_375,N_9334,N_9384);
nand UO_376 (O_376,N_9700,N_9368);
nor UO_377 (O_377,N_9501,N_9132);
nand UO_378 (O_378,N_9000,N_9448);
and UO_379 (O_379,N_9315,N_9010);
or UO_380 (O_380,N_9481,N_9400);
nand UO_381 (O_381,N_9683,N_9581);
nand UO_382 (O_382,N_9198,N_9779);
and UO_383 (O_383,N_9454,N_9736);
and UO_384 (O_384,N_9506,N_9773);
nor UO_385 (O_385,N_9973,N_9927);
nand UO_386 (O_386,N_9533,N_9341);
and UO_387 (O_387,N_9056,N_9945);
nor UO_388 (O_388,N_9033,N_9500);
nand UO_389 (O_389,N_9422,N_9986);
nand UO_390 (O_390,N_9828,N_9139);
and UO_391 (O_391,N_9948,N_9660);
and UO_392 (O_392,N_9183,N_9097);
nor UO_393 (O_393,N_9042,N_9812);
or UO_394 (O_394,N_9079,N_9799);
nor UO_395 (O_395,N_9135,N_9733);
or UO_396 (O_396,N_9925,N_9001);
or UO_397 (O_397,N_9996,N_9528);
nor UO_398 (O_398,N_9937,N_9313);
nand UO_399 (O_399,N_9008,N_9674);
nand UO_400 (O_400,N_9052,N_9031);
or UO_401 (O_401,N_9636,N_9518);
nand UO_402 (O_402,N_9088,N_9591);
or UO_403 (O_403,N_9432,N_9084);
or UO_404 (O_404,N_9554,N_9653);
or UO_405 (O_405,N_9615,N_9256);
or UO_406 (O_406,N_9742,N_9175);
nand UO_407 (O_407,N_9073,N_9696);
and UO_408 (O_408,N_9021,N_9349);
and UO_409 (O_409,N_9599,N_9380);
and UO_410 (O_410,N_9446,N_9447);
xnor UO_411 (O_411,N_9498,N_9049);
and UO_412 (O_412,N_9839,N_9855);
nor UO_413 (O_413,N_9420,N_9170);
nand UO_414 (O_414,N_9207,N_9686);
and UO_415 (O_415,N_9222,N_9497);
or UO_416 (O_416,N_9386,N_9180);
nand UO_417 (O_417,N_9372,N_9329);
and UO_418 (O_418,N_9379,N_9375);
and UO_419 (O_419,N_9377,N_9577);
and UO_420 (O_420,N_9818,N_9345);
and UO_421 (O_421,N_9704,N_9689);
or UO_422 (O_422,N_9522,N_9549);
nand UO_423 (O_423,N_9598,N_9027);
nor UO_424 (O_424,N_9477,N_9788);
and UO_425 (O_425,N_9661,N_9784);
nand UO_426 (O_426,N_9156,N_9331);
nand UO_427 (O_427,N_9030,N_9346);
nand UO_428 (O_428,N_9611,N_9840);
nand UO_429 (O_429,N_9038,N_9053);
nor UO_430 (O_430,N_9019,N_9576);
xnor UO_431 (O_431,N_9211,N_9584);
nand UO_432 (O_432,N_9536,N_9133);
or UO_433 (O_433,N_9777,N_9868);
or UO_434 (O_434,N_9039,N_9303);
nor UO_435 (O_435,N_9609,N_9209);
nand UO_436 (O_436,N_9800,N_9206);
nand UO_437 (O_437,N_9192,N_9453);
nand UO_438 (O_438,N_9066,N_9750);
or UO_439 (O_439,N_9594,N_9634);
and UO_440 (O_440,N_9376,N_9705);
or UO_441 (O_441,N_9124,N_9785);
nand UO_442 (O_442,N_9706,N_9972);
and UO_443 (O_443,N_9306,N_9457);
or UO_444 (O_444,N_9118,N_9425);
nand UO_445 (O_445,N_9371,N_9188);
nor UO_446 (O_446,N_9916,N_9911);
and UO_447 (O_447,N_9817,N_9025);
or UO_448 (O_448,N_9496,N_9467);
xnor UO_449 (O_449,N_9521,N_9516);
and UO_450 (O_450,N_9951,N_9699);
nor UO_451 (O_451,N_9057,N_9022);
or UO_452 (O_452,N_9753,N_9091);
nand UO_453 (O_453,N_9556,N_9354);
nor UO_454 (O_454,N_9439,N_9808);
and UO_455 (O_455,N_9487,N_9228);
and UO_456 (O_456,N_9524,N_9018);
nor UO_457 (O_457,N_9608,N_9552);
nor UO_458 (O_458,N_9444,N_9353);
nor UO_459 (O_459,N_9994,N_9682);
nand UO_460 (O_460,N_9870,N_9548);
or UO_461 (O_461,N_9465,N_9472);
and UO_462 (O_462,N_9551,N_9667);
nand UO_463 (O_463,N_9242,N_9680);
nor UO_464 (O_464,N_9919,N_9296);
or UO_465 (O_465,N_9252,N_9977);
or UO_466 (O_466,N_9017,N_9720);
nor UO_467 (O_467,N_9229,N_9614);
and UO_468 (O_468,N_9068,N_9826);
nor UO_469 (O_469,N_9082,N_9007);
and UO_470 (O_470,N_9985,N_9651);
nor UO_471 (O_471,N_9690,N_9762);
and UO_472 (O_472,N_9414,N_9984);
nor UO_473 (O_473,N_9877,N_9468);
and UO_474 (O_474,N_9237,N_9166);
or UO_475 (O_475,N_9394,N_9871);
nand UO_476 (O_476,N_9260,N_9095);
nor UO_477 (O_477,N_9632,N_9416);
or UO_478 (O_478,N_9096,N_9816);
nand UO_479 (O_479,N_9365,N_9829);
or UO_480 (O_480,N_9956,N_9836);
and UO_481 (O_481,N_9434,N_9040);
nor UO_482 (O_482,N_9684,N_9370);
or UO_483 (O_483,N_9112,N_9841);
or UO_484 (O_484,N_9914,N_9606);
or UO_485 (O_485,N_9823,N_9659);
nor UO_486 (O_486,N_9625,N_9573);
nand UO_487 (O_487,N_9060,N_9732);
nand UO_488 (O_488,N_9456,N_9176);
nand UO_489 (O_489,N_9337,N_9645);
or UO_490 (O_490,N_9382,N_9869);
and UO_491 (O_491,N_9976,N_9559);
and UO_492 (O_492,N_9885,N_9566);
nor UO_493 (O_493,N_9992,N_9317);
nand UO_494 (O_494,N_9899,N_9067);
nand UO_495 (O_495,N_9601,N_9297);
nor UO_496 (O_496,N_9621,N_9363);
nor UO_497 (O_497,N_9905,N_9279);
nor UO_498 (O_498,N_9843,N_9627);
nor UO_499 (O_499,N_9149,N_9171);
nor UO_500 (O_500,N_9342,N_9611);
nand UO_501 (O_501,N_9346,N_9108);
nand UO_502 (O_502,N_9143,N_9922);
or UO_503 (O_503,N_9970,N_9664);
nand UO_504 (O_504,N_9112,N_9755);
or UO_505 (O_505,N_9853,N_9371);
nor UO_506 (O_506,N_9803,N_9851);
and UO_507 (O_507,N_9136,N_9626);
or UO_508 (O_508,N_9478,N_9177);
or UO_509 (O_509,N_9333,N_9447);
nor UO_510 (O_510,N_9391,N_9489);
nand UO_511 (O_511,N_9439,N_9494);
or UO_512 (O_512,N_9275,N_9521);
nor UO_513 (O_513,N_9204,N_9220);
nand UO_514 (O_514,N_9265,N_9378);
or UO_515 (O_515,N_9142,N_9035);
or UO_516 (O_516,N_9675,N_9531);
or UO_517 (O_517,N_9698,N_9411);
nor UO_518 (O_518,N_9797,N_9597);
nand UO_519 (O_519,N_9486,N_9190);
and UO_520 (O_520,N_9782,N_9627);
nand UO_521 (O_521,N_9596,N_9739);
and UO_522 (O_522,N_9745,N_9452);
and UO_523 (O_523,N_9992,N_9426);
and UO_524 (O_524,N_9460,N_9837);
or UO_525 (O_525,N_9413,N_9288);
or UO_526 (O_526,N_9830,N_9422);
or UO_527 (O_527,N_9749,N_9950);
nand UO_528 (O_528,N_9028,N_9807);
nand UO_529 (O_529,N_9746,N_9157);
nor UO_530 (O_530,N_9191,N_9500);
or UO_531 (O_531,N_9081,N_9157);
and UO_532 (O_532,N_9409,N_9799);
nor UO_533 (O_533,N_9145,N_9190);
xnor UO_534 (O_534,N_9207,N_9771);
nor UO_535 (O_535,N_9711,N_9154);
nand UO_536 (O_536,N_9241,N_9270);
and UO_537 (O_537,N_9831,N_9772);
and UO_538 (O_538,N_9798,N_9337);
and UO_539 (O_539,N_9514,N_9786);
nor UO_540 (O_540,N_9942,N_9174);
and UO_541 (O_541,N_9835,N_9636);
xnor UO_542 (O_542,N_9955,N_9182);
and UO_543 (O_543,N_9344,N_9830);
nor UO_544 (O_544,N_9790,N_9709);
and UO_545 (O_545,N_9391,N_9221);
nor UO_546 (O_546,N_9418,N_9810);
and UO_547 (O_547,N_9247,N_9306);
xnor UO_548 (O_548,N_9676,N_9234);
nand UO_549 (O_549,N_9467,N_9874);
and UO_550 (O_550,N_9674,N_9227);
and UO_551 (O_551,N_9593,N_9528);
or UO_552 (O_552,N_9797,N_9643);
and UO_553 (O_553,N_9552,N_9277);
or UO_554 (O_554,N_9488,N_9792);
or UO_555 (O_555,N_9248,N_9672);
and UO_556 (O_556,N_9156,N_9027);
or UO_557 (O_557,N_9975,N_9264);
and UO_558 (O_558,N_9669,N_9311);
xnor UO_559 (O_559,N_9306,N_9582);
nor UO_560 (O_560,N_9392,N_9540);
or UO_561 (O_561,N_9967,N_9332);
nor UO_562 (O_562,N_9683,N_9436);
and UO_563 (O_563,N_9280,N_9726);
and UO_564 (O_564,N_9623,N_9261);
or UO_565 (O_565,N_9234,N_9165);
xnor UO_566 (O_566,N_9486,N_9207);
nand UO_567 (O_567,N_9456,N_9602);
nand UO_568 (O_568,N_9711,N_9760);
nor UO_569 (O_569,N_9318,N_9916);
and UO_570 (O_570,N_9126,N_9530);
or UO_571 (O_571,N_9760,N_9066);
and UO_572 (O_572,N_9854,N_9372);
nand UO_573 (O_573,N_9317,N_9800);
nand UO_574 (O_574,N_9076,N_9876);
nor UO_575 (O_575,N_9681,N_9481);
nand UO_576 (O_576,N_9713,N_9326);
nor UO_577 (O_577,N_9275,N_9843);
xor UO_578 (O_578,N_9158,N_9378);
or UO_579 (O_579,N_9378,N_9474);
nand UO_580 (O_580,N_9842,N_9867);
and UO_581 (O_581,N_9067,N_9143);
nor UO_582 (O_582,N_9331,N_9198);
and UO_583 (O_583,N_9610,N_9638);
nor UO_584 (O_584,N_9449,N_9069);
nor UO_585 (O_585,N_9719,N_9018);
nor UO_586 (O_586,N_9311,N_9756);
or UO_587 (O_587,N_9562,N_9093);
or UO_588 (O_588,N_9485,N_9423);
or UO_589 (O_589,N_9326,N_9773);
and UO_590 (O_590,N_9814,N_9266);
or UO_591 (O_591,N_9085,N_9162);
nand UO_592 (O_592,N_9540,N_9062);
nand UO_593 (O_593,N_9618,N_9606);
nor UO_594 (O_594,N_9121,N_9315);
or UO_595 (O_595,N_9409,N_9545);
and UO_596 (O_596,N_9279,N_9654);
and UO_597 (O_597,N_9106,N_9222);
nor UO_598 (O_598,N_9659,N_9268);
or UO_599 (O_599,N_9294,N_9788);
and UO_600 (O_600,N_9239,N_9670);
nor UO_601 (O_601,N_9032,N_9349);
or UO_602 (O_602,N_9333,N_9475);
and UO_603 (O_603,N_9507,N_9928);
or UO_604 (O_604,N_9988,N_9944);
and UO_605 (O_605,N_9198,N_9983);
or UO_606 (O_606,N_9201,N_9655);
nor UO_607 (O_607,N_9122,N_9593);
nand UO_608 (O_608,N_9185,N_9909);
and UO_609 (O_609,N_9988,N_9282);
nand UO_610 (O_610,N_9255,N_9796);
or UO_611 (O_611,N_9596,N_9648);
nor UO_612 (O_612,N_9151,N_9345);
or UO_613 (O_613,N_9111,N_9215);
nor UO_614 (O_614,N_9339,N_9947);
and UO_615 (O_615,N_9403,N_9491);
and UO_616 (O_616,N_9659,N_9740);
and UO_617 (O_617,N_9962,N_9028);
or UO_618 (O_618,N_9148,N_9677);
or UO_619 (O_619,N_9485,N_9413);
and UO_620 (O_620,N_9956,N_9095);
nor UO_621 (O_621,N_9726,N_9144);
and UO_622 (O_622,N_9117,N_9339);
nand UO_623 (O_623,N_9662,N_9230);
or UO_624 (O_624,N_9109,N_9697);
or UO_625 (O_625,N_9948,N_9998);
nor UO_626 (O_626,N_9285,N_9455);
nor UO_627 (O_627,N_9269,N_9996);
or UO_628 (O_628,N_9750,N_9622);
or UO_629 (O_629,N_9383,N_9625);
xnor UO_630 (O_630,N_9776,N_9471);
nand UO_631 (O_631,N_9029,N_9619);
nor UO_632 (O_632,N_9344,N_9441);
nor UO_633 (O_633,N_9087,N_9438);
nand UO_634 (O_634,N_9402,N_9854);
nand UO_635 (O_635,N_9463,N_9790);
nor UO_636 (O_636,N_9451,N_9005);
nand UO_637 (O_637,N_9926,N_9212);
nor UO_638 (O_638,N_9467,N_9629);
or UO_639 (O_639,N_9991,N_9058);
nor UO_640 (O_640,N_9702,N_9938);
nor UO_641 (O_641,N_9974,N_9671);
or UO_642 (O_642,N_9317,N_9853);
nor UO_643 (O_643,N_9202,N_9837);
nor UO_644 (O_644,N_9697,N_9921);
nor UO_645 (O_645,N_9949,N_9259);
nand UO_646 (O_646,N_9875,N_9913);
nand UO_647 (O_647,N_9533,N_9112);
and UO_648 (O_648,N_9231,N_9974);
nor UO_649 (O_649,N_9097,N_9854);
nor UO_650 (O_650,N_9033,N_9573);
nand UO_651 (O_651,N_9989,N_9289);
nor UO_652 (O_652,N_9306,N_9185);
nor UO_653 (O_653,N_9989,N_9087);
and UO_654 (O_654,N_9312,N_9891);
nor UO_655 (O_655,N_9093,N_9451);
nor UO_656 (O_656,N_9896,N_9330);
or UO_657 (O_657,N_9872,N_9180);
nand UO_658 (O_658,N_9738,N_9417);
and UO_659 (O_659,N_9466,N_9406);
nor UO_660 (O_660,N_9587,N_9676);
or UO_661 (O_661,N_9246,N_9860);
or UO_662 (O_662,N_9244,N_9920);
and UO_663 (O_663,N_9815,N_9185);
or UO_664 (O_664,N_9105,N_9349);
nor UO_665 (O_665,N_9285,N_9922);
nand UO_666 (O_666,N_9395,N_9682);
nand UO_667 (O_667,N_9907,N_9808);
or UO_668 (O_668,N_9401,N_9642);
and UO_669 (O_669,N_9084,N_9198);
nand UO_670 (O_670,N_9955,N_9989);
and UO_671 (O_671,N_9834,N_9924);
nor UO_672 (O_672,N_9241,N_9802);
nor UO_673 (O_673,N_9074,N_9061);
and UO_674 (O_674,N_9207,N_9550);
or UO_675 (O_675,N_9839,N_9956);
nand UO_676 (O_676,N_9708,N_9442);
xnor UO_677 (O_677,N_9046,N_9750);
nand UO_678 (O_678,N_9280,N_9598);
nor UO_679 (O_679,N_9075,N_9032);
nand UO_680 (O_680,N_9655,N_9848);
or UO_681 (O_681,N_9930,N_9989);
nand UO_682 (O_682,N_9209,N_9261);
and UO_683 (O_683,N_9559,N_9881);
or UO_684 (O_684,N_9183,N_9712);
nand UO_685 (O_685,N_9419,N_9793);
or UO_686 (O_686,N_9602,N_9319);
nor UO_687 (O_687,N_9611,N_9320);
nand UO_688 (O_688,N_9920,N_9560);
and UO_689 (O_689,N_9391,N_9648);
or UO_690 (O_690,N_9952,N_9709);
nand UO_691 (O_691,N_9367,N_9102);
nand UO_692 (O_692,N_9468,N_9416);
or UO_693 (O_693,N_9812,N_9353);
or UO_694 (O_694,N_9733,N_9954);
and UO_695 (O_695,N_9703,N_9212);
nor UO_696 (O_696,N_9163,N_9690);
nand UO_697 (O_697,N_9664,N_9392);
nor UO_698 (O_698,N_9389,N_9162);
nand UO_699 (O_699,N_9860,N_9039);
nand UO_700 (O_700,N_9703,N_9687);
or UO_701 (O_701,N_9267,N_9246);
nand UO_702 (O_702,N_9743,N_9095);
and UO_703 (O_703,N_9989,N_9736);
xor UO_704 (O_704,N_9865,N_9167);
nand UO_705 (O_705,N_9009,N_9507);
nor UO_706 (O_706,N_9630,N_9915);
nor UO_707 (O_707,N_9277,N_9386);
nor UO_708 (O_708,N_9795,N_9332);
nand UO_709 (O_709,N_9061,N_9221);
or UO_710 (O_710,N_9795,N_9313);
or UO_711 (O_711,N_9955,N_9627);
xnor UO_712 (O_712,N_9388,N_9632);
nand UO_713 (O_713,N_9744,N_9176);
and UO_714 (O_714,N_9802,N_9305);
nor UO_715 (O_715,N_9043,N_9468);
or UO_716 (O_716,N_9475,N_9557);
nor UO_717 (O_717,N_9232,N_9181);
nor UO_718 (O_718,N_9008,N_9626);
nor UO_719 (O_719,N_9557,N_9712);
nor UO_720 (O_720,N_9338,N_9757);
nor UO_721 (O_721,N_9525,N_9741);
or UO_722 (O_722,N_9498,N_9532);
or UO_723 (O_723,N_9177,N_9189);
nor UO_724 (O_724,N_9138,N_9330);
or UO_725 (O_725,N_9473,N_9852);
nor UO_726 (O_726,N_9798,N_9038);
nand UO_727 (O_727,N_9269,N_9654);
or UO_728 (O_728,N_9128,N_9370);
and UO_729 (O_729,N_9297,N_9237);
nand UO_730 (O_730,N_9523,N_9768);
nand UO_731 (O_731,N_9264,N_9803);
nor UO_732 (O_732,N_9981,N_9139);
and UO_733 (O_733,N_9714,N_9787);
nand UO_734 (O_734,N_9945,N_9019);
nor UO_735 (O_735,N_9392,N_9161);
nand UO_736 (O_736,N_9119,N_9567);
nand UO_737 (O_737,N_9345,N_9349);
or UO_738 (O_738,N_9752,N_9824);
nor UO_739 (O_739,N_9298,N_9781);
or UO_740 (O_740,N_9449,N_9349);
and UO_741 (O_741,N_9618,N_9214);
and UO_742 (O_742,N_9415,N_9775);
nor UO_743 (O_743,N_9390,N_9051);
or UO_744 (O_744,N_9690,N_9523);
nor UO_745 (O_745,N_9913,N_9467);
nand UO_746 (O_746,N_9175,N_9593);
and UO_747 (O_747,N_9822,N_9106);
and UO_748 (O_748,N_9228,N_9858);
nand UO_749 (O_749,N_9435,N_9605);
or UO_750 (O_750,N_9432,N_9344);
nand UO_751 (O_751,N_9755,N_9868);
and UO_752 (O_752,N_9995,N_9257);
or UO_753 (O_753,N_9843,N_9294);
nand UO_754 (O_754,N_9500,N_9423);
or UO_755 (O_755,N_9474,N_9188);
or UO_756 (O_756,N_9550,N_9819);
nor UO_757 (O_757,N_9277,N_9490);
and UO_758 (O_758,N_9004,N_9997);
nand UO_759 (O_759,N_9557,N_9993);
or UO_760 (O_760,N_9439,N_9295);
or UO_761 (O_761,N_9358,N_9171);
nor UO_762 (O_762,N_9384,N_9589);
or UO_763 (O_763,N_9548,N_9919);
nand UO_764 (O_764,N_9716,N_9911);
or UO_765 (O_765,N_9062,N_9614);
nor UO_766 (O_766,N_9467,N_9851);
nand UO_767 (O_767,N_9849,N_9458);
and UO_768 (O_768,N_9838,N_9001);
and UO_769 (O_769,N_9086,N_9902);
nand UO_770 (O_770,N_9092,N_9836);
nor UO_771 (O_771,N_9402,N_9282);
and UO_772 (O_772,N_9431,N_9004);
nand UO_773 (O_773,N_9369,N_9224);
nand UO_774 (O_774,N_9970,N_9568);
nor UO_775 (O_775,N_9849,N_9692);
or UO_776 (O_776,N_9046,N_9747);
nor UO_777 (O_777,N_9936,N_9569);
nand UO_778 (O_778,N_9521,N_9542);
nand UO_779 (O_779,N_9535,N_9063);
or UO_780 (O_780,N_9263,N_9170);
nand UO_781 (O_781,N_9733,N_9596);
and UO_782 (O_782,N_9139,N_9217);
or UO_783 (O_783,N_9463,N_9798);
and UO_784 (O_784,N_9249,N_9186);
or UO_785 (O_785,N_9433,N_9726);
nor UO_786 (O_786,N_9746,N_9732);
and UO_787 (O_787,N_9643,N_9910);
nor UO_788 (O_788,N_9363,N_9423);
or UO_789 (O_789,N_9796,N_9175);
nor UO_790 (O_790,N_9013,N_9142);
and UO_791 (O_791,N_9224,N_9454);
or UO_792 (O_792,N_9458,N_9067);
or UO_793 (O_793,N_9241,N_9791);
or UO_794 (O_794,N_9163,N_9390);
or UO_795 (O_795,N_9992,N_9385);
and UO_796 (O_796,N_9686,N_9057);
and UO_797 (O_797,N_9818,N_9749);
or UO_798 (O_798,N_9586,N_9279);
and UO_799 (O_799,N_9996,N_9980);
nor UO_800 (O_800,N_9736,N_9613);
or UO_801 (O_801,N_9832,N_9463);
or UO_802 (O_802,N_9352,N_9548);
and UO_803 (O_803,N_9699,N_9338);
nor UO_804 (O_804,N_9115,N_9604);
and UO_805 (O_805,N_9791,N_9783);
and UO_806 (O_806,N_9793,N_9243);
nor UO_807 (O_807,N_9946,N_9113);
nor UO_808 (O_808,N_9328,N_9379);
nand UO_809 (O_809,N_9457,N_9363);
nor UO_810 (O_810,N_9952,N_9660);
or UO_811 (O_811,N_9516,N_9372);
nor UO_812 (O_812,N_9320,N_9242);
nor UO_813 (O_813,N_9466,N_9655);
or UO_814 (O_814,N_9372,N_9924);
or UO_815 (O_815,N_9759,N_9963);
and UO_816 (O_816,N_9204,N_9524);
nor UO_817 (O_817,N_9785,N_9841);
nand UO_818 (O_818,N_9610,N_9092);
nand UO_819 (O_819,N_9094,N_9251);
nand UO_820 (O_820,N_9198,N_9024);
nand UO_821 (O_821,N_9981,N_9465);
nor UO_822 (O_822,N_9929,N_9402);
and UO_823 (O_823,N_9386,N_9687);
nand UO_824 (O_824,N_9530,N_9445);
or UO_825 (O_825,N_9031,N_9921);
nand UO_826 (O_826,N_9446,N_9254);
nand UO_827 (O_827,N_9882,N_9824);
nand UO_828 (O_828,N_9514,N_9234);
and UO_829 (O_829,N_9913,N_9745);
or UO_830 (O_830,N_9168,N_9120);
or UO_831 (O_831,N_9567,N_9520);
nor UO_832 (O_832,N_9489,N_9058);
and UO_833 (O_833,N_9262,N_9623);
and UO_834 (O_834,N_9223,N_9209);
nor UO_835 (O_835,N_9528,N_9611);
nor UO_836 (O_836,N_9974,N_9628);
nor UO_837 (O_837,N_9248,N_9165);
and UO_838 (O_838,N_9597,N_9759);
nand UO_839 (O_839,N_9800,N_9638);
xor UO_840 (O_840,N_9360,N_9664);
nor UO_841 (O_841,N_9977,N_9342);
and UO_842 (O_842,N_9749,N_9948);
and UO_843 (O_843,N_9596,N_9258);
or UO_844 (O_844,N_9756,N_9331);
nand UO_845 (O_845,N_9154,N_9755);
and UO_846 (O_846,N_9653,N_9780);
nor UO_847 (O_847,N_9026,N_9924);
and UO_848 (O_848,N_9107,N_9582);
or UO_849 (O_849,N_9237,N_9110);
xor UO_850 (O_850,N_9177,N_9519);
or UO_851 (O_851,N_9034,N_9609);
nand UO_852 (O_852,N_9513,N_9367);
nand UO_853 (O_853,N_9075,N_9842);
nand UO_854 (O_854,N_9946,N_9047);
nor UO_855 (O_855,N_9880,N_9652);
or UO_856 (O_856,N_9159,N_9969);
nand UO_857 (O_857,N_9313,N_9455);
nor UO_858 (O_858,N_9704,N_9618);
or UO_859 (O_859,N_9068,N_9584);
or UO_860 (O_860,N_9395,N_9987);
or UO_861 (O_861,N_9814,N_9647);
nand UO_862 (O_862,N_9276,N_9834);
nand UO_863 (O_863,N_9269,N_9221);
nand UO_864 (O_864,N_9675,N_9449);
nand UO_865 (O_865,N_9951,N_9834);
and UO_866 (O_866,N_9142,N_9546);
nand UO_867 (O_867,N_9707,N_9109);
nand UO_868 (O_868,N_9168,N_9298);
nand UO_869 (O_869,N_9348,N_9806);
and UO_870 (O_870,N_9160,N_9500);
nand UO_871 (O_871,N_9611,N_9758);
nand UO_872 (O_872,N_9992,N_9151);
or UO_873 (O_873,N_9407,N_9151);
nand UO_874 (O_874,N_9338,N_9558);
or UO_875 (O_875,N_9653,N_9183);
nor UO_876 (O_876,N_9040,N_9245);
nand UO_877 (O_877,N_9082,N_9734);
nor UO_878 (O_878,N_9780,N_9399);
or UO_879 (O_879,N_9714,N_9294);
and UO_880 (O_880,N_9196,N_9561);
nor UO_881 (O_881,N_9762,N_9361);
or UO_882 (O_882,N_9284,N_9698);
nor UO_883 (O_883,N_9475,N_9145);
nor UO_884 (O_884,N_9990,N_9109);
nor UO_885 (O_885,N_9131,N_9798);
or UO_886 (O_886,N_9951,N_9084);
and UO_887 (O_887,N_9945,N_9465);
and UO_888 (O_888,N_9348,N_9249);
and UO_889 (O_889,N_9385,N_9504);
nor UO_890 (O_890,N_9952,N_9420);
or UO_891 (O_891,N_9635,N_9442);
nor UO_892 (O_892,N_9950,N_9931);
or UO_893 (O_893,N_9458,N_9931);
nor UO_894 (O_894,N_9130,N_9759);
or UO_895 (O_895,N_9248,N_9192);
nor UO_896 (O_896,N_9116,N_9308);
nor UO_897 (O_897,N_9656,N_9564);
and UO_898 (O_898,N_9705,N_9311);
and UO_899 (O_899,N_9566,N_9240);
and UO_900 (O_900,N_9507,N_9139);
or UO_901 (O_901,N_9129,N_9083);
nor UO_902 (O_902,N_9877,N_9944);
nand UO_903 (O_903,N_9335,N_9274);
nand UO_904 (O_904,N_9044,N_9581);
nor UO_905 (O_905,N_9073,N_9231);
or UO_906 (O_906,N_9076,N_9229);
and UO_907 (O_907,N_9622,N_9712);
or UO_908 (O_908,N_9184,N_9143);
nand UO_909 (O_909,N_9348,N_9835);
or UO_910 (O_910,N_9579,N_9682);
or UO_911 (O_911,N_9080,N_9090);
and UO_912 (O_912,N_9024,N_9936);
or UO_913 (O_913,N_9497,N_9903);
nand UO_914 (O_914,N_9669,N_9394);
nor UO_915 (O_915,N_9432,N_9410);
nand UO_916 (O_916,N_9694,N_9712);
nor UO_917 (O_917,N_9823,N_9689);
nand UO_918 (O_918,N_9083,N_9268);
nand UO_919 (O_919,N_9052,N_9154);
and UO_920 (O_920,N_9950,N_9712);
or UO_921 (O_921,N_9121,N_9007);
or UO_922 (O_922,N_9549,N_9980);
and UO_923 (O_923,N_9937,N_9895);
and UO_924 (O_924,N_9820,N_9071);
nor UO_925 (O_925,N_9057,N_9780);
nand UO_926 (O_926,N_9974,N_9990);
or UO_927 (O_927,N_9041,N_9621);
nand UO_928 (O_928,N_9642,N_9680);
and UO_929 (O_929,N_9100,N_9006);
nor UO_930 (O_930,N_9752,N_9394);
or UO_931 (O_931,N_9396,N_9027);
nand UO_932 (O_932,N_9316,N_9015);
nor UO_933 (O_933,N_9327,N_9459);
nand UO_934 (O_934,N_9323,N_9840);
nor UO_935 (O_935,N_9282,N_9722);
nand UO_936 (O_936,N_9909,N_9921);
and UO_937 (O_937,N_9254,N_9851);
and UO_938 (O_938,N_9613,N_9454);
nor UO_939 (O_939,N_9971,N_9525);
or UO_940 (O_940,N_9315,N_9684);
nand UO_941 (O_941,N_9153,N_9838);
nand UO_942 (O_942,N_9387,N_9127);
nand UO_943 (O_943,N_9041,N_9783);
nand UO_944 (O_944,N_9886,N_9229);
nand UO_945 (O_945,N_9807,N_9516);
nand UO_946 (O_946,N_9881,N_9884);
or UO_947 (O_947,N_9803,N_9021);
nor UO_948 (O_948,N_9762,N_9786);
and UO_949 (O_949,N_9728,N_9338);
and UO_950 (O_950,N_9796,N_9228);
nand UO_951 (O_951,N_9812,N_9022);
nand UO_952 (O_952,N_9640,N_9730);
and UO_953 (O_953,N_9402,N_9592);
and UO_954 (O_954,N_9060,N_9744);
and UO_955 (O_955,N_9228,N_9209);
nand UO_956 (O_956,N_9560,N_9832);
and UO_957 (O_957,N_9680,N_9957);
nor UO_958 (O_958,N_9022,N_9861);
nand UO_959 (O_959,N_9980,N_9072);
and UO_960 (O_960,N_9342,N_9401);
xor UO_961 (O_961,N_9961,N_9115);
and UO_962 (O_962,N_9416,N_9087);
or UO_963 (O_963,N_9868,N_9332);
and UO_964 (O_964,N_9132,N_9404);
and UO_965 (O_965,N_9080,N_9012);
or UO_966 (O_966,N_9947,N_9897);
nand UO_967 (O_967,N_9222,N_9281);
nand UO_968 (O_968,N_9326,N_9354);
nor UO_969 (O_969,N_9016,N_9459);
and UO_970 (O_970,N_9675,N_9257);
and UO_971 (O_971,N_9943,N_9829);
xnor UO_972 (O_972,N_9103,N_9860);
nand UO_973 (O_973,N_9110,N_9798);
nand UO_974 (O_974,N_9906,N_9708);
or UO_975 (O_975,N_9195,N_9802);
nand UO_976 (O_976,N_9632,N_9774);
and UO_977 (O_977,N_9121,N_9292);
nand UO_978 (O_978,N_9269,N_9494);
or UO_979 (O_979,N_9006,N_9212);
and UO_980 (O_980,N_9956,N_9224);
nand UO_981 (O_981,N_9669,N_9759);
nand UO_982 (O_982,N_9619,N_9792);
or UO_983 (O_983,N_9986,N_9453);
nand UO_984 (O_984,N_9182,N_9374);
nand UO_985 (O_985,N_9099,N_9565);
and UO_986 (O_986,N_9718,N_9055);
nand UO_987 (O_987,N_9737,N_9651);
nand UO_988 (O_988,N_9383,N_9465);
and UO_989 (O_989,N_9445,N_9816);
nor UO_990 (O_990,N_9743,N_9913);
nand UO_991 (O_991,N_9733,N_9043);
nand UO_992 (O_992,N_9262,N_9566);
and UO_993 (O_993,N_9096,N_9881);
nor UO_994 (O_994,N_9886,N_9185);
or UO_995 (O_995,N_9583,N_9384);
nor UO_996 (O_996,N_9883,N_9588);
and UO_997 (O_997,N_9505,N_9628);
xor UO_998 (O_998,N_9808,N_9992);
or UO_999 (O_999,N_9619,N_9799);
nor UO_1000 (O_1000,N_9023,N_9420);
xor UO_1001 (O_1001,N_9477,N_9123);
or UO_1002 (O_1002,N_9495,N_9509);
and UO_1003 (O_1003,N_9145,N_9363);
and UO_1004 (O_1004,N_9617,N_9936);
or UO_1005 (O_1005,N_9697,N_9074);
nor UO_1006 (O_1006,N_9686,N_9822);
or UO_1007 (O_1007,N_9894,N_9799);
nand UO_1008 (O_1008,N_9616,N_9091);
and UO_1009 (O_1009,N_9317,N_9753);
nand UO_1010 (O_1010,N_9806,N_9872);
nand UO_1011 (O_1011,N_9371,N_9115);
and UO_1012 (O_1012,N_9492,N_9245);
or UO_1013 (O_1013,N_9860,N_9371);
nor UO_1014 (O_1014,N_9044,N_9489);
and UO_1015 (O_1015,N_9715,N_9838);
xor UO_1016 (O_1016,N_9281,N_9963);
or UO_1017 (O_1017,N_9136,N_9059);
or UO_1018 (O_1018,N_9587,N_9358);
nand UO_1019 (O_1019,N_9899,N_9803);
or UO_1020 (O_1020,N_9057,N_9680);
and UO_1021 (O_1021,N_9157,N_9695);
xor UO_1022 (O_1022,N_9686,N_9096);
or UO_1023 (O_1023,N_9305,N_9810);
and UO_1024 (O_1024,N_9450,N_9484);
nor UO_1025 (O_1025,N_9424,N_9391);
nor UO_1026 (O_1026,N_9757,N_9207);
xnor UO_1027 (O_1027,N_9270,N_9045);
nand UO_1028 (O_1028,N_9409,N_9334);
and UO_1029 (O_1029,N_9878,N_9836);
and UO_1030 (O_1030,N_9590,N_9071);
or UO_1031 (O_1031,N_9059,N_9030);
nand UO_1032 (O_1032,N_9908,N_9108);
and UO_1033 (O_1033,N_9626,N_9453);
nand UO_1034 (O_1034,N_9751,N_9715);
nand UO_1035 (O_1035,N_9454,N_9896);
nor UO_1036 (O_1036,N_9736,N_9469);
and UO_1037 (O_1037,N_9762,N_9415);
or UO_1038 (O_1038,N_9024,N_9151);
nand UO_1039 (O_1039,N_9823,N_9342);
and UO_1040 (O_1040,N_9890,N_9663);
nor UO_1041 (O_1041,N_9084,N_9234);
nor UO_1042 (O_1042,N_9979,N_9088);
and UO_1043 (O_1043,N_9583,N_9788);
and UO_1044 (O_1044,N_9596,N_9530);
and UO_1045 (O_1045,N_9044,N_9689);
nand UO_1046 (O_1046,N_9350,N_9537);
nand UO_1047 (O_1047,N_9212,N_9974);
nand UO_1048 (O_1048,N_9841,N_9199);
or UO_1049 (O_1049,N_9054,N_9661);
or UO_1050 (O_1050,N_9356,N_9415);
or UO_1051 (O_1051,N_9222,N_9011);
nor UO_1052 (O_1052,N_9052,N_9541);
and UO_1053 (O_1053,N_9245,N_9917);
nand UO_1054 (O_1054,N_9053,N_9054);
nor UO_1055 (O_1055,N_9183,N_9036);
nand UO_1056 (O_1056,N_9677,N_9590);
xnor UO_1057 (O_1057,N_9094,N_9567);
nand UO_1058 (O_1058,N_9895,N_9225);
and UO_1059 (O_1059,N_9681,N_9077);
and UO_1060 (O_1060,N_9562,N_9964);
nor UO_1061 (O_1061,N_9801,N_9715);
nand UO_1062 (O_1062,N_9195,N_9764);
nor UO_1063 (O_1063,N_9400,N_9733);
nor UO_1064 (O_1064,N_9510,N_9003);
or UO_1065 (O_1065,N_9435,N_9385);
and UO_1066 (O_1066,N_9743,N_9863);
nand UO_1067 (O_1067,N_9605,N_9945);
and UO_1068 (O_1068,N_9577,N_9450);
nor UO_1069 (O_1069,N_9961,N_9397);
and UO_1070 (O_1070,N_9701,N_9119);
and UO_1071 (O_1071,N_9666,N_9399);
and UO_1072 (O_1072,N_9880,N_9955);
nor UO_1073 (O_1073,N_9045,N_9150);
or UO_1074 (O_1074,N_9168,N_9335);
nand UO_1075 (O_1075,N_9014,N_9299);
and UO_1076 (O_1076,N_9924,N_9802);
or UO_1077 (O_1077,N_9320,N_9270);
nor UO_1078 (O_1078,N_9042,N_9259);
nor UO_1079 (O_1079,N_9201,N_9611);
nand UO_1080 (O_1080,N_9404,N_9309);
nand UO_1081 (O_1081,N_9467,N_9217);
and UO_1082 (O_1082,N_9176,N_9588);
nand UO_1083 (O_1083,N_9581,N_9612);
xnor UO_1084 (O_1084,N_9265,N_9724);
or UO_1085 (O_1085,N_9764,N_9749);
or UO_1086 (O_1086,N_9689,N_9657);
nand UO_1087 (O_1087,N_9413,N_9987);
and UO_1088 (O_1088,N_9912,N_9009);
or UO_1089 (O_1089,N_9254,N_9463);
or UO_1090 (O_1090,N_9311,N_9376);
xnor UO_1091 (O_1091,N_9998,N_9320);
nor UO_1092 (O_1092,N_9111,N_9745);
nand UO_1093 (O_1093,N_9042,N_9045);
or UO_1094 (O_1094,N_9121,N_9900);
nand UO_1095 (O_1095,N_9699,N_9672);
nor UO_1096 (O_1096,N_9468,N_9369);
or UO_1097 (O_1097,N_9507,N_9492);
nand UO_1098 (O_1098,N_9362,N_9506);
and UO_1099 (O_1099,N_9970,N_9723);
or UO_1100 (O_1100,N_9932,N_9055);
or UO_1101 (O_1101,N_9910,N_9476);
and UO_1102 (O_1102,N_9311,N_9032);
or UO_1103 (O_1103,N_9993,N_9314);
nand UO_1104 (O_1104,N_9856,N_9941);
nor UO_1105 (O_1105,N_9925,N_9363);
nand UO_1106 (O_1106,N_9848,N_9486);
nand UO_1107 (O_1107,N_9587,N_9796);
nor UO_1108 (O_1108,N_9219,N_9460);
nor UO_1109 (O_1109,N_9457,N_9178);
and UO_1110 (O_1110,N_9595,N_9599);
or UO_1111 (O_1111,N_9017,N_9944);
nand UO_1112 (O_1112,N_9725,N_9403);
and UO_1113 (O_1113,N_9117,N_9510);
and UO_1114 (O_1114,N_9215,N_9887);
nand UO_1115 (O_1115,N_9289,N_9144);
nand UO_1116 (O_1116,N_9952,N_9000);
nor UO_1117 (O_1117,N_9294,N_9104);
nor UO_1118 (O_1118,N_9874,N_9799);
and UO_1119 (O_1119,N_9650,N_9074);
xor UO_1120 (O_1120,N_9618,N_9671);
or UO_1121 (O_1121,N_9087,N_9852);
nor UO_1122 (O_1122,N_9558,N_9874);
or UO_1123 (O_1123,N_9292,N_9396);
nor UO_1124 (O_1124,N_9466,N_9481);
and UO_1125 (O_1125,N_9313,N_9351);
nor UO_1126 (O_1126,N_9660,N_9909);
or UO_1127 (O_1127,N_9960,N_9116);
nand UO_1128 (O_1128,N_9746,N_9418);
or UO_1129 (O_1129,N_9506,N_9557);
xnor UO_1130 (O_1130,N_9677,N_9530);
xor UO_1131 (O_1131,N_9534,N_9879);
and UO_1132 (O_1132,N_9323,N_9226);
nand UO_1133 (O_1133,N_9313,N_9922);
nor UO_1134 (O_1134,N_9743,N_9716);
and UO_1135 (O_1135,N_9319,N_9855);
or UO_1136 (O_1136,N_9191,N_9619);
and UO_1137 (O_1137,N_9328,N_9764);
nor UO_1138 (O_1138,N_9940,N_9331);
and UO_1139 (O_1139,N_9595,N_9322);
nand UO_1140 (O_1140,N_9695,N_9249);
or UO_1141 (O_1141,N_9306,N_9153);
nor UO_1142 (O_1142,N_9259,N_9846);
or UO_1143 (O_1143,N_9944,N_9965);
nor UO_1144 (O_1144,N_9048,N_9514);
nand UO_1145 (O_1145,N_9483,N_9870);
or UO_1146 (O_1146,N_9675,N_9493);
and UO_1147 (O_1147,N_9791,N_9362);
and UO_1148 (O_1148,N_9762,N_9320);
nand UO_1149 (O_1149,N_9107,N_9515);
or UO_1150 (O_1150,N_9170,N_9117);
and UO_1151 (O_1151,N_9878,N_9780);
nand UO_1152 (O_1152,N_9996,N_9835);
or UO_1153 (O_1153,N_9108,N_9632);
and UO_1154 (O_1154,N_9797,N_9910);
or UO_1155 (O_1155,N_9144,N_9315);
nor UO_1156 (O_1156,N_9316,N_9813);
nand UO_1157 (O_1157,N_9429,N_9215);
xnor UO_1158 (O_1158,N_9782,N_9697);
nand UO_1159 (O_1159,N_9621,N_9587);
or UO_1160 (O_1160,N_9237,N_9147);
nor UO_1161 (O_1161,N_9552,N_9066);
or UO_1162 (O_1162,N_9379,N_9389);
or UO_1163 (O_1163,N_9304,N_9245);
nor UO_1164 (O_1164,N_9195,N_9547);
xnor UO_1165 (O_1165,N_9298,N_9616);
nand UO_1166 (O_1166,N_9501,N_9299);
nand UO_1167 (O_1167,N_9340,N_9097);
nand UO_1168 (O_1168,N_9428,N_9644);
nand UO_1169 (O_1169,N_9920,N_9829);
nand UO_1170 (O_1170,N_9344,N_9623);
or UO_1171 (O_1171,N_9877,N_9972);
or UO_1172 (O_1172,N_9358,N_9300);
or UO_1173 (O_1173,N_9621,N_9167);
nand UO_1174 (O_1174,N_9428,N_9939);
nor UO_1175 (O_1175,N_9043,N_9431);
and UO_1176 (O_1176,N_9278,N_9286);
or UO_1177 (O_1177,N_9988,N_9098);
nand UO_1178 (O_1178,N_9430,N_9580);
and UO_1179 (O_1179,N_9700,N_9209);
or UO_1180 (O_1180,N_9405,N_9629);
or UO_1181 (O_1181,N_9615,N_9795);
nor UO_1182 (O_1182,N_9607,N_9005);
and UO_1183 (O_1183,N_9553,N_9334);
nor UO_1184 (O_1184,N_9635,N_9378);
nor UO_1185 (O_1185,N_9114,N_9991);
nor UO_1186 (O_1186,N_9759,N_9375);
nor UO_1187 (O_1187,N_9402,N_9191);
nor UO_1188 (O_1188,N_9764,N_9048);
nor UO_1189 (O_1189,N_9740,N_9609);
or UO_1190 (O_1190,N_9140,N_9825);
and UO_1191 (O_1191,N_9817,N_9860);
nand UO_1192 (O_1192,N_9451,N_9196);
xnor UO_1193 (O_1193,N_9951,N_9467);
nand UO_1194 (O_1194,N_9963,N_9019);
nor UO_1195 (O_1195,N_9474,N_9923);
nand UO_1196 (O_1196,N_9230,N_9890);
and UO_1197 (O_1197,N_9026,N_9606);
xor UO_1198 (O_1198,N_9480,N_9185);
nand UO_1199 (O_1199,N_9777,N_9774);
nand UO_1200 (O_1200,N_9471,N_9394);
nor UO_1201 (O_1201,N_9618,N_9799);
or UO_1202 (O_1202,N_9116,N_9681);
nor UO_1203 (O_1203,N_9275,N_9978);
and UO_1204 (O_1204,N_9323,N_9057);
xnor UO_1205 (O_1205,N_9082,N_9172);
and UO_1206 (O_1206,N_9368,N_9399);
nand UO_1207 (O_1207,N_9485,N_9433);
or UO_1208 (O_1208,N_9354,N_9480);
nand UO_1209 (O_1209,N_9997,N_9514);
or UO_1210 (O_1210,N_9665,N_9047);
nand UO_1211 (O_1211,N_9958,N_9022);
nand UO_1212 (O_1212,N_9157,N_9607);
nor UO_1213 (O_1213,N_9600,N_9638);
and UO_1214 (O_1214,N_9329,N_9142);
or UO_1215 (O_1215,N_9227,N_9701);
or UO_1216 (O_1216,N_9411,N_9965);
xor UO_1217 (O_1217,N_9070,N_9827);
nand UO_1218 (O_1218,N_9032,N_9422);
nand UO_1219 (O_1219,N_9836,N_9897);
or UO_1220 (O_1220,N_9378,N_9045);
nand UO_1221 (O_1221,N_9574,N_9013);
nand UO_1222 (O_1222,N_9481,N_9775);
and UO_1223 (O_1223,N_9217,N_9617);
and UO_1224 (O_1224,N_9707,N_9907);
nor UO_1225 (O_1225,N_9384,N_9868);
and UO_1226 (O_1226,N_9614,N_9295);
nand UO_1227 (O_1227,N_9444,N_9190);
and UO_1228 (O_1228,N_9637,N_9491);
and UO_1229 (O_1229,N_9181,N_9580);
and UO_1230 (O_1230,N_9024,N_9666);
nor UO_1231 (O_1231,N_9521,N_9074);
or UO_1232 (O_1232,N_9289,N_9028);
nor UO_1233 (O_1233,N_9939,N_9626);
and UO_1234 (O_1234,N_9853,N_9363);
nor UO_1235 (O_1235,N_9475,N_9144);
or UO_1236 (O_1236,N_9582,N_9489);
nor UO_1237 (O_1237,N_9194,N_9009);
nand UO_1238 (O_1238,N_9869,N_9843);
and UO_1239 (O_1239,N_9613,N_9587);
or UO_1240 (O_1240,N_9693,N_9183);
xor UO_1241 (O_1241,N_9686,N_9257);
nand UO_1242 (O_1242,N_9544,N_9192);
nand UO_1243 (O_1243,N_9648,N_9303);
and UO_1244 (O_1244,N_9767,N_9533);
or UO_1245 (O_1245,N_9922,N_9630);
or UO_1246 (O_1246,N_9656,N_9544);
and UO_1247 (O_1247,N_9203,N_9022);
nor UO_1248 (O_1248,N_9779,N_9654);
nor UO_1249 (O_1249,N_9079,N_9781);
nor UO_1250 (O_1250,N_9632,N_9913);
or UO_1251 (O_1251,N_9145,N_9968);
nor UO_1252 (O_1252,N_9727,N_9507);
nor UO_1253 (O_1253,N_9784,N_9476);
nor UO_1254 (O_1254,N_9767,N_9764);
nand UO_1255 (O_1255,N_9526,N_9337);
nand UO_1256 (O_1256,N_9238,N_9907);
or UO_1257 (O_1257,N_9106,N_9363);
nand UO_1258 (O_1258,N_9783,N_9327);
nor UO_1259 (O_1259,N_9257,N_9873);
nand UO_1260 (O_1260,N_9205,N_9599);
nor UO_1261 (O_1261,N_9115,N_9023);
or UO_1262 (O_1262,N_9965,N_9185);
and UO_1263 (O_1263,N_9877,N_9992);
xnor UO_1264 (O_1264,N_9951,N_9011);
nor UO_1265 (O_1265,N_9454,N_9368);
or UO_1266 (O_1266,N_9955,N_9176);
nor UO_1267 (O_1267,N_9607,N_9911);
nor UO_1268 (O_1268,N_9606,N_9559);
and UO_1269 (O_1269,N_9700,N_9160);
and UO_1270 (O_1270,N_9046,N_9660);
nand UO_1271 (O_1271,N_9229,N_9693);
nor UO_1272 (O_1272,N_9202,N_9466);
nor UO_1273 (O_1273,N_9747,N_9512);
or UO_1274 (O_1274,N_9735,N_9113);
nand UO_1275 (O_1275,N_9149,N_9359);
nand UO_1276 (O_1276,N_9344,N_9466);
xnor UO_1277 (O_1277,N_9382,N_9027);
nor UO_1278 (O_1278,N_9783,N_9966);
nand UO_1279 (O_1279,N_9031,N_9296);
or UO_1280 (O_1280,N_9608,N_9343);
and UO_1281 (O_1281,N_9378,N_9315);
and UO_1282 (O_1282,N_9712,N_9812);
nand UO_1283 (O_1283,N_9624,N_9303);
or UO_1284 (O_1284,N_9383,N_9842);
xnor UO_1285 (O_1285,N_9377,N_9278);
and UO_1286 (O_1286,N_9401,N_9757);
nand UO_1287 (O_1287,N_9074,N_9818);
and UO_1288 (O_1288,N_9553,N_9240);
nand UO_1289 (O_1289,N_9569,N_9973);
nand UO_1290 (O_1290,N_9099,N_9411);
nor UO_1291 (O_1291,N_9793,N_9465);
nor UO_1292 (O_1292,N_9418,N_9301);
nand UO_1293 (O_1293,N_9192,N_9624);
nor UO_1294 (O_1294,N_9061,N_9034);
and UO_1295 (O_1295,N_9890,N_9281);
or UO_1296 (O_1296,N_9731,N_9779);
nand UO_1297 (O_1297,N_9589,N_9591);
nand UO_1298 (O_1298,N_9667,N_9127);
or UO_1299 (O_1299,N_9931,N_9047);
and UO_1300 (O_1300,N_9776,N_9836);
or UO_1301 (O_1301,N_9504,N_9307);
and UO_1302 (O_1302,N_9083,N_9590);
xor UO_1303 (O_1303,N_9814,N_9784);
nand UO_1304 (O_1304,N_9337,N_9611);
or UO_1305 (O_1305,N_9434,N_9609);
or UO_1306 (O_1306,N_9198,N_9613);
and UO_1307 (O_1307,N_9837,N_9071);
or UO_1308 (O_1308,N_9840,N_9187);
nand UO_1309 (O_1309,N_9002,N_9451);
nor UO_1310 (O_1310,N_9854,N_9715);
nand UO_1311 (O_1311,N_9989,N_9437);
or UO_1312 (O_1312,N_9831,N_9007);
or UO_1313 (O_1313,N_9202,N_9421);
or UO_1314 (O_1314,N_9275,N_9133);
and UO_1315 (O_1315,N_9411,N_9321);
nor UO_1316 (O_1316,N_9522,N_9592);
and UO_1317 (O_1317,N_9763,N_9590);
nor UO_1318 (O_1318,N_9689,N_9231);
nand UO_1319 (O_1319,N_9551,N_9474);
nor UO_1320 (O_1320,N_9789,N_9363);
or UO_1321 (O_1321,N_9827,N_9351);
and UO_1322 (O_1322,N_9265,N_9488);
or UO_1323 (O_1323,N_9134,N_9478);
or UO_1324 (O_1324,N_9770,N_9127);
and UO_1325 (O_1325,N_9189,N_9080);
or UO_1326 (O_1326,N_9798,N_9595);
nor UO_1327 (O_1327,N_9319,N_9623);
or UO_1328 (O_1328,N_9614,N_9990);
nor UO_1329 (O_1329,N_9368,N_9929);
or UO_1330 (O_1330,N_9995,N_9823);
and UO_1331 (O_1331,N_9896,N_9644);
nor UO_1332 (O_1332,N_9967,N_9582);
and UO_1333 (O_1333,N_9820,N_9703);
nor UO_1334 (O_1334,N_9401,N_9795);
nor UO_1335 (O_1335,N_9620,N_9199);
nand UO_1336 (O_1336,N_9205,N_9149);
or UO_1337 (O_1337,N_9249,N_9040);
and UO_1338 (O_1338,N_9704,N_9783);
nor UO_1339 (O_1339,N_9785,N_9973);
nor UO_1340 (O_1340,N_9648,N_9872);
or UO_1341 (O_1341,N_9275,N_9273);
nand UO_1342 (O_1342,N_9245,N_9335);
nor UO_1343 (O_1343,N_9945,N_9836);
or UO_1344 (O_1344,N_9605,N_9385);
and UO_1345 (O_1345,N_9536,N_9778);
nor UO_1346 (O_1346,N_9120,N_9907);
or UO_1347 (O_1347,N_9024,N_9197);
nor UO_1348 (O_1348,N_9033,N_9659);
nand UO_1349 (O_1349,N_9052,N_9387);
nand UO_1350 (O_1350,N_9919,N_9719);
nor UO_1351 (O_1351,N_9702,N_9810);
and UO_1352 (O_1352,N_9641,N_9825);
or UO_1353 (O_1353,N_9844,N_9696);
or UO_1354 (O_1354,N_9037,N_9657);
nor UO_1355 (O_1355,N_9074,N_9341);
nand UO_1356 (O_1356,N_9331,N_9038);
or UO_1357 (O_1357,N_9646,N_9084);
nor UO_1358 (O_1358,N_9809,N_9717);
nand UO_1359 (O_1359,N_9525,N_9881);
nor UO_1360 (O_1360,N_9962,N_9487);
nand UO_1361 (O_1361,N_9569,N_9926);
or UO_1362 (O_1362,N_9805,N_9492);
or UO_1363 (O_1363,N_9967,N_9850);
nor UO_1364 (O_1364,N_9884,N_9855);
nand UO_1365 (O_1365,N_9409,N_9253);
or UO_1366 (O_1366,N_9132,N_9546);
and UO_1367 (O_1367,N_9716,N_9625);
or UO_1368 (O_1368,N_9636,N_9418);
nand UO_1369 (O_1369,N_9760,N_9607);
and UO_1370 (O_1370,N_9289,N_9395);
nor UO_1371 (O_1371,N_9266,N_9423);
nand UO_1372 (O_1372,N_9727,N_9814);
nand UO_1373 (O_1373,N_9787,N_9404);
and UO_1374 (O_1374,N_9724,N_9661);
or UO_1375 (O_1375,N_9908,N_9690);
nand UO_1376 (O_1376,N_9381,N_9420);
or UO_1377 (O_1377,N_9113,N_9124);
and UO_1378 (O_1378,N_9953,N_9496);
or UO_1379 (O_1379,N_9174,N_9717);
and UO_1380 (O_1380,N_9689,N_9494);
nand UO_1381 (O_1381,N_9865,N_9594);
or UO_1382 (O_1382,N_9643,N_9471);
nor UO_1383 (O_1383,N_9548,N_9522);
nand UO_1384 (O_1384,N_9448,N_9165);
and UO_1385 (O_1385,N_9539,N_9135);
and UO_1386 (O_1386,N_9215,N_9441);
nor UO_1387 (O_1387,N_9122,N_9934);
nor UO_1388 (O_1388,N_9836,N_9144);
and UO_1389 (O_1389,N_9224,N_9431);
and UO_1390 (O_1390,N_9807,N_9225);
nand UO_1391 (O_1391,N_9694,N_9027);
nand UO_1392 (O_1392,N_9809,N_9423);
and UO_1393 (O_1393,N_9588,N_9148);
and UO_1394 (O_1394,N_9773,N_9036);
nor UO_1395 (O_1395,N_9884,N_9710);
nand UO_1396 (O_1396,N_9033,N_9622);
or UO_1397 (O_1397,N_9951,N_9662);
and UO_1398 (O_1398,N_9888,N_9277);
or UO_1399 (O_1399,N_9627,N_9902);
nand UO_1400 (O_1400,N_9096,N_9703);
nand UO_1401 (O_1401,N_9011,N_9803);
xnor UO_1402 (O_1402,N_9464,N_9246);
and UO_1403 (O_1403,N_9617,N_9790);
or UO_1404 (O_1404,N_9581,N_9097);
or UO_1405 (O_1405,N_9553,N_9137);
nor UO_1406 (O_1406,N_9331,N_9141);
nand UO_1407 (O_1407,N_9649,N_9223);
nand UO_1408 (O_1408,N_9524,N_9994);
nor UO_1409 (O_1409,N_9804,N_9411);
nand UO_1410 (O_1410,N_9498,N_9385);
nor UO_1411 (O_1411,N_9084,N_9971);
and UO_1412 (O_1412,N_9927,N_9461);
nor UO_1413 (O_1413,N_9990,N_9057);
nor UO_1414 (O_1414,N_9181,N_9526);
nor UO_1415 (O_1415,N_9104,N_9372);
nand UO_1416 (O_1416,N_9534,N_9253);
nor UO_1417 (O_1417,N_9150,N_9851);
and UO_1418 (O_1418,N_9646,N_9188);
nand UO_1419 (O_1419,N_9052,N_9265);
nor UO_1420 (O_1420,N_9019,N_9388);
and UO_1421 (O_1421,N_9026,N_9693);
xnor UO_1422 (O_1422,N_9799,N_9445);
nor UO_1423 (O_1423,N_9184,N_9149);
nor UO_1424 (O_1424,N_9725,N_9133);
xor UO_1425 (O_1425,N_9591,N_9614);
and UO_1426 (O_1426,N_9753,N_9373);
nor UO_1427 (O_1427,N_9497,N_9329);
nand UO_1428 (O_1428,N_9734,N_9257);
and UO_1429 (O_1429,N_9373,N_9954);
nand UO_1430 (O_1430,N_9205,N_9311);
or UO_1431 (O_1431,N_9965,N_9261);
nor UO_1432 (O_1432,N_9864,N_9430);
nand UO_1433 (O_1433,N_9195,N_9474);
and UO_1434 (O_1434,N_9168,N_9943);
nand UO_1435 (O_1435,N_9131,N_9573);
nor UO_1436 (O_1436,N_9478,N_9909);
and UO_1437 (O_1437,N_9222,N_9375);
or UO_1438 (O_1438,N_9606,N_9239);
nor UO_1439 (O_1439,N_9694,N_9758);
or UO_1440 (O_1440,N_9332,N_9878);
and UO_1441 (O_1441,N_9280,N_9509);
or UO_1442 (O_1442,N_9063,N_9163);
xnor UO_1443 (O_1443,N_9915,N_9976);
xnor UO_1444 (O_1444,N_9125,N_9969);
and UO_1445 (O_1445,N_9095,N_9742);
or UO_1446 (O_1446,N_9419,N_9830);
nor UO_1447 (O_1447,N_9799,N_9650);
nand UO_1448 (O_1448,N_9604,N_9317);
nand UO_1449 (O_1449,N_9484,N_9623);
and UO_1450 (O_1450,N_9284,N_9373);
nor UO_1451 (O_1451,N_9012,N_9382);
nor UO_1452 (O_1452,N_9035,N_9701);
nor UO_1453 (O_1453,N_9110,N_9229);
and UO_1454 (O_1454,N_9633,N_9357);
or UO_1455 (O_1455,N_9756,N_9733);
nand UO_1456 (O_1456,N_9325,N_9536);
nor UO_1457 (O_1457,N_9997,N_9674);
and UO_1458 (O_1458,N_9327,N_9121);
nor UO_1459 (O_1459,N_9402,N_9002);
or UO_1460 (O_1460,N_9787,N_9001);
or UO_1461 (O_1461,N_9681,N_9767);
nand UO_1462 (O_1462,N_9564,N_9850);
nor UO_1463 (O_1463,N_9431,N_9535);
or UO_1464 (O_1464,N_9952,N_9461);
nor UO_1465 (O_1465,N_9839,N_9844);
or UO_1466 (O_1466,N_9431,N_9202);
nand UO_1467 (O_1467,N_9863,N_9716);
nand UO_1468 (O_1468,N_9662,N_9163);
or UO_1469 (O_1469,N_9020,N_9663);
and UO_1470 (O_1470,N_9506,N_9224);
or UO_1471 (O_1471,N_9639,N_9143);
or UO_1472 (O_1472,N_9073,N_9241);
or UO_1473 (O_1473,N_9146,N_9684);
and UO_1474 (O_1474,N_9860,N_9598);
nand UO_1475 (O_1475,N_9705,N_9544);
and UO_1476 (O_1476,N_9427,N_9667);
or UO_1477 (O_1477,N_9436,N_9282);
and UO_1478 (O_1478,N_9540,N_9634);
nor UO_1479 (O_1479,N_9680,N_9421);
nand UO_1480 (O_1480,N_9206,N_9683);
nor UO_1481 (O_1481,N_9209,N_9590);
or UO_1482 (O_1482,N_9328,N_9400);
nand UO_1483 (O_1483,N_9679,N_9024);
or UO_1484 (O_1484,N_9945,N_9225);
xnor UO_1485 (O_1485,N_9582,N_9294);
nor UO_1486 (O_1486,N_9764,N_9084);
xor UO_1487 (O_1487,N_9266,N_9836);
nor UO_1488 (O_1488,N_9624,N_9867);
or UO_1489 (O_1489,N_9127,N_9587);
or UO_1490 (O_1490,N_9559,N_9878);
nor UO_1491 (O_1491,N_9598,N_9815);
nor UO_1492 (O_1492,N_9551,N_9037);
or UO_1493 (O_1493,N_9326,N_9918);
and UO_1494 (O_1494,N_9757,N_9102);
and UO_1495 (O_1495,N_9259,N_9870);
nand UO_1496 (O_1496,N_9220,N_9702);
and UO_1497 (O_1497,N_9061,N_9544);
nand UO_1498 (O_1498,N_9597,N_9146);
nand UO_1499 (O_1499,N_9533,N_9386);
endmodule