module basic_1000_10000_1500_2_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5002,N_5003,N_5005,N_5006,N_5007,N_5009,N_5011,N_5012,N_5014,N_5016,N_5017,N_5018,N_5020,N_5024,N_5025,N_5026,N_5029,N_5032,N_5033,N_5037,N_5038,N_5040,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5049,N_5050,N_5053,N_5056,N_5058,N_5062,N_5063,N_5064,N_5065,N_5066,N_5068,N_5069,N_5070,N_5071,N_5072,N_5076,N_5078,N_5079,N_5080,N_5082,N_5083,N_5086,N_5087,N_5090,N_5092,N_5093,N_5095,N_5097,N_5098,N_5103,N_5105,N_5106,N_5107,N_5108,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5119,N_5120,N_5122,N_5124,N_5125,N_5126,N_5129,N_5132,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5143,N_5144,N_5145,N_5147,N_5149,N_5151,N_5152,N_5153,N_5155,N_5156,N_5159,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5177,N_5179,N_5180,N_5181,N_5183,N_5186,N_5187,N_5188,N_5189,N_5192,N_5193,N_5195,N_5196,N_5198,N_5199,N_5200,N_5202,N_5204,N_5205,N_5206,N_5207,N_5209,N_5210,N_5212,N_5213,N_5215,N_5216,N_5219,N_5221,N_5226,N_5229,N_5231,N_5232,N_5234,N_5235,N_5236,N_5237,N_5238,N_5240,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5251,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5261,N_5262,N_5263,N_5266,N_5267,N_5272,N_5273,N_5274,N_5278,N_5279,N_5280,N_5281,N_5284,N_5285,N_5286,N_5287,N_5288,N_5290,N_5294,N_5296,N_5297,N_5298,N_5301,N_5303,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5313,N_5315,N_5318,N_5321,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5333,N_5337,N_5341,N_5342,N_5343,N_5344,N_5345,N_5347,N_5348,N_5349,N_5353,N_5355,N_5361,N_5362,N_5363,N_5364,N_5366,N_5367,N_5369,N_5371,N_5372,N_5373,N_5374,N_5376,N_5377,N_5378,N_5379,N_5380,N_5383,N_5386,N_5387,N_5389,N_5392,N_5395,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5405,N_5406,N_5407,N_5409,N_5413,N_5414,N_5415,N_5416,N_5418,N_5424,N_5425,N_5430,N_5432,N_5433,N_5435,N_5436,N_5437,N_5441,N_5443,N_5444,N_5445,N_5446,N_5447,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5460,N_5462,N_5463,N_5466,N_5467,N_5468,N_5469,N_5475,N_5476,N_5477,N_5482,N_5483,N_5484,N_5486,N_5490,N_5491,N_5493,N_5495,N_5496,N_5497,N_5498,N_5500,N_5504,N_5510,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5519,N_5520,N_5522,N_5523,N_5524,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5535,N_5538,N_5540,N_5541,N_5542,N_5546,N_5547,N_5548,N_5550,N_5551,N_5552,N_5553,N_5554,N_5557,N_5558,N_5559,N_5561,N_5562,N_5563,N_5564,N_5566,N_5567,N_5570,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5579,N_5581,N_5584,N_5585,N_5586,N_5587,N_5588,N_5591,N_5593,N_5596,N_5598,N_5600,N_5601,N_5602,N_5604,N_5605,N_5610,N_5611,N_5612,N_5613,N_5614,N_5616,N_5618,N_5619,N_5623,N_5625,N_5626,N_5627,N_5629,N_5631,N_5632,N_5633,N_5635,N_5636,N_5637,N_5638,N_5639,N_5641,N_5643,N_5644,N_5647,N_5649,N_5650,N_5652,N_5654,N_5655,N_5657,N_5659,N_5660,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5674,N_5676,N_5677,N_5678,N_5680,N_5681,N_5682,N_5686,N_5687,N_5689,N_5691,N_5693,N_5694,N_5695,N_5696,N_5699,N_5704,N_5705,N_5706,N_5709,N_5710,N_5714,N_5715,N_5720,N_5721,N_5723,N_5725,N_5726,N_5728,N_5729,N_5731,N_5733,N_5734,N_5736,N_5739,N_5741,N_5746,N_5748,N_5750,N_5751,N_5752,N_5755,N_5756,N_5757,N_5758,N_5760,N_5761,N_5762,N_5765,N_5768,N_5769,N_5771,N_5772,N_5774,N_5775,N_5776,N_5778,N_5780,N_5781,N_5782,N_5785,N_5786,N_5787,N_5789,N_5792,N_5793,N_5794,N_5795,N_5797,N_5798,N_5800,N_5801,N_5802,N_5804,N_5805,N_5806,N_5808,N_5811,N_5813,N_5814,N_5815,N_5816,N_5817,N_5819,N_5821,N_5823,N_5825,N_5826,N_5827,N_5828,N_5829,N_5834,N_5836,N_5839,N_5840,N_5841,N_5843,N_5845,N_5847,N_5848,N_5849,N_5850,N_5853,N_5857,N_5858,N_5860,N_5862,N_5863,N_5864,N_5865,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5876,N_5880,N_5882,N_5883,N_5884,N_5885,N_5886,N_5889,N_5890,N_5891,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5904,N_5905,N_5908,N_5910,N_5911,N_5912,N_5917,N_5919,N_5921,N_5923,N_5924,N_5926,N_5927,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5946,N_5948,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5960,N_5961,N_5964,N_5965,N_5966,N_5967,N_5968,N_5971,N_5972,N_5973,N_5974,N_5976,N_5977,N_5980,N_5981,N_5982,N_5986,N_5988,N_5989,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_6001,N_6002,N_6003,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6016,N_6018,N_6019,N_6020,N_6023,N_6024,N_6026,N_6027,N_6029,N_6031,N_6032,N_6033,N_6038,N_6039,N_6041,N_6042,N_6043,N_6045,N_6047,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6062,N_6063,N_6064,N_6068,N_6069,N_6072,N_6073,N_6074,N_6075,N_6077,N_6078,N_6079,N_6080,N_6081,N_6083,N_6086,N_6087,N_6091,N_6092,N_6093,N_6095,N_6100,N_6103,N_6104,N_6107,N_6109,N_6112,N_6113,N_6114,N_6116,N_6117,N_6118,N_6120,N_6121,N_6123,N_6124,N_6125,N_6127,N_6128,N_6129,N_6132,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6149,N_6151,N_6153,N_6154,N_6157,N_6158,N_6159,N_6160,N_6162,N_6164,N_6166,N_6168,N_6171,N_6172,N_6173,N_6174,N_6178,N_6179,N_6182,N_6184,N_6185,N_6186,N_6187,N_6191,N_6192,N_6193,N_6194,N_6195,N_6198,N_6199,N_6200,N_6202,N_6203,N_6204,N_6205,N_6208,N_6209,N_6211,N_6212,N_6215,N_6216,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6227,N_6228,N_6231,N_6232,N_6233,N_6234,N_6235,N_6239,N_6240,N_6242,N_6245,N_6246,N_6247,N_6249,N_6250,N_6251,N_6253,N_6254,N_6255,N_6256,N_6260,N_6264,N_6265,N_6266,N_6269,N_6270,N_6273,N_6276,N_6277,N_6278,N_6279,N_6280,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6298,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6308,N_6317,N_6319,N_6320,N_6321,N_6324,N_6325,N_6326,N_6327,N_6334,N_6338,N_6340,N_6341,N_6342,N_6343,N_6344,N_6346,N_6347,N_6349,N_6350,N_6351,N_6354,N_6356,N_6358,N_6359,N_6360,N_6361,N_6362,N_6364,N_6366,N_6367,N_6370,N_6372,N_6374,N_6375,N_6378,N_6381,N_6387,N_6390,N_6392,N_6394,N_6396,N_6398,N_6400,N_6401,N_6402,N_6406,N_6409,N_6410,N_6412,N_6414,N_6415,N_6416,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6427,N_6428,N_6429,N_6430,N_6434,N_6440,N_6443,N_6447,N_6448,N_6450,N_6453,N_6454,N_6455,N_6456,N_6457,N_6459,N_6461,N_6463,N_6464,N_6467,N_6469,N_6470,N_6471,N_6472,N_6477,N_6478,N_6479,N_6480,N_6483,N_6484,N_6485,N_6493,N_6494,N_6496,N_6498,N_6499,N_6501,N_6502,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6516,N_6517,N_6523,N_6524,N_6525,N_6526,N_6527,N_6529,N_6530,N_6532,N_6533,N_6534,N_6535,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6553,N_6556,N_6558,N_6559,N_6560,N_6562,N_6563,N_6565,N_6567,N_6568,N_6571,N_6573,N_6574,N_6576,N_6577,N_6578,N_6579,N_6582,N_6583,N_6584,N_6586,N_6587,N_6588,N_6590,N_6592,N_6594,N_6596,N_6597,N_6598,N_6599,N_6600,N_6603,N_6604,N_6605,N_6611,N_6612,N_6614,N_6615,N_6616,N_6617,N_6619,N_6620,N_6623,N_6624,N_6625,N_6626,N_6627,N_6629,N_6631,N_6634,N_6635,N_6636,N_6639,N_6640,N_6641,N_6643,N_6649,N_6650,N_6651,N_6652,N_6654,N_6655,N_6656,N_6657,N_6658,N_6660,N_6661,N_6662,N_6663,N_6665,N_6668,N_6670,N_6674,N_6677,N_6678,N_6680,N_6681,N_6682,N_6684,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6696,N_6697,N_6698,N_6699,N_6700,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6711,N_6712,N_6713,N_6714,N_6716,N_6718,N_6719,N_6720,N_6721,N_6722,N_6724,N_6725,N_6727,N_6729,N_6730,N_6732,N_6733,N_6735,N_6736,N_6737,N_6739,N_6741,N_6742,N_6743,N_6744,N_6746,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6755,N_6756,N_6757,N_6758,N_6759,N_6761,N_6765,N_6769,N_6770,N_6772,N_6774,N_6776,N_6777,N_6779,N_6780,N_6781,N_6783,N_6786,N_6792,N_6794,N_6795,N_6796,N_6800,N_6802,N_6803,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6814,N_6815,N_6816,N_6817,N_6824,N_6825,N_6830,N_6831,N_6832,N_6834,N_6835,N_6836,N_6837,N_6838,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6850,N_6851,N_6853,N_6855,N_6857,N_6859,N_6860,N_6862,N_6863,N_6864,N_6865,N_6866,N_6868,N_6871,N_6873,N_6876,N_6877,N_6878,N_6883,N_6885,N_6887,N_6888,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6897,N_6899,N_6900,N_6901,N_6902,N_6904,N_6905,N_6911,N_6919,N_6920,N_6921,N_6922,N_6924,N_6925,N_6930,N_6931,N_6935,N_6937,N_6939,N_6940,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6958,N_6959,N_6960,N_6962,N_6963,N_6964,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6986,N_6987,N_6988,N_6990,N_6993,N_6997,N_6999,N_7001,N_7002,N_7004,N_7006,N_7007,N_7011,N_7012,N_7013,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7023,N_7024,N_7026,N_7027,N_7030,N_7032,N_7033,N_7034,N_7037,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7047,N_7048,N_7050,N_7051,N_7053,N_7054,N_7055,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7067,N_7070,N_7071,N_7072,N_7074,N_7076,N_7077,N_7079,N_7080,N_7082,N_7084,N_7085,N_7087,N_7088,N_7090,N_7093,N_7094,N_7095,N_7098,N_7100,N_7101,N_7103,N_7104,N_7105,N_7106,N_7108,N_7111,N_7112,N_7114,N_7116,N_7117,N_7118,N_7119,N_7120,N_7125,N_7126,N_7127,N_7129,N_7130,N_7132,N_7134,N_7135,N_7138,N_7139,N_7140,N_7141,N_7145,N_7146,N_7147,N_7148,N_7150,N_7151,N_7155,N_7158,N_7160,N_7162,N_7166,N_7167,N_7170,N_7171,N_7172,N_7173,N_7174,N_7176,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7187,N_7188,N_7192,N_7193,N_7194,N_7195,N_7196,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7210,N_7212,N_7214,N_7215,N_7217,N_7218,N_7220,N_7221,N_7223,N_7224,N_7228,N_7231,N_7232,N_7233,N_7235,N_7236,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7246,N_7250,N_7253,N_7255,N_7256,N_7257,N_7258,N_7260,N_7261,N_7262,N_7266,N_7267,N_7269,N_7270,N_7271,N_7272,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7284,N_7285,N_7286,N_7288,N_7291,N_7292,N_7293,N_7294,N_7297,N_7298,N_7300,N_7302,N_7303,N_7306,N_7307,N_7308,N_7310,N_7313,N_7315,N_7316,N_7317,N_7318,N_7320,N_7321,N_7322,N_7323,N_7324,N_7326,N_7327,N_7329,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7343,N_7344,N_7345,N_7348,N_7350,N_7351,N_7352,N_7353,N_7356,N_7360,N_7361,N_7364,N_7365,N_7367,N_7368,N_7369,N_7372,N_7373,N_7375,N_7376,N_7377,N_7380,N_7383,N_7384,N_7386,N_7387,N_7388,N_7391,N_7393,N_7395,N_7398,N_7400,N_7402,N_7403,N_7404,N_7406,N_7407,N_7408,N_7411,N_7412,N_7416,N_7418,N_7419,N_7420,N_7423,N_7426,N_7427,N_7431,N_7433,N_7434,N_7436,N_7438,N_7441,N_7442,N_7443,N_7444,N_7445,N_7450,N_7458,N_7459,N_7460,N_7461,N_7463,N_7464,N_7465,N_7468,N_7469,N_7470,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7488,N_7490,N_7491,N_7499,N_7500,N_7505,N_7509,N_7510,N_7513,N_7514,N_7515,N_7516,N_7518,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7529,N_7530,N_7531,N_7535,N_7536,N_7539,N_7541,N_7542,N_7543,N_7544,N_7548,N_7549,N_7552,N_7554,N_7556,N_7557,N_7558,N_7560,N_7562,N_7564,N_7565,N_7567,N_7569,N_7571,N_7572,N_7576,N_7578,N_7580,N_7583,N_7586,N_7588,N_7592,N_7593,N_7594,N_7597,N_7598,N_7599,N_7601,N_7602,N_7604,N_7605,N_7606,N_7610,N_7613,N_7614,N_7618,N_7620,N_7621,N_7624,N_7625,N_7628,N_7632,N_7634,N_7639,N_7641,N_7642,N_7643,N_7648,N_7650,N_7651,N_7652,N_7653,N_7656,N_7657,N_7658,N_7660,N_7661,N_7662,N_7664,N_7665,N_7670,N_7671,N_7672,N_7673,N_7675,N_7676,N_7677,N_7679,N_7680,N_7681,N_7682,N_7684,N_7685,N_7687,N_7688,N_7689,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7699,N_7701,N_7702,N_7703,N_7707,N_7709,N_7710,N_7713,N_7717,N_7719,N_7720,N_7723,N_7726,N_7728,N_7734,N_7736,N_7737,N_7739,N_7740,N_7741,N_7746,N_7748,N_7749,N_7751,N_7752,N_7753,N_7755,N_7756,N_7760,N_7762,N_7767,N_7768,N_7769,N_7770,N_7771,N_7775,N_7776,N_7780,N_7783,N_7785,N_7786,N_7789,N_7792,N_7793,N_7795,N_7796,N_7799,N_7800,N_7801,N_7802,N_7804,N_7805,N_7806,N_7807,N_7808,N_7810,N_7812,N_7815,N_7816,N_7818,N_7819,N_7821,N_7822,N_7824,N_7825,N_7828,N_7829,N_7830,N_7834,N_7835,N_7837,N_7838,N_7839,N_7842,N_7844,N_7845,N_7846,N_7847,N_7848,N_7850,N_7851,N_7852,N_7854,N_7855,N_7857,N_7858,N_7860,N_7861,N_7862,N_7863,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7872,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7885,N_7886,N_7887,N_7889,N_7893,N_7895,N_7896,N_7897,N_7899,N_7900,N_7901,N_7903,N_7904,N_7905,N_7906,N_7910,N_7911,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7920,N_7922,N_7923,N_7925,N_7927,N_7928,N_7929,N_7931,N_7932,N_7933,N_7935,N_7938,N_7939,N_7940,N_7941,N_7942,N_7945,N_7949,N_7950,N_7956,N_7957,N_7959,N_7965,N_7966,N_7968,N_7969,N_7973,N_7975,N_7976,N_7977,N_7979,N_7980,N_7981,N_7983,N_7984,N_7986,N_7988,N_7990,N_7992,N_7993,N_7994,N_7995,N_7996,N_7998,N_8000,N_8001,N_8003,N_8006,N_8007,N_8008,N_8009,N_8010,N_8012,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8021,N_8023,N_8025,N_8026,N_8027,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8039,N_8040,N_8041,N_8043,N_8044,N_8046,N_8047,N_8049,N_8050,N_8051,N_8052,N_8053,N_8056,N_8057,N_8058,N_8059,N_8060,N_8062,N_8063,N_8065,N_8066,N_8068,N_8069,N_8074,N_8076,N_8077,N_8078,N_8081,N_8083,N_8084,N_8085,N_8086,N_8087,N_8091,N_8094,N_8095,N_8098,N_8099,N_8100,N_8101,N_8103,N_8105,N_8106,N_8108,N_8109,N_8110,N_8112,N_8114,N_8115,N_8117,N_8119,N_8121,N_8123,N_8124,N_8125,N_8128,N_8130,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8139,N_8144,N_8145,N_8146,N_8147,N_8152,N_8157,N_8158,N_8160,N_8161,N_8163,N_8165,N_8171,N_8172,N_8173,N_8175,N_8176,N_8178,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8202,N_8203,N_8204,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8222,N_8223,N_8224,N_8227,N_8228,N_8229,N_8232,N_8234,N_8236,N_8237,N_8239,N_8240,N_8243,N_8244,N_8248,N_8249,N_8251,N_8253,N_8254,N_8258,N_8259,N_8260,N_8262,N_8264,N_8265,N_8268,N_8269,N_8271,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8283,N_8287,N_8291,N_8292,N_8295,N_8297,N_8298,N_8301,N_8306,N_8307,N_8309,N_8310,N_8312,N_8313,N_8314,N_8315,N_8318,N_8320,N_8322,N_8324,N_8325,N_8327,N_8331,N_8332,N_8334,N_8336,N_8337,N_8338,N_8339,N_8342,N_8343,N_8345,N_8346,N_8348,N_8349,N_8350,N_8352,N_8354,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8363,N_8364,N_8369,N_8370,N_8374,N_8376,N_8377,N_8379,N_8383,N_8385,N_8386,N_8387,N_8389,N_8393,N_8394,N_8397,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8407,N_8408,N_8409,N_8412,N_8413,N_8414,N_8416,N_8417,N_8418,N_8421,N_8422,N_8423,N_8425,N_8427,N_8428,N_8429,N_8430,N_8432,N_8433,N_8434,N_8435,N_8436,N_8438,N_8439,N_8442,N_8443,N_8444,N_8445,N_8446,N_8448,N_8449,N_8450,N_8451,N_8452,N_8456,N_8458,N_8459,N_8460,N_8461,N_8465,N_8466,N_8467,N_8469,N_8471,N_8473,N_8479,N_8480,N_8482,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8491,N_8496,N_8500,N_8501,N_8504,N_8505,N_8509,N_8511,N_8512,N_8514,N_8517,N_8518,N_8519,N_8521,N_8523,N_8524,N_8525,N_8526,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8539,N_8540,N_8541,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8552,N_8556,N_8558,N_8559,N_8560,N_8562,N_8564,N_8566,N_8567,N_8568,N_8569,N_8570,N_8572,N_8573,N_8575,N_8578,N_8580,N_8582,N_8584,N_8585,N_8586,N_8588,N_8589,N_8592,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8605,N_8608,N_8609,N_8610,N_8612,N_8613,N_8615,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8627,N_8628,N_8629,N_8630,N_8631,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8646,N_8648,N_8649,N_8651,N_8652,N_8653,N_8655,N_8656,N_8657,N_8659,N_8663,N_8664,N_8665,N_8666,N_8667,N_8669,N_8670,N_8671,N_8676,N_8679,N_8681,N_8682,N_8683,N_8684,N_8685,N_8688,N_8689,N_8693,N_8698,N_8699,N_8701,N_8707,N_8708,N_8709,N_8711,N_8712,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8726,N_8727,N_8730,N_8733,N_8734,N_8735,N_8736,N_8740,N_8741,N_8742,N_8743,N_8744,N_8747,N_8748,N_8751,N_8752,N_8753,N_8755,N_8756,N_8757,N_8758,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8772,N_8773,N_8775,N_8776,N_8777,N_8780,N_8782,N_8783,N_8786,N_8787,N_8788,N_8790,N_8791,N_8792,N_8795,N_8796,N_8797,N_8799,N_8800,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8818,N_8819,N_8821,N_8822,N_8823,N_8829,N_8830,N_8831,N_8832,N_8836,N_8841,N_8843,N_8844,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8858,N_8859,N_8860,N_8861,N_8866,N_8867,N_8869,N_8870,N_8871,N_8875,N_8876,N_8877,N_8878,N_8879,N_8881,N_8884,N_8885,N_8886,N_8887,N_8890,N_8891,N_8892,N_8894,N_8897,N_8898,N_8899,N_8902,N_8906,N_8907,N_8909,N_8912,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8926,N_8930,N_8933,N_8934,N_8935,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8944,N_8945,N_8946,N_8948,N_8950,N_8951,N_8953,N_8954,N_8955,N_8956,N_8958,N_8959,N_8960,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8969,N_8970,N_8971,N_8975,N_8977,N_8979,N_8980,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8992,N_8993,N_8994,N_8995,N_8996,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9007,N_9008,N_9010,N_9011,N_9013,N_9015,N_9024,N_9025,N_9026,N_9027,N_9029,N_9030,N_9031,N_9033,N_9035,N_9036,N_9038,N_9040,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9053,N_9060,N_9061,N_9064,N_9065,N_9067,N_9069,N_9070,N_9071,N_9072,N_9074,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9088,N_9089,N_9091,N_9092,N_9093,N_9094,N_9096,N_9097,N_9099,N_9100,N_9101,N_9103,N_9104,N_9106,N_9107,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9116,N_9118,N_9119,N_9120,N_9121,N_9123,N_9124,N_9125,N_9126,N_9127,N_9129,N_9133,N_9134,N_9135,N_9137,N_9139,N_9141,N_9142,N_9144,N_9145,N_9146,N_9147,N_9149,N_9152,N_9154,N_9155,N_9158,N_9161,N_9162,N_9163,N_9164,N_9165,N_9167,N_9168,N_9172,N_9173,N_9174,N_9175,N_9178,N_9179,N_9180,N_9183,N_9186,N_9187,N_9189,N_9195,N_9200,N_9202,N_9203,N_9206,N_9207,N_9209,N_9210,N_9213,N_9214,N_9216,N_9221,N_9222,N_9223,N_9227,N_9231,N_9234,N_9235,N_9237,N_9238,N_9242,N_9245,N_9247,N_9248,N_9252,N_9253,N_9255,N_9256,N_9258,N_9259,N_9260,N_9261,N_9263,N_9264,N_9265,N_9266,N_9267,N_9269,N_9270,N_9272,N_9275,N_9278,N_9280,N_9281,N_9282,N_9283,N_9285,N_9289,N_9290,N_9292,N_9294,N_9295,N_9296,N_9298,N_9299,N_9300,N_9301,N_9303,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9315,N_9316,N_9317,N_9318,N_9321,N_9322,N_9324,N_9325,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9336,N_9337,N_9339,N_9341,N_9342,N_9345,N_9348,N_9349,N_9351,N_9353,N_9354,N_9355,N_9360,N_9361,N_9364,N_9365,N_9366,N_9369,N_9370,N_9371,N_9373,N_9375,N_9376,N_9377,N_9379,N_9381,N_9382,N_9388,N_9390,N_9395,N_9397,N_9401,N_9403,N_9405,N_9408,N_9409,N_9410,N_9411,N_9413,N_9414,N_9417,N_9420,N_9421,N_9424,N_9425,N_9426,N_9427,N_9428,N_9430,N_9431,N_9435,N_9436,N_9437,N_9439,N_9444,N_9445,N_9447,N_9449,N_9451,N_9452,N_9455,N_9456,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9465,N_9469,N_9474,N_9476,N_9478,N_9482,N_9483,N_9484,N_9486,N_9488,N_9489,N_9490,N_9491,N_9493,N_9494,N_9495,N_9498,N_9499,N_9500,N_9501,N_9503,N_9504,N_9505,N_9506,N_9508,N_9509,N_9510,N_9511,N_9512,N_9514,N_9518,N_9521,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9531,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9540,N_9541,N_9542,N_9543,N_9544,N_9546,N_9547,N_9549,N_9550,N_9551,N_9552,N_9553,N_9558,N_9559,N_9561,N_9562,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9571,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9585,N_9588,N_9590,N_9594,N_9596,N_9600,N_9605,N_9607,N_9608,N_9610,N_9612,N_9613,N_9614,N_9615,N_9616,N_9618,N_9621,N_9626,N_9627,N_9629,N_9633,N_9634,N_9636,N_9637,N_9638,N_9639,N_9641,N_9642,N_9643,N_9645,N_9646,N_9648,N_9649,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9662,N_9663,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9672,N_9673,N_9675,N_9679,N_9680,N_9681,N_9682,N_9684,N_9685,N_9686,N_9687,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9696,N_9698,N_9699,N_9701,N_9704,N_9705,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9715,N_9716,N_9717,N_9718,N_9719,N_9721,N_9724,N_9725,N_9727,N_9728,N_9737,N_9739,N_9740,N_9741,N_9743,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9757,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9767,N_9771,N_9772,N_9777,N_9779,N_9781,N_9784,N_9785,N_9786,N_9787,N_9788,N_9791,N_9793,N_9794,N_9797,N_9800,N_9803,N_9804,N_9805,N_9807,N_9808,N_9809,N_9811,N_9814,N_9816,N_9817,N_9818,N_9820,N_9821,N_9822,N_9825,N_9826,N_9827,N_9830,N_9831,N_9832,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9842,N_9843,N_9845,N_9847,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9856,N_9857,N_9859,N_9860,N_9865,N_9866,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9878,N_9879,N_9881,N_9883,N_9884,N_9885,N_9886,N_9887,N_9890,N_9892,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9903,N_9904,N_9905,N_9907,N_9909,N_9910,N_9912,N_9913,N_9914,N_9915,N_9917,N_9919,N_9920,N_9922,N_9923,N_9925,N_9927,N_9931,N_9932,N_9933,N_9934,N_9937,N_9940,N_9941,N_9945,N_9947,N_9949,N_9951,N_9952,N_9953,N_9954,N_9956,N_9957,N_9959,N_9961,N_9963,N_9965,N_9966,N_9967,N_9968,N_9969,N_9971,N_9972,N_9976,N_9977,N_9978,N_9980,N_9982,N_9984,N_9986,N_9987,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9999;
xnor U0 (N_0,In_250,In_919);
nor U1 (N_1,In_133,In_541);
nor U2 (N_2,In_800,In_635);
and U3 (N_3,In_535,In_963);
nor U4 (N_4,In_3,In_164);
or U5 (N_5,In_20,In_586);
nand U6 (N_6,In_490,In_663);
or U7 (N_7,In_654,In_391);
and U8 (N_8,In_634,In_448);
nor U9 (N_9,In_820,In_273);
nor U10 (N_10,In_5,In_503);
nor U11 (N_11,In_386,In_486);
or U12 (N_12,In_18,In_776);
and U13 (N_13,In_153,In_210);
nor U14 (N_14,In_242,In_304);
nand U15 (N_15,In_425,In_353);
nor U16 (N_16,In_642,In_840);
nand U17 (N_17,In_687,In_804);
xnor U18 (N_18,In_315,In_599);
xnor U19 (N_19,In_990,In_430);
nand U20 (N_20,In_884,In_505);
or U21 (N_21,In_621,In_213);
nor U22 (N_22,In_548,In_893);
or U23 (N_23,In_674,In_936);
xor U24 (N_24,In_516,In_773);
or U25 (N_25,In_596,In_724);
and U26 (N_26,In_131,In_461);
and U27 (N_27,In_441,In_581);
nor U28 (N_28,In_246,In_366);
nand U29 (N_29,In_392,In_137);
or U30 (N_30,In_514,In_98);
xor U31 (N_31,In_338,In_54);
nand U32 (N_32,In_385,In_382);
or U33 (N_33,In_829,In_428);
or U34 (N_34,In_355,In_127);
nor U35 (N_35,In_523,In_595);
and U36 (N_36,In_746,In_194);
nor U37 (N_37,In_288,In_331);
and U38 (N_38,In_653,In_563);
or U39 (N_39,In_381,In_55);
or U40 (N_40,In_286,In_670);
nor U41 (N_41,In_732,In_429);
and U42 (N_42,In_705,In_843);
or U43 (N_43,In_7,In_301);
xnor U44 (N_44,In_664,In_142);
nor U45 (N_45,In_313,In_260);
and U46 (N_46,In_717,In_43);
nand U47 (N_47,In_601,In_460);
or U48 (N_48,In_178,In_584);
nand U49 (N_49,In_302,In_45);
nand U50 (N_50,In_512,In_4);
nand U51 (N_51,In_684,In_110);
or U52 (N_52,In_940,In_193);
and U53 (N_53,In_998,In_58);
or U54 (N_54,In_417,In_408);
nor U55 (N_55,In_332,In_423);
nand U56 (N_56,In_855,In_52);
xor U57 (N_57,In_587,In_256);
nor U58 (N_58,In_731,In_658);
or U59 (N_59,In_585,In_309);
or U60 (N_60,In_147,In_934);
or U61 (N_61,In_853,In_583);
nor U62 (N_62,In_442,In_868);
nand U63 (N_63,In_798,In_76);
and U64 (N_64,In_36,In_343);
and U65 (N_65,In_463,In_368);
or U66 (N_66,In_867,In_96);
nand U67 (N_67,In_565,In_220);
and U68 (N_68,In_668,In_680);
xnor U69 (N_69,In_825,In_190);
or U70 (N_70,In_140,In_292);
nor U71 (N_71,In_501,In_721);
nand U72 (N_72,In_413,In_28);
or U73 (N_73,In_44,In_645);
nor U74 (N_74,In_966,In_434);
and U75 (N_75,In_768,In_784);
xnor U76 (N_76,In_561,In_470);
nand U77 (N_77,In_443,In_606);
xor U78 (N_78,In_907,In_613);
nor U79 (N_79,In_239,In_822);
or U80 (N_80,In_277,In_232);
and U81 (N_81,In_949,In_556);
or U82 (N_82,In_830,In_667);
nand U83 (N_83,In_754,In_981);
or U84 (N_84,In_276,In_787);
xor U85 (N_85,In_412,In_376);
or U86 (N_86,In_219,In_150);
nand U87 (N_87,In_504,In_805);
and U88 (N_88,In_396,In_719);
nor U89 (N_89,In_83,In_706);
nand U90 (N_90,In_681,In_553);
or U91 (N_91,In_802,In_749);
nand U92 (N_92,In_708,In_729);
nor U93 (N_93,In_812,In_701);
nand U94 (N_94,In_121,In_351);
and U95 (N_95,In_437,In_471);
or U96 (N_96,In_290,In_115);
xnor U97 (N_97,In_593,In_818);
nor U98 (N_98,In_515,In_559);
nor U99 (N_99,In_750,In_475);
or U100 (N_100,In_679,In_326);
nand U101 (N_101,In_165,In_577);
nor U102 (N_102,In_502,In_569);
or U103 (N_103,In_212,In_207);
or U104 (N_104,In_864,In_499);
xnor U105 (N_105,In_252,In_143);
nor U106 (N_106,In_325,In_828);
or U107 (N_107,In_965,In_821);
nor U108 (N_108,In_298,In_100);
nand U109 (N_109,In_106,In_50);
xnor U110 (N_110,In_904,In_925);
or U111 (N_111,In_69,In_689);
nand U112 (N_112,In_259,In_712);
and U113 (N_113,In_216,In_330);
and U114 (N_114,In_878,In_957);
nand U115 (N_115,In_780,In_967);
nand U116 (N_116,In_94,In_415);
and U117 (N_117,In_92,In_467);
and U118 (N_118,In_874,In_474);
xor U119 (N_119,In_384,In_192);
and U120 (N_120,In_937,In_163);
or U121 (N_121,In_543,In_342);
or U122 (N_122,In_209,In_540);
or U123 (N_123,In_402,In_972);
xor U124 (N_124,In_751,In_638);
and U125 (N_125,In_988,In_579);
and U126 (N_126,In_615,In_880);
and U127 (N_127,In_57,In_611);
and U128 (N_128,In_699,In_319);
xor U129 (N_129,In_660,In_155);
and U130 (N_130,In_51,In_995);
or U131 (N_131,In_9,In_123);
nand U132 (N_132,In_172,In_973);
or U133 (N_133,In_694,In_624);
nand U134 (N_134,In_419,In_335);
or U135 (N_135,In_234,In_617);
nand U136 (N_136,In_267,In_803);
nand U137 (N_137,In_1,In_145);
nand U138 (N_138,In_418,In_608);
nand U139 (N_139,In_400,In_598);
nor U140 (N_140,In_347,In_930);
or U141 (N_141,In_77,In_589);
nand U142 (N_142,In_727,In_865);
nor U143 (N_143,In_819,In_378);
nand U144 (N_144,In_592,In_462);
nor U145 (N_145,In_861,In_375);
nand U146 (N_146,In_745,In_258);
or U147 (N_147,In_836,In_785);
nor U148 (N_148,In_170,In_275);
xnor U149 (N_149,In_85,In_198);
xnor U150 (N_150,In_683,In_328);
nor U151 (N_151,In_648,In_520);
xor U152 (N_152,In_139,In_926);
xnor U153 (N_153,In_436,In_126);
and U154 (N_154,In_394,In_446);
nand U155 (N_155,In_824,In_715);
nor U156 (N_156,In_756,In_237);
and U157 (N_157,In_488,In_775);
or U158 (N_158,In_726,In_336);
and U159 (N_159,In_612,In_66);
and U160 (N_160,In_445,In_703);
or U161 (N_161,In_0,In_734);
xnor U162 (N_162,In_112,In_901);
nand U163 (N_163,In_90,In_823);
nand U164 (N_164,In_892,In_360);
nand U165 (N_165,In_883,In_716);
nand U166 (N_166,In_591,In_32);
nand U167 (N_167,In_380,In_558);
or U168 (N_168,In_424,In_295);
nand U169 (N_169,In_594,In_568);
xor U170 (N_170,In_103,In_969);
xor U171 (N_171,In_196,In_269);
nand U172 (N_172,In_566,In_68);
nand U173 (N_173,In_690,In_320);
or U174 (N_174,In_24,In_265);
nor U175 (N_175,In_280,In_793);
and U176 (N_176,In_984,In_813);
or U177 (N_177,In_204,In_493);
xor U178 (N_178,In_607,In_151);
or U179 (N_179,In_468,In_377);
and U180 (N_180,In_317,In_796);
and U181 (N_181,In_809,In_911);
xnor U182 (N_182,In_225,In_346);
and U183 (N_183,In_946,In_903);
nand U184 (N_184,In_910,In_420);
xnor U185 (N_185,In_801,In_134);
and U186 (N_186,In_233,In_405);
and U187 (N_187,In_261,In_114);
nor U188 (N_188,In_158,In_497);
xor U189 (N_189,In_955,In_154);
or U190 (N_190,In_455,In_238);
or U191 (N_191,In_482,In_469);
nand U192 (N_192,In_622,In_152);
nor U193 (N_193,In_923,In_383);
or U194 (N_194,In_950,In_177);
and U195 (N_195,In_53,In_920);
and U196 (N_196,In_19,In_310);
xnor U197 (N_197,In_842,In_171);
nand U198 (N_198,In_922,In_677);
nor U199 (N_199,In_673,In_846);
and U200 (N_200,In_120,In_167);
nor U201 (N_201,In_244,In_827);
or U202 (N_202,In_831,In_691);
nand U203 (N_203,In_480,In_144);
and U204 (N_204,In_976,In_929);
nand U205 (N_205,In_248,In_199);
or U206 (N_206,In_464,In_270);
xnor U207 (N_207,In_21,In_156);
or U208 (N_208,In_637,In_928);
xor U209 (N_209,In_580,In_859);
or U210 (N_210,In_851,In_38);
and U211 (N_211,In_241,In_839);
xor U212 (N_212,In_725,In_974);
or U213 (N_213,In_27,In_125);
nand U214 (N_214,In_697,In_743);
and U215 (N_215,In_254,In_870);
nor U216 (N_216,In_747,In_771);
nor U217 (N_217,In_539,In_647);
nand U218 (N_218,In_40,In_485);
nor U219 (N_219,In_882,In_266);
or U220 (N_220,In_181,In_856);
and U221 (N_221,In_61,In_941);
and U222 (N_222,In_849,In_649);
and U223 (N_223,In_274,In_47);
nor U224 (N_224,In_666,In_411);
nand U225 (N_225,In_426,In_627);
and U226 (N_226,In_682,In_14);
or U227 (N_227,In_772,In_980);
and U228 (N_228,In_404,In_958);
and U229 (N_229,In_174,In_834);
and U230 (N_230,In_761,In_959);
or U231 (N_231,In_961,In_932);
or U232 (N_232,In_487,In_432);
and U233 (N_233,In_473,In_105);
and U234 (N_234,In_327,In_217);
and U235 (N_235,In_902,In_46);
or U236 (N_236,In_372,In_183);
nand U237 (N_237,In_169,In_73);
or U238 (N_238,In_102,In_887);
nor U239 (N_239,In_264,In_202);
nand U240 (N_240,In_308,In_625);
nor U241 (N_241,In_449,In_996);
nor U242 (N_242,In_365,In_816);
and U243 (N_243,In_844,In_989);
and U244 (N_244,In_531,In_945);
or U245 (N_245,In_733,In_547);
or U246 (N_246,In_221,In_953);
nand U247 (N_247,In_42,In_511);
nor U248 (N_248,In_713,In_696);
and U249 (N_249,In_86,In_354);
and U250 (N_250,In_116,In_435);
or U251 (N_251,In_362,In_885);
nand U252 (N_252,In_709,In_453);
nand U253 (N_253,In_550,In_909);
nand U254 (N_254,In_906,In_857);
xor U255 (N_255,In_530,In_492);
or U256 (N_256,In_337,In_519);
nor U257 (N_257,In_281,In_296);
nor U258 (N_258,In_186,In_597);
and U259 (N_259,In_552,In_80);
and U260 (N_260,In_675,In_466);
or U261 (N_261,In_847,In_321);
nand U262 (N_262,In_191,In_15);
nor U263 (N_263,In_588,In_769);
nand U264 (N_264,In_364,In_282);
nand U265 (N_265,In_350,In_791);
nand U266 (N_266,In_837,In_939);
nor U267 (N_267,In_763,In_977);
nor U268 (N_268,In_549,In_799);
nand U269 (N_269,In_740,In_875);
or U270 (N_270,In_189,In_722);
or U271 (N_271,In_214,In_529);
nor U272 (N_272,In_444,In_723);
and U273 (N_273,In_104,In_860);
xnor U274 (N_274,In_532,In_924);
or U275 (N_275,In_498,In_95);
and U276 (N_276,In_452,In_367);
or U277 (N_277,In_245,In_574);
nand U278 (N_278,In_287,In_111);
or U279 (N_279,In_333,In_56);
nand U280 (N_280,In_927,In_454);
and U281 (N_281,In_863,In_91);
xnor U282 (N_282,In_915,In_669);
nand U283 (N_283,In_971,In_869);
or U284 (N_284,In_149,In_390);
or U285 (N_285,In_26,In_345);
or U286 (N_286,In_833,In_401);
nand U287 (N_287,In_176,In_852);
and U288 (N_288,In_711,In_358);
nor U289 (N_289,In_741,In_873);
or U290 (N_290,In_753,In_630);
xnor U291 (N_291,In_182,In_900);
nand U292 (N_292,In_693,In_421);
nand U293 (N_293,In_369,In_166);
nand U294 (N_294,In_628,In_952);
and U295 (N_295,In_916,In_465);
nand U296 (N_296,In_278,In_71);
or U297 (N_297,In_807,In_293);
xor U298 (N_298,In_399,In_510);
or U299 (N_299,In_704,In_67);
or U300 (N_300,In_742,In_982);
nand U301 (N_301,In_113,In_616);
or U302 (N_302,In_70,In_243);
nand U303 (N_303,In_921,In_618);
and U304 (N_304,In_665,In_636);
or U305 (N_305,In_477,In_25);
xor U306 (N_306,In_757,In_554);
and U307 (N_307,In_59,In_895);
nand U308 (N_308,In_748,In_789);
and U309 (N_309,In_656,In_10);
nor U310 (N_310,In_23,In_536);
nand U311 (N_311,In_605,In_294);
nor U312 (N_312,In_999,In_12);
and U313 (N_313,In_912,In_758);
nand U314 (N_314,In_373,In_218);
nor U315 (N_315,In_129,In_792);
nor U316 (N_316,In_513,In_271);
or U317 (N_317,In_947,In_251);
or U318 (N_318,In_978,In_406);
and U319 (N_319,In_652,In_544);
xor U320 (N_320,In_324,In_983);
nand U321 (N_321,In_457,In_600);
or U322 (N_322,In_815,In_570);
nand U323 (N_323,In_227,In_363);
or U324 (N_324,In_744,In_135);
nand U325 (N_325,In_307,In_279);
xor U326 (N_326,In_890,In_13);
nand U327 (N_327,In_943,In_956);
nand U328 (N_328,In_604,In_838);
nand U329 (N_329,In_179,In_714);
and U330 (N_330,In_22,In_555);
xnor U331 (N_331,In_872,In_311);
xor U332 (N_332,In_894,In_93);
nor U333 (N_333,In_908,In_187);
nand U334 (N_334,In_388,In_986);
and U335 (N_335,In_99,In_215);
nor U336 (N_336,In_707,In_289);
or U337 (N_337,In_898,In_272);
xor U338 (N_338,In_759,In_889);
nand U339 (N_339,In_357,In_942);
and U340 (N_340,In_688,In_397);
or U341 (N_341,In_695,In_334);
nand U342 (N_342,In_74,In_879);
or U343 (N_343,In_284,In_546);
and U344 (N_344,In_948,In_557);
nor U345 (N_345,In_795,In_678);
nor U346 (N_346,In_180,In_63);
or U347 (N_347,In_283,In_30);
xnor U348 (N_348,In_130,In_231);
or U349 (N_349,In_205,In_409);
or U350 (N_350,In_938,In_542);
or U351 (N_351,In_291,In_854);
or U352 (N_352,In_632,In_479);
and U353 (N_353,In_814,In_779);
nor U354 (N_354,In_657,In_760);
xnor U355 (N_355,In_808,In_109);
and U356 (N_356,In_300,In_933);
xor U357 (N_357,In_136,In_571);
or U358 (N_358,In_175,In_146);
nor U359 (N_359,In_886,In_782);
nor U360 (N_360,In_702,In_602);
or U361 (N_361,In_371,In_728);
nand U362 (N_362,In_676,In_262);
nor U363 (N_363,In_229,In_159);
nor U364 (N_364,In_459,In_75);
xor U365 (N_365,In_484,In_806);
nor U366 (N_366,In_440,In_528);
and U367 (N_367,In_438,In_395);
and U368 (N_368,In_81,In_49);
xor U369 (N_369,In_609,In_562);
nor U370 (N_370,In_496,In_764);
nand U371 (N_371,In_370,In_157);
and U372 (N_372,In_97,In_379);
and U373 (N_373,In_788,In_876);
nor U374 (N_374,In_2,In_456);
nand U375 (N_375,In_877,In_521);
or U376 (N_376,In_686,In_817);
and U377 (N_377,In_619,In_348);
nand U378 (N_378,In_640,In_564);
or U379 (N_379,In_11,In_850);
nor U380 (N_380,In_810,In_845);
nor U381 (N_381,In_551,In_89);
and U382 (N_382,In_235,In_299);
nand U383 (N_383,In_344,In_314);
nand U384 (N_384,In_361,In_603);
or U385 (N_385,In_662,In_794);
or U386 (N_386,In_862,In_848);
nor U387 (N_387,In_646,In_905);
nand U388 (N_388,In_770,In_573);
nor U389 (N_389,In_576,In_935);
and U390 (N_390,In_951,In_34);
and U391 (N_391,In_79,In_671);
or U392 (N_392,In_33,In_718);
nor U393 (N_393,In_8,In_507);
nand U394 (N_394,In_352,In_832);
nand U395 (N_395,In_422,In_897);
or U396 (N_396,In_82,In_161);
xor U397 (N_397,In_954,In_88);
nor U398 (N_398,In_458,In_478);
or U399 (N_399,In_913,In_141);
xor U400 (N_400,In_781,In_672);
nor U401 (N_401,In_650,In_720);
nor U402 (N_402,In_305,In_590);
or U403 (N_403,In_506,In_329);
or U404 (N_404,In_917,In_962);
nand U405 (N_405,In_427,In_626);
nand U406 (N_406,In_944,In_623);
nor U407 (N_407,In_871,In_450);
nand U408 (N_408,In_633,In_107);
nand U409 (N_409,In_29,In_64);
xnor U410 (N_410,In_960,In_483);
nand U411 (N_411,In_629,In_527);
and U412 (N_412,In_651,In_692);
nor U413 (N_413,In_866,In_858);
nor U414 (N_414,In_964,In_525);
nand U415 (N_415,In_997,In_774);
xor U416 (N_416,In_572,In_389);
nor U417 (N_417,In_341,In_374);
nor U418 (N_418,In_783,In_78);
and U419 (N_419,In_979,In_200);
nand U420 (N_420,In_968,In_398);
nor U421 (N_421,In_698,In_644);
xnor U422 (N_422,In_247,In_881);
nor U423 (N_423,In_407,In_359);
and U424 (N_424,In_451,In_811);
nor U425 (N_425,In_236,In_62);
xor U426 (N_426,In_318,In_518);
nor U427 (N_427,In_567,In_263);
and U428 (N_428,In_228,In_985);
xnor U429 (N_429,In_117,In_891);
nor U430 (N_430,In_303,In_762);
nor U431 (N_431,In_610,In_35);
nor U432 (N_432,In_655,In_777);
nand U433 (N_433,In_184,In_160);
nor U434 (N_434,In_433,In_316);
nand U435 (N_435,In_240,In_72);
nor U436 (N_436,In_737,In_339);
or U437 (N_437,In_124,In_918);
nand U438 (N_438,In_201,In_306);
nor U439 (N_439,In_835,In_6);
nor U440 (N_440,In_403,In_992);
nor U441 (N_441,In_533,In_101);
nor U442 (N_442,In_118,In_500);
and U443 (N_443,In_439,In_766);
nand U444 (N_444,In_323,In_195);
and U445 (N_445,In_987,In_730);
and U446 (N_446,In_537,In_765);
nor U447 (N_447,In_710,In_48);
and U448 (N_448,In_39,In_108);
and U449 (N_449,In_416,In_138);
nand U450 (N_450,In_211,In_223);
or U451 (N_451,In_203,In_489);
nand U452 (N_452,In_255,In_224);
xor U453 (N_453,In_132,In_841);
and U454 (N_454,In_188,In_931);
and U455 (N_455,In_285,In_643);
nor U456 (N_456,In_826,In_970);
xnor U457 (N_457,In_975,In_495);
xnor U458 (N_458,In_522,In_393);
xor U459 (N_459,In_340,In_631);
nand U460 (N_460,In_387,In_752);
nor U461 (N_461,In_122,In_168);
xnor U462 (N_462,In_60,In_797);
nand U463 (N_463,In_517,In_767);
nor U464 (N_464,In_700,In_206);
nor U465 (N_465,In_230,In_491);
nor U466 (N_466,In_37,In_659);
nor U467 (N_467,In_582,In_534);
nand U468 (N_468,In_739,In_560);
nor U469 (N_469,In_65,In_509);
nand U470 (N_470,In_268,In_162);
or U471 (N_471,In_31,In_755);
nor U472 (N_472,In_322,In_778);
nand U473 (N_473,In_16,In_993);
nor U474 (N_474,In_410,In_526);
and U475 (N_475,In_84,In_297);
or U476 (N_476,In_148,In_257);
or U477 (N_477,In_356,In_249);
nor U478 (N_478,In_620,In_476);
nand U479 (N_479,In_197,In_226);
xnor U480 (N_480,In_472,In_790);
nand U481 (N_481,In_914,In_738);
or U482 (N_482,In_524,In_538);
xor U483 (N_483,In_614,In_208);
and U484 (N_484,In_639,In_508);
nand U485 (N_485,In_431,In_888);
or U486 (N_486,In_494,In_899);
or U487 (N_487,In_735,In_41);
nor U488 (N_488,In_173,In_641);
and U489 (N_489,In_896,In_253);
nand U490 (N_490,In_185,In_736);
nor U491 (N_491,In_414,In_119);
or U492 (N_492,In_575,In_786);
nor U493 (N_493,In_481,In_578);
or U494 (N_494,In_17,In_685);
nand U495 (N_495,In_991,In_312);
and U496 (N_496,In_87,In_349);
nor U497 (N_497,In_994,In_128);
or U498 (N_498,In_447,In_222);
or U499 (N_499,In_545,In_661);
nand U500 (N_500,In_63,In_494);
and U501 (N_501,In_23,In_411);
nand U502 (N_502,In_808,In_393);
nor U503 (N_503,In_454,In_355);
or U504 (N_504,In_922,In_246);
nand U505 (N_505,In_231,In_482);
xor U506 (N_506,In_482,In_86);
and U507 (N_507,In_603,In_994);
nand U508 (N_508,In_710,In_430);
and U509 (N_509,In_737,In_304);
nand U510 (N_510,In_406,In_30);
or U511 (N_511,In_899,In_880);
xor U512 (N_512,In_564,In_69);
nand U513 (N_513,In_424,In_419);
nand U514 (N_514,In_707,In_800);
nor U515 (N_515,In_401,In_483);
xnor U516 (N_516,In_897,In_791);
and U517 (N_517,In_971,In_402);
or U518 (N_518,In_143,In_514);
nand U519 (N_519,In_796,In_316);
or U520 (N_520,In_755,In_914);
or U521 (N_521,In_408,In_241);
or U522 (N_522,In_910,In_534);
or U523 (N_523,In_455,In_705);
nor U524 (N_524,In_978,In_315);
nor U525 (N_525,In_893,In_482);
or U526 (N_526,In_924,In_734);
xor U527 (N_527,In_683,In_407);
nand U528 (N_528,In_773,In_948);
or U529 (N_529,In_574,In_957);
nor U530 (N_530,In_160,In_270);
nand U531 (N_531,In_236,In_435);
xor U532 (N_532,In_96,In_288);
and U533 (N_533,In_692,In_956);
nand U534 (N_534,In_276,In_39);
and U535 (N_535,In_562,In_599);
and U536 (N_536,In_378,In_653);
nand U537 (N_537,In_538,In_509);
xnor U538 (N_538,In_807,In_903);
nor U539 (N_539,In_251,In_219);
nand U540 (N_540,In_268,In_109);
nor U541 (N_541,In_343,In_474);
nor U542 (N_542,In_887,In_385);
and U543 (N_543,In_932,In_286);
nand U544 (N_544,In_917,In_947);
xor U545 (N_545,In_126,In_462);
nor U546 (N_546,In_158,In_978);
xnor U547 (N_547,In_438,In_563);
nor U548 (N_548,In_825,In_894);
nand U549 (N_549,In_783,In_808);
or U550 (N_550,In_879,In_945);
nand U551 (N_551,In_269,In_150);
xnor U552 (N_552,In_810,In_137);
nand U553 (N_553,In_142,In_996);
nand U554 (N_554,In_227,In_925);
nor U555 (N_555,In_529,In_352);
or U556 (N_556,In_155,In_710);
or U557 (N_557,In_713,In_193);
or U558 (N_558,In_980,In_423);
or U559 (N_559,In_144,In_973);
nor U560 (N_560,In_767,In_264);
or U561 (N_561,In_714,In_197);
xor U562 (N_562,In_690,In_735);
nor U563 (N_563,In_182,In_39);
nor U564 (N_564,In_742,In_913);
nor U565 (N_565,In_845,In_372);
nor U566 (N_566,In_758,In_439);
nor U567 (N_567,In_255,In_46);
xnor U568 (N_568,In_811,In_559);
and U569 (N_569,In_196,In_882);
or U570 (N_570,In_407,In_513);
xor U571 (N_571,In_782,In_36);
xnor U572 (N_572,In_668,In_437);
or U573 (N_573,In_768,In_834);
nand U574 (N_574,In_878,In_130);
nor U575 (N_575,In_396,In_225);
or U576 (N_576,In_727,In_151);
nand U577 (N_577,In_849,In_129);
nand U578 (N_578,In_262,In_567);
and U579 (N_579,In_234,In_334);
nor U580 (N_580,In_929,In_106);
nor U581 (N_581,In_345,In_32);
and U582 (N_582,In_344,In_389);
nand U583 (N_583,In_850,In_855);
or U584 (N_584,In_130,In_442);
or U585 (N_585,In_931,In_315);
and U586 (N_586,In_144,In_987);
and U587 (N_587,In_925,In_649);
nand U588 (N_588,In_488,In_84);
or U589 (N_589,In_480,In_339);
nand U590 (N_590,In_983,In_206);
xnor U591 (N_591,In_87,In_748);
and U592 (N_592,In_329,In_57);
nand U593 (N_593,In_652,In_123);
nand U594 (N_594,In_145,In_593);
nand U595 (N_595,In_33,In_654);
or U596 (N_596,In_123,In_190);
nand U597 (N_597,In_343,In_228);
and U598 (N_598,In_527,In_265);
or U599 (N_599,In_686,In_795);
nand U600 (N_600,In_586,In_83);
and U601 (N_601,In_835,In_645);
nor U602 (N_602,In_282,In_531);
or U603 (N_603,In_765,In_619);
nand U604 (N_604,In_420,In_441);
and U605 (N_605,In_401,In_166);
and U606 (N_606,In_530,In_170);
nand U607 (N_607,In_177,In_983);
and U608 (N_608,In_243,In_830);
nor U609 (N_609,In_259,In_291);
or U610 (N_610,In_407,In_326);
nor U611 (N_611,In_807,In_299);
xor U612 (N_612,In_987,In_167);
or U613 (N_613,In_532,In_379);
or U614 (N_614,In_404,In_81);
or U615 (N_615,In_764,In_862);
nand U616 (N_616,In_747,In_661);
and U617 (N_617,In_805,In_37);
and U618 (N_618,In_954,In_207);
or U619 (N_619,In_626,In_237);
or U620 (N_620,In_769,In_115);
or U621 (N_621,In_65,In_483);
and U622 (N_622,In_133,In_583);
or U623 (N_623,In_692,In_7);
nor U624 (N_624,In_149,In_421);
and U625 (N_625,In_535,In_302);
nand U626 (N_626,In_981,In_949);
or U627 (N_627,In_942,In_414);
and U628 (N_628,In_516,In_152);
nor U629 (N_629,In_467,In_342);
nand U630 (N_630,In_47,In_786);
nand U631 (N_631,In_426,In_525);
xnor U632 (N_632,In_915,In_786);
and U633 (N_633,In_234,In_503);
and U634 (N_634,In_684,In_309);
nand U635 (N_635,In_195,In_34);
nor U636 (N_636,In_815,In_937);
nor U637 (N_637,In_237,In_227);
nor U638 (N_638,In_568,In_704);
or U639 (N_639,In_932,In_706);
nand U640 (N_640,In_355,In_485);
or U641 (N_641,In_477,In_383);
and U642 (N_642,In_929,In_189);
or U643 (N_643,In_355,In_611);
or U644 (N_644,In_461,In_517);
nand U645 (N_645,In_176,In_355);
nor U646 (N_646,In_750,In_98);
nand U647 (N_647,In_622,In_259);
nand U648 (N_648,In_212,In_985);
or U649 (N_649,In_697,In_55);
or U650 (N_650,In_31,In_642);
or U651 (N_651,In_330,In_962);
nor U652 (N_652,In_375,In_622);
or U653 (N_653,In_27,In_592);
nor U654 (N_654,In_385,In_305);
nor U655 (N_655,In_699,In_997);
and U656 (N_656,In_218,In_766);
and U657 (N_657,In_4,In_401);
and U658 (N_658,In_946,In_6);
and U659 (N_659,In_889,In_476);
nand U660 (N_660,In_84,In_230);
and U661 (N_661,In_971,In_611);
and U662 (N_662,In_384,In_806);
or U663 (N_663,In_684,In_178);
nor U664 (N_664,In_553,In_803);
nor U665 (N_665,In_363,In_813);
nor U666 (N_666,In_26,In_292);
nor U667 (N_667,In_527,In_216);
nand U668 (N_668,In_290,In_273);
nor U669 (N_669,In_496,In_842);
nor U670 (N_670,In_503,In_122);
xor U671 (N_671,In_243,In_122);
nand U672 (N_672,In_20,In_60);
and U673 (N_673,In_784,In_857);
or U674 (N_674,In_683,In_156);
nand U675 (N_675,In_507,In_924);
xnor U676 (N_676,In_407,In_857);
nand U677 (N_677,In_654,In_337);
or U678 (N_678,In_253,In_34);
nand U679 (N_679,In_41,In_130);
nand U680 (N_680,In_654,In_945);
nand U681 (N_681,In_42,In_667);
nand U682 (N_682,In_525,In_459);
xnor U683 (N_683,In_350,In_716);
nand U684 (N_684,In_732,In_433);
nor U685 (N_685,In_697,In_298);
nand U686 (N_686,In_258,In_589);
nand U687 (N_687,In_999,In_984);
or U688 (N_688,In_489,In_959);
nor U689 (N_689,In_452,In_172);
xor U690 (N_690,In_832,In_348);
nand U691 (N_691,In_364,In_221);
nand U692 (N_692,In_538,In_566);
or U693 (N_693,In_595,In_569);
and U694 (N_694,In_380,In_699);
and U695 (N_695,In_487,In_407);
nor U696 (N_696,In_806,In_267);
nor U697 (N_697,In_315,In_720);
nor U698 (N_698,In_825,In_63);
and U699 (N_699,In_430,In_718);
or U700 (N_700,In_894,In_775);
or U701 (N_701,In_76,In_706);
nand U702 (N_702,In_426,In_89);
nand U703 (N_703,In_988,In_138);
nand U704 (N_704,In_478,In_103);
nand U705 (N_705,In_280,In_173);
nand U706 (N_706,In_372,In_235);
xnor U707 (N_707,In_375,In_686);
and U708 (N_708,In_791,In_547);
and U709 (N_709,In_975,In_637);
or U710 (N_710,In_922,In_865);
and U711 (N_711,In_735,In_780);
nor U712 (N_712,In_671,In_695);
nand U713 (N_713,In_947,In_73);
or U714 (N_714,In_821,In_826);
and U715 (N_715,In_480,In_332);
and U716 (N_716,In_756,In_346);
and U717 (N_717,In_431,In_407);
and U718 (N_718,In_289,In_480);
nor U719 (N_719,In_784,In_245);
xor U720 (N_720,In_674,In_497);
nor U721 (N_721,In_684,In_227);
or U722 (N_722,In_321,In_653);
nor U723 (N_723,In_161,In_677);
nand U724 (N_724,In_83,In_121);
nand U725 (N_725,In_61,In_255);
and U726 (N_726,In_674,In_770);
nor U727 (N_727,In_462,In_773);
or U728 (N_728,In_767,In_366);
nand U729 (N_729,In_370,In_122);
and U730 (N_730,In_340,In_148);
or U731 (N_731,In_656,In_582);
nor U732 (N_732,In_371,In_984);
nand U733 (N_733,In_426,In_42);
nor U734 (N_734,In_871,In_354);
or U735 (N_735,In_474,In_23);
xor U736 (N_736,In_82,In_710);
nand U737 (N_737,In_975,In_871);
nor U738 (N_738,In_820,In_798);
and U739 (N_739,In_596,In_676);
xor U740 (N_740,In_792,In_286);
or U741 (N_741,In_905,In_569);
or U742 (N_742,In_764,In_564);
or U743 (N_743,In_639,In_174);
or U744 (N_744,In_958,In_686);
or U745 (N_745,In_207,In_467);
nand U746 (N_746,In_97,In_780);
or U747 (N_747,In_247,In_55);
or U748 (N_748,In_194,In_38);
and U749 (N_749,In_229,In_742);
and U750 (N_750,In_537,In_89);
or U751 (N_751,In_579,In_151);
nor U752 (N_752,In_463,In_761);
nor U753 (N_753,In_597,In_711);
nor U754 (N_754,In_915,In_26);
and U755 (N_755,In_943,In_617);
nand U756 (N_756,In_816,In_19);
nand U757 (N_757,In_782,In_831);
and U758 (N_758,In_227,In_949);
nand U759 (N_759,In_764,In_387);
nand U760 (N_760,In_267,In_714);
nand U761 (N_761,In_199,In_343);
and U762 (N_762,In_232,In_158);
nand U763 (N_763,In_346,In_674);
nor U764 (N_764,In_970,In_245);
or U765 (N_765,In_133,In_603);
or U766 (N_766,In_471,In_350);
nand U767 (N_767,In_779,In_460);
nand U768 (N_768,In_779,In_787);
and U769 (N_769,In_544,In_759);
or U770 (N_770,In_495,In_284);
nand U771 (N_771,In_601,In_323);
and U772 (N_772,In_719,In_446);
nand U773 (N_773,In_574,In_658);
nor U774 (N_774,In_927,In_317);
xor U775 (N_775,In_563,In_21);
and U776 (N_776,In_937,In_540);
nor U777 (N_777,In_700,In_816);
xnor U778 (N_778,In_585,In_113);
nor U779 (N_779,In_542,In_236);
or U780 (N_780,In_461,In_336);
or U781 (N_781,In_316,In_399);
and U782 (N_782,In_197,In_68);
nand U783 (N_783,In_979,In_978);
and U784 (N_784,In_756,In_535);
nor U785 (N_785,In_107,In_706);
nand U786 (N_786,In_806,In_898);
and U787 (N_787,In_650,In_284);
nor U788 (N_788,In_486,In_945);
and U789 (N_789,In_798,In_422);
and U790 (N_790,In_380,In_790);
or U791 (N_791,In_43,In_791);
and U792 (N_792,In_142,In_739);
and U793 (N_793,In_134,In_689);
nor U794 (N_794,In_519,In_52);
or U795 (N_795,In_332,In_508);
or U796 (N_796,In_776,In_364);
nand U797 (N_797,In_359,In_513);
nor U798 (N_798,In_768,In_553);
nand U799 (N_799,In_766,In_936);
or U800 (N_800,In_634,In_865);
or U801 (N_801,In_59,In_821);
nand U802 (N_802,In_596,In_632);
or U803 (N_803,In_550,In_317);
or U804 (N_804,In_80,In_237);
or U805 (N_805,In_142,In_349);
and U806 (N_806,In_822,In_805);
nand U807 (N_807,In_601,In_68);
nand U808 (N_808,In_455,In_732);
nor U809 (N_809,In_355,In_959);
and U810 (N_810,In_151,In_5);
nor U811 (N_811,In_219,In_284);
or U812 (N_812,In_99,In_951);
nor U813 (N_813,In_432,In_704);
xor U814 (N_814,In_725,In_829);
nand U815 (N_815,In_629,In_147);
and U816 (N_816,In_837,In_458);
nand U817 (N_817,In_56,In_537);
and U818 (N_818,In_524,In_726);
or U819 (N_819,In_813,In_756);
and U820 (N_820,In_954,In_878);
and U821 (N_821,In_288,In_222);
nor U822 (N_822,In_308,In_697);
and U823 (N_823,In_435,In_213);
xor U824 (N_824,In_905,In_158);
nand U825 (N_825,In_679,In_774);
xor U826 (N_826,In_552,In_888);
nand U827 (N_827,In_221,In_567);
and U828 (N_828,In_708,In_905);
xnor U829 (N_829,In_376,In_712);
and U830 (N_830,In_728,In_684);
nor U831 (N_831,In_442,In_737);
or U832 (N_832,In_19,In_225);
nor U833 (N_833,In_896,In_304);
nor U834 (N_834,In_803,In_27);
nand U835 (N_835,In_531,In_473);
nand U836 (N_836,In_88,In_633);
nand U837 (N_837,In_928,In_113);
nor U838 (N_838,In_657,In_962);
or U839 (N_839,In_759,In_556);
nand U840 (N_840,In_183,In_221);
nor U841 (N_841,In_183,In_279);
nand U842 (N_842,In_844,In_983);
and U843 (N_843,In_321,In_782);
nand U844 (N_844,In_798,In_893);
or U845 (N_845,In_364,In_632);
and U846 (N_846,In_550,In_377);
nor U847 (N_847,In_545,In_498);
or U848 (N_848,In_13,In_250);
nor U849 (N_849,In_50,In_311);
or U850 (N_850,In_680,In_22);
nor U851 (N_851,In_397,In_21);
or U852 (N_852,In_121,In_580);
or U853 (N_853,In_184,In_425);
xnor U854 (N_854,In_583,In_932);
and U855 (N_855,In_924,In_299);
nand U856 (N_856,In_28,In_323);
nor U857 (N_857,In_795,In_351);
or U858 (N_858,In_98,In_85);
or U859 (N_859,In_822,In_451);
nand U860 (N_860,In_289,In_32);
or U861 (N_861,In_861,In_874);
or U862 (N_862,In_964,In_284);
nor U863 (N_863,In_431,In_986);
and U864 (N_864,In_80,In_465);
and U865 (N_865,In_480,In_297);
or U866 (N_866,In_513,In_302);
and U867 (N_867,In_951,In_55);
nor U868 (N_868,In_435,In_45);
and U869 (N_869,In_738,In_868);
nand U870 (N_870,In_911,In_516);
nor U871 (N_871,In_29,In_583);
and U872 (N_872,In_101,In_950);
or U873 (N_873,In_467,In_5);
xor U874 (N_874,In_51,In_611);
nor U875 (N_875,In_854,In_15);
and U876 (N_876,In_7,In_659);
and U877 (N_877,In_836,In_363);
xor U878 (N_878,In_290,In_954);
nor U879 (N_879,In_715,In_99);
or U880 (N_880,In_714,In_90);
and U881 (N_881,In_162,In_751);
and U882 (N_882,In_864,In_575);
and U883 (N_883,In_894,In_782);
or U884 (N_884,In_804,In_644);
nor U885 (N_885,In_122,In_463);
nor U886 (N_886,In_505,In_688);
nor U887 (N_887,In_317,In_348);
or U888 (N_888,In_999,In_561);
and U889 (N_889,In_682,In_384);
nand U890 (N_890,In_529,In_990);
nor U891 (N_891,In_71,In_521);
or U892 (N_892,In_9,In_42);
and U893 (N_893,In_575,In_506);
nand U894 (N_894,In_841,In_657);
and U895 (N_895,In_757,In_490);
and U896 (N_896,In_796,In_667);
nor U897 (N_897,In_915,In_902);
xnor U898 (N_898,In_745,In_479);
nor U899 (N_899,In_985,In_159);
and U900 (N_900,In_405,In_933);
xor U901 (N_901,In_546,In_232);
xor U902 (N_902,In_169,In_990);
nand U903 (N_903,In_951,In_272);
nor U904 (N_904,In_635,In_908);
or U905 (N_905,In_255,In_830);
xnor U906 (N_906,In_177,In_718);
nand U907 (N_907,In_510,In_743);
nand U908 (N_908,In_255,In_340);
xor U909 (N_909,In_351,In_589);
nor U910 (N_910,In_325,In_181);
nand U911 (N_911,In_794,In_90);
and U912 (N_912,In_493,In_393);
and U913 (N_913,In_950,In_526);
nor U914 (N_914,In_836,In_151);
or U915 (N_915,In_63,In_869);
nor U916 (N_916,In_347,In_387);
and U917 (N_917,In_694,In_157);
nor U918 (N_918,In_477,In_81);
nor U919 (N_919,In_85,In_526);
and U920 (N_920,In_919,In_628);
or U921 (N_921,In_981,In_80);
xor U922 (N_922,In_527,In_156);
or U923 (N_923,In_567,In_697);
nor U924 (N_924,In_563,In_464);
and U925 (N_925,In_582,In_216);
nand U926 (N_926,In_812,In_804);
or U927 (N_927,In_607,In_659);
nor U928 (N_928,In_215,In_607);
and U929 (N_929,In_284,In_430);
nor U930 (N_930,In_230,In_605);
and U931 (N_931,In_963,In_896);
or U932 (N_932,In_280,In_8);
or U933 (N_933,In_268,In_247);
or U934 (N_934,In_868,In_962);
nor U935 (N_935,In_165,In_588);
or U936 (N_936,In_897,In_420);
nand U937 (N_937,In_996,In_238);
nand U938 (N_938,In_836,In_519);
nor U939 (N_939,In_400,In_680);
or U940 (N_940,In_822,In_3);
and U941 (N_941,In_783,In_528);
nor U942 (N_942,In_205,In_873);
nand U943 (N_943,In_186,In_273);
and U944 (N_944,In_750,In_55);
nor U945 (N_945,In_624,In_935);
nand U946 (N_946,In_203,In_793);
nand U947 (N_947,In_206,In_101);
or U948 (N_948,In_83,In_733);
nand U949 (N_949,In_298,In_165);
nand U950 (N_950,In_949,In_344);
nand U951 (N_951,In_644,In_860);
xor U952 (N_952,In_185,In_64);
xor U953 (N_953,In_968,In_857);
nand U954 (N_954,In_330,In_188);
nand U955 (N_955,In_329,In_581);
and U956 (N_956,In_574,In_505);
nor U957 (N_957,In_142,In_629);
or U958 (N_958,In_997,In_230);
nor U959 (N_959,In_254,In_285);
nand U960 (N_960,In_316,In_552);
and U961 (N_961,In_450,In_514);
xor U962 (N_962,In_998,In_561);
nand U963 (N_963,In_158,In_471);
nor U964 (N_964,In_333,In_254);
or U965 (N_965,In_875,In_244);
nor U966 (N_966,In_989,In_704);
and U967 (N_967,In_614,In_247);
nor U968 (N_968,In_890,In_559);
nand U969 (N_969,In_308,In_482);
nor U970 (N_970,In_312,In_514);
xor U971 (N_971,In_551,In_4);
xnor U972 (N_972,In_602,In_28);
nor U973 (N_973,In_655,In_379);
nand U974 (N_974,In_979,In_920);
nor U975 (N_975,In_437,In_944);
and U976 (N_976,In_317,In_968);
or U977 (N_977,In_109,In_954);
and U978 (N_978,In_945,In_437);
and U979 (N_979,In_319,In_780);
nand U980 (N_980,In_718,In_728);
xnor U981 (N_981,In_291,In_813);
and U982 (N_982,In_484,In_107);
and U983 (N_983,In_247,In_611);
nand U984 (N_984,In_690,In_507);
and U985 (N_985,In_435,In_697);
nor U986 (N_986,In_615,In_356);
nand U987 (N_987,In_182,In_339);
or U988 (N_988,In_108,In_247);
nand U989 (N_989,In_422,In_88);
or U990 (N_990,In_449,In_321);
nor U991 (N_991,In_908,In_711);
xnor U992 (N_992,In_819,In_215);
nand U993 (N_993,In_758,In_559);
or U994 (N_994,In_185,In_779);
nand U995 (N_995,In_787,In_37);
xor U996 (N_996,In_903,In_337);
and U997 (N_997,In_552,In_456);
and U998 (N_998,In_491,In_69);
nand U999 (N_999,In_893,In_757);
and U1000 (N_1000,In_173,In_492);
nand U1001 (N_1001,In_302,In_464);
nor U1002 (N_1002,In_820,In_271);
or U1003 (N_1003,In_412,In_558);
or U1004 (N_1004,In_614,In_17);
and U1005 (N_1005,In_757,In_801);
and U1006 (N_1006,In_223,In_159);
nand U1007 (N_1007,In_655,In_250);
or U1008 (N_1008,In_359,In_821);
nor U1009 (N_1009,In_379,In_435);
nor U1010 (N_1010,In_839,In_332);
nor U1011 (N_1011,In_778,In_463);
nor U1012 (N_1012,In_312,In_526);
nand U1013 (N_1013,In_215,In_527);
xor U1014 (N_1014,In_969,In_35);
or U1015 (N_1015,In_742,In_793);
or U1016 (N_1016,In_534,In_331);
xor U1017 (N_1017,In_595,In_942);
or U1018 (N_1018,In_36,In_309);
or U1019 (N_1019,In_375,In_495);
nor U1020 (N_1020,In_995,In_690);
nand U1021 (N_1021,In_876,In_472);
or U1022 (N_1022,In_101,In_471);
and U1023 (N_1023,In_988,In_171);
and U1024 (N_1024,In_670,In_256);
and U1025 (N_1025,In_289,In_912);
nand U1026 (N_1026,In_812,In_367);
or U1027 (N_1027,In_620,In_731);
or U1028 (N_1028,In_159,In_79);
or U1029 (N_1029,In_34,In_885);
nand U1030 (N_1030,In_290,In_19);
and U1031 (N_1031,In_900,In_297);
nor U1032 (N_1032,In_811,In_970);
nand U1033 (N_1033,In_640,In_807);
nor U1034 (N_1034,In_430,In_218);
and U1035 (N_1035,In_857,In_310);
nor U1036 (N_1036,In_826,In_477);
or U1037 (N_1037,In_965,In_978);
nand U1038 (N_1038,In_934,In_543);
nand U1039 (N_1039,In_704,In_68);
nor U1040 (N_1040,In_694,In_360);
and U1041 (N_1041,In_305,In_587);
or U1042 (N_1042,In_994,In_850);
nand U1043 (N_1043,In_534,In_176);
nor U1044 (N_1044,In_700,In_119);
and U1045 (N_1045,In_989,In_548);
and U1046 (N_1046,In_180,In_961);
nand U1047 (N_1047,In_736,In_27);
nor U1048 (N_1048,In_645,In_217);
nand U1049 (N_1049,In_601,In_41);
or U1050 (N_1050,In_708,In_864);
nor U1051 (N_1051,In_236,In_589);
and U1052 (N_1052,In_436,In_892);
nand U1053 (N_1053,In_563,In_99);
or U1054 (N_1054,In_655,In_483);
nand U1055 (N_1055,In_42,In_299);
nor U1056 (N_1056,In_711,In_263);
and U1057 (N_1057,In_68,In_162);
nand U1058 (N_1058,In_699,In_89);
nand U1059 (N_1059,In_492,In_28);
or U1060 (N_1060,In_830,In_709);
and U1061 (N_1061,In_817,In_269);
or U1062 (N_1062,In_944,In_805);
nand U1063 (N_1063,In_365,In_452);
nand U1064 (N_1064,In_651,In_795);
nor U1065 (N_1065,In_689,In_188);
xnor U1066 (N_1066,In_82,In_312);
nand U1067 (N_1067,In_474,In_720);
or U1068 (N_1068,In_727,In_469);
nor U1069 (N_1069,In_908,In_871);
or U1070 (N_1070,In_334,In_725);
or U1071 (N_1071,In_468,In_897);
nor U1072 (N_1072,In_804,In_231);
or U1073 (N_1073,In_981,In_450);
nand U1074 (N_1074,In_674,In_955);
nor U1075 (N_1075,In_810,In_190);
or U1076 (N_1076,In_948,In_792);
nor U1077 (N_1077,In_811,In_935);
xor U1078 (N_1078,In_272,In_251);
or U1079 (N_1079,In_573,In_705);
nand U1080 (N_1080,In_268,In_726);
or U1081 (N_1081,In_610,In_427);
nand U1082 (N_1082,In_83,In_11);
and U1083 (N_1083,In_59,In_233);
or U1084 (N_1084,In_516,In_150);
nor U1085 (N_1085,In_537,In_126);
and U1086 (N_1086,In_417,In_622);
nand U1087 (N_1087,In_442,In_755);
or U1088 (N_1088,In_185,In_708);
or U1089 (N_1089,In_509,In_118);
and U1090 (N_1090,In_709,In_247);
xor U1091 (N_1091,In_305,In_536);
and U1092 (N_1092,In_785,In_267);
and U1093 (N_1093,In_781,In_60);
or U1094 (N_1094,In_446,In_892);
xor U1095 (N_1095,In_578,In_814);
and U1096 (N_1096,In_696,In_220);
nor U1097 (N_1097,In_685,In_675);
or U1098 (N_1098,In_732,In_93);
nand U1099 (N_1099,In_189,In_179);
nor U1100 (N_1100,In_232,In_56);
and U1101 (N_1101,In_633,In_76);
xor U1102 (N_1102,In_50,In_739);
and U1103 (N_1103,In_917,In_59);
nor U1104 (N_1104,In_795,In_558);
xnor U1105 (N_1105,In_284,In_464);
nand U1106 (N_1106,In_771,In_637);
nor U1107 (N_1107,In_152,In_958);
and U1108 (N_1108,In_28,In_665);
nand U1109 (N_1109,In_16,In_581);
or U1110 (N_1110,In_799,In_932);
nand U1111 (N_1111,In_428,In_882);
or U1112 (N_1112,In_856,In_133);
or U1113 (N_1113,In_531,In_745);
nor U1114 (N_1114,In_69,In_837);
or U1115 (N_1115,In_725,In_872);
or U1116 (N_1116,In_21,In_371);
and U1117 (N_1117,In_931,In_293);
nand U1118 (N_1118,In_542,In_624);
nor U1119 (N_1119,In_503,In_112);
nor U1120 (N_1120,In_348,In_840);
xor U1121 (N_1121,In_808,In_76);
and U1122 (N_1122,In_393,In_626);
xor U1123 (N_1123,In_563,In_51);
nor U1124 (N_1124,In_109,In_856);
or U1125 (N_1125,In_318,In_363);
nand U1126 (N_1126,In_692,In_115);
or U1127 (N_1127,In_884,In_440);
nand U1128 (N_1128,In_691,In_503);
or U1129 (N_1129,In_837,In_184);
or U1130 (N_1130,In_560,In_643);
and U1131 (N_1131,In_630,In_267);
xnor U1132 (N_1132,In_574,In_522);
nor U1133 (N_1133,In_408,In_103);
or U1134 (N_1134,In_81,In_218);
nor U1135 (N_1135,In_373,In_288);
nor U1136 (N_1136,In_122,In_244);
nand U1137 (N_1137,In_873,In_55);
nand U1138 (N_1138,In_217,In_757);
nand U1139 (N_1139,In_814,In_310);
or U1140 (N_1140,In_81,In_949);
or U1141 (N_1141,In_793,In_171);
nand U1142 (N_1142,In_531,In_854);
nor U1143 (N_1143,In_917,In_494);
nor U1144 (N_1144,In_560,In_71);
xor U1145 (N_1145,In_881,In_753);
and U1146 (N_1146,In_317,In_562);
nand U1147 (N_1147,In_908,In_589);
or U1148 (N_1148,In_103,In_729);
and U1149 (N_1149,In_596,In_513);
nand U1150 (N_1150,In_95,In_81);
xnor U1151 (N_1151,In_793,In_695);
and U1152 (N_1152,In_928,In_658);
nor U1153 (N_1153,In_809,In_649);
nor U1154 (N_1154,In_208,In_889);
nor U1155 (N_1155,In_110,In_405);
nand U1156 (N_1156,In_562,In_924);
and U1157 (N_1157,In_86,In_952);
xnor U1158 (N_1158,In_403,In_551);
and U1159 (N_1159,In_562,In_512);
nor U1160 (N_1160,In_21,In_583);
and U1161 (N_1161,In_43,In_787);
nor U1162 (N_1162,In_976,In_868);
nand U1163 (N_1163,In_368,In_912);
xnor U1164 (N_1164,In_478,In_351);
nand U1165 (N_1165,In_734,In_483);
and U1166 (N_1166,In_567,In_351);
nor U1167 (N_1167,In_634,In_983);
or U1168 (N_1168,In_271,In_601);
or U1169 (N_1169,In_24,In_480);
or U1170 (N_1170,In_788,In_203);
or U1171 (N_1171,In_12,In_402);
or U1172 (N_1172,In_71,In_5);
or U1173 (N_1173,In_239,In_600);
or U1174 (N_1174,In_673,In_270);
nor U1175 (N_1175,In_1,In_184);
nor U1176 (N_1176,In_992,In_27);
nand U1177 (N_1177,In_540,In_63);
or U1178 (N_1178,In_803,In_918);
nand U1179 (N_1179,In_290,In_749);
or U1180 (N_1180,In_355,In_503);
xnor U1181 (N_1181,In_9,In_898);
nand U1182 (N_1182,In_853,In_224);
or U1183 (N_1183,In_948,In_277);
nand U1184 (N_1184,In_911,In_134);
nor U1185 (N_1185,In_174,In_661);
nand U1186 (N_1186,In_605,In_631);
or U1187 (N_1187,In_865,In_556);
nor U1188 (N_1188,In_184,In_886);
nand U1189 (N_1189,In_3,In_498);
nor U1190 (N_1190,In_630,In_273);
or U1191 (N_1191,In_863,In_930);
nand U1192 (N_1192,In_669,In_818);
or U1193 (N_1193,In_544,In_462);
nor U1194 (N_1194,In_442,In_89);
nand U1195 (N_1195,In_418,In_982);
nor U1196 (N_1196,In_784,In_763);
nor U1197 (N_1197,In_847,In_635);
nor U1198 (N_1198,In_928,In_36);
xor U1199 (N_1199,In_308,In_679);
nand U1200 (N_1200,In_987,In_352);
nand U1201 (N_1201,In_404,In_591);
nor U1202 (N_1202,In_17,In_506);
nor U1203 (N_1203,In_753,In_899);
and U1204 (N_1204,In_399,In_144);
nor U1205 (N_1205,In_84,In_491);
or U1206 (N_1206,In_885,In_927);
and U1207 (N_1207,In_754,In_258);
and U1208 (N_1208,In_720,In_376);
nand U1209 (N_1209,In_389,In_232);
nand U1210 (N_1210,In_865,In_623);
nand U1211 (N_1211,In_325,In_787);
or U1212 (N_1212,In_441,In_617);
and U1213 (N_1213,In_646,In_109);
or U1214 (N_1214,In_512,In_709);
nor U1215 (N_1215,In_174,In_744);
xnor U1216 (N_1216,In_139,In_333);
and U1217 (N_1217,In_414,In_777);
nor U1218 (N_1218,In_517,In_410);
and U1219 (N_1219,In_588,In_956);
nand U1220 (N_1220,In_653,In_760);
nand U1221 (N_1221,In_85,In_474);
or U1222 (N_1222,In_572,In_375);
and U1223 (N_1223,In_501,In_993);
and U1224 (N_1224,In_82,In_491);
and U1225 (N_1225,In_543,In_883);
and U1226 (N_1226,In_587,In_498);
or U1227 (N_1227,In_822,In_894);
or U1228 (N_1228,In_446,In_307);
nand U1229 (N_1229,In_965,In_165);
or U1230 (N_1230,In_274,In_153);
nand U1231 (N_1231,In_275,In_196);
xnor U1232 (N_1232,In_386,In_831);
or U1233 (N_1233,In_216,In_102);
or U1234 (N_1234,In_448,In_501);
xor U1235 (N_1235,In_182,In_930);
or U1236 (N_1236,In_574,In_837);
or U1237 (N_1237,In_249,In_422);
or U1238 (N_1238,In_497,In_212);
nor U1239 (N_1239,In_764,In_574);
and U1240 (N_1240,In_934,In_876);
or U1241 (N_1241,In_534,In_700);
and U1242 (N_1242,In_139,In_193);
nor U1243 (N_1243,In_8,In_632);
or U1244 (N_1244,In_103,In_564);
nor U1245 (N_1245,In_764,In_38);
nor U1246 (N_1246,In_279,In_84);
nor U1247 (N_1247,In_512,In_650);
and U1248 (N_1248,In_441,In_207);
nor U1249 (N_1249,In_688,In_226);
or U1250 (N_1250,In_894,In_409);
nor U1251 (N_1251,In_52,In_280);
or U1252 (N_1252,In_652,In_802);
and U1253 (N_1253,In_925,In_726);
or U1254 (N_1254,In_283,In_261);
nor U1255 (N_1255,In_195,In_408);
and U1256 (N_1256,In_832,In_531);
and U1257 (N_1257,In_844,In_93);
and U1258 (N_1258,In_6,In_971);
or U1259 (N_1259,In_435,In_810);
and U1260 (N_1260,In_291,In_469);
or U1261 (N_1261,In_248,In_776);
and U1262 (N_1262,In_741,In_773);
xor U1263 (N_1263,In_322,In_443);
nor U1264 (N_1264,In_48,In_66);
nor U1265 (N_1265,In_61,In_532);
or U1266 (N_1266,In_920,In_714);
nor U1267 (N_1267,In_429,In_254);
or U1268 (N_1268,In_817,In_683);
nand U1269 (N_1269,In_168,In_622);
or U1270 (N_1270,In_458,In_705);
nor U1271 (N_1271,In_486,In_460);
nor U1272 (N_1272,In_785,In_874);
xnor U1273 (N_1273,In_273,In_468);
nand U1274 (N_1274,In_656,In_921);
or U1275 (N_1275,In_962,In_894);
nor U1276 (N_1276,In_522,In_960);
or U1277 (N_1277,In_710,In_915);
xor U1278 (N_1278,In_48,In_492);
nand U1279 (N_1279,In_19,In_467);
nand U1280 (N_1280,In_555,In_42);
and U1281 (N_1281,In_16,In_690);
or U1282 (N_1282,In_475,In_420);
or U1283 (N_1283,In_670,In_647);
nor U1284 (N_1284,In_996,In_691);
or U1285 (N_1285,In_967,In_590);
nand U1286 (N_1286,In_894,In_353);
nand U1287 (N_1287,In_126,In_746);
and U1288 (N_1288,In_680,In_493);
nor U1289 (N_1289,In_714,In_516);
nand U1290 (N_1290,In_97,In_169);
nand U1291 (N_1291,In_241,In_532);
nand U1292 (N_1292,In_313,In_945);
and U1293 (N_1293,In_730,In_504);
and U1294 (N_1294,In_589,In_724);
nor U1295 (N_1295,In_158,In_372);
nor U1296 (N_1296,In_515,In_304);
and U1297 (N_1297,In_961,In_283);
or U1298 (N_1298,In_558,In_503);
nand U1299 (N_1299,In_799,In_582);
nand U1300 (N_1300,In_285,In_147);
nand U1301 (N_1301,In_322,In_620);
and U1302 (N_1302,In_409,In_955);
nand U1303 (N_1303,In_261,In_490);
nor U1304 (N_1304,In_572,In_346);
nand U1305 (N_1305,In_501,In_710);
xor U1306 (N_1306,In_533,In_169);
and U1307 (N_1307,In_88,In_196);
nor U1308 (N_1308,In_144,In_44);
xnor U1309 (N_1309,In_509,In_622);
nand U1310 (N_1310,In_269,In_37);
nor U1311 (N_1311,In_334,In_690);
and U1312 (N_1312,In_494,In_49);
nor U1313 (N_1313,In_506,In_569);
or U1314 (N_1314,In_17,In_476);
or U1315 (N_1315,In_61,In_780);
nor U1316 (N_1316,In_853,In_622);
nor U1317 (N_1317,In_67,In_101);
or U1318 (N_1318,In_365,In_723);
xor U1319 (N_1319,In_558,In_798);
and U1320 (N_1320,In_627,In_247);
or U1321 (N_1321,In_829,In_37);
or U1322 (N_1322,In_130,In_571);
and U1323 (N_1323,In_664,In_538);
or U1324 (N_1324,In_176,In_418);
and U1325 (N_1325,In_637,In_638);
or U1326 (N_1326,In_679,In_950);
nand U1327 (N_1327,In_180,In_637);
nand U1328 (N_1328,In_546,In_921);
and U1329 (N_1329,In_397,In_391);
and U1330 (N_1330,In_981,In_386);
xor U1331 (N_1331,In_760,In_322);
or U1332 (N_1332,In_537,In_42);
nand U1333 (N_1333,In_960,In_154);
nor U1334 (N_1334,In_396,In_751);
nor U1335 (N_1335,In_93,In_497);
or U1336 (N_1336,In_828,In_269);
nand U1337 (N_1337,In_84,In_95);
nor U1338 (N_1338,In_110,In_917);
nor U1339 (N_1339,In_625,In_138);
or U1340 (N_1340,In_423,In_788);
nand U1341 (N_1341,In_338,In_399);
nor U1342 (N_1342,In_981,In_993);
nor U1343 (N_1343,In_161,In_21);
nand U1344 (N_1344,In_605,In_271);
xor U1345 (N_1345,In_795,In_298);
nand U1346 (N_1346,In_563,In_663);
nor U1347 (N_1347,In_73,In_222);
nor U1348 (N_1348,In_528,In_766);
or U1349 (N_1349,In_11,In_764);
xor U1350 (N_1350,In_300,In_457);
or U1351 (N_1351,In_5,In_0);
nor U1352 (N_1352,In_991,In_91);
and U1353 (N_1353,In_86,In_252);
and U1354 (N_1354,In_448,In_386);
nor U1355 (N_1355,In_298,In_662);
or U1356 (N_1356,In_481,In_417);
nor U1357 (N_1357,In_252,In_140);
xor U1358 (N_1358,In_716,In_491);
nor U1359 (N_1359,In_318,In_761);
xnor U1360 (N_1360,In_869,In_873);
or U1361 (N_1361,In_792,In_79);
nor U1362 (N_1362,In_48,In_620);
nor U1363 (N_1363,In_5,In_516);
or U1364 (N_1364,In_596,In_378);
or U1365 (N_1365,In_677,In_943);
nand U1366 (N_1366,In_7,In_785);
nand U1367 (N_1367,In_155,In_604);
nor U1368 (N_1368,In_995,In_45);
nand U1369 (N_1369,In_498,In_165);
nand U1370 (N_1370,In_777,In_860);
or U1371 (N_1371,In_608,In_474);
nor U1372 (N_1372,In_437,In_279);
nor U1373 (N_1373,In_696,In_830);
nor U1374 (N_1374,In_504,In_32);
xor U1375 (N_1375,In_309,In_11);
or U1376 (N_1376,In_950,In_479);
xnor U1377 (N_1377,In_851,In_471);
and U1378 (N_1378,In_448,In_32);
nor U1379 (N_1379,In_422,In_13);
or U1380 (N_1380,In_182,In_640);
nand U1381 (N_1381,In_533,In_641);
nand U1382 (N_1382,In_783,In_229);
nor U1383 (N_1383,In_911,In_384);
or U1384 (N_1384,In_84,In_105);
or U1385 (N_1385,In_928,In_552);
xnor U1386 (N_1386,In_567,In_953);
nor U1387 (N_1387,In_719,In_892);
nand U1388 (N_1388,In_477,In_864);
xor U1389 (N_1389,In_490,In_433);
nor U1390 (N_1390,In_84,In_971);
nand U1391 (N_1391,In_848,In_781);
nand U1392 (N_1392,In_209,In_653);
and U1393 (N_1393,In_746,In_63);
and U1394 (N_1394,In_304,In_838);
nor U1395 (N_1395,In_775,In_146);
nand U1396 (N_1396,In_117,In_713);
nand U1397 (N_1397,In_820,In_536);
nand U1398 (N_1398,In_558,In_308);
nand U1399 (N_1399,In_765,In_213);
or U1400 (N_1400,In_658,In_480);
xor U1401 (N_1401,In_445,In_794);
or U1402 (N_1402,In_230,In_337);
nand U1403 (N_1403,In_555,In_936);
nor U1404 (N_1404,In_470,In_737);
xnor U1405 (N_1405,In_454,In_907);
nand U1406 (N_1406,In_725,In_904);
or U1407 (N_1407,In_55,In_25);
or U1408 (N_1408,In_299,In_902);
nor U1409 (N_1409,In_672,In_408);
and U1410 (N_1410,In_816,In_715);
xor U1411 (N_1411,In_252,In_262);
or U1412 (N_1412,In_923,In_162);
and U1413 (N_1413,In_951,In_768);
or U1414 (N_1414,In_589,In_118);
nand U1415 (N_1415,In_395,In_642);
or U1416 (N_1416,In_687,In_831);
and U1417 (N_1417,In_431,In_398);
nand U1418 (N_1418,In_132,In_109);
nand U1419 (N_1419,In_156,In_895);
nor U1420 (N_1420,In_327,In_301);
or U1421 (N_1421,In_33,In_371);
and U1422 (N_1422,In_988,In_319);
xor U1423 (N_1423,In_844,In_536);
nor U1424 (N_1424,In_662,In_959);
and U1425 (N_1425,In_962,In_92);
nand U1426 (N_1426,In_513,In_881);
xor U1427 (N_1427,In_301,In_431);
nand U1428 (N_1428,In_366,In_264);
nor U1429 (N_1429,In_827,In_454);
nand U1430 (N_1430,In_49,In_675);
or U1431 (N_1431,In_37,In_23);
nand U1432 (N_1432,In_691,In_719);
nor U1433 (N_1433,In_283,In_194);
nand U1434 (N_1434,In_594,In_11);
and U1435 (N_1435,In_79,In_626);
nor U1436 (N_1436,In_571,In_68);
and U1437 (N_1437,In_1,In_954);
or U1438 (N_1438,In_990,In_281);
nand U1439 (N_1439,In_161,In_496);
and U1440 (N_1440,In_762,In_43);
nor U1441 (N_1441,In_298,In_718);
nor U1442 (N_1442,In_88,In_396);
nor U1443 (N_1443,In_919,In_716);
and U1444 (N_1444,In_981,In_331);
and U1445 (N_1445,In_414,In_176);
or U1446 (N_1446,In_373,In_762);
and U1447 (N_1447,In_540,In_533);
nor U1448 (N_1448,In_295,In_552);
or U1449 (N_1449,In_387,In_528);
and U1450 (N_1450,In_687,In_359);
or U1451 (N_1451,In_725,In_117);
and U1452 (N_1452,In_236,In_134);
or U1453 (N_1453,In_43,In_963);
xnor U1454 (N_1454,In_962,In_286);
nor U1455 (N_1455,In_777,In_301);
or U1456 (N_1456,In_269,In_49);
nand U1457 (N_1457,In_469,In_966);
nand U1458 (N_1458,In_439,In_805);
nand U1459 (N_1459,In_478,In_26);
and U1460 (N_1460,In_148,In_780);
nor U1461 (N_1461,In_653,In_119);
and U1462 (N_1462,In_680,In_639);
and U1463 (N_1463,In_93,In_711);
and U1464 (N_1464,In_279,In_775);
nor U1465 (N_1465,In_898,In_504);
or U1466 (N_1466,In_852,In_796);
nand U1467 (N_1467,In_563,In_751);
xnor U1468 (N_1468,In_75,In_489);
and U1469 (N_1469,In_368,In_726);
nor U1470 (N_1470,In_280,In_53);
nand U1471 (N_1471,In_230,In_931);
xor U1472 (N_1472,In_351,In_396);
and U1473 (N_1473,In_829,In_248);
or U1474 (N_1474,In_129,In_177);
or U1475 (N_1475,In_599,In_584);
or U1476 (N_1476,In_7,In_448);
nor U1477 (N_1477,In_210,In_620);
or U1478 (N_1478,In_51,In_986);
and U1479 (N_1479,In_689,In_58);
nor U1480 (N_1480,In_702,In_446);
or U1481 (N_1481,In_776,In_641);
xor U1482 (N_1482,In_95,In_513);
and U1483 (N_1483,In_531,In_875);
or U1484 (N_1484,In_296,In_430);
nand U1485 (N_1485,In_265,In_504);
and U1486 (N_1486,In_678,In_968);
and U1487 (N_1487,In_472,In_46);
or U1488 (N_1488,In_265,In_123);
nand U1489 (N_1489,In_437,In_37);
or U1490 (N_1490,In_421,In_170);
nand U1491 (N_1491,In_125,In_569);
or U1492 (N_1492,In_567,In_639);
nor U1493 (N_1493,In_862,In_469);
nor U1494 (N_1494,In_459,In_880);
nor U1495 (N_1495,In_624,In_718);
or U1496 (N_1496,In_248,In_957);
nand U1497 (N_1497,In_920,In_932);
and U1498 (N_1498,In_383,In_348);
nand U1499 (N_1499,In_901,In_823);
nor U1500 (N_1500,In_392,In_425);
xnor U1501 (N_1501,In_122,In_711);
nor U1502 (N_1502,In_150,In_943);
xnor U1503 (N_1503,In_820,In_30);
xor U1504 (N_1504,In_462,In_124);
and U1505 (N_1505,In_324,In_854);
xnor U1506 (N_1506,In_981,In_998);
nor U1507 (N_1507,In_903,In_847);
and U1508 (N_1508,In_542,In_56);
nor U1509 (N_1509,In_594,In_572);
and U1510 (N_1510,In_339,In_72);
nand U1511 (N_1511,In_974,In_550);
and U1512 (N_1512,In_197,In_805);
nor U1513 (N_1513,In_754,In_950);
nand U1514 (N_1514,In_540,In_258);
nor U1515 (N_1515,In_906,In_565);
nor U1516 (N_1516,In_992,In_874);
nand U1517 (N_1517,In_31,In_908);
and U1518 (N_1518,In_117,In_948);
or U1519 (N_1519,In_626,In_395);
nand U1520 (N_1520,In_97,In_183);
and U1521 (N_1521,In_920,In_30);
nor U1522 (N_1522,In_83,In_159);
nand U1523 (N_1523,In_869,In_446);
and U1524 (N_1524,In_688,In_673);
nand U1525 (N_1525,In_769,In_256);
and U1526 (N_1526,In_913,In_968);
and U1527 (N_1527,In_809,In_209);
nand U1528 (N_1528,In_166,In_771);
nand U1529 (N_1529,In_948,In_227);
xor U1530 (N_1530,In_537,In_152);
or U1531 (N_1531,In_338,In_482);
nand U1532 (N_1532,In_737,In_124);
and U1533 (N_1533,In_555,In_544);
or U1534 (N_1534,In_875,In_722);
xnor U1535 (N_1535,In_38,In_894);
nor U1536 (N_1536,In_552,In_723);
and U1537 (N_1537,In_891,In_887);
xnor U1538 (N_1538,In_404,In_575);
xnor U1539 (N_1539,In_246,In_681);
nor U1540 (N_1540,In_81,In_898);
nand U1541 (N_1541,In_477,In_445);
and U1542 (N_1542,In_367,In_859);
nor U1543 (N_1543,In_398,In_392);
nor U1544 (N_1544,In_171,In_64);
and U1545 (N_1545,In_311,In_948);
nand U1546 (N_1546,In_463,In_315);
and U1547 (N_1547,In_231,In_458);
and U1548 (N_1548,In_937,In_26);
or U1549 (N_1549,In_586,In_364);
and U1550 (N_1550,In_601,In_695);
and U1551 (N_1551,In_262,In_605);
nand U1552 (N_1552,In_885,In_655);
or U1553 (N_1553,In_639,In_734);
nand U1554 (N_1554,In_451,In_653);
xor U1555 (N_1555,In_709,In_524);
nand U1556 (N_1556,In_148,In_574);
nor U1557 (N_1557,In_817,In_705);
or U1558 (N_1558,In_205,In_356);
and U1559 (N_1559,In_373,In_1);
or U1560 (N_1560,In_875,In_507);
or U1561 (N_1561,In_193,In_437);
nand U1562 (N_1562,In_747,In_154);
nor U1563 (N_1563,In_545,In_695);
nand U1564 (N_1564,In_769,In_929);
or U1565 (N_1565,In_319,In_869);
or U1566 (N_1566,In_901,In_936);
nand U1567 (N_1567,In_975,In_541);
nor U1568 (N_1568,In_451,In_192);
and U1569 (N_1569,In_268,In_517);
nor U1570 (N_1570,In_78,In_541);
nand U1571 (N_1571,In_179,In_218);
xnor U1572 (N_1572,In_282,In_69);
and U1573 (N_1573,In_874,In_72);
or U1574 (N_1574,In_850,In_425);
and U1575 (N_1575,In_615,In_96);
and U1576 (N_1576,In_521,In_167);
and U1577 (N_1577,In_869,In_376);
and U1578 (N_1578,In_753,In_202);
nand U1579 (N_1579,In_108,In_444);
nor U1580 (N_1580,In_546,In_747);
and U1581 (N_1581,In_915,In_883);
or U1582 (N_1582,In_614,In_130);
and U1583 (N_1583,In_577,In_284);
and U1584 (N_1584,In_48,In_378);
and U1585 (N_1585,In_959,In_89);
nand U1586 (N_1586,In_709,In_189);
and U1587 (N_1587,In_383,In_182);
nor U1588 (N_1588,In_160,In_225);
and U1589 (N_1589,In_547,In_776);
xnor U1590 (N_1590,In_879,In_790);
or U1591 (N_1591,In_792,In_897);
nor U1592 (N_1592,In_829,In_933);
or U1593 (N_1593,In_602,In_874);
xor U1594 (N_1594,In_215,In_886);
nand U1595 (N_1595,In_795,In_279);
nand U1596 (N_1596,In_509,In_950);
nor U1597 (N_1597,In_689,In_791);
nor U1598 (N_1598,In_393,In_2);
or U1599 (N_1599,In_10,In_420);
and U1600 (N_1600,In_793,In_298);
or U1601 (N_1601,In_652,In_668);
nor U1602 (N_1602,In_697,In_814);
and U1603 (N_1603,In_416,In_740);
nor U1604 (N_1604,In_854,In_63);
nand U1605 (N_1605,In_660,In_456);
and U1606 (N_1606,In_416,In_102);
or U1607 (N_1607,In_843,In_507);
or U1608 (N_1608,In_116,In_167);
xnor U1609 (N_1609,In_402,In_8);
nor U1610 (N_1610,In_861,In_741);
xnor U1611 (N_1611,In_890,In_476);
nand U1612 (N_1612,In_492,In_666);
nor U1613 (N_1613,In_645,In_596);
nand U1614 (N_1614,In_456,In_606);
and U1615 (N_1615,In_172,In_361);
xor U1616 (N_1616,In_451,In_948);
and U1617 (N_1617,In_530,In_716);
or U1618 (N_1618,In_297,In_293);
nor U1619 (N_1619,In_263,In_197);
nor U1620 (N_1620,In_389,In_187);
and U1621 (N_1621,In_42,In_81);
nand U1622 (N_1622,In_791,In_494);
and U1623 (N_1623,In_780,In_713);
or U1624 (N_1624,In_442,In_670);
or U1625 (N_1625,In_833,In_162);
xnor U1626 (N_1626,In_84,In_784);
and U1627 (N_1627,In_133,In_267);
nand U1628 (N_1628,In_190,In_416);
nor U1629 (N_1629,In_258,In_356);
nand U1630 (N_1630,In_788,In_984);
nor U1631 (N_1631,In_599,In_147);
xnor U1632 (N_1632,In_124,In_227);
or U1633 (N_1633,In_575,In_867);
and U1634 (N_1634,In_958,In_477);
and U1635 (N_1635,In_759,In_139);
and U1636 (N_1636,In_692,In_942);
or U1637 (N_1637,In_606,In_304);
or U1638 (N_1638,In_704,In_222);
or U1639 (N_1639,In_109,In_587);
nand U1640 (N_1640,In_390,In_704);
and U1641 (N_1641,In_849,In_269);
nand U1642 (N_1642,In_258,In_822);
nand U1643 (N_1643,In_661,In_213);
and U1644 (N_1644,In_52,In_781);
nor U1645 (N_1645,In_484,In_970);
and U1646 (N_1646,In_521,In_839);
and U1647 (N_1647,In_328,In_26);
nor U1648 (N_1648,In_431,In_806);
xnor U1649 (N_1649,In_560,In_951);
or U1650 (N_1650,In_779,In_374);
xor U1651 (N_1651,In_0,In_562);
and U1652 (N_1652,In_991,In_283);
or U1653 (N_1653,In_309,In_222);
nand U1654 (N_1654,In_344,In_164);
nor U1655 (N_1655,In_184,In_994);
and U1656 (N_1656,In_660,In_761);
nand U1657 (N_1657,In_151,In_662);
or U1658 (N_1658,In_847,In_732);
nand U1659 (N_1659,In_788,In_654);
nand U1660 (N_1660,In_772,In_44);
and U1661 (N_1661,In_981,In_719);
and U1662 (N_1662,In_106,In_194);
nand U1663 (N_1663,In_366,In_836);
and U1664 (N_1664,In_199,In_593);
or U1665 (N_1665,In_851,In_492);
xnor U1666 (N_1666,In_58,In_647);
xor U1667 (N_1667,In_332,In_65);
and U1668 (N_1668,In_968,In_577);
nand U1669 (N_1669,In_252,In_634);
and U1670 (N_1670,In_997,In_205);
nand U1671 (N_1671,In_402,In_897);
nand U1672 (N_1672,In_993,In_840);
nand U1673 (N_1673,In_496,In_518);
nand U1674 (N_1674,In_620,In_585);
or U1675 (N_1675,In_327,In_806);
and U1676 (N_1676,In_794,In_231);
and U1677 (N_1677,In_61,In_910);
nand U1678 (N_1678,In_407,In_165);
nand U1679 (N_1679,In_483,In_963);
and U1680 (N_1680,In_615,In_291);
nor U1681 (N_1681,In_73,In_211);
and U1682 (N_1682,In_343,In_663);
and U1683 (N_1683,In_731,In_382);
nand U1684 (N_1684,In_852,In_936);
nand U1685 (N_1685,In_342,In_835);
nor U1686 (N_1686,In_655,In_565);
and U1687 (N_1687,In_993,In_283);
nor U1688 (N_1688,In_60,In_374);
nor U1689 (N_1689,In_799,In_465);
nand U1690 (N_1690,In_681,In_469);
nand U1691 (N_1691,In_842,In_876);
or U1692 (N_1692,In_550,In_701);
nand U1693 (N_1693,In_906,In_34);
and U1694 (N_1694,In_555,In_153);
xnor U1695 (N_1695,In_187,In_982);
nand U1696 (N_1696,In_162,In_406);
nor U1697 (N_1697,In_174,In_796);
and U1698 (N_1698,In_534,In_172);
nand U1699 (N_1699,In_375,In_198);
or U1700 (N_1700,In_279,In_712);
and U1701 (N_1701,In_969,In_257);
and U1702 (N_1702,In_989,In_838);
and U1703 (N_1703,In_687,In_62);
nand U1704 (N_1704,In_485,In_253);
nand U1705 (N_1705,In_574,In_603);
nor U1706 (N_1706,In_100,In_566);
nand U1707 (N_1707,In_321,In_163);
xnor U1708 (N_1708,In_193,In_212);
and U1709 (N_1709,In_75,In_453);
and U1710 (N_1710,In_687,In_357);
nor U1711 (N_1711,In_80,In_173);
or U1712 (N_1712,In_96,In_700);
and U1713 (N_1713,In_381,In_618);
nand U1714 (N_1714,In_391,In_681);
or U1715 (N_1715,In_664,In_534);
nor U1716 (N_1716,In_341,In_974);
nand U1717 (N_1717,In_601,In_456);
and U1718 (N_1718,In_329,In_119);
or U1719 (N_1719,In_915,In_631);
nand U1720 (N_1720,In_926,In_94);
and U1721 (N_1721,In_841,In_891);
and U1722 (N_1722,In_637,In_954);
and U1723 (N_1723,In_149,In_633);
and U1724 (N_1724,In_224,In_318);
nand U1725 (N_1725,In_448,In_955);
nand U1726 (N_1726,In_180,In_908);
nor U1727 (N_1727,In_17,In_807);
nand U1728 (N_1728,In_788,In_678);
and U1729 (N_1729,In_530,In_788);
nand U1730 (N_1730,In_683,In_602);
or U1731 (N_1731,In_428,In_137);
and U1732 (N_1732,In_45,In_963);
nand U1733 (N_1733,In_477,In_89);
nand U1734 (N_1734,In_25,In_705);
nand U1735 (N_1735,In_516,In_226);
or U1736 (N_1736,In_504,In_634);
nand U1737 (N_1737,In_333,In_255);
nor U1738 (N_1738,In_76,In_6);
nand U1739 (N_1739,In_406,In_174);
nand U1740 (N_1740,In_326,In_859);
nor U1741 (N_1741,In_198,In_736);
or U1742 (N_1742,In_364,In_804);
nor U1743 (N_1743,In_982,In_543);
xor U1744 (N_1744,In_347,In_78);
xor U1745 (N_1745,In_690,In_11);
nand U1746 (N_1746,In_520,In_795);
or U1747 (N_1747,In_543,In_475);
xor U1748 (N_1748,In_365,In_937);
and U1749 (N_1749,In_234,In_844);
nor U1750 (N_1750,In_659,In_930);
or U1751 (N_1751,In_452,In_412);
nor U1752 (N_1752,In_842,In_408);
or U1753 (N_1753,In_232,In_601);
and U1754 (N_1754,In_768,In_214);
xor U1755 (N_1755,In_92,In_723);
and U1756 (N_1756,In_759,In_781);
nor U1757 (N_1757,In_257,In_915);
nand U1758 (N_1758,In_578,In_710);
xor U1759 (N_1759,In_673,In_85);
nand U1760 (N_1760,In_247,In_871);
or U1761 (N_1761,In_341,In_546);
and U1762 (N_1762,In_653,In_640);
xnor U1763 (N_1763,In_994,In_230);
nand U1764 (N_1764,In_858,In_61);
nor U1765 (N_1765,In_538,In_514);
and U1766 (N_1766,In_976,In_282);
and U1767 (N_1767,In_284,In_532);
nand U1768 (N_1768,In_984,In_882);
and U1769 (N_1769,In_670,In_770);
or U1770 (N_1770,In_817,In_511);
nand U1771 (N_1771,In_559,In_583);
nor U1772 (N_1772,In_856,In_397);
or U1773 (N_1773,In_425,In_106);
nand U1774 (N_1774,In_379,In_950);
or U1775 (N_1775,In_370,In_194);
xnor U1776 (N_1776,In_534,In_535);
nand U1777 (N_1777,In_655,In_932);
and U1778 (N_1778,In_609,In_155);
xor U1779 (N_1779,In_755,In_318);
or U1780 (N_1780,In_43,In_254);
xor U1781 (N_1781,In_174,In_699);
or U1782 (N_1782,In_158,In_666);
and U1783 (N_1783,In_783,In_671);
nor U1784 (N_1784,In_881,In_413);
or U1785 (N_1785,In_449,In_205);
and U1786 (N_1786,In_556,In_134);
or U1787 (N_1787,In_132,In_901);
xor U1788 (N_1788,In_987,In_889);
or U1789 (N_1789,In_17,In_652);
or U1790 (N_1790,In_999,In_867);
or U1791 (N_1791,In_910,In_756);
nand U1792 (N_1792,In_8,In_940);
nor U1793 (N_1793,In_308,In_298);
nand U1794 (N_1794,In_355,In_733);
and U1795 (N_1795,In_205,In_348);
nor U1796 (N_1796,In_843,In_116);
or U1797 (N_1797,In_146,In_229);
or U1798 (N_1798,In_480,In_100);
or U1799 (N_1799,In_763,In_927);
or U1800 (N_1800,In_624,In_973);
nor U1801 (N_1801,In_157,In_336);
or U1802 (N_1802,In_288,In_718);
nor U1803 (N_1803,In_51,In_898);
nand U1804 (N_1804,In_472,In_598);
or U1805 (N_1805,In_791,In_258);
or U1806 (N_1806,In_134,In_647);
or U1807 (N_1807,In_271,In_875);
xnor U1808 (N_1808,In_922,In_83);
nor U1809 (N_1809,In_873,In_384);
xnor U1810 (N_1810,In_921,In_705);
nand U1811 (N_1811,In_496,In_752);
nand U1812 (N_1812,In_663,In_721);
nand U1813 (N_1813,In_218,In_879);
nand U1814 (N_1814,In_125,In_249);
and U1815 (N_1815,In_692,In_961);
or U1816 (N_1816,In_672,In_125);
or U1817 (N_1817,In_886,In_144);
and U1818 (N_1818,In_746,In_893);
xnor U1819 (N_1819,In_263,In_454);
nor U1820 (N_1820,In_523,In_101);
or U1821 (N_1821,In_721,In_131);
nand U1822 (N_1822,In_574,In_204);
nand U1823 (N_1823,In_21,In_928);
and U1824 (N_1824,In_400,In_354);
nor U1825 (N_1825,In_260,In_301);
and U1826 (N_1826,In_802,In_30);
xnor U1827 (N_1827,In_286,In_922);
nand U1828 (N_1828,In_26,In_914);
nor U1829 (N_1829,In_760,In_876);
nand U1830 (N_1830,In_100,In_980);
or U1831 (N_1831,In_939,In_813);
nand U1832 (N_1832,In_922,In_281);
nor U1833 (N_1833,In_319,In_151);
or U1834 (N_1834,In_422,In_239);
nor U1835 (N_1835,In_309,In_145);
nand U1836 (N_1836,In_120,In_992);
nand U1837 (N_1837,In_951,In_733);
or U1838 (N_1838,In_401,In_429);
and U1839 (N_1839,In_434,In_487);
nor U1840 (N_1840,In_395,In_940);
nor U1841 (N_1841,In_739,In_210);
nor U1842 (N_1842,In_225,In_550);
nor U1843 (N_1843,In_292,In_642);
and U1844 (N_1844,In_226,In_420);
or U1845 (N_1845,In_8,In_901);
or U1846 (N_1846,In_113,In_464);
nor U1847 (N_1847,In_400,In_606);
nor U1848 (N_1848,In_9,In_515);
xnor U1849 (N_1849,In_324,In_707);
and U1850 (N_1850,In_639,In_98);
and U1851 (N_1851,In_591,In_520);
and U1852 (N_1852,In_948,In_454);
and U1853 (N_1853,In_59,In_41);
nor U1854 (N_1854,In_581,In_725);
and U1855 (N_1855,In_60,In_712);
nand U1856 (N_1856,In_811,In_563);
nor U1857 (N_1857,In_190,In_849);
nor U1858 (N_1858,In_581,In_396);
or U1859 (N_1859,In_85,In_867);
nor U1860 (N_1860,In_798,In_752);
nor U1861 (N_1861,In_259,In_165);
or U1862 (N_1862,In_100,In_269);
nor U1863 (N_1863,In_115,In_597);
or U1864 (N_1864,In_763,In_148);
nand U1865 (N_1865,In_927,In_787);
or U1866 (N_1866,In_284,In_998);
nor U1867 (N_1867,In_656,In_47);
nor U1868 (N_1868,In_35,In_274);
nor U1869 (N_1869,In_810,In_527);
nand U1870 (N_1870,In_170,In_400);
and U1871 (N_1871,In_920,In_569);
nand U1872 (N_1872,In_326,In_391);
xor U1873 (N_1873,In_446,In_171);
and U1874 (N_1874,In_939,In_518);
nand U1875 (N_1875,In_795,In_608);
and U1876 (N_1876,In_788,In_674);
nand U1877 (N_1877,In_964,In_952);
xnor U1878 (N_1878,In_239,In_260);
and U1879 (N_1879,In_804,In_778);
nor U1880 (N_1880,In_412,In_844);
nand U1881 (N_1881,In_30,In_674);
nor U1882 (N_1882,In_942,In_339);
or U1883 (N_1883,In_935,In_966);
nand U1884 (N_1884,In_531,In_34);
or U1885 (N_1885,In_233,In_918);
or U1886 (N_1886,In_293,In_113);
xor U1887 (N_1887,In_522,In_298);
or U1888 (N_1888,In_734,In_5);
nand U1889 (N_1889,In_715,In_185);
xnor U1890 (N_1890,In_15,In_640);
nand U1891 (N_1891,In_828,In_523);
nor U1892 (N_1892,In_32,In_415);
or U1893 (N_1893,In_471,In_426);
and U1894 (N_1894,In_594,In_657);
nand U1895 (N_1895,In_804,In_407);
nor U1896 (N_1896,In_561,In_190);
nor U1897 (N_1897,In_162,In_965);
or U1898 (N_1898,In_422,In_655);
nor U1899 (N_1899,In_457,In_722);
or U1900 (N_1900,In_416,In_16);
or U1901 (N_1901,In_378,In_87);
nor U1902 (N_1902,In_945,In_930);
nor U1903 (N_1903,In_715,In_160);
or U1904 (N_1904,In_164,In_303);
or U1905 (N_1905,In_655,In_466);
or U1906 (N_1906,In_428,In_159);
nand U1907 (N_1907,In_436,In_886);
nand U1908 (N_1908,In_413,In_922);
nand U1909 (N_1909,In_842,In_483);
or U1910 (N_1910,In_352,In_439);
and U1911 (N_1911,In_968,In_896);
nand U1912 (N_1912,In_538,In_334);
nor U1913 (N_1913,In_151,In_773);
nand U1914 (N_1914,In_343,In_214);
and U1915 (N_1915,In_204,In_935);
nor U1916 (N_1916,In_21,In_979);
or U1917 (N_1917,In_643,In_836);
nand U1918 (N_1918,In_212,In_128);
xor U1919 (N_1919,In_361,In_946);
nand U1920 (N_1920,In_774,In_829);
nand U1921 (N_1921,In_533,In_557);
nor U1922 (N_1922,In_817,In_320);
nor U1923 (N_1923,In_600,In_420);
xor U1924 (N_1924,In_861,In_14);
nand U1925 (N_1925,In_309,In_661);
nand U1926 (N_1926,In_111,In_554);
nor U1927 (N_1927,In_461,In_582);
nor U1928 (N_1928,In_116,In_930);
and U1929 (N_1929,In_893,In_662);
nor U1930 (N_1930,In_755,In_389);
and U1931 (N_1931,In_435,In_13);
or U1932 (N_1932,In_364,In_614);
or U1933 (N_1933,In_48,In_509);
nand U1934 (N_1934,In_294,In_320);
and U1935 (N_1935,In_935,In_670);
and U1936 (N_1936,In_365,In_184);
and U1937 (N_1937,In_712,In_366);
nand U1938 (N_1938,In_111,In_275);
and U1939 (N_1939,In_381,In_556);
and U1940 (N_1940,In_450,In_318);
or U1941 (N_1941,In_764,In_817);
or U1942 (N_1942,In_587,In_541);
nand U1943 (N_1943,In_92,In_155);
nor U1944 (N_1944,In_694,In_74);
nor U1945 (N_1945,In_764,In_643);
nand U1946 (N_1946,In_795,In_509);
and U1947 (N_1947,In_547,In_315);
or U1948 (N_1948,In_415,In_692);
or U1949 (N_1949,In_398,In_450);
or U1950 (N_1950,In_614,In_756);
and U1951 (N_1951,In_557,In_888);
and U1952 (N_1952,In_233,In_88);
nor U1953 (N_1953,In_188,In_834);
and U1954 (N_1954,In_463,In_59);
xor U1955 (N_1955,In_381,In_78);
nand U1956 (N_1956,In_100,In_67);
or U1957 (N_1957,In_811,In_458);
nand U1958 (N_1958,In_73,In_835);
or U1959 (N_1959,In_11,In_855);
and U1960 (N_1960,In_516,In_344);
nand U1961 (N_1961,In_836,In_271);
xor U1962 (N_1962,In_991,In_435);
nor U1963 (N_1963,In_581,In_792);
and U1964 (N_1964,In_693,In_187);
or U1965 (N_1965,In_816,In_970);
nand U1966 (N_1966,In_504,In_361);
nor U1967 (N_1967,In_769,In_979);
nor U1968 (N_1968,In_326,In_623);
nand U1969 (N_1969,In_479,In_240);
nand U1970 (N_1970,In_700,In_222);
or U1971 (N_1971,In_462,In_680);
nor U1972 (N_1972,In_658,In_347);
and U1973 (N_1973,In_863,In_492);
nand U1974 (N_1974,In_379,In_734);
nand U1975 (N_1975,In_277,In_678);
nand U1976 (N_1976,In_341,In_138);
and U1977 (N_1977,In_116,In_62);
or U1978 (N_1978,In_534,In_608);
nand U1979 (N_1979,In_384,In_712);
nor U1980 (N_1980,In_683,In_173);
nor U1981 (N_1981,In_717,In_217);
xor U1982 (N_1982,In_891,In_78);
nand U1983 (N_1983,In_950,In_669);
nand U1984 (N_1984,In_796,In_528);
or U1985 (N_1985,In_791,In_105);
xor U1986 (N_1986,In_368,In_1);
or U1987 (N_1987,In_80,In_176);
nor U1988 (N_1988,In_643,In_785);
nand U1989 (N_1989,In_369,In_690);
nor U1990 (N_1990,In_144,In_660);
or U1991 (N_1991,In_149,In_239);
nor U1992 (N_1992,In_315,In_339);
and U1993 (N_1993,In_414,In_118);
nor U1994 (N_1994,In_500,In_451);
and U1995 (N_1995,In_521,In_564);
nand U1996 (N_1996,In_538,In_289);
and U1997 (N_1997,In_850,In_436);
nor U1998 (N_1998,In_459,In_305);
nor U1999 (N_1999,In_790,In_743);
nor U2000 (N_2000,In_166,In_99);
nand U2001 (N_2001,In_528,In_819);
and U2002 (N_2002,In_228,In_928);
nor U2003 (N_2003,In_448,In_430);
or U2004 (N_2004,In_632,In_994);
and U2005 (N_2005,In_651,In_213);
and U2006 (N_2006,In_829,In_307);
nor U2007 (N_2007,In_87,In_734);
nor U2008 (N_2008,In_529,In_202);
nor U2009 (N_2009,In_237,In_243);
nand U2010 (N_2010,In_558,In_363);
nor U2011 (N_2011,In_166,In_640);
nor U2012 (N_2012,In_814,In_148);
nand U2013 (N_2013,In_136,In_493);
nor U2014 (N_2014,In_715,In_505);
or U2015 (N_2015,In_40,In_208);
and U2016 (N_2016,In_765,In_895);
and U2017 (N_2017,In_504,In_881);
nor U2018 (N_2018,In_24,In_290);
xor U2019 (N_2019,In_833,In_565);
and U2020 (N_2020,In_556,In_380);
nor U2021 (N_2021,In_315,In_826);
nand U2022 (N_2022,In_306,In_687);
nor U2023 (N_2023,In_162,In_485);
or U2024 (N_2024,In_505,In_925);
xnor U2025 (N_2025,In_708,In_714);
nor U2026 (N_2026,In_307,In_104);
and U2027 (N_2027,In_60,In_682);
or U2028 (N_2028,In_225,In_590);
or U2029 (N_2029,In_607,In_722);
or U2030 (N_2030,In_974,In_60);
and U2031 (N_2031,In_999,In_754);
xnor U2032 (N_2032,In_286,In_697);
xor U2033 (N_2033,In_63,In_122);
xor U2034 (N_2034,In_492,In_269);
xnor U2035 (N_2035,In_233,In_356);
nor U2036 (N_2036,In_941,In_203);
and U2037 (N_2037,In_490,In_311);
nand U2038 (N_2038,In_470,In_15);
or U2039 (N_2039,In_927,In_277);
and U2040 (N_2040,In_773,In_251);
nand U2041 (N_2041,In_455,In_347);
nor U2042 (N_2042,In_503,In_217);
and U2043 (N_2043,In_39,In_652);
or U2044 (N_2044,In_88,In_629);
or U2045 (N_2045,In_87,In_31);
and U2046 (N_2046,In_475,In_324);
nor U2047 (N_2047,In_823,In_474);
and U2048 (N_2048,In_132,In_162);
xor U2049 (N_2049,In_149,In_227);
xor U2050 (N_2050,In_951,In_510);
or U2051 (N_2051,In_564,In_357);
xnor U2052 (N_2052,In_159,In_173);
or U2053 (N_2053,In_277,In_160);
nand U2054 (N_2054,In_405,In_871);
and U2055 (N_2055,In_559,In_94);
or U2056 (N_2056,In_821,In_24);
and U2057 (N_2057,In_556,In_789);
and U2058 (N_2058,In_592,In_769);
nor U2059 (N_2059,In_255,In_623);
and U2060 (N_2060,In_833,In_837);
and U2061 (N_2061,In_34,In_463);
nand U2062 (N_2062,In_256,In_96);
nand U2063 (N_2063,In_644,In_637);
nor U2064 (N_2064,In_260,In_98);
nor U2065 (N_2065,In_752,In_907);
xor U2066 (N_2066,In_590,In_262);
and U2067 (N_2067,In_364,In_894);
and U2068 (N_2068,In_271,In_549);
or U2069 (N_2069,In_541,In_928);
and U2070 (N_2070,In_483,In_500);
and U2071 (N_2071,In_682,In_549);
nor U2072 (N_2072,In_636,In_343);
xnor U2073 (N_2073,In_313,In_431);
nor U2074 (N_2074,In_105,In_440);
nand U2075 (N_2075,In_542,In_6);
nand U2076 (N_2076,In_439,In_491);
xor U2077 (N_2077,In_313,In_251);
nor U2078 (N_2078,In_869,In_183);
nor U2079 (N_2079,In_455,In_538);
or U2080 (N_2080,In_908,In_299);
nor U2081 (N_2081,In_403,In_155);
and U2082 (N_2082,In_158,In_276);
nand U2083 (N_2083,In_236,In_967);
nor U2084 (N_2084,In_543,In_394);
nand U2085 (N_2085,In_402,In_488);
or U2086 (N_2086,In_698,In_815);
xnor U2087 (N_2087,In_759,In_486);
or U2088 (N_2088,In_363,In_587);
nor U2089 (N_2089,In_371,In_51);
nand U2090 (N_2090,In_950,In_146);
and U2091 (N_2091,In_173,In_883);
and U2092 (N_2092,In_24,In_464);
or U2093 (N_2093,In_22,In_512);
and U2094 (N_2094,In_167,In_608);
nor U2095 (N_2095,In_885,In_593);
nor U2096 (N_2096,In_70,In_596);
nand U2097 (N_2097,In_897,In_571);
or U2098 (N_2098,In_866,In_362);
or U2099 (N_2099,In_220,In_15);
xnor U2100 (N_2100,In_724,In_156);
and U2101 (N_2101,In_311,In_868);
xor U2102 (N_2102,In_19,In_502);
nand U2103 (N_2103,In_968,In_148);
xnor U2104 (N_2104,In_272,In_78);
or U2105 (N_2105,In_245,In_861);
nor U2106 (N_2106,In_617,In_327);
or U2107 (N_2107,In_300,In_424);
nand U2108 (N_2108,In_647,In_249);
and U2109 (N_2109,In_468,In_633);
nand U2110 (N_2110,In_640,In_462);
and U2111 (N_2111,In_321,In_581);
nand U2112 (N_2112,In_410,In_507);
xor U2113 (N_2113,In_566,In_562);
or U2114 (N_2114,In_114,In_985);
nor U2115 (N_2115,In_143,In_804);
nand U2116 (N_2116,In_626,In_144);
nand U2117 (N_2117,In_401,In_616);
nor U2118 (N_2118,In_178,In_108);
or U2119 (N_2119,In_963,In_674);
and U2120 (N_2120,In_57,In_173);
or U2121 (N_2121,In_30,In_439);
and U2122 (N_2122,In_430,In_729);
and U2123 (N_2123,In_629,In_293);
and U2124 (N_2124,In_614,In_854);
xnor U2125 (N_2125,In_155,In_916);
and U2126 (N_2126,In_721,In_926);
and U2127 (N_2127,In_579,In_837);
nand U2128 (N_2128,In_481,In_859);
nand U2129 (N_2129,In_216,In_770);
nor U2130 (N_2130,In_21,In_765);
nand U2131 (N_2131,In_591,In_356);
nand U2132 (N_2132,In_905,In_928);
nand U2133 (N_2133,In_483,In_168);
nor U2134 (N_2134,In_488,In_838);
or U2135 (N_2135,In_152,In_746);
nand U2136 (N_2136,In_73,In_82);
and U2137 (N_2137,In_801,In_883);
and U2138 (N_2138,In_152,In_0);
nor U2139 (N_2139,In_381,In_377);
xor U2140 (N_2140,In_506,In_35);
and U2141 (N_2141,In_18,In_581);
nand U2142 (N_2142,In_928,In_437);
nand U2143 (N_2143,In_280,In_54);
and U2144 (N_2144,In_926,In_360);
or U2145 (N_2145,In_832,In_488);
nor U2146 (N_2146,In_209,In_565);
and U2147 (N_2147,In_569,In_129);
nand U2148 (N_2148,In_405,In_385);
or U2149 (N_2149,In_208,In_848);
nand U2150 (N_2150,In_574,In_630);
or U2151 (N_2151,In_371,In_466);
or U2152 (N_2152,In_36,In_755);
or U2153 (N_2153,In_645,In_900);
nand U2154 (N_2154,In_892,In_139);
nor U2155 (N_2155,In_513,In_850);
nand U2156 (N_2156,In_463,In_858);
nand U2157 (N_2157,In_432,In_625);
or U2158 (N_2158,In_423,In_294);
or U2159 (N_2159,In_725,In_980);
and U2160 (N_2160,In_370,In_982);
or U2161 (N_2161,In_691,In_875);
or U2162 (N_2162,In_586,In_693);
or U2163 (N_2163,In_874,In_78);
nor U2164 (N_2164,In_29,In_376);
nand U2165 (N_2165,In_379,In_256);
nand U2166 (N_2166,In_789,In_366);
and U2167 (N_2167,In_804,In_350);
nand U2168 (N_2168,In_844,In_600);
and U2169 (N_2169,In_703,In_268);
and U2170 (N_2170,In_242,In_840);
and U2171 (N_2171,In_375,In_786);
and U2172 (N_2172,In_345,In_78);
nor U2173 (N_2173,In_465,In_851);
nor U2174 (N_2174,In_611,In_404);
nand U2175 (N_2175,In_559,In_181);
nand U2176 (N_2176,In_441,In_700);
and U2177 (N_2177,In_844,In_373);
or U2178 (N_2178,In_114,In_881);
and U2179 (N_2179,In_162,In_34);
nand U2180 (N_2180,In_224,In_797);
xnor U2181 (N_2181,In_443,In_762);
nor U2182 (N_2182,In_485,In_849);
nor U2183 (N_2183,In_181,In_938);
nor U2184 (N_2184,In_679,In_930);
nand U2185 (N_2185,In_418,In_828);
and U2186 (N_2186,In_255,In_590);
nor U2187 (N_2187,In_48,In_297);
or U2188 (N_2188,In_303,In_161);
or U2189 (N_2189,In_129,In_622);
xor U2190 (N_2190,In_87,In_289);
nor U2191 (N_2191,In_760,In_984);
or U2192 (N_2192,In_964,In_121);
nand U2193 (N_2193,In_233,In_986);
nor U2194 (N_2194,In_934,In_7);
and U2195 (N_2195,In_911,In_589);
nand U2196 (N_2196,In_974,In_450);
nand U2197 (N_2197,In_233,In_355);
nor U2198 (N_2198,In_660,In_733);
xnor U2199 (N_2199,In_510,In_87);
and U2200 (N_2200,In_333,In_785);
nor U2201 (N_2201,In_895,In_34);
and U2202 (N_2202,In_692,In_419);
or U2203 (N_2203,In_643,In_913);
nor U2204 (N_2204,In_86,In_299);
and U2205 (N_2205,In_687,In_449);
and U2206 (N_2206,In_913,In_175);
or U2207 (N_2207,In_921,In_280);
nor U2208 (N_2208,In_705,In_104);
nand U2209 (N_2209,In_715,In_242);
and U2210 (N_2210,In_804,In_718);
nor U2211 (N_2211,In_93,In_465);
nand U2212 (N_2212,In_718,In_886);
nand U2213 (N_2213,In_433,In_824);
and U2214 (N_2214,In_329,In_38);
nand U2215 (N_2215,In_717,In_203);
nand U2216 (N_2216,In_470,In_429);
nand U2217 (N_2217,In_684,In_260);
nand U2218 (N_2218,In_850,In_302);
xor U2219 (N_2219,In_924,In_116);
nor U2220 (N_2220,In_268,In_231);
or U2221 (N_2221,In_742,In_345);
and U2222 (N_2222,In_326,In_792);
or U2223 (N_2223,In_908,In_147);
nand U2224 (N_2224,In_788,In_729);
xnor U2225 (N_2225,In_74,In_350);
nor U2226 (N_2226,In_460,In_667);
xor U2227 (N_2227,In_288,In_860);
nand U2228 (N_2228,In_865,In_442);
nand U2229 (N_2229,In_954,In_945);
nand U2230 (N_2230,In_232,In_728);
or U2231 (N_2231,In_726,In_442);
nor U2232 (N_2232,In_109,In_801);
nand U2233 (N_2233,In_636,In_246);
xnor U2234 (N_2234,In_306,In_111);
and U2235 (N_2235,In_44,In_816);
or U2236 (N_2236,In_505,In_88);
xnor U2237 (N_2237,In_30,In_121);
nor U2238 (N_2238,In_76,In_940);
nor U2239 (N_2239,In_755,In_325);
or U2240 (N_2240,In_114,In_511);
or U2241 (N_2241,In_153,In_691);
nor U2242 (N_2242,In_291,In_380);
nand U2243 (N_2243,In_595,In_733);
nor U2244 (N_2244,In_350,In_87);
or U2245 (N_2245,In_18,In_43);
nor U2246 (N_2246,In_836,In_308);
and U2247 (N_2247,In_987,In_618);
and U2248 (N_2248,In_352,In_219);
nand U2249 (N_2249,In_236,In_358);
and U2250 (N_2250,In_716,In_114);
and U2251 (N_2251,In_879,In_770);
nand U2252 (N_2252,In_403,In_23);
and U2253 (N_2253,In_313,In_908);
nand U2254 (N_2254,In_115,In_551);
nand U2255 (N_2255,In_556,In_419);
or U2256 (N_2256,In_42,In_398);
xor U2257 (N_2257,In_361,In_680);
xnor U2258 (N_2258,In_330,In_627);
nor U2259 (N_2259,In_934,In_641);
nor U2260 (N_2260,In_692,In_243);
nand U2261 (N_2261,In_346,In_418);
nand U2262 (N_2262,In_194,In_204);
and U2263 (N_2263,In_239,In_505);
xor U2264 (N_2264,In_499,In_463);
and U2265 (N_2265,In_478,In_553);
nor U2266 (N_2266,In_170,In_922);
nor U2267 (N_2267,In_981,In_598);
nor U2268 (N_2268,In_896,In_814);
and U2269 (N_2269,In_393,In_263);
xor U2270 (N_2270,In_98,In_888);
nor U2271 (N_2271,In_551,In_795);
or U2272 (N_2272,In_418,In_67);
xnor U2273 (N_2273,In_172,In_52);
nand U2274 (N_2274,In_626,In_387);
and U2275 (N_2275,In_863,In_965);
or U2276 (N_2276,In_90,In_395);
xor U2277 (N_2277,In_655,In_392);
or U2278 (N_2278,In_946,In_630);
nor U2279 (N_2279,In_346,In_490);
nand U2280 (N_2280,In_313,In_885);
nor U2281 (N_2281,In_196,In_733);
nor U2282 (N_2282,In_759,In_314);
and U2283 (N_2283,In_777,In_975);
nand U2284 (N_2284,In_315,In_351);
or U2285 (N_2285,In_882,In_761);
nor U2286 (N_2286,In_61,In_804);
nor U2287 (N_2287,In_61,In_173);
nor U2288 (N_2288,In_481,In_820);
nand U2289 (N_2289,In_40,In_7);
and U2290 (N_2290,In_364,In_991);
nand U2291 (N_2291,In_687,In_47);
and U2292 (N_2292,In_476,In_414);
nor U2293 (N_2293,In_159,In_655);
nand U2294 (N_2294,In_295,In_473);
or U2295 (N_2295,In_474,In_959);
or U2296 (N_2296,In_212,In_771);
nor U2297 (N_2297,In_522,In_844);
and U2298 (N_2298,In_631,In_70);
nand U2299 (N_2299,In_728,In_173);
nand U2300 (N_2300,In_69,In_446);
and U2301 (N_2301,In_885,In_904);
xor U2302 (N_2302,In_113,In_550);
or U2303 (N_2303,In_556,In_813);
nor U2304 (N_2304,In_552,In_973);
nand U2305 (N_2305,In_424,In_463);
or U2306 (N_2306,In_963,In_374);
nor U2307 (N_2307,In_912,In_443);
nor U2308 (N_2308,In_352,In_615);
nand U2309 (N_2309,In_324,In_343);
or U2310 (N_2310,In_961,In_608);
nand U2311 (N_2311,In_376,In_963);
xnor U2312 (N_2312,In_671,In_737);
or U2313 (N_2313,In_44,In_192);
or U2314 (N_2314,In_535,In_764);
xor U2315 (N_2315,In_975,In_716);
or U2316 (N_2316,In_994,In_316);
xnor U2317 (N_2317,In_714,In_813);
xor U2318 (N_2318,In_686,In_77);
and U2319 (N_2319,In_884,In_328);
nand U2320 (N_2320,In_816,In_400);
nand U2321 (N_2321,In_695,In_744);
nor U2322 (N_2322,In_326,In_475);
and U2323 (N_2323,In_662,In_758);
and U2324 (N_2324,In_961,In_39);
nand U2325 (N_2325,In_968,In_181);
or U2326 (N_2326,In_694,In_950);
or U2327 (N_2327,In_502,In_254);
or U2328 (N_2328,In_419,In_70);
nand U2329 (N_2329,In_474,In_346);
and U2330 (N_2330,In_235,In_141);
or U2331 (N_2331,In_345,In_454);
xor U2332 (N_2332,In_490,In_877);
and U2333 (N_2333,In_150,In_714);
xnor U2334 (N_2334,In_184,In_706);
xor U2335 (N_2335,In_225,In_530);
xnor U2336 (N_2336,In_749,In_187);
nand U2337 (N_2337,In_528,In_328);
nand U2338 (N_2338,In_131,In_267);
nor U2339 (N_2339,In_280,In_48);
or U2340 (N_2340,In_132,In_248);
nor U2341 (N_2341,In_462,In_873);
nand U2342 (N_2342,In_282,In_244);
nor U2343 (N_2343,In_895,In_214);
nor U2344 (N_2344,In_209,In_688);
and U2345 (N_2345,In_551,In_992);
and U2346 (N_2346,In_846,In_723);
xor U2347 (N_2347,In_414,In_906);
or U2348 (N_2348,In_93,In_845);
xor U2349 (N_2349,In_688,In_358);
xor U2350 (N_2350,In_452,In_767);
nor U2351 (N_2351,In_502,In_382);
xor U2352 (N_2352,In_779,In_826);
and U2353 (N_2353,In_21,In_902);
and U2354 (N_2354,In_802,In_425);
nand U2355 (N_2355,In_156,In_613);
and U2356 (N_2356,In_680,In_690);
nand U2357 (N_2357,In_510,In_315);
or U2358 (N_2358,In_719,In_393);
and U2359 (N_2359,In_14,In_713);
nor U2360 (N_2360,In_848,In_548);
xnor U2361 (N_2361,In_67,In_998);
and U2362 (N_2362,In_824,In_757);
and U2363 (N_2363,In_705,In_687);
or U2364 (N_2364,In_836,In_763);
nor U2365 (N_2365,In_630,In_952);
xor U2366 (N_2366,In_683,In_426);
or U2367 (N_2367,In_224,In_599);
or U2368 (N_2368,In_139,In_802);
or U2369 (N_2369,In_275,In_660);
nand U2370 (N_2370,In_601,In_654);
and U2371 (N_2371,In_621,In_806);
xor U2372 (N_2372,In_431,In_457);
or U2373 (N_2373,In_930,In_121);
or U2374 (N_2374,In_610,In_211);
nand U2375 (N_2375,In_788,In_863);
and U2376 (N_2376,In_872,In_382);
nor U2377 (N_2377,In_774,In_980);
nand U2378 (N_2378,In_633,In_682);
nand U2379 (N_2379,In_149,In_951);
and U2380 (N_2380,In_367,In_537);
or U2381 (N_2381,In_851,In_69);
nand U2382 (N_2382,In_332,In_372);
or U2383 (N_2383,In_245,In_780);
or U2384 (N_2384,In_894,In_951);
or U2385 (N_2385,In_983,In_871);
xor U2386 (N_2386,In_792,In_542);
and U2387 (N_2387,In_398,In_128);
nor U2388 (N_2388,In_495,In_35);
or U2389 (N_2389,In_436,In_334);
and U2390 (N_2390,In_644,In_875);
nor U2391 (N_2391,In_419,In_802);
or U2392 (N_2392,In_439,In_725);
nand U2393 (N_2393,In_225,In_516);
nor U2394 (N_2394,In_297,In_564);
xor U2395 (N_2395,In_862,In_699);
and U2396 (N_2396,In_685,In_909);
nand U2397 (N_2397,In_704,In_121);
or U2398 (N_2398,In_426,In_316);
nand U2399 (N_2399,In_119,In_920);
xnor U2400 (N_2400,In_894,In_765);
nand U2401 (N_2401,In_409,In_482);
nand U2402 (N_2402,In_768,In_227);
nand U2403 (N_2403,In_850,In_780);
and U2404 (N_2404,In_768,In_992);
nor U2405 (N_2405,In_910,In_509);
nor U2406 (N_2406,In_214,In_460);
and U2407 (N_2407,In_330,In_807);
or U2408 (N_2408,In_482,In_27);
nand U2409 (N_2409,In_275,In_63);
or U2410 (N_2410,In_118,In_176);
or U2411 (N_2411,In_903,In_526);
and U2412 (N_2412,In_967,In_571);
or U2413 (N_2413,In_632,In_674);
nand U2414 (N_2414,In_877,In_414);
and U2415 (N_2415,In_363,In_518);
nor U2416 (N_2416,In_276,In_729);
or U2417 (N_2417,In_958,In_304);
nand U2418 (N_2418,In_532,In_19);
xor U2419 (N_2419,In_936,In_254);
and U2420 (N_2420,In_494,In_479);
or U2421 (N_2421,In_168,In_573);
nor U2422 (N_2422,In_817,In_500);
nand U2423 (N_2423,In_200,In_243);
xnor U2424 (N_2424,In_315,In_730);
and U2425 (N_2425,In_490,In_366);
or U2426 (N_2426,In_675,In_222);
xnor U2427 (N_2427,In_770,In_545);
nand U2428 (N_2428,In_997,In_216);
or U2429 (N_2429,In_307,In_628);
or U2430 (N_2430,In_710,In_770);
or U2431 (N_2431,In_670,In_718);
and U2432 (N_2432,In_128,In_894);
or U2433 (N_2433,In_765,In_129);
or U2434 (N_2434,In_656,In_459);
or U2435 (N_2435,In_18,In_287);
nor U2436 (N_2436,In_968,In_252);
or U2437 (N_2437,In_991,In_878);
nor U2438 (N_2438,In_310,In_417);
or U2439 (N_2439,In_99,In_88);
nand U2440 (N_2440,In_669,In_193);
xor U2441 (N_2441,In_868,In_287);
xnor U2442 (N_2442,In_673,In_808);
nor U2443 (N_2443,In_300,In_731);
and U2444 (N_2444,In_678,In_144);
nand U2445 (N_2445,In_876,In_431);
nor U2446 (N_2446,In_421,In_967);
nor U2447 (N_2447,In_443,In_33);
nand U2448 (N_2448,In_162,In_876);
nor U2449 (N_2449,In_557,In_43);
and U2450 (N_2450,In_840,In_134);
nand U2451 (N_2451,In_945,In_103);
or U2452 (N_2452,In_825,In_810);
nor U2453 (N_2453,In_394,In_623);
nand U2454 (N_2454,In_336,In_978);
and U2455 (N_2455,In_646,In_680);
and U2456 (N_2456,In_141,In_940);
xnor U2457 (N_2457,In_374,In_840);
and U2458 (N_2458,In_922,In_404);
or U2459 (N_2459,In_884,In_292);
nor U2460 (N_2460,In_372,In_829);
nor U2461 (N_2461,In_921,In_854);
and U2462 (N_2462,In_855,In_406);
and U2463 (N_2463,In_528,In_750);
or U2464 (N_2464,In_413,In_19);
or U2465 (N_2465,In_701,In_930);
or U2466 (N_2466,In_273,In_344);
and U2467 (N_2467,In_350,In_553);
or U2468 (N_2468,In_961,In_797);
xnor U2469 (N_2469,In_857,In_222);
and U2470 (N_2470,In_360,In_341);
nor U2471 (N_2471,In_417,In_896);
nor U2472 (N_2472,In_175,In_487);
nor U2473 (N_2473,In_33,In_79);
nor U2474 (N_2474,In_225,In_279);
xor U2475 (N_2475,In_400,In_93);
and U2476 (N_2476,In_565,In_170);
nand U2477 (N_2477,In_137,In_639);
nor U2478 (N_2478,In_892,In_386);
or U2479 (N_2479,In_128,In_98);
and U2480 (N_2480,In_918,In_283);
nand U2481 (N_2481,In_813,In_850);
and U2482 (N_2482,In_563,In_352);
nor U2483 (N_2483,In_830,In_930);
nand U2484 (N_2484,In_189,In_303);
or U2485 (N_2485,In_949,In_897);
and U2486 (N_2486,In_630,In_397);
or U2487 (N_2487,In_72,In_859);
xnor U2488 (N_2488,In_234,In_170);
nor U2489 (N_2489,In_247,In_798);
and U2490 (N_2490,In_906,In_958);
or U2491 (N_2491,In_703,In_450);
nor U2492 (N_2492,In_172,In_123);
and U2493 (N_2493,In_845,In_665);
nand U2494 (N_2494,In_662,In_640);
nor U2495 (N_2495,In_116,In_274);
nand U2496 (N_2496,In_155,In_283);
nand U2497 (N_2497,In_384,In_926);
xnor U2498 (N_2498,In_667,In_416);
nor U2499 (N_2499,In_929,In_257);
or U2500 (N_2500,In_52,In_265);
nor U2501 (N_2501,In_244,In_6);
nor U2502 (N_2502,In_517,In_717);
or U2503 (N_2503,In_433,In_423);
and U2504 (N_2504,In_441,In_779);
xor U2505 (N_2505,In_640,In_503);
or U2506 (N_2506,In_308,In_219);
nor U2507 (N_2507,In_994,In_139);
or U2508 (N_2508,In_643,In_515);
and U2509 (N_2509,In_616,In_839);
nand U2510 (N_2510,In_248,In_638);
nand U2511 (N_2511,In_639,In_379);
nand U2512 (N_2512,In_341,In_184);
nand U2513 (N_2513,In_297,In_922);
or U2514 (N_2514,In_269,In_356);
nor U2515 (N_2515,In_500,In_357);
and U2516 (N_2516,In_396,In_754);
nand U2517 (N_2517,In_873,In_425);
xnor U2518 (N_2518,In_920,In_919);
or U2519 (N_2519,In_884,In_862);
or U2520 (N_2520,In_387,In_669);
and U2521 (N_2521,In_960,In_318);
nand U2522 (N_2522,In_474,In_857);
or U2523 (N_2523,In_838,In_30);
nor U2524 (N_2524,In_757,In_17);
xor U2525 (N_2525,In_66,In_143);
or U2526 (N_2526,In_359,In_895);
or U2527 (N_2527,In_244,In_215);
and U2528 (N_2528,In_714,In_89);
and U2529 (N_2529,In_332,In_632);
or U2530 (N_2530,In_615,In_711);
and U2531 (N_2531,In_69,In_861);
nor U2532 (N_2532,In_774,In_407);
nand U2533 (N_2533,In_936,In_357);
and U2534 (N_2534,In_771,In_93);
nor U2535 (N_2535,In_167,In_890);
or U2536 (N_2536,In_843,In_30);
and U2537 (N_2537,In_432,In_718);
and U2538 (N_2538,In_150,In_524);
and U2539 (N_2539,In_167,In_492);
nand U2540 (N_2540,In_524,In_365);
nor U2541 (N_2541,In_844,In_59);
nand U2542 (N_2542,In_533,In_155);
nand U2543 (N_2543,In_752,In_572);
nor U2544 (N_2544,In_878,In_797);
nor U2545 (N_2545,In_20,In_653);
or U2546 (N_2546,In_863,In_262);
or U2547 (N_2547,In_489,In_313);
nor U2548 (N_2548,In_991,In_270);
nand U2549 (N_2549,In_243,In_697);
or U2550 (N_2550,In_370,In_609);
xor U2551 (N_2551,In_47,In_527);
nand U2552 (N_2552,In_433,In_285);
nor U2553 (N_2553,In_75,In_766);
or U2554 (N_2554,In_864,In_881);
and U2555 (N_2555,In_616,In_877);
nand U2556 (N_2556,In_887,In_239);
or U2557 (N_2557,In_849,In_553);
nor U2558 (N_2558,In_843,In_969);
nand U2559 (N_2559,In_782,In_413);
or U2560 (N_2560,In_797,In_368);
and U2561 (N_2561,In_350,In_579);
xor U2562 (N_2562,In_538,In_157);
nand U2563 (N_2563,In_136,In_303);
nand U2564 (N_2564,In_7,In_885);
and U2565 (N_2565,In_3,In_428);
and U2566 (N_2566,In_467,In_632);
and U2567 (N_2567,In_947,In_182);
xnor U2568 (N_2568,In_636,In_428);
nor U2569 (N_2569,In_870,In_905);
and U2570 (N_2570,In_112,In_482);
nand U2571 (N_2571,In_25,In_458);
and U2572 (N_2572,In_713,In_996);
nor U2573 (N_2573,In_293,In_829);
and U2574 (N_2574,In_522,In_389);
nand U2575 (N_2575,In_183,In_954);
or U2576 (N_2576,In_838,In_684);
and U2577 (N_2577,In_523,In_198);
nand U2578 (N_2578,In_356,In_878);
or U2579 (N_2579,In_995,In_176);
or U2580 (N_2580,In_891,In_959);
and U2581 (N_2581,In_430,In_720);
or U2582 (N_2582,In_664,In_880);
nor U2583 (N_2583,In_340,In_97);
nand U2584 (N_2584,In_179,In_677);
nand U2585 (N_2585,In_390,In_614);
and U2586 (N_2586,In_179,In_401);
or U2587 (N_2587,In_416,In_7);
nand U2588 (N_2588,In_858,In_651);
nand U2589 (N_2589,In_66,In_445);
xnor U2590 (N_2590,In_686,In_832);
nor U2591 (N_2591,In_776,In_13);
and U2592 (N_2592,In_850,In_23);
nand U2593 (N_2593,In_631,In_933);
nor U2594 (N_2594,In_553,In_783);
or U2595 (N_2595,In_464,In_736);
nand U2596 (N_2596,In_817,In_772);
nand U2597 (N_2597,In_495,In_334);
and U2598 (N_2598,In_653,In_509);
and U2599 (N_2599,In_597,In_178);
or U2600 (N_2600,In_0,In_184);
nor U2601 (N_2601,In_339,In_611);
nand U2602 (N_2602,In_320,In_518);
and U2603 (N_2603,In_498,In_716);
and U2604 (N_2604,In_162,In_362);
nor U2605 (N_2605,In_933,In_91);
xor U2606 (N_2606,In_992,In_450);
nand U2607 (N_2607,In_459,In_279);
nand U2608 (N_2608,In_754,In_849);
nor U2609 (N_2609,In_859,In_656);
or U2610 (N_2610,In_839,In_61);
and U2611 (N_2611,In_294,In_949);
and U2612 (N_2612,In_470,In_34);
nand U2613 (N_2613,In_14,In_599);
or U2614 (N_2614,In_591,In_928);
nor U2615 (N_2615,In_970,In_41);
and U2616 (N_2616,In_557,In_857);
xnor U2617 (N_2617,In_37,In_915);
nor U2618 (N_2618,In_165,In_576);
or U2619 (N_2619,In_821,In_148);
or U2620 (N_2620,In_877,In_860);
and U2621 (N_2621,In_298,In_331);
xnor U2622 (N_2622,In_318,In_382);
nor U2623 (N_2623,In_22,In_818);
or U2624 (N_2624,In_180,In_330);
nand U2625 (N_2625,In_490,In_131);
nand U2626 (N_2626,In_737,In_128);
nand U2627 (N_2627,In_789,In_990);
nand U2628 (N_2628,In_204,In_587);
nand U2629 (N_2629,In_601,In_606);
nand U2630 (N_2630,In_154,In_462);
or U2631 (N_2631,In_879,In_319);
nor U2632 (N_2632,In_404,In_820);
or U2633 (N_2633,In_689,In_258);
nor U2634 (N_2634,In_913,In_845);
nand U2635 (N_2635,In_85,In_777);
nor U2636 (N_2636,In_699,In_107);
and U2637 (N_2637,In_760,In_450);
nor U2638 (N_2638,In_998,In_350);
and U2639 (N_2639,In_811,In_404);
nand U2640 (N_2640,In_574,In_853);
nand U2641 (N_2641,In_59,In_204);
and U2642 (N_2642,In_144,In_350);
nand U2643 (N_2643,In_233,In_491);
xor U2644 (N_2644,In_227,In_319);
or U2645 (N_2645,In_254,In_658);
nor U2646 (N_2646,In_75,In_885);
or U2647 (N_2647,In_283,In_951);
or U2648 (N_2648,In_603,In_583);
or U2649 (N_2649,In_983,In_453);
or U2650 (N_2650,In_66,In_313);
and U2651 (N_2651,In_287,In_616);
nor U2652 (N_2652,In_321,In_205);
nand U2653 (N_2653,In_343,In_627);
nor U2654 (N_2654,In_427,In_444);
or U2655 (N_2655,In_302,In_543);
or U2656 (N_2656,In_516,In_239);
nand U2657 (N_2657,In_335,In_78);
or U2658 (N_2658,In_451,In_798);
and U2659 (N_2659,In_564,In_760);
and U2660 (N_2660,In_245,In_589);
and U2661 (N_2661,In_880,In_596);
nor U2662 (N_2662,In_780,In_812);
nor U2663 (N_2663,In_281,In_583);
nor U2664 (N_2664,In_864,In_844);
nor U2665 (N_2665,In_728,In_315);
and U2666 (N_2666,In_210,In_643);
xnor U2667 (N_2667,In_347,In_499);
and U2668 (N_2668,In_841,In_274);
xnor U2669 (N_2669,In_381,In_127);
or U2670 (N_2670,In_3,In_69);
xnor U2671 (N_2671,In_219,In_483);
nor U2672 (N_2672,In_540,In_340);
or U2673 (N_2673,In_715,In_170);
or U2674 (N_2674,In_134,In_486);
nor U2675 (N_2675,In_888,In_877);
and U2676 (N_2676,In_685,In_373);
nand U2677 (N_2677,In_83,In_707);
nor U2678 (N_2678,In_804,In_744);
nand U2679 (N_2679,In_179,In_74);
nor U2680 (N_2680,In_181,In_184);
nor U2681 (N_2681,In_298,In_136);
and U2682 (N_2682,In_676,In_333);
nor U2683 (N_2683,In_919,In_326);
and U2684 (N_2684,In_618,In_114);
nand U2685 (N_2685,In_634,In_862);
or U2686 (N_2686,In_465,In_807);
nand U2687 (N_2687,In_594,In_19);
nand U2688 (N_2688,In_498,In_152);
or U2689 (N_2689,In_740,In_559);
and U2690 (N_2690,In_234,In_282);
and U2691 (N_2691,In_710,In_181);
nor U2692 (N_2692,In_637,In_588);
or U2693 (N_2693,In_557,In_539);
nor U2694 (N_2694,In_313,In_31);
nor U2695 (N_2695,In_161,In_413);
nand U2696 (N_2696,In_160,In_929);
or U2697 (N_2697,In_310,In_154);
and U2698 (N_2698,In_338,In_546);
and U2699 (N_2699,In_403,In_246);
or U2700 (N_2700,In_705,In_578);
xor U2701 (N_2701,In_178,In_260);
or U2702 (N_2702,In_801,In_607);
xnor U2703 (N_2703,In_968,In_822);
nand U2704 (N_2704,In_929,In_8);
nand U2705 (N_2705,In_898,In_700);
and U2706 (N_2706,In_677,In_405);
and U2707 (N_2707,In_84,In_78);
and U2708 (N_2708,In_254,In_123);
nor U2709 (N_2709,In_917,In_985);
nand U2710 (N_2710,In_158,In_972);
and U2711 (N_2711,In_101,In_191);
and U2712 (N_2712,In_221,In_749);
nor U2713 (N_2713,In_475,In_869);
nor U2714 (N_2714,In_453,In_303);
xor U2715 (N_2715,In_888,In_441);
and U2716 (N_2716,In_108,In_246);
nor U2717 (N_2717,In_965,In_495);
nand U2718 (N_2718,In_593,In_207);
xnor U2719 (N_2719,In_313,In_666);
and U2720 (N_2720,In_324,In_975);
nor U2721 (N_2721,In_893,In_851);
xor U2722 (N_2722,In_752,In_475);
nor U2723 (N_2723,In_890,In_382);
nand U2724 (N_2724,In_471,In_713);
nand U2725 (N_2725,In_758,In_859);
and U2726 (N_2726,In_293,In_481);
nor U2727 (N_2727,In_711,In_767);
and U2728 (N_2728,In_4,In_529);
and U2729 (N_2729,In_863,In_443);
nor U2730 (N_2730,In_270,In_95);
and U2731 (N_2731,In_262,In_171);
nand U2732 (N_2732,In_714,In_654);
xor U2733 (N_2733,In_579,In_373);
xnor U2734 (N_2734,In_958,In_518);
and U2735 (N_2735,In_63,In_685);
nor U2736 (N_2736,In_944,In_276);
and U2737 (N_2737,In_622,In_719);
nor U2738 (N_2738,In_530,In_293);
xor U2739 (N_2739,In_98,In_227);
or U2740 (N_2740,In_344,In_783);
nand U2741 (N_2741,In_278,In_553);
and U2742 (N_2742,In_22,In_257);
or U2743 (N_2743,In_613,In_417);
or U2744 (N_2744,In_156,In_334);
xor U2745 (N_2745,In_49,In_350);
nor U2746 (N_2746,In_605,In_79);
or U2747 (N_2747,In_305,In_23);
nor U2748 (N_2748,In_512,In_835);
and U2749 (N_2749,In_253,In_855);
nand U2750 (N_2750,In_957,In_5);
nand U2751 (N_2751,In_354,In_346);
and U2752 (N_2752,In_120,In_381);
nor U2753 (N_2753,In_145,In_228);
and U2754 (N_2754,In_868,In_709);
nand U2755 (N_2755,In_860,In_714);
or U2756 (N_2756,In_550,In_40);
nor U2757 (N_2757,In_787,In_427);
nand U2758 (N_2758,In_611,In_251);
nand U2759 (N_2759,In_8,In_985);
nand U2760 (N_2760,In_330,In_646);
nand U2761 (N_2761,In_821,In_401);
or U2762 (N_2762,In_702,In_603);
and U2763 (N_2763,In_522,In_226);
nand U2764 (N_2764,In_351,In_992);
nor U2765 (N_2765,In_920,In_571);
nor U2766 (N_2766,In_403,In_278);
or U2767 (N_2767,In_983,In_744);
xor U2768 (N_2768,In_475,In_973);
and U2769 (N_2769,In_993,In_119);
nor U2770 (N_2770,In_355,In_633);
xnor U2771 (N_2771,In_721,In_69);
and U2772 (N_2772,In_494,In_567);
and U2773 (N_2773,In_468,In_658);
or U2774 (N_2774,In_14,In_6);
or U2775 (N_2775,In_748,In_977);
and U2776 (N_2776,In_551,In_501);
nor U2777 (N_2777,In_62,In_510);
nand U2778 (N_2778,In_690,In_891);
and U2779 (N_2779,In_302,In_862);
and U2780 (N_2780,In_474,In_863);
nand U2781 (N_2781,In_391,In_410);
and U2782 (N_2782,In_633,In_899);
nor U2783 (N_2783,In_762,In_622);
and U2784 (N_2784,In_101,In_333);
or U2785 (N_2785,In_552,In_984);
or U2786 (N_2786,In_401,In_12);
nand U2787 (N_2787,In_480,In_501);
nor U2788 (N_2788,In_226,In_78);
nor U2789 (N_2789,In_526,In_521);
nor U2790 (N_2790,In_348,In_195);
or U2791 (N_2791,In_721,In_382);
or U2792 (N_2792,In_845,In_3);
nand U2793 (N_2793,In_2,In_609);
and U2794 (N_2794,In_685,In_481);
or U2795 (N_2795,In_626,In_771);
and U2796 (N_2796,In_103,In_462);
nand U2797 (N_2797,In_403,In_834);
or U2798 (N_2798,In_201,In_667);
xor U2799 (N_2799,In_797,In_881);
or U2800 (N_2800,In_444,In_509);
or U2801 (N_2801,In_544,In_521);
nor U2802 (N_2802,In_568,In_907);
nor U2803 (N_2803,In_32,In_656);
and U2804 (N_2804,In_321,In_143);
nor U2805 (N_2805,In_521,In_794);
or U2806 (N_2806,In_449,In_751);
nor U2807 (N_2807,In_980,In_643);
and U2808 (N_2808,In_270,In_463);
nor U2809 (N_2809,In_701,In_63);
nor U2810 (N_2810,In_652,In_837);
or U2811 (N_2811,In_20,In_468);
nand U2812 (N_2812,In_305,In_274);
nor U2813 (N_2813,In_398,In_731);
nand U2814 (N_2814,In_795,In_961);
and U2815 (N_2815,In_433,In_598);
and U2816 (N_2816,In_834,In_780);
and U2817 (N_2817,In_922,In_421);
nor U2818 (N_2818,In_84,In_306);
or U2819 (N_2819,In_843,In_628);
nand U2820 (N_2820,In_255,In_596);
xnor U2821 (N_2821,In_392,In_63);
nor U2822 (N_2822,In_728,In_554);
or U2823 (N_2823,In_100,In_278);
or U2824 (N_2824,In_887,In_3);
nand U2825 (N_2825,In_63,In_697);
and U2826 (N_2826,In_491,In_157);
nand U2827 (N_2827,In_741,In_65);
or U2828 (N_2828,In_320,In_321);
nand U2829 (N_2829,In_715,In_786);
nand U2830 (N_2830,In_251,In_499);
nand U2831 (N_2831,In_747,In_967);
and U2832 (N_2832,In_114,In_734);
nor U2833 (N_2833,In_484,In_780);
nor U2834 (N_2834,In_155,In_269);
or U2835 (N_2835,In_664,In_184);
or U2836 (N_2836,In_182,In_278);
nand U2837 (N_2837,In_379,In_452);
nor U2838 (N_2838,In_128,In_442);
and U2839 (N_2839,In_867,In_627);
nor U2840 (N_2840,In_681,In_256);
nor U2841 (N_2841,In_964,In_110);
xor U2842 (N_2842,In_261,In_952);
or U2843 (N_2843,In_348,In_521);
or U2844 (N_2844,In_245,In_71);
nand U2845 (N_2845,In_561,In_964);
nand U2846 (N_2846,In_314,In_472);
and U2847 (N_2847,In_584,In_585);
and U2848 (N_2848,In_928,In_758);
and U2849 (N_2849,In_798,In_608);
nor U2850 (N_2850,In_755,In_925);
or U2851 (N_2851,In_48,In_229);
xnor U2852 (N_2852,In_646,In_949);
nor U2853 (N_2853,In_724,In_337);
and U2854 (N_2854,In_868,In_805);
and U2855 (N_2855,In_828,In_350);
and U2856 (N_2856,In_471,In_628);
nor U2857 (N_2857,In_729,In_649);
nor U2858 (N_2858,In_748,In_881);
and U2859 (N_2859,In_241,In_932);
xnor U2860 (N_2860,In_187,In_519);
nand U2861 (N_2861,In_826,In_405);
nand U2862 (N_2862,In_210,In_462);
and U2863 (N_2863,In_848,In_739);
nor U2864 (N_2864,In_624,In_984);
and U2865 (N_2865,In_702,In_254);
nor U2866 (N_2866,In_737,In_822);
nand U2867 (N_2867,In_565,In_186);
or U2868 (N_2868,In_958,In_413);
nand U2869 (N_2869,In_861,In_926);
and U2870 (N_2870,In_345,In_669);
and U2871 (N_2871,In_484,In_500);
nand U2872 (N_2872,In_336,In_5);
nor U2873 (N_2873,In_858,In_414);
and U2874 (N_2874,In_9,In_709);
xnor U2875 (N_2875,In_931,In_756);
and U2876 (N_2876,In_125,In_788);
and U2877 (N_2877,In_477,In_124);
nor U2878 (N_2878,In_303,In_315);
nand U2879 (N_2879,In_97,In_898);
nand U2880 (N_2880,In_628,In_781);
and U2881 (N_2881,In_320,In_881);
and U2882 (N_2882,In_584,In_908);
nand U2883 (N_2883,In_61,In_511);
nand U2884 (N_2884,In_327,In_271);
or U2885 (N_2885,In_77,In_793);
or U2886 (N_2886,In_291,In_639);
nand U2887 (N_2887,In_194,In_501);
or U2888 (N_2888,In_462,In_957);
or U2889 (N_2889,In_7,In_989);
or U2890 (N_2890,In_73,In_625);
nor U2891 (N_2891,In_73,In_116);
and U2892 (N_2892,In_838,In_863);
nor U2893 (N_2893,In_980,In_234);
xor U2894 (N_2894,In_612,In_475);
nand U2895 (N_2895,In_351,In_622);
or U2896 (N_2896,In_774,In_477);
xnor U2897 (N_2897,In_992,In_225);
or U2898 (N_2898,In_156,In_717);
or U2899 (N_2899,In_361,In_465);
or U2900 (N_2900,In_699,In_538);
xor U2901 (N_2901,In_369,In_143);
nor U2902 (N_2902,In_697,In_291);
and U2903 (N_2903,In_639,In_587);
or U2904 (N_2904,In_486,In_657);
nand U2905 (N_2905,In_188,In_261);
or U2906 (N_2906,In_416,In_260);
nand U2907 (N_2907,In_605,In_237);
nor U2908 (N_2908,In_742,In_700);
or U2909 (N_2909,In_776,In_20);
and U2910 (N_2910,In_303,In_46);
nand U2911 (N_2911,In_78,In_497);
xnor U2912 (N_2912,In_117,In_1);
xnor U2913 (N_2913,In_507,In_156);
nor U2914 (N_2914,In_932,In_940);
or U2915 (N_2915,In_588,In_855);
xor U2916 (N_2916,In_436,In_226);
nand U2917 (N_2917,In_271,In_761);
nand U2918 (N_2918,In_803,In_896);
or U2919 (N_2919,In_24,In_348);
nor U2920 (N_2920,In_104,In_58);
nor U2921 (N_2921,In_298,In_894);
nor U2922 (N_2922,In_143,In_932);
and U2923 (N_2923,In_404,In_74);
or U2924 (N_2924,In_469,In_33);
nand U2925 (N_2925,In_180,In_223);
xnor U2926 (N_2926,In_597,In_595);
nand U2927 (N_2927,In_470,In_995);
nor U2928 (N_2928,In_358,In_85);
nand U2929 (N_2929,In_499,In_586);
xnor U2930 (N_2930,In_848,In_271);
or U2931 (N_2931,In_223,In_984);
or U2932 (N_2932,In_120,In_657);
and U2933 (N_2933,In_764,In_860);
nand U2934 (N_2934,In_838,In_849);
nand U2935 (N_2935,In_600,In_752);
or U2936 (N_2936,In_54,In_860);
and U2937 (N_2937,In_991,In_949);
and U2938 (N_2938,In_872,In_641);
or U2939 (N_2939,In_470,In_287);
and U2940 (N_2940,In_228,In_792);
nand U2941 (N_2941,In_185,In_882);
and U2942 (N_2942,In_825,In_764);
nand U2943 (N_2943,In_627,In_351);
xor U2944 (N_2944,In_238,In_584);
nor U2945 (N_2945,In_346,In_429);
xor U2946 (N_2946,In_958,In_16);
and U2947 (N_2947,In_125,In_15);
nor U2948 (N_2948,In_854,In_817);
nor U2949 (N_2949,In_936,In_145);
nand U2950 (N_2950,In_593,In_371);
or U2951 (N_2951,In_89,In_497);
or U2952 (N_2952,In_108,In_232);
or U2953 (N_2953,In_606,In_944);
and U2954 (N_2954,In_975,In_819);
nand U2955 (N_2955,In_786,In_602);
nor U2956 (N_2956,In_974,In_987);
or U2957 (N_2957,In_237,In_285);
nand U2958 (N_2958,In_264,In_46);
xor U2959 (N_2959,In_303,In_696);
and U2960 (N_2960,In_862,In_88);
or U2961 (N_2961,In_125,In_419);
nand U2962 (N_2962,In_274,In_691);
nand U2963 (N_2963,In_265,In_226);
or U2964 (N_2964,In_440,In_548);
or U2965 (N_2965,In_640,In_115);
or U2966 (N_2966,In_589,In_776);
nand U2967 (N_2967,In_225,In_632);
and U2968 (N_2968,In_205,In_706);
or U2969 (N_2969,In_79,In_640);
nor U2970 (N_2970,In_416,In_784);
or U2971 (N_2971,In_798,In_485);
nor U2972 (N_2972,In_349,In_62);
nand U2973 (N_2973,In_459,In_402);
or U2974 (N_2974,In_446,In_917);
nor U2975 (N_2975,In_118,In_316);
nor U2976 (N_2976,In_414,In_730);
nor U2977 (N_2977,In_477,In_853);
and U2978 (N_2978,In_902,In_71);
nand U2979 (N_2979,In_380,In_423);
nor U2980 (N_2980,In_600,In_897);
nor U2981 (N_2981,In_425,In_458);
or U2982 (N_2982,In_803,In_742);
or U2983 (N_2983,In_430,In_796);
or U2984 (N_2984,In_209,In_564);
and U2985 (N_2985,In_695,In_43);
nand U2986 (N_2986,In_444,In_148);
nand U2987 (N_2987,In_555,In_615);
nor U2988 (N_2988,In_490,In_750);
nand U2989 (N_2989,In_570,In_911);
and U2990 (N_2990,In_174,In_610);
nand U2991 (N_2991,In_286,In_766);
nor U2992 (N_2992,In_196,In_342);
and U2993 (N_2993,In_280,In_540);
nand U2994 (N_2994,In_11,In_576);
xnor U2995 (N_2995,In_933,In_426);
nand U2996 (N_2996,In_785,In_782);
nand U2997 (N_2997,In_703,In_636);
nor U2998 (N_2998,In_851,In_175);
nand U2999 (N_2999,In_79,In_812);
and U3000 (N_3000,In_560,In_678);
and U3001 (N_3001,In_555,In_260);
nand U3002 (N_3002,In_943,In_678);
or U3003 (N_3003,In_735,In_159);
nand U3004 (N_3004,In_956,In_771);
and U3005 (N_3005,In_609,In_272);
xnor U3006 (N_3006,In_94,In_450);
and U3007 (N_3007,In_202,In_850);
nand U3008 (N_3008,In_733,In_561);
nor U3009 (N_3009,In_87,In_345);
and U3010 (N_3010,In_918,In_606);
nand U3011 (N_3011,In_169,In_595);
nand U3012 (N_3012,In_287,In_799);
or U3013 (N_3013,In_761,In_270);
nand U3014 (N_3014,In_569,In_660);
nor U3015 (N_3015,In_831,In_883);
or U3016 (N_3016,In_387,In_840);
nor U3017 (N_3017,In_141,In_181);
or U3018 (N_3018,In_643,In_580);
xor U3019 (N_3019,In_221,In_847);
nor U3020 (N_3020,In_851,In_365);
nand U3021 (N_3021,In_467,In_737);
or U3022 (N_3022,In_814,In_281);
and U3023 (N_3023,In_612,In_604);
or U3024 (N_3024,In_804,In_439);
and U3025 (N_3025,In_806,In_246);
and U3026 (N_3026,In_437,In_900);
and U3027 (N_3027,In_444,In_268);
nand U3028 (N_3028,In_979,In_571);
nor U3029 (N_3029,In_777,In_243);
and U3030 (N_3030,In_518,In_721);
and U3031 (N_3031,In_500,In_422);
or U3032 (N_3032,In_525,In_13);
nor U3033 (N_3033,In_581,In_721);
xor U3034 (N_3034,In_76,In_916);
nand U3035 (N_3035,In_19,In_247);
xor U3036 (N_3036,In_384,In_387);
nor U3037 (N_3037,In_215,In_694);
nand U3038 (N_3038,In_459,In_907);
nor U3039 (N_3039,In_223,In_287);
and U3040 (N_3040,In_604,In_669);
nand U3041 (N_3041,In_767,In_605);
nor U3042 (N_3042,In_813,In_879);
nand U3043 (N_3043,In_674,In_273);
nand U3044 (N_3044,In_361,In_416);
and U3045 (N_3045,In_976,In_504);
nand U3046 (N_3046,In_720,In_790);
nor U3047 (N_3047,In_759,In_132);
or U3048 (N_3048,In_506,In_5);
nor U3049 (N_3049,In_394,In_702);
and U3050 (N_3050,In_656,In_695);
and U3051 (N_3051,In_255,In_872);
and U3052 (N_3052,In_619,In_991);
nand U3053 (N_3053,In_66,In_410);
and U3054 (N_3054,In_223,In_819);
nand U3055 (N_3055,In_799,In_852);
and U3056 (N_3056,In_143,In_844);
nand U3057 (N_3057,In_881,In_223);
nand U3058 (N_3058,In_631,In_454);
and U3059 (N_3059,In_168,In_517);
and U3060 (N_3060,In_533,In_852);
nor U3061 (N_3061,In_319,In_194);
nor U3062 (N_3062,In_507,In_695);
or U3063 (N_3063,In_838,In_873);
or U3064 (N_3064,In_712,In_560);
xnor U3065 (N_3065,In_786,In_744);
nand U3066 (N_3066,In_764,In_474);
or U3067 (N_3067,In_305,In_945);
nand U3068 (N_3068,In_675,In_198);
nand U3069 (N_3069,In_628,In_148);
nor U3070 (N_3070,In_476,In_269);
and U3071 (N_3071,In_479,In_118);
nor U3072 (N_3072,In_464,In_764);
nand U3073 (N_3073,In_203,In_499);
xor U3074 (N_3074,In_31,In_415);
and U3075 (N_3075,In_209,In_788);
and U3076 (N_3076,In_28,In_779);
and U3077 (N_3077,In_927,In_566);
or U3078 (N_3078,In_282,In_417);
nand U3079 (N_3079,In_77,In_832);
nor U3080 (N_3080,In_33,In_864);
nor U3081 (N_3081,In_642,In_542);
nor U3082 (N_3082,In_176,In_946);
nand U3083 (N_3083,In_466,In_944);
nor U3084 (N_3084,In_238,In_734);
or U3085 (N_3085,In_132,In_596);
and U3086 (N_3086,In_341,In_793);
nor U3087 (N_3087,In_32,In_564);
nor U3088 (N_3088,In_714,In_363);
nor U3089 (N_3089,In_50,In_534);
or U3090 (N_3090,In_137,In_779);
nor U3091 (N_3091,In_793,In_352);
xnor U3092 (N_3092,In_134,In_359);
nand U3093 (N_3093,In_414,In_755);
nor U3094 (N_3094,In_677,In_106);
or U3095 (N_3095,In_415,In_498);
xnor U3096 (N_3096,In_885,In_811);
nand U3097 (N_3097,In_730,In_148);
nor U3098 (N_3098,In_254,In_226);
nand U3099 (N_3099,In_667,In_963);
and U3100 (N_3100,In_98,In_818);
nand U3101 (N_3101,In_75,In_898);
or U3102 (N_3102,In_50,In_145);
or U3103 (N_3103,In_422,In_326);
nor U3104 (N_3104,In_348,In_323);
or U3105 (N_3105,In_315,In_434);
nor U3106 (N_3106,In_156,In_984);
and U3107 (N_3107,In_86,In_161);
and U3108 (N_3108,In_978,In_785);
or U3109 (N_3109,In_158,In_791);
or U3110 (N_3110,In_819,In_88);
or U3111 (N_3111,In_471,In_111);
nor U3112 (N_3112,In_261,In_903);
and U3113 (N_3113,In_295,In_951);
xor U3114 (N_3114,In_18,In_515);
nor U3115 (N_3115,In_446,In_339);
xor U3116 (N_3116,In_414,In_974);
or U3117 (N_3117,In_272,In_992);
nand U3118 (N_3118,In_801,In_250);
nor U3119 (N_3119,In_510,In_435);
xnor U3120 (N_3120,In_310,In_984);
or U3121 (N_3121,In_579,In_161);
nor U3122 (N_3122,In_585,In_906);
and U3123 (N_3123,In_519,In_614);
or U3124 (N_3124,In_386,In_577);
nand U3125 (N_3125,In_70,In_656);
nor U3126 (N_3126,In_913,In_458);
and U3127 (N_3127,In_379,In_293);
nand U3128 (N_3128,In_923,In_233);
or U3129 (N_3129,In_681,In_707);
nor U3130 (N_3130,In_93,In_993);
and U3131 (N_3131,In_657,In_835);
and U3132 (N_3132,In_523,In_744);
nand U3133 (N_3133,In_761,In_409);
xnor U3134 (N_3134,In_591,In_710);
and U3135 (N_3135,In_55,In_799);
nand U3136 (N_3136,In_531,In_734);
nand U3137 (N_3137,In_222,In_602);
and U3138 (N_3138,In_904,In_749);
and U3139 (N_3139,In_897,In_529);
or U3140 (N_3140,In_18,In_600);
and U3141 (N_3141,In_212,In_12);
nand U3142 (N_3142,In_468,In_724);
nor U3143 (N_3143,In_123,In_853);
nor U3144 (N_3144,In_614,In_992);
nand U3145 (N_3145,In_934,In_265);
nor U3146 (N_3146,In_825,In_106);
and U3147 (N_3147,In_520,In_337);
nand U3148 (N_3148,In_542,In_582);
nand U3149 (N_3149,In_519,In_707);
and U3150 (N_3150,In_501,In_914);
nand U3151 (N_3151,In_809,In_201);
and U3152 (N_3152,In_956,In_698);
and U3153 (N_3153,In_727,In_813);
and U3154 (N_3154,In_993,In_903);
xnor U3155 (N_3155,In_653,In_457);
nor U3156 (N_3156,In_545,In_637);
nor U3157 (N_3157,In_353,In_482);
and U3158 (N_3158,In_739,In_752);
or U3159 (N_3159,In_446,In_186);
nand U3160 (N_3160,In_676,In_663);
and U3161 (N_3161,In_581,In_406);
nand U3162 (N_3162,In_328,In_86);
and U3163 (N_3163,In_551,In_123);
or U3164 (N_3164,In_770,In_321);
xor U3165 (N_3165,In_731,In_72);
nor U3166 (N_3166,In_458,In_927);
nand U3167 (N_3167,In_815,In_84);
nor U3168 (N_3168,In_936,In_340);
and U3169 (N_3169,In_806,In_336);
nor U3170 (N_3170,In_879,In_427);
and U3171 (N_3171,In_446,In_823);
nand U3172 (N_3172,In_483,In_878);
nand U3173 (N_3173,In_458,In_821);
xnor U3174 (N_3174,In_484,In_651);
nand U3175 (N_3175,In_282,In_63);
or U3176 (N_3176,In_842,In_454);
or U3177 (N_3177,In_913,In_54);
nand U3178 (N_3178,In_266,In_585);
or U3179 (N_3179,In_836,In_743);
xnor U3180 (N_3180,In_492,In_925);
and U3181 (N_3181,In_795,In_879);
or U3182 (N_3182,In_849,In_832);
nand U3183 (N_3183,In_843,In_146);
nor U3184 (N_3184,In_842,In_156);
xnor U3185 (N_3185,In_606,In_271);
nand U3186 (N_3186,In_941,In_11);
nor U3187 (N_3187,In_738,In_322);
nor U3188 (N_3188,In_659,In_821);
nand U3189 (N_3189,In_639,In_471);
or U3190 (N_3190,In_531,In_478);
nand U3191 (N_3191,In_777,In_425);
or U3192 (N_3192,In_307,In_562);
and U3193 (N_3193,In_597,In_10);
nand U3194 (N_3194,In_570,In_63);
nand U3195 (N_3195,In_112,In_440);
nor U3196 (N_3196,In_713,In_77);
nand U3197 (N_3197,In_55,In_586);
nor U3198 (N_3198,In_445,In_590);
and U3199 (N_3199,In_928,In_318);
nand U3200 (N_3200,In_111,In_110);
nor U3201 (N_3201,In_105,In_560);
and U3202 (N_3202,In_823,In_820);
nor U3203 (N_3203,In_54,In_29);
nor U3204 (N_3204,In_794,In_749);
nor U3205 (N_3205,In_817,In_312);
and U3206 (N_3206,In_743,In_887);
and U3207 (N_3207,In_175,In_422);
or U3208 (N_3208,In_892,In_656);
xnor U3209 (N_3209,In_3,In_584);
xor U3210 (N_3210,In_366,In_215);
and U3211 (N_3211,In_611,In_489);
or U3212 (N_3212,In_159,In_418);
nor U3213 (N_3213,In_19,In_987);
nor U3214 (N_3214,In_801,In_497);
and U3215 (N_3215,In_710,In_267);
and U3216 (N_3216,In_905,In_598);
nand U3217 (N_3217,In_381,In_926);
nor U3218 (N_3218,In_610,In_46);
xor U3219 (N_3219,In_211,In_812);
nand U3220 (N_3220,In_298,In_458);
nor U3221 (N_3221,In_466,In_885);
and U3222 (N_3222,In_293,In_438);
nor U3223 (N_3223,In_522,In_812);
nor U3224 (N_3224,In_137,In_925);
or U3225 (N_3225,In_575,In_89);
and U3226 (N_3226,In_973,In_920);
or U3227 (N_3227,In_454,In_473);
nand U3228 (N_3228,In_286,In_476);
nor U3229 (N_3229,In_947,In_227);
nor U3230 (N_3230,In_902,In_471);
or U3231 (N_3231,In_646,In_976);
nand U3232 (N_3232,In_705,In_481);
or U3233 (N_3233,In_74,In_794);
nor U3234 (N_3234,In_24,In_712);
nor U3235 (N_3235,In_701,In_453);
or U3236 (N_3236,In_819,In_502);
xnor U3237 (N_3237,In_688,In_155);
nor U3238 (N_3238,In_745,In_911);
or U3239 (N_3239,In_690,In_464);
and U3240 (N_3240,In_641,In_103);
nand U3241 (N_3241,In_781,In_789);
or U3242 (N_3242,In_843,In_138);
and U3243 (N_3243,In_981,In_492);
xor U3244 (N_3244,In_897,In_321);
nor U3245 (N_3245,In_828,In_897);
nand U3246 (N_3246,In_963,In_437);
xnor U3247 (N_3247,In_886,In_371);
xnor U3248 (N_3248,In_630,In_234);
xor U3249 (N_3249,In_280,In_74);
nor U3250 (N_3250,In_356,In_848);
nor U3251 (N_3251,In_738,In_469);
or U3252 (N_3252,In_455,In_231);
and U3253 (N_3253,In_600,In_997);
nand U3254 (N_3254,In_44,In_776);
and U3255 (N_3255,In_543,In_626);
or U3256 (N_3256,In_627,In_575);
nor U3257 (N_3257,In_359,In_363);
or U3258 (N_3258,In_370,In_123);
nor U3259 (N_3259,In_790,In_39);
or U3260 (N_3260,In_62,In_571);
or U3261 (N_3261,In_744,In_392);
nand U3262 (N_3262,In_735,In_9);
nand U3263 (N_3263,In_879,In_947);
or U3264 (N_3264,In_570,In_210);
nand U3265 (N_3265,In_634,In_256);
and U3266 (N_3266,In_350,In_854);
nor U3267 (N_3267,In_661,In_349);
and U3268 (N_3268,In_437,In_336);
nor U3269 (N_3269,In_264,In_895);
or U3270 (N_3270,In_251,In_767);
nor U3271 (N_3271,In_999,In_373);
nand U3272 (N_3272,In_769,In_489);
nor U3273 (N_3273,In_313,In_941);
xor U3274 (N_3274,In_812,In_125);
and U3275 (N_3275,In_275,In_264);
nand U3276 (N_3276,In_884,In_395);
and U3277 (N_3277,In_672,In_83);
nand U3278 (N_3278,In_161,In_813);
or U3279 (N_3279,In_788,In_318);
nand U3280 (N_3280,In_676,In_53);
or U3281 (N_3281,In_791,In_943);
nand U3282 (N_3282,In_620,In_734);
nand U3283 (N_3283,In_721,In_861);
xor U3284 (N_3284,In_756,In_244);
and U3285 (N_3285,In_924,In_972);
nor U3286 (N_3286,In_440,In_666);
or U3287 (N_3287,In_581,In_462);
nor U3288 (N_3288,In_67,In_601);
nand U3289 (N_3289,In_955,In_879);
and U3290 (N_3290,In_326,In_215);
or U3291 (N_3291,In_385,In_262);
or U3292 (N_3292,In_95,In_848);
or U3293 (N_3293,In_520,In_958);
or U3294 (N_3294,In_900,In_63);
nor U3295 (N_3295,In_629,In_791);
nand U3296 (N_3296,In_824,In_816);
nor U3297 (N_3297,In_932,In_934);
nand U3298 (N_3298,In_940,In_632);
nand U3299 (N_3299,In_186,In_308);
nor U3300 (N_3300,In_795,In_446);
xor U3301 (N_3301,In_85,In_441);
nand U3302 (N_3302,In_149,In_889);
nand U3303 (N_3303,In_852,In_939);
or U3304 (N_3304,In_793,In_493);
nor U3305 (N_3305,In_717,In_774);
and U3306 (N_3306,In_399,In_167);
and U3307 (N_3307,In_424,In_522);
nor U3308 (N_3308,In_352,In_330);
or U3309 (N_3309,In_329,In_55);
or U3310 (N_3310,In_788,In_133);
or U3311 (N_3311,In_247,In_923);
and U3312 (N_3312,In_960,In_569);
nor U3313 (N_3313,In_977,In_156);
and U3314 (N_3314,In_486,In_823);
xnor U3315 (N_3315,In_121,In_300);
nand U3316 (N_3316,In_577,In_345);
and U3317 (N_3317,In_377,In_423);
nand U3318 (N_3318,In_410,In_22);
or U3319 (N_3319,In_333,In_923);
and U3320 (N_3320,In_949,In_524);
and U3321 (N_3321,In_419,In_409);
nand U3322 (N_3322,In_570,In_669);
nand U3323 (N_3323,In_809,In_189);
nor U3324 (N_3324,In_528,In_521);
nor U3325 (N_3325,In_417,In_564);
or U3326 (N_3326,In_505,In_172);
and U3327 (N_3327,In_451,In_265);
or U3328 (N_3328,In_321,In_237);
or U3329 (N_3329,In_623,In_448);
and U3330 (N_3330,In_774,In_248);
nand U3331 (N_3331,In_773,In_988);
xnor U3332 (N_3332,In_500,In_25);
and U3333 (N_3333,In_328,In_111);
nand U3334 (N_3334,In_236,In_981);
or U3335 (N_3335,In_529,In_902);
and U3336 (N_3336,In_440,In_252);
xnor U3337 (N_3337,In_104,In_824);
or U3338 (N_3338,In_579,In_63);
xor U3339 (N_3339,In_50,In_726);
and U3340 (N_3340,In_945,In_882);
and U3341 (N_3341,In_813,In_910);
nor U3342 (N_3342,In_781,In_209);
or U3343 (N_3343,In_410,In_737);
nand U3344 (N_3344,In_956,In_723);
or U3345 (N_3345,In_968,In_399);
nor U3346 (N_3346,In_456,In_165);
and U3347 (N_3347,In_732,In_615);
nor U3348 (N_3348,In_949,In_195);
nand U3349 (N_3349,In_60,In_965);
and U3350 (N_3350,In_177,In_329);
and U3351 (N_3351,In_839,In_722);
nand U3352 (N_3352,In_589,In_913);
and U3353 (N_3353,In_613,In_450);
xnor U3354 (N_3354,In_382,In_662);
nor U3355 (N_3355,In_897,In_282);
nand U3356 (N_3356,In_349,In_387);
nor U3357 (N_3357,In_449,In_585);
and U3358 (N_3358,In_2,In_9);
nand U3359 (N_3359,In_547,In_175);
or U3360 (N_3360,In_939,In_343);
and U3361 (N_3361,In_647,In_282);
or U3362 (N_3362,In_2,In_275);
nor U3363 (N_3363,In_247,In_209);
nor U3364 (N_3364,In_459,In_390);
nand U3365 (N_3365,In_811,In_974);
nand U3366 (N_3366,In_677,In_899);
nor U3367 (N_3367,In_347,In_844);
nand U3368 (N_3368,In_786,In_107);
or U3369 (N_3369,In_837,In_655);
xor U3370 (N_3370,In_640,In_488);
nor U3371 (N_3371,In_902,In_603);
nand U3372 (N_3372,In_428,In_572);
nor U3373 (N_3373,In_451,In_186);
and U3374 (N_3374,In_507,In_740);
xnor U3375 (N_3375,In_249,In_587);
nor U3376 (N_3376,In_283,In_490);
nor U3377 (N_3377,In_673,In_632);
and U3378 (N_3378,In_517,In_100);
or U3379 (N_3379,In_683,In_612);
or U3380 (N_3380,In_968,In_565);
or U3381 (N_3381,In_328,In_725);
nor U3382 (N_3382,In_817,In_140);
xor U3383 (N_3383,In_394,In_774);
nand U3384 (N_3384,In_273,In_650);
or U3385 (N_3385,In_340,In_72);
and U3386 (N_3386,In_689,In_607);
and U3387 (N_3387,In_70,In_442);
xnor U3388 (N_3388,In_656,In_503);
or U3389 (N_3389,In_82,In_916);
or U3390 (N_3390,In_54,In_191);
and U3391 (N_3391,In_395,In_904);
or U3392 (N_3392,In_136,In_578);
or U3393 (N_3393,In_830,In_792);
xor U3394 (N_3394,In_905,In_311);
nand U3395 (N_3395,In_678,In_732);
and U3396 (N_3396,In_482,In_701);
nor U3397 (N_3397,In_390,In_262);
nand U3398 (N_3398,In_10,In_305);
and U3399 (N_3399,In_554,In_335);
or U3400 (N_3400,In_354,In_719);
or U3401 (N_3401,In_482,In_355);
xor U3402 (N_3402,In_145,In_749);
and U3403 (N_3403,In_455,In_336);
and U3404 (N_3404,In_266,In_674);
or U3405 (N_3405,In_954,In_257);
or U3406 (N_3406,In_887,In_524);
and U3407 (N_3407,In_907,In_927);
and U3408 (N_3408,In_234,In_309);
or U3409 (N_3409,In_440,In_712);
nor U3410 (N_3410,In_306,In_972);
nor U3411 (N_3411,In_396,In_632);
nor U3412 (N_3412,In_190,In_378);
or U3413 (N_3413,In_720,In_496);
xnor U3414 (N_3414,In_479,In_793);
and U3415 (N_3415,In_373,In_87);
nor U3416 (N_3416,In_963,In_567);
nand U3417 (N_3417,In_917,In_188);
or U3418 (N_3418,In_758,In_441);
nor U3419 (N_3419,In_298,In_299);
nand U3420 (N_3420,In_933,In_993);
nor U3421 (N_3421,In_450,In_835);
or U3422 (N_3422,In_795,In_303);
or U3423 (N_3423,In_724,In_532);
nand U3424 (N_3424,In_150,In_33);
and U3425 (N_3425,In_254,In_109);
nand U3426 (N_3426,In_76,In_427);
and U3427 (N_3427,In_19,In_796);
nand U3428 (N_3428,In_600,In_549);
or U3429 (N_3429,In_525,In_732);
and U3430 (N_3430,In_968,In_514);
nor U3431 (N_3431,In_619,In_290);
nand U3432 (N_3432,In_110,In_125);
and U3433 (N_3433,In_932,In_330);
nand U3434 (N_3434,In_597,In_420);
and U3435 (N_3435,In_206,In_222);
nor U3436 (N_3436,In_489,In_227);
xor U3437 (N_3437,In_197,In_150);
or U3438 (N_3438,In_713,In_187);
nor U3439 (N_3439,In_366,In_698);
nor U3440 (N_3440,In_761,In_88);
nand U3441 (N_3441,In_641,In_826);
nand U3442 (N_3442,In_31,In_183);
nand U3443 (N_3443,In_639,In_195);
xnor U3444 (N_3444,In_866,In_980);
or U3445 (N_3445,In_817,In_922);
or U3446 (N_3446,In_844,In_842);
xor U3447 (N_3447,In_814,In_277);
nor U3448 (N_3448,In_529,In_483);
nor U3449 (N_3449,In_137,In_749);
nor U3450 (N_3450,In_368,In_975);
or U3451 (N_3451,In_928,In_844);
and U3452 (N_3452,In_804,In_55);
nor U3453 (N_3453,In_891,In_172);
and U3454 (N_3454,In_537,In_954);
nor U3455 (N_3455,In_124,In_770);
nand U3456 (N_3456,In_51,In_399);
nor U3457 (N_3457,In_458,In_263);
or U3458 (N_3458,In_736,In_818);
nor U3459 (N_3459,In_525,In_567);
nor U3460 (N_3460,In_681,In_88);
nand U3461 (N_3461,In_877,In_541);
nand U3462 (N_3462,In_528,In_187);
and U3463 (N_3463,In_21,In_677);
nor U3464 (N_3464,In_485,In_285);
and U3465 (N_3465,In_105,In_397);
nand U3466 (N_3466,In_92,In_660);
nor U3467 (N_3467,In_12,In_315);
and U3468 (N_3468,In_893,In_527);
nand U3469 (N_3469,In_877,In_906);
and U3470 (N_3470,In_213,In_951);
xnor U3471 (N_3471,In_628,In_211);
nor U3472 (N_3472,In_5,In_147);
and U3473 (N_3473,In_67,In_183);
nand U3474 (N_3474,In_761,In_834);
xor U3475 (N_3475,In_586,In_152);
and U3476 (N_3476,In_912,In_658);
xnor U3477 (N_3477,In_123,In_331);
nor U3478 (N_3478,In_280,In_32);
nor U3479 (N_3479,In_481,In_393);
nand U3480 (N_3480,In_623,In_716);
nor U3481 (N_3481,In_482,In_236);
and U3482 (N_3482,In_265,In_931);
nand U3483 (N_3483,In_520,In_430);
xor U3484 (N_3484,In_497,In_667);
nand U3485 (N_3485,In_464,In_368);
nand U3486 (N_3486,In_264,In_811);
or U3487 (N_3487,In_387,In_951);
nor U3488 (N_3488,In_883,In_157);
nand U3489 (N_3489,In_183,In_710);
xnor U3490 (N_3490,In_384,In_143);
nand U3491 (N_3491,In_722,In_940);
nand U3492 (N_3492,In_687,In_391);
nor U3493 (N_3493,In_442,In_513);
xor U3494 (N_3494,In_378,In_110);
xnor U3495 (N_3495,In_696,In_74);
nor U3496 (N_3496,In_299,In_936);
nand U3497 (N_3497,In_644,In_324);
nor U3498 (N_3498,In_371,In_432);
nor U3499 (N_3499,In_874,In_201);
or U3500 (N_3500,In_914,In_703);
or U3501 (N_3501,In_191,In_832);
or U3502 (N_3502,In_148,In_700);
and U3503 (N_3503,In_655,In_463);
nor U3504 (N_3504,In_459,In_269);
nand U3505 (N_3505,In_446,In_278);
nand U3506 (N_3506,In_166,In_704);
and U3507 (N_3507,In_421,In_205);
or U3508 (N_3508,In_100,In_426);
nand U3509 (N_3509,In_537,In_206);
nor U3510 (N_3510,In_66,In_550);
nand U3511 (N_3511,In_788,In_434);
or U3512 (N_3512,In_79,In_619);
nand U3513 (N_3513,In_203,In_373);
and U3514 (N_3514,In_196,In_635);
and U3515 (N_3515,In_423,In_103);
nand U3516 (N_3516,In_297,In_41);
xnor U3517 (N_3517,In_378,In_66);
or U3518 (N_3518,In_916,In_275);
xor U3519 (N_3519,In_518,In_663);
nor U3520 (N_3520,In_72,In_379);
xor U3521 (N_3521,In_594,In_630);
nor U3522 (N_3522,In_92,In_716);
and U3523 (N_3523,In_598,In_319);
and U3524 (N_3524,In_291,In_235);
and U3525 (N_3525,In_104,In_589);
nand U3526 (N_3526,In_413,In_942);
or U3527 (N_3527,In_421,In_803);
nor U3528 (N_3528,In_25,In_460);
or U3529 (N_3529,In_975,In_286);
xor U3530 (N_3530,In_817,In_409);
nor U3531 (N_3531,In_106,In_179);
nand U3532 (N_3532,In_151,In_38);
nor U3533 (N_3533,In_892,In_409);
and U3534 (N_3534,In_945,In_606);
nand U3535 (N_3535,In_174,In_88);
or U3536 (N_3536,In_781,In_242);
nand U3537 (N_3537,In_270,In_244);
and U3538 (N_3538,In_423,In_607);
or U3539 (N_3539,In_786,In_476);
and U3540 (N_3540,In_26,In_3);
or U3541 (N_3541,In_664,In_832);
or U3542 (N_3542,In_454,In_622);
xnor U3543 (N_3543,In_929,In_159);
nand U3544 (N_3544,In_839,In_850);
nor U3545 (N_3545,In_489,In_766);
and U3546 (N_3546,In_10,In_977);
and U3547 (N_3547,In_552,In_330);
or U3548 (N_3548,In_166,In_503);
and U3549 (N_3549,In_118,In_984);
nand U3550 (N_3550,In_652,In_190);
nor U3551 (N_3551,In_258,In_598);
and U3552 (N_3552,In_732,In_364);
nor U3553 (N_3553,In_747,In_92);
nand U3554 (N_3554,In_9,In_957);
nand U3555 (N_3555,In_858,In_831);
nor U3556 (N_3556,In_637,In_829);
and U3557 (N_3557,In_331,In_250);
or U3558 (N_3558,In_906,In_304);
xor U3559 (N_3559,In_906,In_927);
nand U3560 (N_3560,In_248,In_67);
and U3561 (N_3561,In_198,In_573);
nor U3562 (N_3562,In_995,In_61);
xor U3563 (N_3563,In_102,In_929);
nand U3564 (N_3564,In_30,In_164);
or U3565 (N_3565,In_132,In_872);
xnor U3566 (N_3566,In_284,In_584);
nor U3567 (N_3567,In_244,In_397);
xnor U3568 (N_3568,In_322,In_651);
and U3569 (N_3569,In_275,In_767);
xor U3570 (N_3570,In_69,In_71);
nand U3571 (N_3571,In_848,In_388);
and U3572 (N_3572,In_577,In_404);
nor U3573 (N_3573,In_128,In_949);
or U3574 (N_3574,In_917,In_391);
nor U3575 (N_3575,In_219,In_190);
and U3576 (N_3576,In_248,In_768);
nor U3577 (N_3577,In_837,In_94);
nand U3578 (N_3578,In_241,In_126);
or U3579 (N_3579,In_393,In_673);
nor U3580 (N_3580,In_580,In_959);
nand U3581 (N_3581,In_38,In_694);
nor U3582 (N_3582,In_511,In_72);
and U3583 (N_3583,In_850,In_771);
or U3584 (N_3584,In_394,In_960);
nor U3585 (N_3585,In_119,In_652);
nand U3586 (N_3586,In_904,In_737);
or U3587 (N_3587,In_556,In_158);
nand U3588 (N_3588,In_908,In_719);
nand U3589 (N_3589,In_994,In_499);
nand U3590 (N_3590,In_554,In_574);
xor U3591 (N_3591,In_4,In_581);
or U3592 (N_3592,In_765,In_67);
and U3593 (N_3593,In_264,In_377);
nor U3594 (N_3594,In_689,In_173);
nand U3595 (N_3595,In_601,In_374);
nor U3596 (N_3596,In_784,In_106);
or U3597 (N_3597,In_74,In_410);
nand U3598 (N_3598,In_196,In_368);
or U3599 (N_3599,In_678,In_120);
nand U3600 (N_3600,In_679,In_39);
nor U3601 (N_3601,In_152,In_488);
and U3602 (N_3602,In_205,In_71);
nand U3603 (N_3603,In_911,In_590);
or U3604 (N_3604,In_855,In_81);
nand U3605 (N_3605,In_609,In_394);
nand U3606 (N_3606,In_866,In_616);
nor U3607 (N_3607,In_919,In_185);
nand U3608 (N_3608,In_9,In_21);
nor U3609 (N_3609,In_897,In_622);
nor U3610 (N_3610,In_690,In_613);
or U3611 (N_3611,In_87,In_663);
and U3612 (N_3612,In_750,In_379);
xor U3613 (N_3613,In_430,In_958);
and U3614 (N_3614,In_636,In_605);
nor U3615 (N_3615,In_8,In_799);
and U3616 (N_3616,In_487,In_147);
xor U3617 (N_3617,In_139,In_124);
nand U3618 (N_3618,In_363,In_691);
nand U3619 (N_3619,In_920,In_175);
or U3620 (N_3620,In_326,In_314);
nand U3621 (N_3621,In_289,In_403);
and U3622 (N_3622,In_202,In_206);
or U3623 (N_3623,In_525,In_161);
nand U3624 (N_3624,In_869,In_670);
xnor U3625 (N_3625,In_116,In_69);
or U3626 (N_3626,In_822,In_977);
nand U3627 (N_3627,In_562,In_448);
and U3628 (N_3628,In_47,In_532);
or U3629 (N_3629,In_766,In_207);
and U3630 (N_3630,In_753,In_940);
nor U3631 (N_3631,In_545,In_679);
or U3632 (N_3632,In_332,In_562);
or U3633 (N_3633,In_958,In_528);
nor U3634 (N_3634,In_290,In_288);
or U3635 (N_3635,In_662,In_747);
and U3636 (N_3636,In_909,In_168);
xor U3637 (N_3637,In_520,In_471);
nand U3638 (N_3638,In_720,In_717);
and U3639 (N_3639,In_903,In_684);
or U3640 (N_3640,In_741,In_421);
or U3641 (N_3641,In_886,In_451);
nor U3642 (N_3642,In_447,In_9);
and U3643 (N_3643,In_975,In_891);
or U3644 (N_3644,In_696,In_803);
or U3645 (N_3645,In_793,In_818);
and U3646 (N_3646,In_927,In_818);
nor U3647 (N_3647,In_130,In_937);
or U3648 (N_3648,In_549,In_99);
nand U3649 (N_3649,In_47,In_997);
nand U3650 (N_3650,In_901,In_878);
or U3651 (N_3651,In_175,In_347);
and U3652 (N_3652,In_928,In_808);
xnor U3653 (N_3653,In_972,In_124);
xor U3654 (N_3654,In_485,In_423);
and U3655 (N_3655,In_553,In_464);
or U3656 (N_3656,In_377,In_841);
nor U3657 (N_3657,In_302,In_23);
nor U3658 (N_3658,In_617,In_414);
nor U3659 (N_3659,In_13,In_703);
and U3660 (N_3660,In_696,In_500);
nand U3661 (N_3661,In_303,In_819);
nor U3662 (N_3662,In_143,In_497);
nand U3663 (N_3663,In_580,In_448);
and U3664 (N_3664,In_341,In_624);
nand U3665 (N_3665,In_277,In_881);
or U3666 (N_3666,In_176,In_102);
nor U3667 (N_3667,In_781,In_353);
nand U3668 (N_3668,In_50,In_819);
or U3669 (N_3669,In_217,In_568);
nand U3670 (N_3670,In_753,In_193);
or U3671 (N_3671,In_491,In_263);
nand U3672 (N_3672,In_272,In_121);
or U3673 (N_3673,In_784,In_868);
or U3674 (N_3674,In_500,In_936);
nor U3675 (N_3675,In_279,In_233);
nor U3676 (N_3676,In_876,In_184);
and U3677 (N_3677,In_709,In_874);
and U3678 (N_3678,In_63,In_652);
nand U3679 (N_3679,In_973,In_914);
or U3680 (N_3680,In_570,In_6);
nor U3681 (N_3681,In_219,In_871);
nand U3682 (N_3682,In_908,In_655);
nor U3683 (N_3683,In_285,In_551);
or U3684 (N_3684,In_125,In_682);
nor U3685 (N_3685,In_660,In_763);
or U3686 (N_3686,In_403,In_882);
nor U3687 (N_3687,In_188,In_170);
and U3688 (N_3688,In_394,In_833);
nor U3689 (N_3689,In_249,In_769);
nand U3690 (N_3690,In_271,In_179);
or U3691 (N_3691,In_645,In_743);
and U3692 (N_3692,In_518,In_20);
or U3693 (N_3693,In_590,In_892);
or U3694 (N_3694,In_601,In_462);
nor U3695 (N_3695,In_599,In_641);
nor U3696 (N_3696,In_335,In_470);
nand U3697 (N_3697,In_825,In_226);
nand U3698 (N_3698,In_50,In_521);
or U3699 (N_3699,In_874,In_999);
nand U3700 (N_3700,In_958,In_473);
and U3701 (N_3701,In_642,In_139);
and U3702 (N_3702,In_191,In_612);
or U3703 (N_3703,In_943,In_919);
and U3704 (N_3704,In_487,In_60);
and U3705 (N_3705,In_617,In_77);
and U3706 (N_3706,In_566,In_3);
nand U3707 (N_3707,In_158,In_565);
nand U3708 (N_3708,In_269,In_223);
and U3709 (N_3709,In_235,In_441);
xnor U3710 (N_3710,In_23,In_35);
or U3711 (N_3711,In_682,In_910);
nor U3712 (N_3712,In_439,In_343);
nand U3713 (N_3713,In_678,In_311);
or U3714 (N_3714,In_585,In_420);
nand U3715 (N_3715,In_315,In_930);
and U3716 (N_3716,In_702,In_163);
and U3717 (N_3717,In_370,In_704);
or U3718 (N_3718,In_584,In_885);
nor U3719 (N_3719,In_675,In_577);
and U3720 (N_3720,In_503,In_552);
nand U3721 (N_3721,In_487,In_844);
or U3722 (N_3722,In_487,In_554);
nor U3723 (N_3723,In_944,In_320);
nor U3724 (N_3724,In_213,In_703);
nand U3725 (N_3725,In_14,In_609);
and U3726 (N_3726,In_549,In_978);
or U3727 (N_3727,In_875,In_910);
nand U3728 (N_3728,In_359,In_262);
and U3729 (N_3729,In_725,In_49);
nand U3730 (N_3730,In_994,In_253);
nand U3731 (N_3731,In_758,In_957);
or U3732 (N_3732,In_889,In_51);
nor U3733 (N_3733,In_736,In_746);
nor U3734 (N_3734,In_952,In_174);
or U3735 (N_3735,In_685,In_148);
xnor U3736 (N_3736,In_461,In_317);
nor U3737 (N_3737,In_187,In_905);
and U3738 (N_3738,In_892,In_108);
and U3739 (N_3739,In_696,In_557);
xnor U3740 (N_3740,In_69,In_685);
xnor U3741 (N_3741,In_603,In_42);
or U3742 (N_3742,In_471,In_92);
nand U3743 (N_3743,In_249,In_879);
or U3744 (N_3744,In_617,In_958);
and U3745 (N_3745,In_533,In_928);
nor U3746 (N_3746,In_152,In_969);
nor U3747 (N_3747,In_698,In_782);
nor U3748 (N_3748,In_724,In_822);
or U3749 (N_3749,In_540,In_213);
and U3750 (N_3750,In_367,In_249);
nand U3751 (N_3751,In_650,In_589);
nor U3752 (N_3752,In_658,In_634);
nand U3753 (N_3753,In_526,In_721);
and U3754 (N_3754,In_181,In_42);
or U3755 (N_3755,In_835,In_775);
nor U3756 (N_3756,In_556,In_552);
or U3757 (N_3757,In_569,In_431);
nor U3758 (N_3758,In_692,In_368);
and U3759 (N_3759,In_670,In_951);
and U3760 (N_3760,In_914,In_864);
nand U3761 (N_3761,In_360,In_60);
or U3762 (N_3762,In_6,In_879);
nor U3763 (N_3763,In_440,In_360);
nor U3764 (N_3764,In_386,In_93);
nor U3765 (N_3765,In_791,In_261);
xnor U3766 (N_3766,In_340,In_877);
or U3767 (N_3767,In_109,In_198);
or U3768 (N_3768,In_36,In_562);
nor U3769 (N_3769,In_4,In_130);
xor U3770 (N_3770,In_440,In_228);
and U3771 (N_3771,In_53,In_330);
and U3772 (N_3772,In_585,In_414);
xnor U3773 (N_3773,In_574,In_681);
and U3774 (N_3774,In_535,In_515);
xnor U3775 (N_3775,In_849,In_693);
xor U3776 (N_3776,In_959,In_41);
nor U3777 (N_3777,In_393,In_614);
and U3778 (N_3778,In_100,In_927);
and U3779 (N_3779,In_906,In_577);
nand U3780 (N_3780,In_368,In_486);
nand U3781 (N_3781,In_747,In_782);
nor U3782 (N_3782,In_850,In_124);
or U3783 (N_3783,In_960,In_41);
and U3784 (N_3784,In_144,In_518);
or U3785 (N_3785,In_659,In_640);
nor U3786 (N_3786,In_264,In_551);
nand U3787 (N_3787,In_556,In_892);
or U3788 (N_3788,In_859,In_781);
nor U3789 (N_3789,In_662,In_720);
and U3790 (N_3790,In_459,In_903);
nor U3791 (N_3791,In_140,In_557);
nor U3792 (N_3792,In_875,In_473);
nand U3793 (N_3793,In_641,In_231);
nor U3794 (N_3794,In_741,In_769);
nor U3795 (N_3795,In_750,In_767);
or U3796 (N_3796,In_979,In_428);
nand U3797 (N_3797,In_609,In_532);
or U3798 (N_3798,In_102,In_788);
xnor U3799 (N_3799,In_971,In_831);
nor U3800 (N_3800,In_144,In_800);
nor U3801 (N_3801,In_846,In_877);
or U3802 (N_3802,In_929,In_41);
and U3803 (N_3803,In_698,In_228);
and U3804 (N_3804,In_888,In_65);
nand U3805 (N_3805,In_324,In_546);
nor U3806 (N_3806,In_506,In_79);
xnor U3807 (N_3807,In_860,In_67);
xnor U3808 (N_3808,In_373,In_175);
or U3809 (N_3809,In_501,In_338);
and U3810 (N_3810,In_536,In_425);
nor U3811 (N_3811,In_901,In_86);
nor U3812 (N_3812,In_563,In_32);
and U3813 (N_3813,In_576,In_665);
or U3814 (N_3814,In_111,In_45);
nor U3815 (N_3815,In_988,In_993);
or U3816 (N_3816,In_211,In_820);
nor U3817 (N_3817,In_550,In_800);
and U3818 (N_3818,In_788,In_373);
and U3819 (N_3819,In_215,In_149);
and U3820 (N_3820,In_221,In_81);
and U3821 (N_3821,In_609,In_504);
or U3822 (N_3822,In_346,In_511);
or U3823 (N_3823,In_455,In_897);
nor U3824 (N_3824,In_256,In_942);
or U3825 (N_3825,In_358,In_355);
nor U3826 (N_3826,In_433,In_226);
nand U3827 (N_3827,In_634,In_229);
xnor U3828 (N_3828,In_385,In_951);
or U3829 (N_3829,In_642,In_673);
and U3830 (N_3830,In_140,In_389);
nor U3831 (N_3831,In_857,In_313);
or U3832 (N_3832,In_820,In_137);
nor U3833 (N_3833,In_88,In_605);
nand U3834 (N_3834,In_806,In_505);
or U3835 (N_3835,In_713,In_806);
xnor U3836 (N_3836,In_365,In_703);
and U3837 (N_3837,In_120,In_439);
nor U3838 (N_3838,In_520,In_448);
or U3839 (N_3839,In_511,In_234);
or U3840 (N_3840,In_745,In_385);
or U3841 (N_3841,In_446,In_246);
and U3842 (N_3842,In_573,In_835);
nor U3843 (N_3843,In_430,In_960);
or U3844 (N_3844,In_610,In_999);
nand U3845 (N_3845,In_863,In_893);
or U3846 (N_3846,In_670,In_311);
and U3847 (N_3847,In_425,In_207);
nor U3848 (N_3848,In_171,In_350);
or U3849 (N_3849,In_75,In_840);
nor U3850 (N_3850,In_964,In_880);
nand U3851 (N_3851,In_21,In_858);
or U3852 (N_3852,In_76,In_578);
and U3853 (N_3853,In_950,In_972);
or U3854 (N_3854,In_502,In_480);
or U3855 (N_3855,In_292,In_990);
nand U3856 (N_3856,In_760,In_811);
nand U3857 (N_3857,In_942,In_861);
xnor U3858 (N_3858,In_532,In_694);
nand U3859 (N_3859,In_383,In_302);
xor U3860 (N_3860,In_22,In_566);
and U3861 (N_3861,In_308,In_469);
nand U3862 (N_3862,In_841,In_157);
and U3863 (N_3863,In_65,In_936);
xnor U3864 (N_3864,In_125,In_982);
or U3865 (N_3865,In_646,In_835);
or U3866 (N_3866,In_455,In_710);
or U3867 (N_3867,In_523,In_504);
nand U3868 (N_3868,In_162,In_815);
nor U3869 (N_3869,In_285,In_790);
nor U3870 (N_3870,In_241,In_349);
and U3871 (N_3871,In_316,In_600);
nor U3872 (N_3872,In_874,In_775);
nor U3873 (N_3873,In_362,In_391);
nor U3874 (N_3874,In_706,In_701);
nand U3875 (N_3875,In_260,In_149);
nor U3876 (N_3876,In_301,In_676);
nor U3877 (N_3877,In_156,In_564);
and U3878 (N_3878,In_658,In_893);
xor U3879 (N_3879,In_89,In_94);
nor U3880 (N_3880,In_893,In_521);
and U3881 (N_3881,In_824,In_20);
nor U3882 (N_3882,In_781,In_951);
or U3883 (N_3883,In_733,In_739);
and U3884 (N_3884,In_687,In_565);
xnor U3885 (N_3885,In_978,In_580);
nor U3886 (N_3886,In_661,In_356);
nand U3887 (N_3887,In_619,In_598);
nor U3888 (N_3888,In_327,In_912);
nor U3889 (N_3889,In_949,In_84);
and U3890 (N_3890,In_908,In_515);
nand U3891 (N_3891,In_217,In_623);
xor U3892 (N_3892,In_989,In_716);
and U3893 (N_3893,In_182,In_571);
or U3894 (N_3894,In_420,In_222);
and U3895 (N_3895,In_38,In_108);
and U3896 (N_3896,In_871,In_24);
or U3897 (N_3897,In_770,In_294);
xnor U3898 (N_3898,In_150,In_525);
and U3899 (N_3899,In_461,In_389);
and U3900 (N_3900,In_636,In_894);
and U3901 (N_3901,In_287,In_61);
and U3902 (N_3902,In_518,In_97);
and U3903 (N_3903,In_556,In_88);
or U3904 (N_3904,In_950,In_724);
or U3905 (N_3905,In_180,In_769);
and U3906 (N_3906,In_265,In_932);
or U3907 (N_3907,In_743,In_446);
nand U3908 (N_3908,In_227,In_300);
nand U3909 (N_3909,In_501,In_363);
or U3910 (N_3910,In_280,In_861);
and U3911 (N_3911,In_505,In_887);
nor U3912 (N_3912,In_3,In_455);
xor U3913 (N_3913,In_217,In_469);
nor U3914 (N_3914,In_246,In_308);
nor U3915 (N_3915,In_258,In_581);
xnor U3916 (N_3916,In_836,In_593);
and U3917 (N_3917,In_957,In_834);
xor U3918 (N_3918,In_962,In_538);
nand U3919 (N_3919,In_370,In_917);
and U3920 (N_3920,In_348,In_0);
nor U3921 (N_3921,In_879,In_389);
nor U3922 (N_3922,In_220,In_819);
or U3923 (N_3923,In_20,In_944);
nand U3924 (N_3924,In_152,In_150);
nand U3925 (N_3925,In_987,In_757);
and U3926 (N_3926,In_871,In_92);
and U3927 (N_3927,In_474,In_0);
or U3928 (N_3928,In_497,In_1);
nor U3929 (N_3929,In_730,In_358);
nor U3930 (N_3930,In_105,In_908);
nor U3931 (N_3931,In_988,In_199);
or U3932 (N_3932,In_720,In_90);
and U3933 (N_3933,In_260,In_335);
nand U3934 (N_3934,In_398,In_810);
nor U3935 (N_3935,In_583,In_699);
nand U3936 (N_3936,In_390,In_941);
and U3937 (N_3937,In_545,In_641);
and U3938 (N_3938,In_942,In_352);
xor U3939 (N_3939,In_461,In_796);
nor U3940 (N_3940,In_826,In_630);
nand U3941 (N_3941,In_994,In_461);
nand U3942 (N_3942,In_282,In_909);
nand U3943 (N_3943,In_467,In_729);
and U3944 (N_3944,In_79,In_693);
and U3945 (N_3945,In_623,In_221);
and U3946 (N_3946,In_402,In_956);
or U3947 (N_3947,In_382,In_588);
nor U3948 (N_3948,In_277,In_87);
or U3949 (N_3949,In_166,In_20);
or U3950 (N_3950,In_574,In_627);
and U3951 (N_3951,In_951,In_195);
and U3952 (N_3952,In_172,In_884);
xnor U3953 (N_3953,In_911,In_86);
and U3954 (N_3954,In_177,In_888);
nor U3955 (N_3955,In_41,In_999);
nor U3956 (N_3956,In_657,In_747);
xor U3957 (N_3957,In_374,In_176);
or U3958 (N_3958,In_364,In_212);
or U3959 (N_3959,In_960,In_551);
or U3960 (N_3960,In_476,In_207);
nor U3961 (N_3961,In_875,In_757);
nor U3962 (N_3962,In_613,In_868);
nand U3963 (N_3963,In_206,In_131);
and U3964 (N_3964,In_812,In_489);
or U3965 (N_3965,In_983,In_133);
nor U3966 (N_3966,In_67,In_923);
nand U3967 (N_3967,In_563,In_822);
and U3968 (N_3968,In_720,In_792);
and U3969 (N_3969,In_137,In_298);
or U3970 (N_3970,In_389,In_235);
nand U3971 (N_3971,In_307,In_673);
or U3972 (N_3972,In_642,In_857);
nor U3973 (N_3973,In_959,In_723);
nand U3974 (N_3974,In_998,In_282);
nor U3975 (N_3975,In_621,In_958);
and U3976 (N_3976,In_768,In_353);
and U3977 (N_3977,In_134,In_982);
nand U3978 (N_3978,In_333,In_195);
nor U3979 (N_3979,In_920,In_610);
nand U3980 (N_3980,In_164,In_826);
and U3981 (N_3981,In_624,In_161);
and U3982 (N_3982,In_333,In_33);
and U3983 (N_3983,In_250,In_374);
and U3984 (N_3984,In_99,In_77);
and U3985 (N_3985,In_777,In_907);
or U3986 (N_3986,In_518,In_710);
nor U3987 (N_3987,In_214,In_318);
and U3988 (N_3988,In_106,In_735);
nand U3989 (N_3989,In_939,In_698);
nor U3990 (N_3990,In_810,In_920);
nand U3991 (N_3991,In_301,In_402);
and U3992 (N_3992,In_198,In_392);
nand U3993 (N_3993,In_779,In_538);
nor U3994 (N_3994,In_688,In_535);
xor U3995 (N_3995,In_811,In_940);
nor U3996 (N_3996,In_939,In_162);
xor U3997 (N_3997,In_431,In_871);
nand U3998 (N_3998,In_231,In_317);
nor U3999 (N_3999,In_465,In_667);
nand U4000 (N_4000,In_881,In_732);
or U4001 (N_4001,In_4,In_108);
and U4002 (N_4002,In_307,In_148);
nand U4003 (N_4003,In_758,In_917);
and U4004 (N_4004,In_495,In_446);
xnor U4005 (N_4005,In_450,In_603);
nor U4006 (N_4006,In_895,In_757);
nor U4007 (N_4007,In_288,In_783);
and U4008 (N_4008,In_618,In_928);
nor U4009 (N_4009,In_731,In_294);
and U4010 (N_4010,In_80,In_47);
and U4011 (N_4011,In_71,In_647);
xor U4012 (N_4012,In_637,In_859);
or U4013 (N_4013,In_484,In_418);
nor U4014 (N_4014,In_974,In_937);
xor U4015 (N_4015,In_595,In_948);
and U4016 (N_4016,In_81,In_242);
and U4017 (N_4017,In_387,In_824);
or U4018 (N_4018,In_112,In_288);
or U4019 (N_4019,In_140,In_78);
nand U4020 (N_4020,In_834,In_749);
or U4021 (N_4021,In_821,In_72);
and U4022 (N_4022,In_867,In_27);
and U4023 (N_4023,In_496,In_409);
and U4024 (N_4024,In_282,In_772);
nor U4025 (N_4025,In_571,In_56);
and U4026 (N_4026,In_433,In_136);
nor U4027 (N_4027,In_887,In_54);
nand U4028 (N_4028,In_535,In_781);
nor U4029 (N_4029,In_503,In_184);
nor U4030 (N_4030,In_202,In_31);
or U4031 (N_4031,In_915,In_941);
nand U4032 (N_4032,In_485,In_287);
or U4033 (N_4033,In_953,In_648);
and U4034 (N_4034,In_530,In_663);
and U4035 (N_4035,In_749,In_972);
or U4036 (N_4036,In_490,In_608);
or U4037 (N_4037,In_457,In_659);
or U4038 (N_4038,In_685,In_639);
or U4039 (N_4039,In_806,In_800);
xnor U4040 (N_4040,In_127,In_318);
and U4041 (N_4041,In_594,In_198);
xnor U4042 (N_4042,In_663,In_463);
nor U4043 (N_4043,In_404,In_843);
and U4044 (N_4044,In_27,In_516);
nor U4045 (N_4045,In_990,In_157);
or U4046 (N_4046,In_985,In_591);
or U4047 (N_4047,In_515,In_54);
nand U4048 (N_4048,In_755,In_628);
or U4049 (N_4049,In_514,In_760);
or U4050 (N_4050,In_384,In_268);
and U4051 (N_4051,In_670,In_828);
nor U4052 (N_4052,In_582,In_602);
and U4053 (N_4053,In_490,In_555);
and U4054 (N_4054,In_46,In_394);
or U4055 (N_4055,In_64,In_234);
nand U4056 (N_4056,In_967,In_427);
and U4057 (N_4057,In_425,In_669);
or U4058 (N_4058,In_984,In_323);
nor U4059 (N_4059,In_317,In_151);
nor U4060 (N_4060,In_714,In_129);
or U4061 (N_4061,In_474,In_262);
nor U4062 (N_4062,In_975,In_865);
nor U4063 (N_4063,In_244,In_748);
nor U4064 (N_4064,In_152,In_454);
nand U4065 (N_4065,In_304,In_918);
or U4066 (N_4066,In_783,In_252);
or U4067 (N_4067,In_453,In_149);
and U4068 (N_4068,In_463,In_244);
and U4069 (N_4069,In_2,In_173);
nand U4070 (N_4070,In_218,In_975);
nor U4071 (N_4071,In_367,In_259);
nand U4072 (N_4072,In_888,In_299);
or U4073 (N_4073,In_549,In_779);
nand U4074 (N_4074,In_524,In_420);
and U4075 (N_4075,In_65,In_865);
and U4076 (N_4076,In_307,In_398);
and U4077 (N_4077,In_593,In_202);
nand U4078 (N_4078,In_40,In_858);
nand U4079 (N_4079,In_653,In_166);
and U4080 (N_4080,In_524,In_20);
nand U4081 (N_4081,In_847,In_165);
nor U4082 (N_4082,In_749,In_82);
nand U4083 (N_4083,In_915,In_826);
and U4084 (N_4084,In_396,In_465);
nand U4085 (N_4085,In_694,In_325);
or U4086 (N_4086,In_417,In_74);
and U4087 (N_4087,In_733,In_983);
and U4088 (N_4088,In_787,In_301);
or U4089 (N_4089,In_117,In_45);
and U4090 (N_4090,In_563,In_29);
nand U4091 (N_4091,In_284,In_889);
nand U4092 (N_4092,In_213,In_555);
nand U4093 (N_4093,In_774,In_351);
and U4094 (N_4094,In_162,In_513);
xor U4095 (N_4095,In_255,In_215);
nor U4096 (N_4096,In_354,In_449);
or U4097 (N_4097,In_187,In_149);
nor U4098 (N_4098,In_516,In_805);
nor U4099 (N_4099,In_523,In_536);
nand U4100 (N_4100,In_948,In_513);
nand U4101 (N_4101,In_6,In_941);
nand U4102 (N_4102,In_787,In_958);
nor U4103 (N_4103,In_967,In_662);
nor U4104 (N_4104,In_818,In_960);
nand U4105 (N_4105,In_276,In_991);
nor U4106 (N_4106,In_874,In_133);
and U4107 (N_4107,In_870,In_268);
and U4108 (N_4108,In_520,In_716);
and U4109 (N_4109,In_121,In_312);
nor U4110 (N_4110,In_218,In_85);
xor U4111 (N_4111,In_816,In_7);
or U4112 (N_4112,In_520,In_892);
nand U4113 (N_4113,In_441,In_682);
and U4114 (N_4114,In_675,In_469);
xnor U4115 (N_4115,In_694,In_194);
or U4116 (N_4116,In_462,In_817);
nor U4117 (N_4117,In_487,In_16);
nand U4118 (N_4118,In_732,In_941);
and U4119 (N_4119,In_402,In_281);
nand U4120 (N_4120,In_232,In_265);
nor U4121 (N_4121,In_942,In_340);
xnor U4122 (N_4122,In_793,In_66);
or U4123 (N_4123,In_555,In_322);
nand U4124 (N_4124,In_7,In_131);
nand U4125 (N_4125,In_765,In_90);
xnor U4126 (N_4126,In_56,In_810);
nand U4127 (N_4127,In_870,In_70);
or U4128 (N_4128,In_397,In_962);
or U4129 (N_4129,In_977,In_519);
nand U4130 (N_4130,In_419,In_49);
or U4131 (N_4131,In_132,In_579);
nor U4132 (N_4132,In_97,In_8);
nor U4133 (N_4133,In_303,In_141);
and U4134 (N_4134,In_860,In_793);
nand U4135 (N_4135,In_385,In_973);
nor U4136 (N_4136,In_770,In_996);
nor U4137 (N_4137,In_796,In_257);
or U4138 (N_4138,In_553,In_737);
or U4139 (N_4139,In_388,In_439);
nand U4140 (N_4140,In_714,In_220);
xnor U4141 (N_4141,In_421,In_806);
nand U4142 (N_4142,In_773,In_787);
nand U4143 (N_4143,In_936,In_960);
nor U4144 (N_4144,In_634,In_271);
and U4145 (N_4145,In_891,In_49);
and U4146 (N_4146,In_313,In_16);
and U4147 (N_4147,In_42,In_798);
or U4148 (N_4148,In_555,In_236);
and U4149 (N_4149,In_903,In_342);
nor U4150 (N_4150,In_543,In_906);
nand U4151 (N_4151,In_278,In_557);
nor U4152 (N_4152,In_218,In_659);
nand U4153 (N_4153,In_503,In_319);
and U4154 (N_4154,In_876,In_742);
nor U4155 (N_4155,In_601,In_545);
nor U4156 (N_4156,In_992,In_799);
nor U4157 (N_4157,In_962,In_148);
nand U4158 (N_4158,In_596,In_402);
and U4159 (N_4159,In_717,In_625);
nand U4160 (N_4160,In_740,In_666);
nor U4161 (N_4161,In_939,In_966);
or U4162 (N_4162,In_645,In_490);
nand U4163 (N_4163,In_15,In_339);
nand U4164 (N_4164,In_287,In_38);
nor U4165 (N_4165,In_898,In_520);
nand U4166 (N_4166,In_792,In_711);
nand U4167 (N_4167,In_749,In_580);
and U4168 (N_4168,In_882,In_775);
xnor U4169 (N_4169,In_904,In_712);
xor U4170 (N_4170,In_134,In_326);
and U4171 (N_4171,In_539,In_408);
nor U4172 (N_4172,In_64,In_152);
xnor U4173 (N_4173,In_413,In_473);
and U4174 (N_4174,In_136,In_606);
xor U4175 (N_4175,In_840,In_578);
or U4176 (N_4176,In_22,In_486);
xnor U4177 (N_4177,In_281,In_379);
nand U4178 (N_4178,In_56,In_766);
nor U4179 (N_4179,In_890,In_583);
and U4180 (N_4180,In_642,In_253);
nor U4181 (N_4181,In_912,In_487);
and U4182 (N_4182,In_910,In_252);
or U4183 (N_4183,In_502,In_630);
and U4184 (N_4184,In_535,In_321);
or U4185 (N_4185,In_103,In_446);
xnor U4186 (N_4186,In_453,In_116);
or U4187 (N_4187,In_189,In_337);
nand U4188 (N_4188,In_502,In_59);
nor U4189 (N_4189,In_512,In_338);
and U4190 (N_4190,In_404,In_809);
or U4191 (N_4191,In_325,In_974);
nor U4192 (N_4192,In_914,In_846);
nand U4193 (N_4193,In_685,In_185);
nand U4194 (N_4194,In_539,In_894);
or U4195 (N_4195,In_260,In_868);
nor U4196 (N_4196,In_77,In_727);
or U4197 (N_4197,In_981,In_469);
nor U4198 (N_4198,In_53,In_138);
nand U4199 (N_4199,In_278,In_449);
and U4200 (N_4200,In_699,In_261);
xnor U4201 (N_4201,In_604,In_506);
or U4202 (N_4202,In_346,In_382);
nor U4203 (N_4203,In_310,In_44);
nor U4204 (N_4204,In_952,In_676);
and U4205 (N_4205,In_128,In_249);
and U4206 (N_4206,In_63,In_553);
nor U4207 (N_4207,In_98,In_836);
nand U4208 (N_4208,In_932,In_46);
nor U4209 (N_4209,In_3,In_377);
or U4210 (N_4210,In_773,In_954);
nor U4211 (N_4211,In_406,In_273);
or U4212 (N_4212,In_794,In_304);
or U4213 (N_4213,In_866,In_930);
nor U4214 (N_4214,In_563,In_615);
and U4215 (N_4215,In_674,In_199);
nand U4216 (N_4216,In_641,In_959);
xor U4217 (N_4217,In_887,In_733);
nor U4218 (N_4218,In_795,In_235);
nand U4219 (N_4219,In_772,In_928);
nand U4220 (N_4220,In_294,In_420);
nor U4221 (N_4221,In_511,In_574);
and U4222 (N_4222,In_971,In_139);
nor U4223 (N_4223,In_638,In_584);
xor U4224 (N_4224,In_805,In_895);
xor U4225 (N_4225,In_487,In_171);
or U4226 (N_4226,In_110,In_429);
nand U4227 (N_4227,In_556,In_849);
or U4228 (N_4228,In_594,In_838);
and U4229 (N_4229,In_43,In_849);
or U4230 (N_4230,In_214,In_452);
or U4231 (N_4231,In_76,In_647);
or U4232 (N_4232,In_507,In_856);
xor U4233 (N_4233,In_363,In_616);
nor U4234 (N_4234,In_396,In_482);
nor U4235 (N_4235,In_938,In_656);
and U4236 (N_4236,In_983,In_944);
nor U4237 (N_4237,In_404,In_992);
nand U4238 (N_4238,In_257,In_11);
nor U4239 (N_4239,In_476,In_564);
nor U4240 (N_4240,In_40,In_973);
nor U4241 (N_4241,In_632,In_375);
nand U4242 (N_4242,In_47,In_211);
or U4243 (N_4243,In_87,In_505);
nand U4244 (N_4244,In_826,In_705);
nor U4245 (N_4245,In_761,In_503);
nor U4246 (N_4246,In_694,In_927);
nor U4247 (N_4247,In_872,In_353);
or U4248 (N_4248,In_23,In_525);
nor U4249 (N_4249,In_330,In_761);
nand U4250 (N_4250,In_795,In_502);
nand U4251 (N_4251,In_831,In_470);
nor U4252 (N_4252,In_148,In_260);
nor U4253 (N_4253,In_39,In_954);
and U4254 (N_4254,In_882,In_461);
xor U4255 (N_4255,In_701,In_134);
or U4256 (N_4256,In_413,In_291);
or U4257 (N_4257,In_692,In_284);
and U4258 (N_4258,In_22,In_844);
and U4259 (N_4259,In_723,In_892);
and U4260 (N_4260,In_526,In_743);
nand U4261 (N_4261,In_248,In_485);
and U4262 (N_4262,In_912,In_651);
nor U4263 (N_4263,In_197,In_439);
and U4264 (N_4264,In_692,In_801);
and U4265 (N_4265,In_293,In_702);
nand U4266 (N_4266,In_690,In_873);
nand U4267 (N_4267,In_699,In_987);
nand U4268 (N_4268,In_418,In_838);
nor U4269 (N_4269,In_939,In_156);
nand U4270 (N_4270,In_859,In_374);
and U4271 (N_4271,In_582,In_315);
nand U4272 (N_4272,In_472,In_612);
nand U4273 (N_4273,In_734,In_774);
xor U4274 (N_4274,In_771,In_690);
nand U4275 (N_4275,In_242,In_933);
nor U4276 (N_4276,In_403,In_806);
or U4277 (N_4277,In_9,In_289);
nor U4278 (N_4278,In_617,In_135);
or U4279 (N_4279,In_583,In_887);
nand U4280 (N_4280,In_635,In_890);
nor U4281 (N_4281,In_141,In_610);
nand U4282 (N_4282,In_861,In_432);
and U4283 (N_4283,In_936,In_608);
nor U4284 (N_4284,In_90,In_771);
nor U4285 (N_4285,In_999,In_489);
or U4286 (N_4286,In_340,In_117);
and U4287 (N_4287,In_157,In_299);
and U4288 (N_4288,In_498,In_293);
and U4289 (N_4289,In_949,In_288);
nor U4290 (N_4290,In_530,In_310);
or U4291 (N_4291,In_542,In_887);
nand U4292 (N_4292,In_729,In_700);
or U4293 (N_4293,In_229,In_349);
and U4294 (N_4294,In_176,In_880);
nor U4295 (N_4295,In_852,In_998);
or U4296 (N_4296,In_574,In_467);
nor U4297 (N_4297,In_369,In_149);
nand U4298 (N_4298,In_345,In_933);
or U4299 (N_4299,In_220,In_32);
nand U4300 (N_4300,In_137,In_561);
or U4301 (N_4301,In_144,In_185);
nand U4302 (N_4302,In_818,In_857);
nor U4303 (N_4303,In_784,In_833);
nor U4304 (N_4304,In_422,In_640);
nor U4305 (N_4305,In_305,In_328);
or U4306 (N_4306,In_90,In_189);
and U4307 (N_4307,In_113,In_310);
and U4308 (N_4308,In_646,In_125);
and U4309 (N_4309,In_300,In_699);
nand U4310 (N_4310,In_322,In_874);
and U4311 (N_4311,In_578,In_427);
nor U4312 (N_4312,In_854,In_116);
nor U4313 (N_4313,In_650,In_3);
nor U4314 (N_4314,In_741,In_791);
nor U4315 (N_4315,In_761,In_421);
nand U4316 (N_4316,In_491,In_854);
or U4317 (N_4317,In_38,In_658);
or U4318 (N_4318,In_231,In_467);
nand U4319 (N_4319,In_426,In_517);
nor U4320 (N_4320,In_681,In_967);
and U4321 (N_4321,In_921,In_12);
nor U4322 (N_4322,In_647,In_175);
xor U4323 (N_4323,In_767,In_873);
nand U4324 (N_4324,In_594,In_964);
or U4325 (N_4325,In_956,In_232);
or U4326 (N_4326,In_936,In_712);
nand U4327 (N_4327,In_737,In_209);
and U4328 (N_4328,In_327,In_297);
xor U4329 (N_4329,In_610,In_519);
nor U4330 (N_4330,In_551,In_35);
and U4331 (N_4331,In_181,In_130);
xor U4332 (N_4332,In_667,In_76);
nand U4333 (N_4333,In_172,In_219);
nor U4334 (N_4334,In_703,In_909);
nor U4335 (N_4335,In_242,In_42);
or U4336 (N_4336,In_808,In_540);
nand U4337 (N_4337,In_544,In_368);
or U4338 (N_4338,In_174,In_585);
and U4339 (N_4339,In_847,In_11);
and U4340 (N_4340,In_876,In_390);
nand U4341 (N_4341,In_500,In_714);
or U4342 (N_4342,In_103,In_645);
or U4343 (N_4343,In_676,In_290);
and U4344 (N_4344,In_927,In_652);
or U4345 (N_4345,In_745,In_243);
nor U4346 (N_4346,In_6,In_944);
nand U4347 (N_4347,In_602,In_686);
nor U4348 (N_4348,In_686,In_499);
xnor U4349 (N_4349,In_575,In_869);
nor U4350 (N_4350,In_615,In_139);
or U4351 (N_4351,In_184,In_418);
nor U4352 (N_4352,In_302,In_525);
or U4353 (N_4353,In_548,In_805);
nor U4354 (N_4354,In_143,In_908);
nand U4355 (N_4355,In_839,In_303);
and U4356 (N_4356,In_726,In_639);
and U4357 (N_4357,In_586,In_710);
and U4358 (N_4358,In_281,In_12);
or U4359 (N_4359,In_512,In_268);
nor U4360 (N_4360,In_947,In_184);
or U4361 (N_4361,In_896,In_73);
nor U4362 (N_4362,In_371,In_952);
nand U4363 (N_4363,In_710,In_670);
nor U4364 (N_4364,In_825,In_975);
and U4365 (N_4365,In_677,In_437);
or U4366 (N_4366,In_41,In_171);
nor U4367 (N_4367,In_587,In_678);
nand U4368 (N_4368,In_577,In_334);
nor U4369 (N_4369,In_447,In_913);
xor U4370 (N_4370,In_533,In_375);
and U4371 (N_4371,In_838,In_59);
nor U4372 (N_4372,In_236,In_29);
nor U4373 (N_4373,In_61,In_242);
xor U4374 (N_4374,In_997,In_586);
and U4375 (N_4375,In_0,In_206);
or U4376 (N_4376,In_609,In_128);
nor U4377 (N_4377,In_784,In_80);
nand U4378 (N_4378,In_771,In_808);
nand U4379 (N_4379,In_267,In_515);
and U4380 (N_4380,In_728,In_534);
nor U4381 (N_4381,In_419,In_298);
xor U4382 (N_4382,In_706,In_749);
xor U4383 (N_4383,In_589,In_147);
nand U4384 (N_4384,In_279,In_695);
nor U4385 (N_4385,In_130,In_313);
nor U4386 (N_4386,In_823,In_355);
and U4387 (N_4387,In_665,In_683);
nand U4388 (N_4388,In_525,In_934);
and U4389 (N_4389,In_666,In_322);
xnor U4390 (N_4390,In_842,In_843);
and U4391 (N_4391,In_364,In_29);
or U4392 (N_4392,In_80,In_940);
nand U4393 (N_4393,In_529,In_561);
nand U4394 (N_4394,In_721,In_755);
xor U4395 (N_4395,In_853,In_399);
or U4396 (N_4396,In_501,In_851);
nor U4397 (N_4397,In_804,In_663);
xnor U4398 (N_4398,In_202,In_383);
and U4399 (N_4399,In_931,In_206);
and U4400 (N_4400,In_36,In_12);
nor U4401 (N_4401,In_141,In_712);
nor U4402 (N_4402,In_736,In_474);
and U4403 (N_4403,In_362,In_165);
nand U4404 (N_4404,In_210,In_667);
nor U4405 (N_4405,In_688,In_392);
or U4406 (N_4406,In_874,In_79);
xor U4407 (N_4407,In_895,In_539);
nor U4408 (N_4408,In_820,In_433);
or U4409 (N_4409,In_407,In_837);
and U4410 (N_4410,In_305,In_896);
nor U4411 (N_4411,In_532,In_542);
and U4412 (N_4412,In_31,In_711);
nor U4413 (N_4413,In_457,In_387);
xnor U4414 (N_4414,In_282,In_774);
xnor U4415 (N_4415,In_538,In_362);
nand U4416 (N_4416,In_519,In_971);
nor U4417 (N_4417,In_6,In_452);
and U4418 (N_4418,In_264,In_468);
and U4419 (N_4419,In_183,In_821);
nor U4420 (N_4420,In_968,In_238);
and U4421 (N_4421,In_955,In_841);
nand U4422 (N_4422,In_710,In_97);
or U4423 (N_4423,In_467,In_94);
or U4424 (N_4424,In_773,In_367);
or U4425 (N_4425,In_374,In_799);
nand U4426 (N_4426,In_134,In_309);
or U4427 (N_4427,In_702,In_122);
nand U4428 (N_4428,In_204,In_262);
nor U4429 (N_4429,In_322,In_43);
nand U4430 (N_4430,In_437,In_441);
nor U4431 (N_4431,In_358,In_435);
and U4432 (N_4432,In_254,In_655);
and U4433 (N_4433,In_126,In_880);
nand U4434 (N_4434,In_855,In_974);
or U4435 (N_4435,In_694,In_913);
or U4436 (N_4436,In_524,In_769);
and U4437 (N_4437,In_719,In_578);
and U4438 (N_4438,In_802,In_202);
and U4439 (N_4439,In_38,In_293);
or U4440 (N_4440,In_107,In_2);
or U4441 (N_4441,In_87,In_155);
nand U4442 (N_4442,In_267,In_326);
and U4443 (N_4443,In_267,In_793);
and U4444 (N_4444,In_765,In_188);
and U4445 (N_4445,In_580,In_199);
or U4446 (N_4446,In_532,In_253);
and U4447 (N_4447,In_336,In_112);
nor U4448 (N_4448,In_538,In_643);
nand U4449 (N_4449,In_149,In_773);
xnor U4450 (N_4450,In_729,In_979);
or U4451 (N_4451,In_96,In_496);
and U4452 (N_4452,In_177,In_622);
or U4453 (N_4453,In_500,In_860);
or U4454 (N_4454,In_67,In_455);
and U4455 (N_4455,In_848,In_550);
xor U4456 (N_4456,In_476,In_10);
or U4457 (N_4457,In_146,In_295);
nand U4458 (N_4458,In_20,In_883);
and U4459 (N_4459,In_688,In_638);
and U4460 (N_4460,In_37,In_288);
xnor U4461 (N_4461,In_956,In_765);
nor U4462 (N_4462,In_592,In_733);
nand U4463 (N_4463,In_777,In_348);
xor U4464 (N_4464,In_555,In_10);
nor U4465 (N_4465,In_683,In_262);
xnor U4466 (N_4466,In_295,In_143);
nor U4467 (N_4467,In_549,In_153);
or U4468 (N_4468,In_846,In_510);
nand U4469 (N_4469,In_991,In_238);
or U4470 (N_4470,In_522,In_135);
and U4471 (N_4471,In_746,In_865);
nand U4472 (N_4472,In_822,In_337);
nand U4473 (N_4473,In_955,In_397);
or U4474 (N_4474,In_191,In_323);
or U4475 (N_4475,In_717,In_786);
nor U4476 (N_4476,In_619,In_592);
nand U4477 (N_4477,In_227,In_494);
xnor U4478 (N_4478,In_77,In_613);
or U4479 (N_4479,In_615,In_313);
nand U4480 (N_4480,In_160,In_816);
or U4481 (N_4481,In_347,In_11);
nor U4482 (N_4482,In_198,In_637);
nand U4483 (N_4483,In_579,In_147);
nor U4484 (N_4484,In_311,In_317);
nand U4485 (N_4485,In_518,In_700);
xnor U4486 (N_4486,In_286,In_454);
nand U4487 (N_4487,In_746,In_898);
and U4488 (N_4488,In_687,In_982);
nor U4489 (N_4489,In_795,In_806);
and U4490 (N_4490,In_612,In_449);
or U4491 (N_4491,In_1,In_622);
nor U4492 (N_4492,In_880,In_518);
and U4493 (N_4493,In_993,In_923);
xor U4494 (N_4494,In_413,In_533);
xor U4495 (N_4495,In_367,In_964);
or U4496 (N_4496,In_876,In_434);
or U4497 (N_4497,In_852,In_173);
nor U4498 (N_4498,In_10,In_42);
and U4499 (N_4499,In_741,In_833);
or U4500 (N_4500,In_604,In_64);
nand U4501 (N_4501,In_226,In_769);
nor U4502 (N_4502,In_868,In_418);
nand U4503 (N_4503,In_79,In_481);
or U4504 (N_4504,In_600,In_6);
nor U4505 (N_4505,In_410,In_858);
nand U4506 (N_4506,In_246,In_81);
nor U4507 (N_4507,In_941,In_779);
nor U4508 (N_4508,In_544,In_319);
and U4509 (N_4509,In_768,In_241);
and U4510 (N_4510,In_353,In_431);
xnor U4511 (N_4511,In_986,In_138);
nand U4512 (N_4512,In_282,In_448);
nor U4513 (N_4513,In_936,In_994);
xnor U4514 (N_4514,In_576,In_424);
or U4515 (N_4515,In_253,In_924);
or U4516 (N_4516,In_293,In_670);
or U4517 (N_4517,In_599,In_148);
and U4518 (N_4518,In_618,In_38);
and U4519 (N_4519,In_458,In_897);
or U4520 (N_4520,In_780,In_581);
or U4521 (N_4521,In_785,In_380);
and U4522 (N_4522,In_647,In_4);
or U4523 (N_4523,In_435,In_255);
nand U4524 (N_4524,In_361,In_6);
and U4525 (N_4525,In_907,In_520);
and U4526 (N_4526,In_418,In_906);
nand U4527 (N_4527,In_658,In_844);
nor U4528 (N_4528,In_395,In_114);
or U4529 (N_4529,In_428,In_99);
and U4530 (N_4530,In_205,In_533);
nand U4531 (N_4531,In_116,In_392);
or U4532 (N_4532,In_22,In_730);
or U4533 (N_4533,In_689,In_395);
or U4534 (N_4534,In_988,In_761);
and U4535 (N_4535,In_649,In_825);
nor U4536 (N_4536,In_768,In_684);
and U4537 (N_4537,In_418,In_394);
nor U4538 (N_4538,In_330,In_693);
or U4539 (N_4539,In_655,In_56);
nand U4540 (N_4540,In_264,In_228);
or U4541 (N_4541,In_697,In_130);
nand U4542 (N_4542,In_74,In_466);
and U4543 (N_4543,In_661,In_801);
nor U4544 (N_4544,In_994,In_360);
or U4545 (N_4545,In_67,In_801);
and U4546 (N_4546,In_889,In_928);
and U4547 (N_4547,In_47,In_839);
and U4548 (N_4548,In_807,In_759);
or U4549 (N_4549,In_247,In_26);
nor U4550 (N_4550,In_625,In_533);
nand U4551 (N_4551,In_249,In_469);
nand U4552 (N_4552,In_580,In_676);
nor U4553 (N_4553,In_947,In_32);
nand U4554 (N_4554,In_134,In_214);
xnor U4555 (N_4555,In_179,In_893);
nand U4556 (N_4556,In_321,In_769);
and U4557 (N_4557,In_69,In_205);
and U4558 (N_4558,In_939,In_431);
nor U4559 (N_4559,In_121,In_448);
nor U4560 (N_4560,In_156,In_839);
or U4561 (N_4561,In_271,In_924);
or U4562 (N_4562,In_455,In_414);
and U4563 (N_4563,In_812,In_495);
nor U4564 (N_4564,In_273,In_695);
xor U4565 (N_4565,In_720,In_843);
and U4566 (N_4566,In_949,In_257);
and U4567 (N_4567,In_462,In_319);
or U4568 (N_4568,In_536,In_637);
nand U4569 (N_4569,In_867,In_59);
and U4570 (N_4570,In_66,In_203);
or U4571 (N_4571,In_717,In_558);
nand U4572 (N_4572,In_437,In_731);
nor U4573 (N_4573,In_408,In_732);
and U4574 (N_4574,In_758,In_561);
or U4575 (N_4575,In_6,In_920);
and U4576 (N_4576,In_277,In_808);
and U4577 (N_4577,In_472,In_346);
xor U4578 (N_4578,In_351,In_496);
nand U4579 (N_4579,In_230,In_279);
or U4580 (N_4580,In_760,In_743);
and U4581 (N_4581,In_901,In_819);
nor U4582 (N_4582,In_962,In_989);
xor U4583 (N_4583,In_756,In_110);
and U4584 (N_4584,In_447,In_280);
or U4585 (N_4585,In_795,In_309);
nor U4586 (N_4586,In_728,In_631);
nand U4587 (N_4587,In_97,In_497);
and U4588 (N_4588,In_764,In_722);
xnor U4589 (N_4589,In_483,In_762);
xnor U4590 (N_4590,In_33,In_76);
nor U4591 (N_4591,In_11,In_71);
nand U4592 (N_4592,In_799,In_616);
or U4593 (N_4593,In_213,In_569);
or U4594 (N_4594,In_368,In_426);
nand U4595 (N_4595,In_937,In_515);
or U4596 (N_4596,In_83,In_934);
or U4597 (N_4597,In_564,In_784);
or U4598 (N_4598,In_937,In_190);
or U4599 (N_4599,In_10,In_563);
and U4600 (N_4600,In_437,In_141);
nor U4601 (N_4601,In_641,In_2);
and U4602 (N_4602,In_678,In_320);
and U4603 (N_4603,In_356,In_77);
and U4604 (N_4604,In_578,In_345);
nor U4605 (N_4605,In_445,In_340);
nand U4606 (N_4606,In_262,In_400);
or U4607 (N_4607,In_97,In_367);
or U4608 (N_4608,In_296,In_798);
or U4609 (N_4609,In_406,In_314);
or U4610 (N_4610,In_462,In_942);
nand U4611 (N_4611,In_680,In_577);
and U4612 (N_4612,In_260,In_619);
and U4613 (N_4613,In_888,In_802);
or U4614 (N_4614,In_504,In_670);
nand U4615 (N_4615,In_676,In_891);
nor U4616 (N_4616,In_375,In_144);
or U4617 (N_4617,In_52,In_53);
nor U4618 (N_4618,In_880,In_562);
nand U4619 (N_4619,In_561,In_781);
nor U4620 (N_4620,In_999,In_153);
or U4621 (N_4621,In_353,In_355);
and U4622 (N_4622,In_849,In_448);
nor U4623 (N_4623,In_359,In_903);
nand U4624 (N_4624,In_558,In_358);
xor U4625 (N_4625,In_601,In_784);
nor U4626 (N_4626,In_113,In_685);
or U4627 (N_4627,In_627,In_861);
or U4628 (N_4628,In_964,In_696);
and U4629 (N_4629,In_165,In_142);
nand U4630 (N_4630,In_621,In_570);
or U4631 (N_4631,In_475,In_305);
and U4632 (N_4632,In_659,In_576);
or U4633 (N_4633,In_341,In_190);
nand U4634 (N_4634,In_686,In_549);
or U4635 (N_4635,In_409,In_281);
nand U4636 (N_4636,In_265,In_568);
or U4637 (N_4637,In_827,In_143);
or U4638 (N_4638,In_855,In_146);
and U4639 (N_4639,In_608,In_188);
nand U4640 (N_4640,In_442,In_741);
and U4641 (N_4641,In_711,In_600);
nor U4642 (N_4642,In_56,In_323);
and U4643 (N_4643,In_847,In_18);
or U4644 (N_4644,In_822,In_189);
and U4645 (N_4645,In_442,In_472);
nand U4646 (N_4646,In_70,In_83);
nand U4647 (N_4647,In_826,In_803);
or U4648 (N_4648,In_823,In_241);
xnor U4649 (N_4649,In_86,In_273);
or U4650 (N_4650,In_988,In_64);
nor U4651 (N_4651,In_429,In_103);
or U4652 (N_4652,In_803,In_718);
and U4653 (N_4653,In_275,In_326);
nand U4654 (N_4654,In_919,In_463);
nor U4655 (N_4655,In_691,In_919);
or U4656 (N_4656,In_196,In_176);
nor U4657 (N_4657,In_55,In_436);
or U4658 (N_4658,In_17,In_400);
nor U4659 (N_4659,In_885,In_431);
nand U4660 (N_4660,In_198,In_261);
or U4661 (N_4661,In_633,In_239);
nor U4662 (N_4662,In_339,In_71);
nor U4663 (N_4663,In_129,In_490);
and U4664 (N_4664,In_552,In_395);
nand U4665 (N_4665,In_713,In_791);
nand U4666 (N_4666,In_16,In_568);
xnor U4667 (N_4667,In_901,In_391);
or U4668 (N_4668,In_605,In_745);
or U4669 (N_4669,In_934,In_163);
and U4670 (N_4670,In_920,In_922);
nand U4671 (N_4671,In_94,In_424);
or U4672 (N_4672,In_154,In_62);
nand U4673 (N_4673,In_313,In_389);
nor U4674 (N_4674,In_420,In_923);
and U4675 (N_4675,In_504,In_12);
and U4676 (N_4676,In_263,In_193);
nor U4677 (N_4677,In_651,In_221);
and U4678 (N_4678,In_370,In_841);
and U4679 (N_4679,In_332,In_155);
or U4680 (N_4680,In_461,In_707);
nor U4681 (N_4681,In_578,In_185);
nand U4682 (N_4682,In_87,In_371);
and U4683 (N_4683,In_957,In_675);
nor U4684 (N_4684,In_142,In_888);
nand U4685 (N_4685,In_194,In_302);
nor U4686 (N_4686,In_124,In_436);
and U4687 (N_4687,In_734,In_539);
nand U4688 (N_4688,In_859,In_152);
nor U4689 (N_4689,In_148,In_549);
nor U4690 (N_4690,In_900,In_139);
and U4691 (N_4691,In_698,In_365);
nor U4692 (N_4692,In_680,In_134);
and U4693 (N_4693,In_319,In_998);
nor U4694 (N_4694,In_690,In_646);
or U4695 (N_4695,In_151,In_829);
nor U4696 (N_4696,In_926,In_645);
or U4697 (N_4697,In_792,In_740);
xor U4698 (N_4698,In_370,In_62);
nand U4699 (N_4699,In_84,In_926);
and U4700 (N_4700,In_935,In_0);
and U4701 (N_4701,In_642,In_983);
and U4702 (N_4702,In_577,In_710);
nand U4703 (N_4703,In_360,In_590);
nor U4704 (N_4704,In_633,In_267);
or U4705 (N_4705,In_961,In_784);
nor U4706 (N_4706,In_396,In_967);
nand U4707 (N_4707,In_451,In_423);
nor U4708 (N_4708,In_987,In_756);
xor U4709 (N_4709,In_690,In_416);
and U4710 (N_4710,In_84,In_238);
and U4711 (N_4711,In_982,In_303);
nand U4712 (N_4712,In_747,In_425);
nor U4713 (N_4713,In_861,In_804);
nand U4714 (N_4714,In_545,In_865);
or U4715 (N_4715,In_203,In_526);
xnor U4716 (N_4716,In_116,In_747);
nor U4717 (N_4717,In_255,In_632);
and U4718 (N_4718,In_494,In_500);
and U4719 (N_4719,In_314,In_792);
nor U4720 (N_4720,In_568,In_544);
nor U4721 (N_4721,In_518,In_9);
nand U4722 (N_4722,In_853,In_794);
nor U4723 (N_4723,In_602,In_364);
nand U4724 (N_4724,In_0,In_875);
or U4725 (N_4725,In_621,In_168);
nor U4726 (N_4726,In_766,In_416);
and U4727 (N_4727,In_519,In_585);
or U4728 (N_4728,In_598,In_603);
nand U4729 (N_4729,In_303,In_180);
or U4730 (N_4730,In_101,In_956);
nor U4731 (N_4731,In_44,In_814);
or U4732 (N_4732,In_364,In_743);
or U4733 (N_4733,In_623,In_231);
or U4734 (N_4734,In_649,In_842);
and U4735 (N_4735,In_69,In_346);
nor U4736 (N_4736,In_282,In_696);
nand U4737 (N_4737,In_948,In_839);
and U4738 (N_4738,In_470,In_200);
or U4739 (N_4739,In_991,In_661);
and U4740 (N_4740,In_161,In_567);
and U4741 (N_4741,In_189,In_975);
xor U4742 (N_4742,In_805,In_837);
and U4743 (N_4743,In_417,In_143);
and U4744 (N_4744,In_663,In_690);
and U4745 (N_4745,In_707,In_573);
and U4746 (N_4746,In_877,In_402);
or U4747 (N_4747,In_951,In_517);
nor U4748 (N_4748,In_561,In_317);
and U4749 (N_4749,In_128,In_960);
and U4750 (N_4750,In_341,In_792);
nor U4751 (N_4751,In_670,In_933);
nand U4752 (N_4752,In_343,In_787);
nor U4753 (N_4753,In_482,In_45);
nor U4754 (N_4754,In_697,In_675);
nor U4755 (N_4755,In_781,In_921);
nor U4756 (N_4756,In_312,In_383);
xnor U4757 (N_4757,In_88,In_516);
or U4758 (N_4758,In_606,In_496);
or U4759 (N_4759,In_221,In_771);
nor U4760 (N_4760,In_992,In_205);
nand U4761 (N_4761,In_694,In_517);
and U4762 (N_4762,In_275,In_152);
nor U4763 (N_4763,In_696,In_455);
and U4764 (N_4764,In_101,In_330);
nand U4765 (N_4765,In_433,In_622);
nand U4766 (N_4766,In_477,In_141);
nand U4767 (N_4767,In_468,In_947);
or U4768 (N_4768,In_317,In_510);
nor U4769 (N_4769,In_695,In_67);
nand U4770 (N_4770,In_853,In_781);
and U4771 (N_4771,In_610,In_369);
or U4772 (N_4772,In_648,In_635);
or U4773 (N_4773,In_930,In_965);
or U4774 (N_4774,In_793,In_615);
or U4775 (N_4775,In_911,In_447);
or U4776 (N_4776,In_649,In_457);
nor U4777 (N_4777,In_101,In_175);
nand U4778 (N_4778,In_905,In_438);
and U4779 (N_4779,In_335,In_699);
and U4780 (N_4780,In_527,In_317);
nand U4781 (N_4781,In_512,In_793);
nand U4782 (N_4782,In_229,In_288);
nor U4783 (N_4783,In_544,In_58);
and U4784 (N_4784,In_356,In_881);
or U4785 (N_4785,In_606,In_65);
xnor U4786 (N_4786,In_518,In_19);
or U4787 (N_4787,In_207,In_794);
or U4788 (N_4788,In_61,In_947);
and U4789 (N_4789,In_359,In_755);
and U4790 (N_4790,In_645,In_367);
nor U4791 (N_4791,In_866,In_581);
nor U4792 (N_4792,In_289,In_23);
nand U4793 (N_4793,In_660,In_395);
and U4794 (N_4794,In_47,In_596);
xor U4795 (N_4795,In_449,In_874);
or U4796 (N_4796,In_756,In_74);
or U4797 (N_4797,In_8,In_718);
and U4798 (N_4798,In_483,In_806);
nor U4799 (N_4799,In_362,In_625);
or U4800 (N_4800,In_791,In_441);
xnor U4801 (N_4801,In_719,In_85);
nand U4802 (N_4802,In_53,In_395);
and U4803 (N_4803,In_955,In_583);
and U4804 (N_4804,In_249,In_888);
nand U4805 (N_4805,In_940,In_851);
nand U4806 (N_4806,In_328,In_543);
nand U4807 (N_4807,In_466,In_937);
or U4808 (N_4808,In_85,In_720);
nand U4809 (N_4809,In_31,In_132);
and U4810 (N_4810,In_363,In_300);
and U4811 (N_4811,In_366,In_542);
nand U4812 (N_4812,In_207,In_665);
or U4813 (N_4813,In_442,In_188);
and U4814 (N_4814,In_112,In_385);
xor U4815 (N_4815,In_33,In_69);
or U4816 (N_4816,In_552,In_815);
xnor U4817 (N_4817,In_831,In_430);
nor U4818 (N_4818,In_9,In_450);
or U4819 (N_4819,In_758,In_99);
nor U4820 (N_4820,In_979,In_39);
and U4821 (N_4821,In_279,In_865);
or U4822 (N_4822,In_56,In_790);
or U4823 (N_4823,In_634,In_411);
or U4824 (N_4824,In_891,In_579);
nor U4825 (N_4825,In_785,In_647);
nand U4826 (N_4826,In_638,In_648);
nand U4827 (N_4827,In_81,In_172);
nand U4828 (N_4828,In_13,In_678);
and U4829 (N_4829,In_832,In_194);
nand U4830 (N_4830,In_346,In_758);
nor U4831 (N_4831,In_121,In_447);
and U4832 (N_4832,In_506,In_383);
or U4833 (N_4833,In_205,In_195);
xor U4834 (N_4834,In_805,In_402);
nand U4835 (N_4835,In_615,In_679);
or U4836 (N_4836,In_933,In_696);
nor U4837 (N_4837,In_597,In_868);
nand U4838 (N_4838,In_166,In_913);
nor U4839 (N_4839,In_72,In_935);
nand U4840 (N_4840,In_597,In_175);
and U4841 (N_4841,In_633,In_234);
or U4842 (N_4842,In_563,In_641);
and U4843 (N_4843,In_948,In_185);
nor U4844 (N_4844,In_317,In_829);
nand U4845 (N_4845,In_322,In_150);
and U4846 (N_4846,In_642,In_891);
and U4847 (N_4847,In_736,In_826);
nand U4848 (N_4848,In_258,In_976);
or U4849 (N_4849,In_685,In_457);
and U4850 (N_4850,In_184,In_771);
xnor U4851 (N_4851,In_742,In_9);
nor U4852 (N_4852,In_573,In_782);
and U4853 (N_4853,In_246,In_83);
nor U4854 (N_4854,In_12,In_60);
nand U4855 (N_4855,In_278,In_95);
nand U4856 (N_4856,In_783,In_516);
or U4857 (N_4857,In_532,In_741);
nor U4858 (N_4858,In_942,In_119);
nand U4859 (N_4859,In_442,In_907);
nand U4860 (N_4860,In_809,In_191);
and U4861 (N_4861,In_156,In_126);
and U4862 (N_4862,In_970,In_234);
xor U4863 (N_4863,In_402,In_917);
nor U4864 (N_4864,In_638,In_171);
xnor U4865 (N_4865,In_183,In_981);
or U4866 (N_4866,In_946,In_462);
nor U4867 (N_4867,In_402,In_445);
nor U4868 (N_4868,In_556,In_96);
and U4869 (N_4869,In_46,In_703);
xnor U4870 (N_4870,In_770,In_156);
and U4871 (N_4871,In_950,In_987);
xnor U4872 (N_4872,In_114,In_52);
or U4873 (N_4873,In_10,In_199);
xnor U4874 (N_4874,In_867,In_67);
or U4875 (N_4875,In_666,In_914);
and U4876 (N_4876,In_796,In_641);
xnor U4877 (N_4877,In_874,In_93);
or U4878 (N_4878,In_880,In_937);
or U4879 (N_4879,In_66,In_469);
nor U4880 (N_4880,In_943,In_345);
or U4881 (N_4881,In_484,In_781);
or U4882 (N_4882,In_83,In_205);
xnor U4883 (N_4883,In_261,In_857);
nand U4884 (N_4884,In_413,In_985);
and U4885 (N_4885,In_824,In_727);
xnor U4886 (N_4886,In_181,In_905);
nand U4887 (N_4887,In_207,In_789);
or U4888 (N_4888,In_96,In_684);
nand U4889 (N_4889,In_119,In_812);
xor U4890 (N_4890,In_491,In_140);
nor U4891 (N_4891,In_353,In_917);
or U4892 (N_4892,In_960,In_145);
or U4893 (N_4893,In_168,In_591);
or U4894 (N_4894,In_423,In_182);
nor U4895 (N_4895,In_25,In_702);
and U4896 (N_4896,In_806,In_958);
xnor U4897 (N_4897,In_750,In_389);
or U4898 (N_4898,In_196,In_870);
nor U4899 (N_4899,In_558,In_382);
or U4900 (N_4900,In_301,In_829);
nor U4901 (N_4901,In_162,In_482);
or U4902 (N_4902,In_302,In_622);
and U4903 (N_4903,In_843,In_157);
and U4904 (N_4904,In_121,In_535);
or U4905 (N_4905,In_786,In_929);
and U4906 (N_4906,In_699,In_190);
nor U4907 (N_4907,In_214,In_368);
and U4908 (N_4908,In_973,In_987);
nand U4909 (N_4909,In_637,In_424);
and U4910 (N_4910,In_873,In_52);
and U4911 (N_4911,In_928,In_483);
nor U4912 (N_4912,In_68,In_689);
nor U4913 (N_4913,In_298,In_388);
nor U4914 (N_4914,In_309,In_268);
nor U4915 (N_4915,In_110,In_829);
or U4916 (N_4916,In_167,In_854);
or U4917 (N_4917,In_733,In_337);
and U4918 (N_4918,In_768,In_535);
nor U4919 (N_4919,In_971,In_774);
and U4920 (N_4920,In_861,In_594);
and U4921 (N_4921,In_481,In_18);
nand U4922 (N_4922,In_18,In_826);
nor U4923 (N_4923,In_517,In_823);
nand U4924 (N_4924,In_455,In_693);
nor U4925 (N_4925,In_482,In_432);
nor U4926 (N_4926,In_324,In_674);
nor U4927 (N_4927,In_140,In_392);
nor U4928 (N_4928,In_321,In_470);
or U4929 (N_4929,In_234,In_741);
and U4930 (N_4930,In_517,In_412);
or U4931 (N_4931,In_337,In_254);
nand U4932 (N_4932,In_39,In_224);
nand U4933 (N_4933,In_6,In_345);
or U4934 (N_4934,In_163,In_939);
nor U4935 (N_4935,In_520,In_316);
or U4936 (N_4936,In_666,In_380);
or U4937 (N_4937,In_991,In_158);
nand U4938 (N_4938,In_687,In_177);
or U4939 (N_4939,In_357,In_374);
or U4940 (N_4940,In_873,In_897);
and U4941 (N_4941,In_91,In_388);
or U4942 (N_4942,In_59,In_567);
or U4943 (N_4943,In_628,In_286);
or U4944 (N_4944,In_803,In_892);
and U4945 (N_4945,In_957,In_489);
nand U4946 (N_4946,In_224,In_97);
or U4947 (N_4947,In_815,In_684);
xnor U4948 (N_4948,In_908,In_124);
or U4949 (N_4949,In_39,In_238);
and U4950 (N_4950,In_709,In_836);
and U4951 (N_4951,In_647,In_169);
nor U4952 (N_4952,In_384,In_576);
or U4953 (N_4953,In_898,In_294);
or U4954 (N_4954,In_357,In_636);
and U4955 (N_4955,In_346,In_49);
or U4956 (N_4956,In_232,In_453);
xor U4957 (N_4957,In_293,In_667);
xor U4958 (N_4958,In_984,In_920);
or U4959 (N_4959,In_677,In_92);
nand U4960 (N_4960,In_152,In_320);
or U4961 (N_4961,In_276,In_401);
nor U4962 (N_4962,In_931,In_492);
and U4963 (N_4963,In_655,In_760);
xor U4964 (N_4964,In_433,In_579);
nand U4965 (N_4965,In_302,In_42);
or U4966 (N_4966,In_627,In_33);
and U4967 (N_4967,In_460,In_80);
or U4968 (N_4968,In_143,In_127);
or U4969 (N_4969,In_179,In_978);
or U4970 (N_4970,In_507,In_393);
or U4971 (N_4971,In_666,In_501);
nand U4972 (N_4972,In_401,In_81);
and U4973 (N_4973,In_466,In_197);
nand U4974 (N_4974,In_4,In_570);
or U4975 (N_4975,In_351,In_242);
or U4976 (N_4976,In_126,In_175);
nor U4977 (N_4977,In_659,In_430);
nor U4978 (N_4978,In_138,In_128);
and U4979 (N_4979,In_370,In_41);
nor U4980 (N_4980,In_384,In_891);
nand U4981 (N_4981,In_985,In_62);
and U4982 (N_4982,In_633,In_42);
and U4983 (N_4983,In_736,In_340);
and U4984 (N_4984,In_531,In_789);
nand U4985 (N_4985,In_186,In_944);
and U4986 (N_4986,In_210,In_757);
and U4987 (N_4987,In_591,In_794);
or U4988 (N_4988,In_0,In_375);
and U4989 (N_4989,In_795,In_71);
nor U4990 (N_4990,In_233,In_385);
nand U4991 (N_4991,In_946,In_834);
or U4992 (N_4992,In_316,In_449);
nor U4993 (N_4993,In_563,In_773);
or U4994 (N_4994,In_924,In_901);
and U4995 (N_4995,In_427,In_959);
and U4996 (N_4996,In_719,In_811);
nor U4997 (N_4997,In_390,In_989);
nor U4998 (N_4998,In_21,In_141);
nand U4999 (N_4999,In_746,In_596);
or U5000 (N_5000,N_3102,N_872);
or U5001 (N_5001,N_108,N_3694);
or U5002 (N_5002,N_3186,N_1629);
nor U5003 (N_5003,N_814,N_167);
nand U5004 (N_5004,N_2874,N_1203);
and U5005 (N_5005,N_4050,N_4261);
nand U5006 (N_5006,N_3270,N_1292);
and U5007 (N_5007,N_3724,N_3422);
or U5008 (N_5008,N_3906,N_4613);
and U5009 (N_5009,N_917,N_1973);
nand U5010 (N_5010,N_2711,N_2331);
nor U5011 (N_5011,N_1961,N_2721);
nand U5012 (N_5012,N_2825,N_4719);
nand U5013 (N_5013,N_1969,N_2282);
xnor U5014 (N_5014,N_3412,N_3407);
and U5015 (N_5015,N_4020,N_2794);
nor U5016 (N_5016,N_3318,N_2700);
xor U5017 (N_5017,N_2865,N_112);
nand U5018 (N_5018,N_4198,N_3534);
and U5019 (N_5019,N_3925,N_232);
nor U5020 (N_5020,N_3175,N_26);
nor U5021 (N_5021,N_2011,N_1431);
nand U5022 (N_5022,N_3493,N_45);
or U5023 (N_5023,N_3605,N_4589);
nor U5024 (N_5024,N_2276,N_4926);
and U5025 (N_5025,N_1803,N_3178);
and U5026 (N_5026,N_1135,N_3745);
nand U5027 (N_5027,N_2266,N_3599);
nand U5028 (N_5028,N_1596,N_3016);
and U5029 (N_5029,N_113,N_3518);
nor U5030 (N_5030,N_3709,N_3707);
and U5031 (N_5031,N_3688,N_4462);
nand U5032 (N_5032,N_1650,N_2586);
nor U5033 (N_5033,N_3037,N_1792);
nor U5034 (N_5034,N_3877,N_2968);
or U5035 (N_5035,N_4790,N_2800);
nand U5036 (N_5036,N_2490,N_1917);
nand U5037 (N_5037,N_12,N_1702);
and U5038 (N_5038,N_3630,N_576);
xnor U5039 (N_5039,N_1923,N_1414);
nor U5040 (N_5040,N_3683,N_1831);
xor U5041 (N_5041,N_1995,N_1010);
or U5042 (N_5042,N_4944,N_554);
or U5043 (N_5043,N_2294,N_4980);
nor U5044 (N_5044,N_4186,N_157);
or U5045 (N_5045,N_2051,N_4597);
or U5046 (N_5046,N_95,N_3060);
nand U5047 (N_5047,N_3509,N_2879);
nand U5048 (N_5048,N_851,N_4220);
nand U5049 (N_5049,N_2295,N_4939);
xor U5050 (N_5050,N_1574,N_1371);
nand U5051 (N_5051,N_3780,N_898);
and U5052 (N_5052,N_3800,N_2569);
or U5053 (N_5053,N_886,N_1685);
or U5054 (N_5054,N_2081,N_4494);
nand U5055 (N_5055,N_330,N_227);
nand U5056 (N_5056,N_4952,N_3212);
or U5057 (N_5057,N_4160,N_3655);
or U5058 (N_5058,N_130,N_4617);
or U5059 (N_5059,N_3863,N_4463);
nor U5060 (N_5060,N_3606,N_468);
nor U5061 (N_5061,N_573,N_2430);
nor U5062 (N_5062,N_1339,N_2324);
xor U5063 (N_5063,N_1535,N_1784);
nand U5064 (N_5064,N_4507,N_1);
or U5065 (N_5065,N_2252,N_4084);
nor U5066 (N_5066,N_3841,N_4741);
and U5067 (N_5067,N_129,N_2418);
and U5068 (N_5068,N_4841,N_4769);
nor U5069 (N_5069,N_4139,N_1937);
xor U5070 (N_5070,N_3446,N_3512);
nor U5071 (N_5071,N_1074,N_1821);
nand U5072 (N_5072,N_1948,N_813);
and U5073 (N_5073,N_632,N_3849);
and U5074 (N_5074,N_3919,N_451);
xor U5075 (N_5075,N_1694,N_4179);
nand U5076 (N_5076,N_1418,N_2053);
nor U5077 (N_5077,N_3762,N_3380);
or U5078 (N_5078,N_4510,N_2082);
and U5079 (N_5079,N_4716,N_4620);
nor U5080 (N_5080,N_581,N_4073);
or U5081 (N_5081,N_3007,N_392);
nor U5082 (N_5082,N_2519,N_217);
or U5083 (N_5083,N_4820,N_3144);
nor U5084 (N_5084,N_2254,N_1172);
nand U5085 (N_5085,N_1982,N_2801);
or U5086 (N_5086,N_561,N_958);
nor U5087 (N_5087,N_1857,N_2579);
xnor U5088 (N_5088,N_3337,N_490);
and U5089 (N_5089,N_2540,N_1660);
nor U5090 (N_5090,N_571,N_4700);
xor U5091 (N_5091,N_2936,N_3379);
or U5092 (N_5092,N_4253,N_744);
and U5093 (N_5093,N_4149,N_2894);
and U5094 (N_5094,N_1706,N_2609);
xor U5095 (N_5095,N_2042,N_1711);
or U5096 (N_5096,N_2610,N_32);
nand U5097 (N_5097,N_976,N_3131);
or U5098 (N_5098,N_3190,N_2957);
xor U5099 (N_5099,N_2173,N_3262);
nand U5100 (N_5100,N_2376,N_4235);
nand U5101 (N_5101,N_1163,N_4001);
and U5102 (N_5102,N_890,N_1868);
and U5103 (N_5103,N_3842,N_1176);
or U5104 (N_5104,N_3558,N_2256);
nor U5105 (N_5105,N_1173,N_4935);
or U5106 (N_5106,N_4779,N_193);
and U5107 (N_5107,N_2654,N_2262);
nand U5108 (N_5108,N_2336,N_3503);
or U5109 (N_5109,N_3818,N_4246);
nor U5110 (N_5110,N_1737,N_1394);
nor U5111 (N_5111,N_656,N_4512);
and U5112 (N_5112,N_3888,N_4975);
or U5113 (N_5113,N_2204,N_2299);
nand U5114 (N_5114,N_962,N_4257);
nor U5115 (N_5115,N_1206,N_4749);
xnor U5116 (N_5116,N_196,N_497);
nor U5117 (N_5117,N_1497,N_1318);
nand U5118 (N_5118,N_2682,N_927);
and U5119 (N_5119,N_307,N_1362);
nand U5120 (N_5120,N_2064,N_1168);
nor U5121 (N_5121,N_1966,N_655);
nor U5122 (N_5122,N_251,N_3438);
and U5123 (N_5123,N_4730,N_3961);
nor U5124 (N_5124,N_3740,N_3561);
nor U5125 (N_5125,N_2691,N_4519);
nor U5126 (N_5126,N_3361,N_206);
nor U5127 (N_5127,N_2175,N_187);
or U5128 (N_5128,N_3875,N_1395);
or U5129 (N_5129,N_4872,N_3426);
or U5130 (N_5130,N_1117,N_2161);
nor U5131 (N_5131,N_1048,N_4013);
nor U5132 (N_5132,N_4919,N_4207);
nand U5133 (N_5133,N_30,N_987);
nand U5134 (N_5134,N_1107,N_198);
nor U5135 (N_5135,N_3880,N_4039);
xor U5136 (N_5136,N_714,N_4969);
and U5137 (N_5137,N_250,N_849);
nor U5138 (N_5138,N_1090,N_3417);
nor U5139 (N_5139,N_1126,N_1007);
or U5140 (N_5140,N_2284,N_671);
and U5141 (N_5141,N_87,N_2697);
nor U5142 (N_5142,N_1445,N_3205);
nand U5143 (N_5143,N_1401,N_4717);
or U5144 (N_5144,N_2828,N_267);
or U5145 (N_5145,N_549,N_3492);
nor U5146 (N_5146,N_4292,N_1481);
nor U5147 (N_5147,N_841,N_382);
nor U5148 (N_5148,N_4671,N_104);
nor U5149 (N_5149,N_919,N_4782);
xor U5150 (N_5150,N_163,N_4166);
and U5151 (N_5151,N_4351,N_244);
or U5152 (N_5152,N_3506,N_2308);
and U5153 (N_5153,N_147,N_425);
nand U5154 (N_5154,N_1558,N_826);
and U5155 (N_5155,N_1960,N_3309);
nor U5156 (N_5156,N_1125,N_4865);
nor U5157 (N_5157,N_2673,N_3794);
nand U5158 (N_5158,N_2991,N_2988);
and U5159 (N_5159,N_4454,N_4214);
nor U5160 (N_5160,N_1536,N_4009);
nor U5161 (N_5161,N_4051,N_4727);
nor U5162 (N_5162,N_2456,N_1734);
nand U5163 (N_5163,N_2333,N_915);
and U5164 (N_5164,N_4352,N_2970);
and U5165 (N_5165,N_2612,N_242);
nor U5166 (N_5166,N_3408,N_1249);
xnor U5167 (N_5167,N_46,N_679);
nor U5168 (N_5168,N_766,N_3069);
or U5169 (N_5169,N_4541,N_4855);
or U5170 (N_5170,N_1120,N_786);
nand U5171 (N_5171,N_2311,N_4338);
or U5172 (N_5172,N_2489,N_1407);
nor U5173 (N_5173,N_346,N_2655);
xnor U5174 (N_5174,N_1907,N_4864);
nand U5175 (N_5175,N_3308,N_558);
nor U5176 (N_5176,N_1199,N_2242);
and U5177 (N_5177,N_2237,N_4079);
and U5178 (N_5178,N_295,N_4918);
nor U5179 (N_5179,N_4602,N_2117);
or U5180 (N_5180,N_162,N_2850);
nor U5181 (N_5181,N_1712,N_4100);
or U5182 (N_5182,N_752,N_4335);
nor U5183 (N_5183,N_527,N_3944);
or U5184 (N_5184,N_4890,N_1511);
nand U5185 (N_5185,N_2103,N_2361);
nand U5186 (N_5186,N_4773,N_2961);
or U5187 (N_5187,N_1128,N_1326);
or U5188 (N_5188,N_2594,N_2791);
nand U5189 (N_5189,N_4995,N_3654);
xnor U5190 (N_5190,N_4049,N_722);
or U5191 (N_5191,N_2537,N_4469);
nor U5192 (N_5192,N_1940,N_2492);
or U5193 (N_5193,N_4204,N_3592);
or U5194 (N_5194,N_2509,N_694);
and U5195 (N_5195,N_4448,N_609);
xnor U5196 (N_5196,N_2057,N_4345);
or U5197 (N_5197,N_3844,N_2575);
xnor U5198 (N_5198,N_386,N_1698);
nor U5199 (N_5199,N_3404,N_973);
xnor U5200 (N_5200,N_3381,N_3428);
nand U5201 (N_5201,N_2293,N_690);
nor U5202 (N_5202,N_1827,N_4892);
xnor U5203 (N_5203,N_1597,N_4284);
or U5204 (N_5204,N_1462,N_4453);
xnor U5205 (N_5205,N_4319,N_3276);
nand U5206 (N_5206,N_218,N_1210);
and U5207 (N_5207,N_4112,N_4907);
nand U5208 (N_5208,N_4687,N_3964);
xor U5209 (N_5209,N_3536,N_2368);
nor U5210 (N_5210,N_4118,N_1240);
xnor U5211 (N_5211,N_2249,N_831);
or U5212 (N_5212,N_4847,N_4533);
xnor U5213 (N_5213,N_1467,N_4333);
xnor U5214 (N_5214,N_2595,N_1305);
xor U5215 (N_5215,N_824,N_2317);
or U5216 (N_5216,N_3808,N_2208);
or U5217 (N_5217,N_3706,N_80);
nand U5218 (N_5218,N_4997,N_3315);
nand U5219 (N_5219,N_2468,N_1520);
or U5220 (N_5220,N_4406,N_3195);
nor U5221 (N_5221,N_3923,N_1179);
xor U5222 (N_5222,N_2760,N_621);
and U5223 (N_5223,N_525,N_3570);
and U5224 (N_5224,N_799,N_3858);
nor U5225 (N_5225,N_3832,N_3301);
nand U5226 (N_5226,N_2954,N_4609);
nand U5227 (N_5227,N_509,N_2104);
or U5228 (N_5228,N_1278,N_3343);
nor U5229 (N_5229,N_4663,N_1646);
or U5230 (N_5230,N_3608,N_4422);
nand U5231 (N_5231,N_1002,N_3513);
nor U5232 (N_5232,N_668,N_4960);
xnor U5233 (N_5233,N_4684,N_1833);
nand U5234 (N_5234,N_4571,N_178);
nor U5235 (N_5235,N_4954,N_1483);
xor U5236 (N_5236,N_1012,N_1582);
and U5237 (N_5237,N_42,N_3817);
and U5238 (N_5238,N_4317,N_4313);
nor U5239 (N_5239,N_3391,N_1461);
and U5240 (N_5240,N_3348,N_4818);
nand U5241 (N_5241,N_291,N_2137);
xnor U5242 (N_5242,N_4817,N_109);
or U5243 (N_5243,N_2320,N_3731);
and U5244 (N_5244,N_1083,N_420);
or U5245 (N_5245,N_3192,N_3960);
nand U5246 (N_5246,N_1096,N_3109);
and U5247 (N_5247,N_2883,N_731);
or U5248 (N_5248,N_321,N_2561);
or U5249 (N_5249,N_4807,N_4056);
nand U5250 (N_5250,N_599,N_3411);
or U5251 (N_5251,N_3983,N_3331);
nand U5252 (N_5252,N_3631,N_3073);
nor U5253 (N_5253,N_3202,N_3458);
nor U5254 (N_5254,N_1681,N_4029);
nand U5255 (N_5255,N_4635,N_2375);
nor U5256 (N_5256,N_2600,N_1277);
or U5257 (N_5257,N_3734,N_177);
and U5258 (N_5258,N_4413,N_3702);
and U5259 (N_5259,N_2822,N_4178);
and U5260 (N_5260,N_2693,N_1436);
and U5261 (N_5261,N_243,N_1018);
or U5262 (N_5262,N_2934,N_3632);
xnor U5263 (N_5263,N_1599,N_829);
nand U5264 (N_5264,N_3003,N_723);
xor U5265 (N_5265,N_1755,N_3161);
nor U5266 (N_5266,N_1251,N_2386);
nand U5267 (N_5267,N_417,N_1617);
or U5268 (N_5268,N_3194,N_2426);
and U5269 (N_5269,N_1241,N_4083);
and U5270 (N_5270,N_710,N_3779);
nor U5271 (N_5271,N_811,N_3671);
or U5272 (N_5272,N_1109,N_2189);
or U5273 (N_5273,N_1196,N_1219);
nor U5274 (N_5274,N_3074,N_4738);
or U5275 (N_5275,N_2166,N_334);
or U5276 (N_5276,N_4608,N_904);
and U5277 (N_5277,N_2010,N_3292);
nor U5278 (N_5278,N_3157,N_2974);
or U5279 (N_5279,N_4685,N_4189);
nand U5280 (N_5280,N_3299,N_3722);
xor U5281 (N_5281,N_4374,N_2488);
nor U5282 (N_5282,N_3966,N_4366);
xnor U5283 (N_5283,N_4213,N_1990);
or U5284 (N_5284,N_102,N_2515);
nor U5285 (N_5285,N_3120,N_2170);
or U5286 (N_5286,N_4707,N_3350);
nand U5287 (N_5287,N_3826,N_760);
or U5288 (N_5288,N_1841,N_3902);
nand U5289 (N_5289,N_28,N_340);
or U5290 (N_5290,N_471,N_279);
or U5291 (N_5291,N_2888,N_2842);
nand U5292 (N_5292,N_4300,N_4670);
nor U5293 (N_5293,N_1986,N_2583);
nand U5294 (N_5294,N_3303,N_2660);
nor U5295 (N_5295,N_2843,N_2578);
nor U5296 (N_5296,N_900,N_770);
and U5297 (N_5297,N_3134,N_2159);
nand U5298 (N_5298,N_4269,N_3837);
or U5299 (N_5299,N_3839,N_812);
nor U5300 (N_5300,N_4812,N_2710);
nand U5301 (N_5301,N_3203,N_560);
and U5302 (N_5302,N_593,N_4611);
nand U5303 (N_5303,N_60,N_1032);
xor U5304 (N_5304,N_3383,N_2824);
nand U5305 (N_5305,N_2587,N_2931);
and U5306 (N_5306,N_3965,N_352);
nor U5307 (N_5307,N_1656,N_362);
nor U5308 (N_5308,N_3742,N_2555);
nand U5309 (N_5309,N_3240,N_90);
nor U5310 (N_5310,N_4874,N_2724);
nand U5311 (N_5311,N_4423,N_3065);
nor U5312 (N_5312,N_4479,N_2482);
nor U5313 (N_5313,N_3133,N_2350);
nor U5314 (N_5314,N_2347,N_4880);
nor U5315 (N_5315,N_1570,N_1603);
nand U5316 (N_5316,N_4516,N_3444);
nand U5317 (N_5317,N_1636,N_2154);
nand U5318 (N_5318,N_1188,N_3653);
or U5319 (N_5319,N_3810,N_2054);
nand U5320 (N_5320,N_4535,N_1863);
or U5321 (N_5321,N_1337,N_1189);
nor U5322 (N_5322,N_3633,N_2596);
or U5323 (N_5323,N_4254,N_2613);
nand U5324 (N_5324,N_455,N_780);
nand U5325 (N_5325,N_536,N_1814);
xor U5326 (N_5326,N_3886,N_771);
nand U5327 (N_5327,N_4552,N_4408);
or U5328 (N_5328,N_3012,N_3545);
xnor U5329 (N_5329,N_2434,N_4403);
nand U5330 (N_5330,N_2813,N_2698);
nand U5331 (N_5331,N_1268,N_467);
or U5332 (N_5332,N_488,N_1524);
nor U5333 (N_5333,N_2562,N_4389);
or U5334 (N_5334,N_2549,N_951);
nand U5335 (N_5335,N_4973,N_4848);
nand U5336 (N_5336,N_4175,N_3788);
or U5337 (N_5337,N_4304,N_2754);
nor U5338 (N_5338,N_2184,N_2378);
nor U5339 (N_5339,N_3862,N_3256);
and U5340 (N_5340,N_720,N_3048);
nor U5341 (N_5341,N_1137,N_1084);
and U5342 (N_5342,N_843,N_4053);
nand U5343 (N_5343,N_2097,N_972);
or U5344 (N_5344,N_4043,N_70);
nand U5345 (N_5345,N_3751,N_1218);
and U5346 (N_5346,N_4770,N_3972);
nor U5347 (N_5347,N_27,N_1106);
or U5348 (N_5348,N_4409,N_4583);
or U5349 (N_5349,N_1983,N_4068);
nand U5350 (N_5350,N_1770,N_1024);
and U5351 (N_5351,N_1740,N_1951);
xnor U5352 (N_5352,N_2845,N_4721);
nor U5353 (N_5353,N_3713,N_3845);
or U5354 (N_5354,N_4776,N_689);
and U5355 (N_5355,N_2436,N_2025);
and U5356 (N_5356,N_4612,N_4775);
nand U5357 (N_5357,N_2169,N_3791);
nand U5358 (N_5358,N_4638,N_4110);
or U5359 (N_5359,N_3141,N_4481);
and U5360 (N_5360,N_4237,N_4850);
nand U5361 (N_5361,N_4802,N_4391);
nand U5362 (N_5362,N_1458,N_199);
nand U5363 (N_5363,N_442,N_2326);
nor U5364 (N_5364,N_2499,N_961);
or U5365 (N_5365,N_134,N_75);
nand U5366 (N_5366,N_4265,N_2152);
or U5367 (N_5367,N_3040,N_1115);
nand U5368 (N_5368,N_1092,N_3311);
or U5369 (N_5369,N_1543,N_4165);
or U5370 (N_5370,N_4250,N_3621);
nor U5371 (N_5371,N_4236,N_1040);
or U5372 (N_5372,N_1170,N_3782);
nand U5373 (N_5373,N_4968,N_4966);
and U5374 (N_5374,N_1864,N_4930);
and U5375 (N_5375,N_1512,N_3449);
and U5376 (N_5376,N_1064,N_1667);
or U5377 (N_5377,N_3191,N_4393);
or U5378 (N_5378,N_3868,N_2639);
nand U5379 (N_5379,N_1585,N_138);
or U5380 (N_5380,N_4295,N_1213);
or U5381 (N_5381,N_132,N_4579);
nand U5382 (N_5382,N_4696,N_4285);
and U5383 (N_5383,N_3319,N_550);
or U5384 (N_5384,N_2965,N_3386);
or U5385 (N_5385,N_2038,N_15);
nand U5386 (N_5386,N_4526,N_4244);
nor U5387 (N_5387,N_4574,N_981);
or U5388 (N_5388,N_1771,N_2742);
and U5389 (N_5389,N_889,N_4724);
nor U5390 (N_5390,N_207,N_706);
nand U5391 (N_5391,N_4645,N_4396);
or U5392 (N_5392,N_3281,N_2558);
and U5393 (N_5393,N_1510,N_2390);
nor U5394 (N_5394,N_1503,N_4065);
nor U5395 (N_5395,N_2958,N_4953);
nand U5396 (N_5396,N_1579,N_1099);
and U5397 (N_5397,N_4761,N_3406);
or U5398 (N_5398,N_2358,N_1642);
and U5399 (N_5399,N_670,N_4844);
and U5400 (N_5400,N_29,N_4998);
and U5401 (N_5401,N_4281,N_630);
nor U5402 (N_5402,N_1915,N_1386);
nor U5403 (N_5403,N_197,N_640);
nand U5404 (N_5404,N_472,N_538);
and U5405 (N_5405,N_411,N_1297);
and U5406 (N_5406,N_4920,N_4542);
or U5407 (N_5407,N_2315,N_1521);
nor U5408 (N_5408,N_3847,N_3106);
and U5409 (N_5409,N_4825,N_4537);
nand U5410 (N_5410,N_2534,N_3882);
and U5411 (N_5411,N_4098,N_2628);
nor U5412 (N_5412,N_3593,N_4852);
or U5413 (N_5413,N_1914,N_309);
or U5414 (N_5414,N_4756,N_2484);
nand U5415 (N_5415,N_1364,N_4725);
nand U5416 (N_5416,N_778,N_1062);
nor U5417 (N_5417,N_2199,N_2381);
nor U5418 (N_5418,N_3483,N_1586);
or U5419 (N_5419,N_2155,N_4411);
or U5420 (N_5420,N_2120,N_3660);
nor U5421 (N_5421,N_1367,N_4965);
and U5422 (N_5422,N_4266,N_4087);
xnor U5423 (N_5423,N_128,N_820);
nand U5424 (N_5424,N_4651,N_3129);
and U5425 (N_5425,N_1112,N_3812);
xnor U5426 (N_5426,N_1728,N_1081);
or U5427 (N_5427,N_4233,N_4977);
nor U5428 (N_5428,N_1250,N_551);
nand U5429 (N_5429,N_2000,N_1225);
and U5430 (N_5430,N_4778,N_3748);
and U5431 (N_5431,N_4373,N_570);
nand U5432 (N_5432,N_2116,N_960);
or U5433 (N_5433,N_686,N_2135);
nor U5434 (N_5434,N_1693,N_1807);
nand U5435 (N_5435,N_3760,N_436);
nor U5436 (N_5436,N_1086,N_4340);
or U5437 (N_5437,N_618,N_2545);
xnor U5438 (N_5438,N_2423,N_450);
nor U5439 (N_5439,N_1194,N_3789);
xor U5440 (N_5440,N_348,N_2061);
and U5441 (N_5441,N_1067,N_1042);
xor U5442 (N_5442,N_3261,N_4227);
and U5443 (N_5443,N_1848,N_1376);
nand U5444 (N_5444,N_4708,N_4249);
or U5445 (N_5445,N_1321,N_413);
nor U5446 (N_5446,N_3777,N_3767);
or U5447 (N_5447,N_769,N_1180);
xor U5448 (N_5448,N_4468,N_3017);
or U5449 (N_5449,N_1254,N_1313);
nand U5450 (N_5450,N_3326,N_3830);
or U5451 (N_5451,N_371,N_4430);
xor U5452 (N_5452,N_3879,N_4681);
xor U5453 (N_5453,N_785,N_574);
or U5454 (N_5454,N_4272,N_3604);
and U5455 (N_5455,N_3486,N_3568);
and U5456 (N_5456,N_72,N_908);
nor U5457 (N_5457,N_2220,N_3434);
or U5458 (N_5458,N_1439,N_3254);
xnor U5459 (N_5459,N_4694,N_2916);
or U5460 (N_5460,N_4455,N_3854);
or U5461 (N_5461,N_4380,N_3388);
and U5462 (N_5462,N_2839,N_3200);
nor U5463 (N_5463,N_2886,N_928);
and U5464 (N_5464,N_1930,N_1900);
nand U5465 (N_5465,N_4706,N_2441);
nand U5466 (N_5466,N_1824,N_2717);
and U5467 (N_5467,N_2876,N_275);
or U5468 (N_5468,N_344,N_98);
or U5469 (N_5469,N_4799,N_2474);
nand U5470 (N_5470,N_4193,N_3353);
and U5471 (N_5471,N_4208,N_3170);
nor U5472 (N_5472,N_94,N_18);
and U5473 (N_5473,N_1427,N_2479);
xor U5474 (N_5474,N_3149,N_3790);
nor U5475 (N_5475,N_4183,N_3980);
and U5476 (N_5476,N_4093,N_4480);
nand U5477 (N_5477,N_20,N_4061);
nand U5478 (N_5478,N_4593,N_2872);
or U5479 (N_5479,N_756,N_2128);
nor U5480 (N_5480,N_3112,N_3378);
and U5481 (N_5481,N_2999,N_1287);
or U5482 (N_5482,N_1036,N_1094);
or U5483 (N_5483,N_3400,N_1013);
or U5484 (N_5484,N_3639,N_4636);
and U5485 (N_5485,N_3652,N_3227);
and U5486 (N_5486,N_611,N_2030);
xnor U5487 (N_5487,N_3597,N_3452);
nor U5488 (N_5488,N_2486,N_2244);
and U5489 (N_5489,N_4127,N_65);
or U5490 (N_5490,N_3667,N_3943);
and U5491 (N_5491,N_4745,N_1361);
nand U5492 (N_5492,N_4339,N_4104);
or U5493 (N_5493,N_3128,N_1370);
nand U5494 (N_5494,N_2933,N_2909);
or U5495 (N_5495,N_257,N_3833);
nand U5496 (N_5496,N_2389,N_3737);
nor U5497 (N_5497,N_1374,N_1046);
nand U5498 (N_5498,N_4999,N_2009);
or U5499 (N_5499,N_873,N_4201);
nand U5500 (N_5500,N_665,N_999);
nand U5501 (N_5501,N_4881,N_647);
xor U5502 (N_5502,N_2790,N_4904);
and U5503 (N_5503,N_1624,N_3682);
or U5504 (N_5504,N_2133,N_4862);
nor U5505 (N_5505,N_2084,N_4003);
and U5506 (N_5506,N_1843,N_2945);
xor U5507 (N_5507,N_5,N_606);
nand U5508 (N_5508,N_855,N_1916);
or U5509 (N_5509,N_2493,N_953);
nor U5510 (N_5510,N_4672,N_3173);
or U5511 (N_5511,N_4558,N_2617);
xnor U5512 (N_5512,N_3497,N_615);
or U5513 (N_5513,N_4364,N_1623);
or U5514 (N_5514,N_2379,N_1159);
xor U5515 (N_5515,N_3101,N_3357);
nor U5516 (N_5516,N_1222,N_314);
or U5517 (N_5517,N_4460,N_2736);
nand U5518 (N_5518,N_838,N_4667);
or U5519 (N_5519,N_4561,N_1175);
or U5520 (N_5520,N_448,N_2538);
nand U5521 (N_5521,N_651,N_1934);
and U5522 (N_5522,N_41,N_1198);
xor U5523 (N_5523,N_759,N_3167);
nor U5524 (N_5524,N_1256,N_3005);
or U5525 (N_5525,N_3123,N_684);
or U5526 (N_5526,N_3773,N_4601);
xnor U5527 (N_5527,N_2121,N_19);
and U5528 (N_5528,N_3974,N_3252);
nor U5529 (N_5529,N_2079,N_1630);
or U5530 (N_5530,N_2321,N_4942);
nand U5531 (N_5531,N_4521,N_4614);
nor U5532 (N_5532,N_2811,N_2953);
nand U5533 (N_5533,N_3453,N_3520);
or U5534 (N_5534,N_4280,N_1116);
and U5535 (N_5535,N_313,N_4699);
or U5536 (N_5536,N_2897,N_600);
and U5537 (N_5537,N_4054,N_423);
nor U5538 (N_5538,N_501,N_1593);
or U5539 (N_5539,N_4606,N_3457);
nand U5540 (N_5540,N_4570,N_2301);
nor U5541 (N_5541,N_3272,N_2623);
and U5542 (N_5542,N_1398,N_1928);
xnor U5543 (N_5543,N_605,N_1557);
nor U5544 (N_5544,N_1860,N_1151);
and U5545 (N_5545,N_1471,N_608);
nor U5546 (N_5546,N_4582,N_2576);
nor U5547 (N_5547,N_764,N_2890);
nand U5548 (N_5548,N_3941,N_775);
nor U5549 (N_5549,N_4135,N_249);
xor U5550 (N_5550,N_1589,N_2840);
or U5551 (N_5551,N_2748,N_1058);
and U5552 (N_5552,N_3217,N_1718);
and U5553 (N_5553,N_2073,N_2525);
nor U5554 (N_5554,N_3027,N_619);
and U5555 (N_5555,N_3853,N_2306);
and U5556 (N_5556,N_2930,N_4922);
nor U5557 (N_5557,N_3776,N_4346);
nand U5558 (N_5558,N_33,N_2193);
nand U5559 (N_5559,N_4649,N_1263);
nor U5560 (N_5560,N_563,N_905);
nor U5561 (N_5561,N_301,N_540);
nor U5562 (N_5562,N_3643,N_2071);
nor U5563 (N_5563,N_897,N_4637);
nand U5564 (N_5564,N_4197,N_2444);
or U5565 (N_5565,N_796,N_2215);
and U5566 (N_5566,N_2732,N_819);
xnor U5567 (N_5567,N_3611,N_2926);
nand U5568 (N_5568,N_4806,N_3650);
xnor U5569 (N_5569,N_659,N_3211);
or U5570 (N_5570,N_24,N_4360);
nor U5571 (N_5571,N_4987,N_2868);
nand U5572 (N_5572,N_1105,N_4734);
nor U5573 (N_5573,N_1154,N_4544);
nor U5574 (N_5574,N_2140,N_4341);
nand U5575 (N_5575,N_4092,N_1992);
xor U5576 (N_5576,N_4177,N_1258);
nand U5577 (N_5577,N_1634,N_4291);
nor U5578 (N_5578,N_2858,N_4529);
or U5579 (N_5579,N_545,N_794);
nand U5580 (N_5580,N_4647,N_827);
xor U5581 (N_5581,N_1678,N_3122);
nor U5582 (N_5582,N_4172,N_1274);
nand U5583 (N_5583,N_4549,N_1588);
xnor U5584 (N_5584,N_2387,N_844);
nor U5585 (N_5585,N_883,N_4082);
or U5586 (N_5586,N_2524,N_3504);
or U5587 (N_5587,N_4884,N_3015);
and U5588 (N_5588,N_332,N_683);
or U5589 (N_5589,N_4897,N_2621);
nor U5590 (N_5590,N_3166,N_3585);
nand U5591 (N_5591,N_4981,N_4140);
nor U5592 (N_5592,N_1576,N_1411);
nor U5593 (N_5593,N_4878,N_2508);
or U5594 (N_5594,N_2437,N_1713);
and U5595 (N_5595,N_1114,N_1476);
or U5596 (N_5596,N_3238,N_2979);
nor U5597 (N_5597,N_788,N_369);
or U5598 (N_5598,N_3110,N_2485);
nand U5599 (N_5599,N_1334,N_4256);
nand U5600 (N_5600,N_3878,N_3344);
or U5601 (N_5601,N_2070,N_3021);
or U5602 (N_5602,N_3447,N_847);
and U5603 (N_5603,N_1939,N_4085);
or U5604 (N_5604,N_4605,N_1244);
nand U5605 (N_5605,N_1788,N_2013);
or U5606 (N_5606,N_3522,N_396);
nor U5607 (N_5607,N_290,N_3646);
nand U5608 (N_5608,N_1356,N_3982);
nand U5609 (N_5609,N_3527,N_3746);
nand U5610 (N_5610,N_225,N_3674);
nand U5611 (N_5611,N_2517,N_4484);
nand U5612 (N_5612,N_433,N_4490);
nor U5613 (N_5613,N_3721,N_742);
nor U5614 (N_5614,N_2629,N_1813);
or U5615 (N_5615,N_2477,N_2904);
or U5616 (N_5616,N_1266,N_4289);
nor U5617 (N_5617,N_1727,N_4870);
nand U5618 (N_5618,N_2755,N_3351);
and U5619 (N_5619,N_3023,N_2459);
nor U5620 (N_5620,N_2867,N_1280);
xnor U5621 (N_5621,N_3011,N_2938);
nor U5622 (N_5622,N_4264,N_1724);
and U5623 (N_5623,N_1767,N_4012);
nand U5624 (N_5624,N_3855,N_2973);
nor U5625 (N_5625,N_14,N_2793);
nand U5626 (N_5626,N_2094,N_1290);
xor U5627 (N_5627,N_1601,N_2785);
nand U5628 (N_5628,N_1905,N_4305);
nor U5629 (N_5629,N_4144,N_1341);
nor U5630 (N_5630,N_1862,N_4368);
xnor U5631 (N_5631,N_473,N_1284);
nor U5632 (N_5632,N_1282,N_9);
or U5633 (N_5633,N_4263,N_2309);
nor U5634 (N_5634,N_2559,N_266);
nand U5635 (N_5635,N_3077,N_3610);
nor U5636 (N_5636,N_4218,N_1399);
and U5637 (N_5637,N_1991,N_2058);
and U5638 (N_5638,N_4122,N_1774);
xnor U5639 (N_5639,N_3993,N_2494);
or U5640 (N_5640,N_4243,N_4639);
nor U5641 (N_5641,N_1098,N_2065);
nand U5642 (N_5642,N_4492,N_1369);
nand U5643 (N_5643,N_2300,N_3168);
and U5644 (N_5644,N_4859,N_4644);
or U5645 (N_5645,N_3924,N_456);
nand U5646 (N_5646,N_62,N_478);
and U5647 (N_5647,N_1267,N_2855);
and U5648 (N_5648,N_3973,N_1078);
and U5649 (N_5649,N_2312,N_3640);
nand U5650 (N_5650,N_2880,N_2977);
and U5651 (N_5651,N_4361,N_203);
nor U5652 (N_5652,N_2279,N_2772);
xnor U5653 (N_5653,N_3577,N_2669);
nor U5654 (N_5654,N_4163,N_3427);
and U5655 (N_5655,N_1902,N_56);
nor U5656 (N_5656,N_3033,N_1621);
nor U5657 (N_5657,N_4398,N_3634);
nor U5658 (N_5658,N_2063,N_424);
nor U5659 (N_5659,N_660,N_3587);
or U5660 (N_5660,N_1644,N_4115);
nand U5661 (N_5661,N_3180,N_1192);
nand U5662 (N_5662,N_2518,N_4499);
or U5663 (N_5663,N_2012,N_3771);
nor U5664 (N_5664,N_4255,N_2510);
and U5665 (N_5665,N_466,N_2234);
xnor U5666 (N_5666,N_3376,N_4641);
nor U5667 (N_5667,N_2251,N_2952);
xnor U5668 (N_5668,N_1981,N_145);
or U5669 (N_5669,N_337,N_2758);
or U5670 (N_5670,N_1491,N_166);
and U5671 (N_5671,N_4202,N_1350);
or U5672 (N_5672,N_3072,N_3926);
nand U5673 (N_5673,N_58,N_280);
xnor U5674 (N_5674,N_1322,N_374);
or U5675 (N_5675,N_4986,N_3541);
nor U5676 (N_5676,N_3364,N_1729);
nand U5677 (N_5677,N_2769,N_4046);
nor U5678 (N_5678,N_3148,N_2531);
nor U5679 (N_5679,N_1400,N_949);
or U5680 (N_5680,N_1820,N_1725);
xor U5681 (N_5681,N_572,N_2792);
or U5682 (N_5682,N_595,N_1133);
nor U5683 (N_5683,N_2941,N_4212);
nand U5684 (N_5684,N_1020,N_2997);
or U5685 (N_5685,N_470,N_1801);
nor U5686 (N_5686,N_965,N_2435);
nand U5687 (N_5687,N_4869,N_2059);
nor U5688 (N_5688,N_607,N_36);
nand U5689 (N_5689,N_3529,N_48);
nand U5690 (N_5690,N_2136,N_4992);
or U5691 (N_5691,N_3712,N_4764);
nand U5692 (N_5692,N_2588,N_3695);
nor U5693 (N_5693,N_4711,N_3582);
nand U5694 (N_5694,N_910,N_1030);
nand U5695 (N_5695,N_1181,N_943);
and U5696 (N_5696,N_3852,N_4772);
nor U5697 (N_5697,N_4701,N_165);
nor U5698 (N_5698,N_2027,N_4511);
nor U5699 (N_5699,N_2983,N_1919);
or U5700 (N_5700,N_1935,N_4548);
and U5701 (N_5701,N_3209,N_3226);
or U5702 (N_5702,N_1684,N_418);
or U5703 (N_5703,N_4662,N_2614);
or U5704 (N_5704,N_717,N_3507);
or U5705 (N_5705,N_1230,N_1312);
and U5706 (N_5706,N_3019,N_4896);
nor U5707 (N_5707,N_1343,N_2568);
nand U5708 (N_5708,N_856,N_4452);
nor U5709 (N_5709,N_2836,N_3020);
nor U5710 (N_5710,N_1070,N_3897);
or U5711 (N_5711,N_3940,N_1806);
nand U5712 (N_5712,N_2304,N_1695);
nand U5713 (N_5713,N_1161,N_461);
xor U5714 (N_5714,N_1095,N_3054);
nor U5715 (N_5715,N_1348,N_1756);
xnor U5716 (N_5716,N_667,N_3750);
nand U5717 (N_5717,N_4314,N_4978);
nand U5718 (N_5718,N_2068,N_4686);
or U5719 (N_5719,N_4230,N_489);
xor U5720 (N_5720,N_4744,N_2147);
nand U5721 (N_5721,N_1904,N_4298);
nand U5722 (N_5722,N_4810,N_1446);
xor U5723 (N_5723,N_3710,N_836);
or U5724 (N_5724,N_482,N_1689);
nor U5725 (N_5725,N_1808,N_2303);
and U5726 (N_5726,N_372,N_339);
nand U5727 (N_5727,N_2779,N_4031);
or U5728 (N_5728,N_1710,N_3258);
or U5729 (N_5729,N_4473,N_3389);
nand U5730 (N_5730,N_1325,N_3756);
nor U5731 (N_5731,N_1856,N_1952);
nand U5732 (N_5732,N_4803,N_1944);
nor U5733 (N_5733,N_4181,N_1138);
nand U5734 (N_5734,N_4485,N_3354);
and U5735 (N_5735,N_4124,N_1690);
xor U5736 (N_5736,N_484,N_4015);
or U5737 (N_5737,N_1202,N_2994);
nand U5738 (N_5738,N_76,N_3233);
nor U5739 (N_5739,N_2406,N_4723);
or U5740 (N_5740,N_3997,N_4943);
nand U5741 (N_5741,N_1954,N_1156);
and U5742 (N_5742,N_1434,N_3214);
and U5743 (N_5743,N_1872,N_2804);
nor U5744 (N_5744,N_3815,N_400);
nor U5745 (N_5745,N_260,N_3636);
nand U5746 (N_5746,N_228,N_3338);
nand U5747 (N_5747,N_4287,N_1167);
nand U5748 (N_5748,N_3086,N_3703);
nand U5749 (N_5749,N_4657,N_4470);
nand U5750 (N_5750,N_1568,N_3693);
nand U5751 (N_5751,N_1223,N_4506);
nor U5752 (N_5752,N_1559,N_3071);
nand U5753 (N_5753,N_4032,N_1027);
nor U5754 (N_5754,N_1858,N_1416);
or U5755 (N_5755,N_1345,N_3843);
xnor U5756 (N_5756,N_3725,N_1486);
or U5757 (N_5757,N_1045,N_2372);
nor U5758 (N_5758,N_3733,N_2626);
and U5759 (N_5759,N_514,N_1751);
nor U5760 (N_5760,N_2431,N_4780);
nor U5761 (N_5761,N_3366,N_4834);
xnor U5762 (N_5762,N_324,N_2420);
and U5763 (N_5763,N_268,N_3010);
or U5764 (N_5764,N_3872,N_3848);
or U5765 (N_5765,N_4369,N_1255);
nor U5766 (N_5766,N_3764,N_2203);
nand U5767 (N_5767,N_636,N_1781);
and U5768 (N_5768,N_1299,N_2248);
nor U5769 (N_5769,N_3874,N_4342);
and U5770 (N_5770,N_1264,N_2696);
nor U5771 (N_5771,N_2781,N_4464);
nor U5772 (N_5772,N_2018,N_388);
or U5773 (N_5773,N_3456,N_2718);
and U5774 (N_5774,N_2074,N_3050);
and U5775 (N_5775,N_3953,N_1798);
nor U5776 (N_5776,N_529,N_491);
nor U5777 (N_5777,N_213,N_4058);
and U5778 (N_5778,N_2505,N_2735);
and U5779 (N_5779,N_4379,N_1472);
or U5780 (N_5780,N_4141,N_4634);
and U5781 (N_5781,N_633,N_719);
and U5782 (N_5782,N_3705,N_4678);
nand U5783 (N_5783,N_2004,N_1044);
nor U5784 (N_5784,N_1785,N_3393);
xor U5785 (N_5785,N_4487,N_399);
nor U5786 (N_5786,N_4883,N_4259);
nor U5787 (N_5787,N_4371,N_1564);
xnor U5788 (N_5788,N_261,N_2138);
or U5789 (N_5789,N_4023,N_2239);
and U5790 (N_5790,N_4221,N_4347);
nor U5791 (N_5791,N_2589,N_3174);
and U5792 (N_5792,N_4785,N_247);
nand U5793 (N_5793,N_3032,N_779);
or U5794 (N_5794,N_4130,N_4827);
or U5795 (N_5795,N_3437,N_4898);
nor U5796 (N_5796,N_1699,N_2856);
or U5797 (N_5797,N_146,N_4839);
and U5798 (N_5798,N_3279,N_4421);
nor U5799 (N_5799,N_918,N_1102);
xor U5800 (N_5800,N_1466,N_1560);
and U5801 (N_5801,N_2241,N_4938);
nor U5802 (N_5802,N_3461,N_1049);
and U5803 (N_5803,N_2424,N_3245);
and U5804 (N_5804,N_3002,N_1265);
or U5805 (N_5805,N_1783,N_4796);
and U5806 (N_5806,N_553,N_3515);
nor U5807 (N_5807,N_1933,N_1023);
nor U5808 (N_5808,N_2190,N_2223);
and U5809 (N_5809,N_2080,N_357);
nand U5810 (N_5810,N_3066,N_523);
or U5811 (N_5811,N_1443,N_1611);
nand U5812 (N_5812,N_1451,N_808);
or U5813 (N_5813,N_1153,N_1243);
nor U5814 (N_5814,N_2544,N_1754);
nor U5815 (N_5815,N_3429,N_4123);
nor U5816 (N_5816,N_2743,N_4382);
and U5817 (N_5817,N_2896,N_2603);
or U5818 (N_5818,N_2928,N_2419);
nor U5819 (N_5819,N_322,N_4607);
nand U5820 (N_5820,N_4590,N_2705);
nand U5821 (N_5821,N_230,N_1009);
and U5822 (N_5822,N_517,N_3285);
xnor U5823 (N_5823,N_853,N_4910);
xnor U5824 (N_5824,N_1082,N_2362);
nor U5825 (N_5825,N_236,N_1573);
or U5826 (N_5826,N_1237,N_1534);
nand U5827 (N_5827,N_3669,N_2853);
nor U5828 (N_5828,N_3945,N_2290);
and U5829 (N_5829,N_4258,N_1272);
nand U5830 (N_5830,N_3816,N_4691);
or U5831 (N_5831,N_2446,N_2164);
and U5832 (N_5832,N_92,N_1759);
nand U5833 (N_5833,N_1304,N_2454);
nand U5834 (N_5834,N_1248,N_765);
or U5835 (N_5835,N_2992,N_1317);
nand U5836 (N_5836,N_3451,N_190);
or U5837 (N_5837,N_4217,N_4180);
or U5838 (N_5838,N_3502,N_2942);
nor U5839 (N_5839,N_1184,N_2440);
xnor U5840 (N_5840,N_3911,N_3365);
and U5841 (N_5841,N_1885,N_2512);
nor U5842 (N_5842,N_2052,N_3130);
and U5843 (N_5843,N_2733,N_4441);
and U5844 (N_5844,N_2330,N_11);
xnor U5845 (N_5845,N_4131,N_906);
and U5846 (N_5846,N_4640,N_1738);
or U5847 (N_5847,N_1875,N_4555);
nand U5848 (N_5848,N_526,N_4914);
or U5849 (N_5849,N_4277,N_214);
nand U5850 (N_5850,N_1390,N_4523);
or U5851 (N_5851,N_4286,N_2149);
and U5852 (N_5852,N_3658,N_675);
nand U5853 (N_5853,N_2670,N_2156);
nor U5854 (N_5854,N_3304,N_2892);
nand U5855 (N_5855,N_2348,N_2943);
nand U5856 (N_5856,N_4472,N_105);
and U5857 (N_5857,N_3907,N_3480);
and U5858 (N_5858,N_2571,N_3524);
or U5859 (N_5859,N_3893,N_2891);
nand U5860 (N_5860,N_2339,N_3732);
or U5861 (N_5861,N_2762,N_1682);
and U5862 (N_5862,N_341,N_4714);
and U5863 (N_5863,N_3537,N_2749);
and U5864 (N_5864,N_1331,N_487);
nor U5865 (N_5865,N_2275,N_2229);
xnor U5866 (N_5866,N_3641,N_4383);
nor U5867 (N_5867,N_956,N_1447);
nor U5868 (N_5868,N_1647,N_661);
and U5869 (N_5869,N_171,N_4386);
nor U5870 (N_5870,N_4483,N_1482);
and U5871 (N_5871,N_3052,N_2955);
nor U5872 (N_5872,N_2766,N_2476);
nand U5873 (N_5873,N_136,N_4991);
nand U5874 (N_5874,N_1575,N_3051);
and U5875 (N_5875,N_1587,N_1651);
nor U5876 (N_5876,N_1257,N_2259);
nand U5877 (N_5877,N_2752,N_1377);
or U5878 (N_5878,N_2037,N_3454);
nor U5879 (N_5879,N_320,N_4486);
nand U5880 (N_5880,N_3799,N_160);
nand U5881 (N_5881,N_800,N_1816);
xnor U5882 (N_5882,N_1591,N_4783);
nor U5883 (N_5883,N_4417,N_1812);
nor U5884 (N_5884,N_2829,N_2863);
nor U5885 (N_5885,N_2851,N_2616);
xnor U5886 (N_5886,N_3987,N_3889);
nor U5887 (N_5887,N_4145,N_2573);
nor U5888 (N_5888,N_4057,N_1429);
and U5889 (N_5889,N_805,N_1949);
nor U5890 (N_5890,N_2923,N_754);
and U5891 (N_5891,N_4071,N_350);
nand U5892 (N_5892,N_3423,N_1177);
nor U5893 (N_5893,N_1652,N_3921);
nor U5894 (N_5894,N_422,N_3155);
or U5895 (N_5895,N_2363,N_2393);
nor U5896 (N_5896,N_1716,N_3692);
nor U5897 (N_5897,N_2,N_4626);
nor U5898 (N_5898,N_3029,N_978);
nor U5899 (N_5899,N_4171,N_743);
nor U5900 (N_5900,N_3241,N_2255);
or U5901 (N_5901,N_863,N_2740);
and U5902 (N_5902,N_107,N_2878);
or U5903 (N_5903,N_2707,N_3387);
or U5904 (N_5904,N_3339,N_2101);
nand U5905 (N_5905,N_4191,N_3282);
and U5906 (N_5906,N_2980,N_3363);
or U5907 (N_5907,N_3752,N_3755);
nand U5908 (N_5908,N_4899,N_2591);
nand U5909 (N_5909,N_1546,N_4276);
xor U5910 (N_5910,N_521,N_3127);
or U5911 (N_5911,N_3970,N_306);
nor U5912 (N_5912,N_4036,N_460);
nor U5913 (N_5913,N_751,N_4911);
or U5914 (N_5914,N_1052,N_3210);
and U5915 (N_5915,N_4224,N_2409);
and U5916 (N_5916,N_4530,N_3781);
nand U5917 (N_5917,N_859,N_2449);
and U5918 (N_5918,N_3649,N_3784);
nand U5919 (N_5919,N_4787,N_1607);
nand U5920 (N_5920,N_3699,N_1004);
nand U5921 (N_5921,N_4751,N_4121);
and U5922 (N_5922,N_3159,N_3169);
nor U5923 (N_5923,N_932,N_4358);
nor U5924 (N_5924,N_1413,N_1307);
nor U5925 (N_5925,N_4988,N_3890);
or U5926 (N_5926,N_4384,N_1011);
and U5927 (N_5927,N_3316,N_2471);
xor U5928 (N_5928,N_3567,N_1245);
xor U5929 (N_5929,N_3717,N_1772);
nand U5930 (N_5930,N_3793,N_1519);
xor U5931 (N_5931,N_4002,N_4136);
and U5932 (N_5932,N_205,N_4161);
and U5933 (N_5933,N_2768,N_3257);
and U5934 (N_5934,N_4427,N_1789);
nor U5935 (N_5935,N_499,N_1594);
nor U5936 (N_5936,N_3385,N_2319);
and U5937 (N_5937,N_2134,N_53);
or U5938 (N_5938,N_4324,N_2922);
nand U5939 (N_5939,N_4909,N_1802);
or U5940 (N_5940,N_4886,N_1351);
or U5941 (N_5941,N_4742,N_2092);
or U5942 (N_5942,N_3589,N_4777);
or U5943 (N_5943,N_4929,N_93);
and U5944 (N_5944,N_4429,N_1613);
nor U5945 (N_5945,N_333,N_1971);
and U5946 (N_5946,N_2355,N_2286);
or U5947 (N_5947,N_4027,N_1505);
and U5948 (N_5948,N_1675,N_2115);
nor U5949 (N_5949,N_4419,N_2548);
nor U5950 (N_5950,N_989,N_3154);
xnor U5951 (N_5951,N_2808,N_1396);
nor U5952 (N_5952,N_1659,N_583);
and U5953 (N_5953,N_749,N_2050);
nor U5954 (N_5954,N_2438,N_3521);
and U5955 (N_5955,N_994,N_3111);
and U5956 (N_5956,N_480,N_1851);
or U5957 (N_5957,N_404,N_3553);
nand U5958 (N_5958,N_2651,N_1822);
or U5959 (N_5959,N_3121,N_4106);
nor U5960 (N_5960,N_4908,N_4072);
or U5961 (N_5961,N_2144,N_944);
nand U5962 (N_5962,N_2212,N_4648);
xor U5963 (N_5963,N_2676,N_1388);
xor U5964 (N_5964,N_2044,N_2278);
and U5965 (N_5965,N_2844,N_4856);
or U5966 (N_5966,N_957,N_2318);
and U5967 (N_5967,N_4435,N_3229);
nor U5968 (N_5968,N_903,N_4633);
nand U5969 (N_5969,N_2713,N_3260);
xnor U5970 (N_5970,N_4418,N_318);
nand U5971 (N_5971,N_3424,N_3728);
and U5972 (N_5972,N_1308,N_2196);
nand U5973 (N_5973,N_3540,N_3335);
nor U5974 (N_5974,N_4906,N_1166);
nor U5975 (N_5975,N_1974,N_476);
and U5976 (N_5976,N_2981,N_2706);
nor U5977 (N_5977,N_4893,N_3549);
and U5978 (N_5978,N_4704,N_3749);
nor U5979 (N_5979,N_2783,N_1253);
and U5980 (N_5980,N_2738,N_3346);
nor U5981 (N_5981,N_3951,N_1441);
nand U5982 (N_5982,N_4327,N_1545);
nor U5983 (N_5983,N_2690,N_1477);
nor U5984 (N_5984,N_4566,N_1604);
nor U5985 (N_5985,N_188,N_4066);
nand U5986 (N_5986,N_4185,N_3820);
or U5987 (N_5987,N_3811,N_2139);
nor U5988 (N_5988,N_2704,N_4019);
nand U5989 (N_5989,N_4320,N_4821);
nor U5990 (N_5990,N_4832,N_2774);
nand U5991 (N_5991,N_542,N_414);
or U5992 (N_5992,N_1119,N_1275);
nor U5993 (N_5993,N_4842,N_293);
and U5994 (N_5994,N_1422,N_148);
nor U5995 (N_5995,N_4117,N_3362);
or U5996 (N_5996,N_1238,N_1402);
nand U5997 (N_5997,N_830,N_1506);
or U5998 (N_5998,N_2826,N_3419);
and U5999 (N_5999,N_2467,N_643);
xnor U6000 (N_6000,N_3609,N_8);
nor U6001 (N_6001,N_4591,N_782);
and U6002 (N_6002,N_4504,N_3330);
nand U6003 (N_6003,N_3952,N_2109);
nor U6004 (N_6004,N_1522,N_533);
or U6005 (N_6005,N_1687,N_1876);
nor U6006 (N_6006,N_1686,N_1542);
or U6007 (N_6007,N_3491,N_3594);
xnor U6008 (N_6008,N_3176,N_530);
nor U6009 (N_6009,N_677,N_3691);
and U6010 (N_6010,N_1214,N_1205);
or U6011 (N_6011,N_556,N_4594);
nor U6012 (N_6012,N_4307,N_2302);
or U6013 (N_6013,N_2877,N_1869);
nor U6014 (N_6014,N_4567,N_4045);
and U6015 (N_6015,N_51,N_3367);
xnor U6016 (N_6016,N_4038,N_2967);
and U6017 (N_6017,N_584,N_3876);
nor U6018 (N_6018,N_4182,N_175);
nor U6019 (N_6019,N_790,N_4080);
nand U6020 (N_6020,N_84,N_1959);
and U6021 (N_6021,N_1878,N_398);
or U6022 (N_6022,N_3137,N_3648);
or U6023 (N_6023,N_4090,N_4424);
and U6024 (N_6024,N_2323,N_2127);
or U6025 (N_6025,N_3004,N_1926);
nand U6026 (N_6026,N_4426,N_1676);
and U6027 (N_6027,N_3091,N_3555);
and U6028 (N_6028,N_846,N_2066);
nand U6029 (N_6029,N_237,N_2374);
and U6030 (N_6030,N_2172,N_3526);
xor U6031 (N_6031,N_50,N_930);
and U6032 (N_6032,N_3283,N_4581);
nor U6033 (N_6033,N_2351,N_2307);
nand U6034 (N_6034,N_2847,N_1005);
xor U6035 (N_6035,N_204,N_4040);
and U6036 (N_6036,N_4375,N_438);
nand U6037 (N_6037,N_4885,N_952);
and U6038 (N_6038,N_3581,N_252);
nor U6039 (N_6039,N_3477,N_3904);
nor U6040 (N_6040,N_477,N_277);
nor U6041 (N_6041,N_241,N_1556);
or U6042 (N_6042,N_2370,N_2394);
nand U6043 (N_6043,N_733,N_1910);
and U6044 (N_6044,N_2580,N_4321);
nand U6045 (N_6045,N_3627,N_3183);
or U6046 (N_6046,N_143,N_3059);
nor U6047 (N_6047,N_1421,N_200);
nor U6048 (N_6048,N_4211,N_1666);
nor U6049 (N_6049,N_3635,N_1259);
and U6050 (N_6050,N_991,N_2183);
and U6051 (N_6051,N_1295,N_170);
or U6052 (N_6052,N_2949,N_4069);
and U6053 (N_6053,N_2240,N_865);
or U6054 (N_6054,N_2686,N_1976);
nand U6055 (N_6055,N_1641,N_2209);
nor U6056 (N_6056,N_1664,N_1958);
and U6057 (N_6057,N_3601,N_984);
or U6058 (N_6058,N_1453,N_492);
xor U6059 (N_6059,N_462,N_3062);
nand U6060 (N_6060,N_67,N_2633);
nor U6061 (N_6061,N_57,N_1145);
nor U6062 (N_6062,N_2784,N_4894);
and U6063 (N_6063,N_316,N_2296);
or U6064 (N_6064,N_2422,N_2167);
xnor U6065 (N_6065,N_3894,N_1479);
or U6066 (N_6066,N_4900,N_4365);
nor U6067 (N_6067,N_936,N_2346);
xnor U6068 (N_6068,N_935,N_397);
and U6069 (N_6069,N_1281,N_4828);
and U6070 (N_6070,N_1247,N_783);
nand U6071 (N_6071,N_3979,N_283);
or U6072 (N_6072,N_1886,N_3726);
nand U6073 (N_6073,N_3698,N_1366);
nand U6074 (N_6074,N_3711,N_3228);
nor U6075 (N_6075,N_1987,N_3340);
nor U6076 (N_6076,N_1883,N_3929);
or U6077 (N_6077,N_650,N_4948);
or U6078 (N_6078,N_447,N_4746);
nand U6079 (N_6079,N_3948,N_4575);
or U6080 (N_6080,N_4436,N_1513);
and U6081 (N_6081,N_3913,N_3617);
nand U6082 (N_6082,N_1019,N_4921);
and U6083 (N_6083,N_1124,N_3470);
nor U6084 (N_6084,N_1384,N_3761);
xnor U6085 (N_6085,N_4829,N_1221);
nor U6086 (N_6086,N_1925,N_945);
nor U6087 (N_6087,N_1452,N_4405);
nor U6088 (N_6088,N_3095,N_2036);
or U6089 (N_6089,N_673,N_4134);
nor U6090 (N_6090,N_577,N_1895);
nand U6091 (N_6091,N_4748,N_99);
nor U6092 (N_6092,N_520,N_375);
nand U6093 (N_6093,N_3000,N_1246);
or U6094 (N_6094,N_1160,N_3370);
xor U6095 (N_6095,N_1977,N_216);
or U6096 (N_6096,N_444,N_1953);
nor U6097 (N_6097,N_613,N_2543);
and U6098 (N_6098,N_2496,N_3628);
or U6099 (N_6099,N_3390,N_4397);
and U6100 (N_6100,N_3266,N_3838);
or U6101 (N_6101,N_3831,N_3094);
and U6102 (N_6102,N_2273,N_3432);
nand U6103 (N_6103,N_3489,N_2095);
or U6104 (N_6104,N_503,N_3939);
nand U6105 (N_6105,N_4293,N_4113);
or U6106 (N_6106,N_2597,N_4798);
or U6107 (N_6107,N_2529,N_4703);
nand U6108 (N_6108,N_3867,N_2818);
xor U6109 (N_6109,N_3488,N_971);
nand U6110 (N_6110,N_4103,N_4963);
nor U6111 (N_6111,N_2069,N_543);
nor U6112 (N_6112,N_4632,N_125);
nor U6113 (N_6113,N_4478,N_3576);
nor U6114 (N_6114,N_3672,N_688);
or U6115 (N_6115,N_4322,N_4016);
nand U6116 (N_6116,N_950,N_3207);
nor U6117 (N_6117,N_3108,N_1674);
nor U6118 (N_6118,N_2465,N_2971);
nand U6119 (N_6119,N_4860,N_85);
nor U6120 (N_6120,N_4420,N_2960);
xor U6121 (N_6121,N_4194,N_2763);
xor U6122 (N_6122,N_2247,N_3359);
nor U6123 (N_6123,N_59,N_439);
nor U6124 (N_6124,N_2834,N_2773);
and U6125 (N_6125,N_4162,N_2253);
nor U6126 (N_6126,N_575,N_1749);
nand U6127 (N_6127,N_3253,N_1201);
nor U6128 (N_6128,N_3999,N_2948);
or U6129 (N_6129,N_297,N_3034);
or U6130 (N_6130,N_1335,N_1484);
or U6131 (N_6131,N_3936,N_938);
and U6132 (N_6132,N_1932,N_3783);
or U6133 (N_6133,N_2429,N_4042);
nand U6134 (N_6134,N_768,N_3116);
xor U6135 (N_6135,N_3996,N_4546);
nor U6136 (N_6136,N_1891,N_459);
or U6137 (N_6137,N_1565,N_1985);
nor U6138 (N_6138,N_4312,N_666);
nor U6139 (N_6139,N_3840,N_1968);
and U6140 (N_6140,N_3243,N_966);
nor U6141 (N_6141,N_2481,N_631);
and U6142 (N_6142,N_569,N_587);
and U6143 (N_6143,N_748,N_1967);
and U6144 (N_6144,N_512,N_4627);
and U6145 (N_6145,N_3156,N_256);
and U6146 (N_6146,N_1164,N_3061);
or U6147 (N_6147,N_1487,N_2866);
and U6148 (N_6148,N_2906,N_638);
and U6149 (N_6149,N_4524,N_825);
xor U6150 (N_6150,N_1739,N_343);
or U6151 (N_6151,N_3946,N_746);
nor U6152 (N_6152,N_721,N_1504);
nand U6153 (N_6153,N_1212,N_209);
nor U6154 (N_6154,N_2605,N_96);
xnor U6155 (N_6155,N_1001,N_3992);
or U6156 (N_6156,N_6,N_2231);
nor U6157 (N_6157,N_2959,N_101);
nand U6158 (N_6158,N_4086,N_2198);
nor U6159 (N_6159,N_3464,N_852);
and U6160 (N_6160,N_4927,N_548);
nand U6161 (N_6161,N_3224,N_3622);
nor U6162 (N_6162,N_1627,N_3778);
or U6163 (N_6163,N_390,N_2106);
nor U6164 (N_6164,N_955,N_1127);
nand U6165 (N_6165,N_1229,N_921);
and U6166 (N_6166,N_1185,N_4585);
xnor U6167 (N_6167,N_304,N_1139);
nand U6168 (N_6168,N_299,N_2099);
xnor U6169 (N_6169,N_127,N_1191);
nand U6170 (N_6170,N_3495,N_3753);
nand U6171 (N_6171,N_4308,N_2464);
nand U6172 (N_6172,N_4006,N_2265);
nor U6173 (N_6173,N_922,N_3689);
and U6174 (N_6174,N_1368,N_2397);
or U6175 (N_6175,N_2530,N_3696);
or U6176 (N_6176,N_2383,N_2618);
and U6177 (N_6177,N_3162,N_1865);
and U6178 (N_6178,N_0,N_4353);
nor U6179 (N_6179,N_3164,N_894);
or U6180 (N_6180,N_1752,N_192);
or U6181 (N_6181,N_179,N_2536);
and U6182 (N_6182,N_911,N_4781);
and U6183 (N_6183,N_4089,N_2745);
and U6184 (N_6184,N_1765,N_515);
xor U6185 (N_6185,N_2457,N_4795);
or U6186 (N_6186,N_4520,N_4941);
nand U6187 (N_6187,N_3105,N_3371);
nor U6188 (N_6188,N_4030,N_1392);
nand U6189 (N_6189,N_3334,N_912);
and U6190 (N_6190,N_2408,N_3158);
and U6191 (N_6191,N_4915,N_286);
or U6192 (N_6192,N_255,N_874);
nand U6193 (N_6193,N_2604,N_454);
nand U6194 (N_6194,N_4290,N_692);
xor U6195 (N_6195,N_1298,N_626);
and U6196 (N_6196,N_3985,N_3001);
or U6197 (N_6197,N_1957,N_3686);
or U6198 (N_6198,N_496,N_2230);
nor U6199 (N_6199,N_2898,N_4508);
and U6200 (N_6200,N_1053,N_2432);
xnor U6201 (N_6201,N_1464,N_2023);
nand U6202 (N_6202,N_697,N_552);
nand U6203 (N_6203,N_588,N_728);
and U6204 (N_6204,N_4536,N_1606);
and U6205 (N_6205,N_726,N_1679);
and U6206 (N_6206,N_210,N_1104);
and U6207 (N_6207,N_61,N_1147);
or U6208 (N_6208,N_1635,N_3554);
xnor U6209 (N_6209,N_2414,N_564);
or U6210 (N_6210,N_421,N_292);
or U6211 (N_6211,N_2819,N_763);
nor U6212 (N_6212,N_3616,N_3510);
or U6213 (N_6213,N_1584,N_81);
and U6214 (N_6214,N_4495,N_2837);
nand U6215 (N_6215,N_2956,N_3455);
nor U6216 (N_6216,N_2527,N_2016);
nor U6217 (N_6217,N_3600,N_1420);
nand U6218 (N_6218,N_377,N_2715);
nor U6219 (N_6219,N_1683,N_1360);
xor U6220 (N_6220,N_2641,N_3280);
xnor U6221 (N_6221,N_1498,N_2357);
nor U6222 (N_6222,N_1723,N_3197);
xnor U6223 (N_6223,N_4325,N_2523);
or U6224 (N_6224,N_2862,N_1410);
and U6225 (N_6225,N_31,N_2181);
nand U6226 (N_6226,N_3971,N_3327);
or U6227 (N_6227,N_1577,N_931);
or U6228 (N_6228,N_4296,N_4081);
nand U6229 (N_6229,N_4150,N_1310);
or U6230 (N_6230,N_1269,N_2907);
and U6231 (N_6231,N_298,N_1435);
and U6232 (N_6232,N_704,N_1236);
or U6233 (N_6233,N_2475,N_3647);
nor U6234 (N_6234,N_2124,N_3538);
nand U6235 (N_6235,N_993,N_1743);
or U6236 (N_6236,N_4867,N_934);
or U6237 (N_6237,N_3221,N_3250);
xnor U6238 (N_6238,N_155,N_1609);
and U6239 (N_6239,N_21,N_2542);
or U6240 (N_6240,N_1029,N_4376);
nor U6241 (N_6241,N_708,N_1826);
nand U6242 (N_6242,N_3273,N_2407);
nand U6243 (N_6243,N_4275,N_3096);
nor U6244 (N_6244,N_1123,N_4240);
and U6245 (N_6245,N_1879,N_4332);
or U6246 (N_6246,N_2123,N_3834);
xor U6247 (N_6247,N_233,N_2716);
nand U6248 (N_6248,N_367,N_4562);
nor U6249 (N_6249,N_3297,N_4288);
nand U6250 (N_6250,N_4395,N_3264);
nand U6251 (N_6251,N_1747,N_1996);
and U6252 (N_6252,N_4951,N_2995);
or U6253 (N_6253,N_4316,N_4005);
and U6254 (N_6254,N_1301,N_4569);
nand U6255 (N_6255,N_4840,N_1358);
or U6256 (N_6256,N_2143,N_4167);
nand U6257 (N_6257,N_1130,N_2765);
nand U6258 (N_6258,N_4964,N_3950);
or U6259 (N_6259,N_510,N_941);
nor U6260 (N_6260,N_2391,N_1786);
nand U6261 (N_6261,N_458,N_1088);
nor U6262 (N_6262,N_2802,N_4982);
nand U6263 (N_6263,N_338,N_4568);
xnor U6264 (N_6264,N_1837,N_678);
or U6265 (N_6265,N_1726,N_1532);
nand U6266 (N_6266,N_3064,N_69);
or U6267 (N_6267,N_3892,N_2108);
nand U6268 (N_6268,N_1344,N_1551);
or U6269 (N_6269,N_2039,N_331);
or U6270 (N_6270,N_834,N_2246);
nor U6271 (N_6271,N_2060,N_4);
nor U6272 (N_6272,N_2969,N_1796);
nand U6273 (N_6273,N_3900,N_262);
or U6274 (N_6274,N_3079,N_4062);
nor U6275 (N_6275,N_1888,N_4912);
nand U6276 (N_6276,N_1884,N_2944);
or U6277 (N_6277,N_4753,N_2727);
or U6278 (N_6278,N_2987,N_741);
or U6279 (N_6279,N_1994,N_288);
nand U6280 (N_6280,N_1182,N_3918);
and U6281 (N_6281,N_4577,N_4766);
nor U6282 (N_6282,N_1662,N_2750);
and U6283 (N_6283,N_4835,N_1567);
or U6284 (N_6284,N_793,N_1025);
or U6285 (N_6285,N_3720,N_4618);
xnor U6286 (N_6286,N_2367,N_914);
nor U6287 (N_6287,N_144,N_3152);
nand U6288 (N_6288,N_2921,N_2984);
nor U6289 (N_6289,N_822,N_4876);
nor U6290 (N_6290,N_3070,N_3165);
nor U6291 (N_6291,N_789,N_3927);
and U6292 (N_6292,N_1533,N_3172);
nand U6293 (N_6293,N_4532,N_968);
or U6294 (N_6294,N_3312,N_1279);
and U6295 (N_6295,N_870,N_3560);
nor U6296 (N_6296,N_3198,N_1041);
nand U6297 (N_6297,N_2049,N_2918);
and U6298 (N_6298,N_3916,N_1979);
nand U6299 (N_6299,N_3901,N_4153);
and U6300 (N_6300,N_1889,N_2258);
nor U6301 (N_6301,N_38,N_1758);
and U6302 (N_6302,N_4475,N_1972);
nor U6303 (N_6303,N_4654,N_2550);
or U6304 (N_6304,N_806,N_2541);
and U6305 (N_6305,N_4688,N_287);
and U6306 (N_6306,N_2035,N_3602);
or U6307 (N_6307,N_2630,N_3508);
and U6308 (N_6308,N_3150,N_4004);
and U6309 (N_6309,N_4354,N_1073);
nand U6310 (N_6310,N_2107,N_850);
or U6311 (N_6311,N_4014,N_3516);
nor U6312 (N_6312,N_2089,N_4128);
nand U6313 (N_6313,N_2380,N_1887);
nor U6314 (N_6314,N_804,N_117);
or U6315 (N_6315,N_3496,N_4595);
xor U6316 (N_6316,N_381,N_3201);
nand U6317 (N_6317,N_4048,N_1964);
nor U6318 (N_6318,N_135,N_528);
or U6319 (N_6319,N_580,N_3666);
nand U6320 (N_6320,N_3917,N_2034);
xnor U6321 (N_6321,N_2213,N_1703);
nor U6322 (N_6322,N_3659,N_226);
and U6323 (N_6323,N_933,N_2160);
or U6324 (N_6324,N_1643,N_2041);
or U6325 (N_6325,N_1720,N_3277);
or U6326 (N_6326,N_3739,N_3730);
and U6327 (N_6327,N_3676,N_1818);
or U6328 (N_6328,N_4035,N_2153);
nand U6329 (N_6329,N_823,N_40);
nand U6330 (N_6330,N_88,N_4022);
nor U6331 (N_6331,N_3860,N_1750);
nand U6332 (N_6332,N_4450,N_3991);
nor U6333 (N_6333,N_2382,N_4522);
or U6334 (N_6334,N_2741,N_2884);
nor U6335 (N_6335,N_4983,N_3823);
nand U6336 (N_6336,N_875,N_2570);
or U6337 (N_6337,N_3075,N_1372);
nand U6338 (N_6338,N_2105,N_4278);
nand U6339 (N_6339,N_3543,N_4598);
and U6340 (N_6340,N_2615,N_1688);
or U6341 (N_6341,N_2267,N_880);
nand U6342 (N_6342,N_1293,N_1286);
nand U6343 (N_6343,N_4849,N_1921);
nor U6344 (N_6344,N_465,N_3535);
nand U6345 (N_6345,N_2197,N_2096);
or U6346 (N_6346,N_133,N_1819);
nor U6347 (N_6347,N_3374,N_44);
nand U6348 (N_6348,N_3296,N_954);
nand U6349 (N_6349,N_2338,N_142);
nand U6350 (N_6350,N_118,N_4695);
nand U6351 (N_6351,N_2889,N_412);
and U6352 (N_6352,N_2083,N_1553);
and U6353 (N_6353,N_2206,N_1975);
xor U6354 (N_6354,N_3532,N_4967);
or U6355 (N_6355,N_1309,N_3684);
nor U6356 (N_6356,N_1672,N_1291);
nor U6357 (N_6357,N_393,N_882);
or U6358 (N_6358,N_3539,N_2905);
nand U6359 (N_6359,N_1753,N_3043);
nand U6360 (N_6360,N_940,N_1332);
or U6361 (N_6361,N_1942,N_4705);
nand U6362 (N_6362,N_4573,N_876);
nand U6363 (N_6363,N_2413,N_3714);
nor U6364 (N_6364,N_79,N_2656);
or U6365 (N_6365,N_4851,N_3384);
nand U6366 (N_6366,N_3861,N_712);
nor U6367 (N_6367,N_1839,N_2757);
or U6368 (N_6368,N_2687,N_4650);
nor U6369 (N_6369,N_3883,N_727);
or U6370 (N_6370,N_2497,N_2998);
nand U6371 (N_6371,N_555,N_3747);
nor U6372 (N_6372,N_4710,N_4273);
nand U6373 (N_6373,N_3729,N_700);
xnor U6374 (N_6374,N_3030,N_625);
nand U6375 (N_6375,N_2910,N_4152);
and U6376 (N_6376,N_4459,N_758);
and U6377 (N_6377,N_3930,N_559);
or U6378 (N_6378,N_1998,N_2635);
xnor U6379 (N_6379,N_3038,N_3754);
and U6380 (N_6380,N_3935,N_807);
or U6381 (N_6381,N_4105,N_1871);
nor U6382 (N_6382,N_2817,N_1076);
xor U6383 (N_6383,N_3236,N_2250);
and U6384 (N_6384,N_1707,N_358);
nor U6385 (N_6385,N_4328,N_1387);
and U6386 (N_6386,N_506,N_2917);
nor U6387 (N_6387,N_1795,N_1552);
and U6388 (N_6388,N_797,N_4985);
nand U6389 (N_6389,N_4096,N_2002);
and U6390 (N_6390,N_4622,N_1525);
or U6391 (N_6391,N_1475,N_1746);
xor U6392 (N_6392,N_1132,N_3459);
and U6393 (N_6393,N_1924,N_2297);
nand U6394 (N_6394,N_1142,N_2996);
and U6395 (N_6395,N_4271,N_2264);
and U6396 (N_6396,N_3595,N_4200);
and U6397 (N_6397,N_699,N_1661);
and U6398 (N_6398,N_1050,N_4184);
or U6399 (N_6399,N_4946,N_4133);
nand U6400 (N_6400,N_1605,N_3409);
nand U6401 (N_6401,N_1999,N_116);
or U6402 (N_6402,N_1978,N_2701);
or U6403 (N_6403,N_767,N_1463);
or U6404 (N_6404,N_1766,N_3321);
nand U6405 (N_6405,N_431,N_4170);
xor U6406 (N_6406,N_1817,N_405);
and U6407 (N_6407,N_2478,N_2776);
nand U6408 (N_6408,N_3629,N_2448);
nor U6409 (N_6409,N_4343,N_1031);
or U6410 (N_6410,N_596,N_1566);
nor U6411 (N_6411,N_3377,N_3573);
and U6412 (N_6412,N_1777,N_2722);
and U6413 (N_6413,N_2780,N_2033);
nand U6414 (N_6414,N_1850,N_4094);
and U6415 (N_6415,N_4996,N_1357);
or U6416 (N_6416,N_2986,N_871);
or U6417 (N_6417,N_354,N_3525);
or U6418 (N_6418,N_2725,N_4400);
nand U6419 (N_6419,N_4425,N_3775);
nor U6420 (N_6420,N_3967,N_4143);
and U6421 (N_6421,N_248,N_2129);
xnor U6422 (N_6422,N_3870,N_1333);
nand U6423 (N_6423,N_3213,N_4956);
nand U6424 (N_6424,N_676,N_282);
xor U6425 (N_6425,N_3638,N_235);
and U6426 (N_6426,N_1853,N_278);
or U6427 (N_6427,N_308,N_4303);
nor U6428 (N_6428,N_2132,N_2385);
nor U6429 (N_6429,N_3938,N_4556);
nand U6430 (N_6430,N_2557,N_1468);
and U6431 (N_6431,N_4924,N_2261);
xor U6432 (N_6432,N_4990,N_3439);
and U6433 (N_6433,N_2920,N_828);
nand U6434 (N_6434,N_4786,N_702);
nand U6435 (N_6435,N_1793,N_2171);
nor U6436 (N_6436,N_345,N_1490);
and U6437 (N_6437,N_2720,N_3373);
nor U6438 (N_6438,N_1764,N_4060);
and U6439 (N_6439,N_4958,N_963);
nor U6440 (N_6440,N_942,N_2712);
or U6441 (N_6441,N_106,N_4517);
nor U6442 (N_6442,N_1838,N_380);
nor U6443 (N_6443,N_1148,N_2340);
nor U6444 (N_6444,N_4563,N_2398);
nor U6445 (N_6445,N_3082,N_3287);
nand U6446 (N_6446,N_1633,N_2373);
and U6447 (N_6447,N_959,N_4971);
xnor U6448 (N_6448,N_792,N_4513);
nand U6449 (N_6449,N_1149,N_997);
nand U6450 (N_6450,N_4456,N_259);
nor U6451 (N_6451,N_4252,N_801);
or U6452 (N_6452,N_2985,N_3099);
xnor U6453 (N_6453,N_1336,N_2859);
nor U6454 (N_6454,N_3290,N_4610);
nor U6455 (N_6455,N_4156,N_734);
or U6456 (N_6456,N_590,N_347);
nand U6457 (N_6457,N_3341,N_370);
nor U6458 (N_6458,N_1669,N_4437);
or U6459 (N_6459,N_896,N_2803);
or U6460 (N_6460,N_725,N_3796);
nand U6461 (N_6461,N_2210,N_1296);
nor U6462 (N_6462,N_3765,N_1289);
and U6463 (N_6463,N_4173,N_1457);
and U6464 (N_6464,N_578,N_2445);
nor U6465 (N_6465,N_3836,N_3528);
or U6466 (N_6466,N_2114,N_1195);
nand U6467 (N_6467,N_4891,N_401);
or U6468 (N_6468,N_2821,N_1499);
xor U6469 (N_6469,N_620,N_3246);
xor U6470 (N_6470,N_2337,N_4599);
and U6471 (N_6471,N_1550,N_2728);
nor U6472 (N_6472,N_4270,N_240);
or U6473 (N_6473,N_1454,N_3396);
nand U6474 (N_6474,N_3550,N_3807);
nand U6475 (N_6475,N_672,N_2221);
nor U6476 (N_6476,N_3009,N_1854);
nor U6477 (N_6477,N_3564,N_740);
nor U6478 (N_6478,N_4600,N_263);
nor U6479 (N_6479,N_4501,N_4311);
xor U6480 (N_6480,N_2593,N_2551);
and U6481 (N_6481,N_475,N_3219);
or U6482 (N_6482,N_2458,N_220);
or U6483 (N_6483,N_3546,N_366);
or U6484 (N_6484,N_2565,N_3107);
nand U6485 (N_6485,N_4074,N_403);
nor U6486 (N_6486,N_3124,N_4097);
nand U6487 (N_6487,N_4349,N_2849);
nand U6488 (N_6488,N_2885,N_3959);
or U6489 (N_6489,N_360,N_1450);
and U6490 (N_6490,N_22,N_2365);
nand U6491 (N_6491,N_795,N_1423);
or U6492 (N_6492,N_3445,N_383);
xor U6493 (N_6493,N_777,N_3618);
nor U6494 (N_6494,N_3557,N_1721);
nand U6495 (N_6495,N_1037,N_4931);
or U6496 (N_6496,N_4458,N_2450);
nand U6497 (N_6497,N_2388,N_2685);
and U6498 (N_6498,N_17,N_2055);
and U6499 (N_6499,N_4889,N_231);
xnor U6500 (N_6500,N_1645,N_1294);
nor U6501 (N_6501,N_2864,N_4539);
nand U6502 (N_6502,N_4330,N_4102);
nor U6503 (N_6503,N_1549,N_4107);
or U6504 (N_6504,N_1022,N_3145);
nand U6505 (N_6505,N_2657,N_3394);
or U6506 (N_6506,N_4348,N_63);
and U6507 (N_6507,N_3322,N_1733);
and U6508 (N_6508,N_3181,N_434);
and U6509 (N_6509,N_3530,N_4538);
xor U6510 (N_6510,N_4120,N_4932);
nand U6511 (N_6511,N_16,N_4656);
or U6512 (N_6512,N_2702,N_2908);
xor U6513 (N_6513,N_4010,N_1283);
and U6514 (N_6514,N_1363,N_2119);
nand U6515 (N_6515,N_3104,N_253);
nor U6516 (N_6516,N_1171,N_878);
and U6517 (N_6517,N_2224,N_2648);
nand U6518 (N_6518,N_323,N_2421);
nand U6519 (N_6519,N_1455,N_2416);
xnor U6520 (N_6520,N_1252,N_3795);
nand U6521 (N_6521,N_305,N_4628);
nand U6522 (N_6522,N_4972,N_3956);
nand U6523 (N_6523,N_1157,N_522);
and U6524 (N_6524,N_4587,N_3465);
or U6525 (N_6525,N_4947,N_1091);
nor U6526 (N_6526,N_1207,N_2903);
xnor U6527 (N_6527,N_77,N_4718);
nor U6528 (N_6528,N_4588,N_435);
nor U6529 (N_6529,N_1649,N_2798);
and U6530 (N_6530,N_2681,N_2146);
xnor U6531 (N_6531,N_2226,N_189);
nand U6532 (N_6532,N_3851,N_4059);
nand U6533 (N_6533,N_3981,N_1572);
and U6534 (N_6534,N_591,N_4789);
or U6535 (N_6535,N_4387,N_4025);
or U6536 (N_6536,N_507,N_2405);
nand U6537 (N_6537,N_4757,N_4551);
nand U6538 (N_6538,N_1051,N_2976);
nor U6539 (N_6539,N_2364,N_4344);
and U6540 (N_6540,N_1300,N_1485);
nand U6541 (N_6541,N_1174,N_3358);
nor U6542 (N_6542,N_3440,N_4363);
or U6543 (N_6543,N_270,N_4119);
or U6544 (N_6544,N_907,N_761);
or U6545 (N_6545,N_2314,N_4381);
xnor U6546 (N_6546,N_2546,N_3478);
or U6547 (N_6547,N_3118,N_3103);
and U6548 (N_6548,N_2782,N_4808);
and U6549 (N_6549,N_3995,N_2535);
xnor U6550 (N_6550,N_2902,N_3887);
nor U6551 (N_6551,N_384,N_2217);
nor U6552 (N_6552,N_2652,N_623);
nand U6553 (N_6553,N_4740,N_718);
and U6554 (N_6554,N_3668,N_4416);
nand U6555 (N_6555,N_4514,N_3313);
xnor U6556 (N_6556,N_3328,N_124);
nand U6557 (N_6557,N_4616,N_3677);
and U6558 (N_6558,N_1047,N_1473);
or U6559 (N_6559,N_3523,N_3036);
nor U6560 (N_6560,N_2360,N_3248);
nor U6561 (N_6561,N_4658,N_998);
or U6562 (N_6562,N_669,N_1507);
nor U6563 (N_6563,N_1873,N_1700);
and U6564 (N_6564,N_4584,N_4125);
xor U6565 (N_6565,N_4326,N_3864);
and U6566 (N_6566,N_4114,N_4132);
or U6567 (N_6567,N_567,N_1616);
nand U6568 (N_6568,N_3908,N_3500);
xor U6569 (N_6569,N_4370,N_2377);
and U6570 (N_6570,N_3563,N_1352);
nor U6571 (N_6571,N_1782,N_3469);
or U6572 (N_6572,N_2871,N_410);
nand U6573 (N_6573,N_3644,N_3884);
nand U6574 (N_6574,N_937,N_1162);
and U6575 (N_6575,N_2827,N_3575);
nand U6576 (N_6576,N_3013,N_325);
or U6577 (N_6577,N_842,N_342);
nand U6578 (N_6578,N_153,N_566);
or U6579 (N_6579,N_4895,N_3687);
nor U6580 (N_6580,N_2947,N_3903);
xnor U6581 (N_6581,N_3247,N_2201);
and U6582 (N_6582,N_2662,N_2077);
or U6583 (N_6583,N_2371,N_1319);
nand U6584 (N_6584,N_1515,N_1913);
or U6585 (N_6585,N_1554,N_2913);
nor U6586 (N_6586,N_3046,N_868);
nand U6587 (N_6587,N_427,N_4169);
and U6588 (N_6588,N_3768,N_4949);
nand U6589 (N_6589,N_3230,N_1920);
nand U6590 (N_6590,N_3598,N_1663);
nor U6591 (N_6591,N_1320,N_601);
nor U6592 (N_6592,N_3583,N_3143);
nor U6593 (N_6593,N_2015,N_1430);
and U6594 (N_6594,N_913,N_4845);
and U6595 (N_6595,N_463,N_1544);
or U6596 (N_6596,N_4329,N_1260);
xnor U6597 (N_6597,N_628,N_3895);
nor U6598 (N_6598,N_2384,N_815);
or U6599 (N_6599,N_4357,N_1997);
or U6600 (N_6600,N_864,N_1054);
nand U6601 (N_6601,N_1152,N_867);
nand U6602 (N_6602,N_3533,N_3163);
nand U6603 (N_6603,N_2684,N_4428);
or U6604 (N_6604,N_4359,N_3835);
or U6605 (N_6605,N_2592,N_681);
or U6606 (N_6606,N_990,N_2008);
and U6607 (N_6607,N_3295,N_4076);
nor U6608 (N_6608,N_4028,N_1830);
and U6609 (N_6609,N_3920,N_1608);
nand U6610 (N_6610,N_4572,N_4819);
or U6611 (N_6611,N_3237,N_1489);
xnor U6612 (N_6612,N_3905,N_3462);
or U6613 (N_6613,N_586,N_49);
or U6614 (N_6614,N_3024,N_4267);
and U6615 (N_6615,N_4676,N_2032);
nand U6616 (N_6616,N_3662,N_1980);
or U6617 (N_6617,N_474,N_3196);
nand U6618 (N_6618,N_201,N_13);
nand U6619 (N_6619,N_100,N_1110);
or U6620 (N_6620,N_3399,N_78);
and U6621 (N_6621,N_2841,N_68);
or U6622 (N_6622,N_2899,N_4467);
nand U6623 (N_6623,N_4203,N_544);
nand U6624 (N_6624,N_2341,N_1908);
or U6625 (N_6625,N_2703,N_4247);
nor U6626 (N_6626,N_687,N_254);
or U6627 (N_6627,N_2024,N_854);
nand U6628 (N_6628,N_123,N_610);
or U6629 (N_6629,N_1840,N_4242);
or U6630 (N_6630,N_4108,N_1970);
nand U6631 (N_6631,N_169,N_2665);
or U6632 (N_6632,N_495,N_336);
and U6633 (N_6633,N_3661,N_602);
or U6634 (N_6634,N_4631,N_4116);
or U6635 (N_6635,N_353,N_4937);
nand U6636 (N_6636,N_3022,N_4596);
and U6637 (N_6637,N_4697,N_2502);
or U6638 (N_6638,N_39,N_4350);
nor U6639 (N_6639,N_2305,N_505);
and U6640 (N_6640,N_2566,N_2001);
nor U6641 (N_6641,N_1474,N_2521);
nand U6642 (N_6642,N_848,N_2914);
nand U6643 (N_6643,N_4017,N_3588);
and U6644 (N_6644,N_1121,N_2937);
nor U6645 (N_6645,N_110,N_557);
nand U6646 (N_6646,N_4461,N_977);
nor U6647 (N_6647,N_1034,N_1744);
nor U6648 (N_6648,N_2962,N_2227);
nand U6649 (N_6649,N_1741,N_3206);
nand U6650 (N_6650,N_817,N_408);
xnor U6651 (N_6651,N_493,N_3663);
or U6652 (N_6652,N_406,N_653);
or U6653 (N_6653,N_2787,N_4477);
and U6654 (N_6654,N_1527,N_327);
xor U6655 (N_6655,N_89,N_271);
or U6656 (N_6656,N_641,N_4111);
nor U6657 (N_6657,N_4955,N_3097);
nor U6658 (N_6658,N_126,N_4936);
nor U6659 (N_6659,N_707,N_2007);
nand U6660 (N_6660,N_1823,N_3787);
nand U6661 (N_6661,N_3498,N_2356);
nor U6662 (N_6662,N_2708,N_4216);
and U6663 (N_6663,N_1947,N_2915);
nand U6664 (N_6664,N_4199,N_1516);
nor U6665 (N_6665,N_1140,N_1093);
nor U6666 (N_6666,N_3302,N_3067);
xor U6667 (N_6667,N_4301,N_3579);
or U6668 (N_6668,N_3809,N_4669);
or U6669 (N_6669,N_2148,N_1035);
xor U6670 (N_6670,N_3571,N_1929);
or U6671 (N_6671,N_186,N_4129);
and U6672 (N_6672,N_3320,N_2466);
or U6673 (N_6673,N_1671,N_2833);
and U6674 (N_6674,N_4509,N_513);
xnor U6675 (N_6675,N_4337,N_4078);
xnor U6676 (N_6676,N_1261,N_2554);
xor U6677 (N_6677,N_598,N_453);
nand U6678 (N_6678,N_83,N_2526);
nand U6679 (N_6679,N_4934,N_3801);
nor U6680 (N_6680,N_4752,N_1187);
and U6681 (N_6681,N_3140,N_2329);
nor U6682 (N_6682,N_3517,N_2719);
and U6683 (N_6683,N_1941,N_2503);
and U6684 (N_6684,N_1760,N_2924);
or U6685 (N_6685,N_4805,N_4174);
xnor U6686 (N_6686,N_4310,N_589);
or U6687 (N_6687,N_4306,N_3947);
and U6688 (N_6688,N_3160,N_3612);
xnor U6689 (N_6689,N_86,N_1097);
and U6690 (N_6690,N_4154,N_273);
nor U6691 (N_6691,N_1639,N_3490);
or U6692 (N_6692,N_1065,N_1442);
and U6693 (N_6693,N_3954,N_1165);
nand U6694 (N_6694,N_1118,N_328);
xor U6695 (N_6695,N_1912,N_646);
nand U6696 (N_6696,N_2404,N_862);
and U6697 (N_6697,N_1021,N_2730);
xnor U6698 (N_6698,N_4126,N_4712);
nand U6699 (N_6699,N_4241,N_2590);
nand U6700 (N_6700,N_3824,N_4728);
xnor U6701 (N_6701,N_4438,N_4629);
and U6702 (N_6702,N_1242,N_10);
and U6703 (N_6703,N_3332,N_3873);
nand U6704 (N_6704,N_2400,N_2598);
nor U6705 (N_6705,N_1963,N_3542);
nand U6706 (N_6706,N_445,N_866);
nor U6707 (N_6707,N_4713,N_3076);
or U6708 (N_6708,N_1654,N_774);
or U6709 (N_6709,N_4729,N_1668);
and U6710 (N_6710,N_3990,N_2744);
xnor U6711 (N_6711,N_221,N_74);
or U6712 (N_6712,N_173,N_1805);
nor U6713 (N_6713,N_534,N_2395);
nor U6714 (N_6714,N_4219,N_3562);
xor U6715 (N_6715,N_3620,N_3132);
and U6716 (N_6716,N_3117,N_1200);
nor U6717 (N_6717,N_3418,N_4518);
nor U6718 (N_6718,N_3986,N_2642);
and U6719 (N_6719,N_3063,N_1405);
nand U6720 (N_6720,N_3265,N_1867);
nand U6721 (N_6721,N_4873,N_315);
nand U6722 (N_6722,N_452,N_2006);
or U6723 (N_6723,N_2607,N_4801);
or U6724 (N_6724,N_2870,N_1501);
nor U6725 (N_6725,N_4260,N_4367);
or U6726 (N_6726,N_3263,N_1470);
and U6727 (N_6727,N_64,N_103);
xor U6728 (N_6728,N_3035,N_326);
nand U6729 (N_6729,N_2122,N_3735);
nor U6730 (N_6730,N_1103,N_183);
or U6731 (N_6731,N_1811,N_3184);
and U6732 (N_6732,N_4439,N_1480);
or U6733 (N_6733,N_709,N_2402);
or U6734 (N_6734,N_498,N_2411);
or U6735 (N_6735,N_703,N_239);
xnor U6736 (N_6736,N_161,N_1614);
nand U6737 (N_6737,N_4693,N_1108);
nor U6738 (N_6738,N_3179,N_4077);
and U6739 (N_6739,N_4547,N_4765);
and U6740 (N_6740,N_2245,N_3284);
nand U6741 (N_6741,N_3822,N_3255);
or U6742 (N_6742,N_983,N_215);
or U6743 (N_6743,N_1425,N_2451);
nor U6744 (N_6744,N_4151,N_1488);
nor U6745 (N_6745,N_272,N_2672);
nor U6746 (N_6746,N_2522,N_3623);
or U6747 (N_6747,N_1404,N_616);
nand U6748 (N_6748,N_1657,N_3624);
and U6749 (N_6749,N_1111,N_164);
or U6750 (N_6750,N_3670,N_809);
nand U6751 (N_6751,N_3998,N_4646);
xnor U6752 (N_6752,N_3087,N_916);
nor U6753 (N_6753,N_3435,N_2313);
xnor U6754 (N_6754,N_3402,N_644);
nand U6755 (N_6755,N_1769,N_1598);
nor U6756 (N_6756,N_1100,N_2932);
nor U6757 (N_6757,N_3395,N_2236);
or U6758 (N_6758,N_184,N_4528);
nor U6759 (N_6759,N_1880,N_627);
or U6760 (N_6760,N_1539,N_3673);
or U6761 (N_6761,N_1155,N_2563);
nor U6762 (N_6762,N_4709,N_3239);
nor U6763 (N_6763,N_2667,N_629);
nor U6764 (N_6764,N_4767,N_464);
nand U6765 (N_6765,N_419,N_2113);
xnor U6766 (N_6766,N_2040,N_3473);
or U6767 (N_6767,N_2699,N_3548);
nand U6768 (N_6768,N_1583,N_1849);
nand U6769 (N_6769,N_1060,N_2975);
nand U6770 (N_6770,N_1773,N_546);
or U6771 (N_6771,N_724,N_3306);
xnor U6772 (N_6772,N_1768,N_899);
xor U6773 (N_6773,N_2463,N_1285);
or U6774 (N_6774,N_974,N_592);
and U6775 (N_6775,N_1215,N_4315);
xor U6776 (N_6776,N_1017,N_4279);
or U6777 (N_6777,N_3,N_2281);
and U6778 (N_6778,N_3922,N_4768);
or U6779 (N_6779,N_1059,N_2664);
or U6780 (N_6780,N_222,N_4412);
xor U6781 (N_6781,N_4385,N_4168);
nor U6782 (N_6782,N_4804,N_3018);
and U6783 (N_6783,N_594,N_3937);
and U6784 (N_6784,N_3479,N_1943);
and U6785 (N_6785,N_3797,N_1380);
and U6786 (N_6786,N_3431,N_861);
nor U6787 (N_6787,N_4372,N_149);
or U6788 (N_6788,N_1581,N_3718);
nor U6789 (N_6789,N_4336,N_3416);
and U6790 (N_6790,N_1209,N_4491);
and U6791 (N_6791,N_2552,N_1893);
and U6792 (N_6792,N_1794,N_4564);
xnor U6793 (N_6793,N_4238,N_2274);
or U6794 (N_6794,N_1705,N_698);
or U6795 (N_6795,N_1731,N_1217);
and U6796 (N_6796,N_1531,N_2325);
and U6797 (N_6797,N_4702,N_3614);
or U6798 (N_6798,N_1592,N_3300);
and U6799 (N_6799,N_4545,N_4159);
nand U6800 (N_6800,N_4737,N_1950);
or U6801 (N_6801,N_378,N_637);
nand U6802 (N_6802,N_1089,N_2625);
and U6803 (N_6803,N_705,N_1776);
and U6804 (N_6804,N_234,N_219);
or U6805 (N_6805,N_2797,N_1397);
or U6806 (N_6806,N_1620,N_4604);
or U6807 (N_6807,N_4816,N_3146);
or U6808 (N_6808,N_1612,N_131);
nand U6809 (N_6809,N_1432,N_4489);
and U6810 (N_6810,N_3559,N_4493);
and U6811 (N_6811,N_3850,N_3235);
nor U6812 (N_6812,N_2900,N_3859);
or U6813 (N_6813,N_3885,N_654);
nand U6814 (N_6814,N_4052,N_4560);
nand U6815 (N_6815,N_888,N_4026);
and U6816 (N_6816,N_4465,N_747);
nand U6817 (N_6817,N_4195,N_716);
or U6818 (N_6818,N_2192,N_1508);
or U6819 (N_6819,N_3267,N_3881);
nor U6820 (N_6820,N_2511,N_3403);
nand U6821 (N_6821,N_1722,N_3727);
or U6822 (N_6822,N_3293,N_4692);
and U6823 (N_6823,N_3433,N_3805);
or U6824 (N_6824,N_1984,N_2901);
nor U6825 (N_6825,N_25,N_1354);
and U6826 (N_6826,N_3415,N_2126);
or U6827 (N_6827,N_3323,N_762);
or U6828 (N_6828,N_4209,N_4444);
or U6829 (N_6829,N_1409,N_885);
xor U6830 (N_6830,N_3819,N_97);
or U6831 (N_6831,N_1890,N_923);
and U6832 (N_6832,N_504,N_1892);
xor U6833 (N_6833,N_4309,N_2835);
or U6834 (N_6834,N_4743,N_3142);
xnor U6835 (N_6835,N_1730,N_2157);
and U6836 (N_6836,N_2335,N_1437);
and U6837 (N_6837,N_3085,N_4488);
or U6838 (N_6838,N_1965,N_2982);
nand U6839 (N_6839,N_2764,N_1809);
xor U6840 (N_6840,N_428,N_1193);
or U6841 (N_6841,N_4101,N_3821);
nand U6842 (N_6842,N_511,N_1719);
and U6843 (N_6843,N_4624,N_787);
nor U6844 (N_6844,N_1600,N_3171);
nor U6845 (N_6845,N_1962,N_4534);
xnor U6846 (N_6846,N_441,N_3222);
or U6847 (N_6847,N_3484,N_4916);
and U6848 (N_6848,N_2823,N_2473);
and U6849 (N_6849,N_4148,N_4760);
and U6850 (N_6850,N_2125,N_1896);
or U6851 (N_6851,N_2141,N_1406);
and U6852 (N_6852,N_3080,N_3398);
xor U6853 (N_6853,N_329,N_1538);
nand U6854 (N_6854,N_2410,N_23);
xnor U6855 (N_6855,N_269,N_4540);
nor U6856 (N_6856,N_2232,N_4355);
or U6857 (N_6857,N_2547,N_3933);
nand U6858 (N_6858,N_73,N_4362);
nand U6859 (N_6859,N_4505,N_2447);
nand U6860 (N_6860,N_2940,N_3467);
xnor U6861 (N_6861,N_4793,N_2925);
nand U6862 (N_6862,N_4008,N_1615);
nor U6863 (N_6863,N_845,N_2425);
nor U6864 (N_6864,N_2218,N_4302);
and U6865 (N_6865,N_4222,N_1349);
nand U6866 (N_6866,N_3039,N_3975);
xor U6867 (N_6867,N_4826,N_1365);
and U6868 (N_6868,N_1993,N_1419);
nand U6869 (N_6869,N_3147,N_3397);
or U6870 (N_6870,N_1517,N_1378);
xnor U6871 (N_6871,N_2163,N_4044);
nand U6872 (N_6872,N_4007,N_860);
nand U6873 (N_6873,N_2644,N_2854);
nor U6874 (N_6874,N_2110,N_71);
xnor U6875 (N_6875,N_3664,N_2283);
nor U6876 (N_6876,N_1186,N_3471);
and U6877 (N_6877,N_407,N_3769);
or U6878 (N_6878,N_1866,N_614);
nor U6879 (N_6879,N_2342,N_4531);
nor U6880 (N_6880,N_3014,N_1144);
and U6881 (N_6881,N_4075,N_1158);
or U6882 (N_6882,N_4099,N_3008);
and U6883 (N_6883,N_1898,N_2366);
or U6884 (N_6884,N_3325,N_1626);
nand U6885 (N_6885,N_1459,N_449);
nor U6886 (N_6886,N_4735,N_4414);
and U6887 (N_6887,N_2946,N_3078);
nor U6888 (N_6888,N_2327,N_1080);
or U6889 (N_6889,N_802,N_2500);
xnor U6890 (N_6890,N_1832,N_4146);
and U6891 (N_6891,N_4984,N_1015);
nand U6892 (N_6892,N_639,N_4164);
nand U6893 (N_6893,N_3413,N_2737);
or U6894 (N_6894,N_2287,N_2846);
xor U6895 (N_6895,N_924,N_711);
nor U6896 (N_6896,N_2993,N_2168);
and U6897 (N_6897,N_2093,N_2277);
nand U6898 (N_6898,N_2602,N_1415);
or U6899 (N_6899,N_2640,N_4673);
nand U6900 (N_6900,N_1417,N_3551);
nor U6901 (N_6901,N_4282,N_114);
or U6902 (N_6902,N_996,N_195);
and U6903 (N_6903,N_3766,N_3482);
and U6904 (N_6904,N_1385,N_2553);
or U6905 (N_6905,N_3135,N_246);
and U6906 (N_6906,N_1379,N_3414);
nand U6907 (N_6907,N_4763,N_2796);
xnor U6908 (N_6908,N_4809,N_3569);
nand U6909 (N_6909,N_2043,N_2753);
and U6910 (N_6910,N_1704,N_4457);
and U6911 (N_6911,N_1303,N_2585);
xor U6912 (N_6912,N_4037,N_4064);
nand U6913 (N_6913,N_4680,N_1495);
nor U6914 (N_6914,N_1129,N_1262);
and U6915 (N_6915,N_2759,N_3499);
nor U6916 (N_6916,N_4901,N_3481);
xnor U6917 (N_6917,N_156,N_2709);
xor U6918 (N_6918,N_2650,N_1456);
or U6919 (N_6919,N_229,N_4846);
nand U6920 (N_6920,N_1077,N_2848);
and U6921 (N_6921,N_3651,N_4831);
nand U6922 (N_6922,N_3685,N_1075);
or U6923 (N_6923,N_1190,N_3278);
nand U6924 (N_6924,N_4655,N_2131);
nand U6925 (N_6925,N_3138,N_1855);
nor U6926 (N_6926,N_2291,N_2504);
nand U6927 (N_6927,N_3041,N_2353);
nand U6928 (N_6928,N_1804,N_2634);
or U6929 (N_6929,N_970,N_2182);
and U6930 (N_6930,N_3083,N_3049);
nand U6931 (N_6931,N_946,N_738);
nand U6932 (N_6932,N_4771,N_1424);
nor U6933 (N_6933,N_4525,N_982);
or U6934 (N_6934,N_4000,N_1235);
nor U6935 (N_6935,N_3757,N_784);
nand U6936 (N_6936,N_1273,N_1220);
nor U6937 (N_6937,N_1197,N_281);
or U6938 (N_6938,N_2599,N_3053);
nand U6939 (N_6939,N_3244,N_3188);
or U6940 (N_6940,N_901,N_363);
or U6941 (N_6941,N_2316,N_4471);
and U6942 (N_6942,N_4733,N_4994);
or U6943 (N_6943,N_4274,N_3828);
and U6944 (N_6944,N_3591,N_485);
nand U6945 (N_6945,N_2150,N_4157);
or U6946 (N_6946,N_296,N_2875);
and U6947 (N_6947,N_2677,N_3436);
nand U6948 (N_6948,N_4854,N_2238);
nor U6949 (N_6949,N_1569,N_4497);
nand U6950 (N_6950,N_840,N_3708);
or U6951 (N_6951,N_2887,N_2048);
nor U6952 (N_6952,N_440,N_2873);
nand U6953 (N_6953,N_1701,N_4239);
or U6954 (N_6954,N_3026,N_2520);
or U6955 (N_6955,N_3310,N_1610);
nand U6956 (N_6956,N_4500,N_1757);
nand U6957 (N_6957,N_3665,N_877);
and U6958 (N_6958,N_2581,N_1066);
and U6959 (N_6959,N_1311,N_3177);
or U6960 (N_6960,N_3909,N_4091);
xnor U6961 (N_6961,N_4449,N_3914);
and U6962 (N_6962,N_2228,N_1618);
xnor U6963 (N_6963,N_2627,N_3324);
nor U6964 (N_6964,N_1894,N_4502);
nor U6965 (N_6965,N_47,N_4565);
or U6966 (N_6966,N_4137,N_1061);
nor U6967 (N_6967,N_3298,N_2675);
and U6968 (N_6968,N_3294,N_2653);
or U6969 (N_6969,N_3274,N_2455);
nand U6970 (N_6970,N_4668,N_3472);
and U6971 (N_6971,N_3092,N_4402);
nand U6972 (N_6972,N_3590,N_389);
nor U6973 (N_6973,N_773,N_2022);
and U6974 (N_6974,N_1502,N_2692);
and U6975 (N_6975,N_2619,N_2838);
nand U6976 (N_6976,N_2403,N_2778);
and U6977 (N_6977,N_1347,N_4674);
xor U6978 (N_6978,N_1665,N_1478);
nor U6979 (N_6979,N_1526,N_1528);
nor U6980 (N_6980,N_1697,N_3090);
nand U6981 (N_6981,N_2624,N_265);
xor U6982 (N_6982,N_1518,N_2659);
or U6983 (N_6983,N_3225,N_1842);
and U6984 (N_6984,N_4903,N_1761);
or U6985 (N_6985,N_3619,N_3678);
nand U6986 (N_6986,N_4021,N_2513);
nor U6987 (N_6987,N_2789,N_1658);
xor U6988 (N_6988,N_1653,N_2683);
and U6989 (N_6989,N_159,N_753);
and U6990 (N_6990,N_4033,N_4377);
xor U6991 (N_6991,N_1799,N_3798);
xor U6992 (N_6992,N_4445,N_4945);
and U6993 (N_6993,N_4788,N_3487);
and U6994 (N_6994,N_3976,N_4675);
or U6995 (N_6995,N_1448,N_1632);
xnor U6996 (N_6996,N_4957,N_3584);
nand U6997 (N_6997,N_2694,N_4677);
nand U6998 (N_6998,N_832,N_1016);
nand U6999 (N_6999,N_4830,N_1329);
nand U7000 (N_7000,N_2285,N_3204);
nor U7001 (N_7001,N_2026,N_4248);
or U7002 (N_7002,N_1938,N_2637);
and U7003 (N_7003,N_3803,N_2645);
nor U7004 (N_7004,N_3544,N_3349);
and U7005 (N_7005,N_1338,N_1373);
nor U7006 (N_7006,N_837,N_2666);
or U7007 (N_7007,N_902,N_2028);
and U7008 (N_7008,N_4392,N_486);
and U7009 (N_7009,N_4482,N_3153);
xnor U7010 (N_7010,N_1440,N_1714);
nor U7011 (N_7011,N_1134,N_1625);
xnor U7012 (N_7012,N_2158,N_2085);
nand U7013 (N_7013,N_3759,N_140);
nor U7014 (N_7014,N_415,N_3126);
or U7015 (N_7015,N_2567,N_4925);
nand U7016 (N_7016,N_2674,N_4758);
nor U7017 (N_7017,N_1797,N_4088);
and U7018 (N_7018,N_1692,N_409);
xor U7019 (N_7019,N_1316,N_2560);
nor U7020 (N_7020,N_893,N_518);
and U7021 (N_7021,N_1874,N_1906);
and U7022 (N_7022,N_929,N_565);
and U7023 (N_7023,N_3058,N_2019);
nand U7024 (N_7024,N_4811,N_4251);
and U7025 (N_7025,N_1079,N_2334);
and U7026 (N_7026,N_2086,N_4206);
nor U7027 (N_7027,N_1000,N_4331);
nand U7028 (N_7028,N_1033,N_202);
nand U7029 (N_7029,N_1224,N_4630);
nor U7030 (N_7030,N_2263,N_4190);
or U7031 (N_7031,N_920,N_2288);
xnor U7032 (N_7032,N_1327,N_3910);
nor U7033 (N_7033,N_457,N_4615);
nor U7034 (N_7034,N_969,N_4902);
and U7035 (N_7035,N_4578,N_1101);
or U7036 (N_7036,N_1956,N_500);
nor U7037 (N_7037,N_2214,N_750);
or U7038 (N_7038,N_2714,N_3962);
nor U7039 (N_7039,N_4660,N_3392);
and U7040 (N_7040,N_2176,N_2142);
nor U7041 (N_7041,N_2747,N_1901);
nor U7042 (N_7042,N_4720,N_4559);
nand U7043 (N_7043,N_212,N_2202);
nor U7044 (N_7044,N_701,N_1691);
nand U7045 (N_7045,N_2532,N_4868);
and U7046 (N_7046,N_4446,N_3307);
nor U7047 (N_7047,N_294,N_284);
and U7048 (N_7048,N_979,N_2501);
nor U7049 (N_7049,N_3891,N_311);
nor U7050 (N_7050,N_1208,N_2111);
nand U7051 (N_7051,N_3421,N_541);
nor U7052 (N_7052,N_3565,N_879);
nor U7053 (N_7053,N_2729,N_1828);
xnor U7054 (N_7054,N_680,N_2087);
nor U7055 (N_7055,N_4979,N_1493);
or U7056 (N_7056,N_4232,N_1324);
nand U7057 (N_7057,N_3215,N_443);
nor U7058 (N_7058,N_224,N_2225);
and U7059 (N_7059,N_1870,N_4474);
or U7060 (N_7060,N_3441,N_2200);
xnor U7061 (N_7061,N_317,N_3723);
nor U7062 (N_7062,N_4070,N_1709);
or U7063 (N_7063,N_158,N_3566);
nor U7064 (N_7064,N_483,N_2539);
or U7065 (N_7065,N_1085,N_3697);
nor U7066 (N_7066,N_967,N_1673);
nand U7067 (N_7067,N_2584,N_4586);
and U7068 (N_7068,N_3289,N_537);
nor U7069 (N_7069,N_3113,N_4205);
and U7070 (N_7070,N_1068,N_1815);
nor U7071 (N_7071,N_3994,N_3744);
or U7072 (N_7072,N_4784,N_4837);
nor U7073 (N_7073,N_3955,N_2606);
xor U7074 (N_7074,N_2091,N_2556);
and U7075 (N_7075,N_2211,N_735);
or U7076 (N_7076,N_4229,N_4794);
nor U7077 (N_7077,N_3957,N_1790);
nand U7078 (N_7078,N_1233,N_432);
xor U7079 (N_7079,N_1648,N_1514);
nor U7080 (N_7080,N_2831,N_2646);
nor U7081 (N_7081,N_3468,N_1936);
nand U7082 (N_7082,N_1903,N_2029);
nor U7083 (N_7083,N_1340,N_121);
xor U7084 (N_7084,N_585,N_1677);
or U7085 (N_7085,N_4431,N_3410);
and U7086 (N_7086,N_4223,N_2344);
and U7087 (N_7087,N_4755,N_4432);
nand U7088 (N_7088,N_3934,N_3100);
and U7089 (N_7089,N_4665,N_1234);
or U7090 (N_7090,N_1323,N_1696);
nand U7091 (N_7091,N_2770,N_3081);
and U7092 (N_7092,N_1523,N_4698);
nor U7093 (N_7093,N_3430,N_1590);
nand U7094 (N_7094,N_1852,N_1775);
and U7095 (N_7095,N_2861,N_3494);
nand U7096 (N_7096,N_1449,N_3401);
nor U7097 (N_7097,N_755,N_1355);
nand U7098 (N_7098,N_150,N_1026);
or U7099 (N_7099,N_2191,N_3485);
xor U7100 (N_7100,N_1314,N_2345);
nor U7101 (N_7101,N_1183,N_1131);
and U7102 (N_7102,N_3802,N_2222);
nand U7103 (N_7103,N_980,N_3189);
nand U7104 (N_7104,N_429,N_2369);
or U7105 (N_7105,N_2611,N_4814);
nand U7106 (N_7106,N_4792,N_4882);
and U7107 (N_7107,N_2185,N_821);
and U7108 (N_7108,N_3977,N_4215);
and U7109 (N_7109,N_2695,N_3345);
xor U7110 (N_7110,N_4155,N_379);
and U7111 (N_7111,N_2746,N_4245);
nand U7112 (N_7112,N_4722,N_3899);
nand U7113 (N_7113,N_180,N_194);
nand U7114 (N_7114,N_1204,N_1227);
nor U7115 (N_7115,N_1846,N_4823);
or U7116 (N_7116,N_839,N_2622);
nand U7117 (N_7117,N_2814,N_3056);
nand U7118 (N_7118,N_2658,N_3505);
nand U7119 (N_7119,N_4813,N_3741);
nor U7120 (N_7120,N_1911,N_696);
and U7121 (N_7121,N_3915,N_2528);
and U7122 (N_7122,N_985,N_939);
nand U7123 (N_7123,N_4498,N_3259);
and U7124 (N_7124,N_2076,N_1780);
nand U7125 (N_7125,N_3269,N_3251);
nand U7126 (N_7126,N_2332,N_4047);
nor U7127 (N_7127,N_3405,N_2810);
and U7128 (N_7128,N_2668,N_3637);
and U7129 (N_7129,N_2322,N_122);
or U7130 (N_7130,N_3928,N_1638);
or U7131 (N_7131,N_3603,N_547);
xnor U7132 (N_7132,N_3675,N_1779);
or U7133 (N_7133,N_2912,N_2433);
nand U7134 (N_7134,N_385,N_3305);
xnor U7135 (N_7135,N_2349,N_4550);
nand U7136 (N_7136,N_2978,N_2014);
nor U7137 (N_7137,N_1547,N_4933);
nor U7138 (N_7138,N_4861,N_3045);
nand U7139 (N_7139,N_3846,N_2472);
nand U7140 (N_7140,N_2939,N_4732);
xnor U7141 (N_7141,N_3089,N_1778);
nor U7142 (N_7142,N_1602,N_4736);
nor U7143 (N_7143,N_276,N_1571);
and U7144 (N_7144,N_2812,N_4838);
nor U7145 (N_7145,N_2815,N_3136);
nand U7146 (N_7146,N_3119,N_3268);
nor U7147 (N_7147,N_2194,N_3988);
nor U7148 (N_7148,N_3690,N_4664);
or U7149 (N_7149,N_3774,N_3057);
xnor U7150 (N_7150,N_2632,N_3626);
and U7151 (N_7151,N_2461,N_2495);
nor U7152 (N_7152,N_355,N_4928);
nor U7153 (N_7153,N_285,N_1882);
nand U7154 (N_7154,N_3372,N_776);
and U7155 (N_7155,N_437,N_4739);
nand U7156 (N_7156,N_3501,N_2820);
nor U7157 (N_7157,N_4871,N_909);
xor U7158 (N_7158,N_2452,N_1931);
or U7159 (N_7159,N_4791,N_2734);
or U7160 (N_7160,N_2396,N_373);
xor U7161 (N_7161,N_3736,N_1748);
nand U7162 (N_7162,N_4095,N_1655);
or U7163 (N_7163,N_223,N_2972);
nor U7164 (N_7164,N_3958,N_3360);
and U7165 (N_7165,N_4415,N_649);
xor U7166 (N_7166,N_1353,N_303);
nand U7167 (N_7167,N_1791,N_532);
xnor U7168 (N_7168,N_4970,N_3514);
nor U7169 (N_7169,N_2178,N_3700);
and U7170 (N_7170,N_4824,N_835);
and U7171 (N_7171,N_2643,N_2507);
nor U7172 (N_7172,N_2564,N_682);
nor U7173 (N_7173,N_66,N_597);
nand U7174 (N_7174,N_3042,N_4503);
and U7175 (N_7175,N_238,N_4879);
or U7176 (N_7176,N_3288,N_3475);
and U7177 (N_7177,N_2533,N_2443);
nor U7178 (N_7178,N_111,N_1433);
or U7179 (N_7179,N_645,N_2188);
and U7180 (N_7180,N_1509,N_2678);
and U7181 (N_7181,N_3314,N_3679);
nand U7182 (N_7182,N_3375,N_1006);
xnor U7183 (N_7183,N_365,N_1637);
xor U7184 (N_7184,N_4877,N_3231);
and U7185 (N_7185,N_4962,N_37);
or U7186 (N_7186,N_2270,N_1063);
or U7187 (N_7187,N_4989,N_2767);
nor U7188 (N_7188,N_2679,N_3291);
or U7189 (N_7189,N_3716,N_3047);
or U7190 (N_7190,N_172,N_579);
nand U7191 (N_7191,N_1563,N_664);
or U7192 (N_7192,N_4619,N_652);
nor U7193 (N_7193,N_2469,N_3804);
and U7194 (N_7194,N_1628,N_2442);
nand U7195 (N_7195,N_4866,N_2756);
nand U7196 (N_7196,N_2964,N_4603);
and U7197 (N_7197,N_858,N_1403);
nor U7198 (N_7198,N_4394,N_3931);
nor U7199 (N_7199,N_2268,N_1460);
or U7200 (N_7200,N_3613,N_791);
nand U7201 (N_7201,N_479,N_181);
nor U7202 (N_7202,N_2572,N_1359);
or U7203 (N_7203,N_2354,N_1038);
and U7204 (N_7204,N_151,N_2857);
and U7205 (N_7205,N_4228,N_2427);
nor U7206 (N_7206,N_2663,N_289);
or U7207 (N_7207,N_975,N_1955);
and U7208 (N_7208,N_516,N_798);
or U7209 (N_7209,N_1346,N_1548);
or U7210 (N_7210,N_3088,N_4496);
nand U7211 (N_7211,N_2195,N_2777);
xnor U7212 (N_7212,N_4940,N_4858);
nor U7213 (N_7213,N_4063,N_335);
nor U7214 (N_7214,N_4442,N_736);
nor U7215 (N_7215,N_4399,N_635);
and U7216 (N_7216,N_137,N_2392);
or U7217 (N_7217,N_1122,N_4959);
or U7218 (N_7218,N_3680,N_1302);
nor U7219 (N_7219,N_2174,N_1945);
and U7220 (N_7220,N_3978,N_4800);
nor U7221 (N_7221,N_2205,N_349);
nor U7222 (N_7222,N_356,N_4527);
nor U7223 (N_7223,N_4434,N_964);
xor U7224 (N_7224,N_4262,N_1276);
nor U7225 (N_7225,N_2359,N_3806);
nand U7226 (N_7226,N_141,N_119);
nor U7227 (N_7227,N_4683,N_772);
and U7228 (N_7228,N_781,N_4815);
or U7229 (N_7229,N_2017,N_1927);
or U7230 (N_7230,N_4682,N_426);
nor U7231 (N_7231,N_2731,N_3356);
and U7232 (N_7232,N_2514,N_4466);
or U7233 (N_7233,N_895,N_1494);
nand U7234 (N_7234,N_2462,N_1072);
nand U7235 (N_7235,N_1909,N_1763);
or U7236 (N_7236,N_2399,N_4356);
nor U7237 (N_7237,N_2577,N_3866);
and U7238 (N_7238,N_4690,N_2216);
and U7239 (N_7239,N_2739,N_1008);
xor U7240 (N_7240,N_174,N_3216);
and U7241 (N_7241,N_1810,N_4294);
nand U7242 (N_7242,N_3615,N_715);
or U7243 (N_7243,N_3580,N_1069);
xor U7244 (N_7244,N_3355,N_2483);
and U7245 (N_7245,N_1845,N_1228);
xnor U7246 (N_7246,N_4234,N_2830);
nand U7247 (N_7247,N_891,N_4404);
nand U7248 (N_7248,N_502,N_2165);
nand U7249 (N_7249,N_3333,N_1742);
xor U7250 (N_7250,N_1787,N_139);
or U7251 (N_7251,N_674,N_4652);
nand U7252 (N_7252,N_2428,N_4443);
nor U7253 (N_7253,N_1028,N_2805);
and U7254 (N_7254,N_1496,N_1071);
nand U7255 (N_7255,N_2151,N_1391);
or U7256 (N_7256,N_2003,N_3382);
nand U7257 (N_7257,N_4857,N_3151);
and U7258 (N_7258,N_4158,N_2145);
nand U7259 (N_7259,N_3625,N_4378);
nand U7260 (N_7260,N_1231,N_1465);
nor U7261 (N_7261,N_1444,N_1622);
nand U7262 (N_7262,N_1835,N_2788);
xor U7263 (N_7263,N_3220,N_2860);
nand U7264 (N_7264,N_4515,N_3450);
and U7265 (N_7265,N_2601,N_3574);
and U7266 (N_7266,N_1578,N_494);
nor U7267 (N_7267,N_3552,N_120);
and U7268 (N_7268,N_4974,N_4283);
nand U7269 (N_7269,N_816,N_617);
xor U7270 (N_7270,N_3352,N_3336);
nor U7271 (N_7271,N_2636,N_4554);
or U7272 (N_7272,N_3984,N_3187);
nor U7273 (N_7273,N_3763,N_3813);
nor U7274 (N_7274,N_2723,N_925);
or U7275 (N_7275,N_4011,N_3963);
nor U7276 (N_7276,N_3448,N_4623);
xnor U7277 (N_7277,N_430,N_4863);
and U7278 (N_7278,N_4905,N_1918);
nor U7279 (N_7279,N_1881,N_4323);
or U7280 (N_7280,N_258,N_1014);
nand U7281 (N_7281,N_634,N_2470);
or U7282 (N_7282,N_926,N_691);
nor U7283 (N_7283,N_4643,N_2989);
and U7284 (N_7284,N_154,N_508);
or U7285 (N_7285,N_2233,N_1555);
nor U7286 (N_7286,N_4750,N_3949);
or U7287 (N_7287,N_3657,N_395);
and U7288 (N_7288,N_2417,N_2098);
nand U7289 (N_7289,N_857,N_3420);
nor U7290 (N_7290,N_264,N_2574);
and U7291 (N_7291,N_2869,N_4731);
or U7292 (N_7292,N_1239,N_4923);
or U7293 (N_7293,N_1383,N_3989);
nor U7294 (N_7294,N_4196,N_693);
and U7295 (N_7295,N_2235,N_3474);
xor U7296 (N_7296,N_4390,N_319);
and U7297 (N_7297,N_4993,N_3125);
and U7298 (N_7298,N_2480,N_3942);
or U7299 (N_7299,N_3743,N_185);
nand U7300 (N_7300,N_3232,N_535);
or U7301 (N_7301,N_4642,N_1211);
and U7302 (N_7302,N_603,N_1178);
nor U7303 (N_7303,N_2806,N_2688);
nand U7304 (N_7304,N_3006,N_1438);
nand U7305 (N_7305,N_3578,N_4759);
nand U7306 (N_7306,N_1389,N_3093);
and U7307 (N_7307,N_2257,N_3865);
nor U7308 (N_7308,N_2608,N_4192);
and U7309 (N_7309,N_2816,N_947);
and U7310 (N_7310,N_2950,N_2882);
nand U7311 (N_7311,N_1861,N_1382);
or U7312 (N_7312,N_1541,N_3856);
or U7313 (N_7313,N_3969,N_1829);
and U7314 (N_7314,N_3869,N_3115);
nor U7315 (N_7315,N_2412,N_2807);
or U7316 (N_7316,N_3249,N_1469);
or U7317 (N_7317,N_2180,N_1342);
and U7318 (N_7318,N_359,N_4226);
and U7319 (N_7319,N_245,N_2893);
or U7320 (N_7320,N_1288,N_3814);
nor U7321 (N_7321,N_992,N_211);
nor U7322 (N_7322,N_4299,N_803);
or U7323 (N_7323,N_4797,N_2352);
nor U7324 (N_7324,N_2963,N_3556);
nor U7325 (N_7325,N_3199,N_4557);
nor U7326 (N_7326,N_4451,N_810);
nand U7327 (N_7327,N_3825,N_4187);
nor U7328 (N_7328,N_4754,N_4188);
and U7329 (N_7329,N_3511,N_1922);
or U7330 (N_7330,N_469,N_4822);
nor U7331 (N_7331,N_52,N_2516);
and U7332 (N_7332,N_833,N_3932);
or U7333 (N_7333,N_191,N_3519);
and U7334 (N_7334,N_1492,N_3317);
or U7335 (N_7335,N_1715,N_2771);
or U7336 (N_7336,N_3871,N_1537);
nor U7337 (N_7337,N_2280,N_3114);
or U7338 (N_7338,N_416,N_1836);
or U7339 (N_7339,N_986,N_3572);
nand U7340 (N_7340,N_82,N_2795);
or U7341 (N_7341,N_2638,N_35);
xor U7342 (N_7342,N_4318,N_3185);
nand U7343 (N_7343,N_4888,N_624);
and U7344 (N_7344,N_4024,N_1381);
nand U7345 (N_7345,N_1619,N_2031);
or U7346 (N_7346,N_1003,N_3025);
nor U7347 (N_7347,N_519,N_1113);
xnor U7348 (N_7348,N_2881,N_364);
and U7349 (N_7349,N_3715,N_1087);
or U7350 (N_7350,N_2799,N_1762);
or U7351 (N_7351,N_3968,N_2020);
xor U7352 (N_7352,N_1169,N_4176);
nand U7353 (N_7353,N_351,N_2047);
nand U7354 (N_7354,N_2269,N_1150);
and U7355 (N_7355,N_3286,N_622);
or U7356 (N_7356,N_4055,N_1393);
nand U7357 (N_7357,N_152,N_2895);
and U7358 (N_7358,N_4225,N_4592);
or U7359 (N_7359,N_2046,N_869);
nand U7360 (N_7360,N_3681,N_3218);
and U7361 (N_7361,N_4715,N_3704);
and U7362 (N_7362,N_4976,N_1270);
nor U7363 (N_7363,N_3701,N_2075);
nand U7364 (N_7364,N_115,N_568);
nand U7365 (N_7365,N_3329,N_2186);
xor U7366 (N_7366,N_2775,N_2726);
or U7367 (N_7367,N_2498,N_582);
nand U7368 (N_7368,N_3656,N_1717);
nand U7369 (N_7369,N_2067,N_4553);
and U7370 (N_7370,N_376,N_1500);
xor U7371 (N_7371,N_1834,N_737);
nor U7372 (N_7372,N_2271,N_168);
nor U7373 (N_7373,N_4917,N_1988);
and U7374 (N_7374,N_739,N_4661);
nor U7375 (N_7375,N_2649,N_4913);
and U7376 (N_7376,N_3369,N_3772);
nand U7377 (N_7377,N_2187,N_732);
and U7378 (N_7378,N_34,N_2460);
or U7379 (N_7379,N_4142,N_3898);
and U7380 (N_7380,N_3098,N_176);
nand U7381 (N_7381,N_1375,N_2272);
nand U7382 (N_7382,N_2207,N_2130);
or U7383 (N_7383,N_685,N_4447);
nand U7384 (N_7384,N_4950,N_2852);
or U7385 (N_7385,N_54,N_2689);
nor U7386 (N_7386,N_4653,N_2680);
or U7387 (N_7387,N_745,N_3242);
nor U7388 (N_7388,N_3829,N_531);
xnor U7389 (N_7389,N_2661,N_4401);
or U7390 (N_7390,N_2487,N_2292);
nor U7391 (N_7391,N_2260,N_3347);
xnor U7392 (N_7392,N_2118,N_2298);
and U7393 (N_7393,N_1412,N_3466);
and U7394 (N_7394,N_1141,N_1315);
nand U7395 (N_7395,N_4388,N_2045);
nor U7396 (N_7396,N_3271,N_300);
nor U7397 (N_7397,N_3785,N_995);
nor U7398 (N_7398,N_1561,N_4268);
nand U7399 (N_7399,N_3547,N_3084);
or U7400 (N_7400,N_2062,N_2671);
nand U7401 (N_7401,N_2506,N_3275);
or U7402 (N_7402,N_2056,N_2832);
xor U7403 (N_7403,N_3031,N_1271);
or U7404 (N_7404,N_1226,N_1736);
or U7405 (N_7405,N_1899,N_3368);
or U7406 (N_7406,N_1670,N_4679);
nand U7407 (N_7407,N_3896,N_4836);
xnor U7408 (N_7408,N_612,N_1330);
nor U7409 (N_7409,N_648,N_4476);
and U7410 (N_7410,N_4041,N_4625);
nand U7411 (N_7411,N_387,N_2310);
nor U7412 (N_7412,N_695,N_663);
nor U7413 (N_7413,N_642,N_446);
nor U7414 (N_7414,N_3193,N_1946);
nor U7415 (N_7415,N_757,N_2219);
nor U7416 (N_7416,N_4875,N_1989);
nand U7417 (N_7417,N_3827,N_4407);
xor U7418 (N_7418,N_884,N_562);
and U7419 (N_7419,N_948,N_1540);
nor U7420 (N_7420,N_1146,N_3642);
and U7421 (N_7421,N_1057,N_3442);
xnor U7422 (N_7422,N_3463,N_4018);
or U7423 (N_7423,N_4109,N_3607);
or U7424 (N_7424,N_2179,N_604);
or U7425 (N_7425,N_4334,N_730);
nor U7426 (N_7426,N_4833,N_729);
nor U7427 (N_7427,N_988,N_1825);
and U7428 (N_7428,N_3139,N_368);
or U7429 (N_7429,N_2935,N_402);
xnor U7430 (N_7430,N_4659,N_1680);
xor U7431 (N_7431,N_3758,N_3208);
or U7432 (N_7432,N_4689,N_3068);
nand U7433 (N_7433,N_2401,N_4621);
and U7434 (N_7434,N_2966,N_4410);
nor U7435 (N_7435,N_3786,N_3531);
nand U7436 (N_7436,N_2090,N_3738);
nand U7437 (N_7437,N_4747,N_2021);
and U7438 (N_7438,N_2919,N_2647);
or U7439 (N_7439,N_4034,N_524);
xor U7440 (N_7440,N_1800,N_274);
nor U7441 (N_7441,N_312,N_391);
xnor U7442 (N_7442,N_2951,N_4843);
nor U7443 (N_7443,N_1595,N_3857);
or U7444 (N_7444,N_4576,N_1056);
xor U7445 (N_7445,N_4543,N_2453);
nor U7446 (N_7446,N_4138,N_657);
or U7447 (N_7447,N_2751,N_1039);
or U7448 (N_7448,N_2809,N_361);
or U7449 (N_7449,N_3770,N_4853);
xor U7450 (N_7450,N_91,N_3425);
and U7451 (N_7451,N_818,N_1897);
nand U7452 (N_7452,N_3342,N_4147);
and U7453 (N_7453,N_713,N_2929);
and U7454 (N_7454,N_887,N_1143);
nand U7455 (N_7455,N_1306,N_55);
nor U7456 (N_7456,N_3719,N_2415);
nor U7457 (N_7457,N_1426,N_1745);
nor U7458 (N_7458,N_1580,N_2100);
and U7459 (N_7459,N_1328,N_2761);
and U7460 (N_7460,N_1232,N_310);
and U7461 (N_7461,N_4440,N_3912);
nand U7462 (N_7462,N_1055,N_892);
nor U7463 (N_7463,N_2582,N_3055);
or U7464 (N_7464,N_394,N_1428);
or U7465 (N_7465,N_1562,N_4887);
nor U7466 (N_7466,N_2927,N_3792);
and U7467 (N_7467,N_2102,N_481);
nand U7468 (N_7468,N_7,N_182);
nand U7469 (N_7469,N_3586,N_2786);
and U7470 (N_7470,N_2005,N_3223);
or U7471 (N_7471,N_662,N_1735);
xnor U7472 (N_7472,N_1136,N_2289);
or U7473 (N_7473,N_1631,N_1732);
nand U7474 (N_7474,N_4726,N_3596);
and U7475 (N_7475,N_1216,N_2328);
and U7476 (N_7476,N_4580,N_3182);
nor U7477 (N_7477,N_4961,N_2343);
or U7478 (N_7478,N_3443,N_4297);
or U7479 (N_7479,N_2620,N_302);
or U7480 (N_7480,N_3460,N_3028);
nor U7481 (N_7481,N_1640,N_3044);
nand U7482 (N_7482,N_1708,N_658);
or U7483 (N_7483,N_4231,N_4762);
and U7484 (N_7484,N_4067,N_2078);
or U7485 (N_7485,N_3645,N_2177);
or U7486 (N_7486,N_43,N_1530);
nand U7487 (N_7487,N_2911,N_1043);
nor U7488 (N_7488,N_1408,N_1859);
xor U7489 (N_7489,N_4210,N_1847);
and U7490 (N_7490,N_2088,N_3476);
or U7491 (N_7491,N_2243,N_2162);
or U7492 (N_7492,N_2072,N_1529);
xor U7493 (N_7493,N_881,N_3234);
nor U7494 (N_7494,N_4666,N_2112);
or U7495 (N_7495,N_2439,N_1877);
nand U7496 (N_7496,N_2631,N_2491);
nor U7497 (N_7497,N_539,N_4433);
nor U7498 (N_7498,N_2990,N_1844);
nand U7499 (N_7499,N_4774,N_208);
nand U7500 (N_7500,N_2474,N_195);
nor U7501 (N_7501,N_2882,N_369);
or U7502 (N_7502,N_3816,N_638);
and U7503 (N_7503,N_506,N_3712);
nor U7504 (N_7504,N_3559,N_1092);
xnor U7505 (N_7505,N_4469,N_3311);
and U7506 (N_7506,N_4698,N_2574);
nor U7507 (N_7507,N_4646,N_2020);
and U7508 (N_7508,N_4675,N_4235);
or U7509 (N_7509,N_2774,N_786);
nand U7510 (N_7510,N_2645,N_4919);
or U7511 (N_7511,N_2626,N_4345);
or U7512 (N_7512,N_330,N_4508);
nor U7513 (N_7513,N_816,N_4328);
xnor U7514 (N_7514,N_3438,N_4438);
nand U7515 (N_7515,N_3339,N_2825);
xor U7516 (N_7516,N_335,N_140);
and U7517 (N_7517,N_4146,N_3955);
nor U7518 (N_7518,N_2631,N_4612);
and U7519 (N_7519,N_4941,N_578);
nand U7520 (N_7520,N_4795,N_1782);
or U7521 (N_7521,N_1481,N_1636);
xnor U7522 (N_7522,N_2337,N_4307);
nor U7523 (N_7523,N_4397,N_684);
and U7524 (N_7524,N_1717,N_4047);
nand U7525 (N_7525,N_335,N_4758);
nor U7526 (N_7526,N_4486,N_1078);
nor U7527 (N_7527,N_978,N_3143);
and U7528 (N_7528,N_4613,N_4295);
and U7529 (N_7529,N_3713,N_3881);
xnor U7530 (N_7530,N_613,N_4743);
nor U7531 (N_7531,N_184,N_3998);
xnor U7532 (N_7532,N_3498,N_2297);
nor U7533 (N_7533,N_1088,N_1430);
nand U7534 (N_7534,N_2141,N_1097);
or U7535 (N_7535,N_2008,N_604);
nand U7536 (N_7536,N_1766,N_530);
or U7537 (N_7537,N_4702,N_2749);
nor U7538 (N_7538,N_1675,N_967);
nor U7539 (N_7539,N_479,N_1940);
nand U7540 (N_7540,N_735,N_3387);
and U7541 (N_7541,N_2353,N_4924);
and U7542 (N_7542,N_4352,N_2334);
and U7543 (N_7543,N_3005,N_2701);
nor U7544 (N_7544,N_1760,N_2987);
and U7545 (N_7545,N_3334,N_3866);
and U7546 (N_7546,N_438,N_4859);
or U7547 (N_7547,N_3877,N_3297);
and U7548 (N_7548,N_4592,N_3314);
xnor U7549 (N_7549,N_927,N_2168);
nor U7550 (N_7550,N_1127,N_2006);
and U7551 (N_7551,N_954,N_1691);
and U7552 (N_7552,N_654,N_1667);
nand U7553 (N_7553,N_450,N_4691);
or U7554 (N_7554,N_1358,N_1162);
nor U7555 (N_7555,N_3504,N_2657);
nand U7556 (N_7556,N_1578,N_1566);
or U7557 (N_7557,N_4971,N_4436);
and U7558 (N_7558,N_2239,N_4223);
nor U7559 (N_7559,N_2688,N_4055);
and U7560 (N_7560,N_1242,N_664);
nand U7561 (N_7561,N_3666,N_1606);
and U7562 (N_7562,N_3652,N_1603);
nor U7563 (N_7563,N_1121,N_2171);
nand U7564 (N_7564,N_1717,N_3601);
or U7565 (N_7565,N_3507,N_1059);
and U7566 (N_7566,N_3260,N_2881);
or U7567 (N_7567,N_4150,N_1729);
nor U7568 (N_7568,N_3443,N_4424);
nand U7569 (N_7569,N_2962,N_4392);
and U7570 (N_7570,N_382,N_1450);
nor U7571 (N_7571,N_523,N_2422);
nor U7572 (N_7572,N_2813,N_3608);
or U7573 (N_7573,N_3276,N_1045);
xnor U7574 (N_7574,N_4590,N_2662);
or U7575 (N_7575,N_2805,N_568);
and U7576 (N_7576,N_1477,N_1125);
nor U7577 (N_7577,N_4742,N_438);
and U7578 (N_7578,N_1771,N_973);
or U7579 (N_7579,N_1870,N_4973);
nand U7580 (N_7580,N_4361,N_3507);
and U7581 (N_7581,N_1663,N_2671);
xor U7582 (N_7582,N_3753,N_3743);
and U7583 (N_7583,N_3887,N_2031);
or U7584 (N_7584,N_2718,N_4760);
and U7585 (N_7585,N_1787,N_306);
or U7586 (N_7586,N_1362,N_3923);
and U7587 (N_7587,N_261,N_1173);
nand U7588 (N_7588,N_4809,N_1757);
nand U7589 (N_7589,N_4785,N_2278);
nand U7590 (N_7590,N_4251,N_2977);
nor U7591 (N_7591,N_2098,N_1500);
and U7592 (N_7592,N_1212,N_4622);
or U7593 (N_7593,N_1386,N_2977);
nor U7594 (N_7594,N_4943,N_3594);
nor U7595 (N_7595,N_2480,N_4072);
nor U7596 (N_7596,N_2228,N_1728);
and U7597 (N_7597,N_4205,N_2849);
and U7598 (N_7598,N_1103,N_3132);
xor U7599 (N_7599,N_486,N_2644);
or U7600 (N_7600,N_3364,N_1075);
or U7601 (N_7601,N_938,N_3854);
or U7602 (N_7602,N_3838,N_1316);
and U7603 (N_7603,N_1608,N_3997);
or U7604 (N_7604,N_533,N_4258);
and U7605 (N_7605,N_4417,N_179);
or U7606 (N_7606,N_3957,N_2230);
and U7607 (N_7607,N_2181,N_130);
xor U7608 (N_7608,N_2976,N_3631);
nor U7609 (N_7609,N_3394,N_555);
nand U7610 (N_7610,N_3562,N_1782);
and U7611 (N_7611,N_997,N_2767);
nand U7612 (N_7612,N_2447,N_1975);
nor U7613 (N_7613,N_2714,N_4579);
nand U7614 (N_7614,N_2873,N_3785);
nand U7615 (N_7615,N_3359,N_905);
or U7616 (N_7616,N_3778,N_3683);
xor U7617 (N_7617,N_1921,N_2385);
nand U7618 (N_7618,N_682,N_4983);
nor U7619 (N_7619,N_2239,N_4400);
or U7620 (N_7620,N_469,N_3373);
nor U7621 (N_7621,N_4598,N_3309);
nand U7622 (N_7622,N_4539,N_732);
nand U7623 (N_7623,N_4779,N_1828);
nor U7624 (N_7624,N_1988,N_4324);
nor U7625 (N_7625,N_1303,N_4856);
and U7626 (N_7626,N_4946,N_3895);
and U7627 (N_7627,N_49,N_2590);
xnor U7628 (N_7628,N_668,N_3270);
nand U7629 (N_7629,N_289,N_4507);
nand U7630 (N_7630,N_4161,N_4978);
and U7631 (N_7631,N_1151,N_3865);
nor U7632 (N_7632,N_302,N_1658);
or U7633 (N_7633,N_1457,N_2089);
or U7634 (N_7634,N_368,N_3605);
xnor U7635 (N_7635,N_1410,N_1682);
and U7636 (N_7636,N_839,N_4171);
or U7637 (N_7637,N_262,N_1883);
or U7638 (N_7638,N_3043,N_3770);
nand U7639 (N_7639,N_1752,N_3722);
and U7640 (N_7640,N_4618,N_4462);
or U7641 (N_7641,N_2239,N_4027);
nand U7642 (N_7642,N_4762,N_3093);
nor U7643 (N_7643,N_2669,N_4076);
or U7644 (N_7644,N_4031,N_2969);
xor U7645 (N_7645,N_3182,N_447);
nand U7646 (N_7646,N_3777,N_4832);
and U7647 (N_7647,N_2017,N_2113);
xor U7648 (N_7648,N_3198,N_773);
and U7649 (N_7649,N_2719,N_1865);
nor U7650 (N_7650,N_2529,N_4960);
nor U7651 (N_7651,N_4838,N_3417);
nor U7652 (N_7652,N_2112,N_3400);
or U7653 (N_7653,N_527,N_1906);
xnor U7654 (N_7654,N_1445,N_3544);
or U7655 (N_7655,N_559,N_4899);
and U7656 (N_7656,N_3,N_3173);
nand U7657 (N_7657,N_4077,N_4646);
and U7658 (N_7658,N_2996,N_1326);
nor U7659 (N_7659,N_2529,N_411);
nor U7660 (N_7660,N_3242,N_2800);
nor U7661 (N_7661,N_1317,N_314);
nand U7662 (N_7662,N_4180,N_3919);
and U7663 (N_7663,N_2827,N_273);
and U7664 (N_7664,N_2128,N_1362);
and U7665 (N_7665,N_53,N_3036);
nand U7666 (N_7666,N_534,N_1817);
nor U7667 (N_7667,N_1057,N_582);
and U7668 (N_7668,N_3322,N_2252);
and U7669 (N_7669,N_4783,N_4012);
or U7670 (N_7670,N_3726,N_2753);
or U7671 (N_7671,N_586,N_2731);
nor U7672 (N_7672,N_4226,N_262);
xnor U7673 (N_7673,N_4130,N_3126);
nand U7674 (N_7674,N_1370,N_2082);
nand U7675 (N_7675,N_4898,N_3702);
or U7676 (N_7676,N_416,N_2701);
and U7677 (N_7677,N_1158,N_4055);
or U7678 (N_7678,N_322,N_1895);
nor U7679 (N_7679,N_2752,N_3133);
xnor U7680 (N_7680,N_2961,N_3269);
xor U7681 (N_7681,N_3050,N_3954);
xor U7682 (N_7682,N_2225,N_3494);
and U7683 (N_7683,N_1945,N_2813);
or U7684 (N_7684,N_2067,N_4294);
nand U7685 (N_7685,N_1079,N_1313);
xor U7686 (N_7686,N_36,N_3187);
or U7687 (N_7687,N_2752,N_673);
nor U7688 (N_7688,N_3687,N_3744);
and U7689 (N_7689,N_4887,N_2053);
or U7690 (N_7690,N_568,N_2766);
nor U7691 (N_7691,N_2547,N_3382);
xor U7692 (N_7692,N_4854,N_2634);
or U7693 (N_7693,N_4125,N_4151);
xnor U7694 (N_7694,N_688,N_3894);
or U7695 (N_7695,N_3708,N_3511);
and U7696 (N_7696,N_4268,N_541);
nor U7697 (N_7697,N_2078,N_4420);
and U7698 (N_7698,N_3671,N_3814);
nand U7699 (N_7699,N_758,N_3918);
xnor U7700 (N_7700,N_4835,N_4848);
nor U7701 (N_7701,N_3696,N_1782);
or U7702 (N_7702,N_1991,N_3558);
nor U7703 (N_7703,N_2496,N_1602);
or U7704 (N_7704,N_4662,N_3385);
and U7705 (N_7705,N_3425,N_3036);
and U7706 (N_7706,N_1970,N_4861);
xor U7707 (N_7707,N_1270,N_2867);
nor U7708 (N_7708,N_2492,N_1040);
xor U7709 (N_7709,N_1521,N_458);
and U7710 (N_7710,N_4064,N_4991);
nor U7711 (N_7711,N_4988,N_4422);
and U7712 (N_7712,N_3127,N_1083);
nor U7713 (N_7713,N_1069,N_3256);
or U7714 (N_7714,N_1533,N_3213);
or U7715 (N_7715,N_2306,N_1394);
and U7716 (N_7716,N_335,N_4651);
or U7717 (N_7717,N_3982,N_2176);
nand U7718 (N_7718,N_760,N_4930);
xnor U7719 (N_7719,N_1203,N_4934);
nand U7720 (N_7720,N_1177,N_445);
and U7721 (N_7721,N_1345,N_3822);
and U7722 (N_7722,N_216,N_4832);
and U7723 (N_7723,N_3041,N_3771);
and U7724 (N_7724,N_159,N_1041);
and U7725 (N_7725,N_1898,N_4071);
nor U7726 (N_7726,N_727,N_3792);
nor U7727 (N_7727,N_546,N_3567);
nand U7728 (N_7728,N_3650,N_790);
and U7729 (N_7729,N_1041,N_833);
or U7730 (N_7730,N_4048,N_685);
nand U7731 (N_7731,N_4836,N_3808);
xor U7732 (N_7732,N_963,N_2709);
or U7733 (N_7733,N_3405,N_4318);
nor U7734 (N_7734,N_1638,N_4556);
and U7735 (N_7735,N_2997,N_2225);
and U7736 (N_7736,N_4198,N_1229);
xnor U7737 (N_7737,N_953,N_3526);
or U7738 (N_7738,N_3733,N_2667);
and U7739 (N_7739,N_980,N_2550);
nand U7740 (N_7740,N_1905,N_3124);
nand U7741 (N_7741,N_2887,N_1350);
and U7742 (N_7742,N_3589,N_4400);
nor U7743 (N_7743,N_98,N_354);
nor U7744 (N_7744,N_2038,N_2139);
xnor U7745 (N_7745,N_341,N_1257);
nor U7746 (N_7746,N_1175,N_3214);
nor U7747 (N_7747,N_1001,N_1303);
nor U7748 (N_7748,N_684,N_1336);
nor U7749 (N_7749,N_4794,N_603);
nand U7750 (N_7750,N_3761,N_1085);
nand U7751 (N_7751,N_2704,N_4589);
nor U7752 (N_7752,N_3082,N_1150);
or U7753 (N_7753,N_1425,N_1268);
and U7754 (N_7754,N_727,N_2802);
or U7755 (N_7755,N_2444,N_3189);
and U7756 (N_7756,N_1871,N_1484);
or U7757 (N_7757,N_26,N_3260);
nor U7758 (N_7758,N_4652,N_2143);
or U7759 (N_7759,N_4815,N_2664);
xor U7760 (N_7760,N_881,N_1558);
nand U7761 (N_7761,N_3517,N_4654);
nor U7762 (N_7762,N_1892,N_2561);
nor U7763 (N_7763,N_4588,N_1608);
nor U7764 (N_7764,N_3367,N_1652);
nor U7765 (N_7765,N_4553,N_4705);
nand U7766 (N_7766,N_3343,N_3530);
xnor U7767 (N_7767,N_2970,N_871);
nor U7768 (N_7768,N_4612,N_485);
and U7769 (N_7769,N_1708,N_3855);
and U7770 (N_7770,N_4822,N_1246);
nor U7771 (N_7771,N_3961,N_1540);
and U7772 (N_7772,N_4466,N_2472);
nor U7773 (N_7773,N_917,N_3825);
nand U7774 (N_7774,N_3404,N_2101);
nor U7775 (N_7775,N_1199,N_4131);
nand U7776 (N_7776,N_3415,N_4273);
nand U7777 (N_7777,N_782,N_4479);
nand U7778 (N_7778,N_667,N_1314);
and U7779 (N_7779,N_1313,N_3743);
nand U7780 (N_7780,N_4459,N_3319);
nor U7781 (N_7781,N_1409,N_2167);
and U7782 (N_7782,N_3256,N_3430);
nor U7783 (N_7783,N_3638,N_753);
and U7784 (N_7784,N_2207,N_4189);
nor U7785 (N_7785,N_1009,N_570);
nand U7786 (N_7786,N_1092,N_4077);
xnor U7787 (N_7787,N_1742,N_4364);
or U7788 (N_7788,N_98,N_3577);
and U7789 (N_7789,N_233,N_2937);
or U7790 (N_7790,N_942,N_2129);
nor U7791 (N_7791,N_3102,N_904);
or U7792 (N_7792,N_809,N_3715);
or U7793 (N_7793,N_2189,N_1796);
nand U7794 (N_7794,N_1606,N_2700);
and U7795 (N_7795,N_3914,N_3780);
xnor U7796 (N_7796,N_160,N_1319);
nor U7797 (N_7797,N_3403,N_3943);
nand U7798 (N_7798,N_307,N_2075);
nand U7799 (N_7799,N_2281,N_899);
and U7800 (N_7800,N_4191,N_728);
xor U7801 (N_7801,N_791,N_3314);
nor U7802 (N_7802,N_3716,N_4641);
xor U7803 (N_7803,N_3617,N_1348);
nor U7804 (N_7804,N_2201,N_3844);
or U7805 (N_7805,N_2175,N_3009);
and U7806 (N_7806,N_1044,N_1375);
or U7807 (N_7807,N_3856,N_1124);
or U7808 (N_7808,N_2518,N_3168);
and U7809 (N_7809,N_955,N_1390);
and U7810 (N_7810,N_4637,N_3812);
nand U7811 (N_7811,N_4946,N_1731);
nand U7812 (N_7812,N_4754,N_1635);
nand U7813 (N_7813,N_1264,N_2675);
and U7814 (N_7814,N_3874,N_1231);
or U7815 (N_7815,N_3744,N_798);
nand U7816 (N_7816,N_4951,N_3321);
and U7817 (N_7817,N_1254,N_4390);
or U7818 (N_7818,N_4242,N_4335);
or U7819 (N_7819,N_314,N_2922);
nor U7820 (N_7820,N_2386,N_627);
nor U7821 (N_7821,N_4374,N_4205);
nor U7822 (N_7822,N_2041,N_2043);
and U7823 (N_7823,N_4061,N_1627);
xor U7824 (N_7824,N_2179,N_2930);
nor U7825 (N_7825,N_1092,N_606);
and U7826 (N_7826,N_1802,N_339);
nor U7827 (N_7827,N_290,N_387);
nor U7828 (N_7828,N_3710,N_2324);
xnor U7829 (N_7829,N_1108,N_514);
xor U7830 (N_7830,N_2354,N_4771);
nor U7831 (N_7831,N_3677,N_4605);
nand U7832 (N_7832,N_1446,N_2505);
nand U7833 (N_7833,N_2890,N_3530);
nor U7834 (N_7834,N_3255,N_82);
and U7835 (N_7835,N_1402,N_1864);
nand U7836 (N_7836,N_1483,N_785);
nand U7837 (N_7837,N_2337,N_3324);
nor U7838 (N_7838,N_1230,N_1163);
or U7839 (N_7839,N_1164,N_790);
or U7840 (N_7840,N_4202,N_828);
xor U7841 (N_7841,N_1854,N_2981);
nand U7842 (N_7842,N_3926,N_2930);
and U7843 (N_7843,N_1500,N_4652);
nand U7844 (N_7844,N_4896,N_806);
xnor U7845 (N_7845,N_158,N_1604);
nand U7846 (N_7846,N_1693,N_1489);
or U7847 (N_7847,N_56,N_2174);
xor U7848 (N_7848,N_1271,N_213);
or U7849 (N_7849,N_365,N_2810);
nor U7850 (N_7850,N_4620,N_661);
or U7851 (N_7851,N_322,N_2377);
nand U7852 (N_7852,N_4348,N_14);
nand U7853 (N_7853,N_39,N_3520);
or U7854 (N_7854,N_1201,N_3841);
nor U7855 (N_7855,N_511,N_1997);
nor U7856 (N_7856,N_1259,N_1119);
or U7857 (N_7857,N_1762,N_2923);
nor U7858 (N_7858,N_628,N_2520);
nor U7859 (N_7859,N_2700,N_1654);
and U7860 (N_7860,N_602,N_3913);
or U7861 (N_7861,N_1648,N_1814);
nand U7862 (N_7862,N_4750,N_3545);
or U7863 (N_7863,N_3889,N_666);
or U7864 (N_7864,N_4467,N_3000);
nand U7865 (N_7865,N_2471,N_1687);
nor U7866 (N_7866,N_1255,N_4164);
nor U7867 (N_7867,N_321,N_814);
and U7868 (N_7868,N_645,N_1875);
nor U7869 (N_7869,N_3079,N_1581);
nand U7870 (N_7870,N_4670,N_1180);
xnor U7871 (N_7871,N_4415,N_2587);
nand U7872 (N_7872,N_4976,N_68);
nor U7873 (N_7873,N_172,N_3175);
nor U7874 (N_7874,N_859,N_3647);
and U7875 (N_7875,N_4543,N_4931);
or U7876 (N_7876,N_3834,N_3576);
nor U7877 (N_7877,N_1794,N_1842);
or U7878 (N_7878,N_2146,N_2732);
or U7879 (N_7879,N_1579,N_4510);
nand U7880 (N_7880,N_4848,N_3894);
nor U7881 (N_7881,N_4648,N_3384);
nand U7882 (N_7882,N_1614,N_2444);
nor U7883 (N_7883,N_3742,N_743);
and U7884 (N_7884,N_3656,N_1628);
nor U7885 (N_7885,N_1083,N_1445);
and U7886 (N_7886,N_4771,N_1636);
nand U7887 (N_7887,N_34,N_240);
nor U7888 (N_7888,N_1155,N_2733);
nand U7889 (N_7889,N_4597,N_4322);
xnor U7890 (N_7890,N_4151,N_681);
and U7891 (N_7891,N_3765,N_3924);
nand U7892 (N_7892,N_1271,N_1538);
and U7893 (N_7893,N_1051,N_3103);
or U7894 (N_7894,N_3987,N_3934);
or U7895 (N_7895,N_4219,N_1160);
or U7896 (N_7896,N_2578,N_1458);
nand U7897 (N_7897,N_2669,N_3438);
and U7898 (N_7898,N_3573,N_849);
nand U7899 (N_7899,N_3299,N_3016);
nor U7900 (N_7900,N_2476,N_176);
and U7901 (N_7901,N_3284,N_1983);
and U7902 (N_7902,N_1762,N_1090);
or U7903 (N_7903,N_2921,N_1885);
or U7904 (N_7904,N_1623,N_1602);
or U7905 (N_7905,N_4283,N_1260);
and U7906 (N_7906,N_435,N_4436);
xnor U7907 (N_7907,N_2807,N_1264);
and U7908 (N_7908,N_4646,N_3585);
nand U7909 (N_7909,N_3459,N_183);
or U7910 (N_7910,N_4324,N_4337);
nor U7911 (N_7911,N_4823,N_2821);
or U7912 (N_7912,N_2898,N_1213);
nor U7913 (N_7913,N_2173,N_2754);
and U7914 (N_7914,N_2384,N_84);
nand U7915 (N_7915,N_903,N_3701);
nand U7916 (N_7916,N_1688,N_3391);
or U7917 (N_7917,N_999,N_213);
and U7918 (N_7918,N_2195,N_497);
nand U7919 (N_7919,N_2815,N_1790);
xor U7920 (N_7920,N_3340,N_3457);
nand U7921 (N_7921,N_1501,N_2876);
and U7922 (N_7922,N_954,N_2595);
and U7923 (N_7923,N_186,N_3211);
nor U7924 (N_7924,N_409,N_2104);
or U7925 (N_7925,N_2411,N_4339);
or U7926 (N_7926,N_3923,N_3956);
nor U7927 (N_7927,N_2703,N_3036);
nor U7928 (N_7928,N_1299,N_1672);
nor U7929 (N_7929,N_2798,N_1896);
nor U7930 (N_7930,N_439,N_2079);
nor U7931 (N_7931,N_4350,N_1779);
nor U7932 (N_7932,N_3018,N_122);
or U7933 (N_7933,N_4909,N_4591);
and U7934 (N_7934,N_2056,N_4816);
and U7935 (N_7935,N_3949,N_2566);
nor U7936 (N_7936,N_1548,N_3415);
nor U7937 (N_7937,N_4099,N_3502);
nor U7938 (N_7938,N_1395,N_3686);
nand U7939 (N_7939,N_1548,N_1265);
nor U7940 (N_7940,N_4614,N_1155);
nand U7941 (N_7941,N_3995,N_3186);
and U7942 (N_7942,N_3675,N_1855);
or U7943 (N_7943,N_2636,N_1643);
nand U7944 (N_7944,N_2396,N_1286);
nand U7945 (N_7945,N_4699,N_4298);
or U7946 (N_7946,N_3236,N_4801);
or U7947 (N_7947,N_2057,N_3149);
nor U7948 (N_7948,N_3123,N_2448);
and U7949 (N_7949,N_148,N_3407);
or U7950 (N_7950,N_4560,N_4473);
nor U7951 (N_7951,N_2388,N_4734);
nand U7952 (N_7952,N_217,N_2405);
nor U7953 (N_7953,N_2532,N_3321);
nand U7954 (N_7954,N_2288,N_1098);
nor U7955 (N_7955,N_3743,N_3774);
or U7956 (N_7956,N_2420,N_892);
or U7957 (N_7957,N_512,N_2421);
nand U7958 (N_7958,N_2787,N_3708);
or U7959 (N_7959,N_4993,N_834);
nor U7960 (N_7960,N_922,N_4395);
and U7961 (N_7961,N_1644,N_2410);
nor U7962 (N_7962,N_614,N_1849);
xnor U7963 (N_7963,N_3142,N_3426);
nor U7964 (N_7964,N_4649,N_2188);
nand U7965 (N_7965,N_1509,N_2173);
nor U7966 (N_7966,N_4199,N_423);
and U7967 (N_7967,N_1105,N_1422);
or U7968 (N_7968,N_1420,N_3666);
nor U7969 (N_7969,N_1099,N_89);
nor U7970 (N_7970,N_4178,N_4877);
and U7971 (N_7971,N_3206,N_2512);
nand U7972 (N_7972,N_4479,N_618);
and U7973 (N_7973,N_1947,N_2711);
nor U7974 (N_7974,N_3531,N_1921);
or U7975 (N_7975,N_2461,N_4040);
nor U7976 (N_7976,N_3326,N_3685);
nor U7977 (N_7977,N_1730,N_2010);
and U7978 (N_7978,N_4070,N_2162);
and U7979 (N_7979,N_4555,N_2965);
or U7980 (N_7980,N_2925,N_1117);
or U7981 (N_7981,N_4722,N_133);
nor U7982 (N_7982,N_3033,N_855);
nand U7983 (N_7983,N_2836,N_4249);
and U7984 (N_7984,N_2870,N_4673);
xnor U7985 (N_7985,N_4378,N_414);
or U7986 (N_7986,N_3552,N_1775);
or U7987 (N_7987,N_4382,N_1374);
or U7988 (N_7988,N_1875,N_2282);
nand U7989 (N_7989,N_96,N_1349);
nand U7990 (N_7990,N_621,N_3215);
and U7991 (N_7991,N_555,N_2429);
and U7992 (N_7992,N_4911,N_2909);
and U7993 (N_7993,N_2180,N_3940);
nand U7994 (N_7994,N_4379,N_3896);
and U7995 (N_7995,N_1054,N_3193);
and U7996 (N_7996,N_4963,N_1377);
nand U7997 (N_7997,N_3665,N_4549);
nand U7998 (N_7998,N_4569,N_923);
nor U7999 (N_7999,N_2748,N_2281);
and U8000 (N_8000,N_1008,N_3100);
or U8001 (N_8001,N_1874,N_1369);
xnor U8002 (N_8002,N_4850,N_221);
or U8003 (N_8003,N_2109,N_561);
nor U8004 (N_8004,N_2923,N_2500);
nand U8005 (N_8005,N_2052,N_905);
and U8006 (N_8006,N_2465,N_2973);
xnor U8007 (N_8007,N_3548,N_358);
and U8008 (N_8008,N_3591,N_4247);
and U8009 (N_8009,N_3066,N_2299);
or U8010 (N_8010,N_3,N_4982);
nor U8011 (N_8011,N_4458,N_2020);
nand U8012 (N_8012,N_1298,N_4119);
nor U8013 (N_8013,N_3960,N_3676);
xor U8014 (N_8014,N_844,N_1875);
or U8015 (N_8015,N_2559,N_1436);
nor U8016 (N_8016,N_4175,N_1841);
or U8017 (N_8017,N_1131,N_1647);
xor U8018 (N_8018,N_3527,N_2946);
and U8019 (N_8019,N_4288,N_2938);
and U8020 (N_8020,N_2810,N_676);
nor U8021 (N_8021,N_3449,N_4703);
nor U8022 (N_8022,N_2713,N_1709);
nor U8023 (N_8023,N_4963,N_1609);
nand U8024 (N_8024,N_214,N_305);
or U8025 (N_8025,N_4524,N_672);
or U8026 (N_8026,N_1258,N_3159);
and U8027 (N_8027,N_109,N_1645);
or U8028 (N_8028,N_2670,N_596);
or U8029 (N_8029,N_1837,N_2177);
nor U8030 (N_8030,N_1892,N_3258);
nor U8031 (N_8031,N_839,N_4045);
nand U8032 (N_8032,N_3758,N_553);
nand U8033 (N_8033,N_242,N_1782);
nand U8034 (N_8034,N_1136,N_1321);
or U8035 (N_8035,N_3029,N_286);
nor U8036 (N_8036,N_3874,N_807);
and U8037 (N_8037,N_3497,N_1050);
nand U8038 (N_8038,N_2538,N_2553);
nand U8039 (N_8039,N_3424,N_597);
nor U8040 (N_8040,N_4278,N_94);
nand U8041 (N_8041,N_4157,N_3314);
or U8042 (N_8042,N_1582,N_3400);
nor U8043 (N_8043,N_290,N_4978);
or U8044 (N_8044,N_3632,N_2887);
and U8045 (N_8045,N_3230,N_1076);
and U8046 (N_8046,N_2018,N_1983);
nor U8047 (N_8047,N_998,N_1691);
and U8048 (N_8048,N_875,N_2257);
and U8049 (N_8049,N_1409,N_3055);
and U8050 (N_8050,N_3714,N_4708);
nand U8051 (N_8051,N_148,N_2628);
nand U8052 (N_8052,N_238,N_412);
or U8053 (N_8053,N_3718,N_546);
or U8054 (N_8054,N_3814,N_3853);
nand U8055 (N_8055,N_775,N_540);
nor U8056 (N_8056,N_2746,N_4647);
nand U8057 (N_8057,N_3094,N_4546);
and U8058 (N_8058,N_3188,N_989);
nand U8059 (N_8059,N_3393,N_349);
xnor U8060 (N_8060,N_3435,N_4139);
nor U8061 (N_8061,N_1620,N_4946);
nor U8062 (N_8062,N_4241,N_4609);
xor U8063 (N_8063,N_3126,N_3060);
nor U8064 (N_8064,N_2618,N_3549);
or U8065 (N_8065,N_4776,N_1464);
nand U8066 (N_8066,N_213,N_1078);
and U8067 (N_8067,N_2843,N_1783);
and U8068 (N_8068,N_194,N_2144);
nand U8069 (N_8069,N_4984,N_3441);
and U8070 (N_8070,N_4488,N_3278);
nor U8071 (N_8071,N_2542,N_218);
and U8072 (N_8072,N_2650,N_4684);
and U8073 (N_8073,N_734,N_4833);
nor U8074 (N_8074,N_2985,N_3947);
nand U8075 (N_8075,N_4489,N_3215);
xor U8076 (N_8076,N_2898,N_712);
or U8077 (N_8077,N_3109,N_3647);
or U8078 (N_8078,N_3868,N_18);
xor U8079 (N_8079,N_3722,N_1463);
or U8080 (N_8080,N_2802,N_4422);
or U8081 (N_8081,N_1094,N_3790);
nor U8082 (N_8082,N_627,N_2800);
and U8083 (N_8083,N_3473,N_1397);
and U8084 (N_8084,N_99,N_2274);
nor U8085 (N_8085,N_937,N_2902);
nand U8086 (N_8086,N_2652,N_3899);
or U8087 (N_8087,N_61,N_4320);
or U8088 (N_8088,N_1525,N_2876);
xor U8089 (N_8089,N_3233,N_3585);
or U8090 (N_8090,N_528,N_4970);
and U8091 (N_8091,N_279,N_4878);
or U8092 (N_8092,N_867,N_3317);
nand U8093 (N_8093,N_3612,N_67);
nor U8094 (N_8094,N_1610,N_3667);
nor U8095 (N_8095,N_395,N_3268);
or U8096 (N_8096,N_384,N_605);
xor U8097 (N_8097,N_4518,N_1072);
nand U8098 (N_8098,N_944,N_466);
or U8099 (N_8099,N_2294,N_1752);
nand U8100 (N_8100,N_3702,N_1665);
or U8101 (N_8101,N_4523,N_3667);
xor U8102 (N_8102,N_3898,N_1506);
nor U8103 (N_8103,N_4347,N_653);
or U8104 (N_8104,N_1320,N_2101);
nor U8105 (N_8105,N_4048,N_2714);
and U8106 (N_8106,N_778,N_3066);
and U8107 (N_8107,N_4848,N_1248);
nor U8108 (N_8108,N_1815,N_2649);
nand U8109 (N_8109,N_4203,N_4041);
nand U8110 (N_8110,N_3556,N_3131);
or U8111 (N_8111,N_1393,N_2140);
and U8112 (N_8112,N_3452,N_4978);
and U8113 (N_8113,N_492,N_3279);
nand U8114 (N_8114,N_4076,N_4275);
or U8115 (N_8115,N_4765,N_41);
xor U8116 (N_8116,N_2464,N_1164);
and U8117 (N_8117,N_380,N_3239);
nand U8118 (N_8118,N_3425,N_3552);
or U8119 (N_8119,N_655,N_3883);
nor U8120 (N_8120,N_2228,N_3896);
nand U8121 (N_8121,N_2669,N_1366);
nor U8122 (N_8122,N_2722,N_1568);
nand U8123 (N_8123,N_3840,N_1427);
nand U8124 (N_8124,N_2116,N_1453);
or U8125 (N_8125,N_539,N_4764);
nand U8126 (N_8126,N_16,N_357);
nand U8127 (N_8127,N_3202,N_555);
nand U8128 (N_8128,N_544,N_3326);
and U8129 (N_8129,N_1008,N_3901);
and U8130 (N_8130,N_161,N_4645);
and U8131 (N_8131,N_3071,N_420);
and U8132 (N_8132,N_3048,N_1636);
and U8133 (N_8133,N_163,N_3823);
nand U8134 (N_8134,N_3340,N_4555);
nor U8135 (N_8135,N_2420,N_1870);
and U8136 (N_8136,N_3434,N_1182);
or U8137 (N_8137,N_3130,N_3977);
nand U8138 (N_8138,N_3314,N_415);
or U8139 (N_8139,N_154,N_951);
or U8140 (N_8140,N_203,N_219);
nand U8141 (N_8141,N_4065,N_1676);
and U8142 (N_8142,N_417,N_2216);
or U8143 (N_8143,N_2982,N_1432);
nand U8144 (N_8144,N_2673,N_2885);
or U8145 (N_8145,N_2600,N_1910);
or U8146 (N_8146,N_297,N_4745);
xnor U8147 (N_8147,N_668,N_4462);
nor U8148 (N_8148,N_313,N_4639);
and U8149 (N_8149,N_609,N_245);
and U8150 (N_8150,N_186,N_4987);
or U8151 (N_8151,N_1829,N_1536);
nor U8152 (N_8152,N_1056,N_395);
or U8153 (N_8153,N_4884,N_3706);
and U8154 (N_8154,N_2803,N_2412);
nor U8155 (N_8155,N_2231,N_3318);
and U8156 (N_8156,N_1312,N_1576);
or U8157 (N_8157,N_409,N_1759);
nor U8158 (N_8158,N_3905,N_4367);
nand U8159 (N_8159,N_1442,N_2862);
nor U8160 (N_8160,N_924,N_4600);
and U8161 (N_8161,N_799,N_2173);
nor U8162 (N_8162,N_1895,N_1863);
xor U8163 (N_8163,N_1175,N_4528);
and U8164 (N_8164,N_3466,N_755);
nand U8165 (N_8165,N_4738,N_242);
nor U8166 (N_8166,N_4903,N_1688);
nor U8167 (N_8167,N_3889,N_4359);
and U8168 (N_8168,N_349,N_2954);
nand U8169 (N_8169,N_2614,N_4694);
or U8170 (N_8170,N_4460,N_3834);
xor U8171 (N_8171,N_4912,N_4950);
nand U8172 (N_8172,N_4173,N_2502);
nor U8173 (N_8173,N_2536,N_2217);
xor U8174 (N_8174,N_238,N_1557);
nand U8175 (N_8175,N_1619,N_410);
or U8176 (N_8176,N_4199,N_2143);
and U8177 (N_8177,N_1747,N_3989);
nor U8178 (N_8178,N_4086,N_1518);
nor U8179 (N_8179,N_3758,N_4261);
or U8180 (N_8180,N_3127,N_3133);
or U8181 (N_8181,N_843,N_611);
and U8182 (N_8182,N_1893,N_1928);
nand U8183 (N_8183,N_2573,N_4200);
xor U8184 (N_8184,N_2843,N_4611);
nor U8185 (N_8185,N_3838,N_2915);
or U8186 (N_8186,N_1652,N_2845);
nor U8187 (N_8187,N_2423,N_2871);
xor U8188 (N_8188,N_2238,N_3526);
nor U8189 (N_8189,N_1088,N_4191);
nand U8190 (N_8190,N_2506,N_2446);
nor U8191 (N_8191,N_4999,N_2917);
and U8192 (N_8192,N_2153,N_2694);
or U8193 (N_8193,N_4000,N_2868);
and U8194 (N_8194,N_1066,N_1009);
and U8195 (N_8195,N_2307,N_2367);
xor U8196 (N_8196,N_4491,N_1900);
nand U8197 (N_8197,N_3104,N_4736);
nor U8198 (N_8198,N_784,N_1759);
nor U8199 (N_8199,N_4950,N_3989);
xnor U8200 (N_8200,N_3887,N_2678);
and U8201 (N_8201,N_4274,N_4359);
nor U8202 (N_8202,N_1460,N_3126);
and U8203 (N_8203,N_685,N_997);
nor U8204 (N_8204,N_1900,N_3359);
xor U8205 (N_8205,N_2940,N_1393);
nand U8206 (N_8206,N_462,N_354);
or U8207 (N_8207,N_3575,N_4769);
and U8208 (N_8208,N_1649,N_922);
or U8209 (N_8209,N_494,N_4225);
or U8210 (N_8210,N_2707,N_4355);
xor U8211 (N_8211,N_4089,N_642);
or U8212 (N_8212,N_633,N_315);
xnor U8213 (N_8213,N_4038,N_752);
nand U8214 (N_8214,N_3672,N_4998);
and U8215 (N_8215,N_3720,N_3576);
nand U8216 (N_8216,N_134,N_3777);
or U8217 (N_8217,N_882,N_2606);
and U8218 (N_8218,N_2584,N_704);
or U8219 (N_8219,N_484,N_4627);
or U8220 (N_8220,N_541,N_4293);
or U8221 (N_8221,N_4614,N_137);
nand U8222 (N_8222,N_1803,N_4494);
or U8223 (N_8223,N_3694,N_1811);
nor U8224 (N_8224,N_2820,N_274);
or U8225 (N_8225,N_2024,N_1245);
nand U8226 (N_8226,N_872,N_803);
or U8227 (N_8227,N_3404,N_3832);
nand U8228 (N_8228,N_3521,N_4385);
nand U8229 (N_8229,N_4565,N_4452);
nand U8230 (N_8230,N_400,N_4963);
xnor U8231 (N_8231,N_3537,N_3372);
xor U8232 (N_8232,N_2297,N_729);
or U8233 (N_8233,N_1810,N_2212);
nor U8234 (N_8234,N_969,N_4293);
nand U8235 (N_8235,N_4727,N_681);
nor U8236 (N_8236,N_3098,N_952);
nand U8237 (N_8237,N_2350,N_504);
nor U8238 (N_8238,N_3846,N_4538);
nand U8239 (N_8239,N_4208,N_50);
nand U8240 (N_8240,N_893,N_4022);
or U8241 (N_8241,N_844,N_296);
or U8242 (N_8242,N_4553,N_2964);
and U8243 (N_8243,N_3433,N_2594);
nand U8244 (N_8244,N_2713,N_4293);
nand U8245 (N_8245,N_3974,N_4403);
nor U8246 (N_8246,N_4285,N_3546);
nand U8247 (N_8247,N_3206,N_3888);
nand U8248 (N_8248,N_3009,N_2848);
or U8249 (N_8249,N_2794,N_4593);
nor U8250 (N_8250,N_4141,N_4795);
and U8251 (N_8251,N_939,N_4964);
nand U8252 (N_8252,N_562,N_3794);
nand U8253 (N_8253,N_2130,N_4214);
or U8254 (N_8254,N_1882,N_3);
nand U8255 (N_8255,N_1883,N_1710);
nor U8256 (N_8256,N_808,N_4832);
and U8257 (N_8257,N_1734,N_2169);
and U8258 (N_8258,N_3485,N_2773);
or U8259 (N_8259,N_1493,N_2110);
nor U8260 (N_8260,N_3005,N_3594);
nand U8261 (N_8261,N_3116,N_1828);
or U8262 (N_8262,N_3,N_106);
or U8263 (N_8263,N_83,N_2309);
and U8264 (N_8264,N_1884,N_2454);
xor U8265 (N_8265,N_3765,N_57);
or U8266 (N_8266,N_4174,N_2183);
nand U8267 (N_8267,N_153,N_226);
nor U8268 (N_8268,N_2261,N_263);
or U8269 (N_8269,N_4068,N_999);
and U8270 (N_8270,N_3686,N_2920);
xnor U8271 (N_8271,N_136,N_1369);
nand U8272 (N_8272,N_3689,N_834);
and U8273 (N_8273,N_1577,N_1333);
nor U8274 (N_8274,N_535,N_770);
and U8275 (N_8275,N_1047,N_1879);
nand U8276 (N_8276,N_4155,N_1858);
and U8277 (N_8277,N_1168,N_4238);
xor U8278 (N_8278,N_474,N_1303);
xnor U8279 (N_8279,N_3704,N_921);
nor U8280 (N_8280,N_3830,N_1144);
nand U8281 (N_8281,N_1180,N_251);
xor U8282 (N_8282,N_2518,N_1997);
and U8283 (N_8283,N_4168,N_1507);
and U8284 (N_8284,N_749,N_4972);
nand U8285 (N_8285,N_735,N_2701);
and U8286 (N_8286,N_4234,N_913);
nor U8287 (N_8287,N_3525,N_1588);
nand U8288 (N_8288,N_888,N_1318);
nand U8289 (N_8289,N_1059,N_2346);
or U8290 (N_8290,N_3677,N_1942);
nand U8291 (N_8291,N_291,N_775);
and U8292 (N_8292,N_1104,N_4914);
nand U8293 (N_8293,N_4503,N_3271);
nand U8294 (N_8294,N_1206,N_3710);
and U8295 (N_8295,N_4494,N_1425);
and U8296 (N_8296,N_294,N_4463);
or U8297 (N_8297,N_38,N_3050);
xor U8298 (N_8298,N_3951,N_353);
and U8299 (N_8299,N_1749,N_383);
xor U8300 (N_8300,N_1096,N_3375);
and U8301 (N_8301,N_3919,N_2866);
or U8302 (N_8302,N_2215,N_4653);
xor U8303 (N_8303,N_3058,N_4911);
nor U8304 (N_8304,N_4742,N_112);
or U8305 (N_8305,N_1084,N_3939);
nor U8306 (N_8306,N_4284,N_2137);
nor U8307 (N_8307,N_983,N_874);
or U8308 (N_8308,N_2586,N_1487);
and U8309 (N_8309,N_4058,N_3127);
or U8310 (N_8310,N_1843,N_3731);
and U8311 (N_8311,N_2105,N_2583);
nor U8312 (N_8312,N_2241,N_4832);
nor U8313 (N_8313,N_232,N_3181);
and U8314 (N_8314,N_2508,N_1164);
nand U8315 (N_8315,N_3474,N_782);
or U8316 (N_8316,N_760,N_3075);
nand U8317 (N_8317,N_4439,N_2764);
and U8318 (N_8318,N_3471,N_4781);
xor U8319 (N_8319,N_1762,N_4408);
and U8320 (N_8320,N_937,N_3502);
or U8321 (N_8321,N_1035,N_2560);
nand U8322 (N_8322,N_714,N_443);
nor U8323 (N_8323,N_3472,N_111);
xnor U8324 (N_8324,N_2370,N_4584);
or U8325 (N_8325,N_3386,N_3044);
xnor U8326 (N_8326,N_2127,N_1419);
nand U8327 (N_8327,N_4931,N_4476);
nor U8328 (N_8328,N_2342,N_1448);
or U8329 (N_8329,N_1983,N_1114);
or U8330 (N_8330,N_2815,N_3504);
nand U8331 (N_8331,N_1402,N_200);
xnor U8332 (N_8332,N_4908,N_353);
nand U8333 (N_8333,N_2727,N_4908);
and U8334 (N_8334,N_1253,N_4067);
xnor U8335 (N_8335,N_630,N_2133);
nand U8336 (N_8336,N_2147,N_674);
xnor U8337 (N_8337,N_553,N_2954);
and U8338 (N_8338,N_2521,N_645);
nand U8339 (N_8339,N_3418,N_1736);
nand U8340 (N_8340,N_2115,N_3803);
nand U8341 (N_8341,N_1422,N_1039);
nor U8342 (N_8342,N_893,N_4729);
or U8343 (N_8343,N_616,N_4390);
or U8344 (N_8344,N_153,N_118);
nor U8345 (N_8345,N_4115,N_1289);
or U8346 (N_8346,N_2341,N_4701);
or U8347 (N_8347,N_3198,N_1567);
nand U8348 (N_8348,N_1609,N_4168);
and U8349 (N_8349,N_3612,N_3765);
or U8350 (N_8350,N_1399,N_3868);
and U8351 (N_8351,N_1313,N_2891);
nor U8352 (N_8352,N_2020,N_4074);
or U8353 (N_8353,N_946,N_4220);
or U8354 (N_8354,N_3317,N_4768);
nand U8355 (N_8355,N_1992,N_3782);
nor U8356 (N_8356,N_3232,N_1920);
or U8357 (N_8357,N_3196,N_1858);
nor U8358 (N_8358,N_4883,N_4543);
or U8359 (N_8359,N_421,N_616);
xor U8360 (N_8360,N_2264,N_2524);
and U8361 (N_8361,N_4196,N_520);
or U8362 (N_8362,N_1112,N_1069);
nor U8363 (N_8363,N_2964,N_3135);
or U8364 (N_8364,N_304,N_466);
nand U8365 (N_8365,N_2258,N_1966);
and U8366 (N_8366,N_2202,N_2439);
and U8367 (N_8367,N_391,N_2954);
nor U8368 (N_8368,N_2673,N_1185);
xor U8369 (N_8369,N_1838,N_4645);
nand U8370 (N_8370,N_1826,N_3072);
and U8371 (N_8371,N_344,N_1887);
nor U8372 (N_8372,N_2938,N_4870);
nor U8373 (N_8373,N_2282,N_2426);
or U8374 (N_8374,N_1338,N_2957);
and U8375 (N_8375,N_4077,N_4671);
nor U8376 (N_8376,N_3486,N_2685);
and U8377 (N_8377,N_3861,N_3642);
nand U8378 (N_8378,N_4761,N_2525);
nor U8379 (N_8379,N_563,N_3973);
nand U8380 (N_8380,N_2081,N_446);
nor U8381 (N_8381,N_2134,N_261);
nand U8382 (N_8382,N_2797,N_1223);
or U8383 (N_8383,N_2031,N_3664);
and U8384 (N_8384,N_236,N_1040);
and U8385 (N_8385,N_2136,N_2076);
or U8386 (N_8386,N_2869,N_3681);
or U8387 (N_8387,N_1037,N_2668);
nand U8388 (N_8388,N_4314,N_4289);
and U8389 (N_8389,N_3392,N_4377);
nor U8390 (N_8390,N_3337,N_3847);
nor U8391 (N_8391,N_3496,N_1972);
or U8392 (N_8392,N_3202,N_1678);
xor U8393 (N_8393,N_236,N_4278);
nand U8394 (N_8394,N_525,N_3969);
nor U8395 (N_8395,N_3497,N_4250);
nor U8396 (N_8396,N_4491,N_1057);
or U8397 (N_8397,N_1707,N_1307);
nor U8398 (N_8398,N_2060,N_983);
and U8399 (N_8399,N_3005,N_4193);
nor U8400 (N_8400,N_1621,N_88);
nand U8401 (N_8401,N_4016,N_1059);
nor U8402 (N_8402,N_2857,N_1741);
nor U8403 (N_8403,N_932,N_444);
nor U8404 (N_8404,N_4895,N_114);
xor U8405 (N_8405,N_4183,N_4724);
nand U8406 (N_8406,N_2669,N_1738);
nand U8407 (N_8407,N_1919,N_1391);
and U8408 (N_8408,N_382,N_2513);
or U8409 (N_8409,N_1694,N_1546);
and U8410 (N_8410,N_2701,N_925);
xnor U8411 (N_8411,N_2468,N_3010);
nand U8412 (N_8412,N_4968,N_875);
nor U8413 (N_8413,N_1297,N_4394);
nor U8414 (N_8414,N_3115,N_1635);
nor U8415 (N_8415,N_1474,N_1911);
nor U8416 (N_8416,N_1805,N_1166);
xor U8417 (N_8417,N_4229,N_1681);
and U8418 (N_8418,N_3884,N_1103);
and U8419 (N_8419,N_1395,N_185);
nand U8420 (N_8420,N_4690,N_918);
nor U8421 (N_8421,N_4576,N_2180);
or U8422 (N_8422,N_1647,N_3542);
xor U8423 (N_8423,N_3466,N_4469);
and U8424 (N_8424,N_4897,N_4483);
nor U8425 (N_8425,N_3949,N_4185);
nand U8426 (N_8426,N_1542,N_4368);
nor U8427 (N_8427,N_4652,N_2055);
nand U8428 (N_8428,N_3147,N_676);
nor U8429 (N_8429,N_2304,N_3474);
xnor U8430 (N_8430,N_3136,N_450);
nor U8431 (N_8431,N_233,N_4372);
and U8432 (N_8432,N_4990,N_2830);
and U8433 (N_8433,N_3614,N_1874);
and U8434 (N_8434,N_1858,N_1759);
nand U8435 (N_8435,N_2344,N_4108);
nand U8436 (N_8436,N_440,N_2446);
nor U8437 (N_8437,N_2851,N_2104);
and U8438 (N_8438,N_4541,N_3405);
nand U8439 (N_8439,N_556,N_2914);
nand U8440 (N_8440,N_53,N_1319);
or U8441 (N_8441,N_4129,N_1989);
and U8442 (N_8442,N_1903,N_3790);
or U8443 (N_8443,N_1616,N_3304);
nand U8444 (N_8444,N_3261,N_4210);
nand U8445 (N_8445,N_475,N_1781);
nor U8446 (N_8446,N_3933,N_2251);
and U8447 (N_8447,N_2562,N_1753);
or U8448 (N_8448,N_743,N_3370);
and U8449 (N_8449,N_2263,N_1161);
xnor U8450 (N_8450,N_921,N_1755);
or U8451 (N_8451,N_2084,N_4840);
nor U8452 (N_8452,N_2037,N_3642);
nor U8453 (N_8453,N_427,N_1710);
nand U8454 (N_8454,N_4956,N_798);
or U8455 (N_8455,N_2811,N_3405);
nor U8456 (N_8456,N_2909,N_3359);
nand U8457 (N_8457,N_4148,N_752);
xnor U8458 (N_8458,N_1857,N_1866);
nand U8459 (N_8459,N_531,N_802);
or U8460 (N_8460,N_4053,N_3312);
and U8461 (N_8461,N_3793,N_131);
or U8462 (N_8462,N_4490,N_1406);
xor U8463 (N_8463,N_272,N_2538);
nand U8464 (N_8464,N_3074,N_984);
xnor U8465 (N_8465,N_1569,N_1128);
or U8466 (N_8466,N_1229,N_535);
nand U8467 (N_8467,N_854,N_4199);
nand U8468 (N_8468,N_2019,N_3390);
nor U8469 (N_8469,N_4494,N_1144);
or U8470 (N_8470,N_4476,N_3382);
nor U8471 (N_8471,N_1223,N_1528);
and U8472 (N_8472,N_1113,N_3197);
and U8473 (N_8473,N_2809,N_2684);
or U8474 (N_8474,N_2839,N_1013);
or U8475 (N_8475,N_1226,N_2199);
nand U8476 (N_8476,N_3004,N_1441);
and U8477 (N_8477,N_2748,N_328);
and U8478 (N_8478,N_3866,N_3045);
xnor U8479 (N_8479,N_336,N_2283);
or U8480 (N_8480,N_1143,N_3019);
and U8481 (N_8481,N_1051,N_2245);
nor U8482 (N_8482,N_1865,N_3931);
and U8483 (N_8483,N_4663,N_3533);
or U8484 (N_8484,N_1758,N_2981);
nand U8485 (N_8485,N_3440,N_4076);
and U8486 (N_8486,N_4565,N_792);
xnor U8487 (N_8487,N_4972,N_357);
or U8488 (N_8488,N_865,N_2251);
nor U8489 (N_8489,N_1603,N_4450);
xnor U8490 (N_8490,N_4509,N_2417);
or U8491 (N_8491,N_2759,N_2105);
or U8492 (N_8492,N_1504,N_193);
and U8493 (N_8493,N_777,N_4427);
nor U8494 (N_8494,N_1228,N_1786);
or U8495 (N_8495,N_4787,N_4747);
and U8496 (N_8496,N_239,N_1884);
and U8497 (N_8497,N_674,N_1287);
nand U8498 (N_8498,N_3123,N_918);
and U8499 (N_8499,N_909,N_2743);
and U8500 (N_8500,N_2769,N_2228);
xor U8501 (N_8501,N_2282,N_45);
and U8502 (N_8502,N_1760,N_637);
xnor U8503 (N_8503,N_4137,N_3441);
and U8504 (N_8504,N_436,N_2851);
nand U8505 (N_8505,N_4796,N_221);
and U8506 (N_8506,N_3378,N_758);
and U8507 (N_8507,N_3400,N_4934);
nor U8508 (N_8508,N_823,N_662);
or U8509 (N_8509,N_740,N_3592);
and U8510 (N_8510,N_122,N_3014);
xor U8511 (N_8511,N_2827,N_2747);
nand U8512 (N_8512,N_3925,N_1428);
nand U8513 (N_8513,N_4335,N_3790);
and U8514 (N_8514,N_1233,N_2348);
nand U8515 (N_8515,N_2532,N_2711);
nand U8516 (N_8516,N_4497,N_2982);
nor U8517 (N_8517,N_2357,N_2076);
xnor U8518 (N_8518,N_3479,N_3151);
and U8519 (N_8519,N_1652,N_4055);
and U8520 (N_8520,N_4813,N_4166);
and U8521 (N_8521,N_1490,N_3556);
nand U8522 (N_8522,N_3707,N_1497);
and U8523 (N_8523,N_821,N_4805);
or U8524 (N_8524,N_3016,N_4269);
and U8525 (N_8525,N_1923,N_957);
or U8526 (N_8526,N_597,N_3438);
or U8527 (N_8527,N_1683,N_2359);
or U8528 (N_8528,N_4979,N_2078);
xor U8529 (N_8529,N_4930,N_2261);
and U8530 (N_8530,N_930,N_1175);
or U8531 (N_8531,N_1155,N_1119);
xor U8532 (N_8532,N_1641,N_4947);
nand U8533 (N_8533,N_839,N_3151);
and U8534 (N_8534,N_4929,N_173);
or U8535 (N_8535,N_2621,N_4626);
and U8536 (N_8536,N_3539,N_1313);
and U8537 (N_8537,N_4211,N_4422);
nand U8538 (N_8538,N_873,N_811);
or U8539 (N_8539,N_968,N_2339);
nor U8540 (N_8540,N_823,N_340);
xnor U8541 (N_8541,N_2134,N_2292);
nand U8542 (N_8542,N_1256,N_3676);
nor U8543 (N_8543,N_1035,N_2023);
nor U8544 (N_8544,N_4021,N_4373);
or U8545 (N_8545,N_4804,N_822);
xnor U8546 (N_8546,N_418,N_2876);
or U8547 (N_8547,N_953,N_1597);
nand U8548 (N_8548,N_1262,N_328);
or U8549 (N_8549,N_71,N_1859);
and U8550 (N_8550,N_833,N_4012);
and U8551 (N_8551,N_4399,N_2675);
nand U8552 (N_8552,N_768,N_3120);
or U8553 (N_8553,N_4041,N_1588);
and U8554 (N_8554,N_3689,N_4010);
or U8555 (N_8555,N_532,N_1770);
or U8556 (N_8556,N_3473,N_1391);
or U8557 (N_8557,N_4908,N_3922);
or U8558 (N_8558,N_2006,N_2197);
and U8559 (N_8559,N_140,N_1146);
or U8560 (N_8560,N_768,N_3486);
nand U8561 (N_8561,N_4953,N_2568);
xnor U8562 (N_8562,N_4276,N_4069);
and U8563 (N_8563,N_4870,N_4635);
nand U8564 (N_8564,N_2393,N_4626);
or U8565 (N_8565,N_369,N_3467);
nor U8566 (N_8566,N_3383,N_1172);
or U8567 (N_8567,N_3844,N_198);
nand U8568 (N_8568,N_2651,N_606);
and U8569 (N_8569,N_1097,N_3333);
or U8570 (N_8570,N_4034,N_3940);
nor U8571 (N_8571,N_1034,N_2773);
nor U8572 (N_8572,N_4752,N_2219);
or U8573 (N_8573,N_1561,N_2801);
or U8574 (N_8574,N_4665,N_3416);
or U8575 (N_8575,N_4005,N_4884);
nand U8576 (N_8576,N_463,N_4234);
or U8577 (N_8577,N_2003,N_384);
nand U8578 (N_8578,N_4582,N_3531);
nand U8579 (N_8579,N_1361,N_1812);
nor U8580 (N_8580,N_2407,N_2363);
or U8581 (N_8581,N_3267,N_897);
nor U8582 (N_8582,N_1636,N_4065);
or U8583 (N_8583,N_1068,N_639);
nor U8584 (N_8584,N_2114,N_4560);
nor U8585 (N_8585,N_3748,N_3803);
and U8586 (N_8586,N_108,N_1630);
and U8587 (N_8587,N_2154,N_3606);
and U8588 (N_8588,N_738,N_3299);
or U8589 (N_8589,N_3015,N_2750);
xor U8590 (N_8590,N_4549,N_3004);
nand U8591 (N_8591,N_2241,N_1392);
nand U8592 (N_8592,N_2797,N_4703);
or U8593 (N_8593,N_3854,N_198);
and U8594 (N_8594,N_979,N_270);
nand U8595 (N_8595,N_4914,N_3506);
or U8596 (N_8596,N_227,N_4767);
nor U8597 (N_8597,N_3558,N_3304);
nor U8598 (N_8598,N_2979,N_4147);
nor U8599 (N_8599,N_1230,N_3354);
nor U8600 (N_8600,N_3226,N_4486);
xnor U8601 (N_8601,N_1710,N_405);
or U8602 (N_8602,N_3396,N_4495);
xor U8603 (N_8603,N_4899,N_1808);
nor U8604 (N_8604,N_46,N_1277);
or U8605 (N_8605,N_3133,N_1944);
and U8606 (N_8606,N_3616,N_4735);
nand U8607 (N_8607,N_557,N_3615);
and U8608 (N_8608,N_286,N_956);
and U8609 (N_8609,N_808,N_4325);
nor U8610 (N_8610,N_2933,N_1218);
nor U8611 (N_8611,N_712,N_2473);
or U8612 (N_8612,N_1152,N_4723);
or U8613 (N_8613,N_2686,N_1601);
nand U8614 (N_8614,N_3472,N_154);
or U8615 (N_8615,N_1870,N_1096);
nor U8616 (N_8616,N_4984,N_463);
or U8617 (N_8617,N_3191,N_3582);
and U8618 (N_8618,N_1060,N_4094);
nor U8619 (N_8619,N_3085,N_1899);
and U8620 (N_8620,N_4383,N_3786);
or U8621 (N_8621,N_3932,N_4234);
and U8622 (N_8622,N_3393,N_2429);
and U8623 (N_8623,N_4903,N_196);
or U8624 (N_8624,N_4467,N_4204);
xor U8625 (N_8625,N_408,N_1313);
and U8626 (N_8626,N_572,N_3158);
and U8627 (N_8627,N_1049,N_4661);
nand U8628 (N_8628,N_3206,N_3231);
nand U8629 (N_8629,N_2064,N_3167);
nand U8630 (N_8630,N_4563,N_741);
and U8631 (N_8631,N_4949,N_1113);
or U8632 (N_8632,N_3146,N_2270);
xnor U8633 (N_8633,N_4686,N_3341);
and U8634 (N_8634,N_1902,N_1942);
and U8635 (N_8635,N_1163,N_1111);
nor U8636 (N_8636,N_2050,N_2);
nand U8637 (N_8637,N_1055,N_4398);
and U8638 (N_8638,N_570,N_1406);
or U8639 (N_8639,N_1282,N_1254);
xor U8640 (N_8640,N_3978,N_910);
nor U8641 (N_8641,N_4344,N_4955);
nor U8642 (N_8642,N_4139,N_1943);
or U8643 (N_8643,N_4660,N_4516);
nand U8644 (N_8644,N_3644,N_2237);
nand U8645 (N_8645,N_4918,N_4152);
nor U8646 (N_8646,N_4686,N_163);
nand U8647 (N_8647,N_3879,N_3878);
or U8648 (N_8648,N_3769,N_3488);
and U8649 (N_8649,N_3955,N_4604);
and U8650 (N_8650,N_3,N_397);
or U8651 (N_8651,N_3988,N_706);
nor U8652 (N_8652,N_4070,N_118);
and U8653 (N_8653,N_2046,N_3854);
and U8654 (N_8654,N_3049,N_3106);
nand U8655 (N_8655,N_3423,N_2969);
and U8656 (N_8656,N_4605,N_913);
xnor U8657 (N_8657,N_551,N_3272);
and U8658 (N_8658,N_3444,N_60);
nand U8659 (N_8659,N_4387,N_2997);
nand U8660 (N_8660,N_1081,N_3946);
and U8661 (N_8661,N_263,N_3811);
nor U8662 (N_8662,N_842,N_3242);
and U8663 (N_8663,N_3508,N_3313);
nand U8664 (N_8664,N_1703,N_378);
nand U8665 (N_8665,N_4983,N_2772);
xor U8666 (N_8666,N_3173,N_1510);
and U8667 (N_8667,N_791,N_740);
and U8668 (N_8668,N_4977,N_2895);
or U8669 (N_8669,N_3853,N_2633);
or U8670 (N_8670,N_1023,N_4594);
nor U8671 (N_8671,N_1454,N_431);
nor U8672 (N_8672,N_1003,N_3030);
nor U8673 (N_8673,N_547,N_4627);
and U8674 (N_8674,N_3097,N_1249);
and U8675 (N_8675,N_4820,N_1878);
and U8676 (N_8676,N_4084,N_2518);
or U8677 (N_8677,N_2006,N_1698);
or U8678 (N_8678,N_4533,N_2351);
xor U8679 (N_8679,N_3357,N_3583);
and U8680 (N_8680,N_2775,N_2907);
xnor U8681 (N_8681,N_3451,N_633);
and U8682 (N_8682,N_630,N_3156);
and U8683 (N_8683,N_290,N_660);
nand U8684 (N_8684,N_3184,N_1688);
or U8685 (N_8685,N_1555,N_598);
nand U8686 (N_8686,N_1807,N_1831);
xnor U8687 (N_8687,N_2093,N_2838);
nor U8688 (N_8688,N_563,N_3658);
nor U8689 (N_8689,N_2236,N_4501);
and U8690 (N_8690,N_4043,N_3054);
and U8691 (N_8691,N_3126,N_3918);
and U8692 (N_8692,N_2170,N_3762);
nor U8693 (N_8693,N_1203,N_3455);
and U8694 (N_8694,N_2596,N_1539);
xnor U8695 (N_8695,N_4381,N_247);
nor U8696 (N_8696,N_463,N_3047);
xnor U8697 (N_8697,N_576,N_2420);
and U8698 (N_8698,N_3975,N_852);
and U8699 (N_8699,N_3279,N_260);
xnor U8700 (N_8700,N_879,N_2894);
and U8701 (N_8701,N_2518,N_3954);
or U8702 (N_8702,N_1182,N_3639);
and U8703 (N_8703,N_2170,N_2320);
nand U8704 (N_8704,N_2352,N_3499);
xnor U8705 (N_8705,N_1852,N_4059);
or U8706 (N_8706,N_104,N_2748);
and U8707 (N_8707,N_1160,N_1881);
and U8708 (N_8708,N_3776,N_4459);
or U8709 (N_8709,N_2083,N_3395);
nor U8710 (N_8710,N_2905,N_2383);
or U8711 (N_8711,N_2692,N_2528);
nand U8712 (N_8712,N_1369,N_1194);
and U8713 (N_8713,N_3346,N_3084);
or U8714 (N_8714,N_1644,N_3892);
nand U8715 (N_8715,N_924,N_3518);
or U8716 (N_8716,N_4976,N_3149);
or U8717 (N_8717,N_4880,N_4492);
nor U8718 (N_8718,N_1193,N_4572);
xor U8719 (N_8719,N_3513,N_3575);
nor U8720 (N_8720,N_33,N_2113);
nor U8721 (N_8721,N_4511,N_3257);
nand U8722 (N_8722,N_4935,N_1697);
nor U8723 (N_8723,N_3869,N_2734);
and U8724 (N_8724,N_4776,N_3893);
or U8725 (N_8725,N_3901,N_611);
xnor U8726 (N_8726,N_3151,N_1558);
xnor U8727 (N_8727,N_407,N_1993);
and U8728 (N_8728,N_1330,N_899);
and U8729 (N_8729,N_3606,N_2566);
and U8730 (N_8730,N_2573,N_3852);
nor U8731 (N_8731,N_3533,N_1962);
and U8732 (N_8732,N_3119,N_2960);
nand U8733 (N_8733,N_1865,N_2167);
nand U8734 (N_8734,N_908,N_4021);
nand U8735 (N_8735,N_2359,N_2156);
xor U8736 (N_8736,N_1038,N_194);
nor U8737 (N_8737,N_2937,N_816);
and U8738 (N_8738,N_1990,N_4859);
and U8739 (N_8739,N_3969,N_3127);
nand U8740 (N_8740,N_3565,N_4223);
nor U8741 (N_8741,N_2116,N_2686);
and U8742 (N_8742,N_3131,N_1719);
nand U8743 (N_8743,N_1282,N_521);
or U8744 (N_8744,N_3289,N_4632);
and U8745 (N_8745,N_2725,N_2971);
and U8746 (N_8746,N_3130,N_4578);
nand U8747 (N_8747,N_1601,N_2445);
and U8748 (N_8748,N_1092,N_3309);
xor U8749 (N_8749,N_4276,N_2682);
nor U8750 (N_8750,N_2851,N_2692);
nand U8751 (N_8751,N_471,N_1884);
nand U8752 (N_8752,N_633,N_3031);
nand U8753 (N_8753,N_3722,N_2508);
or U8754 (N_8754,N_2270,N_935);
or U8755 (N_8755,N_1121,N_3266);
nor U8756 (N_8756,N_3181,N_1941);
or U8757 (N_8757,N_2613,N_196);
xor U8758 (N_8758,N_1200,N_4928);
xnor U8759 (N_8759,N_3690,N_1484);
nand U8760 (N_8760,N_2362,N_212);
or U8761 (N_8761,N_1533,N_375);
nand U8762 (N_8762,N_2018,N_1769);
nand U8763 (N_8763,N_2185,N_4954);
nand U8764 (N_8764,N_4290,N_2384);
nor U8765 (N_8765,N_4645,N_1600);
xnor U8766 (N_8766,N_4844,N_818);
nand U8767 (N_8767,N_1803,N_2563);
or U8768 (N_8768,N_1055,N_658);
nand U8769 (N_8769,N_3002,N_2292);
and U8770 (N_8770,N_2935,N_4524);
and U8771 (N_8771,N_3817,N_791);
and U8772 (N_8772,N_3892,N_2420);
nor U8773 (N_8773,N_2787,N_3110);
nor U8774 (N_8774,N_4685,N_2734);
nor U8775 (N_8775,N_3070,N_4140);
or U8776 (N_8776,N_2145,N_4317);
and U8777 (N_8777,N_4601,N_3951);
nor U8778 (N_8778,N_424,N_4899);
or U8779 (N_8779,N_1389,N_1808);
nand U8780 (N_8780,N_589,N_4023);
or U8781 (N_8781,N_2127,N_4735);
or U8782 (N_8782,N_4368,N_2041);
nand U8783 (N_8783,N_2611,N_2941);
or U8784 (N_8784,N_3829,N_1905);
and U8785 (N_8785,N_1438,N_3531);
xnor U8786 (N_8786,N_3,N_4509);
nand U8787 (N_8787,N_2,N_1432);
nor U8788 (N_8788,N_2026,N_2658);
or U8789 (N_8789,N_3752,N_535);
xnor U8790 (N_8790,N_3891,N_4127);
and U8791 (N_8791,N_4778,N_3841);
nand U8792 (N_8792,N_651,N_1215);
or U8793 (N_8793,N_915,N_2980);
nor U8794 (N_8794,N_3736,N_154);
nand U8795 (N_8795,N_1291,N_3085);
or U8796 (N_8796,N_4917,N_4561);
and U8797 (N_8797,N_2214,N_3343);
nor U8798 (N_8798,N_2989,N_1513);
nand U8799 (N_8799,N_1647,N_4628);
nand U8800 (N_8800,N_4519,N_2516);
and U8801 (N_8801,N_4659,N_1371);
and U8802 (N_8802,N_2514,N_4332);
and U8803 (N_8803,N_3012,N_4767);
and U8804 (N_8804,N_2788,N_1355);
nor U8805 (N_8805,N_1367,N_4234);
or U8806 (N_8806,N_3864,N_324);
nor U8807 (N_8807,N_4932,N_4220);
xor U8808 (N_8808,N_121,N_2409);
or U8809 (N_8809,N_3822,N_86);
nand U8810 (N_8810,N_4909,N_3035);
nor U8811 (N_8811,N_2948,N_1226);
nor U8812 (N_8812,N_299,N_718);
nand U8813 (N_8813,N_3719,N_1291);
nor U8814 (N_8814,N_2817,N_410);
nand U8815 (N_8815,N_2294,N_731);
and U8816 (N_8816,N_1200,N_4422);
nand U8817 (N_8817,N_3006,N_4987);
xnor U8818 (N_8818,N_1676,N_2780);
nand U8819 (N_8819,N_2965,N_1401);
and U8820 (N_8820,N_1209,N_3652);
or U8821 (N_8821,N_1825,N_3003);
nor U8822 (N_8822,N_714,N_4477);
or U8823 (N_8823,N_330,N_1551);
nand U8824 (N_8824,N_1860,N_1212);
nor U8825 (N_8825,N_2690,N_3295);
nor U8826 (N_8826,N_2271,N_4845);
and U8827 (N_8827,N_3344,N_1129);
nand U8828 (N_8828,N_3299,N_23);
nor U8829 (N_8829,N_516,N_867);
nor U8830 (N_8830,N_3726,N_4198);
xnor U8831 (N_8831,N_342,N_2783);
or U8832 (N_8832,N_1639,N_2229);
and U8833 (N_8833,N_2292,N_3267);
nor U8834 (N_8834,N_3773,N_3817);
and U8835 (N_8835,N_3499,N_516);
or U8836 (N_8836,N_2253,N_298);
nand U8837 (N_8837,N_1526,N_3511);
nand U8838 (N_8838,N_521,N_4254);
and U8839 (N_8839,N_2844,N_4214);
or U8840 (N_8840,N_3984,N_3382);
or U8841 (N_8841,N_3280,N_3479);
and U8842 (N_8842,N_4367,N_2487);
and U8843 (N_8843,N_2063,N_2064);
nor U8844 (N_8844,N_3485,N_249);
nand U8845 (N_8845,N_4237,N_4499);
and U8846 (N_8846,N_4824,N_731);
nand U8847 (N_8847,N_133,N_95);
nand U8848 (N_8848,N_1959,N_3784);
xor U8849 (N_8849,N_1055,N_2759);
and U8850 (N_8850,N_3440,N_4786);
nand U8851 (N_8851,N_4011,N_2626);
nor U8852 (N_8852,N_3558,N_3742);
nor U8853 (N_8853,N_4598,N_2549);
or U8854 (N_8854,N_4538,N_352);
xnor U8855 (N_8855,N_1215,N_2436);
nor U8856 (N_8856,N_869,N_1576);
or U8857 (N_8857,N_545,N_2659);
or U8858 (N_8858,N_2448,N_1311);
and U8859 (N_8859,N_4127,N_4831);
xor U8860 (N_8860,N_1527,N_2730);
or U8861 (N_8861,N_1253,N_4031);
nand U8862 (N_8862,N_1788,N_1400);
nor U8863 (N_8863,N_125,N_374);
nand U8864 (N_8864,N_4769,N_970);
or U8865 (N_8865,N_3725,N_1355);
and U8866 (N_8866,N_3629,N_1866);
nand U8867 (N_8867,N_223,N_145);
nor U8868 (N_8868,N_1167,N_1317);
or U8869 (N_8869,N_3735,N_1531);
xor U8870 (N_8870,N_3502,N_2618);
nand U8871 (N_8871,N_3693,N_2771);
or U8872 (N_8872,N_1388,N_1659);
nand U8873 (N_8873,N_813,N_2864);
and U8874 (N_8874,N_1446,N_1068);
nor U8875 (N_8875,N_4560,N_4139);
and U8876 (N_8876,N_771,N_1956);
or U8877 (N_8877,N_1038,N_1054);
nand U8878 (N_8878,N_791,N_4566);
and U8879 (N_8879,N_1247,N_4262);
or U8880 (N_8880,N_1416,N_1834);
nand U8881 (N_8881,N_1239,N_4604);
nand U8882 (N_8882,N_4974,N_1841);
nor U8883 (N_8883,N_1535,N_3194);
or U8884 (N_8884,N_4947,N_3495);
and U8885 (N_8885,N_92,N_3167);
and U8886 (N_8886,N_573,N_1449);
and U8887 (N_8887,N_4460,N_429);
and U8888 (N_8888,N_4552,N_1436);
and U8889 (N_8889,N_285,N_2010);
or U8890 (N_8890,N_734,N_1619);
or U8891 (N_8891,N_4964,N_1561);
nand U8892 (N_8892,N_3340,N_2407);
and U8893 (N_8893,N_813,N_298);
nand U8894 (N_8894,N_1552,N_2496);
and U8895 (N_8895,N_2752,N_3749);
and U8896 (N_8896,N_514,N_2607);
nand U8897 (N_8897,N_869,N_2736);
nor U8898 (N_8898,N_1122,N_1966);
and U8899 (N_8899,N_778,N_2340);
or U8900 (N_8900,N_2966,N_2012);
or U8901 (N_8901,N_2792,N_33);
and U8902 (N_8902,N_786,N_1663);
or U8903 (N_8903,N_4768,N_8);
nor U8904 (N_8904,N_3363,N_3358);
or U8905 (N_8905,N_4337,N_2832);
nand U8906 (N_8906,N_3348,N_586);
nor U8907 (N_8907,N_1601,N_2018);
xor U8908 (N_8908,N_1683,N_4700);
nand U8909 (N_8909,N_871,N_599);
nor U8910 (N_8910,N_3320,N_64);
nor U8911 (N_8911,N_1972,N_1061);
nand U8912 (N_8912,N_3738,N_4727);
and U8913 (N_8913,N_526,N_670);
and U8914 (N_8914,N_2432,N_1403);
or U8915 (N_8915,N_2940,N_1909);
and U8916 (N_8916,N_73,N_1068);
and U8917 (N_8917,N_1602,N_4554);
nand U8918 (N_8918,N_2070,N_1311);
nor U8919 (N_8919,N_3296,N_971);
nand U8920 (N_8920,N_349,N_645);
nand U8921 (N_8921,N_2391,N_4384);
or U8922 (N_8922,N_4709,N_4768);
or U8923 (N_8923,N_4025,N_2454);
nor U8924 (N_8924,N_2283,N_3672);
and U8925 (N_8925,N_4513,N_955);
nand U8926 (N_8926,N_220,N_1245);
or U8927 (N_8927,N_4061,N_3398);
or U8928 (N_8928,N_3257,N_1830);
xor U8929 (N_8929,N_398,N_3492);
xnor U8930 (N_8930,N_3141,N_1741);
and U8931 (N_8931,N_2627,N_1321);
nor U8932 (N_8932,N_3090,N_4782);
or U8933 (N_8933,N_4967,N_2278);
nor U8934 (N_8934,N_52,N_2965);
nor U8935 (N_8935,N_3330,N_2781);
or U8936 (N_8936,N_1387,N_1336);
or U8937 (N_8937,N_1370,N_2013);
nor U8938 (N_8938,N_2094,N_4230);
nor U8939 (N_8939,N_1506,N_3525);
or U8940 (N_8940,N_4615,N_3347);
and U8941 (N_8941,N_2685,N_3330);
nand U8942 (N_8942,N_253,N_2529);
and U8943 (N_8943,N_2512,N_1367);
nor U8944 (N_8944,N_1275,N_53);
nor U8945 (N_8945,N_2753,N_723);
and U8946 (N_8946,N_2669,N_3761);
nand U8947 (N_8947,N_4241,N_1903);
or U8948 (N_8948,N_4394,N_442);
xnor U8949 (N_8949,N_1829,N_3351);
or U8950 (N_8950,N_4988,N_3268);
or U8951 (N_8951,N_1087,N_4427);
and U8952 (N_8952,N_2926,N_1265);
or U8953 (N_8953,N_849,N_4113);
or U8954 (N_8954,N_2620,N_267);
nor U8955 (N_8955,N_2967,N_2878);
and U8956 (N_8956,N_3635,N_3589);
and U8957 (N_8957,N_386,N_124);
nand U8958 (N_8958,N_2490,N_4380);
xor U8959 (N_8959,N_2968,N_551);
xor U8960 (N_8960,N_4814,N_1478);
and U8961 (N_8961,N_2880,N_4731);
nor U8962 (N_8962,N_4812,N_442);
nand U8963 (N_8963,N_3274,N_3407);
xor U8964 (N_8964,N_2201,N_4626);
nand U8965 (N_8965,N_3805,N_567);
and U8966 (N_8966,N_4958,N_3291);
nor U8967 (N_8967,N_1158,N_4065);
or U8968 (N_8968,N_1426,N_3019);
xnor U8969 (N_8969,N_679,N_2975);
nand U8970 (N_8970,N_1207,N_4179);
and U8971 (N_8971,N_1920,N_227);
and U8972 (N_8972,N_3564,N_4069);
and U8973 (N_8973,N_940,N_4442);
or U8974 (N_8974,N_1267,N_4988);
nor U8975 (N_8975,N_3978,N_2782);
nand U8976 (N_8976,N_3249,N_3881);
and U8977 (N_8977,N_2552,N_3510);
nand U8978 (N_8978,N_4806,N_3011);
nor U8979 (N_8979,N_918,N_1579);
xnor U8980 (N_8980,N_585,N_2132);
nor U8981 (N_8981,N_271,N_690);
and U8982 (N_8982,N_4376,N_4637);
nor U8983 (N_8983,N_643,N_403);
nor U8984 (N_8984,N_2191,N_4714);
or U8985 (N_8985,N_3872,N_4580);
or U8986 (N_8986,N_1818,N_689);
nor U8987 (N_8987,N_3788,N_1269);
nand U8988 (N_8988,N_271,N_646);
nand U8989 (N_8989,N_1744,N_1420);
nor U8990 (N_8990,N_4177,N_4781);
nand U8991 (N_8991,N_2118,N_3231);
or U8992 (N_8992,N_204,N_2108);
and U8993 (N_8993,N_3002,N_2877);
nor U8994 (N_8994,N_2460,N_4698);
or U8995 (N_8995,N_586,N_3609);
and U8996 (N_8996,N_1448,N_989);
nand U8997 (N_8997,N_4494,N_3704);
or U8998 (N_8998,N_1945,N_2320);
nand U8999 (N_8999,N_4968,N_1822);
nand U9000 (N_9000,N_4132,N_3423);
nand U9001 (N_9001,N_2973,N_993);
nand U9002 (N_9002,N_2431,N_3698);
nor U9003 (N_9003,N_2715,N_4636);
nand U9004 (N_9004,N_612,N_1373);
nand U9005 (N_9005,N_1036,N_1153);
and U9006 (N_9006,N_1017,N_678);
nor U9007 (N_9007,N_3372,N_701);
and U9008 (N_9008,N_1616,N_1760);
nand U9009 (N_9009,N_1876,N_2377);
nor U9010 (N_9010,N_2802,N_2179);
nor U9011 (N_9011,N_4802,N_2464);
or U9012 (N_9012,N_4079,N_3518);
nand U9013 (N_9013,N_2897,N_1291);
or U9014 (N_9014,N_3667,N_1300);
or U9015 (N_9015,N_3172,N_1335);
or U9016 (N_9016,N_1332,N_1526);
nand U9017 (N_9017,N_3106,N_2460);
and U9018 (N_9018,N_2246,N_3289);
and U9019 (N_9019,N_4499,N_3509);
nand U9020 (N_9020,N_4247,N_4766);
and U9021 (N_9021,N_1052,N_4081);
nor U9022 (N_9022,N_4333,N_3761);
nor U9023 (N_9023,N_3965,N_2354);
nor U9024 (N_9024,N_1106,N_963);
or U9025 (N_9025,N_1529,N_4472);
and U9026 (N_9026,N_4287,N_734);
or U9027 (N_9027,N_4308,N_804);
nor U9028 (N_9028,N_4357,N_2607);
nor U9029 (N_9029,N_4643,N_3288);
and U9030 (N_9030,N_4724,N_2754);
and U9031 (N_9031,N_2768,N_1061);
nand U9032 (N_9032,N_392,N_3315);
or U9033 (N_9033,N_4914,N_1123);
nor U9034 (N_9034,N_4652,N_2096);
nand U9035 (N_9035,N_4852,N_3481);
nor U9036 (N_9036,N_2423,N_334);
nor U9037 (N_9037,N_4368,N_2936);
and U9038 (N_9038,N_4738,N_3404);
nor U9039 (N_9039,N_439,N_786);
nor U9040 (N_9040,N_3720,N_2545);
and U9041 (N_9041,N_1179,N_3245);
nand U9042 (N_9042,N_37,N_4750);
nand U9043 (N_9043,N_2795,N_1295);
or U9044 (N_9044,N_1302,N_4033);
nand U9045 (N_9045,N_353,N_2852);
or U9046 (N_9046,N_3929,N_2192);
and U9047 (N_9047,N_749,N_1268);
or U9048 (N_9048,N_2636,N_4607);
nor U9049 (N_9049,N_12,N_2801);
nor U9050 (N_9050,N_4746,N_2192);
nor U9051 (N_9051,N_98,N_3676);
nand U9052 (N_9052,N_3089,N_4417);
and U9053 (N_9053,N_2498,N_728);
nor U9054 (N_9054,N_4356,N_4277);
and U9055 (N_9055,N_513,N_431);
nor U9056 (N_9056,N_43,N_4349);
and U9057 (N_9057,N_1249,N_2241);
nand U9058 (N_9058,N_168,N_4476);
or U9059 (N_9059,N_547,N_112);
or U9060 (N_9060,N_4544,N_1176);
nand U9061 (N_9061,N_860,N_4660);
nor U9062 (N_9062,N_4923,N_2134);
and U9063 (N_9063,N_1986,N_751);
and U9064 (N_9064,N_319,N_2163);
xor U9065 (N_9065,N_932,N_3729);
and U9066 (N_9066,N_2722,N_1134);
nor U9067 (N_9067,N_50,N_1378);
and U9068 (N_9068,N_823,N_4715);
and U9069 (N_9069,N_2121,N_4623);
xnor U9070 (N_9070,N_4631,N_1804);
or U9071 (N_9071,N_581,N_1161);
nor U9072 (N_9072,N_167,N_1447);
nor U9073 (N_9073,N_2715,N_2671);
nor U9074 (N_9074,N_918,N_272);
nand U9075 (N_9075,N_1284,N_1745);
or U9076 (N_9076,N_2358,N_4420);
xnor U9077 (N_9077,N_3369,N_4470);
or U9078 (N_9078,N_4952,N_50);
and U9079 (N_9079,N_2324,N_4553);
and U9080 (N_9080,N_2426,N_258);
or U9081 (N_9081,N_314,N_4728);
or U9082 (N_9082,N_3460,N_512);
and U9083 (N_9083,N_2508,N_1760);
nor U9084 (N_9084,N_171,N_4926);
and U9085 (N_9085,N_2780,N_3448);
nor U9086 (N_9086,N_2515,N_4628);
nand U9087 (N_9087,N_4725,N_4024);
and U9088 (N_9088,N_1822,N_13);
nand U9089 (N_9089,N_1419,N_373);
nor U9090 (N_9090,N_2232,N_2538);
nand U9091 (N_9091,N_3074,N_4290);
xor U9092 (N_9092,N_945,N_2984);
or U9093 (N_9093,N_4249,N_4822);
nor U9094 (N_9094,N_658,N_1349);
nand U9095 (N_9095,N_4082,N_3911);
nand U9096 (N_9096,N_721,N_4319);
or U9097 (N_9097,N_2013,N_1976);
xnor U9098 (N_9098,N_762,N_311);
nor U9099 (N_9099,N_3652,N_3604);
or U9100 (N_9100,N_3358,N_2070);
and U9101 (N_9101,N_2786,N_1523);
xor U9102 (N_9102,N_4132,N_1762);
or U9103 (N_9103,N_4044,N_4503);
nor U9104 (N_9104,N_4760,N_3564);
and U9105 (N_9105,N_4474,N_3148);
nand U9106 (N_9106,N_4027,N_4015);
and U9107 (N_9107,N_4,N_1329);
nand U9108 (N_9108,N_109,N_4538);
or U9109 (N_9109,N_3851,N_4660);
nand U9110 (N_9110,N_3437,N_3612);
nor U9111 (N_9111,N_1694,N_837);
nor U9112 (N_9112,N_1222,N_1968);
xor U9113 (N_9113,N_3304,N_3994);
or U9114 (N_9114,N_3606,N_2307);
nand U9115 (N_9115,N_340,N_4348);
and U9116 (N_9116,N_2236,N_2422);
or U9117 (N_9117,N_2428,N_2970);
nand U9118 (N_9118,N_4297,N_386);
nand U9119 (N_9119,N_4528,N_1785);
or U9120 (N_9120,N_1759,N_28);
nor U9121 (N_9121,N_246,N_537);
nor U9122 (N_9122,N_2355,N_3893);
and U9123 (N_9123,N_3059,N_4008);
xnor U9124 (N_9124,N_3532,N_1856);
and U9125 (N_9125,N_3478,N_2837);
or U9126 (N_9126,N_2991,N_1267);
nand U9127 (N_9127,N_4631,N_1791);
nor U9128 (N_9128,N_934,N_226);
or U9129 (N_9129,N_2963,N_1);
xnor U9130 (N_9130,N_4491,N_4060);
xor U9131 (N_9131,N_3443,N_1773);
nand U9132 (N_9132,N_1171,N_2732);
or U9133 (N_9133,N_340,N_3248);
or U9134 (N_9134,N_1459,N_4500);
nor U9135 (N_9135,N_3977,N_2425);
or U9136 (N_9136,N_1875,N_3554);
or U9137 (N_9137,N_4975,N_2035);
nand U9138 (N_9138,N_2597,N_2251);
or U9139 (N_9139,N_1253,N_4937);
nor U9140 (N_9140,N_4038,N_263);
xnor U9141 (N_9141,N_1764,N_1155);
nor U9142 (N_9142,N_250,N_4506);
or U9143 (N_9143,N_1473,N_4875);
nand U9144 (N_9144,N_118,N_4383);
nand U9145 (N_9145,N_285,N_884);
nor U9146 (N_9146,N_1220,N_4558);
nor U9147 (N_9147,N_2063,N_2486);
and U9148 (N_9148,N_1525,N_4403);
nand U9149 (N_9149,N_3013,N_2770);
nor U9150 (N_9150,N_1914,N_3684);
and U9151 (N_9151,N_416,N_1310);
nand U9152 (N_9152,N_3877,N_3451);
and U9153 (N_9153,N_2485,N_1722);
nand U9154 (N_9154,N_4476,N_2020);
or U9155 (N_9155,N_3868,N_3556);
nand U9156 (N_9156,N_4975,N_1302);
and U9157 (N_9157,N_2884,N_2358);
nor U9158 (N_9158,N_4167,N_4627);
nand U9159 (N_9159,N_2106,N_4664);
xor U9160 (N_9160,N_4066,N_146);
nor U9161 (N_9161,N_2305,N_4645);
or U9162 (N_9162,N_1895,N_3181);
nand U9163 (N_9163,N_3575,N_2908);
or U9164 (N_9164,N_2161,N_3597);
nand U9165 (N_9165,N_2442,N_1710);
nand U9166 (N_9166,N_2951,N_2731);
nand U9167 (N_9167,N_2880,N_4459);
or U9168 (N_9168,N_584,N_2116);
nor U9169 (N_9169,N_3950,N_98);
nor U9170 (N_9170,N_4399,N_3622);
xor U9171 (N_9171,N_2514,N_334);
nor U9172 (N_9172,N_2835,N_286);
and U9173 (N_9173,N_1638,N_124);
and U9174 (N_9174,N_38,N_4844);
nand U9175 (N_9175,N_4387,N_4943);
or U9176 (N_9176,N_2426,N_2086);
nand U9177 (N_9177,N_4652,N_268);
and U9178 (N_9178,N_4123,N_2266);
and U9179 (N_9179,N_4996,N_1229);
xor U9180 (N_9180,N_489,N_3653);
and U9181 (N_9181,N_3143,N_479);
nor U9182 (N_9182,N_3180,N_764);
and U9183 (N_9183,N_2254,N_2018);
or U9184 (N_9184,N_4270,N_1092);
nand U9185 (N_9185,N_3035,N_3440);
and U9186 (N_9186,N_3388,N_614);
xor U9187 (N_9187,N_2719,N_2527);
and U9188 (N_9188,N_2958,N_1);
xnor U9189 (N_9189,N_1977,N_4051);
nor U9190 (N_9190,N_2479,N_1649);
and U9191 (N_9191,N_4323,N_4611);
nor U9192 (N_9192,N_884,N_454);
xor U9193 (N_9193,N_4819,N_3522);
nor U9194 (N_9194,N_1816,N_1465);
nor U9195 (N_9195,N_413,N_2043);
or U9196 (N_9196,N_4496,N_2535);
nand U9197 (N_9197,N_3915,N_634);
nor U9198 (N_9198,N_1727,N_551);
xnor U9199 (N_9199,N_1223,N_619);
xor U9200 (N_9200,N_361,N_202);
or U9201 (N_9201,N_3738,N_4874);
or U9202 (N_9202,N_2525,N_4300);
nand U9203 (N_9203,N_266,N_1123);
nor U9204 (N_9204,N_3295,N_1384);
or U9205 (N_9205,N_2497,N_740);
nand U9206 (N_9206,N_830,N_4335);
and U9207 (N_9207,N_1431,N_4068);
nor U9208 (N_9208,N_1364,N_569);
and U9209 (N_9209,N_3532,N_4430);
nand U9210 (N_9210,N_4761,N_4471);
nor U9211 (N_9211,N_880,N_3904);
or U9212 (N_9212,N_3672,N_4403);
and U9213 (N_9213,N_1485,N_375);
nand U9214 (N_9214,N_2351,N_4276);
nor U9215 (N_9215,N_3199,N_3484);
nand U9216 (N_9216,N_740,N_4502);
or U9217 (N_9217,N_478,N_1619);
nor U9218 (N_9218,N_1863,N_4389);
xor U9219 (N_9219,N_3477,N_3097);
and U9220 (N_9220,N_143,N_2006);
or U9221 (N_9221,N_4236,N_1712);
and U9222 (N_9222,N_1508,N_3799);
xnor U9223 (N_9223,N_568,N_1790);
or U9224 (N_9224,N_3522,N_3240);
and U9225 (N_9225,N_1552,N_1966);
nor U9226 (N_9226,N_988,N_3344);
nand U9227 (N_9227,N_3095,N_1271);
or U9228 (N_9228,N_1445,N_3773);
and U9229 (N_9229,N_822,N_3975);
or U9230 (N_9230,N_412,N_2398);
or U9231 (N_9231,N_4791,N_2170);
nor U9232 (N_9232,N_4255,N_686);
nand U9233 (N_9233,N_3040,N_424);
or U9234 (N_9234,N_4242,N_4672);
nand U9235 (N_9235,N_1629,N_2138);
and U9236 (N_9236,N_1510,N_88);
or U9237 (N_9237,N_1377,N_1780);
nand U9238 (N_9238,N_1501,N_4876);
xnor U9239 (N_9239,N_1922,N_2779);
or U9240 (N_9240,N_3994,N_307);
or U9241 (N_9241,N_975,N_2981);
and U9242 (N_9242,N_3549,N_4776);
or U9243 (N_9243,N_2826,N_2524);
nand U9244 (N_9244,N_2857,N_2134);
or U9245 (N_9245,N_218,N_4761);
and U9246 (N_9246,N_1543,N_449);
nand U9247 (N_9247,N_1967,N_2192);
xor U9248 (N_9248,N_4462,N_4673);
nand U9249 (N_9249,N_3984,N_3483);
and U9250 (N_9250,N_4439,N_3097);
nand U9251 (N_9251,N_1076,N_470);
and U9252 (N_9252,N_4454,N_280);
or U9253 (N_9253,N_2562,N_1858);
and U9254 (N_9254,N_1877,N_1318);
or U9255 (N_9255,N_871,N_294);
or U9256 (N_9256,N_3965,N_1540);
nor U9257 (N_9257,N_2902,N_1493);
nand U9258 (N_9258,N_3215,N_799);
and U9259 (N_9259,N_2619,N_4098);
or U9260 (N_9260,N_975,N_3013);
nand U9261 (N_9261,N_1454,N_4418);
nor U9262 (N_9262,N_3714,N_3213);
or U9263 (N_9263,N_4704,N_1554);
or U9264 (N_9264,N_954,N_3528);
and U9265 (N_9265,N_4694,N_1660);
or U9266 (N_9266,N_1300,N_914);
nor U9267 (N_9267,N_2347,N_3456);
and U9268 (N_9268,N_4941,N_2939);
xnor U9269 (N_9269,N_4775,N_2829);
nand U9270 (N_9270,N_3203,N_4812);
and U9271 (N_9271,N_2520,N_2139);
or U9272 (N_9272,N_1248,N_2646);
xnor U9273 (N_9273,N_4391,N_3627);
nor U9274 (N_9274,N_1476,N_3288);
nand U9275 (N_9275,N_1300,N_3709);
or U9276 (N_9276,N_3834,N_4393);
and U9277 (N_9277,N_297,N_3695);
and U9278 (N_9278,N_3360,N_894);
nand U9279 (N_9279,N_3616,N_4481);
nor U9280 (N_9280,N_1229,N_367);
and U9281 (N_9281,N_2016,N_4067);
nor U9282 (N_9282,N_2509,N_4429);
and U9283 (N_9283,N_514,N_3431);
or U9284 (N_9284,N_3887,N_1184);
or U9285 (N_9285,N_2134,N_2899);
xor U9286 (N_9286,N_2503,N_2317);
or U9287 (N_9287,N_4082,N_1927);
nor U9288 (N_9288,N_2364,N_241);
and U9289 (N_9289,N_1100,N_3916);
nor U9290 (N_9290,N_1674,N_4943);
or U9291 (N_9291,N_3998,N_4181);
or U9292 (N_9292,N_3977,N_1210);
nand U9293 (N_9293,N_1615,N_2757);
nor U9294 (N_9294,N_702,N_3068);
nand U9295 (N_9295,N_1919,N_3201);
nor U9296 (N_9296,N_4208,N_2360);
or U9297 (N_9297,N_1336,N_3108);
or U9298 (N_9298,N_17,N_1636);
nand U9299 (N_9299,N_2763,N_2561);
and U9300 (N_9300,N_4026,N_1391);
xor U9301 (N_9301,N_2120,N_1640);
or U9302 (N_9302,N_2746,N_1042);
nor U9303 (N_9303,N_4678,N_1752);
and U9304 (N_9304,N_327,N_2452);
xor U9305 (N_9305,N_4296,N_1764);
or U9306 (N_9306,N_4597,N_2586);
or U9307 (N_9307,N_4165,N_1786);
nor U9308 (N_9308,N_1803,N_1075);
and U9309 (N_9309,N_4728,N_4754);
nor U9310 (N_9310,N_3216,N_3924);
nand U9311 (N_9311,N_4292,N_1024);
and U9312 (N_9312,N_319,N_786);
nor U9313 (N_9313,N_1329,N_176);
and U9314 (N_9314,N_3520,N_2346);
nand U9315 (N_9315,N_126,N_2422);
xnor U9316 (N_9316,N_3029,N_4311);
and U9317 (N_9317,N_2682,N_3524);
xor U9318 (N_9318,N_293,N_2407);
nand U9319 (N_9319,N_3143,N_1845);
nand U9320 (N_9320,N_4276,N_3420);
nand U9321 (N_9321,N_84,N_1049);
and U9322 (N_9322,N_240,N_2583);
or U9323 (N_9323,N_324,N_2358);
and U9324 (N_9324,N_636,N_2103);
xnor U9325 (N_9325,N_398,N_3078);
and U9326 (N_9326,N_2258,N_2455);
and U9327 (N_9327,N_2309,N_4848);
or U9328 (N_9328,N_3686,N_1327);
or U9329 (N_9329,N_4467,N_3768);
nand U9330 (N_9330,N_4258,N_3784);
or U9331 (N_9331,N_4143,N_1254);
nand U9332 (N_9332,N_652,N_2661);
nor U9333 (N_9333,N_3753,N_2707);
and U9334 (N_9334,N_1977,N_987);
nor U9335 (N_9335,N_2139,N_651);
nor U9336 (N_9336,N_491,N_3329);
xnor U9337 (N_9337,N_4967,N_4484);
nor U9338 (N_9338,N_2015,N_2461);
or U9339 (N_9339,N_29,N_4277);
or U9340 (N_9340,N_2258,N_3551);
and U9341 (N_9341,N_4456,N_4266);
and U9342 (N_9342,N_796,N_1219);
nor U9343 (N_9343,N_1843,N_3645);
nor U9344 (N_9344,N_1074,N_558);
or U9345 (N_9345,N_3843,N_616);
or U9346 (N_9346,N_4980,N_1266);
xor U9347 (N_9347,N_3986,N_3129);
and U9348 (N_9348,N_1662,N_192);
nor U9349 (N_9349,N_4868,N_731);
xnor U9350 (N_9350,N_4730,N_4264);
nor U9351 (N_9351,N_1727,N_400);
and U9352 (N_9352,N_629,N_546);
or U9353 (N_9353,N_1310,N_1363);
xnor U9354 (N_9354,N_4904,N_1111);
nor U9355 (N_9355,N_1855,N_3078);
or U9356 (N_9356,N_2843,N_3173);
nor U9357 (N_9357,N_2343,N_625);
nor U9358 (N_9358,N_4643,N_1123);
nand U9359 (N_9359,N_1532,N_867);
xnor U9360 (N_9360,N_1645,N_3512);
and U9361 (N_9361,N_4530,N_2783);
or U9362 (N_9362,N_239,N_1483);
xnor U9363 (N_9363,N_2799,N_9);
nand U9364 (N_9364,N_3177,N_1156);
or U9365 (N_9365,N_3441,N_3153);
or U9366 (N_9366,N_3142,N_958);
nand U9367 (N_9367,N_3805,N_262);
nor U9368 (N_9368,N_2760,N_179);
or U9369 (N_9369,N_3921,N_4248);
nor U9370 (N_9370,N_4238,N_1942);
and U9371 (N_9371,N_95,N_2575);
nor U9372 (N_9372,N_2267,N_4664);
and U9373 (N_9373,N_1430,N_787);
or U9374 (N_9374,N_4824,N_4835);
or U9375 (N_9375,N_477,N_1660);
nor U9376 (N_9376,N_4,N_1240);
or U9377 (N_9377,N_33,N_892);
or U9378 (N_9378,N_1583,N_2950);
nor U9379 (N_9379,N_2743,N_72);
nor U9380 (N_9380,N_683,N_2269);
nand U9381 (N_9381,N_1602,N_2465);
or U9382 (N_9382,N_2946,N_136);
and U9383 (N_9383,N_4661,N_4547);
and U9384 (N_9384,N_1011,N_3201);
or U9385 (N_9385,N_804,N_4079);
or U9386 (N_9386,N_306,N_4558);
and U9387 (N_9387,N_4994,N_3716);
nand U9388 (N_9388,N_4399,N_678);
xor U9389 (N_9389,N_1665,N_908);
nor U9390 (N_9390,N_4726,N_236);
nand U9391 (N_9391,N_3237,N_4171);
or U9392 (N_9392,N_3573,N_973);
nand U9393 (N_9393,N_200,N_2456);
nor U9394 (N_9394,N_299,N_156);
and U9395 (N_9395,N_3298,N_898);
nand U9396 (N_9396,N_2294,N_304);
nor U9397 (N_9397,N_2104,N_831);
and U9398 (N_9398,N_3248,N_1331);
nor U9399 (N_9399,N_2952,N_2074);
or U9400 (N_9400,N_2692,N_541);
nand U9401 (N_9401,N_2261,N_2152);
nor U9402 (N_9402,N_3802,N_3772);
and U9403 (N_9403,N_1596,N_2031);
nor U9404 (N_9404,N_4893,N_4237);
and U9405 (N_9405,N_2532,N_2772);
or U9406 (N_9406,N_4978,N_2335);
nor U9407 (N_9407,N_20,N_3944);
and U9408 (N_9408,N_9,N_293);
nor U9409 (N_9409,N_429,N_3794);
and U9410 (N_9410,N_1609,N_939);
and U9411 (N_9411,N_4700,N_3924);
nor U9412 (N_9412,N_2451,N_2059);
or U9413 (N_9413,N_4720,N_2800);
nand U9414 (N_9414,N_1002,N_929);
nand U9415 (N_9415,N_4463,N_3665);
or U9416 (N_9416,N_4246,N_4315);
nor U9417 (N_9417,N_3975,N_100);
xnor U9418 (N_9418,N_4432,N_224);
nand U9419 (N_9419,N_2755,N_4880);
xor U9420 (N_9420,N_488,N_4025);
xor U9421 (N_9421,N_1972,N_4459);
nor U9422 (N_9422,N_56,N_308);
xnor U9423 (N_9423,N_651,N_4021);
nor U9424 (N_9424,N_4187,N_1434);
or U9425 (N_9425,N_3596,N_772);
nor U9426 (N_9426,N_2022,N_3185);
or U9427 (N_9427,N_2645,N_3345);
nand U9428 (N_9428,N_2780,N_2200);
xor U9429 (N_9429,N_453,N_586);
nand U9430 (N_9430,N_3189,N_269);
and U9431 (N_9431,N_3398,N_2621);
nor U9432 (N_9432,N_2329,N_121);
xor U9433 (N_9433,N_3316,N_4536);
or U9434 (N_9434,N_3949,N_3370);
nor U9435 (N_9435,N_731,N_4508);
and U9436 (N_9436,N_3550,N_1785);
or U9437 (N_9437,N_686,N_3565);
and U9438 (N_9438,N_4440,N_2272);
nand U9439 (N_9439,N_1330,N_4322);
nand U9440 (N_9440,N_802,N_104);
or U9441 (N_9441,N_126,N_2521);
nor U9442 (N_9442,N_1708,N_1577);
or U9443 (N_9443,N_50,N_2207);
nand U9444 (N_9444,N_325,N_202);
nor U9445 (N_9445,N_4623,N_602);
nor U9446 (N_9446,N_2527,N_4222);
or U9447 (N_9447,N_1077,N_539);
nand U9448 (N_9448,N_4349,N_761);
or U9449 (N_9449,N_3172,N_353);
nor U9450 (N_9450,N_1956,N_1280);
nand U9451 (N_9451,N_4766,N_2826);
nand U9452 (N_9452,N_1681,N_3858);
xor U9453 (N_9453,N_596,N_3513);
and U9454 (N_9454,N_2760,N_2682);
and U9455 (N_9455,N_4604,N_2301);
and U9456 (N_9456,N_3146,N_684);
nor U9457 (N_9457,N_766,N_588);
or U9458 (N_9458,N_4139,N_4466);
or U9459 (N_9459,N_2475,N_4554);
or U9460 (N_9460,N_922,N_166);
nand U9461 (N_9461,N_2439,N_2);
and U9462 (N_9462,N_2058,N_857);
nand U9463 (N_9463,N_3480,N_1388);
or U9464 (N_9464,N_3418,N_3672);
nand U9465 (N_9465,N_1558,N_4289);
and U9466 (N_9466,N_1555,N_2788);
or U9467 (N_9467,N_629,N_724);
nor U9468 (N_9468,N_1116,N_4098);
xnor U9469 (N_9469,N_2202,N_488);
and U9470 (N_9470,N_1347,N_4611);
nand U9471 (N_9471,N_768,N_3744);
or U9472 (N_9472,N_4221,N_3626);
nor U9473 (N_9473,N_2803,N_3803);
and U9474 (N_9474,N_4464,N_4230);
or U9475 (N_9475,N_2788,N_2991);
nor U9476 (N_9476,N_2068,N_3111);
nor U9477 (N_9477,N_2116,N_3620);
and U9478 (N_9478,N_4204,N_864);
or U9479 (N_9479,N_437,N_3991);
or U9480 (N_9480,N_2654,N_1866);
and U9481 (N_9481,N_2637,N_1576);
nor U9482 (N_9482,N_4413,N_4531);
or U9483 (N_9483,N_1527,N_1437);
and U9484 (N_9484,N_198,N_4805);
nand U9485 (N_9485,N_2306,N_3243);
or U9486 (N_9486,N_1057,N_1588);
nor U9487 (N_9487,N_3168,N_2521);
nor U9488 (N_9488,N_4859,N_3318);
xnor U9489 (N_9489,N_315,N_1103);
or U9490 (N_9490,N_1540,N_1304);
nand U9491 (N_9491,N_4930,N_2175);
nor U9492 (N_9492,N_4650,N_3784);
xor U9493 (N_9493,N_3969,N_4463);
nand U9494 (N_9494,N_4317,N_393);
nor U9495 (N_9495,N_4626,N_3416);
or U9496 (N_9496,N_2915,N_96);
or U9497 (N_9497,N_3889,N_1160);
nand U9498 (N_9498,N_2690,N_2254);
nor U9499 (N_9499,N_4758,N_2332);
or U9500 (N_9500,N_3013,N_2579);
or U9501 (N_9501,N_3583,N_1986);
and U9502 (N_9502,N_4087,N_3436);
or U9503 (N_9503,N_2621,N_2177);
and U9504 (N_9504,N_4575,N_2345);
xor U9505 (N_9505,N_1617,N_621);
nor U9506 (N_9506,N_1809,N_74);
and U9507 (N_9507,N_4923,N_3647);
and U9508 (N_9508,N_173,N_4104);
or U9509 (N_9509,N_3176,N_3822);
nand U9510 (N_9510,N_1955,N_3411);
and U9511 (N_9511,N_630,N_2015);
nor U9512 (N_9512,N_982,N_530);
or U9513 (N_9513,N_994,N_2520);
nand U9514 (N_9514,N_3457,N_2207);
xor U9515 (N_9515,N_3519,N_250);
nand U9516 (N_9516,N_753,N_3472);
and U9517 (N_9517,N_982,N_4192);
or U9518 (N_9518,N_1796,N_1244);
xor U9519 (N_9519,N_1120,N_1811);
and U9520 (N_9520,N_985,N_162);
and U9521 (N_9521,N_4639,N_1064);
nand U9522 (N_9522,N_916,N_2539);
xor U9523 (N_9523,N_3608,N_2340);
and U9524 (N_9524,N_3929,N_632);
nand U9525 (N_9525,N_4971,N_715);
nand U9526 (N_9526,N_395,N_1054);
nand U9527 (N_9527,N_3252,N_2807);
and U9528 (N_9528,N_1325,N_4189);
nand U9529 (N_9529,N_2412,N_4980);
or U9530 (N_9530,N_4654,N_4008);
nand U9531 (N_9531,N_2675,N_2359);
and U9532 (N_9532,N_2730,N_3102);
and U9533 (N_9533,N_2092,N_4348);
and U9534 (N_9534,N_4238,N_3898);
nand U9535 (N_9535,N_963,N_2968);
nor U9536 (N_9536,N_1597,N_797);
or U9537 (N_9537,N_4821,N_4355);
nand U9538 (N_9538,N_4381,N_1213);
or U9539 (N_9539,N_2748,N_597);
nor U9540 (N_9540,N_1194,N_883);
or U9541 (N_9541,N_675,N_2140);
xnor U9542 (N_9542,N_4234,N_4187);
and U9543 (N_9543,N_4923,N_4382);
and U9544 (N_9544,N_570,N_65);
nor U9545 (N_9545,N_4516,N_3201);
and U9546 (N_9546,N_1345,N_1298);
or U9547 (N_9547,N_3646,N_4194);
nor U9548 (N_9548,N_3276,N_1841);
and U9549 (N_9549,N_910,N_653);
and U9550 (N_9550,N_4655,N_3298);
and U9551 (N_9551,N_4846,N_1458);
or U9552 (N_9552,N_4522,N_3672);
xnor U9553 (N_9553,N_4318,N_4607);
nand U9554 (N_9554,N_1404,N_3326);
nand U9555 (N_9555,N_3360,N_2018);
nor U9556 (N_9556,N_1344,N_2102);
nor U9557 (N_9557,N_1974,N_3496);
nor U9558 (N_9558,N_4359,N_3672);
or U9559 (N_9559,N_2890,N_2833);
nand U9560 (N_9560,N_4840,N_4465);
nand U9561 (N_9561,N_1637,N_219);
nand U9562 (N_9562,N_4967,N_1593);
nor U9563 (N_9563,N_919,N_936);
xor U9564 (N_9564,N_4161,N_239);
nor U9565 (N_9565,N_2046,N_629);
and U9566 (N_9566,N_2032,N_3145);
nand U9567 (N_9567,N_4512,N_3661);
and U9568 (N_9568,N_797,N_1749);
or U9569 (N_9569,N_1821,N_984);
nand U9570 (N_9570,N_813,N_1055);
or U9571 (N_9571,N_2965,N_2276);
nor U9572 (N_9572,N_750,N_3945);
and U9573 (N_9573,N_410,N_1750);
and U9574 (N_9574,N_3205,N_493);
nand U9575 (N_9575,N_3621,N_3);
xor U9576 (N_9576,N_2367,N_173);
and U9577 (N_9577,N_1288,N_3221);
and U9578 (N_9578,N_826,N_4684);
xnor U9579 (N_9579,N_3682,N_2273);
nor U9580 (N_9580,N_988,N_2525);
nand U9581 (N_9581,N_456,N_1767);
nand U9582 (N_9582,N_2014,N_2393);
or U9583 (N_9583,N_1060,N_448);
nand U9584 (N_9584,N_202,N_1890);
nand U9585 (N_9585,N_2446,N_2328);
nand U9586 (N_9586,N_4461,N_2692);
or U9587 (N_9587,N_4012,N_425);
nand U9588 (N_9588,N_1516,N_2702);
nor U9589 (N_9589,N_4279,N_2567);
or U9590 (N_9590,N_839,N_1806);
or U9591 (N_9591,N_359,N_4801);
nor U9592 (N_9592,N_3323,N_4815);
nand U9593 (N_9593,N_2391,N_141);
nand U9594 (N_9594,N_250,N_1774);
nor U9595 (N_9595,N_221,N_3871);
or U9596 (N_9596,N_81,N_2982);
and U9597 (N_9597,N_3632,N_1283);
and U9598 (N_9598,N_2142,N_1475);
xnor U9599 (N_9599,N_783,N_3541);
or U9600 (N_9600,N_961,N_1902);
or U9601 (N_9601,N_1295,N_3892);
or U9602 (N_9602,N_2917,N_602);
or U9603 (N_9603,N_1297,N_2417);
xnor U9604 (N_9604,N_4360,N_2310);
nand U9605 (N_9605,N_4782,N_4195);
and U9606 (N_9606,N_4997,N_4876);
or U9607 (N_9607,N_1159,N_3016);
nor U9608 (N_9608,N_3183,N_990);
or U9609 (N_9609,N_3559,N_2706);
nand U9610 (N_9610,N_2926,N_1126);
nor U9611 (N_9611,N_1213,N_170);
nor U9612 (N_9612,N_4914,N_4361);
xnor U9613 (N_9613,N_1635,N_2083);
nor U9614 (N_9614,N_1333,N_4106);
or U9615 (N_9615,N_3237,N_2399);
and U9616 (N_9616,N_3475,N_372);
and U9617 (N_9617,N_3953,N_1737);
and U9618 (N_9618,N_3314,N_821);
nor U9619 (N_9619,N_1945,N_4083);
nor U9620 (N_9620,N_2035,N_4024);
nand U9621 (N_9621,N_4439,N_137);
or U9622 (N_9622,N_3479,N_1725);
nor U9623 (N_9623,N_1931,N_2763);
and U9624 (N_9624,N_541,N_2280);
nor U9625 (N_9625,N_357,N_1773);
and U9626 (N_9626,N_1146,N_4387);
nor U9627 (N_9627,N_3721,N_339);
nand U9628 (N_9628,N_4709,N_3633);
nand U9629 (N_9629,N_4372,N_1655);
or U9630 (N_9630,N_4964,N_904);
nor U9631 (N_9631,N_3002,N_3405);
nor U9632 (N_9632,N_1613,N_2187);
and U9633 (N_9633,N_3295,N_894);
nor U9634 (N_9634,N_3124,N_1644);
or U9635 (N_9635,N_4311,N_2264);
and U9636 (N_9636,N_3767,N_3026);
nand U9637 (N_9637,N_487,N_3736);
nor U9638 (N_9638,N_3105,N_2978);
nor U9639 (N_9639,N_223,N_4091);
nand U9640 (N_9640,N_796,N_4496);
nor U9641 (N_9641,N_49,N_2439);
nand U9642 (N_9642,N_4825,N_874);
or U9643 (N_9643,N_2102,N_2665);
or U9644 (N_9644,N_1685,N_4967);
and U9645 (N_9645,N_4519,N_3324);
xnor U9646 (N_9646,N_269,N_4830);
nand U9647 (N_9647,N_1404,N_4574);
and U9648 (N_9648,N_1779,N_3812);
nand U9649 (N_9649,N_3976,N_3594);
or U9650 (N_9650,N_1427,N_1055);
nand U9651 (N_9651,N_4253,N_769);
or U9652 (N_9652,N_4352,N_2981);
nand U9653 (N_9653,N_754,N_2711);
or U9654 (N_9654,N_768,N_4641);
or U9655 (N_9655,N_3167,N_1059);
and U9656 (N_9656,N_4269,N_3863);
and U9657 (N_9657,N_3552,N_1908);
nor U9658 (N_9658,N_4311,N_2713);
and U9659 (N_9659,N_3861,N_589);
nor U9660 (N_9660,N_1213,N_4118);
and U9661 (N_9661,N_4098,N_4033);
nor U9662 (N_9662,N_1061,N_3913);
or U9663 (N_9663,N_1613,N_2776);
or U9664 (N_9664,N_2114,N_2343);
and U9665 (N_9665,N_2367,N_4982);
and U9666 (N_9666,N_488,N_1723);
nand U9667 (N_9667,N_1103,N_2539);
nand U9668 (N_9668,N_3535,N_3910);
or U9669 (N_9669,N_1357,N_836);
nand U9670 (N_9670,N_4519,N_3945);
or U9671 (N_9671,N_2449,N_1019);
or U9672 (N_9672,N_2408,N_962);
or U9673 (N_9673,N_1071,N_3178);
xnor U9674 (N_9674,N_191,N_535);
nor U9675 (N_9675,N_867,N_4842);
and U9676 (N_9676,N_3859,N_900);
nand U9677 (N_9677,N_3888,N_2789);
nor U9678 (N_9678,N_3875,N_2238);
and U9679 (N_9679,N_4829,N_1198);
nand U9680 (N_9680,N_696,N_3941);
nor U9681 (N_9681,N_4465,N_4635);
nand U9682 (N_9682,N_2496,N_4939);
and U9683 (N_9683,N_4846,N_3723);
nor U9684 (N_9684,N_2473,N_835);
nand U9685 (N_9685,N_4828,N_3220);
nor U9686 (N_9686,N_2573,N_2176);
and U9687 (N_9687,N_576,N_929);
nand U9688 (N_9688,N_4404,N_660);
and U9689 (N_9689,N_166,N_4200);
and U9690 (N_9690,N_3134,N_4895);
and U9691 (N_9691,N_2700,N_3762);
and U9692 (N_9692,N_4349,N_1288);
nand U9693 (N_9693,N_156,N_705);
and U9694 (N_9694,N_2296,N_3157);
or U9695 (N_9695,N_4157,N_1088);
nor U9696 (N_9696,N_2347,N_3013);
xnor U9697 (N_9697,N_3314,N_1077);
or U9698 (N_9698,N_4408,N_2042);
or U9699 (N_9699,N_4316,N_3212);
xor U9700 (N_9700,N_3636,N_986);
nor U9701 (N_9701,N_3284,N_238);
and U9702 (N_9702,N_4542,N_1640);
nor U9703 (N_9703,N_4882,N_1850);
and U9704 (N_9704,N_53,N_19);
and U9705 (N_9705,N_3130,N_3168);
or U9706 (N_9706,N_2890,N_3670);
nor U9707 (N_9707,N_1863,N_3337);
or U9708 (N_9708,N_4763,N_1563);
nand U9709 (N_9709,N_761,N_4851);
and U9710 (N_9710,N_352,N_4271);
nand U9711 (N_9711,N_2807,N_2838);
nand U9712 (N_9712,N_3064,N_753);
nand U9713 (N_9713,N_1043,N_1096);
and U9714 (N_9714,N_2150,N_2299);
and U9715 (N_9715,N_1187,N_2105);
nand U9716 (N_9716,N_621,N_2679);
and U9717 (N_9717,N_87,N_2738);
xnor U9718 (N_9718,N_4488,N_121);
nand U9719 (N_9719,N_530,N_4602);
nor U9720 (N_9720,N_1356,N_987);
and U9721 (N_9721,N_2872,N_846);
or U9722 (N_9722,N_292,N_2874);
or U9723 (N_9723,N_1968,N_2563);
nand U9724 (N_9724,N_3270,N_41);
nor U9725 (N_9725,N_2692,N_4617);
xnor U9726 (N_9726,N_3421,N_1524);
nand U9727 (N_9727,N_870,N_3998);
or U9728 (N_9728,N_3288,N_4893);
nand U9729 (N_9729,N_318,N_2888);
nand U9730 (N_9730,N_2531,N_563);
nor U9731 (N_9731,N_4040,N_2755);
and U9732 (N_9732,N_172,N_4829);
nor U9733 (N_9733,N_4020,N_841);
nor U9734 (N_9734,N_156,N_2255);
and U9735 (N_9735,N_895,N_3257);
and U9736 (N_9736,N_1397,N_4270);
nor U9737 (N_9737,N_4523,N_860);
and U9738 (N_9738,N_4509,N_4214);
nand U9739 (N_9739,N_558,N_3653);
and U9740 (N_9740,N_3687,N_4050);
nand U9741 (N_9741,N_29,N_4344);
and U9742 (N_9742,N_1717,N_1814);
or U9743 (N_9743,N_4487,N_245);
nand U9744 (N_9744,N_365,N_1434);
xor U9745 (N_9745,N_4520,N_41);
nor U9746 (N_9746,N_1070,N_4603);
nand U9747 (N_9747,N_3479,N_156);
nor U9748 (N_9748,N_1612,N_3773);
nand U9749 (N_9749,N_743,N_1247);
and U9750 (N_9750,N_4919,N_2386);
and U9751 (N_9751,N_4642,N_4362);
and U9752 (N_9752,N_2286,N_643);
nand U9753 (N_9753,N_3893,N_3766);
or U9754 (N_9754,N_2862,N_1636);
nand U9755 (N_9755,N_1769,N_3501);
xnor U9756 (N_9756,N_1145,N_280);
nand U9757 (N_9757,N_1875,N_1549);
nand U9758 (N_9758,N_4501,N_828);
or U9759 (N_9759,N_3838,N_2599);
nand U9760 (N_9760,N_4454,N_4951);
and U9761 (N_9761,N_499,N_4081);
nor U9762 (N_9762,N_4296,N_4941);
xor U9763 (N_9763,N_3038,N_1614);
or U9764 (N_9764,N_1665,N_731);
nor U9765 (N_9765,N_4958,N_1420);
xor U9766 (N_9766,N_60,N_2066);
or U9767 (N_9767,N_62,N_2116);
nor U9768 (N_9768,N_4930,N_4497);
nand U9769 (N_9769,N_2192,N_3327);
and U9770 (N_9770,N_3967,N_1342);
and U9771 (N_9771,N_4415,N_4145);
nor U9772 (N_9772,N_1111,N_4056);
and U9773 (N_9773,N_1464,N_3744);
and U9774 (N_9774,N_4409,N_4700);
and U9775 (N_9775,N_319,N_4124);
nand U9776 (N_9776,N_1365,N_1394);
xnor U9777 (N_9777,N_2793,N_3168);
nor U9778 (N_9778,N_4935,N_4853);
nor U9779 (N_9779,N_3360,N_4806);
xor U9780 (N_9780,N_2010,N_4865);
or U9781 (N_9781,N_4062,N_4700);
nor U9782 (N_9782,N_3278,N_4563);
and U9783 (N_9783,N_4678,N_1214);
or U9784 (N_9784,N_2425,N_4798);
or U9785 (N_9785,N_1269,N_3281);
nand U9786 (N_9786,N_42,N_1026);
nand U9787 (N_9787,N_4991,N_3975);
and U9788 (N_9788,N_1810,N_2620);
xnor U9789 (N_9789,N_61,N_3807);
or U9790 (N_9790,N_3398,N_4838);
and U9791 (N_9791,N_1152,N_2000);
nor U9792 (N_9792,N_3193,N_3320);
and U9793 (N_9793,N_4642,N_1529);
nand U9794 (N_9794,N_3930,N_2363);
xor U9795 (N_9795,N_4584,N_4560);
nor U9796 (N_9796,N_824,N_933);
or U9797 (N_9797,N_4784,N_4367);
or U9798 (N_9798,N_3682,N_2352);
or U9799 (N_9799,N_2576,N_151);
and U9800 (N_9800,N_2364,N_1240);
nor U9801 (N_9801,N_4902,N_4786);
or U9802 (N_9802,N_440,N_1786);
or U9803 (N_9803,N_2740,N_4309);
nand U9804 (N_9804,N_985,N_2194);
and U9805 (N_9805,N_2428,N_2104);
and U9806 (N_9806,N_1248,N_2713);
nor U9807 (N_9807,N_4020,N_190);
or U9808 (N_9808,N_3305,N_3383);
nor U9809 (N_9809,N_4131,N_4471);
and U9810 (N_9810,N_20,N_3656);
or U9811 (N_9811,N_683,N_3664);
and U9812 (N_9812,N_1134,N_3576);
nor U9813 (N_9813,N_4187,N_491);
xnor U9814 (N_9814,N_2204,N_4289);
and U9815 (N_9815,N_421,N_4567);
xnor U9816 (N_9816,N_4261,N_1902);
nand U9817 (N_9817,N_3389,N_4835);
and U9818 (N_9818,N_1776,N_2548);
or U9819 (N_9819,N_108,N_3918);
and U9820 (N_9820,N_3006,N_201);
and U9821 (N_9821,N_4788,N_1974);
or U9822 (N_9822,N_2147,N_3978);
or U9823 (N_9823,N_4744,N_4152);
and U9824 (N_9824,N_3196,N_850);
or U9825 (N_9825,N_2068,N_4352);
xor U9826 (N_9826,N_933,N_831);
nor U9827 (N_9827,N_3505,N_2759);
or U9828 (N_9828,N_2775,N_2639);
or U9829 (N_9829,N_431,N_577);
and U9830 (N_9830,N_3528,N_4950);
nor U9831 (N_9831,N_4083,N_665);
and U9832 (N_9832,N_1074,N_4220);
and U9833 (N_9833,N_4360,N_3099);
or U9834 (N_9834,N_1756,N_974);
nor U9835 (N_9835,N_4338,N_3302);
nand U9836 (N_9836,N_616,N_4548);
nand U9837 (N_9837,N_3249,N_1090);
nor U9838 (N_9838,N_3674,N_1025);
or U9839 (N_9839,N_3197,N_1883);
nand U9840 (N_9840,N_4723,N_4052);
nand U9841 (N_9841,N_2612,N_207);
and U9842 (N_9842,N_4769,N_640);
nand U9843 (N_9843,N_4289,N_222);
nor U9844 (N_9844,N_548,N_2457);
nor U9845 (N_9845,N_3252,N_2307);
or U9846 (N_9846,N_1791,N_1470);
nand U9847 (N_9847,N_4121,N_1380);
and U9848 (N_9848,N_2072,N_2400);
and U9849 (N_9849,N_3130,N_402);
and U9850 (N_9850,N_1762,N_3943);
xor U9851 (N_9851,N_711,N_283);
or U9852 (N_9852,N_1886,N_2299);
nor U9853 (N_9853,N_3059,N_3382);
xor U9854 (N_9854,N_3886,N_2056);
nor U9855 (N_9855,N_3935,N_2626);
or U9856 (N_9856,N_949,N_2803);
nand U9857 (N_9857,N_811,N_3331);
nor U9858 (N_9858,N_1504,N_1824);
or U9859 (N_9859,N_2349,N_1493);
nor U9860 (N_9860,N_2520,N_2465);
or U9861 (N_9861,N_984,N_757);
and U9862 (N_9862,N_1951,N_3136);
or U9863 (N_9863,N_1644,N_1214);
nand U9864 (N_9864,N_4997,N_3121);
nor U9865 (N_9865,N_1327,N_4606);
or U9866 (N_9866,N_2942,N_2391);
xnor U9867 (N_9867,N_1673,N_4011);
and U9868 (N_9868,N_2921,N_1844);
xnor U9869 (N_9869,N_3370,N_2798);
nor U9870 (N_9870,N_1111,N_3225);
or U9871 (N_9871,N_2773,N_4749);
or U9872 (N_9872,N_3000,N_2585);
and U9873 (N_9873,N_4764,N_3747);
nand U9874 (N_9874,N_2077,N_1894);
and U9875 (N_9875,N_4976,N_1791);
nor U9876 (N_9876,N_3906,N_1948);
nor U9877 (N_9877,N_2196,N_321);
or U9878 (N_9878,N_570,N_514);
nor U9879 (N_9879,N_4920,N_3554);
and U9880 (N_9880,N_1775,N_2986);
nand U9881 (N_9881,N_961,N_1970);
nor U9882 (N_9882,N_4208,N_2192);
nor U9883 (N_9883,N_3803,N_1156);
nor U9884 (N_9884,N_1548,N_932);
nor U9885 (N_9885,N_1074,N_1129);
nor U9886 (N_9886,N_3272,N_530);
or U9887 (N_9887,N_877,N_3370);
nand U9888 (N_9888,N_2290,N_3943);
xnor U9889 (N_9889,N_3047,N_1644);
nor U9890 (N_9890,N_2592,N_3746);
nand U9891 (N_9891,N_125,N_1163);
xnor U9892 (N_9892,N_1823,N_4506);
and U9893 (N_9893,N_1861,N_1993);
nor U9894 (N_9894,N_395,N_3561);
and U9895 (N_9895,N_118,N_1715);
and U9896 (N_9896,N_1021,N_3515);
nand U9897 (N_9897,N_4001,N_2958);
nor U9898 (N_9898,N_4433,N_2602);
and U9899 (N_9899,N_4208,N_1129);
and U9900 (N_9900,N_3926,N_461);
nand U9901 (N_9901,N_4602,N_1738);
xor U9902 (N_9902,N_4805,N_3252);
and U9903 (N_9903,N_1696,N_4295);
nand U9904 (N_9904,N_4540,N_3734);
nor U9905 (N_9905,N_741,N_3608);
nand U9906 (N_9906,N_139,N_3484);
and U9907 (N_9907,N_3711,N_2915);
or U9908 (N_9908,N_1595,N_469);
xnor U9909 (N_9909,N_560,N_1293);
or U9910 (N_9910,N_124,N_2542);
nand U9911 (N_9911,N_1571,N_1440);
nor U9912 (N_9912,N_1535,N_4392);
nand U9913 (N_9913,N_3992,N_3132);
nand U9914 (N_9914,N_908,N_2936);
and U9915 (N_9915,N_1892,N_450);
and U9916 (N_9916,N_1096,N_484);
nor U9917 (N_9917,N_4531,N_2884);
or U9918 (N_9918,N_2603,N_4859);
nand U9919 (N_9919,N_104,N_2980);
or U9920 (N_9920,N_2584,N_3069);
and U9921 (N_9921,N_268,N_1941);
and U9922 (N_9922,N_1309,N_3207);
or U9923 (N_9923,N_863,N_2483);
or U9924 (N_9924,N_3830,N_4544);
or U9925 (N_9925,N_2184,N_3612);
or U9926 (N_9926,N_3863,N_3592);
nand U9927 (N_9927,N_4146,N_1720);
and U9928 (N_9928,N_2263,N_2409);
and U9929 (N_9929,N_2639,N_3633);
or U9930 (N_9930,N_2737,N_723);
nand U9931 (N_9931,N_1812,N_2087);
or U9932 (N_9932,N_4477,N_94);
and U9933 (N_9933,N_3800,N_2399);
nand U9934 (N_9934,N_1043,N_858);
xor U9935 (N_9935,N_2994,N_2182);
nand U9936 (N_9936,N_3589,N_1370);
nand U9937 (N_9937,N_395,N_746);
nor U9938 (N_9938,N_7,N_98);
or U9939 (N_9939,N_2369,N_1290);
nand U9940 (N_9940,N_3208,N_746);
and U9941 (N_9941,N_1879,N_1700);
nand U9942 (N_9942,N_1271,N_2946);
nor U9943 (N_9943,N_2439,N_3637);
nor U9944 (N_9944,N_4285,N_2191);
nor U9945 (N_9945,N_3371,N_14);
or U9946 (N_9946,N_752,N_2694);
xnor U9947 (N_9947,N_1700,N_2018);
nand U9948 (N_9948,N_3964,N_370);
xnor U9949 (N_9949,N_14,N_2281);
nor U9950 (N_9950,N_2584,N_4427);
or U9951 (N_9951,N_2853,N_3617);
or U9952 (N_9952,N_1520,N_2890);
nand U9953 (N_9953,N_452,N_1801);
nand U9954 (N_9954,N_1279,N_3850);
nand U9955 (N_9955,N_862,N_1593);
and U9956 (N_9956,N_344,N_3993);
or U9957 (N_9957,N_381,N_4572);
xor U9958 (N_9958,N_551,N_892);
nor U9959 (N_9959,N_2228,N_4778);
nand U9960 (N_9960,N_4781,N_2980);
nand U9961 (N_9961,N_664,N_4050);
nand U9962 (N_9962,N_4395,N_4557);
and U9963 (N_9963,N_3162,N_3574);
nor U9964 (N_9964,N_4614,N_2360);
xor U9965 (N_9965,N_4276,N_396);
or U9966 (N_9966,N_3695,N_2229);
nor U9967 (N_9967,N_3615,N_1807);
nor U9968 (N_9968,N_577,N_4157);
or U9969 (N_9969,N_2706,N_3406);
nor U9970 (N_9970,N_2112,N_4649);
nand U9971 (N_9971,N_2231,N_3903);
and U9972 (N_9972,N_4854,N_2771);
xnor U9973 (N_9973,N_3607,N_4159);
or U9974 (N_9974,N_406,N_4094);
nand U9975 (N_9975,N_4953,N_615);
and U9976 (N_9976,N_4057,N_552);
and U9977 (N_9977,N_2263,N_1004);
nand U9978 (N_9978,N_2564,N_2409);
and U9979 (N_9979,N_4624,N_2562);
or U9980 (N_9980,N_2874,N_1115);
nor U9981 (N_9981,N_4621,N_3279);
or U9982 (N_9982,N_1573,N_1486);
nor U9983 (N_9983,N_2562,N_2241);
and U9984 (N_9984,N_1913,N_2235);
nand U9985 (N_9985,N_4591,N_1580);
nand U9986 (N_9986,N_2927,N_735);
nor U9987 (N_9987,N_4607,N_3364);
xor U9988 (N_9988,N_1067,N_2052);
nand U9989 (N_9989,N_3637,N_1489);
and U9990 (N_9990,N_2161,N_1980);
nor U9991 (N_9991,N_1481,N_3027);
xor U9992 (N_9992,N_4659,N_299);
xnor U9993 (N_9993,N_2449,N_1185);
nand U9994 (N_9994,N_3218,N_413);
and U9995 (N_9995,N_2871,N_3269);
and U9996 (N_9996,N_893,N_2033);
xor U9997 (N_9997,N_3246,N_3525);
xor U9998 (N_9998,N_4772,N_1098);
xor U9999 (N_9999,N_3975,N_1078);
nand UO_0 (O_0,N_6233,N_6347);
or UO_1 (O_1,N_6963,N_5110);
nor UO_2 (O_2,N_9649,N_9213);
nand UO_3 (O_3,N_9001,N_7050);
nor UO_4 (O_4,N_7246,N_8018);
or UO_5 (O_5,N_5840,N_7193);
nor UO_6 (O_6,N_8724,N_9966);
and UO_7 (O_7,N_8387,N_7624);
nand UO_8 (O_8,N_6523,N_6242);
or UO_9 (O_9,N_7539,N_5042);
or UO_10 (O_10,N_9331,N_5567);
and UO_11 (O_11,N_9126,N_5193);
and UO_12 (O_12,N_6144,N_6807);
and UO_13 (O_13,N_5172,N_7652);
and UO_14 (O_14,N_6305,N_8176);
and UO_15 (O_15,N_6149,N_9762);
nand UO_16 (O_16,N_7364,N_6394);
nand UO_17 (O_17,N_7920,N_9642);
xnor UO_18 (O_18,N_7253,N_6966);
xnor UO_19 (O_19,N_7650,N_8134);
nand UO_20 (O_20,N_7866,N_6107);
nor UO_21 (O_21,N_9919,N_8074);
nor UO_22 (O_22,N_7641,N_5050);
and UO_23 (O_23,N_5923,N_5558);
nand UO_24 (O_24,N_7728,N_7179);
nor UO_25 (O_25,N_8940,N_8734);
xnor UO_26 (O_26,N_9997,N_5237);
nor UO_27 (O_27,N_5958,N_5699);
and UO_28 (O_28,N_6450,N_6951);
and UO_29 (O_29,N_6042,N_6095);
or UO_30 (O_30,N_9296,N_5937);
nand UO_31 (O_31,N_5795,N_6945);
nor UO_32 (O_32,N_8283,N_7444);
nor UO_33 (O_33,N_6264,N_5857);
xnor UO_34 (O_34,N_5090,N_5538);
xor UO_35 (O_35,N_6863,N_8133);
or UO_36 (O_36,N_5025,N_7542);
nor UO_37 (O_37,N_9749,N_9596);
or UO_38 (O_38,N_5259,N_8336);
or UO_39 (O_39,N_7187,N_6499);
nand UO_40 (O_40,N_7344,N_5244);
nand UO_41 (O_41,N_7118,N_9345);
nor UO_42 (O_42,N_5955,N_7291);
nand UO_43 (O_43,N_9060,N_5587);
nor UO_44 (O_44,N_8777,N_5136);
nor UO_45 (O_45,N_5952,N_6543);
or UO_46 (O_46,N_5513,N_8902);
nand UO_47 (O_47,N_5564,N_6510);
and UO_48 (O_48,N_8651,N_8811);
nand UO_49 (O_49,N_5407,N_8181);
and UO_50 (O_50,N_9659,N_6634);
or UO_51 (O_51,N_7858,N_8369);
nor UO_52 (O_52,N_7445,N_7613);
nand UO_53 (O_53,N_7643,N_8084);
or UO_54 (O_54,N_6302,N_6583);
nand UO_55 (O_55,N_9839,N_6876);
nor UO_56 (O_56,N_6937,N_8689);
nor UO_57 (O_57,N_7662,N_5694);
or UO_58 (O_58,N_5082,N_5931);
nor UO_59 (O_59,N_9079,N_7688);
nor UO_60 (O_60,N_7914,N_9832);
nand UO_61 (O_61,N_8747,N_8898);
and UO_62 (O_62,N_8223,N_6687);
nand UO_63 (O_63,N_6911,N_8852);
nor UO_64 (O_64,N_5720,N_6231);
nor UO_65 (O_65,N_7100,N_8809);
nor UO_66 (O_66,N_6292,N_9259);
nor UO_67 (O_67,N_5003,N_8186);
and UO_68 (O_68,N_9690,N_9490);
nand UO_69 (O_69,N_6136,N_8569);
nand UO_70 (O_70,N_7215,N_9809);
and UO_71 (O_71,N_7047,N_7228);
nand UO_72 (O_72,N_9904,N_7350);
nor UO_73 (O_73,N_6732,N_6772);
or UO_74 (O_74,N_8831,N_7741);
xnor UO_75 (O_75,N_7956,N_9413);
and UO_76 (O_76,N_5843,N_5108);
or UO_77 (O_77,N_6935,N_8767);
and UO_78 (O_78,N_6195,N_6811);
nor UO_79 (O_79,N_9462,N_7239);
or UO_80 (O_80,N_7238,N_5234);
and UO_81 (O_81,N_6887,N_6457);
or UO_82 (O_82,N_6511,N_6984);
and UO_83 (O_83,N_7076,N_7658);
and UO_84 (O_84,N_5775,N_9167);
and UO_85 (O_85,N_5486,N_8788);
or UO_86 (O_86,N_6650,N_9967);
and UO_87 (O_87,N_8733,N_9896);
xor UO_88 (O_88,N_5447,N_9527);
xor UO_89 (O_89,N_6641,N_9816);
nor UO_90 (O_90,N_9540,N_6529);
or UO_91 (O_91,N_7702,N_8795);
nor UO_92 (O_92,N_9264,N_8436);
and UO_93 (O_93,N_8450,N_6260);
or UO_94 (O_94,N_5669,N_6629);
nand UO_95 (O_95,N_8103,N_8469);
or UO_96 (O_96,N_9033,N_5800);
nor UO_97 (O_97,N_9835,N_9025);
and UO_98 (O_98,N_6317,N_9751);
nand UO_99 (O_99,N_8679,N_5965);
and UO_100 (O_100,N_8548,N_7693);
or UO_101 (O_101,N_8467,N_6008);
xnor UO_102 (O_102,N_5076,N_5369);
nand UO_103 (O_103,N_6892,N_6429);
xnor UO_104 (O_104,N_7233,N_6412);
nand UO_105 (O_105,N_6205,N_6453);
nand UO_106 (O_106,N_5238,N_5263);
nor UO_107 (O_107,N_6454,N_5313);
nand UO_108 (O_108,N_6587,N_6840);
and UO_109 (O_109,N_9843,N_5198);
and UO_110 (O_110,N_6422,N_9147);
nor UO_111 (O_111,N_9491,N_8589);
nor UO_112 (O_112,N_6558,N_6537);
nor UO_113 (O_113,N_5596,N_7170);
and UO_114 (O_114,N_8933,N_5348);
xor UO_115 (O_115,N_7876,N_9685);
nand UO_116 (O_116,N_8764,N_6501);
and UO_117 (O_117,N_8434,N_6577);
xor UO_118 (O_118,N_7996,N_6448);
nor UO_119 (O_119,N_5554,N_8234);
nor UO_120 (O_120,N_9000,N_9849);
xor UO_121 (O_121,N_9111,N_5574);
nand UO_122 (O_122,N_7021,N_8858);
and UO_123 (O_123,N_5155,N_9183);
nor UO_124 (O_124,N_9306,N_8615);
or UO_125 (O_125,N_8822,N_7896);
xnor UO_126 (O_126,N_9684,N_8253);
or UO_127 (O_127,N_8715,N_9546);
and UO_128 (O_128,N_6100,N_6300);
and UO_129 (O_129,N_5748,N_9237);
nand UO_130 (O_130,N_9077,N_5444);
xnor UO_131 (O_131,N_7194,N_6981);
nor UO_132 (O_132,N_6635,N_7556);
and UO_133 (O_133,N_6921,N_8370);
or UO_134 (O_134,N_8519,N_7525);
or UO_135 (O_135,N_8033,N_9460);
or UO_136 (O_136,N_7391,N_9741);
nand UO_137 (O_137,N_7995,N_7292);
or UO_138 (O_138,N_5403,N_9875);
or UO_139 (O_139,N_5776,N_9542);
nand UO_140 (O_140,N_7682,N_5927);
and UO_141 (O_141,N_8271,N_5891);
or UO_142 (O_142,N_9847,N_5288);
and UO_143 (O_143,N_9370,N_9837);
and UO_144 (O_144,N_9784,N_7785);
nand UO_145 (O_145,N_6954,N_6249);
or UO_146 (O_146,N_5677,N_9838);
and UO_147 (O_147,N_8807,N_9100);
and UO_148 (O_148,N_8295,N_7340);
xnor UO_149 (O_149,N_9903,N_9421);
or UO_150 (O_150,N_8608,N_7001);
or UO_151 (O_151,N_9989,N_8053);
and UO_152 (O_152,N_5941,N_8984);
or UO_153 (O_153,N_5546,N_8646);
nand UO_154 (O_154,N_6513,N_5138);
nor UO_155 (O_155,N_5167,N_8435);
nand UO_156 (O_156,N_9892,N_9234);
nand UO_157 (O_157,N_7042,N_8009);
or UO_158 (O_158,N_7530,N_8622);
xor UO_159 (O_159,N_9821,N_7199);
nor UO_160 (O_160,N_7565,N_6924);
or UO_161 (O_161,N_9349,N_9670);
or UO_162 (O_162,N_7368,N_7882);
nor UO_163 (O_163,N_7842,N_7336);
and UO_164 (O_164,N_8443,N_7656);
or UO_165 (O_165,N_9566,N_9952);
and UO_166 (O_166,N_7147,N_7386);
nand UO_167 (O_167,N_6350,N_7294);
and UO_168 (O_168,N_7030,N_9092);
nor UO_169 (O_169,N_9764,N_8776);
or UO_170 (O_170,N_7016,N_7862);
or UO_171 (O_171,N_5966,N_8240);
and UO_172 (O_172,N_6222,N_9027);
and UO_173 (O_173,N_6392,N_6409);
and UO_174 (O_174,N_6157,N_6809);
and UO_175 (O_175,N_5229,N_7002);
and UO_176 (O_176,N_9528,N_8983);
and UO_177 (O_177,N_9728,N_5200);
nor UO_178 (O_178,N_7007,N_9002);
nor UO_179 (O_179,N_8031,N_5672);
xnor UO_180 (O_180,N_7033,N_5813);
and UO_181 (O_181,N_5255,N_6187);
xor UO_182 (O_182,N_8956,N_5612);
or UO_183 (O_183,N_5165,N_5910);
or UO_184 (O_184,N_6192,N_8787);
nand UO_185 (O_185,N_8083,N_8964);
nor UO_186 (O_186,N_8057,N_7310);
nor UO_187 (O_187,N_6118,N_6172);
nand UO_188 (O_188,N_5151,N_8325);
nand UO_189 (O_189,N_5926,N_5441);
nand UO_190 (O_190,N_6883,N_7320);
or UO_191 (O_191,N_6087,N_6662);
and UO_192 (O_192,N_7975,N_9752);
and UO_193 (O_193,N_9836,N_6571);
nor UO_194 (O_194,N_6737,N_7262);
nand UO_195 (O_195,N_8386,N_9610);
and UO_196 (O_196,N_8717,N_6725);
and UO_197 (O_197,N_5933,N_5548);
and UO_198 (O_198,N_8194,N_5632);
or UO_199 (O_199,N_6204,N_7628);
and UO_200 (O_200,N_7061,N_8460);
xnor UO_201 (O_201,N_7271,N_7775);
nand UO_202 (O_202,N_8743,N_9294);
and UO_203 (O_203,N_9484,N_8015);
nand UO_204 (O_204,N_6120,N_8324);
nand UO_205 (O_205,N_6020,N_6166);
xor UO_206 (O_206,N_9494,N_7383);
nor UO_207 (O_207,N_5251,N_7172);
or UO_208 (O_208,N_6138,N_6711);
and UO_209 (O_209,N_6419,N_8549);
nand UO_210 (O_210,N_9687,N_8292);
or UO_211 (O_211,N_5671,N_7488);
xnor UO_212 (O_212,N_7303,N_8707);
xnor UO_213 (O_213,N_7734,N_5466);
nor UO_214 (O_214,N_8596,N_9870);
nand UO_215 (O_215,N_5280,N_6256);
nand UO_216 (O_216,N_8228,N_9743);
xor UO_217 (O_217,N_8394,N_9080);
or UO_218 (O_218,N_8275,N_9552);
nor UO_219 (O_219,N_8123,N_9104);
nand UO_220 (O_220,N_7618,N_5541);
or UO_221 (O_221,N_6294,N_7904);
or UO_222 (O_222,N_6406,N_7925);
nand UO_223 (O_223,N_6534,N_8364);
nor UO_224 (O_224,N_6123,N_5802);
and UO_225 (O_225,N_9322,N_9124);
and UO_226 (O_226,N_6019,N_5604);
and UO_227 (O_227,N_8035,N_7796);
nor UO_228 (O_228,N_9885,N_6524);
and UO_229 (O_229,N_9763,N_7878);
and UO_230 (O_230,N_5452,N_7436);
and UO_231 (O_231,N_5493,N_8514);
or UO_232 (O_232,N_5159,N_8185);
or UO_233 (O_233,N_8236,N_8318);
xor UO_234 (O_234,N_8887,N_5638);
xor UO_235 (O_235,N_8060,N_9097);
or UO_236 (O_236,N_7070,N_9895);
xor UO_237 (O_237,N_9679,N_5723);
or UO_238 (O_238,N_7969,N_9558);
nor UO_239 (O_239,N_6857,N_8756);
nor UO_240 (O_240,N_9614,N_9564);
and UO_241 (O_241,N_6029,N_9616);
and UO_242 (O_242,N_7442,N_7088);
nand UO_243 (O_243,N_6532,N_9607);
and UO_244 (O_244,N_8393,N_8528);
or UO_245 (O_245,N_9689,N_5588);
nand UO_246 (O_246,N_9879,N_6940);
nor UO_247 (O_247,N_9216,N_6199);
nor UO_248 (O_248,N_5815,N_7214);
xor UO_249 (O_249,N_7675,N_8836);
or UO_250 (O_250,N_8613,N_8212);
xor UO_251 (O_251,N_6401,N_5654);
or UO_252 (O_252,N_8017,N_9329);
xor UO_253 (O_253,N_6855,N_7017);
and UO_254 (O_254,N_8575,N_6428);
nor UO_255 (O_255,N_6375,N_9361);
nor UO_256 (O_256,N_7983,N_9065);
nor UO_257 (O_257,N_8379,N_7242);
and UO_258 (O_258,N_9529,N_6817);
and UO_259 (O_259,N_5186,N_5409);
xor UO_260 (O_260,N_8881,N_8923);
and UO_261 (O_261,N_6194,N_8975);
nand UO_262 (O_262,N_6001,N_6722);
or UO_263 (O_263,N_9083,N_9501);
and UO_264 (O_264,N_7111,N_8782);
xnor UO_265 (O_265,N_8558,N_9164);
nand UO_266 (O_266,N_7282,N_8969);
nand UO_267 (O_267,N_9686,N_9961);
xnor UO_268 (O_268,N_5559,N_5132);
or UO_269 (O_269,N_9506,N_9834);
xor UO_270 (O_270,N_5014,N_9580);
nor UO_271 (O_271,N_9980,N_9049);
nand UO_272 (O_272,N_9074,N_5333);
nand UO_273 (O_273,N_7288,N_9760);
nor UO_274 (O_274,N_9585,N_7523);
or UO_275 (O_275,N_6145,N_6421);
nor UO_276 (O_276,N_6549,N_9754);
or UO_277 (O_277,N_8313,N_7148);
nand UO_278 (O_278,N_9737,N_8327);
and UO_279 (O_279,N_6539,N_8334);
nor UO_280 (O_280,N_5032,N_8545);
nor UO_281 (O_281,N_5741,N_8529);
or UO_282 (O_282,N_9524,N_5455);
nor UO_283 (O_283,N_6779,N_7255);
nand UO_284 (O_284,N_9854,N_7648);
xor UO_285 (O_285,N_6496,N_6751);
nor UO_286 (O_286,N_9909,N_7929);
nand UO_287 (O_287,N_7767,N_6893);
and UO_288 (O_288,N_6663,N_7544);
or UO_289 (O_289,N_5367,N_6573);
or UO_290 (O_290,N_8309,N_5460);
or UO_291 (O_291,N_9200,N_6498);
or UO_292 (O_292,N_8585,N_7418);
or UO_293 (O_293,N_7673,N_5153);
xnor UO_294 (O_294,N_7135,N_9038);
or UO_295 (O_295,N_7019,N_9269);
and UO_296 (O_296,N_8486,N_9787);
nand UO_297 (O_297,N_8866,N_5971);
nor UO_298 (O_298,N_8178,N_8588);
nand UO_299 (O_299,N_7776,N_7657);
nor UO_300 (O_300,N_9543,N_9458);
and UO_301 (O_301,N_6387,N_8030);
nor UO_302 (O_302,N_6075,N_6901);
or UO_303 (O_303,N_8422,N_8012);
or UO_304 (O_304,N_6324,N_8278);
and UO_305 (O_305,N_5213,N_6692);
nand UO_306 (O_306,N_7388,N_9195);
and UO_307 (O_307,N_5865,N_6699);
nand UO_308 (O_308,N_7339,N_7258);
and UO_309 (O_309,N_6011,N_9500);
xnor UO_310 (O_310,N_9639,N_6542);
or UO_311 (O_311,N_7132,N_8192);
nand UO_312 (O_312,N_8670,N_9015);
nand UO_313 (O_313,N_5063,N_5143);
xor UO_314 (O_314,N_7402,N_7063);
nor UO_315 (O_315,N_6796,N_6007);
nand UO_316 (O_316,N_9050,N_9094);
nand UO_317 (O_317,N_5477,N_8564);
xor UO_318 (O_318,N_8830,N_9781);
or UO_319 (O_319,N_5387,N_5667);
nand UO_320 (O_320,N_8119,N_8312);
nand UO_321 (O_321,N_5120,N_7491);
nor UO_322 (O_322,N_7510,N_9845);
nand UO_323 (O_323,N_9669,N_7529);
and UO_324 (O_324,N_7792,N_6560);
and UO_325 (O_325,N_6919,N_5219);
nand UO_326 (O_326,N_8461,N_6812);
or UO_327 (O_327,N_6851,N_7183);
or UO_328 (O_328,N_6582,N_8348);
and UO_329 (O_329,N_6069,N_9089);
nor UO_330 (O_330,N_6620,N_7760);
or UO_331 (O_331,N_8269,N_6198);
or UO_332 (O_332,N_9653,N_6735);
and UO_333 (O_333,N_9410,N_9852);
nor UO_334 (O_334,N_9113,N_9675);
nor UO_335 (O_335,N_5884,N_8572);
nand UO_336 (O_336,N_5192,N_9452);
or UO_337 (O_337,N_5994,N_9162);
and UO_338 (O_338,N_5305,N_8306);
nor UO_339 (O_339,N_7610,N_7981);
nor UO_340 (O_340,N_5633,N_8451);
nand UO_341 (O_341,N_9129,N_9655);
nand UO_342 (O_342,N_8444,N_6266);
nand UO_343 (O_343,N_6153,N_9811);
nor UO_344 (O_344,N_9794,N_8652);
and UO_345 (O_345,N_6372,N_9910);
and UO_346 (O_346,N_9785,N_9526);
nor UO_347 (O_347,N_7893,N_7653);
and UO_348 (O_348,N_5982,N_7783);
nor UO_349 (O_349,N_9654,N_7771);
nand UO_350 (O_350,N_7267,N_8560);
xor UO_351 (O_351,N_8930,N_9648);
and UO_352 (O_352,N_6151,N_9665);
or UO_353 (O_353,N_6006,N_6721);
nand UO_354 (O_354,N_9588,N_8955);
nand UO_355 (O_355,N_5079,N_6182);
and UO_356 (O_356,N_6415,N_6173);
or UO_357 (O_357,N_9099,N_6289);
or UO_358 (O_358,N_8741,N_9408);
or UO_359 (O_359,N_9403,N_9656);
and UO_360 (O_360,N_5938,N_7828);
xor UO_361 (O_361,N_7478,N_6739);
or UO_362 (O_362,N_8721,N_8511);
nand UO_363 (O_363,N_7101,N_9692);
nand UO_364 (O_364,N_8112,N_5324);
and UO_365 (O_365,N_7514,N_5344);
nand UO_366 (O_366,N_6698,N_8720);
nor UO_367 (O_367,N_9913,N_8331);
nor UO_368 (O_368,N_8049,N_9459);
nand UO_369 (O_369,N_8445,N_5326);
nand UO_370 (O_370,N_5017,N_8101);
or UO_371 (O_371,N_7210,N_8688);
xnor UO_372 (O_372,N_8595,N_7240);
nand UO_373 (O_373,N_5798,N_9076);
nor UO_374 (O_374,N_9982,N_7810);
and UO_375 (O_375,N_8465,N_9375);
nand UO_376 (O_376,N_7071,N_5093);
or UO_377 (O_377,N_5562,N_7689);
or UO_378 (O_378,N_9626,N_9145);
nor UO_379 (O_379,N_7945,N_5614);
or UO_380 (O_380,N_5180,N_9289);
nand UO_381 (O_381,N_7155,N_5418);
and UO_382 (O_382,N_9629,N_8000);
or UO_383 (O_383,N_6548,N_8990);
nand UO_384 (O_384,N_7762,N_9920);
xor UO_385 (O_385,N_7586,N_5092);
and UO_386 (O_386,N_8100,N_5202);
nand UO_387 (O_387,N_9444,N_7150);
xnor UO_388 (O_388,N_5207,N_7348);
or UO_389 (O_389,N_6086,N_9710);
nor UO_390 (O_390,N_8813,N_8859);
and UO_391 (O_391,N_7808,N_6273);
nor UO_392 (O_392,N_9231,N_6154);
nand UO_393 (O_393,N_5049,N_6969);
nor UO_394 (O_394,N_6340,N_8171);
xor UO_395 (O_395,N_7800,N_8517);
nor UO_396 (O_396,N_9698,N_7940);
nor UO_397 (O_397,N_7064,N_6041);
and UO_398 (O_398,N_8473,N_6398);
nor UO_399 (O_399,N_8220,N_5378);
and UO_400 (O_400,N_7837,N_6805);
nand UO_401 (O_401,N_6427,N_8922);
nand UO_402 (O_402,N_6143,N_7661);
or UO_403 (O_403,N_8428,N_6038);
and UO_404 (O_404,N_6031,N_8360);
or UO_405 (O_405,N_8222,N_6137);
and UO_406 (O_406,N_6269,N_9210);
and UO_407 (O_407,N_5635,N_6765);
or UO_408 (O_408,N_6783,N_9334);
and UO_409 (O_409,N_8280,N_9712);
xor UO_410 (O_410,N_8907,N_8132);
nand UO_411 (O_411,N_6424,N_9544);
nand UO_412 (O_412,N_9932,N_9426);
and UO_413 (O_413,N_9341,N_5801);
xor UO_414 (O_414,N_7011,N_8877);
nor UO_415 (O_415,N_6276,N_6600);
or UO_416 (O_416,N_5248,N_5561);
xnor UO_417 (O_417,N_7112,N_7965);
xor UO_418 (O_418,N_5631,N_6980);
and UO_419 (O_419,N_6990,N_6636);
nor UO_420 (O_420,N_6733,N_5870);
or UO_421 (O_421,N_8537,N_7855);
nand UO_422 (O_422,N_9779,N_7679);
nor UO_423 (O_423,N_6493,N_6533);
and UO_424 (O_424,N_9949,N_5957);
nand UO_425 (O_425,N_6624,N_8485);
nor UO_426 (O_426,N_5321,N_8642);
nor UO_427 (O_427,N_7202,N_7910);
and UO_428 (O_428,N_7883,N_5789);
or UO_429 (O_429,N_8438,N_5246);
nand UO_430 (O_430,N_9514,N_8617);
nand UO_431 (O_431,N_9914,N_8909);
nor UO_432 (O_432,N_6174,N_6178);
nand UO_433 (O_433,N_7521,N_9353);
and UO_434 (O_434,N_5586,N_6565);
and UO_435 (O_435,N_7463,N_7020);
and UO_436 (O_436,N_6649,N_5078);
or UO_437 (O_437,N_6232,N_6400);
xor UO_438 (O_438,N_5935,N_8408);
or UO_439 (O_439,N_9525,N_5896);
or UO_440 (O_440,N_8383,N_6251);
nand UO_441 (O_441,N_8052,N_9069);
and UO_442 (O_442,N_5819,N_7140);
nor UO_443 (O_443,N_9152,N_8584);
nand UO_444 (O_444,N_9174,N_5593);
nor UO_445 (O_445,N_9272,N_9551);
xnor UO_446 (O_446,N_7053,N_5976);
xnor UO_447 (O_447,N_9965,N_8891);
or UO_448 (O_448,N_7875,N_8685);
or UO_449 (O_449,N_6303,N_5341);
and UO_450 (O_450,N_7752,N_7173);
or UO_451 (O_451,N_8203,N_7901);
or UO_452 (O_452,N_7280,N_6931);
and UO_453 (O_453,N_8641,N_9667);
nand UO_454 (O_454,N_6838,N_8980);
nor UO_455 (O_455,N_7373,N_6009);
or UO_456 (O_456,N_8751,N_7933);
nor UO_457 (O_457,N_8260,N_8796);
nor UO_458 (O_458,N_9971,N_9575);
nor UO_459 (O_459,N_8346,N_8124);
nor UO_460 (O_460,N_8570,N_6139);
and UO_461 (O_461,N_9004,N_8742);
nor UO_462 (O_462,N_7162,N_5171);
xnor UO_463 (O_463,N_5760,N_9651);
and UO_464 (O_464,N_8417,N_8301);
nor UO_465 (O_465,N_7554,N_7988);
or UO_466 (O_466,N_6865,N_7839);
nand UO_467 (O_467,N_7748,N_9569);
or UO_468 (O_468,N_7835,N_5785);
and UO_469 (O_469,N_5517,N_7632);
xor UO_470 (O_470,N_8135,N_9621);
nor UO_471 (O_471,N_9425,N_5827);
or UO_472 (O_472,N_9409,N_6544);
or UO_473 (O_473,N_6227,N_8712);
or UO_474 (O_474,N_7324,N_9461);
or UO_475 (O_475,N_8197,N_9084);
and UO_476 (O_476,N_9937,N_7302);
xor UO_477 (O_477,N_8482,N_7713);
and UO_478 (O_478,N_5644,N_8546);
and UO_479 (O_479,N_5179,N_5682);
nand UO_480 (O_480,N_8948,N_7804);
or UO_481 (O_481,N_7129,N_5307);
nor UO_482 (O_482,N_9820,N_8165);
nand UO_483 (O_483,N_5437,N_6470);
nor UO_484 (O_484,N_8003,N_8849);
or UO_485 (O_485,N_6665,N_7278);
or UO_486 (O_486,N_5889,N_6670);
nand UO_487 (O_487,N_5363,N_8043);
nor UO_488 (O_488,N_5662,N_9715);
nor UO_489 (O_489,N_6342,N_6832);
nand UO_490 (O_490,N_8047,N_9405);
nand UO_491 (O_491,N_7308,N_9993);
nand UO_492 (O_492,N_9746,N_5376);
nor UO_493 (O_493,N_5894,N_8586);
and UO_494 (O_494,N_8338,N_6081);
and UO_495 (O_495,N_9576,N_9144);
and UO_496 (O_496,N_9652,N_5649);
or UO_497 (O_497,N_7720,N_6525);
nor UO_498 (O_498,N_6605,N_7372);
nor UO_499 (O_499,N_9947,N_6517);
nor UO_500 (O_500,N_5318,N_8268);
nand UO_501 (O_501,N_6456,N_5973);
nor UO_502 (O_502,N_8198,N_9010);
nor UO_503 (O_503,N_9646,N_9482);
nor UO_504 (O_504,N_6678,N_5361);
nand UO_505 (O_505,N_6512,N_6270);
and UO_506 (O_506,N_5847,N_7353);
nand UO_507 (O_507,N_7094,N_9633);
xor UO_508 (O_508,N_6899,N_7369);
nor UO_509 (O_509,N_9376,N_7322);
xor UO_510 (O_510,N_7034,N_8970);
or UO_511 (O_511,N_7158,N_6247);
xnor UO_512 (O_512,N_9934,N_5111);
or UO_513 (O_513,N_9850,N_5600);
or UO_514 (O_514,N_6999,N_5446);
and UO_515 (O_515,N_9562,N_5940);
nor UO_516 (O_516,N_5774,N_7376);
nand UO_517 (O_517,N_5823,N_6396);
and UO_518 (O_518,N_7881,N_9578);
nor UO_519 (O_519,N_6900,N_8580);
nor UO_520 (O_520,N_9222,N_5849);
nand UO_521 (O_521,N_6640,N_6661);
or UO_522 (O_522,N_7516,N_9282);
nand UO_523 (O_523,N_5284,N_7692);
and UO_524 (O_524,N_5695,N_5535);
and UO_525 (O_525,N_9207,N_7329);
and UO_526 (O_526,N_7103,N_5401);
nand UO_527 (O_527,N_7077,N_7846);
or UO_528 (O_528,N_7949,N_7968);
nand UO_529 (O_529,N_8345,N_5515);
and UO_530 (O_530,N_9328,N_9005);
nor UO_531 (O_531,N_7182,N_6112);
and UO_532 (O_532,N_5400,N_9660);
and UO_533 (O_533,N_6440,N_8433);
or UO_534 (O_534,N_5825,N_7588);
nor UO_535 (O_535,N_9512,N_9146);
nor UO_536 (O_536,N_7923,N_8963);
nand UO_537 (O_537,N_8977,N_5904);
nor UO_538 (O_538,N_5960,N_8648);
nand UO_539 (O_539,N_8105,N_5834);
nor UO_540 (O_540,N_6410,N_5221);
or UO_541 (O_541,N_9594,N_5147);
and UO_542 (O_542,N_8357,N_7106);
nor UO_543 (O_543,N_8001,N_9242);
or UO_544 (O_544,N_6939,N_5886);
and UO_545 (O_545,N_7286,N_7195);
nor UO_546 (O_546,N_6727,N_6741);
nand UO_547 (O_547,N_6024,N_5911);
or UO_548 (O_548,N_7205,N_9086);
nand UO_549 (O_549,N_6810,N_8491);
nand UO_550 (O_550,N_9897,N_8783);
xor UO_551 (O_551,N_7780,N_9876);
or UO_552 (O_552,N_8912,N_8279);
nor UO_553 (O_553,N_9972,N_5523);
xor UO_554 (O_554,N_8117,N_7151);
or UO_555 (O_555,N_6657,N_9381);
nand UO_556 (O_556,N_8439,N_7043);
or UO_557 (O_557,N_9355,N_5793);
or UO_558 (O_558,N_5618,N_8291);
nor UO_559 (O_559,N_7356,N_9933);
nand UO_560 (O_560,N_6878,N_8536);
nor UO_561 (O_561,N_5585,N_8027);
xor UO_562 (O_562,N_7270,N_7895);
nand UO_563 (O_563,N_5750,N_5728);
or UO_564 (O_564,N_5433,N_6689);
or UO_565 (O_565,N_8693,N_8244);
or UO_566 (O_566,N_5681,N_5380);
nand UO_567 (O_567,N_7395,N_7768);
nor UO_568 (O_568,N_6218,N_6977);
nand UO_569 (O_569,N_8500,N_9807);
nor UO_570 (O_570,N_5848,N_9186);
and UO_571 (O_571,N_7105,N_7830);
xnor UO_572 (O_572,N_6891,N_5379);
and UO_573 (O_573,N_5686,N_8986);
and UO_574 (O_574,N_8146,N_5853);
nor UO_575 (O_575,N_7473,N_8085);
or UO_576 (O_576,N_5373,N_6079);
nand UO_577 (O_577,N_8711,N_6220);
xor UO_578 (O_578,N_6658,N_9247);
and UO_579 (O_579,N_7979,N_5839);
or UO_580 (O_580,N_9072,N_7479);
nand UO_581 (O_581,N_8215,N_5721);
or UO_582 (O_582,N_5254,N_5715);
and UO_583 (O_583,N_7726,N_9003);
or UO_584 (O_584,N_8844,N_9275);
nand UO_585 (O_585,N_6093,N_8640);
nand UO_586 (O_586,N_7816,N_6703);
or UO_587 (O_587,N_7986,N_9536);
nand UO_588 (O_588,N_8934,N_5162);
nand UO_589 (O_589,N_9040,N_5902);
and UO_590 (O_590,N_5140,N_5808);
or UO_591 (O_591,N_7108,N_5974);
nand UO_592 (O_592,N_5236,N_8582);
or UO_593 (O_593,N_6842,N_9379);
or UO_594 (O_594,N_6979,N_7642);
or UO_595 (O_595,N_8056,N_6835);
and UO_596 (O_596,N_5303,N_9940);
and UO_597 (O_597,N_7387,N_7880);
or UO_598 (O_598,N_7477,N_8541);
nand UO_599 (O_599,N_8656,N_6091);
nand UO_600 (O_600,N_9777,N_7939);
nand UO_601 (O_601,N_6655,N_7931);
or UO_602 (O_602,N_9008,N_6830);
or UO_603 (O_603,N_7801,N_5115);
and UO_604 (O_604,N_6135,N_7206);
or UO_605 (O_605,N_6364,N_7054);
nand UO_606 (O_606,N_9725,N_8157);
nor UO_607 (O_607,N_6535,N_7695);
or UO_608 (O_608,N_7786,N_9627);
and UO_609 (O_609,N_7178,N_5921);
and UO_610 (O_610,N_7959,N_7857);
and UO_611 (O_611,N_8025,N_9523);
and UO_612 (O_612,N_7404,N_6724);
nor UO_613 (O_613,N_7526,N_9371);
nand UO_614 (O_614,N_7799,N_8039);
nand UO_615 (O_615,N_8069,N_6825);
or UO_616 (O_616,N_6293,N_6894);
nor UO_617 (O_617,N_6134,N_9505);
nand UO_618 (O_618,N_7879,N_7621);
or UO_619 (O_619,N_8917,N_7217);
and UO_620 (O_620,N_9071,N_9324);
and UO_621 (O_621,N_8402,N_6253);
nand UO_622 (O_622,N_8619,N_6402);
or UO_623 (O_623,N_5757,N_6039);
nand UO_624 (O_624,N_7074,N_9694);
nor UO_625 (O_625,N_7973,N_8427);
or UO_626 (O_626,N_9959,N_8609);
nand UO_627 (O_627,N_6349,N_7045);
nand UO_628 (O_628,N_8144,N_8152);
and UO_629 (O_629,N_8994,N_5040);
nand UO_630 (O_630,N_5540,N_6547);
nor UO_631 (O_631,N_5414,N_9814);
or UO_632 (O_632,N_9978,N_8389);
and UO_633 (O_633,N_9537,N_8878);
xor UO_634 (O_634,N_5787,N_8518);
or UO_635 (O_635,N_9704,N_7326);
nor UO_636 (O_636,N_5995,N_9791);
xnor UO_637 (O_637,N_5392,N_9351);
or UO_638 (O_638,N_8137,N_5591);
nand UO_639 (O_639,N_5850,N_8636);
nand UO_640 (O_640,N_7458,N_7441);
or UO_641 (O_641,N_8871,N_6978);
nor UO_642 (O_642,N_7597,N_5817);
and UO_643 (O_643,N_9808,N_5037);
nor UO_644 (O_644,N_8109,N_7367);
nand UO_645 (O_645,N_9135,N_8310);
and UO_646 (O_646,N_8987,N_7023);
and UO_647 (O_647,N_9175,N_6077);
and UO_648 (O_648,N_7104,N_7412);
nand UO_649 (O_649,N_8339,N_7966);
and UO_650 (O_650,N_6750,N_5946);
nor UO_651 (O_651,N_7360,N_7235);
nor UO_652 (O_652,N_9360,N_5570);
or UO_653 (O_653,N_6986,N_5768);
and UO_654 (O_654,N_7026,N_6062);
nand UO_655 (O_655,N_9890,N_7685);
or UO_656 (O_656,N_8332,N_5530);
and UO_657 (O_657,N_9202,N_8629);
nand UO_658 (O_658,N_5177,N_6485);
nand UO_659 (O_659,N_8921,N_7802);
nor UO_660 (O_660,N_8051,N_8535);
nor UO_661 (O_661,N_5897,N_8254);
nor UO_662 (O_662,N_5895,N_5828);
nor UO_663 (O_663,N_9463,N_7701);
nor UO_664 (O_664,N_9036,N_9303);
nor UO_665 (O_665,N_7594,N_8669);
or UO_666 (O_666,N_6971,N_7560);
nor UO_667 (O_667,N_6902,N_7055);
nand UO_668 (O_668,N_7851,N_8769);
or UO_669 (O_669,N_6325,N_8512);
nand UO_670 (O_670,N_7352,N_7006);
nor UO_671 (O_671,N_5860,N_6203);
nor UO_672 (O_672,N_6925,N_6743);
and UO_673 (O_673,N_8065,N_6834);
nand UO_674 (O_674,N_7845,N_9803);
nand UO_675 (O_675,N_6568,N_6803);
nand UO_676 (O_676,N_8125,N_7138);
nand UO_677 (O_677,N_6083,N_8699);
and UO_678 (O_678,N_9747,N_6562);
and UO_679 (O_679,N_6612,N_5944);
nand UO_680 (O_680,N_7013,N_5967);
nor UO_681 (O_681,N_6623,N_6526);
xor UO_682 (O_682,N_9078,N_5125);
xnor UO_683 (O_683,N_8799,N_5287);
xnor UO_684 (O_684,N_8846,N_9865);
and UO_685 (O_685,N_9680,N_7717);
and UO_686 (O_686,N_8924,N_6224);
nand UO_687 (O_687,N_6749,N_5105);
nand UO_688 (O_688,N_8322,N_5024);
nand UO_689 (O_689,N_7821,N_7927);
and UO_690 (O_690,N_6012,N_5124);
and UO_691 (O_691,N_6228,N_7736);
xnor UO_692 (O_692,N_7543,N_8766);
xnor UO_693 (O_693,N_5516,N_5687);
nor UO_694 (O_694,N_8989,N_9395);
xnor UO_695 (O_695,N_7941,N_6471);
nand UO_696 (O_696,N_8276,N_6890);
or UO_697 (O_697,N_8915,N_7795);
or UO_698 (O_698,N_9103,N_7284);
nor UO_699 (O_699,N_5166,N_8399);
nand UO_700 (O_700,N_5482,N_6546);
xnor UO_701 (O_701,N_9299,N_8412);
and UO_702 (O_702,N_8655,N_5371);
or UO_703 (O_703,N_6378,N_6358);
or UO_704 (O_704,N_8735,N_8653);
nand UO_705 (O_705,N_5231,N_7490);
or UO_706 (O_706,N_9553,N_9534);
and UO_707 (O_707,N_9101,N_7564);
or UO_708 (O_708,N_9107,N_6507);
xor UO_709 (O_709,N_8361,N_8791);
or UO_710 (O_710,N_7464,N_8202);
nand UO_711 (O_711,N_8627,N_6576);
nand UO_712 (O_712,N_7384,N_6104);
nand UO_713 (O_713,N_7697,N_8034);
nand UO_714 (O_714,N_8219,N_8573);
nand UO_715 (O_715,N_6381,N_6972);
nand UO_716 (O_716,N_8163,N_5069);
and UO_717 (O_717,N_5816,N_7232);
or UO_718 (O_718,N_8068,N_6758);
and UO_719 (O_719,N_8139,N_6944);
and UO_720 (O_720,N_6284,N_7990);
and UO_721 (O_721,N_8945,N_9579);
and UO_722 (O_722,N_9786,N_8114);
nor UO_723 (O_723,N_5664,N_5383);
and UO_724 (O_724,N_6117,N_5898);
or UO_725 (O_725,N_9705,N_6514);
xnor UO_726 (O_726,N_7212,N_6604);
and UO_727 (O_727,N_6988,N_6704);
and UO_728 (O_728,N_7861,N_9336);
nand UO_729 (O_729,N_6506,N_6594);
xor UO_730 (O_730,N_6016,N_9701);
or UO_731 (O_731,N_5413,N_9945);
nand UO_732 (O_732,N_6344,N_5660);
or UO_733 (O_733,N_7950,N_9662);
xor UO_734 (O_734,N_7306,N_5113);
or UO_735 (O_735,N_5432,N_9573);
and UO_736 (O_736,N_5794,N_6351);
and UO_737 (O_737,N_8726,N_6074);
xnor UO_738 (O_738,N_8297,N_8821);
and UO_739 (O_739,N_7272,N_7236);
nor UO_740 (O_740,N_5529,N_9280);
nor UO_741 (O_741,N_5056,N_8145);
xnor UO_742 (O_742,N_9771,N_9317);
and UO_743 (O_743,N_6125,N_8532);
and UO_744 (O_744,N_8521,N_8358);
nand UO_745 (O_745,N_7203,N_9859);
and UO_746 (O_746,N_6987,N_6023);
nor UO_747 (O_747,N_6147,N_9825);
and UO_748 (O_748,N_5389,N_9887);
nor UO_749 (O_749,N_7605,N_7470);
nor UO_750 (O_750,N_6245,N_6463);
and UO_751 (O_751,N_5993,N_5215);
nor UO_752 (O_752,N_9681,N_9047);
or UO_753 (O_753,N_5007,N_5531);
or UO_754 (O_754,N_8182,N_9091);
nand UO_755 (O_755,N_7218,N_8853);
xor UO_756 (O_756,N_5209,N_9957);
and UO_757 (O_757,N_5435,N_5919);
and UO_758 (O_758,N_7549,N_6319);
or UO_759 (O_759,N_6430,N_5908);
or UO_760 (O_760,N_7869,N_9830);
nand UO_761 (O_761,N_7018,N_8967);
nor UO_762 (O_762,N_5980,N_5939);
and UO_763 (O_763,N_9445,N_7377);
or UO_764 (O_764,N_7250,N_6997);
and UO_765 (O_765,N_8806,N_6553);
nand UO_766 (O_766,N_6208,N_9206);
xor UO_767 (O_767,N_8078,N_8894);
nor UO_768 (O_768,N_8946,N_5996);
nand UO_769 (O_769,N_9179,N_8610);
nor UO_770 (O_770,N_5758,N_5782);
nand UO_771 (O_771,N_9600,N_5424);
or UO_772 (O_772,N_9538,N_8966);
or UO_773 (O_773,N_9871,N_9451);
xor UO_774 (O_774,N_6808,N_8768);
xnor UO_775 (O_775,N_6866,N_8935);
nor UO_776 (O_776,N_5261,N_5325);
nand UO_777 (O_777,N_9154,N_9968);
and UO_778 (O_778,N_7812,N_9898);
and UO_779 (O_779,N_9605,N_9590);
or UO_780 (O_780,N_9325,N_5680);
nand UO_781 (O_781,N_6480,N_8504);
and UO_782 (O_782,N_8638,N_5285);
nor UO_783 (O_783,N_6184,N_6974);
or UO_784 (O_784,N_9634,N_5930);
xor UO_785 (O_785,N_8718,N_9851);
nand UO_786 (O_786,N_7224,N_8920);
nand UO_787 (O_787,N_6516,N_7419);
or UO_788 (O_788,N_7485,N_5726);
or UO_789 (O_789,N_6414,N_9163);
or UO_790 (O_790,N_5065,N_6078);
and UO_791 (O_791,N_5045,N_6246);
nand UO_792 (O_792,N_7578,N_7886);
nand UO_793 (O_793,N_9270,N_5298);
nand UO_794 (O_794,N_6370,N_9772);
nand UO_795 (O_795,N_6278,N_5643);
nand UO_796 (O_796,N_7755,N_7868);
and UO_797 (O_797,N_6423,N_9853);
nand UO_798 (O_798,N_9866,N_9638);
nand UO_799 (O_799,N_8960,N_8213);
nand UO_800 (O_800,N_6179,N_5469);
or UO_801 (O_801,N_8044,N_6509);
nand UO_802 (O_802,N_5637,N_9298);
or UO_803 (O_803,N_5347,N_6559);
and UO_804 (O_804,N_9657,N_8810);
nor UO_805 (O_805,N_5064,N_7139);
or UO_806 (O_806,N_5704,N_7184);
nor UO_807 (O_807,N_8430,N_5187);
or UO_808 (O_808,N_5097,N_9173);
nand UO_809 (O_809,N_6684,N_6051);
or UO_810 (O_810,N_8630,N_5416);
nand UO_811 (O_811,N_7465,N_6255);
xnor UO_812 (O_812,N_8449,N_5175);
or UO_813 (O_813,N_9245,N_6527);
and UO_814 (O_814,N_6952,N_5572);
nor UO_815 (O_815,N_5006,N_7027);
nor UO_816 (O_816,N_5309,N_9488);
nor UO_817 (O_817,N_5315,N_7408);
nand UO_818 (O_818,N_5601,N_6983);
and UO_819 (O_819,N_8773,N_9719);
or UO_820 (O_820,N_9256,N_5310);
and UO_821 (O_821,N_8277,N_8951);
or UO_822 (O_822,N_8649,N_5072);
and UO_823 (O_823,N_9899,N_9260);
nor UO_824 (O_824,N_9437,N_9559);
and UO_825 (O_825,N_5883,N_7844);
nor UO_826 (O_826,N_7117,N_8496);
nand UO_827 (O_827,N_5500,N_7130);
nand UO_828 (O_828,N_8187,N_6730);
nor UO_829 (O_829,N_8631,N_6254);
xor UO_830 (O_830,N_5756,N_8755);
xor UO_831 (O_831,N_9483,N_8136);
nand UO_832 (O_832,N_5858,N_9189);
or UO_833 (O_833,N_5189,N_5869);
and UO_834 (O_834,N_7434,N_5900);
and UO_835 (O_835,N_9449,N_8744);
and UO_836 (O_836,N_8526,N_8716);
nand UO_837 (O_837,N_7915,N_6064);
and UO_838 (O_838,N_9495,N_8456);
nand UO_839 (O_839,N_9498,N_7079);
or UO_840 (O_840,N_9118,N_9666);
and UO_841 (O_841,N_9187,N_6250);
xnor UO_842 (O_842,N_7805,N_5780);
or UO_843 (O_843,N_6279,N_5253);
or UO_844 (O_844,N_5483,N_5491);
nand UO_845 (O_845,N_5752,N_5605);
xnor UO_846 (O_846,N_8819,N_8259);
nand UO_847 (O_847,N_8262,N_8786);
nand UO_848 (O_848,N_5112,N_6656);
nor UO_849 (O_849,N_6367,N_5278);
and UO_850 (O_850,N_7174,N_8173);
or UO_851 (O_851,N_7375,N_9996);
nand UO_852 (O_852,N_8195,N_9757);
and UO_853 (O_853,N_7769,N_6202);
nand UO_854 (O_854,N_7343,N_6660);
or UO_855 (O_855,N_9574,N_8062);
or UO_856 (O_856,N_8765,N_6538);
nand UO_857 (O_857,N_5425,N_5778);
and UO_858 (O_858,N_7012,N_7899);
nand UO_859 (O_859,N_7672,N_5152);
nor UO_860 (O_860,N_9007,N_9333);
xnor UO_861 (O_861,N_5235,N_6141);
and UO_862 (O_862,N_7684,N_8130);
and UO_863 (O_863,N_9307,N_6003);
and UO_864 (O_864,N_7976,N_7935);
nor UO_865 (O_865,N_9990,N_9278);
nand UO_866 (O_866,N_7461,N_9321);
or UO_867 (O_867,N_5514,N_8227);
nand UO_868 (O_868,N_8363,N_5038);
xor UO_869 (O_869,N_8938,N_6993);
nor UO_870 (O_870,N_6590,N_8081);
or UO_871 (O_871,N_6160,N_5893);
and UO_872 (O_872,N_7541,N_5240);
nor UO_873 (O_873,N_6877,N_7625);
xor UO_874 (O_874,N_6770,N_8962);
nand UO_875 (O_875,N_7847,N_8175);
or UO_876 (O_876,N_7739,N_7806);
and UO_877 (O_877,N_8184,N_7872);
xnor UO_878 (O_878,N_7483,N_8941);
nor UO_879 (O_879,N_6073,N_8525);
nor UO_880 (O_880,N_9618,N_7874);
or UO_881 (O_881,N_6748,N_8509);
and UO_882 (O_882,N_6814,N_7829);
and UO_883 (O_883,N_7004,N_8385);
nor UO_884 (O_884,N_8719,N_5557);
or UO_885 (O_885,N_5731,N_8342);
or UO_886 (O_886,N_8530,N_6502);
xor UO_887 (O_887,N_8229,N_5137);
nor UO_888 (O_888,N_6235,N_7185);
xnor UO_889 (O_889,N_9414,N_8612);
and UO_890 (O_890,N_9447,N_6285);
nand UO_891 (O_891,N_7598,N_8046);
nor UO_892 (O_892,N_7687,N_8870);
nor UO_893 (O_893,N_9521,N_7120);
nor UO_894 (O_894,N_5734,N_6459);
nand UO_895 (O_895,N_7361,N_5398);
or UO_896 (O_896,N_8547,N_5454);
or UO_897 (O_897,N_5629,N_6146);
xor UO_898 (O_898,N_7977,N_8007);
and UO_899 (O_899,N_9456,N_8026);
nand UO_900 (O_900,N_6164,N_9636);
nor UO_901 (O_901,N_6614,N_7188);
or UO_902 (O_902,N_8959,N_6859);
or UO_903 (O_903,N_9044,N_5106);
or UO_904 (O_904,N_6777,N_9316);
xor UO_905 (O_905,N_8885,N_8676);
xor UO_906 (O_906,N_8659,N_7327);
and UO_907 (O_907,N_7699,N_9508);
nor UO_908 (O_908,N_6186,N_6185);
nor UO_909 (O_909,N_8727,N_9045);
nor UO_910 (O_910,N_6617,N_8359);
nor UO_911 (O_911,N_8763,N_8016);
and UO_912 (O_912,N_8248,N_7957);
xor UO_913 (O_913,N_6341,N_8562);
or UO_914 (O_914,N_7220,N_6361);
or UO_915 (O_915,N_6716,N_8698);
and UO_916 (O_916,N_6719,N_7854);
or UO_917 (O_917,N_5864,N_9309);
nor UO_918 (O_918,N_6494,N_7338);
nor UO_919 (O_919,N_5977,N_5342);
and UO_920 (O_920,N_9311,N_7499);
nand UO_921 (O_921,N_8183,N_9373);
nand UO_922 (O_922,N_5122,N_8209);
and UO_923 (O_923,N_8723,N_8063);
and UO_924 (O_924,N_6200,N_8050);
nand UO_925 (O_925,N_7905,N_9717);
nor UO_926 (O_926,N_9121,N_5584);
or UO_927 (O_927,N_6366,N_5476);
xnor UO_928 (O_928,N_6054,N_5266);
xor UO_929 (O_929,N_5286,N_8992);
and UO_930 (O_930,N_5693,N_5226);
nor UO_931 (O_931,N_9872,N_5674);
and UO_932 (O_932,N_7406,N_5575);
or UO_933 (O_933,N_8416,N_6158);
nor UO_934 (O_934,N_5279,N_9013);
nand UO_935 (O_935,N_6742,N_5805);
xnor UO_936 (O_936,N_9168,N_5009);
and UO_937 (O_937,N_5566,N_5026);
nand UO_938 (O_938,N_7044,N_5144);
nor UO_939 (O_939,N_7602,N_6578);
nand UO_940 (O_940,N_9258,N_7119);
or UO_941 (O_941,N_5761,N_7298);
and UO_942 (O_942,N_7476,N_5781);
nand UO_943 (O_943,N_8356,N_7166);
nand UO_944 (O_944,N_6697,N_6800);
and UO_945 (O_945,N_8979,N_5170);
or UO_946 (O_946,N_9767,N_9141);
nand UO_947 (O_947,N_9106,N_5098);
and UO_948 (O_948,N_7221,N_6280);
or UO_949 (O_949,N_9748,N_5613);
or UO_950 (O_950,N_6626,N_8592);
xor UO_951 (O_951,N_8566,N_7681);
or UO_952 (O_952,N_9265,N_9999);
nand UO_953 (O_953,N_9907,N_6484);
nand UO_954 (O_954,N_8523,N_5705);
nor UO_955 (O_955,N_6338,N_8815);
and UO_956 (O_956,N_6947,N_7293);
or UO_957 (O_957,N_8916,N_5327);
nor UO_958 (O_958,N_9992,N_9301);
nand UO_959 (O_959,N_7231,N_8298);
nand UO_960 (O_960,N_8550,N_6597);
nand UO_961 (O_961,N_5149,N_8757);
nand UO_962 (O_962,N_6753,N_9342);
nand UO_963 (O_963,N_8459,N_6794);
xnor UO_964 (O_964,N_6464,N_8808);
or UO_965 (O_965,N_9977,N_7753);
nand UO_966 (O_966,N_8258,N_6757);
nand UO_967 (O_967,N_6362,N_8624);
xor UO_968 (O_968,N_5524,N_7522);
or UO_969 (O_969,N_6958,N_6806);
nor UO_970 (O_970,N_7756,N_5256);
nor UO_971 (O_971,N_5058,N_8354);
nand UO_972 (O_972,N_8841,N_9465);
nand UO_973 (O_973,N_5163,N_7431);
nand UO_974 (O_974,N_5611,N_7201);
nor UO_975 (O_975,N_9180,N_9431);
and UO_976 (O_976,N_5655,N_5145);
or UO_977 (O_977,N_6018,N_6447);
or UO_978 (O_978,N_9031,N_9281);
nor UO_979 (O_979,N_7300,N_7922);
nand UO_980 (O_980,N_6109,N_8556);
nand UO_981 (O_981,N_8377,N_5212);
nor UO_982 (O_982,N_5043,N_9026);
nor UO_983 (O_983,N_5551,N_5281);
or UO_984 (O_984,N_9290,N_6681);
or UO_985 (O_985,N_6841,N_5942);
nor UO_986 (O_986,N_5247,N_9550);
or UO_987 (O_987,N_6103,N_6045);
and UO_988 (O_988,N_6072,N_7317);
nor UO_989 (O_989,N_5792,N_5210);
xnor UO_990 (O_990,N_8797,N_9818);
nor UO_991 (O_991,N_8823,N_9976);
nor UO_992 (O_992,N_9953,N_5355);
nor UO_993 (O_993,N_8937,N_5005);
or UO_994 (O_994,N_8995,N_8066);
or UO_995 (O_995,N_5296,N_5739);
nor UO_996 (O_996,N_5573,N_9332);
nand UO_997 (O_997,N_9842,N_6114);
nor UO_998 (O_998,N_6746,N_5262);
or UO_999 (O_999,N_9401,N_5436);
nand UO_1000 (O_1000,N_5199,N_6055);
xnor UO_1001 (O_1001,N_5016,N_6209);
xnor UO_1002 (O_1002,N_8752,N_9941);
nor UO_1003 (O_1003,N_6080,N_6930);
nand UO_1004 (O_1004,N_5456,N_9571);
nor UO_1005 (O_1005,N_5943,N_6295);
or UO_1006 (O_1006,N_8059,N_5188);
xor UO_1007 (O_1007,N_7998,N_6967);
and UO_1008 (O_1008,N_7665,N_6443);
and UO_1009 (O_1009,N_5563,N_9745);
and UO_1010 (O_1010,N_7664,N_6836);
and UO_1011 (O_1011,N_6688,N_9158);
and UO_1012 (O_1012,N_8218,N_7807);
nor UO_1013 (O_1013,N_6905,N_8832);
or UO_1014 (O_1014,N_8722,N_9435);
and UO_1015 (O_1015,N_8534,N_6897);
xor UO_1016 (O_1016,N_7072,N_6720);
nor UO_1017 (O_1017,N_6774,N_8211);
or UO_1018 (O_1018,N_9727,N_9263);
nor UO_1019 (O_1019,N_5659,N_9266);
or UO_1020 (O_1020,N_9531,N_5181);
and UO_1021 (O_1021,N_9788,N_7433);
nor UO_1022 (O_1022,N_7337,N_5689);
nor UO_1023 (O_1023,N_5174,N_9716);
or UO_1024 (O_1024,N_7256,N_9085);
or UO_1025 (O_1025,N_6691,N_5080);
and UO_1026 (O_1026,N_5463,N_8409);
or UO_1027 (O_1027,N_9547,N_8019);
and UO_1028 (O_1028,N_8618,N_8110);
or UO_1029 (O_1029,N_6592,N_8597);
xnor UO_1030 (O_1030,N_6844,N_5126);
nand UO_1031 (O_1031,N_8421,N_9318);
or UO_1032 (O_1032,N_5216,N_5873);
nor UO_1033 (O_1033,N_7824,N_6010);
or UO_1034 (O_1034,N_6868,N_6334);
or UO_1035 (O_1035,N_7651,N_8897);
nor UO_1036 (O_1036,N_8914,N_7877);
xor UO_1037 (O_1037,N_7848,N_5462);
nor UO_1038 (O_1038,N_9178,N_9994);
and UO_1039 (O_1039,N_7145,N_8452);
nand UO_1040 (O_1040,N_6588,N_8848);
or UO_1041 (O_1041,N_5912,N_7815);
and UO_1042 (O_1042,N_7548,N_8740);
and UO_1043 (O_1043,N_7505,N_5245);
xor UO_1044 (O_1044,N_7275,N_9048);
and UO_1045 (O_1045,N_7067,N_9300);
nand UO_1046 (O_1046,N_5652,N_6736);
nand UO_1047 (O_1047,N_5972,N_9369);
and UO_1048 (O_1048,N_9469,N_5062);
or UO_1049 (O_1049,N_9995,N_5691);
nor UO_1050 (O_1050,N_6616,N_7593);
nand UO_1051 (O_1051,N_5610,N_7671);
or UO_1052 (O_1052,N_7680,N_5806);
xnor UO_1053 (O_1053,N_6047,N_9119);
nand UO_1054 (O_1054,N_6904,N_6116);
nor UO_1055 (O_1055,N_7562,N_9070);
and UO_1056 (O_1056,N_7098,N_8708);
nand UO_1057 (O_1057,N_7571,N_7897);
nand UO_1058 (O_1058,N_6596,N_6479);
xor UO_1059 (O_1059,N_8953,N_7460);
nand UO_1060 (O_1060,N_7082,N_5623);
and UO_1061 (O_1061,N_5619,N_6693);
or UO_1062 (O_1062,N_9713,N_5495);
nor UO_1063 (O_1063,N_8224,N_8479);
xor UO_1064 (O_1064,N_9739,N_5663);
nand UO_1065 (O_1065,N_6483,N_8487);
and UO_1066 (O_1066,N_5871,N_5639);
nand UO_1067 (O_1067,N_6563,N_7614);
nor UO_1068 (O_1068,N_9856,N_8639);
nor UO_1069 (O_1069,N_6326,N_6068);
and UO_1070 (O_1070,N_5786,N_5139);
nor UO_1071 (O_1071,N_7903,N_6171);
and UO_1072 (O_1072,N_6652,N_9227);
and UO_1073 (O_1073,N_5329,N_8095);
or UO_1074 (O_1074,N_6586,N_7531);
or UO_1075 (O_1075,N_6853,N_7860);
or UO_1076 (O_1076,N_5012,N_8985);
nand UO_1077 (O_1077,N_9826,N_7420);
nand UO_1078 (O_1078,N_6129,N_7196);
nor UO_1079 (O_1079,N_5002,N_7261);
and UO_1080 (O_1080,N_9873,N_8413);
or UO_1081 (O_1081,N_6718,N_6286);
nand UO_1082 (O_1082,N_7095,N_6002);
nor UO_1083 (O_1083,N_8314,N_5377);
nor UO_1084 (O_1084,N_8621,N_9565);
nor UO_1085 (O_1085,N_8115,N_6540);
and UO_1086 (O_1086,N_9718,N_8442);
and UO_1087 (O_1087,N_7994,N_5876);
nand UO_1088 (O_1088,N_8196,N_5899);
xor UO_1089 (O_1089,N_8249,N_9120);
nand UO_1090 (O_1090,N_9969,N_5337);
nor UO_1091 (O_1091,N_7604,N_5845);
and UO_1092 (O_1092,N_6128,N_5755);
nand UO_1093 (O_1093,N_6359,N_9053);
nand UO_1094 (O_1094,N_5874,N_8121);
nand UO_1095 (O_1095,N_6221,N_5402);
and UO_1096 (O_1096,N_5532,N_9673);
nand UO_1097 (O_1097,N_5714,N_6776);
or UO_1098 (O_1098,N_8701,N_6050);
nand UO_1099 (O_1099,N_5374,N_5641);
nand UO_1100 (O_1100,N_9474,N_6682);
xnor UO_1101 (O_1101,N_9535,N_8287);
nor UO_1102 (O_1102,N_6288,N_7572);
or UO_1103 (O_1103,N_8040,N_5520);
and UO_1104 (O_1104,N_6416,N_9753);
and UO_1105 (O_1105,N_5406,N_7198);
nor UO_1106 (O_1106,N_5308,N_6162);
nor UO_1107 (O_1107,N_8567,N_6756);
xor UO_1108 (O_1108,N_8684,N_9267);
xor UO_1109 (O_1109,N_7620,N_6191);
nand UO_1110 (O_1110,N_6706,N_7469);
or UO_1111 (O_1111,N_9127,N_6211);
nor UO_1112 (O_1112,N_8860,N_9923);
or UO_1113 (O_1113,N_6265,N_6215);
or UO_1114 (O_1114,N_9931,N_5765);
and UO_1115 (O_1115,N_5362,N_9478);
nand UO_1116 (O_1116,N_8758,N_6374);
or UO_1117 (O_1117,N_8792,N_5119);
nor UO_1118 (O_1118,N_9043,N_6053);
and UO_1119 (O_1119,N_9354,N_8939);
and UO_1120 (O_1120,N_6584,N_8251);
nand UO_1121 (O_1121,N_6769,N_5290);
or UO_1122 (O_1122,N_5725,N_7459);
nor UO_1123 (O_1123,N_7176,N_9172);
nand UO_1124 (O_1124,N_6287,N_6530);
nor UO_1125 (O_1125,N_5924,N_5458);
nor UO_1126 (O_1126,N_6124,N_6674);
or UO_1127 (O_1127,N_9125,N_9337);
and UO_1128 (O_1128,N_8400,N_5579);
nor UO_1129 (O_1129,N_8094,N_6946);
or UO_1130 (O_1130,N_6132,N_6982);
and UO_1131 (O_1131,N_6677,N_7639);
nand UO_1132 (O_1132,N_8077,N_6949);
nand UO_1133 (O_1133,N_8403,N_7032);
nand UO_1134 (O_1134,N_6651,N_6964);
nor UO_1135 (O_1135,N_5512,N_5665);
nand UO_1136 (O_1136,N_5018,N_8603);
or UO_1137 (O_1137,N_8307,N_7059);
nor UO_1138 (O_1138,N_9161,N_5991);
xnor UO_1139 (O_1139,N_9922,N_6556);
and UO_1140 (O_1140,N_6700,N_8671);
nor UO_1141 (O_1141,N_9804,N_5882);
nor UO_1142 (O_1142,N_8663,N_5046);
xor UO_1143 (O_1143,N_8232,N_7427);
nand UO_1144 (O_1144,N_6755,N_7850);
or UO_1145 (O_1145,N_9088,N_7580);
and UO_1146 (O_1146,N_5306,N_9388);
or UO_1147 (O_1147,N_7984,N_7403);
and UO_1148 (O_1148,N_5168,N_5156);
or UO_1149 (O_1149,N_7416,N_6005);
xnor UO_1150 (O_1150,N_5498,N_5164);
nor UO_1151 (O_1151,N_8552,N_5841);
nor UO_1152 (O_1152,N_7942,N_8488);
nor UO_1153 (O_1153,N_9800,N_6304);
or UO_1154 (O_1154,N_5273,N_8559);
or UO_1155 (O_1155,N_5475,N_8210);
and UO_1156 (O_1156,N_7863,N_5196);
nor UO_1157 (O_1157,N_5729,N_5364);
nor UO_1158 (O_1158,N_7634,N_5954);
nand UO_1159 (O_1159,N_8906,N_7870);
and UO_1160 (O_1160,N_5141,N_6472);
xnor UO_1161 (O_1161,N_5522,N_9860);
or UO_1162 (O_1162,N_7062,N_8448);
nor UO_1163 (O_1163,N_9759,N_7677);
and UO_1164 (O_1164,N_9709,N_7051);
or UO_1165 (O_1165,N_5863,N_9030);
nor UO_1166 (O_1166,N_6193,N_7707);
or UO_1167 (O_1167,N_6508,N_9116);
xnor UO_1168 (O_1168,N_7141,N_9364);
nand UO_1169 (O_1169,N_9011,N_9509);
and UO_1170 (O_1170,N_9051,N_8879);
nor UO_1171 (O_1171,N_7911,N_7599);
nand UO_1172 (O_1172,N_9951,N_8730);
xnor UO_1173 (O_1173,N_8578,N_8993);
xor UO_1174 (O_1174,N_6477,N_7710);
xnor UO_1175 (O_1175,N_8458,N_8158);
nand UO_1176 (O_1176,N_5769,N_8598);
nand UO_1177 (O_1177,N_7438,N_8023);
nand UO_1178 (O_1178,N_6467,N_8376);
nand UO_1179 (O_1179,N_9637,N_6603);
nor UO_1180 (O_1180,N_5297,N_6579);
nor UO_1181 (O_1181,N_9455,N_9927);
nor UO_1182 (O_1182,N_5948,N_9641);
nand UO_1183 (O_1183,N_8204,N_8818);
nand UO_1184 (O_1184,N_7515,N_5083);
nand UO_1185 (O_1185,N_9137,N_8161);
nor UO_1186 (O_1186,N_6708,N_8965);
and UO_1187 (O_1187,N_8637,N_5625);
and UO_1188 (O_1188,N_7696,N_7980);
and UO_1189 (O_1189,N_5395,N_7670);
or UO_1190 (O_1190,N_6127,N_7558);
and UO_1191 (O_1191,N_5205,N_5968);
nand UO_1192 (O_1192,N_5746,N_6360);
or UO_1193 (O_1193,N_9292,N_8418);
nor UO_1194 (O_1194,N_5602,N_9691);
nor UO_1195 (O_1195,N_8524,N_9499);
nor UO_1196 (O_1196,N_5267,N_7789);
and UO_1197 (O_1197,N_5258,N_9822);
and UO_1198 (O_1198,N_6619,N_9315);
or UO_1199 (O_1199,N_7606,N_5616);
nand UO_1200 (O_1200,N_6962,N_6418);
and UO_1201 (O_1201,N_8772,N_6824);
and UO_1202 (O_1202,N_8899,N_6709);
nor UO_1203 (O_1203,N_6976,N_5445);
and UO_1204 (O_1204,N_7243,N_6434);
or UO_1205 (O_1205,N_6306,N_5709);
nor UO_1206 (O_1206,N_6043,N_8748);
nor UO_1207 (O_1207,N_8008,N_7576);
xor UO_1208 (O_1208,N_9672,N_9134);
and UO_1209 (O_1209,N_6298,N_9096);
xnor UO_1210 (O_1210,N_7126,N_8886);
nand UO_1211 (O_1211,N_7917,N_7281);
or UO_1212 (O_1212,N_8919,N_5195);
nor UO_1213 (O_1213,N_6831,N_8682);
nor UO_1214 (O_1214,N_8568,N_7746);
nor UO_1215 (O_1215,N_9252,N_5510);
nor UO_1216 (O_1216,N_9805,N_6627);
or UO_1217 (O_1217,N_8775,N_7737);
or UO_1218 (O_1218,N_8753,N_9283);
nor UO_1219 (O_1219,N_5762,N_9954);
nand UO_1220 (O_1220,N_7885,N_9285);
nand UO_1221 (O_1221,N_7482,N_5905);
xnor UO_1222 (O_1222,N_8605,N_8600);
or UO_1223 (O_1223,N_6461,N_7351);
or UO_1224 (O_1224,N_5636,N_5666);
nor UO_1225 (O_1225,N_8374,N_6598);
and UO_1226 (O_1226,N_9365,N_7087);
xnor UO_1227 (O_1227,N_9255,N_7307);
xor UO_1228 (O_1228,N_7518,N_9577);
xor UO_1229 (O_1229,N_5457,N_8423);
nor UO_1230 (O_1230,N_9339,N_8446);
nor UO_1231 (O_1231,N_9696,N_5696);
nand UO_1232 (O_1232,N_6953,N_9857);
and UO_1233 (O_1233,N_8320,N_7524);
and UO_1234 (O_1234,N_9881,N_5836);
nor UO_1235 (O_1235,N_6816,N_9663);
nand UO_1236 (O_1236,N_5956,N_6895);
nand UO_1237 (O_1237,N_5173,N_9093);
and UO_1238 (O_1238,N_5986,N_9366);
nand UO_1239 (O_1239,N_8397,N_7269);
xnor UO_1240 (O_1240,N_9348,N_6234);
and UO_1241 (O_1241,N_7037,N_5880);
nand UO_1242 (O_1242,N_8401,N_8407);
or UO_1243 (O_1243,N_7116,N_8243);
nand UO_1244 (O_1244,N_5033,N_6713);
and UO_1245 (O_1245,N_9817,N_7024);
nand UO_1246 (O_1246,N_5011,N_7535);
and UO_1247 (O_1247,N_8736,N_9693);
nand UO_1248 (O_1248,N_5821,N_8264);
nand UO_1249 (O_1249,N_5872,N_9214);
nand UO_1250 (O_1250,N_6654,N_6159);
or UO_1251 (O_1251,N_7918,N_8006);
nor UO_1252 (O_1252,N_5670,N_7703);
and UO_1253 (O_1253,N_7400,N_7279);
or UO_1254 (O_1254,N_5206,N_6802);
and UO_1255 (O_1255,N_7500,N_6420);
and UO_1256 (O_1256,N_6327,N_9765);
nand UO_1257 (O_1257,N_8944,N_5676);
or UO_1258 (O_1258,N_5169,N_7557);
nand UO_1259 (O_1259,N_6168,N_7867);
nor UO_1260 (O_1260,N_5232,N_6033);
xnor UO_1261 (O_1261,N_5343,N_5497);
or UO_1262 (O_1262,N_9248,N_9707);
nor UO_1263 (O_1263,N_6862,N_5751);
nor UO_1264 (O_1264,N_5526,N_5519);
and UO_1265 (O_1265,N_5951,N_9430);
or UO_1266 (O_1266,N_9155,N_8087);
nor UO_1267 (O_1267,N_9209,N_5804);
and UO_1268 (O_1268,N_6469,N_7691);
and UO_1269 (O_1269,N_5453,N_9987);
nor UO_1270 (O_1270,N_5577,N_8014);
nor UO_1271 (O_1271,N_6960,N_8926);
nand UO_1272 (O_1272,N_9149,N_8239);
nor UO_1273 (O_1273,N_6308,N_5647);
nor UO_1274 (O_1274,N_9139,N_6425);
and UO_1275 (O_1275,N_7093,N_6888);
nand UO_1276 (O_1276,N_5988,N_8988);
and UO_1277 (O_1277,N_5934,N_6216);
and UO_1278 (O_1278,N_6729,N_8533);
and UO_1279 (O_1279,N_5349,N_9110);
nor UO_1280 (O_1280,N_6714,N_5885);
and UO_1281 (O_1281,N_8036,N_5528);
or UO_1282 (O_1282,N_8620,N_7481);
nor UO_1283 (O_1283,N_9567,N_7552);
nand UO_1284 (O_1284,N_8942,N_7318);
and UO_1285 (O_1285,N_8091,N_5581);
nand UO_1286 (O_1286,N_7423,N_6973);
nand UO_1287 (O_1287,N_5733,N_5552);
xor UO_1288 (O_1288,N_9894,N_9797);
or UO_1289 (O_1289,N_7321,N_9382);
nand UO_1290 (O_1290,N_7938,N_9489);
or UO_1291 (O_1291,N_5053,N_8664);
nand UO_1292 (O_1292,N_9165,N_5829);
nor UO_1293 (O_1293,N_5547,N_5066);
and UO_1294 (O_1294,N_7192,N_9963);
nor UO_1295 (O_1295,N_9750,N_8489);
or UO_1296 (O_1296,N_8352,N_5706);
or UO_1297 (O_1297,N_7060,N_5430);
and UO_1298 (O_1298,N_8076,N_6873);
nor UO_1299 (O_1299,N_9615,N_8471);
or UO_1300 (O_1300,N_5964,N_7407);
or UO_1301 (O_1301,N_6956,N_9925);
nor UO_1302 (O_1302,N_8890,N_8147);
and UO_1303 (O_1303,N_7276,N_9420);
or UO_1304 (O_1304,N_5862,N_6321);
nand UO_1305 (O_1305,N_7916,N_6343);
nor UO_1306 (O_1306,N_7819,N_6744);
and UO_1307 (O_1307,N_9518,N_9035);
or UO_1308 (O_1308,N_6212,N_6871);
nand UO_1309 (O_1309,N_5550,N_6970);
nor UO_1310 (O_1310,N_7601,N_5020);
and UO_1311 (O_1311,N_9612,N_8160);
and UO_1312 (O_1312,N_6696,N_8602);
nor UO_1313 (O_1313,N_5657,N_7085);
xor UO_1314 (O_1314,N_5932,N_7928);
nor UO_1315 (O_1315,N_5598,N_5047);
or UO_1316 (O_1316,N_8780,N_8010);
and UO_1317 (O_1317,N_8214,N_9956);
nand UO_1318 (O_1318,N_8531,N_5710);
nand UO_1319 (O_1319,N_7723,N_9831);
nor UO_1320 (O_1320,N_8315,N_6850);
xnor UO_1321 (O_1321,N_6752,N_7484);
nand UO_1322 (O_1322,N_9533,N_8884);
or UO_1323 (O_1323,N_8041,N_8484);
nor UO_1324 (O_1324,N_5576,N_7114);
and UO_1325 (O_1325,N_7134,N_9510);
nor UO_1326 (O_1326,N_6625,N_8625);
and UO_1327 (O_1327,N_7513,N_8954);
or UO_1328 (O_1328,N_9986,N_6455);
nor UO_1329 (O_1329,N_5301,N_9874);
xor UO_1330 (O_1330,N_8683,N_5811);
or UO_1331 (O_1331,N_6225,N_6346);
nor UO_1332 (O_1332,N_6959,N_7058);
or UO_1333 (O_1333,N_6680,N_8058);
nor UO_1334 (O_1334,N_8098,N_6277);
or UO_1335 (O_1335,N_7749,N_8128);
nor UO_1336 (O_1336,N_7719,N_7316);
nand UO_1337 (O_1337,N_7127,N_9330);
and UO_1338 (O_1338,N_5243,N_6707);
nor UO_1339 (O_1339,N_7040,N_9295);
nand UO_1340 (O_1340,N_9114,N_9991);
nand UO_1341 (O_1341,N_9427,N_6694);
or UO_1342 (O_1342,N_7694,N_9711);
and UO_1343 (O_1343,N_8404,N_5626);
or UO_1344 (O_1344,N_8217,N_6864);
nand UO_1345 (O_1345,N_8021,N_9417);
nor UO_1346 (O_1346,N_7567,N_9081);
and UO_1347 (O_1347,N_9024,N_5068);
nand UO_1348 (O_1348,N_8623,N_6121);
nand UO_1349 (O_1349,N_7200,N_8099);
nand UO_1350 (O_1350,N_9668,N_5989);
and UO_1351 (O_1351,N_5204,N_6843);
and UO_1352 (O_1352,N_5553,N_8466);
or UO_1353 (O_1353,N_8540,N_9917);
and UO_1354 (O_1354,N_6795,N_5992);
nand UO_1355 (O_1355,N_5484,N_6027);
nor UO_1356 (O_1356,N_7323,N_9377);
nor UO_1357 (O_1357,N_8029,N_5345);
or UO_1358 (O_1358,N_9308,N_9905);
nor UO_1359 (O_1359,N_6845,N_9503);
nand UO_1360 (O_1360,N_8237,N_7266);
and UO_1361 (O_1361,N_6239,N_9884);
nand UO_1362 (O_1362,N_5399,N_6320);
and UO_1363 (O_1363,N_7277,N_8892);
and UO_1364 (O_1364,N_8850,N_5467);
nand UO_1365 (O_1365,N_7913,N_8876);
nor UO_1366 (O_1366,N_5323,N_9109);
or UO_1367 (O_1367,N_7313,N_5496);
nand UO_1368 (O_1368,N_6643,N_5294);
nand UO_1369 (O_1369,N_9912,N_5490);
nand UO_1370 (O_1370,N_5086,N_7171);
nor UO_1371 (O_1371,N_8106,N_8505);
nor UO_1372 (O_1372,N_7380,N_9658);
nand UO_1373 (O_1373,N_7592,N_6955);
xor UO_1374 (O_1374,N_6968,N_7838);
xor UO_1375 (O_1375,N_6837,N_5771);
nor UO_1376 (O_1376,N_9883,N_8800);
or UO_1377 (O_1377,N_8086,N_9504);
and UO_1378 (O_1378,N_8958,N_7709);
nand UO_1379 (O_1379,N_6920,N_5103);
nand UO_1380 (O_1380,N_8869,N_9886);
nor UO_1381 (O_1381,N_7335,N_6550);
or UO_1382 (O_1382,N_8349,N_7393);
or UO_1383 (O_1383,N_5527,N_8714);
nand UO_1384 (O_1384,N_8480,N_9645);
or UO_1385 (O_1385,N_7740,N_5353);
nor UO_1386 (O_1386,N_6142,N_9493);
nor UO_1387 (O_1387,N_8265,N_5328);
nand UO_1388 (O_1388,N_9721,N_5415);
and UO_1389 (O_1389,N_5107,N_9740);
nor UO_1390 (O_1390,N_9827,N_9608);
or UO_1391 (O_1391,N_7825,N_7468);
nor UO_1392 (O_1392,N_9486,N_6092);
nor UO_1393 (O_1393,N_9761,N_7041);
xor UO_1394 (O_1394,N_9643,N_7443);
and UO_1395 (O_1395,N_6759,N_7932);
or UO_1396 (O_1396,N_9253,N_5917);
and UO_1397 (O_1397,N_7992,N_5071);
xor UO_1398 (O_1398,N_9223,N_7223);
or UO_1399 (O_1399,N_6354,N_6574);
nand UO_1400 (O_1400,N_5257,N_9064);
or UO_1401 (O_1401,N_8950,N_6712);
or UO_1402 (O_1402,N_7160,N_7426);
and UO_1403 (O_1403,N_8843,N_9397);
or UO_1404 (O_1404,N_8918,N_9112);
nand UO_1405 (O_1405,N_6615,N_9029);
nand UO_1406 (O_1406,N_9541,N_9915);
nor UO_1407 (O_1407,N_9238,N_7297);
nor UO_1408 (O_1408,N_6705,N_7411);
and UO_1409 (O_1409,N_7676,N_8867);
nor UO_1410 (O_1410,N_7048,N_8337);
and UO_1411 (O_1411,N_9549,N_7852);
nor UO_1412 (O_1412,N_6240,N_7770);
or UO_1413 (O_1413,N_9123,N_6781);
or UO_1414 (O_1414,N_5736,N_7180);
or UO_1415 (O_1415,N_5650,N_7751);
nand UO_1416 (O_1416,N_8709,N_5953);
and UO_1417 (O_1417,N_5901,N_7993);
and UO_1418 (O_1418,N_8816,N_6052);
or UO_1419 (O_1419,N_9561,N_8790);
or UO_1420 (O_1420,N_7285,N_6792);
and UO_1421 (O_1421,N_7900,N_5890);
xnor UO_1422 (O_1422,N_9424,N_5366);
and UO_1423 (O_1423,N_9568,N_6291);
or UO_1424 (O_1424,N_7536,N_8032);
nand UO_1425 (O_1425,N_8667,N_7315);
xor UO_1426 (O_1426,N_9310,N_7889);
and UO_1427 (O_1427,N_7865,N_8814);
xnor UO_1428 (O_1428,N_8108,N_7887);
or UO_1429 (O_1429,N_5386,N_7822);
nor UO_1430 (O_1430,N_8216,N_8350);
and UO_1431 (O_1431,N_5000,N_5961);
xnor UO_1432 (O_1432,N_7583,N_8665);
xnor UO_1433 (O_1433,N_8875,N_6113);
nor UO_1434 (O_1434,N_9436,N_6478);
and UO_1435 (O_1435,N_7084,N_6948);
and UO_1436 (O_1436,N_6639,N_8429);
and UO_1437 (O_1437,N_5372,N_9046);
nand UO_1438 (O_1438,N_7125,N_5272);
or UO_1439 (O_1439,N_8432,N_6599);
or UO_1440 (O_1440,N_8971,N_8998);
nor UO_1441 (O_1441,N_5627,N_7167);
or UO_1442 (O_1442,N_7365,N_9221);
nand UO_1443 (O_1443,N_7527,N_8666);
xor UO_1444 (O_1444,N_8601,N_9511);
and UO_1445 (O_1445,N_8193,N_9613);
nand UO_1446 (O_1446,N_9476,N_5797);
nand UO_1447 (O_1447,N_9439,N_6761);
nand UO_1448 (O_1448,N_5070,N_5274);
and UO_1449 (O_1449,N_5183,N_7818);
nor UO_1450 (O_1450,N_8405,N_6631);
nand UO_1451 (O_1451,N_5443,N_6390);
and UO_1452 (O_1452,N_6301,N_5161);
xnor UO_1453 (O_1453,N_9067,N_5087);
nand UO_1454 (O_1454,N_5468,N_8854);
or UO_1455 (O_1455,N_5814,N_8861);
xnor UO_1456 (O_1456,N_5826,N_7345);
xor UO_1457 (O_1457,N_6786,N_8996);
nand UO_1458 (O_1458,N_5129,N_8343);
nor UO_1459 (O_1459,N_6885,N_8851);
or UO_1460 (O_1460,N_6668,N_9708);
and UO_1461 (O_1461,N_6780,N_5095);
or UO_1462 (O_1462,N_5668,N_9699);
or UO_1463 (O_1463,N_6063,N_5029);
and UO_1464 (O_1464,N_8628,N_8657);
nand UO_1465 (O_1465,N_8425,N_5044);
nand UO_1466 (O_1466,N_7906,N_7660);
nor UO_1467 (O_1467,N_6702,N_6567);
and UO_1468 (O_1468,N_9061,N_5772);
and UO_1469 (O_1469,N_5678,N_7146);
and UO_1470 (O_1470,N_7090,N_7241);
xor UO_1471 (O_1471,N_7793,N_5504);
xor UO_1472 (O_1472,N_6611,N_7450);
or UO_1473 (O_1473,N_9793,N_9682);
nor UO_1474 (O_1474,N_9133,N_5114);
nor UO_1475 (O_1475,N_6815,N_9724);
nand UO_1476 (O_1476,N_8414,N_6545);
xor UO_1477 (O_1477,N_7260,N_8539);
nand UO_1478 (O_1478,N_7080,N_9203);
nand UO_1479 (O_1479,N_7480,N_8681);
and UO_1480 (O_1480,N_6541,N_6026);
nand UO_1481 (O_1481,N_5542,N_9984);
nand UO_1482 (O_1482,N_6296,N_6356);
or UO_1483 (O_1483,N_5405,N_8172);
or UO_1484 (O_1484,N_8501,N_7486);
nand UO_1485 (O_1485,N_7398,N_9142);
nor UO_1486 (O_1486,N_7257,N_7509);
or UO_1487 (O_1487,N_8829,N_8999);
and UO_1488 (O_1488,N_8812,N_7334);
or UO_1489 (O_1489,N_9235,N_9428);
nor UO_1490 (O_1490,N_9082,N_8599);
or UO_1491 (O_1491,N_6032,N_9878);
or UO_1492 (O_1492,N_7474,N_7204);
or UO_1493 (O_1493,N_6219,N_7834);
and UO_1494 (O_1494,N_6860,N_9411);
nand UO_1495 (O_1495,N_7569,N_6922);
and UO_1496 (O_1496,N_6690,N_7475);
and UO_1497 (O_1497,N_5981,N_8847);
xor UO_1498 (O_1498,N_7181,N_9261);
nand UO_1499 (O_1499,N_9390,N_6223);
endmodule