module basic_500_3000_500_5_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_283,In_472);
and U1 (N_1,In_272,In_124);
xor U2 (N_2,In_216,In_46);
and U3 (N_3,In_366,In_249);
nor U4 (N_4,In_68,In_378);
nand U5 (N_5,In_374,In_128);
or U6 (N_6,In_165,In_463);
or U7 (N_7,In_112,In_239);
nand U8 (N_8,In_144,In_414);
nor U9 (N_9,In_85,In_231);
nand U10 (N_10,In_134,In_400);
and U11 (N_11,In_492,In_417);
xor U12 (N_12,In_9,In_304);
xnor U13 (N_13,In_111,In_191);
xnor U14 (N_14,In_260,In_259);
or U15 (N_15,In_172,In_393);
nor U16 (N_16,In_127,In_353);
nor U17 (N_17,In_448,In_402);
nor U18 (N_18,In_13,In_299);
xor U19 (N_19,In_334,In_237);
nor U20 (N_20,In_145,In_398);
xor U21 (N_21,In_479,In_242);
or U22 (N_22,In_88,In_498);
xnor U23 (N_23,In_80,In_411);
nand U24 (N_24,In_291,In_177);
or U25 (N_25,In_332,In_303);
xnor U26 (N_26,In_371,In_485);
or U27 (N_27,In_254,In_157);
or U28 (N_28,In_248,In_445);
nor U29 (N_29,In_358,In_63);
xnor U30 (N_30,In_108,In_208);
and U31 (N_31,In_136,In_269);
nor U32 (N_32,In_125,In_186);
xor U33 (N_33,In_34,In_188);
nor U34 (N_34,In_52,In_71);
nor U35 (N_35,In_11,In_430);
and U36 (N_36,In_65,In_152);
nand U37 (N_37,In_390,In_48);
and U38 (N_38,In_481,In_432);
nand U39 (N_39,In_121,In_78);
nand U40 (N_40,In_97,In_28);
or U41 (N_41,In_343,In_7);
nand U42 (N_42,In_360,In_351);
nand U43 (N_43,In_204,In_91);
nor U44 (N_44,In_163,In_412);
nand U45 (N_45,In_89,In_298);
or U46 (N_46,In_368,In_5);
nor U47 (N_47,In_122,In_442);
xor U48 (N_48,In_262,In_40);
and U49 (N_49,In_168,In_16);
xor U50 (N_50,In_422,In_369);
and U51 (N_51,In_126,In_420);
nand U52 (N_52,In_310,In_483);
and U53 (N_53,In_264,In_350);
and U54 (N_54,In_362,In_293);
or U55 (N_55,In_167,In_473);
and U56 (N_56,In_314,In_154);
and U57 (N_57,In_21,In_289);
and U58 (N_58,In_395,In_123);
nand U59 (N_59,In_443,In_426);
xnor U60 (N_60,In_263,In_215);
or U61 (N_61,In_403,In_45);
nand U62 (N_62,In_312,In_107);
xnor U63 (N_63,In_458,In_243);
or U64 (N_64,In_328,In_138);
nor U65 (N_65,In_4,In_20);
nand U66 (N_66,In_176,In_33);
and U67 (N_67,In_399,In_337);
nor U68 (N_68,In_118,In_179);
or U69 (N_69,In_278,In_211);
nand U70 (N_70,In_363,In_212);
or U71 (N_71,In_347,In_170);
nand U72 (N_72,In_257,In_409);
and U73 (N_73,In_252,In_120);
nand U74 (N_74,In_316,In_244);
and U75 (N_75,In_77,In_427);
nor U76 (N_76,In_413,In_275);
nor U77 (N_77,In_460,In_42);
xor U78 (N_78,In_301,In_333);
nand U79 (N_79,In_18,In_296);
nor U80 (N_80,In_58,In_62);
or U81 (N_81,In_189,In_342);
and U82 (N_82,In_221,In_192);
or U83 (N_83,In_159,In_140);
or U84 (N_84,In_394,In_218);
nand U85 (N_85,In_285,In_341);
xor U86 (N_86,In_266,In_461);
and U87 (N_87,In_219,In_149);
or U88 (N_88,In_475,In_323);
nand U89 (N_89,In_217,In_17);
nor U90 (N_90,In_200,In_339);
nand U91 (N_91,In_222,In_317);
nor U92 (N_92,In_396,In_183);
nand U93 (N_93,In_100,In_130);
nor U94 (N_94,In_169,In_146);
nor U95 (N_95,In_173,In_383);
or U96 (N_96,In_178,In_372);
nand U97 (N_97,In_320,In_84);
nor U98 (N_98,In_497,In_25);
nand U99 (N_99,In_101,In_180);
nand U100 (N_100,In_379,In_478);
or U101 (N_101,In_327,In_205);
or U102 (N_102,In_365,In_69);
and U103 (N_103,In_37,In_86);
nand U104 (N_104,In_367,In_181);
and U105 (N_105,In_446,In_452);
or U106 (N_106,In_486,In_324);
xnor U107 (N_107,In_424,In_29);
nor U108 (N_108,In_82,In_119);
xor U109 (N_109,In_114,In_253);
xnor U110 (N_110,In_433,In_199);
or U111 (N_111,In_19,In_35);
and U112 (N_112,In_440,In_117);
nand U113 (N_113,In_274,In_41);
nor U114 (N_114,In_466,In_354);
or U115 (N_115,In_437,In_271);
xnor U116 (N_116,In_421,In_110);
or U117 (N_117,In_387,In_132);
nor U118 (N_118,In_284,In_76);
nand U119 (N_119,In_464,In_210);
nand U120 (N_120,In_160,In_364);
or U121 (N_121,In_313,In_105);
and U122 (N_122,In_0,In_292);
or U123 (N_123,In_225,In_280);
nor U124 (N_124,In_93,In_309);
nand U125 (N_125,In_406,In_295);
and U126 (N_126,In_397,In_357);
or U127 (N_127,In_197,In_490);
or U128 (N_128,In_36,In_220);
or U129 (N_129,In_330,In_151);
xnor U130 (N_130,In_336,In_75);
nor U131 (N_131,In_175,In_270);
and U132 (N_132,In_213,In_6);
and U133 (N_133,In_235,In_102);
nor U134 (N_134,In_61,In_147);
nor U135 (N_135,In_8,In_247);
and U136 (N_136,In_451,In_245);
and U137 (N_137,In_288,In_407);
nor U138 (N_138,In_322,In_106);
xor U139 (N_139,In_53,In_373);
xnor U140 (N_140,In_315,In_290);
xnor U141 (N_141,In_321,In_480);
or U142 (N_142,In_202,In_92);
nor U143 (N_143,In_455,In_447);
and U144 (N_144,In_352,In_67);
nor U145 (N_145,In_116,In_43);
and U146 (N_146,In_462,In_457);
or U147 (N_147,In_318,In_73);
or U148 (N_148,In_143,In_64);
nand U149 (N_149,In_26,In_223);
nand U150 (N_150,In_431,In_329);
and U151 (N_151,In_236,In_227);
nor U152 (N_152,In_345,In_156);
and U153 (N_153,In_12,In_187);
and U154 (N_154,In_429,In_161);
nand U155 (N_155,In_190,In_418);
or U156 (N_156,In_171,In_94);
xnor U157 (N_157,In_150,In_384);
nor U158 (N_158,In_109,In_1);
and U159 (N_159,In_496,In_453);
or U160 (N_160,In_467,In_95);
xor U161 (N_161,In_404,In_361);
nor U162 (N_162,In_488,In_99);
nand U163 (N_163,In_182,In_349);
or U164 (N_164,In_148,In_70);
nor U165 (N_165,In_87,In_238);
nor U166 (N_166,In_129,In_459);
nor U167 (N_167,In_325,In_436);
nand U168 (N_168,In_196,In_47);
nor U169 (N_169,In_135,In_335);
nand U170 (N_170,In_276,In_306);
xor U171 (N_171,In_392,In_27);
nand U172 (N_172,In_308,In_438);
and U173 (N_173,In_38,In_50);
nor U174 (N_174,In_450,In_224);
and U175 (N_175,In_194,In_305);
nand U176 (N_176,In_319,In_340);
or U177 (N_177,In_302,In_137);
and U178 (N_178,In_142,In_465);
xor U179 (N_179,In_230,In_493);
xnor U180 (N_180,In_434,In_277);
or U181 (N_181,In_233,In_206);
and U182 (N_182,In_416,In_391);
nand U183 (N_183,In_311,In_201);
xor U184 (N_184,In_229,In_435);
nor U185 (N_185,In_24,In_265);
nor U186 (N_186,In_386,In_2);
and U187 (N_187,In_441,In_198);
nor U188 (N_188,In_477,In_256);
nor U189 (N_189,In_56,In_408);
or U190 (N_190,In_419,In_22);
nor U191 (N_191,In_49,In_471);
and U192 (N_192,In_193,In_476);
nor U193 (N_193,In_487,In_428);
nand U194 (N_194,In_258,In_72);
xnor U195 (N_195,In_267,In_331);
nor U196 (N_196,In_282,In_57);
nor U197 (N_197,In_226,In_251);
nand U198 (N_198,In_44,In_166);
nand U199 (N_199,In_415,In_232);
and U200 (N_200,In_185,In_444);
nand U201 (N_201,In_23,In_81);
nor U202 (N_202,In_158,In_385);
nand U203 (N_203,In_74,In_439);
and U204 (N_204,In_405,In_389);
and U205 (N_205,In_98,In_494);
and U206 (N_206,In_113,In_207);
nor U207 (N_207,In_32,In_10);
or U208 (N_208,In_90,In_484);
or U209 (N_209,In_240,In_83);
or U210 (N_210,In_255,In_401);
nor U211 (N_211,In_184,In_54);
nor U212 (N_212,In_30,In_96);
nor U213 (N_213,In_470,In_356);
nand U214 (N_214,In_449,In_468);
and U215 (N_215,In_344,In_326);
nand U216 (N_216,In_456,In_14);
or U217 (N_217,In_499,In_307);
nor U218 (N_218,In_103,In_115);
xnor U219 (N_219,In_382,In_59);
nor U220 (N_220,In_162,In_174);
or U221 (N_221,In_155,In_51);
xnor U222 (N_222,In_246,In_195);
nand U223 (N_223,In_300,In_141);
nor U224 (N_224,In_286,In_268);
or U225 (N_225,In_153,In_474);
nand U226 (N_226,In_491,In_410);
or U227 (N_227,In_250,In_228);
or U228 (N_228,In_15,In_375);
nand U229 (N_229,In_377,In_423);
nand U230 (N_230,In_454,In_489);
or U231 (N_231,In_273,In_380);
nand U232 (N_232,In_60,In_359);
or U233 (N_233,In_469,In_294);
or U234 (N_234,In_79,In_31);
nor U235 (N_235,In_241,In_55);
nor U236 (N_236,In_164,In_482);
or U237 (N_237,In_279,In_139);
and U238 (N_238,In_376,In_425);
nor U239 (N_239,In_209,In_39);
or U240 (N_240,In_355,In_131);
and U241 (N_241,In_66,In_348);
nor U242 (N_242,In_381,In_133);
and U243 (N_243,In_495,In_3);
and U244 (N_244,In_388,In_338);
xnor U245 (N_245,In_261,In_370);
or U246 (N_246,In_297,In_287);
nand U247 (N_247,In_104,In_214);
nor U248 (N_248,In_203,In_346);
nor U249 (N_249,In_234,In_281);
and U250 (N_250,In_50,In_200);
nand U251 (N_251,In_242,In_148);
or U252 (N_252,In_330,In_47);
nand U253 (N_253,In_230,In_208);
or U254 (N_254,In_103,In_297);
nor U255 (N_255,In_64,In_449);
and U256 (N_256,In_373,In_275);
nand U257 (N_257,In_241,In_149);
and U258 (N_258,In_283,In_338);
nand U259 (N_259,In_41,In_280);
or U260 (N_260,In_3,In_171);
and U261 (N_261,In_400,In_408);
and U262 (N_262,In_136,In_491);
and U263 (N_263,In_296,In_85);
and U264 (N_264,In_208,In_75);
nor U265 (N_265,In_248,In_307);
or U266 (N_266,In_216,In_492);
xor U267 (N_267,In_216,In_434);
nor U268 (N_268,In_410,In_199);
xnor U269 (N_269,In_142,In_217);
or U270 (N_270,In_416,In_405);
and U271 (N_271,In_400,In_362);
nor U272 (N_272,In_379,In_313);
nand U273 (N_273,In_483,In_393);
xor U274 (N_274,In_305,In_20);
nor U275 (N_275,In_342,In_294);
nor U276 (N_276,In_486,In_428);
or U277 (N_277,In_84,In_302);
and U278 (N_278,In_94,In_216);
and U279 (N_279,In_204,In_81);
nor U280 (N_280,In_6,In_386);
or U281 (N_281,In_499,In_206);
and U282 (N_282,In_298,In_325);
or U283 (N_283,In_458,In_18);
or U284 (N_284,In_80,In_281);
or U285 (N_285,In_135,In_347);
nor U286 (N_286,In_176,In_397);
nand U287 (N_287,In_434,In_391);
and U288 (N_288,In_306,In_138);
xnor U289 (N_289,In_396,In_34);
or U290 (N_290,In_450,In_53);
or U291 (N_291,In_314,In_443);
and U292 (N_292,In_164,In_429);
nand U293 (N_293,In_477,In_230);
nand U294 (N_294,In_140,In_257);
and U295 (N_295,In_27,In_282);
nor U296 (N_296,In_70,In_162);
and U297 (N_297,In_282,In_242);
xor U298 (N_298,In_69,In_400);
xnor U299 (N_299,In_24,In_397);
nand U300 (N_300,In_25,In_184);
and U301 (N_301,In_164,In_300);
and U302 (N_302,In_76,In_325);
nand U303 (N_303,In_86,In_11);
or U304 (N_304,In_34,In_104);
nand U305 (N_305,In_92,In_475);
or U306 (N_306,In_234,In_173);
xnor U307 (N_307,In_259,In_357);
nand U308 (N_308,In_316,In_30);
nand U309 (N_309,In_29,In_400);
or U310 (N_310,In_422,In_428);
or U311 (N_311,In_258,In_415);
and U312 (N_312,In_91,In_257);
nand U313 (N_313,In_489,In_299);
nor U314 (N_314,In_165,In_260);
xor U315 (N_315,In_156,In_96);
xor U316 (N_316,In_145,In_276);
nand U317 (N_317,In_216,In_237);
nand U318 (N_318,In_386,In_66);
and U319 (N_319,In_378,In_100);
nand U320 (N_320,In_159,In_432);
nor U321 (N_321,In_267,In_193);
or U322 (N_322,In_362,In_84);
or U323 (N_323,In_345,In_331);
or U324 (N_324,In_225,In_327);
nand U325 (N_325,In_151,In_67);
xor U326 (N_326,In_185,In_141);
xor U327 (N_327,In_334,In_402);
nor U328 (N_328,In_66,In_215);
nor U329 (N_329,In_334,In_158);
nand U330 (N_330,In_190,In_368);
nand U331 (N_331,In_204,In_102);
xor U332 (N_332,In_65,In_457);
nor U333 (N_333,In_477,In_157);
nor U334 (N_334,In_472,In_202);
or U335 (N_335,In_29,In_376);
nor U336 (N_336,In_197,In_47);
and U337 (N_337,In_134,In_230);
or U338 (N_338,In_197,In_89);
xor U339 (N_339,In_242,In_212);
nand U340 (N_340,In_23,In_315);
xor U341 (N_341,In_104,In_423);
xor U342 (N_342,In_451,In_466);
and U343 (N_343,In_254,In_48);
xnor U344 (N_344,In_248,In_441);
xor U345 (N_345,In_167,In_417);
nand U346 (N_346,In_98,In_110);
or U347 (N_347,In_333,In_463);
and U348 (N_348,In_418,In_106);
and U349 (N_349,In_493,In_42);
xor U350 (N_350,In_155,In_232);
nand U351 (N_351,In_187,In_459);
or U352 (N_352,In_387,In_92);
nor U353 (N_353,In_349,In_365);
or U354 (N_354,In_177,In_409);
and U355 (N_355,In_193,In_340);
xor U356 (N_356,In_2,In_354);
or U357 (N_357,In_360,In_357);
nand U358 (N_358,In_105,In_489);
nand U359 (N_359,In_428,In_430);
nand U360 (N_360,In_3,In_313);
nor U361 (N_361,In_230,In_138);
and U362 (N_362,In_198,In_115);
xnor U363 (N_363,In_4,In_362);
nor U364 (N_364,In_238,In_69);
or U365 (N_365,In_488,In_478);
xor U366 (N_366,In_126,In_368);
nor U367 (N_367,In_166,In_378);
xnor U368 (N_368,In_378,In_271);
or U369 (N_369,In_294,In_31);
nand U370 (N_370,In_15,In_49);
and U371 (N_371,In_399,In_266);
nor U372 (N_372,In_124,In_0);
and U373 (N_373,In_368,In_198);
and U374 (N_374,In_463,In_420);
nand U375 (N_375,In_42,In_431);
nor U376 (N_376,In_12,In_428);
nand U377 (N_377,In_363,In_484);
nor U378 (N_378,In_106,In_408);
nand U379 (N_379,In_462,In_88);
and U380 (N_380,In_73,In_292);
nor U381 (N_381,In_405,In_409);
and U382 (N_382,In_397,In_41);
or U383 (N_383,In_329,In_323);
or U384 (N_384,In_270,In_435);
and U385 (N_385,In_240,In_20);
and U386 (N_386,In_462,In_295);
nor U387 (N_387,In_244,In_365);
nor U388 (N_388,In_100,In_249);
or U389 (N_389,In_494,In_443);
or U390 (N_390,In_384,In_314);
xor U391 (N_391,In_99,In_213);
xnor U392 (N_392,In_188,In_351);
nor U393 (N_393,In_394,In_413);
and U394 (N_394,In_409,In_255);
nand U395 (N_395,In_80,In_223);
nand U396 (N_396,In_61,In_170);
nor U397 (N_397,In_163,In_71);
or U398 (N_398,In_257,In_386);
or U399 (N_399,In_182,In_329);
nor U400 (N_400,In_450,In_221);
and U401 (N_401,In_8,In_191);
nor U402 (N_402,In_336,In_13);
nor U403 (N_403,In_85,In_318);
or U404 (N_404,In_68,In_96);
nor U405 (N_405,In_43,In_218);
nand U406 (N_406,In_307,In_0);
xor U407 (N_407,In_400,In_253);
nor U408 (N_408,In_207,In_478);
nor U409 (N_409,In_174,In_26);
nand U410 (N_410,In_373,In_177);
and U411 (N_411,In_297,In_54);
nand U412 (N_412,In_240,In_222);
nor U413 (N_413,In_57,In_333);
nor U414 (N_414,In_289,In_238);
xor U415 (N_415,In_138,In_47);
and U416 (N_416,In_31,In_99);
and U417 (N_417,In_16,In_482);
nor U418 (N_418,In_241,In_48);
nand U419 (N_419,In_246,In_120);
and U420 (N_420,In_170,In_340);
and U421 (N_421,In_124,In_137);
nor U422 (N_422,In_124,In_27);
xor U423 (N_423,In_379,In_344);
nor U424 (N_424,In_222,In_287);
and U425 (N_425,In_329,In_222);
and U426 (N_426,In_195,In_1);
xor U427 (N_427,In_496,In_46);
xnor U428 (N_428,In_487,In_237);
or U429 (N_429,In_240,In_141);
and U430 (N_430,In_274,In_474);
or U431 (N_431,In_39,In_84);
or U432 (N_432,In_48,In_293);
and U433 (N_433,In_216,In_172);
or U434 (N_434,In_253,In_160);
or U435 (N_435,In_334,In_289);
and U436 (N_436,In_171,In_462);
nor U437 (N_437,In_217,In_345);
and U438 (N_438,In_254,In_289);
nand U439 (N_439,In_246,In_86);
or U440 (N_440,In_70,In_451);
nand U441 (N_441,In_73,In_468);
nand U442 (N_442,In_390,In_178);
xor U443 (N_443,In_279,In_446);
and U444 (N_444,In_219,In_321);
nand U445 (N_445,In_163,In_80);
nor U446 (N_446,In_62,In_263);
nor U447 (N_447,In_310,In_249);
nor U448 (N_448,In_410,In_68);
nor U449 (N_449,In_4,In_90);
or U450 (N_450,In_146,In_0);
nand U451 (N_451,In_462,In_240);
or U452 (N_452,In_378,In_459);
nand U453 (N_453,In_12,In_475);
and U454 (N_454,In_111,In_221);
nand U455 (N_455,In_389,In_123);
and U456 (N_456,In_344,In_9);
and U457 (N_457,In_85,In_488);
nor U458 (N_458,In_205,In_443);
and U459 (N_459,In_383,In_254);
and U460 (N_460,In_257,In_233);
and U461 (N_461,In_217,In_170);
or U462 (N_462,In_457,In_300);
or U463 (N_463,In_227,In_418);
or U464 (N_464,In_66,In_431);
nand U465 (N_465,In_441,In_485);
nor U466 (N_466,In_172,In_418);
and U467 (N_467,In_448,In_403);
or U468 (N_468,In_325,In_276);
nand U469 (N_469,In_436,In_248);
and U470 (N_470,In_465,In_191);
nor U471 (N_471,In_92,In_439);
and U472 (N_472,In_483,In_158);
nor U473 (N_473,In_39,In_496);
nor U474 (N_474,In_443,In_92);
nor U475 (N_475,In_232,In_366);
xnor U476 (N_476,In_469,In_439);
or U477 (N_477,In_283,In_112);
nand U478 (N_478,In_135,In_11);
nand U479 (N_479,In_356,In_83);
and U480 (N_480,In_138,In_299);
and U481 (N_481,In_196,In_97);
nor U482 (N_482,In_358,In_367);
nand U483 (N_483,In_90,In_242);
and U484 (N_484,In_243,In_67);
nor U485 (N_485,In_10,In_446);
or U486 (N_486,In_326,In_88);
and U487 (N_487,In_450,In_185);
nand U488 (N_488,In_210,In_376);
and U489 (N_489,In_188,In_219);
nand U490 (N_490,In_342,In_245);
or U491 (N_491,In_287,In_141);
nor U492 (N_492,In_292,In_161);
xnor U493 (N_493,In_327,In_497);
xor U494 (N_494,In_150,In_53);
nor U495 (N_495,In_249,In_463);
and U496 (N_496,In_479,In_304);
nand U497 (N_497,In_242,In_413);
nor U498 (N_498,In_321,In_369);
nor U499 (N_499,In_149,In_260);
nand U500 (N_500,In_330,In_391);
or U501 (N_501,In_415,In_436);
nand U502 (N_502,In_279,In_119);
or U503 (N_503,In_15,In_121);
or U504 (N_504,In_227,In_9);
nand U505 (N_505,In_142,In_327);
and U506 (N_506,In_246,In_176);
xnor U507 (N_507,In_448,In_222);
nor U508 (N_508,In_94,In_6);
nor U509 (N_509,In_267,In_59);
nor U510 (N_510,In_86,In_364);
nor U511 (N_511,In_184,In_487);
and U512 (N_512,In_286,In_200);
and U513 (N_513,In_171,In_280);
nor U514 (N_514,In_296,In_52);
nor U515 (N_515,In_259,In_426);
and U516 (N_516,In_380,In_231);
nand U517 (N_517,In_367,In_377);
xnor U518 (N_518,In_192,In_369);
nor U519 (N_519,In_282,In_462);
xnor U520 (N_520,In_356,In_258);
or U521 (N_521,In_461,In_230);
and U522 (N_522,In_224,In_251);
or U523 (N_523,In_152,In_99);
xor U524 (N_524,In_373,In_127);
and U525 (N_525,In_236,In_288);
nand U526 (N_526,In_260,In_339);
nor U527 (N_527,In_54,In_43);
and U528 (N_528,In_176,In_319);
nand U529 (N_529,In_318,In_480);
nor U530 (N_530,In_236,In_305);
nand U531 (N_531,In_103,In_237);
nand U532 (N_532,In_208,In_130);
nand U533 (N_533,In_330,In_387);
nor U534 (N_534,In_361,In_269);
and U535 (N_535,In_87,In_465);
nor U536 (N_536,In_334,In_374);
xor U537 (N_537,In_486,In_288);
nor U538 (N_538,In_17,In_224);
nor U539 (N_539,In_304,In_287);
nand U540 (N_540,In_297,In_331);
nand U541 (N_541,In_311,In_453);
nor U542 (N_542,In_136,In_391);
or U543 (N_543,In_295,In_244);
or U544 (N_544,In_229,In_432);
or U545 (N_545,In_424,In_335);
and U546 (N_546,In_198,In_450);
or U547 (N_547,In_334,In_225);
and U548 (N_548,In_44,In_202);
or U549 (N_549,In_364,In_20);
nand U550 (N_550,In_104,In_481);
and U551 (N_551,In_109,In_242);
or U552 (N_552,In_56,In_110);
nand U553 (N_553,In_172,In_95);
and U554 (N_554,In_19,In_36);
nor U555 (N_555,In_160,In_98);
and U556 (N_556,In_71,In_469);
or U557 (N_557,In_217,In_339);
and U558 (N_558,In_179,In_180);
nand U559 (N_559,In_374,In_367);
and U560 (N_560,In_417,In_205);
xnor U561 (N_561,In_236,In_31);
or U562 (N_562,In_133,In_254);
nor U563 (N_563,In_483,In_372);
nor U564 (N_564,In_122,In_302);
and U565 (N_565,In_72,In_78);
nor U566 (N_566,In_331,In_23);
and U567 (N_567,In_419,In_168);
and U568 (N_568,In_354,In_339);
and U569 (N_569,In_343,In_137);
or U570 (N_570,In_287,In_241);
nand U571 (N_571,In_359,In_246);
or U572 (N_572,In_326,In_69);
xor U573 (N_573,In_47,In_181);
nor U574 (N_574,In_145,In_258);
and U575 (N_575,In_2,In_270);
nor U576 (N_576,In_122,In_164);
nor U577 (N_577,In_39,In_47);
or U578 (N_578,In_154,In_181);
nor U579 (N_579,In_417,In_296);
or U580 (N_580,In_242,In_98);
nor U581 (N_581,In_358,In_103);
or U582 (N_582,In_162,In_66);
and U583 (N_583,In_385,In_157);
xor U584 (N_584,In_170,In_311);
or U585 (N_585,In_101,In_494);
and U586 (N_586,In_153,In_283);
and U587 (N_587,In_440,In_16);
nand U588 (N_588,In_412,In_367);
and U589 (N_589,In_448,In_382);
xnor U590 (N_590,In_433,In_269);
and U591 (N_591,In_125,In_120);
nor U592 (N_592,In_443,In_1);
nor U593 (N_593,In_352,In_477);
nor U594 (N_594,In_422,In_353);
nand U595 (N_595,In_181,In_159);
nor U596 (N_596,In_460,In_8);
and U597 (N_597,In_244,In_411);
nor U598 (N_598,In_446,In_243);
nand U599 (N_599,In_210,In_233);
and U600 (N_600,N_90,N_294);
xnor U601 (N_601,N_388,N_214);
or U602 (N_602,N_217,N_31);
nand U603 (N_603,N_160,N_560);
nand U604 (N_604,N_448,N_304);
and U605 (N_605,N_244,N_377);
or U606 (N_606,N_513,N_189);
or U607 (N_607,N_485,N_148);
nand U608 (N_608,N_393,N_322);
nand U609 (N_609,N_536,N_463);
xor U610 (N_610,N_265,N_120);
nand U611 (N_611,N_79,N_517);
or U612 (N_612,N_230,N_250);
or U613 (N_613,N_238,N_30);
nor U614 (N_614,N_60,N_395);
nand U615 (N_615,N_49,N_42);
xor U616 (N_616,N_479,N_38);
nor U617 (N_617,N_121,N_260);
nand U618 (N_618,N_234,N_391);
nand U619 (N_619,N_241,N_180);
or U620 (N_620,N_23,N_19);
xnor U621 (N_621,N_209,N_116);
or U622 (N_622,N_439,N_429);
and U623 (N_623,N_452,N_422);
nor U624 (N_624,N_298,N_101);
nand U625 (N_625,N_80,N_596);
and U626 (N_626,N_108,N_586);
nand U627 (N_627,N_208,N_53);
nor U628 (N_628,N_130,N_346);
xnor U629 (N_629,N_494,N_276);
or U630 (N_630,N_219,N_18);
nand U631 (N_631,N_275,N_269);
nand U632 (N_632,N_443,N_279);
and U633 (N_633,N_296,N_36);
or U634 (N_634,N_199,N_37);
and U635 (N_635,N_190,N_200);
nand U636 (N_636,N_144,N_595);
xnor U637 (N_637,N_186,N_408);
nand U638 (N_638,N_159,N_593);
xor U639 (N_639,N_548,N_455);
xor U640 (N_640,N_386,N_541);
or U641 (N_641,N_372,N_228);
and U642 (N_642,N_574,N_398);
nor U643 (N_643,N_52,N_585);
and U644 (N_644,N_334,N_415);
xor U645 (N_645,N_515,N_343);
nand U646 (N_646,N_407,N_3);
nand U647 (N_647,N_488,N_430);
and U648 (N_648,N_306,N_232);
and U649 (N_649,N_510,N_51);
nor U650 (N_650,N_198,N_461);
and U651 (N_651,N_17,N_115);
nand U652 (N_652,N_77,N_335);
or U653 (N_653,N_55,N_141);
or U654 (N_654,N_72,N_554);
xor U655 (N_655,N_251,N_272);
and U656 (N_656,N_146,N_182);
nand U657 (N_657,N_454,N_173);
or U658 (N_658,N_290,N_168);
xor U659 (N_659,N_47,N_532);
nor U660 (N_660,N_149,N_352);
xor U661 (N_661,N_555,N_218);
xor U662 (N_662,N_511,N_525);
and U663 (N_663,N_226,N_375);
nand U664 (N_664,N_498,N_259);
xnor U665 (N_665,N_305,N_438);
xor U666 (N_666,N_446,N_458);
or U667 (N_667,N_50,N_414);
nand U668 (N_668,N_124,N_281);
and U669 (N_669,N_462,N_355);
nand U670 (N_670,N_316,N_155);
and U671 (N_671,N_20,N_537);
nor U672 (N_672,N_136,N_210);
nor U673 (N_673,N_167,N_268);
nor U674 (N_674,N_255,N_591);
and U675 (N_675,N_109,N_365);
or U676 (N_676,N_83,N_568);
xnor U677 (N_677,N_431,N_308);
nand U678 (N_678,N_340,N_512);
or U679 (N_679,N_310,N_100);
or U680 (N_680,N_162,N_506);
nor U681 (N_681,N_175,N_399);
nor U682 (N_682,N_564,N_460);
nor U683 (N_683,N_9,N_441);
nor U684 (N_684,N_459,N_318);
and U685 (N_685,N_76,N_261);
nor U686 (N_686,N_363,N_339);
or U687 (N_687,N_206,N_140);
nor U688 (N_688,N_7,N_156);
nor U689 (N_689,N_521,N_153);
xnor U690 (N_690,N_551,N_345);
nor U691 (N_691,N_486,N_93);
and U692 (N_692,N_172,N_91);
and U693 (N_693,N_112,N_196);
or U694 (N_694,N_477,N_361);
nor U695 (N_695,N_371,N_63);
or U696 (N_696,N_464,N_74);
and U697 (N_697,N_347,N_84);
xnor U698 (N_698,N_280,N_553);
nor U699 (N_699,N_292,N_470);
or U700 (N_700,N_505,N_39);
nor U701 (N_701,N_14,N_89);
and U702 (N_702,N_127,N_171);
and U703 (N_703,N_320,N_309);
nand U704 (N_704,N_69,N_263);
nor U705 (N_705,N_192,N_465);
and U706 (N_706,N_475,N_558);
nor U707 (N_707,N_342,N_62);
or U708 (N_708,N_262,N_240);
nor U709 (N_709,N_75,N_557);
nor U710 (N_710,N_125,N_92);
xnor U711 (N_711,N_473,N_170);
nand U712 (N_712,N_594,N_379);
nand U713 (N_713,N_194,N_544);
or U714 (N_714,N_88,N_293);
or U715 (N_715,N_468,N_16);
nand U716 (N_716,N_43,N_2);
nand U717 (N_717,N_289,N_317);
xor U718 (N_718,N_402,N_313);
nand U719 (N_719,N_87,N_221);
nor U720 (N_720,N_71,N_426);
or U721 (N_721,N_56,N_384);
or U722 (N_722,N_97,N_119);
nand U723 (N_723,N_569,N_258);
nand U724 (N_724,N_336,N_562);
or U725 (N_725,N_571,N_507);
xnor U726 (N_726,N_139,N_24);
and U727 (N_727,N_466,N_419);
or U728 (N_728,N_534,N_481);
xor U729 (N_729,N_397,N_231);
nand U730 (N_730,N_270,N_34);
or U731 (N_731,N_392,N_106);
and U732 (N_732,N_535,N_227);
or U733 (N_733,N_110,N_15);
nand U734 (N_734,N_348,N_158);
xor U735 (N_735,N_410,N_191);
or U736 (N_736,N_264,N_400);
xor U737 (N_737,N_54,N_22);
and U738 (N_738,N_599,N_215);
nand U739 (N_739,N_528,N_114);
or U740 (N_740,N_237,N_491);
or U741 (N_741,N_169,N_566);
xor U742 (N_742,N_67,N_394);
xor U743 (N_743,N_185,N_201);
or U744 (N_744,N_444,N_256);
and U745 (N_745,N_418,N_285);
nand U746 (N_746,N_0,N_478);
and U747 (N_747,N_314,N_503);
nand U748 (N_748,N_245,N_366);
and U749 (N_749,N_154,N_500);
and U750 (N_750,N_118,N_423);
nor U751 (N_751,N_300,N_380);
nand U752 (N_752,N_66,N_435);
and U753 (N_753,N_284,N_538);
and U754 (N_754,N_590,N_99);
and U755 (N_755,N_360,N_440);
xnor U756 (N_756,N_563,N_552);
and U757 (N_757,N_273,N_187);
and U758 (N_758,N_572,N_567);
or U759 (N_759,N_483,N_150);
and U760 (N_760,N_518,N_267);
nor U761 (N_761,N_288,N_412);
nor U762 (N_762,N_433,N_331);
or U763 (N_763,N_329,N_376);
or U764 (N_764,N_490,N_103);
or U765 (N_765,N_482,N_195);
or U766 (N_766,N_451,N_223);
xor U767 (N_767,N_70,N_527);
nand U768 (N_768,N_326,N_359);
or U769 (N_769,N_57,N_396);
and U770 (N_770,N_437,N_45);
and U771 (N_771,N_598,N_81);
nor U772 (N_772,N_469,N_225);
nand U773 (N_773,N_246,N_48);
nor U774 (N_774,N_523,N_315);
nand U775 (N_775,N_389,N_416);
and U776 (N_776,N_561,N_592);
nor U777 (N_777,N_94,N_203);
or U778 (N_778,N_28,N_496);
nand U779 (N_779,N_216,N_164);
and U780 (N_780,N_311,N_181);
nand U781 (N_781,N_424,N_577);
nand U782 (N_782,N_220,N_123);
or U783 (N_783,N_447,N_559);
and U784 (N_784,N_539,N_546);
or U785 (N_785,N_236,N_197);
xnor U786 (N_786,N_575,N_579);
or U787 (N_787,N_509,N_13);
or U788 (N_788,N_413,N_550);
or U789 (N_789,N_358,N_492);
nand U790 (N_790,N_420,N_583);
or U791 (N_791,N_565,N_129);
or U792 (N_792,N_1,N_177);
and U793 (N_793,N_282,N_107);
and U794 (N_794,N_202,N_286);
nor U795 (N_795,N_224,N_547);
xnor U796 (N_796,N_243,N_453);
nand U797 (N_797,N_531,N_6);
nor U798 (N_798,N_524,N_530);
xor U799 (N_799,N_341,N_163);
xor U800 (N_800,N_21,N_278);
and U801 (N_801,N_132,N_111);
and U802 (N_802,N_489,N_297);
and U803 (N_803,N_253,N_213);
and U804 (N_804,N_134,N_338);
nand U805 (N_805,N_27,N_307);
or U806 (N_806,N_404,N_549);
or U807 (N_807,N_4,N_117);
nor U808 (N_808,N_248,N_580);
xor U809 (N_809,N_174,N_142);
or U810 (N_810,N_428,N_480);
nand U811 (N_811,N_44,N_8);
nand U812 (N_812,N_312,N_367);
and U813 (N_813,N_337,N_41);
or U814 (N_814,N_301,N_373);
xor U815 (N_815,N_330,N_212);
nand U816 (N_816,N_327,N_122);
and U817 (N_817,N_403,N_233);
and U818 (N_818,N_540,N_46);
nor U819 (N_819,N_325,N_588);
nand U820 (N_820,N_445,N_472);
nand U821 (N_821,N_457,N_229);
or U822 (N_822,N_597,N_133);
and U823 (N_823,N_59,N_434);
or U824 (N_824,N_578,N_369);
and U825 (N_825,N_235,N_61);
or U826 (N_826,N_242,N_157);
nand U827 (N_827,N_105,N_417);
or U828 (N_828,N_128,N_12);
and U829 (N_829,N_176,N_484);
nor U830 (N_830,N_35,N_581);
nand U831 (N_831,N_179,N_249);
nand U832 (N_832,N_135,N_357);
nor U833 (N_833,N_570,N_257);
and U834 (N_834,N_291,N_152);
nor U835 (N_835,N_344,N_436);
nor U836 (N_836,N_96,N_516);
or U837 (N_837,N_529,N_324);
nor U838 (N_838,N_362,N_353);
nand U839 (N_839,N_319,N_302);
and U840 (N_840,N_247,N_274);
nor U841 (N_841,N_350,N_382);
and U842 (N_842,N_26,N_576);
or U843 (N_843,N_456,N_126);
xor U844 (N_844,N_5,N_184);
nor U845 (N_845,N_277,N_165);
and U846 (N_846,N_589,N_421);
or U847 (N_847,N_368,N_587);
or U848 (N_848,N_449,N_113);
or U849 (N_849,N_502,N_499);
nand U850 (N_850,N_328,N_354);
nor U851 (N_851,N_442,N_138);
or U852 (N_852,N_207,N_387);
nor U853 (N_853,N_151,N_98);
nor U854 (N_854,N_432,N_332);
and U855 (N_855,N_239,N_374);
nor U856 (N_856,N_493,N_474);
or U857 (N_857,N_137,N_321);
or U858 (N_858,N_476,N_205);
and U859 (N_859,N_161,N_556);
xnor U860 (N_860,N_364,N_131);
xor U861 (N_861,N_95,N_252);
and U862 (N_862,N_193,N_487);
and U863 (N_863,N_271,N_520);
or U864 (N_864,N_143,N_323);
nand U865 (N_865,N_166,N_545);
nand U866 (N_866,N_102,N_467);
and U867 (N_867,N_333,N_85);
or U868 (N_868,N_378,N_409);
or U869 (N_869,N_211,N_303);
nor U870 (N_870,N_427,N_351);
nor U871 (N_871,N_222,N_370);
nor U872 (N_872,N_33,N_526);
xor U873 (N_873,N_349,N_204);
and U874 (N_874,N_183,N_104);
nand U875 (N_875,N_471,N_582);
nor U876 (N_876,N_584,N_381);
nor U877 (N_877,N_405,N_64);
or U878 (N_878,N_356,N_514);
xor U879 (N_879,N_10,N_522);
and U880 (N_880,N_543,N_542);
xnor U881 (N_881,N_390,N_504);
and U882 (N_882,N_188,N_501);
nand U883 (N_883,N_411,N_573);
nand U884 (N_884,N_254,N_287);
or U885 (N_885,N_68,N_11);
nand U886 (N_886,N_295,N_533);
and U887 (N_887,N_82,N_266);
nand U888 (N_888,N_40,N_406);
nand U889 (N_889,N_147,N_65);
nor U890 (N_890,N_299,N_86);
or U891 (N_891,N_32,N_519);
and U892 (N_892,N_450,N_401);
nor U893 (N_893,N_425,N_283);
and U894 (N_894,N_58,N_29);
nand U895 (N_895,N_78,N_385);
nand U896 (N_896,N_73,N_508);
or U897 (N_897,N_178,N_145);
or U898 (N_898,N_383,N_495);
and U899 (N_899,N_497,N_25);
nor U900 (N_900,N_228,N_400);
or U901 (N_901,N_477,N_290);
or U902 (N_902,N_472,N_284);
xor U903 (N_903,N_285,N_567);
xnor U904 (N_904,N_432,N_112);
nand U905 (N_905,N_359,N_248);
xor U906 (N_906,N_202,N_64);
and U907 (N_907,N_159,N_233);
xnor U908 (N_908,N_341,N_448);
or U909 (N_909,N_91,N_273);
and U910 (N_910,N_397,N_323);
xor U911 (N_911,N_592,N_269);
and U912 (N_912,N_9,N_91);
nor U913 (N_913,N_37,N_252);
and U914 (N_914,N_317,N_515);
nor U915 (N_915,N_405,N_156);
nand U916 (N_916,N_475,N_89);
or U917 (N_917,N_50,N_533);
nor U918 (N_918,N_465,N_449);
and U919 (N_919,N_90,N_386);
nor U920 (N_920,N_181,N_298);
and U921 (N_921,N_148,N_497);
xor U922 (N_922,N_575,N_28);
nand U923 (N_923,N_92,N_526);
and U924 (N_924,N_524,N_289);
nand U925 (N_925,N_427,N_467);
nand U926 (N_926,N_407,N_394);
nor U927 (N_927,N_193,N_269);
nand U928 (N_928,N_433,N_464);
and U929 (N_929,N_424,N_258);
nor U930 (N_930,N_514,N_224);
nor U931 (N_931,N_556,N_433);
and U932 (N_932,N_130,N_69);
and U933 (N_933,N_14,N_2);
and U934 (N_934,N_475,N_150);
nor U935 (N_935,N_519,N_161);
nand U936 (N_936,N_379,N_577);
or U937 (N_937,N_517,N_520);
and U938 (N_938,N_589,N_23);
xnor U939 (N_939,N_398,N_401);
or U940 (N_940,N_544,N_472);
and U941 (N_941,N_120,N_417);
nand U942 (N_942,N_420,N_233);
xor U943 (N_943,N_114,N_370);
nand U944 (N_944,N_198,N_494);
and U945 (N_945,N_429,N_564);
and U946 (N_946,N_392,N_0);
nor U947 (N_947,N_500,N_369);
nor U948 (N_948,N_489,N_408);
nand U949 (N_949,N_51,N_185);
nor U950 (N_950,N_357,N_405);
or U951 (N_951,N_564,N_291);
nand U952 (N_952,N_159,N_460);
and U953 (N_953,N_109,N_56);
and U954 (N_954,N_420,N_228);
xor U955 (N_955,N_464,N_16);
nor U956 (N_956,N_1,N_269);
and U957 (N_957,N_349,N_370);
and U958 (N_958,N_48,N_82);
or U959 (N_959,N_293,N_450);
nand U960 (N_960,N_224,N_341);
or U961 (N_961,N_241,N_415);
and U962 (N_962,N_373,N_147);
nand U963 (N_963,N_592,N_367);
xnor U964 (N_964,N_550,N_299);
or U965 (N_965,N_419,N_58);
nand U966 (N_966,N_76,N_88);
nand U967 (N_967,N_161,N_29);
and U968 (N_968,N_593,N_479);
or U969 (N_969,N_488,N_334);
nor U970 (N_970,N_144,N_590);
nand U971 (N_971,N_426,N_564);
nand U972 (N_972,N_87,N_364);
nand U973 (N_973,N_520,N_119);
xor U974 (N_974,N_449,N_82);
nor U975 (N_975,N_197,N_361);
nor U976 (N_976,N_149,N_505);
or U977 (N_977,N_260,N_245);
and U978 (N_978,N_406,N_424);
nand U979 (N_979,N_203,N_580);
nand U980 (N_980,N_112,N_411);
nand U981 (N_981,N_47,N_120);
nand U982 (N_982,N_451,N_463);
nor U983 (N_983,N_134,N_9);
or U984 (N_984,N_237,N_230);
nor U985 (N_985,N_13,N_382);
or U986 (N_986,N_49,N_338);
or U987 (N_987,N_337,N_16);
nand U988 (N_988,N_3,N_391);
or U989 (N_989,N_430,N_565);
or U990 (N_990,N_192,N_240);
or U991 (N_991,N_389,N_402);
nand U992 (N_992,N_307,N_153);
nand U993 (N_993,N_463,N_296);
and U994 (N_994,N_377,N_120);
or U995 (N_995,N_185,N_84);
and U996 (N_996,N_122,N_13);
and U997 (N_997,N_375,N_497);
nor U998 (N_998,N_266,N_354);
nand U999 (N_999,N_359,N_302);
nand U1000 (N_1000,N_541,N_548);
nor U1001 (N_1001,N_383,N_81);
or U1002 (N_1002,N_294,N_461);
and U1003 (N_1003,N_115,N_485);
nor U1004 (N_1004,N_575,N_229);
and U1005 (N_1005,N_48,N_209);
nand U1006 (N_1006,N_533,N_515);
nand U1007 (N_1007,N_56,N_305);
or U1008 (N_1008,N_455,N_403);
or U1009 (N_1009,N_85,N_15);
and U1010 (N_1010,N_395,N_425);
xnor U1011 (N_1011,N_97,N_210);
nand U1012 (N_1012,N_308,N_172);
nor U1013 (N_1013,N_170,N_587);
and U1014 (N_1014,N_202,N_573);
or U1015 (N_1015,N_546,N_427);
and U1016 (N_1016,N_424,N_529);
and U1017 (N_1017,N_567,N_52);
and U1018 (N_1018,N_156,N_146);
or U1019 (N_1019,N_553,N_365);
and U1020 (N_1020,N_512,N_57);
xnor U1021 (N_1021,N_108,N_125);
nor U1022 (N_1022,N_520,N_0);
and U1023 (N_1023,N_98,N_395);
xor U1024 (N_1024,N_289,N_150);
nand U1025 (N_1025,N_363,N_246);
and U1026 (N_1026,N_184,N_232);
or U1027 (N_1027,N_344,N_188);
or U1028 (N_1028,N_39,N_121);
and U1029 (N_1029,N_336,N_181);
nor U1030 (N_1030,N_115,N_533);
xnor U1031 (N_1031,N_549,N_110);
nor U1032 (N_1032,N_550,N_150);
nor U1033 (N_1033,N_157,N_175);
or U1034 (N_1034,N_403,N_461);
nand U1035 (N_1035,N_599,N_210);
or U1036 (N_1036,N_273,N_232);
nand U1037 (N_1037,N_596,N_82);
or U1038 (N_1038,N_21,N_110);
nand U1039 (N_1039,N_351,N_13);
nor U1040 (N_1040,N_509,N_208);
and U1041 (N_1041,N_380,N_393);
nor U1042 (N_1042,N_451,N_117);
or U1043 (N_1043,N_589,N_407);
nor U1044 (N_1044,N_132,N_552);
and U1045 (N_1045,N_436,N_494);
or U1046 (N_1046,N_376,N_407);
and U1047 (N_1047,N_0,N_591);
or U1048 (N_1048,N_76,N_546);
nor U1049 (N_1049,N_562,N_259);
or U1050 (N_1050,N_222,N_114);
nor U1051 (N_1051,N_566,N_284);
or U1052 (N_1052,N_347,N_579);
or U1053 (N_1053,N_74,N_64);
or U1054 (N_1054,N_257,N_189);
and U1055 (N_1055,N_65,N_159);
nor U1056 (N_1056,N_15,N_494);
nand U1057 (N_1057,N_127,N_434);
nor U1058 (N_1058,N_346,N_587);
and U1059 (N_1059,N_385,N_150);
and U1060 (N_1060,N_19,N_526);
or U1061 (N_1061,N_359,N_458);
nand U1062 (N_1062,N_212,N_413);
nor U1063 (N_1063,N_485,N_129);
or U1064 (N_1064,N_595,N_324);
or U1065 (N_1065,N_236,N_453);
nand U1066 (N_1066,N_58,N_133);
nand U1067 (N_1067,N_258,N_228);
nor U1068 (N_1068,N_477,N_88);
or U1069 (N_1069,N_382,N_52);
or U1070 (N_1070,N_373,N_74);
and U1071 (N_1071,N_5,N_198);
nor U1072 (N_1072,N_101,N_338);
nor U1073 (N_1073,N_237,N_463);
xnor U1074 (N_1074,N_387,N_463);
nand U1075 (N_1075,N_61,N_593);
nor U1076 (N_1076,N_38,N_339);
or U1077 (N_1077,N_594,N_486);
and U1078 (N_1078,N_339,N_109);
nor U1079 (N_1079,N_78,N_20);
nand U1080 (N_1080,N_426,N_428);
or U1081 (N_1081,N_272,N_385);
and U1082 (N_1082,N_128,N_368);
nor U1083 (N_1083,N_63,N_103);
nor U1084 (N_1084,N_341,N_225);
nand U1085 (N_1085,N_228,N_91);
or U1086 (N_1086,N_132,N_498);
nor U1087 (N_1087,N_308,N_513);
xor U1088 (N_1088,N_383,N_394);
xnor U1089 (N_1089,N_566,N_416);
nand U1090 (N_1090,N_327,N_106);
nor U1091 (N_1091,N_331,N_5);
nor U1092 (N_1092,N_105,N_77);
nor U1093 (N_1093,N_306,N_373);
nand U1094 (N_1094,N_422,N_315);
and U1095 (N_1095,N_591,N_557);
nand U1096 (N_1096,N_290,N_63);
and U1097 (N_1097,N_492,N_404);
nand U1098 (N_1098,N_520,N_567);
nand U1099 (N_1099,N_318,N_159);
nand U1100 (N_1100,N_153,N_143);
and U1101 (N_1101,N_544,N_567);
nand U1102 (N_1102,N_288,N_515);
xnor U1103 (N_1103,N_383,N_585);
nor U1104 (N_1104,N_280,N_184);
nor U1105 (N_1105,N_310,N_492);
nand U1106 (N_1106,N_174,N_223);
or U1107 (N_1107,N_110,N_442);
nor U1108 (N_1108,N_593,N_231);
nand U1109 (N_1109,N_27,N_536);
nor U1110 (N_1110,N_347,N_298);
nor U1111 (N_1111,N_459,N_262);
nor U1112 (N_1112,N_515,N_408);
nor U1113 (N_1113,N_485,N_111);
nor U1114 (N_1114,N_455,N_519);
xnor U1115 (N_1115,N_402,N_343);
and U1116 (N_1116,N_550,N_168);
nor U1117 (N_1117,N_141,N_262);
and U1118 (N_1118,N_207,N_518);
nor U1119 (N_1119,N_151,N_35);
nor U1120 (N_1120,N_256,N_403);
or U1121 (N_1121,N_158,N_466);
xor U1122 (N_1122,N_428,N_21);
nand U1123 (N_1123,N_134,N_193);
or U1124 (N_1124,N_538,N_219);
and U1125 (N_1125,N_260,N_430);
or U1126 (N_1126,N_205,N_440);
xor U1127 (N_1127,N_366,N_391);
and U1128 (N_1128,N_43,N_531);
nand U1129 (N_1129,N_119,N_209);
nor U1130 (N_1130,N_169,N_271);
or U1131 (N_1131,N_90,N_599);
nand U1132 (N_1132,N_180,N_63);
nor U1133 (N_1133,N_146,N_437);
nor U1134 (N_1134,N_158,N_596);
nor U1135 (N_1135,N_198,N_363);
and U1136 (N_1136,N_77,N_337);
and U1137 (N_1137,N_412,N_380);
nand U1138 (N_1138,N_305,N_116);
nor U1139 (N_1139,N_334,N_559);
nand U1140 (N_1140,N_133,N_589);
nand U1141 (N_1141,N_526,N_240);
nor U1142 (N_1142,N_7,N_298);
nand U1143 (N_1143,N_470,N_377);
and U1144 (N_1144,N_282,N_581);
nand U1145 (N_1145,N_40,N_145);
nand U1146 (N_1146,N_133,N_182);
and U1147 (N_1147,N_106,N_359);
nor U1148 (N_1148,N_56,N_512);
nor U1149 (N_1149,N_338,N_457);
and U1150 (N_1150,N_7,N_212);
nor U1151 (N_1151,N_362,N_75);
and U1152 (N_1152,N_39,N_472);
nor U1153 (N_1153,N_447,N_97);
or U1154 (N_1154,N_201,N_464);
nand U1155 (N_1155,N_551,N_50);
xnor U1156 (N_1156,N_518,N_52);
nor U1157 (N_1157,N_546,N_60);
nor U1158 (N_1158,N_99,N_92);
and U1159 (N_1159,N_30,N_466);
or U1160 (N_1160,N_82,N_505);
nand U1161 (N_1161,N_388,N_467);
or U1162 (N_1162,N_525,N_440);
nor U1163 (N_1163,N_485,N_390);
or U1164 (N_1164,N_251,N_59);
or U1165 (N_1165,N_4,N_572);
or U1166 (N_1166,N_97,N_395);
or U1167 (N_1167,N_26,N_312);
nand U1168 (N_1168,N_122,N_339);
and U1169 (N_1169,N_353,N_513);
and U1170 (N_1170,N_383,N_519);
nor U1171 (N_1171,N_543,N_579);
or U1172 (N_1172,N_234,N_512);
and U1173 (N_1173,N_134,N_162);
xnor U1174 (N_1174,N_105,N_398);
or U1175 (N_1175,N_539,N_7);
and U1176 (N_1176,N_497,N_106);
and U1177 (N_1177,N_61,N_451);
and U1178 (N_1178,N_5,N_439);
nor U1179 (N_1179,N_266,N_154);
nor U1180 (N_1180,N_359,N_279);
xor U1181 (N_1181,N_490,N_227);
or U1182 (N_1182,N_349,N_117);
and U1183 (N_1183,N_46,N_293);
nand U1184 (N_1184,N_315,N_175);
or U1185 (N_1185,N_259,N_478);
and U1186 (N_1186,N_116,N_569);
and U1187 (N_1187,N_202,N_524);
xnor U1188 (N_1188,N_155,N_363);
and U1189 (N_1189,N_59,N_75);
or U1190 (N_1190,N_473,N_315);
nand U1191 (N_1191,N_460,N_57);
nand U1192 (N_1192,N_312,N_516);
nor U1193 (N_1193,N_482,N_200);
nor U1194 (N_1194,N_41,N_281);
or U1195 (N_1195,N_172,N_335);
or U1196 (N_1196,N_200,N_453);
nand U1197 (N_1197,N_228,N_244);
and U1198 (N_1198,N_177,N_372);
or U1199 (N_1199,N_197,N_384);
xor U1200 (N_1200,N_1018,N_1084);
and U1201 (N_1201,N_894,N_749);
nand U1202 (N_1202,N_1065,N_945);
and U1203 (N_1203,N_831,N_1125);
xnor U1204 (N_1204,N_793,N_991);
nand U1205 (N_1205,N_916,N_1052);
and U1206 (N_1206,N_898,N_988);
or U1207 (N_1207,N_1198,N_690);
nor U1208 (N_1208,N_982,N_997);
nor U1209 (N_1209,N_1031,N_832);
nor U1210 (N_1210,N_817,N_1045);
and U1211 (N_1211,N_860,N_698);
and U1212 (N_1212,N_889,N_910);
nor U1213 (N_1213,N_1121,N_1199);
xor U1214 (N_1214,N_1136,N_1192);
xor U1215 (N_1215,N_932,N_852);
xor U1216 (N_1216,N_963,N_980);
and U1217 (N_1217,N_641,N_699);
nor U1218 (N_1218,N_764,N_752);
nand U1219 (N_1219,N_738,N_1029);
or U1220 (N_1220,N_791,N_790);
nor U1221 (N_1221,N_933,N_1128);
or U1222 (N_1222,N_729,N_723);
xnor U1223 (N_1223,N_1058,N_849);
xor U1224 (N_1224,N_688,N_896);
nand U1225 (N_1225,N_827,N_829);
and U1226 (N_1226,N_1076,N_758);
nand U1227 (N_1227,N_815,N_783);
nand U1228 (N_1228,N_955,N_739);
nand U1229 (N_1229,N_1154,N_1189);
or U1230 (N_1230,N_769,N_984);
xnor U1231 (N_1231,N_661,N_612);
and U1232 (N_1232,N_969,N_838);
nand U1233 (N_1233,N_859,N_744);
xnor U1234 (N_1234,N_1122,N_705);
nand U1235 (N_1235,N_857,N_760);
xnor U1236 (N_1236,N_1069,N_1097);
nor U1237 (N_1237,N_768,N_747);
nor U1238 (N_1238,N_634,N_1176);
and U1239 (N_1239,N_750,N_1126);
and U1240 (N_1240,N_1104,N_950);
and U1241 (N_1241,N_975,N_787);
nor U1242 (N_1242,N_885,N_1183);
nor U1243 (N_1243,N_722,N_998);
nand U1244 (N_1244,N_670,N_850);
nor U1245 (N_1245,N_993,N_1046);
xor U1246 (N_1246,N_702,N_743);
and U1247 (N_1247,N_946,N_856);
nand U1248 (N_1248,N_833,N_708);
and U1249 (N_1249,N_886,N_741);
nand U1250 (N_1250,N_775,N_779);
or U1251 (N_1251,N_620,N_937);
nand U1252 (N_1252,N_754,N_1115);
xnor U1253 (N_1253,N_781,N_610);
or U1254 (N_1254,N_1184,N_732);
or U1255 (N_1255,N_1133,N_1195);
xor U1256 (N_1256,N_1072,N_952);
nand U1257 (N_1257,N_774,N_707);
or U1258 (N_1258,N_989,N_1112);
xor U1259 (N_1259,N_825,N_813);
and U1260 (N_1260,N_746,N_1023);
nor U1261 (N_1261,N_992,N_724);
nor U1262 (N_1262,N_687,N_1147);
and U1263 (N_1263,N_613,N_948);
and U1264 (N_1264,N_865,N_1107);
xor U1265 (N_1265,N_858,N_1061);
and U1266 (N_1266,N_668,N_1186);
xnor U1267 (N_1267,N_1036,N_847);
and U1268 (N_1268,N_1191,N_1078);
nor U1269 (N_1269,N_924,N_1006);
and U1270 (N_1270,N_1012,N_899);
nand U1271 (N_1271,N_805,N_977);
and U1272 (N_1272,N_616,N_1098);
nor U1273 (N_1273,N_1074,N_611);
or U1274 (N_1274,N_1037,N_978);
nor U1275 (N_1275,N_733,N_630);
and U1276 (N_1276,N_962,N_801);
nand U1277 (N_1277,N_936,N_697);
or U1278 (N_1278,N_715,N_1020);
nand U1279 (N_1279,N_1068,N_742);
or U1280 (N_1280,N_1030,N_861);
and U1281 (N_1281,N_1173,N_897);
and U1282 (N_1282,N_682,N_1120);
xor U1283 (N_1283,N_822,N_1049);
nand U1284 (N_1284,N_1146,N_1178);
nor U1285 (N_1285,N_872,N_1063);
and U1286 (N_1286,N_944,N_663);
and U1287 (N_1287,N_1181,N_807);
nand U1288 (N_1288,N_622,N_1132);
or U1289 (N_1289,N_920,N_1040);
xor U1290 (N_1290,N_785,N_953);
and U1291 (N_1291,N_1075,N_915);
nand U1292 (N_1292,N_922,N_776);
and U1293 (N_1293,N_1157,N_911);
nand U1294 (N_1294,N_632,N_864);
nor U1295 (N_1295,N_1057,N_1160);
or U1296 (N_1296,N_1190,N_1105);
or U1297 (N_1297,N_882,N_1130);
xnor U1298 (N_1298,N_674,N_653);
nand U1299 (N_1299,N_1100,N_660);
and U1300 (N_1300,N_1059,N_931);
nand U1301 (N_1301,N_693,N_655);
nor U1302 (N_1302,N_820,N_794);
nor U1303 (N_1303,N_638,N_711);
or U1304 (N_1304,N_996,N_649);
xnor U1305 (N_1305,N_782,N_740);
nor U1306 (N_1306,N_873,N_999);
nand U1307 (N_1307,N_645,N_1153);
nor U1308 (N_1308,N_1127,N_1197);
xnor U1309 (N_1309,N_1110,N_985);
and U1310 (N_1310,N_965,N_600);
nor U1311 (N_1311,N_748,N_907);
or U1312 (N_1312,N_1109,N_1138);
nor U1313 (N_1313,N_935,N_766);
and U1314 (N_1314,N_934,N_617);
and U1315 (N_1315,N_1182,N_680);
and U1316 (N_1316,N_1027,N_631);
nand U1317 (N_1317,N_761,N_713);
and U1318 (N_1318,N_929,N_995);
nor U1319 (N_1319,N_1116,N_796);
and U1320 (N_1320,N_1088,N_1161);
and U1321 (N_1321,N_854,N_951);
or U1322 (N_1322,N_1156,N_1113);
nand U1323 (N_1323,N_710,N_725);
nand U1324 (N_1324,N_973,N_1167);
and U1325 (N_1325,N_1007,N_1079);
or U1326 (N_1326,N_1005,N_1196);
nand U1327 (N_1327,N_971,N_1095);
nand U1328 (N_1328,N_737,N_1148);
and U1329 (N_1329,N_1062,N_1001);
xor U1330 (N_1330,N_1013,N_1086);
and U1331 (N_1331,N_607,N_673);
or U1332 (N_1332,N_770,N_976);
xor U1333 (N_1333,N_1188,N_1170);
nand U1334 (N_1334,N_651,N_1048);
nor U1335 (N_1335,N_666,N_851);
or U1336 (N_1336,N_703,N_875);
nor U1337 (N_1337,N_689,N_621);
nand U1338 (N_1338,N_877,N_974);
nor U1339 (N_1339,N_731,N_837);
nand U1340 (N_1340,N_1083,N_902);
xnor U1341 (N_1341,N_614,N_1093);
or U1342 (N_1342,N_784,N_671);
nand U1343 (N_1343,N_892,N_956);
or U1344 (N_1344,N_1165,N_844);
and U1345 (N_1345,N_1087,N_986);
xor U1346 (N_1346,N_718,N_804);
nand U1347 (N_1347,N_925,N_667);
and U1348 (N_1348,N_1101,N_840);
and U1349 (N_1349,N_765,N_1047);
nand U1350 (N_1350,N_601,N_1108);
xnor U1351 (N_1351,N_762,N_843);
nor U1352 (N_1352,N_818,N_845);
or U1353 (N_1353,N_990,N_695);
xor U1354 (N_1354,N_1016,N_1021);
xor U1355 (N_1355,N_968,N_958);
nor U1356 (N_1356,N_949,N_836);
nand U1357 (N_1357,N_1073,N_706);
nor U1358 (N_1358,N_947,N_1011);
nand U1359 (N_1359,N_1017,N_1090);
or U1360 (N_1360,N_828,N_623);
or U1361 (N_1361,N_772,N_1015);
nor U1362 (N_1362,N_879,N_657);
and U1363 (N_1363,N_830,N_893);
nor U1364 (N_1364,N_692,N_773);
xnor U1365 (N_1365,N_625,N_789);
nor U1366 (N_1366,N_1131,N_903);
or U1367 (N_1367,N_1053,N_756);
and U1368 (N_1368,N_786,N_867);
or U1369 (N_1369,N_928,N_1129);
and U1370 (N_1370,N_778,N_643);
nand U1371 (N_1371,N_834,N_1151);
and U1372 (N_1372,N_1039,N_826);
or U1373 (N_1373,N_771,N_628);
xnor U1374 (N_1374,N_798,N_1174);
or U1375 (N_1375,N_868,N_918);
nor U1376 (N_1376,N_615,N_1091);
and U1377 (N_1377,N_800,N_1043);
and U1378 (N_1378,N_1168,N_639);
and U1379 (N_1379,N_887,N_1042);
and U1380 (N_1380,N_1092,N_862);
nor U1381 (N_1381,N_642,N_1149);
nor U1382 (N_1382,N_1159,N_901);
nand U1383 (N_1383,N_1171,N_717);
or U1384 (N_1384,N_1099,N_913);
xnor U1385 (N_1385,N_1187,N_1067);
xnor U1386 (N_1386,N_633,N_923);
nand U1387 (N_1387,N_987,N_972);
nor U1388 (N_1388,N_635,N_1003);
and U1389 (N_1389,N_1004,N_1185);
nand U1390 (N_1390,N_626,N_881);
nand U1391 (N_1391,N_679,N_909);
nand U1392 (N_1392,N_966,N_1009);
nor U1393 (N_1393,N_957,N_1102);
nand U1394 (N_1394,N_629,N_880);
and U1395 (N_1395,N_811,N_1034);
or U1396 (N_1396,N_1055,N_757);
nor U1397 (N_1397,N_812,N_681);
nand U1398 (N_1398,N_810,N_1145);
nand U1399 (N_1399,N_954,N_914);
nor U1400 (N_1400,N_1119,N_883);
or U1401 (N_1401,N_1158,N_1014);
and U1402 (N_1402,N_700,N_665);
and U1403 (N_1403,N_1169,N_1117);
or U1404 (N_1404,N_619,N_1162);
nor U1405 (N_1405,N_1135,N_792);
nand U1406 (N_1406,N_846,N_927);
or U1407 (N_1407,N_1150,N_606);
and U1408 (N_1408,N_664,N_994);
xor U1409 (N_1409,N_677,N_876);
or U1410 (N_1410,N_719,N_751);
xor U1411 (N_1411,N_735,N_1096);
or U1412 (N_1412,N_1044,N_1033);
nor U1413 (N_1413,N_1028,N_1032);
nor U1414 (N_1414,N_795,N_1035);
and U1415 (N_1415,N_696,N_675);
nor U1416 (N_1416,N_1123,N_835);
nand U1417 (N_1417,N_912,N_608);
and U1418 (N_1418,N_1139,N_809);
nand U1419 (N_1419,N_961,N_839);
nor U1420 (N_1420,N_841,N_1179);
or U1421 (N_1421,N_604,N_802);
and U1422 (N_1422,N_1144,N_658);
or U1423 (N_1423,N_848,N_1025);
xor U1424 (N_1424,N_1141,N_648);
and U1425 (N_1425,N_1124,N_1111);
nor U1426 (N_1426,N_759,N_1118);
nor U1427 (N_1427,N_656,N_669);
and U1428 (N_1428,N_605,N_1163);
nor U1429 (N_1429,N_926,N_1175);
nor U1430 (N_1430,N_808,N_672);
nor U1431 (N_1431,N_942,N_797);
xor U1432 (N_1432,N_728,N_1140);
or U1433 (N_1433,N_959,N_1051);
and U1434 (N_1434,N_755,N_763);
and U1435 (N_1435,N_1082,N_647);
nand U1436 (N_1436,N_1041,N_970);
nand U1437 (N_1437,N_853,N_870);
or U1438 (N_1438,N_1180,N_943);
nand U1439 (N_1439,N_1089,N_1114);
nand U1440 (N_1440,N_866,N_727);
nand U1441 (N_1441,N_676,N_1094);
or U1442 (N_1442,N_803,N_983);
or U1443 (N_1443,N_981,N_1106);
nand U1444 (N_1444,N_694,N_684);
nor U1445 (N_1445,N_788,N_799);
and U1446 (N_1446,N_891,N_1054);
and U1447 (N_1447,N_964,N_1164);
nor U1448 (N_1448,N_709,N_816);
or U1449 (N_1449,N_721,N_678);
or U1450 (N_1450,N_1155,N_753);
and U1451 (N_1451,N_967,N_1050);
nor U1452 (N_1452,N_979,N_842);
nand U1453 (N_1453,N_1019,N_1081);
nor U1454 (N_1454,N_819,N_921);
nor U1455 (N_1455,N_1066,N_736);
or U1456 (N_1456,N_1194,N_659);
nand U1457 (N_1457,N_917,N_691);
nand U1458 (N_1458,N_908,N_603);
or U1459 (N_1459,N_895,N_888);
or U1460 (N_1460,N_1166,N_730);
nor U1461 (N_1461,N_941,N_939);
nand U1462 (N_1462,N_602,N_1137);
nand U1463 (N_1463,N_652,N_701);
nor U1464 (N_1464,N_1002,N_646);
nand U1465 (N_1465,N_1077,N_1024);
nor U1466 (N_1466,N_1071,N_720);
and U1467 (N_1467,N_686,N_636);
nand U1468 (N_1468,N_662,N_704);
and U1469 (N_1469,N_1172,N_734);
and U1470 (N_1470,N_906,N_890);
and U1471 (N_1471,N_1000,N_1038);
or U1472 (N_1472,N_930,N_884);
nand U1473 (N_1473,N_714,N_869);
or U1474 (N_1474,N_627,N_874);
or U1475 (N_1475,N_609,N_823);
nor U1476 (N_1476,N_767,N_640);
and U1477 (N_1477,N_814,N_900);
and U1478 (N_1478,N_1177,N_1080);
or U1479 (N_1479,N_1143,N_855);
or U1480 (N_1480,N_919,N_904);
or U1481 (N_1481,N_871,N_683);
or U1482 (N_1482,N_960,N_1056);
xor U1483 (N_1483,N_1134,N_1026);
or U1484 (N_1484,N_1060,N_940);
nand U1485 (N_1485,N_1064,N_1142);
and U1486 (N_1486,N_644,N_716);
nand U1487 (N_1487,N_685,N_863);
or U1488 (N_1488,N_1193,N_821);
and U1489 (N_1489,N_654,N_780);
and U1490 (N_1490,N_1008,N_878);
nand U1491 (N_1491,N_618,N_650);
nor U1492 (N_1492,N_1152,N_1103);
nor U1493 (N_1493,N_637,N_1022);
and U1494 (N_1494,N_824,N_905);
and U1495 (N_1495,N_1010,N_806);
xnor U1496 (N_1496,N_938,N_1085);
xnor U1497 (N_1497,N_1070,N_712);
nor U1498 (N_1498,N_777,N_624);
or U1499 (N_1499,N_726,N_745);
nor U1500 (N_1500,N_1134,N_1035);
or U1501 (N_1501,N_831,N_788);
nor U1502 (N_1502,N_700,N_1027);
and U1503 (N_1503,N_1143,N_644);
nor U1504 (N_1504,N_839,N_702);
xor U1505 (N_1505,N_916,N_1149);
and U1506 (N_1506,N_934,N_686);
and U1507 (N_1507,N_839,N_844);
and U1508 (N_1508,N_700,N_1141);
xnor U1509 (N_1509,N_1152,N_869);
xor U1510 (N_1510,N_915,N_824);
nand U1511 (N_1511,N_762,N_654);
nand U1512 (N_1512,N_786,N_1027);
or U1513 (N_1513,N_1095,N_641);
or U1514 (N_1514,N_667,N_944);
nand U1515 (N_1515,N_1195,N_712);
nor U1516 (N_1516,N_956,N_1119);
xnor U1517 (N_1517,N_724,N_932);
and U1518 (N_1518,N_1057,N_1049);
and U1519 (N_1519,N_760,N_879);
and U1520 (N_1520,N_1021,N_685);
and U1521 (N_1521,N_885,N_1120);
and U1522 (N_1522,N_779,N_1108);
or U1523 (N_1523,N_926,N_1069);
nand U1524 (N_1524,N_794,N_600);
nor U1525 (N_1525,N_785,N_1029);
nand U1526 (N_1526,N_1028,N_838);
nor U1527 (N_1527,N_866,N_926);
nand U1528 (N_1528,N_790,N_1012);
and U1529 (N_1529,N_1076,N_1182);
or U1530 (N_1530,N_931,N_978);
nor U1531 (N_1531,N_1020,N_1014);
nand U1532 (N_1532,N_1171,N_1030);
or U1533 (N_1533,N_691,N_1133);
or U1534 (N_1534,N_1123,N_600);
and U1535 (N_1535,N_1198,N_1140);
nor U1536 (N_1536,N_942,N_605);
and U1537 (N_1537,N_1194,N_978);
or U1538 (N_1538,N_1005,N_974);
and U1539 (N_1539,N_659,N_832);
xnor U1540 (N_1540,N_807,N_801);
or U1541 (N_1541,N_955,N_1163);
and U1542 (N_1542,N_695,N_776);
nand U1543 (N_1543,N_1059,N_810);
nand U1544 (N_1544,N_929,N_676);
xor U1545 (N_1545,N_1168,N_685);
nand U1546 (N_1546,N_880,N_755);
nand U1547 (N_1547,N_820,N_1004);
or U1548 (N_1548,N_782,N_905);
nor U1549 (N_1549,N_738,N_1090);
xnor U1550 (N_1550,N_899,N_884);
nand U1551 (N_1551,N_1096,N_1050);
nor U1552 (N_1552,N_1076,N_632);
and U1553 (N_1553,N_937,N_1148);
nor U1554 (N_1554,N_989,N_896);
or U1555 (N_1555,N_952,N_897);
or U1556 (N_1556,N_957,N_956);
or U1557 (N_1557,N_844,N_1158);
and U1558 (N_1558,N_808,N_871);
nor U1559 (N_1559,N_882,N_1029);
xor U1560 (N_1560,N_1120,N_1036);
and U1561 (N_1561,N_640,N_717);
nor U1562 (N_1562,N_857,N_770);
and U1563 (N_1563,N_865,N_626);
or U1564 (N_1564,N_1115,N_1168);
or U1565 (N_1565,N_1010,N_974);
and U1566 (N_1566,N_933,N_707);
or U1567 (N_1567,N_1026,N_677);
and U1568 (N_1568,N_872,N_721);
and U1569 (N_1569,N_1116,N_1073);
nor U1570 (N_1570,N_770,N_774);
xnor U1571 (N_1571,N_742,N_952);
nand U1572 (N_1572,N_750,N_888);
or U1573 (N_1573,N_804,N_956);
nand U1574 (N_1574,N_860,N_716);
nand U1575 (N_1575,N_774,N_1154);
or U1576 (N_1576,N_1089,N_694);
or U1577 (N_1577,N_700,N_783);
nand U1578 (N_1578,N_953,N_609);
nand U1579 (N_1579,N_733,N_1068);
and U1580 (N_1580,N_721,N_1040);
nor U1581 (N_1581,N_1027,N_1061);
or U1582 (N_1582,N_991,N_898);
nor U1583 (N_1583,N_996,N_774);
nand U1584 (N_1584,N_974,N_1099);
nor U1585 (N_1585,N_944,N_624);
and U1586 (N_1586,N_1021,N_952);
nor U1587 (N_1587,N_810,N_769);
or U1588 (N_1588,N_903,N_1168);
and U1589 (N_1589,N_1088,N_1078);
nor U1590 (N_1590,N_936,N_915);
nand U1591 (N_1591,N_803,N_775);
and U1592 (N_1592,N_905,N_751);
nand U1593 (N_1593,N_1110,N_1061);
and U1594 (N_1594,N_828,N_662);
nor U1595 (N_1595,N_905,N_904);
nor U1596 (N_1596,N_619,N_1017);
and U1597 (N_1597,N_872,N_791);
xnor U1598 (N_1598,N_971,N_901);
and U1599 (N_1599,N_802,N_1049);
or U1600 (N_1600,N_676,N_1168);
nor U1601 (N_1601,N_991,N_981);
and U1602 (N_1602,N_1076,N_905);
or U1603 (N_1603,N_1011,N_841);
nor U1604 (N_1604,N_980,N_905);
nor U1605 (N_1605,N_810,N_648);
nor U1606 (N_1606,N_1191,N_622);
nor U1607 (N_1607,N_653,N_1185);
or U1608 (N_1608,N_783,N_948);
or U1609 (N_1609,N_1129,N_831);
xor U1610 (N_1610,N_1103,N_803);
nand U1611 (N_1611,N_800,N_799);
or U1612 (N_1612,N_661,N_760);
and U1613 (N_1613,N_1168,N_825);
or U1614 (N_1614,N_640,N_1036);
or U1615 (N_1615,N_1141,N_946);
and U1616 (N_1616,N_1107,N_1136);
and U1617 (N_1617,N_1165,N_1027);
nand U1618 (N_1618,N_1003,N_1049);
nand U1619 (N_1619,N_976,N_1042);
nand U1620 (N_1620,N_1019,N_604);
or U1621 (N_1621,N_617,N_1035);
xor U1622 (N_1622,N_818,N_998);
nor U1623 (N_1623,N_1072,N_732);
nand U1624 (N_1624,N_818,N_779);
and U1625 (N_1625,N_817,N_613);
and U1626 (N_1626,N_769,N_999);
nor U1627 (N_1627,N_609,N_1041);
or U1628 (N_1628,N_1154,N_1085);
nand U1629 (N_1629,N_1021,N_702);
nand U1630 (N_1630,N_619,N_1189);
nor U1631 (N_1631,N_1018,N_1101);
or U1632 (N_1632,N_652,N_733);
nand U1633 (N_1633,N_629,N_1143);
or U1634 (N_1634,N_675,N_1186);
and U1635 (N_1635,N_962,N_964);
or U1636 (N_1636,N_775,N_1157);
nand U1637 (N_1637,N_1051,N_1071);
or U1638 (N_1638,N_1111,N_725);
nand U1639 (N_1639,N_936,N_1005);
xnor U1640 (N_1640,N_650,N_922);
nand U1641 (N_1641,N_899,N_1048);
nand U1642 (N_1642,N_1036,N_902);
nor U1643 (N_1643,N_1134,N_604);
nor U1644 (N_1644,N_938,N_1145);
or U1645 (N_1645,N_1109,N_716);
nor U1646 (N_1646,N_1180,N_1103);
and U1647 (N_1647,N_1044,N_881);
nor U1648 (N_1648,N_1099,N_689);
or U1649 (N_1649,N_1059,N_1035);
and U1650 (N_1650,N_693,N_1065);
and U1651 (N_1651,N_812,N_1106);
nand U1652 (N_1652,N_1132,N_644);
and U1653 (N_1653,N_1081,N_1013);
or U1654 (N_1654,N_1048,N_1015);
and U1655 (N_1655,N_1163,N_633);
and U1656 (N_1656,N_773,N_907);
nor U1657 (N_1657,N_747,N_895);
nor U1658 (N_1658,N_1167,N_1005);
or U1659 (N_1659,N_949,N_840);
and U1660 (N_1660,N_647,N_1116);
nor U1661 (N_1661,N_1056,N_973);
nand U1662 (N_1662,N_1033,N_1192);
nor U1663 (N_1663,N_1034,N_657);
or U1664 (N_1664,N_865,N_1157);
or U1665 (N_1665,N_796,N_618);
and U1666 (N_1666,N_800,N_1098);
or U1667 (N_1667,N_777,N_913);
nor U1668 (N_1668,N_1098,N_610);
and U1669 (N_1669,N_705,N_632);
nand U1670 (N_1670,N_1115,N_651);
nand U1671 (N_1671,N_1180,N_967);
nand U1672 (N_1672,N_879,N_653);
xor U1673 (N_1673,N_761,N_1082);
or U1674 (N_1674,N_767,N_989);
nand U1675 (N_1675,N_966,N_792);
nor U1676 (N_1676,N_1177,N_1109);
and U1677 (N_1677,N_1063,N_1175);
or U1678 (N_1678,N_677,N_1176);
nand U1679 (N_1679,N_645,N_861);
and U1680 (N_1680,N_824,N_937);
or U1681 (N_1681,N_665,N_1124);
or U1682 (N_1682,N_1038,N_630);
and U1683 (N_1683,N_883,N_1164);
and U1684 (N_1684,N_968,N_925);
nand U1685 (N_1685,N_919,N_998);
and U1686 (N_1686,N_875,N_960);
or U1687 (N_1687,N_838,N_710);
nand U1688 (N_1688,N_1089,N_928);
or U1689 (N_1689,N_1128,N_913);
or U1690 (N_1690,N_736,N_613);
xor U1691 (N_1691,N_674,N_706);
and U1692 (N_1692,N_625,N_989);
nor U1693 (N_1693,N_1052,N_1053);
and U1694 (N_1694,N_1048,N_1044);
nor U1695 (N_1695,N_1145,N_1072);
nand U1696 (N_1696,N_652,N_770);
xor U1697 (N_1697,N_1108,N_647);
nand U1698 (N_1698,N_1102,N_1111);
or U1699 (N_1699,N_993,N_1139);
and U1700 (N_1700,N_1154,N_786);
or U1701 (N_1701,N_1004,N_1027);
nor U1702 (N_1702,N_903,N_1192);
or U1703 (N_1703,N_1039,N_819);
or U1704 (N_1704,N_821,N_991);
nor U1705 (N_1705,N_652,N_1180);
and U1706 (N_1706,N_857,N_759);
nor U1707 (N_1707,N_1168,N_830);
and U1708 (N_1708,N_686,N_1107);
and U1709 (N_1709,N_669,N_1015);
nor U1710 (N_1710,N_910,N_1122);
and U1711 (N_1711,N_637,N_770);
nor U1712 (N_1712,N_997,N_941);
nand U1713 (N_1713,N_935,N_645);
nor U1714 (N_1714,N_1163,N_895);
or U1715 (N_1715,N_1000,N_695);
xnor U1716 (N_1716,N_804,N_1087);
nand U1717 (N_1717,N_657,N_931);
or U1718 (N_1718,N_1034,N_637);
or U1719 (N_1719,N_868,N_783);
and U1720 (N_1720,N_724,N_755);
nand U1721 (N_1721,N_1023,N_753);
and U1722 (N_1722,N_859,N_946);
and U1723 (N_1723,N_783,N_967);
nand U1724 (N_1724,N_1018,N_1071);
nor U1725 (N_1725,N_914,N_1176);
or U1726 (N_1726,N_860,N_858);
and U1727 (N_1727,N_875,N_1150);
or U1728 (N_1728,N_1063,N_1197);
xor U1729 (N_1729,N_969,N_1072);
xnor U1730 (N_1730,N_1111,N_1018);
nor U1731 (N_1731,N_1106,N_957);
nor U1732 (N_1732,N_659,N_823);
nor U1733 (N_1733,N_894,N_692);
or U1734 (N_1734,N_1185,N_768);
nand U1735 (N_1735,N_1045,N_1082);
xor U1736 (N_1736,N_1135,N_1063);
or U1737 (N_1737,N_955,N_887);
nor U1738 (N_1738,N_919,N_993);
xnor U1739 (N_1739,N_795,N_987);
and U1740 (N_1740,N_674,N_1084);
nand U1741 (N_1741,N_1181,N_687);
xnor U1742 (N_1742,N_1159,N_1136);
nand U1743 (N_1743,N_1121,N_879);
or U1744 (N_1744,N_1034,N_757);
or U1745 (N_1745,N_1099,N_807);
nand U1746 (N_1746,N_1043,N_1000);
or U1747 (N_1747,N_877,N_1069);
xnor U1748 (N_1748,N_742,N_898);
or U1749 (N_1749,N_905,N_696);
and U1750 (N_1750,N_789,N_835);
xor U1751 (N_1751,N_901,N_655);
or U1752 (N_1752,N_774,N_1061);
or U1753 (N_1753,N_909,N_714);
or U1754 (N_1754,N_840,N_847);
nand U1755 (N_1755,N_1127,N_935);
nand U1756 (N_1756,N_1007,N_1053);
or U1757 (N_1757,N_1166,N_790);
or U1758 (N_1758,N_733,N_743);
or U1759 (N_1759,N_677,N_926);
and U1760 (N_1760,N_1129,N_776);
nand U1761 (N_1761,N_847,N_625);
nand U1762 (N_1762,N_1190,N_885);
or U1763 (N_1763,N_1141,N_738);
nor U1764 (N_1764,N_655,N_686);
nor U1765 (N_1765,N_1069,N_914);
and U1766 (N_1766,N_917,N_1168);
nand U1767 (N_1767,N_1196,N_1188);
or U1768 (N_1768,N_765,N_817);
and U1769 (N_1769,N_827,N_1019);
nand U1770 (N_1770,N_1066,N_1025);
nor U1771 (N_1771,N_808,N_948);
and U1772 (N_1772,N_880,N_796);
and U1773 (N_1773,N_834,N_708);
or U1774 (N_1774,N_1105,N_831);
nand U1775 (N_1775,N_725,N_1027);
and U1776 (N_1776,N_661,N_854);
nor U1777 (N_1777,N_1182,N_682);
nand U1778 (N_1778,N_1181,N_871);
nor U1779 (N_1779,N_825,N_697);
nor U1780 (N_1780,N_1013,N_857);
or U1781 (N_1781,N_1057,N_1110);
nand U1782 (N_1782,N_1008,N_987);
and U1783 (N_1783,N_753,N_914);
and U1784 (N_1784,N_713,N_1062);
and U1785 (N_1785,N_1008,N_616);
or U1786 (N_1786,N_821,N_1199);
or U1787 (N_1787,N_1056,N_826);
nand U1788 (N_1788,N_1059,N_1039);
xor U1789 (N_1789,N_1004,N_903);
nor U1790 (N_1790,N_874,N_728);
or U1791 (N_1791,N_626,N_986);
nor U1792 (N_1792,N_871,N_1102);
nor U1793 (N_1793,N_796,N_1141);
nor U1794 (N_1794,N_1069,N_792);
or U1795 (N_1795,N_642,N_655);
nand U1796 (N_1796,N_638,N_890);
nand U1797 (N_1797,N_658,N_790);
and U1798 (N_1798,N_950,N_974);
xor U1799 (N_1799,N_994,N_894);
nand U1800 (N_1800,N_1416,N_1579);
nand U1801 (N_1801,N_1701,N_1481);
nor U1802 (N_1802,N_1461,N_1388);
nand U1803 (N_1803,N_1747,N_1488);
or U1804 (N_1804,N_1665,N_1402);
nand U1805 (N_1805,N_1492,N_1243);
or U1806 (N_1806,N_1508,N_1353);
and U1807 (N_1807,N_1202,N_1656);
nand U1808 (N_1808,N_1465,N_1386);
and U1809 (N_1809,N_1772,N_1250);
or U1810 (N_1810,N_1329,N_1726);
nand U1811 (N_1811,N_1457,N_1498);
nor U1812 (N_1812,N_1359,N_1373);
or U1813 (N_1813,N_1580,N_1374);
nor U1814 (N_1814,N_1491,N_1438);
or U1815 (N_1815,N_1682,N_1423);
or U1816 (N_1816,N_1332,N_1755);
and U1817 (N_1817,N_1742,N_1697);
nand U1818 (N_1818,N_1437,N_1774);
or U1819 (N_1819,N_1568,N_1396);
nor U1820 (N_1820,N_1661,N_1522);
nor U1821 (N_1821,N_1559,N_1392);
nor U1822 (N_1822,N_1277,N_1748);
and U1823 (N_1823,N_1723,N_1504);
or U1824 (N_1824,N_1229,N_1347);
or U1825 (N_1825,N_1305,N_1535);
nand U1826 (N_1826,N_1647,N_1418);
nor U1827 (N_1827,N_1274,N_1414);
or U1828 (N_1828,N_1589,N_1267);
or U1829 (N_1829,N_1218,N_1345);
or U1830 (N_1830,N_1462,N_1489);
nand U1831 (N_1831,N_1484,N_1474);
and U1832 (N_1832,N_1537,N_1595);
nand U1833 (N_1833,N_1781,N_1735);
and U1834 (N_1834,N_1483,N_1797);
nand U1835 (N_1835,N_1292,N_1238);
and U1836 (N_1836,N_1715,N_1677);
and U1837 (N_1837,N_1658,N_1672);
nand U1838 (N_1838,N_1684,N_1699);
or U1839 (N_1839,N_1338,N_1683);
or U1840 (N_1840,N_1257,N_1317);
and U1841 (N_1841,N_1246,N_1389);
and U1842 (N_1842,N_1371,N_1639);
or U1843 (N_1843,N_1564,N_1517);
nand U1844 (N_1844,N_1585,N_1694);
or U1845 (N_1845,N_1569,N_1527);
nand U1846 (N_1846,N_1577,N_1296);
nand U1847 (N_1847,N_1335,N_1599);
nand U1848 (N_1848,N_1663,N_1224);
nor U1849 (N_1849,N_1350,N_1773);
or U1850 (N_1850,N_1372,N_1744);
nor U1851 (N_1851,N_1566,N_1621);
and U1852 (N_1852,N_1383,N_1709);
nor U1853 (N_1853,N_1429,N_1385);
and U1854 (N_1854,N_1295,N_1512);
or U1855 (N_1855,N_1354,N_1226);
or U1856 (N_1856,N_1320,N_1617);
nand U1857 (N_1857,N_1265,N_1752);
or U1858 (N_1858,N_1601,N_1549);
nand U1859 (N_1859,N_1649,N_1505);
nand U1860 (N_1860,N_1273,N_1209);
nor U1861 (N_1861,N_1328,N_1557);
nor U1862 (N_1862,N_1690,N_1646);
nor U1863 (N_1863,N_1349,N_1252);
or U1864 (N_1864,N_1738,N_1315);
xnor U1865 (N_1865,N_1234,N_1679);
xnor U1866 (N_1866,N_1608,N_1379);
and U1867 (N_1867,N_1361,N_1464);
nand U1868 (N_1868,N_1369,N_1458);
and U1869 (N_1869,N_1763,N_1378);
nor U1870 (N_1870,N_1611,N_1327);
nor U1871 (N_1871,N_1436,N_1572);
nor U1872 (N_1872,N_1479,N_1664);
and U1873 (N_1873,N_1741,N_1757);
nor U1874 (N_1874,N_1563,N_1771);
nor U1875 (N_1875,N_1231,N_1603);
nand U1876 (N_1876,N_1553,N_1310);
nor U1877 (N_1877,N_1318,N_1214);
nor U1878 (N_1878,N_1653,N_1201);
or U1879 (N_1879,N_1263,N_1681);
or U1880 (N_1880,N_1754,N_1625);
xnor U1881 (N_1881,N_1629,N_1669);
xnor U1882 (N_1882,N_1521,N_1552);
nand U1883 (N_1883,N_1666,N_1312);
nor U1884 (N_1884,N_1544,N_1536);
or U1885 (N_1885,N_1671,N_1627);
nor U1886 (N_1886,N_1290,N_1217);
nand U1887 (N_1887,N_1759,N_1430);
and U1888 (N_1888,N_1788,N_1779);
or U1889 (N_1889,N_1390,N_1518);
nor U1890 (N_1890,N_1657,N_1415);
nor U1891 (N_1891,N_1790,N_1322);
and U1892 (N_1892,N_1721,N_1469);
or U1893 (N_1893,N_1323,N_1737);
nand U1894 (N_1894,N_1734,N_1333);
xnor U1895 (N_1895,N_1395,N_1794);
nand U1896 (N_1896,N_1542,N_1729);
and U1897 (N_1897,N_1643,N_1478);
or U1898 (N_1898,N_1344,N_1631);
or U1899 (N_1899,N_1235,N_1460);
nor U1900 (N_1900,N_1583,N_1507);
nor U1901 (N_1901,N_1541,N_1365);
nand U1902 (N_1902,N_1356,N_1545);
nand U1903 (N_1903,N_1792,N_1602);
nand U1904 (N_1904,N_1565,N_1405);
and U1905 (N_1905,N_1482,N_1686);
nand U1906 (N_1906,N_1495,N_1760);
nand U1907 (N_1907,N_1337,N_1219);
or U1908 (N_1908,N_1467,N_1576);
xnor U1909 (N_1909,N_1311,N_1753);
nor U1910 (N_1910,N_1449,N_1300);
or U1911 (N_1911,N_1309,N_1404);
or U1912 (N_1912,N_1427,N_1421);
or U1913 (N_1913,N_1206,N_1299);
nor U1914 (N_1914,N_1503,N_1302);
and U1915 (N_1915,N_1346,N_1357);
or U1916 (N_1916,N_1640,N_1275);
nor U1917 (N_1917,N_1515,N_1348);
nand U1918 (N_1918,N_1710,N_1410);
or U1919 (N_1919,N_1204,N_1780);
and U1920 (N_1920,N_1783,N_1223);
nand U1921 (N_1921,N_1285,N_1447);
and U1922 (N_1922,N_1700,N_1584);
and U1923 (N_1923,N_1225,N_1650);
or U1924 (N_1924,N_1466,N_1502);
xnor U1925 (N_1925,N_1705,N_1413);
nand U1926 (N_1926,N_1698,N_1367);
nand U1927 (N_1927,N_1330,N_1590);
nand U1928 (N_1928,N_1638,N_1662);
nor U1929 (N_1929,N_1432,N_1674);
and U1930 (N_1930,N_1500,N_1615);
or U1931 (N_1931,N_1393,N_1475);
nand U1932 (N_1932,N_1454,N_1546);
and U1933 (N_1933,N_1716,N_1221);
or U1934 (N_1934,N_1336,N_1255);
nor U1935 (N_1935,N_1745,N_1220);
or U1936 (N_1936,N_1613,N_1200);
nand U1937 (N_1937,N_1695,N_1736);
nor U1938 (N_1938,N_1406,N_1494);
nand U1939 (N_1939,N_1499,N_1401);
nand U1940 (N_1940,N_1420,N_1381);
nor U1941 (N_1941,N_1644,N_1708);
nand U1942 (N_1942,N_1795,N_1319);
xnor U1943 (N_1943,N_1713,N_1453);
nand U1944 (N_1944,N_1287,N_1442);
nand U1945 (N_1945,N_1750,N_1408);
nand U1946 (N_1946,N_1487,N_1249);
nor U1947 (N_1947,N_1397,N_1706);
and U1948 (N_1948,N_1270,N_1303);
and U1949 (N_1949,N_1645,N_1548);
and U1950 (N_1950,N_1455,N_1635);
nor U1951 (N_1951,N_1727,N_1703);
nand U1952 (N_1952,N_1384,N_1689);
and U1953 (N_1953,N_1210,N_1516);
nand U1954 (N_1954,N_1283,N_1411);
or U1955 (N_1955,N_1279,N_1463);
or U1956 (N_1956,N_1696,N_1510);
or U1957 (N_1957,N_1417,N_1509);
nand U1958 (N_1958,N_1530,N_1751);
or U1959 (N_1959,N_1775,N_1391);
nand U1960 (N_1960,N_1293,N_1264);
and U1961 (N_1961,N_1778,N_1339);
and U1962 (N_1962,N_1609,N_1620);
nand U1963 (N_1963,N_1693,N_1472);
and U1964 (N_1964,N_1528,N_1366);
xor U1965 (N_1965,N_1343,N_1668);
or U1966 (N_1966,N_1291,N_1237);
or U1967 (N_1967,N_1550,N_1670);
or U1968 (N_1968,N_1426,N_1655);
or U1969 (N_1969,N_1236,N_1450);
nor U1970 (N_1970,N_1746,N_1212);
or U1971 (N_1971,N_1630,N_1262);
xnor U1972 (N_1972,N_1297,N_1796);
nand U1973 (N_1973,N_1574,N_1232);
and U1974 (N_1974,N_1271,N_1364);
nor U1975 (N_1975,N_1524,N_1331);
and U1976 (N_1976,N_1294,N_1251);
or U1977 (N_1977,N_1286,N_1351);
nand U1978 (N_1978,N_1675,N_1586);
nor U1979 (N_1979,N_1731,N_1529);
nand U1980 (N_1980,N_1242,N_1266);
nor U1981 (N_1981,N_1377,N_1387);
and U1982 (N_1982,N_1496,N_1633);
and U1983 (N_1983,N_1648,N_1519);
nor U1984 (N_1984,N_1440,N_1711);
or U1985 (N_1985,N_1468,N_1313);
xnor U1986 (N_1986,N_1445,N_1513);
nand U1987 (N_1987,N_1758,N_1642);
and U1988 (N_1988,N_1203,N_1616);
and U1989 (N_1989,N_1308,N_1636);
and U1990 (N_1990,N_1451,N_1260);
nand U1991 (N_1991,N_1240,N_1687);
and U1992 (N_1992,N_1288,N_1485);
and U1993 (N_1993,N_1362,N_1419);
or U1994 (N_1994,N_1394,N_1480);
nand U1995 (N_1995,N_1626,N_1641);
and U1996 (N_1996,N_1733,N_1592);
or U1997 (N_1997,N_1233,N_1784);
nor U1998 (N_1998,N_1471,N_1720);
nor U1999 (N_1999,N_1600,N_1628);
xor U2000 (N_2000,N_1612,N_1571);
xnor U2001 (N_2001,N_1213,N_1667);
or U2002 (N_2002,N_1446,N_1573);
nand U2003 (N_2003,N_1730,N_1632);
or U2004 (N_2004,N_1749,N_1316);
nand U2005 (N_2005,N_1470,N_1441);
xnor U2006 (N_2006,N_1704,N_1634);
and U2007 (N_2007,N_1651,N_1718);
xor U2008 (N_2008,N_1765,N_1244);
and U2009 (N_2009,N_1761,N_1448);
and U2010 (N_2010,N_1473,N_1567);
or U2011 (N_2011,N_1278,N_1776);
or U2012 (N_2012,N_1591,N_1594);
and U2013 (N_2013,N_1685,N_1298);
nand U2014 (N_2014,N_1743,N_1798);
xnor U2015 (N_2015,N_1767,N_1660);
nor U2016 (N_2016,N_1434,N_1785);
or U2017 (N_2017,N_1547,N_1610);
and U2018 (N_2018,N_1676,N_1248);
nor U2019 (N_2019,N_1654,N_1254);
nor U2020 (N_2020,N_1692,N_1789);
or U2021 (N_2021,N_1324,N_1341);
and U2022 (N_2022,N_1476,N_1422);
nor U2023 (N_2023,N_1272,N_1340);
nor U2024 (N_2024,N_1208,N_1321);
nor U2025 (N_2025,N_1756,N_1301);
nor U2026 (N_2026,N_1725,N_1793);
nand U2027 (N_2027,N_1261,N_1425);
nor U2028 (N_2028,N_1532,N_1289);
nand U2029 (N_2029,N_1614,N_1428);
nor U2030 (N_2030,N_1281,N_1555);
and U2031 (N_2031,N_1358,N_1691);
nand U2032 (N_2032,N_1443,N_1722);
and U2033 (N_2033,N_1493,N_1439);
or U2034 (N_2034,N_1622,N_1712);
nand U2035 (N_2035,N_1412,N_1597);
xnor U2036 (N_2036,N_1538,N_1717);
or U2037 (N_2037,N_1540,N_1375);
and U2038 (N_2038,N_1762,N_1433);
or U2039 (N_2039,N_1370,N_1707);
or U2040 (N_2040,N_1256,N_1604);
nor U2041 (N_2041,N_1562,N_1680);
or U2042 (N_2042,N_1452,N_1239);
xnor U2043 (N_2043,N_1582,N_1216);
nor U2044 (N_2044,N_1307,N_1380);
and U2045 (N_2045,N_1334,N_1306);
and U2046 (N_2046,N_1678,N_1205);
or U2047 (N_2047,N_1253,N_1605);
or U2048 (N_2048,N_1652,N_1570);
nor U2049 (N_2049,N_1786,N_1520);
nor U2050 (N_2050,N_1766,N_1558);
and U2051 (N_2051,N_1247,N_1770);
or U2052 (N_2052,N_1282,N_1526);
or U2053 (N_2053,N_1593,N_1739);
nand U2054 (N_2054,N_1400,N_1561);
and U2055 (N_2055,N_1514,N_1222);
nand U2056 (N_2056,N_1486,N_1740);
and U2057 (N_2057,N_1399,N_1490);
or U2058 (N_2058,N_1523,N_1456);
nand U2059 (N_2059,N_1407,N_1543);
xor U2060 (N_2060,N_1673,N_1598);
nand U2061 (N_2061,N_1304,N_1531);
and U2062 (N_2062,N_1606,N_1782);
and U2063 (N_2063,N_1799,N_1724);
xnor U2064 (N_2064,N_1268,N_1259);
nor U2065 (N_2065,N_1230,N_1241);
and U2066 (N_2066,N_1403,N_1787);
nor U2067 (N_2067,N_1511,N_1326);
nor U2068 (N_2068,N_1276,N_1659);
and U2069 (N_2069,N_1382,N_1363);
nor U2070 (N_2070,N_1714,N_1227);
nor U2071 (N_2071,N_1245,N_1702);
and U2072 (N_2072,N_1284,N_1409);
or U2073 (N_2073,N_1719,N_1325);
or U2074 (N_2074,N_1360,N_1623);
nand U2075 (N_2075,N_1431,N_1587);
or U2076 (N_2076,N_1342,N_1554);
nand U2077 (N_2077,N_1215,N_1578);
nand U2078 (N_2078,N_1791,N_1539);
and U2079 (N_2079,N_1280,N_1768);
and U2080 (N_2080,N_1506,N_1624);
nor U2081 (N_2081,N_1424,N_1777);
nor U2082 (N_2082,N_1444,N_1560);
and U2083 (N_2083,N_1368,N_1732);
nand U2084 (N_2084,N_1501,N_1228);
and U2085 (N_2085,N_1534,N_1637);
or U2086 (N_2086,N_1551,N_1497);
or U2087 (N_2087,N_1314,N_1556);
nor U2088 (N_2088,N_1355,N_1607);
and U2089 (N_2089,N_1525,N_1618);
nor U2090 (N_2090,N_1619,N_1575);
and U2091 (N_2091,N_1211,N_1258);
nand U2092 (N_2092,N_1376,N_1688);
nand U2093 (N_2093,N_1588,N_1769);
xor U2094 (N_2094,N_1398,N_1533);
or U2095 (N_2095,N_1596,N_1477);
and U2096 (N_2096,N_1581,N_1207);
and U2097 (N_2097,N_1728,N_1764);
nand U2098 (N_2098,N_1352,N_1459);
nand U2099 (N_2099,N_1269,N_1435);
and U2100 (N_2100,N_1637,N_1565);
and U2101 (N_2101,N_1411,N_1337);
nand U2102 (N_2102,N_1583,N_1799);
nand U2103 (N_2103,N_1326,N_1518);
and U2104 (N_2104,N_1360,N_1446);
nand U2105 (N_2105,N_1571,N_1613);
nor U2106 (N_2106,N_1745,N_1748);
nand U2107 (N_2107,N_1259,N_1463);
and U2108 (N_2108,N_1505,N_1571);
xnor U2109 (N_2109,N_1564,N_1636);
or U2110 (N_2110,N_1728,N_1716);
or U2111 (N_2111,N_1357,N_1664);
nor U2112 (N_2112,N_1351,N_1432);
nor U2113 (N_2113,N_1322,N_1771);
or U2114 (N_2114,N_1319,N_1584);
or U2115 (N_2115,N_1687,N_1285);
nand U2116 (N_2116,N_1530,N_1239);
or U2117 (N_2117,N_1353,N_1548);
nor U2118 (N_2118,N_1432,N_1610);
or U2119 (N_2119,N_1632,N_1327);
nor U2120 (N_2120,N_1579,N_1553);
nor U2121 (N_2121,N_1256,N_1412);
nand U2122 (N_2122,N_1316,N_1571);
nand U2123 (N_2123,N_1793,N_1438);
or U2124 (N_2124,N_1285,N_1403);
nor U2125 (N_2125,N_1474,N_1627);
nand U2126 (N_2126,N_1349,N_1527);
nor U2127 (N_2127,N_1791,N_1756);
nor U2128 (N_2128,N_1789,N_1221);
and U2129 (N_2129,N_1441,N_1542);
and U2130 (N_2130,N_1220,N_1403);
nand U2131 (N_2131,N_1412,N_1625);
nand U2132 (N_2132,N_1289,N_1652);
and U2133 (N_2133,N_1607,N_1603);
or U2134 (N_2134,N_1331,N_1780);
or U2135 (N_2135,N_1508,N_1738);
nor U2136 (N_2136,N_1280,N_1501);
nand U2137 (N_2137,N_1330,N_1521);
nor U2138 (N_2138,N_1602,N_1455);
nand U2139 (N_2139,N_1280,N_1712);
nand U2140 (N_2140,N_1237,N_1695);
nand U2141 (N_2141,N_1715,N_1779);
nor U2142 (N_2142,N_1498,N_1251);
and U2143 (N_2143,N_1507,N_1496);
nor U2144 (N_2144,N_1538,N_1363);
and U2145 (N_2145,N_1236,N_1409);
nor U2146 (N_2146,N_1325,N_1764);
nor U2147 (N_2147,N_1419,N_1355);
nand U2148 (N_2148,N_1642,N_1647);
and U2149 (N_2149,N_1434,N_1432);
xnor U2150 (N_2150,N_1371,N_1228);
nor U2151 (N_2151,N_1309,N_1623);
xnor U2152 (N_2152,N_1401,N_1323);
and U2153 (N_2153,N_1332,N_1439);
nand U2154 (N_2154,N_1226,N_1309);
xnor U2155 (N_2155,N_1682,N_1675);
nand U2156 (N_2156,N_1306,N_1303);
or U2157 (N_2157,N_1585,N_1459);
and U2158 (N_2158,N_1257,N_1471);
and U2159 (N_2159,N_1505,N_1789);
nor U2160 (N_2160,N_1709,N_1512);
nor U2161 (N_2161,N_1420,N_1336);
nor U2162 (N_2162,N_1494,N_1321);
nor U2163 (N_2163,N_1678,N_1564);
nand U2164 (N_2164,N_1654,N_1568);
and U2165 (N_2165,N_1620,N_1475);
nor U2166 (N_2166,N_1529,N_1623);
or U2167 (N_2167,N_1620,N_1216);
xnor U2168 (N_2168,N_1259,N_1433);
and U2169 (N_2169,N_1669,N_1633);
xnor U2170 (N_2170,N_1587,N_1652);
and U2171 (N_2171,N_1682,N_1584);
nand U2172 (N_2172,N_1528,N_1273);
and U2173 (N_2173,N_1582,N_1559);
nor U2174 (N_2174,N_1420,N_1229);
nand U2175 (N_2175,N_1258,N_1452);
nand U2176 (N_2176,N_1446,N_1436);
or U2177 (N_2177,N_1312,N_1506);
and U2178 (N_2178,N_1574,N_1360);
or U2179 (N_2179,N_1725,N_1460);
and U2180 (N_2180,N_1248,N_1666);
nand U2181 (N_2181,N_1569,N_1799);
nor U2182 (N_2182,N_1559,N_1507);
or U2183 (N_2183,N_1422,N_1744);
and U2184 (N_2184,N_1328,N_1759);
nor U2185 (N_2185,N_1371,N_1342);
nor U2186 (N_2186,N_1486,N_1797);
or U2187 (N_2187,N_1239,N_1406);
or U2188 (N_2188,N_1405,N_1291);
nand U2189 (N_2189,N_1765,N_1276);
and U2190 (N_2190,N_1322,N_1703);
nand U2191 (N_2191,N_1766,N_1427);
or U2192 (N_2192,N_1251,N_1540);
or U2193 (N_2193,N_1287,N_1593);
and U2194 (N_2194,N_1379,N_1421);
nor U2195 (N_2195,N_1312,N_1387);
nand U2196 (N_2196,N_1231,N_1306);
nand U2197 (N_2197,N_1659,N_1682);
nand U2198 (N_2198,N_1541,N_1229);
nor U2199 (N_2199,N_1223,N_1335);
nor U2200 (N_2200,N_1234,N_1239);
xnor U2201 (N_2201,N_1225,N_1201);
nand U2202 (N_2202,N_1224,N_1707);
nor U2203 (N_2203,N_1450,N_1305);
and U2204 (N_2204,N_1320,N_1215);
nor U2205 (N_2205,N_1365,N_1317);
nor U2206 (N_2206,N_1774,N_1544);
and U2207 (N_2207,N_1653,N_1412);
nand U2208 (N_2208,N_1478,N_1640);
or U2209 (N_2209,N_1412,N_1337);
nand U2210 (N_2210,N_1653,N_1313);
or U2211 (N_2211,N_1348,N_1730);
or U2212 (N_2212,N_1468,N_1400);
or U2213 (N_2213,N_1326,N_1232);
or U2214 (N_2214,N_1650,N_1656);
or U2215 (N_2215,N_1239,N_1211);
and U2216 (N_2216,N_1783,N_1640);
nor U2217 (N_2217,N_1659,N_1393);
nand U2218 (N_2218,N_1301,N_1399);
and U2219 (N_2219,N_1341,N_1695);
nand U2220 (N_2220,N_1340,N_1260);
xor U2221 (N_2221,N_1558,N_1753);
nand U2222 (N_2222,N_1475,N_1284);
nand U2223 (N_2223,N_1717,N_1238);
nor U2224 (N_2224,N_1503,N_1677);
or U2225 (N_2225,N_1357,N_1383);
or U2226 (N_2226,N_1584,N_1791);
or U2227 (N_2227,N_1407,N_1553);
nor U2228 (N_2228,N_1515,N_1346);
nand U2229 (N_2229,N_1313,N_1561);
nand U2230 (N_2230,N_1543,N_1270);
and U2231 (N_2231,N_1362,N_1373);
or U2232 (N_2232,N_1710,N_1286);
or U2233 (N_2233,N_1662,N_1731);
xor U2234 (N_2234,N_1573,N_1486);
or U2235 (N_2235,N_1553,N_1670);
and U2236 (N_2236,N_1481,N_1554);
nor U2237 (N_2237,N_1467,N_1769);
nor U2238 (N_2238,N_1352,N_1592);
xnor U2239 (N_2239,N_1536,N_1280);
nor U2240 (N_2240,N_1461,N_1543);
nand U2241 (N_2241,N_1393,N_1376);
nand U2242 (N_2242,N_1641,N_1593);
nor U2243 (N_2243,N_1320,N_1206);
and U2244 (N_2244,N_1738,N_1278);
nand U2245 (N_2245,N_1218,N_1703);
nand U2246 (N_2246,N_1386,N_1403);
nor U2247 (N_2247,N_1693,N_1421);
nor U2248 (N_2248,N_1381,N_1292);
nand U2249 (N_2249,N_1520,N_1730);
nand U2250 (N_2250,N_1273,N_1540);
nand U2251 (N_2251,N_1624,N_1555);
xnor U2252 (N_2252,N_1347,N_1758);
xor U2253 (N_2253,N_1713,N_1228);
or U2254 (N_2254,N_1414,N_1666);
nand U2255 (N_2255,N_1640,N_1633);
nand U2256 (N_2256,N_1519,N_1319);
and U2257 (N_2257,N_1352,N_1618);
xor U2258 (N_2258,N_1341,N_1454);
nor U2259 (N_2259,N_1649,N_1518);
or U2260 (N_2260,N_1757,N_1279);
and U2261 (N_2261,N_1661,N_1440);
or U2262 (N_2262,N_1287,N_1449);
nor U2263 (N_2263,N_1649,N_1324);
and U2264 (N_2264,N_1493,N_1720);
nand U2265 (N_2265,N_1334,N_1456);
xor U2266 (N_2266,N_1609,N_1411);
nor U2267 (N_2267,N_1617,N_1422);
or U2268 (N_2268,N_1263,N_1260);
or U2269 (N_2269,N_1722,N_1424);
and U2270 (N_2270,N_1518,N_1319);
nand U2271 (N_2271,N_1248,N_1706);
and U2272 (N_2272,N_1658,N_1206);
or U2273 (N_2273,N_1656,N_1678);
nor U2274 (N_2274,N_1693,N_1488);
nor U2275 (N_2275,N_1632,N_1287);
nand U2276 (N_2276,N_1358,N_1653);
nor U2277 (N_2277,N_1641,N_1345);
nor U2278 (N_2278,N_1238,N_1212);
nor U2279 (N_2279,N_1321,N_1623);
nand U2280 (N_2280,N_1406,N_1209);
nor U2281 (N_2281,N_1343,N_1722);
and U2282 (N_2282,N_1761,N_1624);
nor U2283 (N_2283,N_1267,N_1749);
nor U2284 (N_2284,N_1222,N_1789);
or U2285 (N_2285,N_1552,N_1240);
or U2286 (N_2286,N_1691,N_1649);
nand U2287 (N_2287,N_1277,N_1787);
nor U2288 (N_2288,N_1621,N_1744);
nand U2289 (N_2289,N_1578,N_1355);
and U2290 (N_2290,N_1646,N_1337);
or U2291 (N_2291,N_1691,N_1654);
nor U2292 (N_2292,N_1507,N_1265);
nand U2293 (N_2293,N_1766,N_1521);
and U2294 (N_2294,N_1656,N_1553);
and U2295 (N_2295,N_1565,N_1487);
and U2296 (N_2296,N_1208,N_1481);
and U2297 (N_2297,N_1739,N_1328);
or U2298 (N_2298,N_1561,N_1696);
nand U2299 (N_2299,N_1722,N_1516);
nor U2300 (N_2300,N_1262,N_1674);
or U2301 (N_2301,N_1538,N_1728);
or U2302 (N_2302,N_1653,N_1462);
or U2303 (N_2303,N_1302,N_1547);
and U2304 (N_2304,N_1688,N_1399);
nor U2305 (N_2305,N_1721,N_1381);
or U2306 (N_2306,N_1460,N_1750);
or U2307 (N_2307,N_1239,N_1278);
nand U2308 (N_2308,N_1358,N_1792);
nand U2309 (N_2309,N_1252,N_1552);
nand U2310 (N_2310,N_1342,N_1399);
nand U2311 (N_2311,N_1610,N_1753);
xnor U2312 (N_2312,N_1363,N_1530);
nand U2313 (N_2313,N_1240,N_1706);
or U2314 (N_2314,N_1289,N_1572);
and U2315 (N_2315,N_1356,N_1583);
or U2316 (N_2316,N_1292,N_1643);
or U2317 (N_2317,N_1242,N_1648);
nor U2318 (N_2318,N_1674,N_1686);
nand U2319 (N_2319,N_1774,N_1682);
or U2320 (N_2320,N_1301,N_1531);
or U2321 (N_2321,N_1427,N_1254);
nand U2322 (N_2322,N_1416,N_1407);
nand U2323 (N_2323,N_1625,N_1291);
xor U2324 (N_2324,N_1355,N_1300);
and U2325 (N_2325,N_1683,N_1511);
and U2326 (N_2326,N_1595,N_1622);
nor U2327 (N_2327,N_1588,N_1790);
nand U2328 (N_2328,N_1583,N_1375);
nor U2329 (N_2329,N_1295,N_1623);
nand U2330 (N_2330,N_1527,N_1219);
or U2331 (N_2331,N_1704,N_1620);
or U2332 (N_2332,N_1292,N_1234);
nand U2333 (N_2333,N_1517,N_1333);
nand U2334 (N_2334,N_1443,N_1589);
and U2335 (N_2335,N_1440,N_1275);
and U2336 (N_2336,N_1484,N_1364);
and U2337 (N_2337,N_1797,N_1737);
and U2338 (N_2338,N_1313,N_1384);
nor U2339 (N_2339,N_1518,N_1260);
or U2340 (N_2340,N_1459,N_1387);
or U2341 (N_2341,N_1338,N_1698);
or U2342 (N_2342,N_1331,N_1249);
and U2343 (N_2343,N_1452,N_1779);
nand U2344 (N_2344,N_1425,N_1245);
nand U2345 (N_2345,N_1411,N_1397);
nand U2346 (N_2346,N_1433,N_1319);
or U2347 (N_2347,N_1294,N_1541);
or U2348 (N_2348,N_1712,N_1460);
xnor U2349 (N_2349,N_1347,N_1310);
nand U2350 (N_2350,N_1409,N_1449);
nand U2351 (N_2351,N_1478,N_1484);
and U2352 (N_2352,N_1780,N_1222);
and U2353 (N_2353,N_1298,N_1295);
xnor U2354 (N_2354,N_1520,N_1311);
nand U2355 (N_2355,N_1776,N_1536);
nand U2356 (N_2356,N_1406,N_1336);
nor U2357 (N_2357,N_1609,N_1396);
nor U2358 (N_2358,N_1347,N_1717);
nor U2359 (N_2359,N_1445,N_1491);
nor U2360 (N_2360,N_1342,N_1585);
and U2361 (N_2361,N_1393,N_1200);
or U2362 (N_2362,N_1226,N_1413);
and U2363 (N_2363,N_1490,N_1509);
and U2364 (N_2364,N_1320,N_1723);
and U2365 (N_2365,N_1490,N_1563);
nor U2366 (N_2366,N_1422,N_1385);
or U2367 (N_2367,N_1351,N_1655);
xor U2368 (N_2368,N_1362,N_1778);
or U2369 (N_2369,N_1477,N_1298);
and U2370 (N_2370,N_1453,N_1704);
nand U2371 (N_2371,N_1496,N_1740);
xnor U2372 (N_2372,N_1790,N_1728);
nand U2373 (N_2373,N_1621,N_1665);
xor U2374 (N_2374,N_1328,N_1274);
and U2375 (N_2375,N_1703,N_1583);
and U2376 (N_2376,N_1449,N_1690);
nor U2377 (N_2377,N_1243,N_1472);
nand U2378 (N_2378,N_1449,N_1650);
and U2379 (N_2379,N_1341,N_1274);
nor U2380 (N_2380,N_1778,N_1502);
or U2381 (N_2381,N_1528,N_1731);
nor U2382 (N_2382,N_1450,N_1276);
and U2383 (N_2383,N_1496,N_1684);
nand U2384 (N_2384,N_1503,N_1257);
or U2385 (N_2385,N_1258,N_1643);
nand U2386 (N_2386,N_1748,N_1466);
nor U2387 (N_2387,N_1397,N_1276);
and U2388 (N_2388,N_1384,N_1771);
or U2389 (N_2389,N_1533,N_1422);
nor U2390 (N_2390,N_1462,N_1435);
nor U2391 (N_2391,N_1731,N_1753);
xnor U2392 (N_2392,N_1375,N_1688);
nor U2393 (N_2393,N_1390,N_1210);
or U2394 (N_2394,N_1355,N_1580);
xor U2395 (N_2395,N_1587,N_1699);
or U2396 (N_2396,N_1613,N_1730);
nor U2397 (N_2397,N_1263,N_1325);
or U2398 (N_2398,N_1438,N_1400);
nand U2399 (N_2399,N_1631,N_1703);
nand U2400 (N_2400,N_1925,N_2385);
and U2401 (N_2401,N_2386,N_2067);
xor U2402 (N_2402,N_1808,N_2027);
nor U2403 (N_2403,N_1974,N_1943);
and U2404 (N_2404,N_2173,N_1989);
or U2405 (N_2405,N_2307,N_1886);
or U2406 (N_2406,N_2202,N_2155);
xnor U2407 (N_2407,N_2298,N_2250);
nor U2408 (N_2408,N_2085,N_2261);
nand U2409 (N_2409,N_1957,N_1815);
or U2410 (N_2410,N_2382,N_2257);
nor U2411 (N_2411,N_2118,N_2256);
or U2412 (N_2412,N_2328,N_2235);
or U2413 (N_2413,N_2295,N_1954);
nor U2414 (N_2414,N_1802,N_2144);
nand U2415 (N_2415,N_2127,N_2342);
nor U2416 (N_2416,N_2076,N_2052);
or U2417 (N_2417,N_2077,N_2188);
nand U2418 (N_2418,N_2061,N_2143);
nand U2419 (N_2419,N_2294,N_2166);
and U2420 (N_2420,N_2090,N_1910);
nand U2421 (N_2421,N_1934,N_2017);
xor U2422 (N_2422,N_2392,N_2369);
and U2423 (N_2423,N_1884,N_2245);
xnor U2424 (N_2424,N_2259,N_2169);
or U2425 (N_2425,N_2038,N_2163);
or U2426 (N_2426,N_2180,N_2326);
nor U2427 (N_2427,N_2226,N_2372);
nor U2428 (N_2428,N_1882,N_2082);
or U2429 (N_2429,N_1898,N_2216);
or U2430 (N_2430,N_2160,N_2083);
or U2431 (N_2431,N_2252,N_2394);
nor U2432 (N_2432,N_1847,N_2348);
and U2433 (N_2433,N_1869,N_2133);
or U2434 (N_2434,N_2079,N_1819);
or U2435 (N_2435,N_1897,N_2305);
or U2436 (N_2436,N_2345,N_2352);
nor U2437 (N_2437,N_2177,N_2266);
or U2438 (N_2438,N_2219,N_2005);
and U2439 (N_2439,N_2162,N_2350);
and U2440 (N_2440,N_1951,N_1827);
nand U2441 (N_2441,N_2103,N_2130);
and U2442 (N_2442,N_2335,N_1903);
or U2443 (N_2443,N_2058,N_2265);
xnor U2444 (N_2444,N_1929,N_1811);
or U2445 (N_2445,N_2009,N_1876);
or U2446 (N_2446,N_2013,N_1829);
and U2447 (N_2447,N_2281,N_2290);
nand U2448 (N_2448,N_2224,N_2153);
nand U2449 (N_2449,N_2093,N_1962);
or U2450 (N_2450,N_1896,N_1870);
nor U2451 (N_2451,N_2107,N_1953);
and U2452 (N_2452,N_2274,N_1880);
and U2453 (N_2453,N_1843,N_1950);
nand U2454 (N_2454,N_1853,N_2152);
or U2455 (N_2455,N_2264,N_2109);
nor U2456 (N_2456,N_1986,N_2278);
and U2457 (N_2457,N_2210,N_1995);
or U2458 (N_2458,N_2240,N_2388);
or U2459 (N_2459,N_2293,N_1997);
nand U2460 (N_2460,N_1902,N_2129);
xnor U2461 (N_2461,N_2139,N_2039);
nand U2462 (N_2462,N_2128,N_2306);
and U2463 (N_2463,N_2292,N_2228);
or U2464 (N_2464,N_1959,N_1981);
nor U2465 (N_2465,N_1883,N_1970);
or U2466 (N_2466,N_2304,N_1872);
nor U2467 (N_2467,N_1801,N_1837);
or U2468 (N_2468,N_1972,N_2189);
nand U2469 (N_2469,N_2333,N_2172);
nand U2470 (N_2470,N_2008,N_1961);
nor U2471 (N_2471,N_2339,N_1823);
or U2472 (N_2472,N_2181,N_2313);
or U2473 (N_2473,N_1889,N_2159);
xnor U2474 (N_2474,N_2195,N_1831);
nor U2475 (N_2475,N_1844,N_1894);
nor U2476 (N_2476,N_1949,N_2078);
nor U2477 (N_2477,N_1914,N_2343);
or U2478 (N_2478,N_2193,N_2336);
nor U2479 (N_2479,N_2065,N_2098);
and U2480 (N_2480,N_2056,N_2397);
nand U2481 (N_2481,N_2223,N_1963);
or U2482 (N_2482,N_2393,N_1906);
nand U2483 (N_2483,N_1893,N_1860);
and U2484 (N_2484,N_2330,N_1965);
xnor U2485 (N_2485,N_1968,N_1891);
nor U2486 (N_2486,N_2251,N_1817);
and U2487 (N_2487,N_2302,N_1851);
and U2488 (N_2488,N_2080,N_1887);
and U2489 (N_2489,N_2001,N_2040);
and U2490 (N_2490,N_2066,N_2045);
xor U2491 (N_2491,N_2316,N_2248);
nand U2492 (N_2492,N_2332,N_1861);
nand U2493 (N_2493,N_2064,N_1878);
and U2494 (N_2494,N_2222,N_2019);
or U2495 (N_2495,N_2396,N_2267);
and U2496 (N_2496,N_1879,N_2362);
nor U2497 (N_2497,N_2011,N_2087);
nor U2498 (N_2498,N_2042,N_2214);
nand U2499 (N_2499,N_2327,N_1885);
or U2500 (N_2500,N_2032,N_1911);
and U2501 (N_2501,N_2025,N_2174);
and U2502 (N_2502,N_2241,N_2319);
nand U2503 (N_2503,N_1900,N_2363);
nand U2504 (N_2504,N_2340,N_2341);
xor U2505 (N_2505,N_2218,N_1812);
nand U2506 (N_2506,N_1818,N_2104);
and U2507 (N_2507,N_2288,N_1816);
and U2508 (N_2508,N_2387,N_2373);
and U2509 (N_2509,N_2151,N_1932);
nand U2510 (N_2510,N_2137,N_2131);
nor U2511 (N_2511,N_2198,N_1945);
xnor U2512 (N_2512,N_1840,N_1998);
and U2513 (N_2513,N_2311,N_2310);
and U2514 (N_2514,N_1821,N_1971);
and U2515 (N_2515,N_2075,N_2149);
nand U2516 (N_2516,N_2207,N_2255);
or U2517 (N_2517,N_1824,N_1807);
xnor U2518 (N_2518,N_2360,N_2334);
nor U2519 (N_2519,N_2054,N_1994);
nand U2520 (N_2520,N_1928,N_2285);
nor U2521 (N_2521,N_2110,N_1852);
or U2522 (N_2522,N_1947,N_2119);
nor U2523 (N_2523,N_2141,N_2276);
nor U2524 (N_2524,N_1996,N_1931);
and U2525 (N_2525,N_2263,N_1956);
or U2526 (N_2526,N_1867,N_2308);
and U2527 (N_2527,N_2003,N_2035);
nor U2528 (N_2528,N_2351,N_1993);
and U2529 (N_2529,N_2323,N_2068);
nor U2530 (N_2530,N_2134,N_2186);
xor U2531 (N_2531,N_2002,N_2142);
and U2532 (N_2532,N_1944,N_2192);
and U2533 (N_2533,N_2246,N_2273);
xnor U2534 (N_2534,N_2121,N_2026);
or U2535 (N_2535,N_1841,N_1845);
nor U2536 (N_2536,N_1985,N_2349);
nand U2537 (N_2537,N_2242,N_1913);
nor U2538 (N_2538,N_1864,N_2234);
xnor U2539 (N_2539,N_2049,N_2395);
nor U2540 (N_2540,N_2232,N_2378);
or U2541 (N_2541,N_2309,N_2043);
and U2542 (N_2542,N_2175,N_2329);
nand U2543 (N_2543,N_2170,N_2016);
or U2544 (N_2544,N_2380,N_1806);
nor U2545 (N_2545,N_2081,N_2086);
nor U2546 (N_2546,N_2070,N_1948);
xnor U2547 (N_2547,N_1909,N_1923);
and U2548 (N_2548,N_2154,N_1834);
or U2549 (N_2549,N_1854,N_2106);
or U2550 (N_2550,N_2053,N_2007);
nor U2551 (N_2551,N_1892,N_2355);
nand U2552 (N_2552,N_2073,N_2354);
xnor U2553 (N_2553,N_1828,N_1877);
nand U2554 (N_2554,N_2145,N_2091);
nor U2555 (N_2555,N_2205,N_2321);
nand U2556 (N_2556,N_1939,N_2074);
nor U2557 (N_2557,N_2185,N_1836);
and U2558 (N_2558,N_2022,N_2399);
nand U2559 (N_2559,N_2200,N_2184);
nand U2560 (N_2560,N_2209,N_2168);
nand U2561 (N_2561,N_1918,N_2359);
and U2562 (N_2562,N_2315,N_1838);
and U2563 (N_2563,N_1935,N_2215);
or U2564 (N_2564,N_2100,N_2024);
nor U2565 (N_2565,N_2135,N_1936);
nand U2566 (N_2566,N_2227,N_2201);
nand U2567 (N_2567,N_2262,N_2161);
nand U2568 (N_2568,N_1907,N_2037);
nand U2569 (N_2569,N_1940,N_1865);
nor U2570 (N_2570,N_2368,N_2033);
and U2571 (N_2571,N_2178,N_2249);
and U2572 (N_2572,N_2004,N_2239);
and U2573 (N_2573,N_1966,N_1875);
nand U2574 (N_2574,N_2020,N_2071);
or U2575 (N_2575,N_1976,N_1983);
or U2576 (N_2576,N_1855,N_2046);
nand U2577 (N_2577,N_2088,N_1846);
and U2578 (N_2578,N_2113,N_2253);
or U2579 (N_2579,N_2112,N_2099);
and U2580 (N_2580,N_2283,N_1857);
xnor U2581 (N_2581,N_2057,N_2125);
nor U2582 (N_2582,N_1924,N_1895);
or U2583 (N_2583,N_2034,N_1922);
and U2584 (N_2584,N_2398,N_2094);
nor U2585 (N_2585,N_2158,N_2062);
and U2586 (N_2586,N_2296,N_2196);
nor U2587 (N_2587,N_1941,N_2291);
nor U2588 (N_2588,N_2370,N_1830);
nor U2589 (N_2589,N_2018,N_2182);
and U2590 (N_2590,N_1826,N_2059);
and U2591 (N_2591,N_2164,N_1871);
nand U2592 (N_2592,N_1952,N_1930);
or U2593 (N_2593,N_2299,N_2337);
xor U2594 (N_2594,N_1937,N_2318);
and U2595 (N_2595,N_2041,N_2006);
or U2596 (N_2596,N_2084,N_2167);
and U2597 (N_2597,N_1866,N_2117);
and U2598 (N_2598,N_2147,N_2187);
nand U2599 (N_2599,N_2384,N_1958);
xnor U2600 (N_2600,N_1863,N_2156);
xor U2601 (N_2601,N_1967,N_2030);
and U2602 (N_2602,N_2199,N_2126);
or U2603 (N_2603,N_2021,N_2069);
nor U2604 (N_2604,N_1835,N_1964);
nand U2605 (N_2605,N_2051,N_2095);
nand U2606 (N_2606,N_2277,N_2374);
and U2607 (N_2607,N_2371,N_2092);
and U2608 (N_2608,N_1955,N_2116);
and U2609 (N_2609,N_1848,N_2282);
and U2610 (N_2610,N_2270,N_2271);
nor U2611 (N_2611,N_2375,N_2379);
nor U2612 (N_2612,N_1987,N_1946);
nand U2613 (N_2613,N_2260,N_1977);
or U2614 (N_2614,N_1908,N_2317);
nor U2615 (N_2615,N_1825,N_1919);
or U2616 (N_2616,N_2391,N_2123);
nand U2617 (N_2617,N_2225,N_2179);
nand U2618 (N_2618,N_1969,N_1990);
and U2619 (N_2619,N_2244,N_2140);
xor U2620 (N_2620,N_2269,N_2383);
and U2621 (N_2621,N_2208,N_2014);
or U2622 (N_2622,N_1978,N_2344);
and U2623 (N_2623,N_2325,N_2108);
or U2624 (N_2624,N_1984,N_2015);
nor U2625 (N_2625,N_2048,N_2365);
nand U2626 (N_2626,N_1800,N_2028);
and U2627 (N_2627,N_1804,N_2115);
and U2628 (N_2628,N_1810,N_2124);
or U2629 (N_2629,N_2314,N_1862);
nor U2630 (N_2630,N_1912,N_1999);
nand U2631 (N_2631,N_2367,N_2194);
and U2632 (N_2632,N_2203,N_2303);
or U2633 (N_2633,N_2217,N_2183);
or U2634 (N_2634,N_2247,N_2221);
xnor U2635 (N_2635,N_1980,N_1933);
and U2636 (N_2636,N_2102,N_1938);
nor U2637 (N_2637,N_1832,N_2331);
nor U2638 (N_2638,N_1988,N_1905);
and U2639 (N_2639,N_2287,N_1842);
and U2640 (N_2640,N_2204,N_2138);
or U2641 (N_2641,N_1822,N_2089);
nand U2642 (N_2642,N_2063,N_2353);
xor U2643 (N_2643,N_2000,N_1859);
nand U2644 (N_2644,N_2230,N_2389);
nand U2645 (N_2645,N_2036,N_2176);
xor U2646 (N_2646,N_1890,N_2010);
nor U2647 (N_2647,N_1820,N_2279);
nand U2648 (N_2648,N_1901,N_1916);
or U2649 (N_2649,N_1888,N_2284);
nand U2650 (N_2650,N_2072,N_2206);
xor U2651 (N_2651,N_2366,N_2324);
nand U2652 (N_2652,N_2229,N_2320);
nor U2653 (N_2653,N_2122,N_2105);
and U2654 (N_2654,N_1850,N_1813);
nand U2655 (N_2655,N_2055,N_2114);
or U2656 (N_2656,N_2212,N_1942);
nand U2657 (N_2657,N_1991,N_2044);
or U2658 (N_2658,N_2150,N_1973);
nor U2659 (N_2659,N_1917,N_2301);
or U2660 (N_2660,N_2101,N_1849);
or U2661 (N_2661,N_1805,N_2157);
or U2662 (N_2662,N_2289,N_1899);
nand U2663 (N_2663,N_1833,N_1982);
nand U2664 (N_2664,N_2233,N_2047);
or U2665 (N_2665,N_2050,N_2280);
and U2666 (N_2666,N_2390,N_2358);
and U2667 (N_2667,N_2197,N_2312);
nor U2668 (N_2668,N_2364,N_2171);
nand U2669 (N_2669,N_2237,N_2097);
and U2670 (N_2670,N_2190,N_1915);
or U2671 (N_2671,N_2213,N_2338);
nor U2672 (N_2672,N_2300,N_1992);
nor U2673 (N_2673,N_2029,N_2357);
and U2674 (N_2674,N_2377,N_2012);
or U2675 (N_2675,N_1814,N_2322);
and U2676 (N_2676,N_2136,N_1803);
and U2677 (N_2677,N_2023,N_1881);
or U2678 (N_2678,N_2120,N_2356);
and U2679 (N_2679,N_2272,N_1979);
nor U2680 (N_2680,N_1926,N_1873);
nor U2681 (N_2681,N_1927,N_1839);
nor U2682 (N_2682,N_1856,N_2381);
xor U2683 (N_2683,N_2220,N_2346);
and U2684 (N_2684,N_2165,N_2268);
xor U2685 (N_2685,N_1960,N_2146);
nor U2686 (N_2686,N_2361,N_2286);
and U2687 (N_2687,N_1975,N_2347);
and U2688 (N_2688,N_2243,N_2275);
and U2689 (N_2689,N_1868,N_2132);
or U2690 (N_2690,N_1809,N_2148);
or U2691 (N_2691,N_1874,N_2236);
nor U2692 (N_2692,N_2238,N_2258);
nor U2693 (N_2693,N_2254,N_1921);
and U2694 (N_2694,N_2231,N_2191);
or U2695 (N_2695,N_1858,N_2060);
nor U2696 (N_2696,N_2211,N_2111);
xor U2697 (N_2697,N_1920,N_2376);
and U2698 (N_2698,N_2096,N_2297);
or U2699 (N_2699,N_2031,N_1904);
xnor U2700 (N_2700,N_2225,N_1844);
or U2701 (N_2701,N_2384,N_2347);
or U2702 (N_2702,N_2388,N_2103);
xnor U2703 (N_2703,N_2124,N_1979);
nand U2704 (N_2704,N_2139,N_1848);
or U2705 (N_2705,N_2123,N_1933);
nor U2706 (N_2706,N_2237,N_2347);
or U2707 (N_2707,N_2357,N_2172);
nand U2708 (N_2708,N_2398,N_2187);
and U2709 (N_2709,N_2025,N_1944);
and U2710 (N_2710,N_2380,N_2332);
xor U2711 (N_2711,N_1875,N_1832);
and U2712 (N_2712,N_1814,N_2238);
nor U2713 (N_2713,N_1918,N_2000);
nand U2714 (N_2714,N_2119,N_2094);
nor U2715 (N_2715,N_2257,N_2005);
and U2716 (N_2716,N_2057,N_1912);
and U2717 (N_2717,N_2357,N_1800);
or U2718 (N_2718,N_2141,N_1816);
and U2719 (N_2719,N_2024,N_2032);
and U2720 (N_2720,N_1805,N_2197);
xor U2721 (N_2721,N_2086,N_2038);
nand U2722 (N_2722,N_2032,N_2185);
nor U2723 (N_2723,N_1937,N_1883);
nor U2724 (N_2724,N_2097,N_1934);
and U2725 (N_2725,N_1929,N_2332);
or U2726 (N_2726,N_2323,N_2339);
nor U2727 (N_2727,N_2221,N_1993);
nand U2728 (N_2728,N_2323,N_2030);
nand U2729 (N_2729,N_1865,N_1859);
nor U2730 (N_2730,N_2075,N_2030);
nor U2731 (N_2731,N_2147,N_2349);
and U2732 (N_2732,N_2372,N_1954);
and U2733 (N_2733,N_2036,N_1842);
nand U2734 (N_2734,N_2116,N_2304);
and U2735 (N_2735,N_2384,N_1899);
and U2736 (N_2736,N_1933,N_2256);
xor U2737 (N_2737,N_2056,N_1941);
nor U2738 (N_2738,N_1955,N_2256);
or U2739 (N_2739,N_2003,N_2046);
and U2740 (N_2740,N_2342,N_1936);
nor U2741 (N_2741,N_1911,N_1877);
nor U2742 (N_2742,N_2004,N_2051);
and U2743 (N_2743,N_2083,N_2081);
nand U2744 (N_2744,N_2346,N_1895);
or U2745 (N_2745,N_2154,N_1814);
or U2746 (N_2746,N_2167,N_2387);
nand U2747 (N_2747,N_1959,N_1909);
nor U2748 (N_2748,N_2384,N_2081);
and U2749 (N_2749,N_2025,N_2080);
nand U2750 (N_2750,N_1913,N_1842);
or U2751 (N_2751,N_1915,N_2130);
nor U2752 (N_2752,N_1917,N_2351);
and U2753 (N_2753,N_1919,N_2193);
xnor U2754 (N_2754,N_1917,N_2370);
nor U2755 (N_2755,N_1827,N_2091);
nand U2756 (N_2756,N_1852,N_2242);
nor U2757 (N_2757,N_1942,N_2055);
nor U2758 (N_2758,N_1829,N_1803);
or U2759 (N_2759,N_2356,N_2330);
nand U2760 (N_2760,N_1815,N_2374);
or U2761 (N_2761,N_2366,N_1838);
nand U2762 (N_2762,N_2364,N_2055);
nor U2763 (N_2763,N_1869,N_1807);
or U2764 (N_2764,N_2186,N_2250);
or U2765 (N_2765,N_1970,N_1872);
or U2766 (N_2766,N_1925,N_2342);
and U2767 (N_2767,N_2251,N_2036);
or U2768 (N_2768,N_1814,N_2048);
nand U2769 (N_2769,N_2377,N_1870);
nand U2770 (N_2770,N_2132,N_2144);
nand U2771 (N_2771,N_2255,N_1880);
and U2772 (N_2772,N_2162,N_2033);
and U2773 (N_2773,N_1947,N_2177);
and U2774 (N_2774,N_2316,N_2147);
nor U2775 (N_2775,N_2339,N_2309);
xor U2776 (N_2776,N_2025,N_2223);
and U2777 (N_2777,N_2059,N_2035);
nor U2778 (N_2778,N_2191,N_2049);
nand U2779 (N_2779,N_2168,N_2225);
nor U2780 (N_2780,N_2119,N_1948);
nor U2781 (N_2781,N_1806,N_2060);
nor U2782 (N_2782,N_2368,N_2152);
and U2783 (N_2783,N_2191,N_1811);
or U2784 (N_2784,N_2052,N_2208);
nand U2785 (N_2785,N_1822,N_1819);
nand U2786 (N_2786,N_1967,N_1845);
or U2787 (N_2787,N_2232,N_2045);
or U2788 (N_2788,N_2300,N_2239);
or U2789 (N_2789,N_2326,N_2298);
or U2790 (N_2790,N_2235,N_1844);
xor U2791 (N_2791,N_2187,N_1828);
nor U2792 (N_2792,N_2327,N_2119);
nand U2793 (N_2793,N_1883,N_2158);
nand U2794 (N_2794,N_2176,N_2311);
nand U2795 (N_2795,N_2102,N_2057);
and U2796 (N_2796,N_2042,N_2204);
nand U2797 (N_2797,N_2104,N_2182);
nor U2798 (N_2798,N_2343,N_2339);
xnor U2799 (N_2799,N_2369,N_1987);
and U2800 (N_2800,N_2197,N_2155);
and U2801 (N_2801,N_2322,N_1809);
xor U2802 (N_2802,N_2223,N_2262);
or U2803 (N_2803,N_2085,N_1817);
nand U2804 (N_2804,N_2156,N_2014);
or U2805 (N_2805,N_2083,N_2032);
or U2806 (N_2806,N_2225,N_2320);
and U2807 (N_2807,N_2244,N_1933);
xor U2808 (N_2808,N_2139,N_2142);
nand U2809 (N_2809,N_2377,N_2365);
and U2810 (N_2810,N_2073,N_2146);
xor U2811 (N_2811,N_2295,N_1942);
and U2812 (N_2812,N_1843,N_2096);
and U2813 (N_2813,N_2338,N_1905);
or U2814 (N_2814,N_2234,N_1926);
or U2815 (N_2815,N_2148,N_2023);
nor U2816 (N_2816,N_1834,N_2004);
and U2817 (N_2817,N_1879,N_2359);
nor U2818 (N_2818,N_2179,N_2054);
nor U2819 (N_2819,N_2175,N_2386);
nand U2820 (N_2820,N_2357,N_2214);
and U2821 (N_2821,N_2119,N_1942);
or U2822 (N_2822,N_2277,N_2007);
nand U2823 (N_2823,N_1875,N_2175);
or U2824 (N_2824,N_2293,N_2398);
xnor U2825 (N_2825,N_2397,N_2200);
and U2826 (N_2826,N_2158,N_1974);
nor U2827 (N_2827,N_2038,N_2368);
nor U2828 (N_2828,N_2136,N_2360);
and U2829 (N_2829,N_1993,N_2275);
and U2830 (N_2830,N_2272,N_2302);
nand U2831 (N_2831,N_2065,N_2158);
or U2832 (N_2832,N_2260,N_2208);
or U2833 (N_2833,N_2251,N_2204);
nand U2834 (N_2834,N_1980,N_1817);
nand U2835 (N_2835,N_1845,N_1953);
or U2836 (N_2836,N_2158,N_2232);
and U2837 (N_2837,N_2352,N_2076);
and U2838 (N_2838,N_2030,N_2236);
or U2839 (N_2839,N_2032,N_2226);
nand U2840 (N_2840,N_2319,N_2361);
xnor U2841 (N_2841,N_2281,N_2239);
nand U2842 (N_2842,N_2079,N_1859);
and U2843 (N_2843,N_2382,N_2183);
nor U2844 (N_2844,N_2353,N_2265);
or U2845 (N_2845,N_2191,N_2051);
and U2846 (N_2846,N_2240,N_1824);
and U2847 (N_2847,N_2333,N_2289);
xor U2848 (N_2848,N_2279,N_2281);
nand U2849 (N_2849,N_2360,N_2176);
nor U2850 (N_2850,N_2265,N_1895);
or U2851 (N_2851,N_2144,N_2317);
or U2852 (N_2852,N_2055,N_2350);
nand U2853 (N_2853,N_2328,N_2311);
xor U2854 (N_2854,N_1970,N_2283);
nor U2855 (N_2855,N_2166,N_2377);
nor U2856 (N_2856,N_2210,N_1885);
or U2857 (N_2857,N_1854,N_2166);
nor U2858 (N_2858,N_2376,N_2136);
nor U2859 (N_2859,N_2297,N_1807);
nor U2860 (N_2860,N_1911,N_2231);
and U2861 (N_2861,N_1845,N_1822);
nand U2862 (N_2862,N_2272,N_2368);
and U2863 (N_2863,N_1804,N_1812);
nor U2864 (N_2864,N_2186,N_1848);
and U2865 (N_2865,N_2323,N_1808);
nor U2866 (N_2866,N_2350,N_2136);
nor U2867 (N_2867,N_2128,N_2167);
nand U2868 (N_2868,N_1802,N_2207);
and U2869 (N_2869,N_2277,N_1842);
nor U2870 (N_2870,N_2178,N_2395);
nor U2871 (N_2871,N_2226,N_2090);
nor U2872 (N_2872,N_2111,N_1895);
nor U2873 (N_2873,N_2060,N_2048);
nor U2874 (N_2874,N_2371,N_2134);
nor U2875 (N_2875,N_1920,N_2224);
nand U2876 (N_2876,N_2366,N_1964);
nor U2877 (N_2877,N_1840,N_2319);
xnor U2878 (N_2878,N_2119,N_2295);
nor U2879 (N_2879,N_1961,N_2176);
nand U2880 (N_2880,N_2127,N_2132);
and U2881 (N_2881,N_2210,N_2130);
and U2882 (N_2882,N_1834,N_2015);
and U2883 (N_2883,N_2104,N_1937);
xor U2884 (N_2884,N_1840,N_1932);
or U2885 (N_2885,N_1836,N_1823);
and U2886 (N_2886,N_1868,N_2114);
nand U2887 (N_2887,N_1912,N_2360);
nor U2888 (N_2888,N_1820,N_2218);
and U2889 (N_2889,N_2108,N_2384);
and U2890 (N_2890,N_2021,N_2379);
and U2891 (N_2891,N_2161,N_2090);
nand U2892 (N_2892,N_1942,N_2299);
nor U2893 (N_2893,N_2199,N_2247);
xnor U2894 (N_2894,N_2060,N_2153);
xnor U2895 (N_2895,N_1815,N_2248);
or U2896 (N_2896,N_2211,N_2253);
nor U2897 (N_2897,N_1940,N_2288);
or U2898 (N_2898,N_2044,N_2340);
nand U2899 (N_2899,N_1974,N_2303);
and U2900 (N_2900,N_1902,N_1949);
nor U2901 (N_2901,N_2044,N_2065);
xor U2902 (N_2902,N_2008,N_2080);
nor U2903 (N_2903,N_2119,N_2364);
xor U2904 (N_2904,N_1946,N_2017);
nand U2905 (N_2905,N_1998,N_2070);
or U2906 (N_2906,N_1974,N_2038);
nand U2907 (N_2907,N_2303,N_2015);
and U2908 (N_2908,N_2274,N_2180);
nor U2909 (N_2909,N_2362,N_2197);
and U2910 (N_2910,N_2151,N_2332);
and U2911 (N_2911,N_2379,N_2208);
or U2912 (N_2912,N_2185,N_1910);
nand U2913 (N_2913,N_2212,N_2181);
xor U2914 (N_2914,N_2291,N_2329);
nor U2915 (N_2915,N_1880,N_2154);
and U2916 (N_2916,N_2329,N_1904);
or U2917 (N_2917,N_1843,N_1898);
or U2918 (N_2918,N_2269,N_2200);
and U2919 (N_2919,N_1996,N_2363);
and U2920 (N_2920,N_2245,N_2088);
or U2921 (N_2921,N_2376,N_2249);
xnor U2922 (N_2922,N_1897,N_2395);
xor U2923 (N_2923,N_2086,N_1922);
xnor U2924 (N_2924,N_1816,N_2217);
and U2925 (N_2925,N_2016,N_2156);
xor U2926 (N_2926,N_1983,N_2372);
or U2927 (N_2927,N_1873,N_2145);
xnor U2928 (N_2928,N_2215,N_2180);
and U2929 (N_2929,N_1901,N_1970);
nand U2930 (N_2930,N_2089,N_1913);
and U2931 (N_2931,N_1878,N_2312);
or U2932 (N_2932,N_2199,N_2390);
or U2933 (N_2933,N_1953,N_1802);
or U2934 (N_2934,N_2347,N_2203);
or U2935 (N_2935,N_1918,N_1943);
and U2936 (N_2936,N_2365,N_2041);
and U2937 (N_2937,N_2358,N_1815);
xor U2938 (N_2938,N_1881,N_2121);
and U2939 (N_2939,N_2057,N_1820);
nand U2940 (N_2940,N_2254,N_2124);
nor U2941 (N_2941,N_2134,N_2031);
nand U2942 (N_2942,N_1837,N_1884);
and U2943 (N_2943,N_2332,N_2224);
and U2944 (N_2944,N_2280,N_2000);
and U2945 (N_2945,N_2087,N_2376);
nor U2946 (N_2946,N_2071,N_2316);
nand U2947 (N_2947,N_2338,N_2099);
xnor U2948 (N_2948,N_2154,N_2259);
and U2949 (N_2949,N_1990,N_1819);
nand U2950 (N_2950,N_1955,N_2391);
or U2951 (N_2951,N_1978,N_2191);
or U2952 (N_2952,N_2296,N_2113);
or U2953 (N_2953,N_1996,N_2099);
and U2954 (N_2954,N_2357,N_2021);
or U2955 (N_2955,N_2200,N_2125);
nor U2956 (N_2956,N_1830,N_1888);
and U2957 (N_2957,N_1980,N_1823);
and U2958 (N_2958,N_2161,N_1873);
and U2959 (N_2959,N_2069,N_2241);
nor U2960 (N_2960,N_2317,N_2100);
xnor U2961 (N_2961,N_2113,N_1916);
nor U2962 (N_2962,N_2166,N_2046);
nand U2963 (N_2963,N_2072,N_2018);
xnor U2964 (N_2964,N_1997,N_2296);
and U2965 (N_2965,N_2157,N_1988);
nand U2966 (N_2966,N_1906,N_2323);
nand U2967 (N_2967,N_2238,N_1989);
and U2968 (N_2968,N_2139,N_1836);
nor U2969 (N_2969,N_2268,N_2364);
xor U2970 (N_2970,N_1852,N_2346);
nand U2971 (N_2971,N_2120,N_2002);
or U2972 (N_2972,N_2092,N_2179);
or U2973 (N_2973,N_1829,N_1841);
and U2974 (N_2974,N_2088,N_2086);
nand U2975 (N_2975,N_2175,N_2071);
xnor U2976 (N_2976,N_1816,N_2111);
nand U2977 (N_2977,N_1949,N_1805);
nand U2978 (N_2978,N_1923,N_2322);
xor U2979 (N_2979,N_2016,N_2280);
and U2980 (N_2980,N_1918,N_1961);
or U2981 (N_2981,N_2157,N_2317);
nor U2982 (N_2982,N_2243,N_1806);
xor U2983 (N_2983,N_1908,N_2185);
and U2984 (N_2984,N_1973,N_2131);
nand U2985 (N_2985,N_1852,N_2131);
nor U2986 (N_2986,N_1864,N_1965);
nand U2987 (N_2987,N_2315,N_1948);
or U2988 (N_2988,N_2099,N_1931);
nand U2989 (N_2989,N_2266,N_2026);
or U2990 (N_2990,N_2109,N_1812);
nand U2991 (N_2991,N_1808,N_2180);
nand U2992 (N_2992,N_2096,N_2000);
and U2993 (N_2993,N_2283,N_2098);
nor U2994 (N_2994,N_2170,N_2166);
or U2995 (N_2995,N_1994,N_1862);
nand U2996 (N_2996,N_2358,N_2114);
nor U2997 (N_2997,N_2051,N_2206);
nand U2998 (N_2998,N_2222,N_1913);
and U2999 (N_2999,N_1978,N_2396);
or UO_0 (O_0,N_2516,N_2632);
or UO_1 (O_1,N_2693,N_2443);
nor UO_2 (O_2,N_2650,N_2688);
nor UO_3 (O_3,N_2512,N_2499);
nor UO_4 (O_4,N_2455,N_2572);
or UO_5 (O_5,N_2825,N_2964);
nor UO_6 (O_6,N_2562,N_2934);
nor UO_7 (O_7,N_2475,N_2445);
nand UO_8 (O_8,N_2916,N_2523);
or UO_9 (O_9,N_2531,N_2416);
nand UO_10 (O_10,N_2878,N_2984);
nand UO_11 (O_11,N_2413,N_2912);
and UO_12 (O_12,N_2943,N_2727);
xnor UO_13 (O_13,N_2755,N_2792);
and UO_14 (O_14,N_2468,N_2911);
nor UO_15 (O_15,N_2621,N_2567);
and UO_16 (O_16,N_2972,N_2850);
nand UO_17 (O_17,N_2954,N_2913);
or UO_18 (O_18,N_2501,N_2645);
nand UO_19 (O_19,N_2986,N_2780);
nand UO_20 (O_20,N_2919,N_2840);
and UO_21 (O_21,N_2432,N_2466);
xor UO_22 (O_22,N_2997,N_2979);
and UO_23 (O_23,N_2791,N_2842);
nor UO_24 (O_24,N_2701,N_2552);
or UO_25 (O_25,N_2960,N_2511);
or UO_26 (O_26,N_2414,N_2594);
and UO_27 (O_27,N_2870,N_2719);
nor UO_28 (O_28,N_2545,N_2444);
nand UO_29 (O_29,N_2918,N_2448);
nand UO_30 (O_30,N_2998,N_2434);
and UO_31 (O_31,N_2408,N_2564);
xnor UO_32 (O_32,N_2436,N_2660);
nor UO_33 (O_33,N_2651,N_2439);
nor UO_34 (O_34,N_2782,N_2771);
or UO_35 (O_35,N_2586,N_2542);
nand UO_36 (O_36,N_2810,N_2653);
nor UO_37 (O_37,N_2822,N_2560);
and UO_38 (O_38,N_2915,N_2988);
nor UO_39 (O_39,N_2429,N_2547);
nor UO_40 (O_40,N_2676,N_2848);
and UO_41 (O_41,N_2697,N_2415);
nand UO_42 (O_42,N_2540,N_2635);
and UO_43 (O_43,N_2607,N_2945);
and UO_44 (O_44,N_2845,N_2853);
or UO_45 (O_45,N_2775,N_2900);
or UO_46 (O_46,N_2488,N_2711);
nor UO_47 (O_47,N_2678,N_2955);
xor UO_48 (O_48,N_2601,N_2865);
or UO_49 (O_49,N_2747,N_2800);
nand UO_50 (O_50,N_2477,N_2731);
nand UO_51 (O_51,N_2734,N_2881);
nand UO_52 (O_52,N_2824,N_2721);
or UO_53 (O_53,N_2610,N_2896);
and UO_54 (O_54,N_2629,N_2811);
xor UO_55 (O_55,N_2830,N_2951);
and UO_56 (O_56,N_2876,N_2879);
and UO_57 (O_57,N_2772,N_2584);
and UO_58 (O_58,N_2626,N_2804);
or UO_59 (O_59,N_2993,N_2614);
and UO_60 (O_60,N_2835,N_2910);
nor UO_61 (O_61,N_2942,N_2941);
and UO_62 (O_62,N_2658,N_2605);
and UO_63 (O_63,N_2832,N_2464);
or UO_64 (O_64,N_2513,N_2901);
or UO_65 (O_65,N_2440,N_2519);
xnor UO_66 (O_66,N_2856,N_2553);
or UO_67 (O_67,N_2767,N_2677);
and UO_68 (O_68,N_2980,N_2597);
nand UO_69 (O_69,N_2683,N_2538);
nand UO_70 (O_70,N_2684,N_2686);
nand UO_71 (O_71,N_2574,N_2816);
and UO_72 (O_72,N_2704,N_2809);
nor UO_73 (O_73,N_2423,N_2409);
or UO_74 (O_74,N_2965,N_2863);
or UO_75 (O_75,N_2671,N_2458);
and UO_76 (O_76,N_2405,N_2999);
nor UO_77 (O_77,N_2819,N_2753);
xnor UO_78 (O_78,N_2533,N_2995);
xor UO_79 (O_79,N_2406,N_2460);
nor UO_80 (O_80,N_2425,N_2655);
nand UO_81 (O_81,N_2478,N_2583);
nor UO_82 (O_82,N_2849,N_2858);
nor UO_83 (O_83,N_2946,N_2764);
or UO_84 (O_84,N_2864,N_2505);
or UO_85 (O_85,N_2723,N_2886);
and UO_86 (O_86,N_2503,N_2426);
or UO_87 (O_87,N_2411,N_2788);
nand UO_88 (O_88,N_2467,N_2748);
nor UO_89 (O_89,N_2654,N_2939);
and UO_90 (O_90,N_2757,N_2797);
xor UO_91 (O_91,N_2469,N_2868);
and UO_92 (O_92,N_2675,N_2948);
and UO_93 (O_93,N_2599,N_2798);
or UO_94 (O_94,N_2787,N_2859);
nand UO_95 (O_95,N_2419,N_2895);
or UO_96 (O_96,N_2861,N_2717);
or UO_97 (O_97,N_2433,N_2722);
and UO_98 (O_98,N_2672,N_2867);
or UO_99 (O_99,N_2575,N_2774);
or UO_100 (O_100,N_2424,N_2839);
or UO_101 (O_101,N_2974,N_2644);
xnor UO_102 (O_102,N_2909,N_2498);
nand UO_103 (O_103,N_2493,N_2925);
or UO_104 (O_104,N_2812,N_2760);
and UO_105 (O_105,N_2823,N_2504);
nand UO_106 (O_106,N_2627,N_2446);
nor UO_107 (O_107,N_2786,N_2496);
nor UO_108 (O_108,N_2462,N_2570);
nor UO_109 (O_109,N_2520,N_2633);
nor UO_110 (O_110,N_2518,N_2818);
nor UO_111 (O_111,N_2647,N_2691);
nand UO_112 (O_112,N_2664,N_2421);
nand UO_113 (O_113,N_2831,N_2991);
and UO_114 (O_114,N_2903,N_2609);
xor UO_115 (O_115,N_2801,N_2779);
or UO_116 (O_116,N_2452,N_2931);
nor UO_117 (O_117,N_2884,N_2451);
and UO_118 (O_118,N_2481,N_2796);
or UO_119 (O_119,N_2932,N_2483);
nand UO_120 (O_120,N_2821,N_2957);
nand UO_121 (O_121,N_2793,N_2985);
and UO_122 (O_122,N_2404,N_2450);
or UO_123 (O_123,N_2714,N_2938);
nor UO_124 (O_124,N_2639,N_2625);
nor UO_125 (O_125,N_2568,N_2852);
nand UO_126 (O_126,N_2975,N_2844);
and UO_127 (O_127,N_2680,N_2412);
and UO_128 (O_128,N_2581,N_2973);
nand UO_129 (O_129,N_2813,N_2927);
and UO_130 (O_130,N_2563,N_2907);
nand UO_131 (O_131,N_2666,N_2785);
and UO_132 (O_132,N_2525,N_2705);
or UO_133 (O_133,N_2698,N_2487);
and UO_134 (O_134,N_2715,N_2659);
or UO_135 (O_135,N_2492,N_2712);
and UO_136 (O_136,N_2739,N_2640);
nand UO_137 (O_137,N_2702,N_2933);
nor UO_138 (O_138,N_2795,N_2978);
nor UO_139 (O_139,N_2790,N_2981);
nand UO_140 (O_140,N_2885,N_2470);
and UO_141 (O_141,N_2578,N_2996);
nor UO_142 (O_142,N_2744,N_2875);
or UO_143 (O_143,N_2762,N_2710);
and UO_144 (O_144,N_2982,N_2490);
and UO_145 (O_145,N_2402,N_2894);
nand UO_146 (O_146,N_2420,N_2846);
xnor UO_147 (O_147,N_2510,N_2992);
nor UO_148 (O_148,N_2541,N_2752);
and UO_149 (O_149,N_2759,N_2828);
nor UO_150 (O_150,N_2604,N_2720);
nand UO_151 (O_151,N_2937,N_2807);
or UO_152 (O_152,N_2930,N_2968);
or UO_153 (O_153,N_2587,N_2620);
or UO_154 (O_154,N_2924,N_2758);
xor UO_155 (O_155,N_2565,N_2606);
nor UO_156 (O_156,N_2642,N_2906);
and UO_157 (O_157,N_2418,N_2517);
and UO_158 (O_158,N_2401,N_2502);
nor UO_159 (O_159,N_2947,N_2732);
nor UO_160 (O_160,N_2904,N_2588);
nor UO_161 (O_161,N_2778,N_2882);
or UO_162 (O_162,N_2579,N_2685);
nor UO_163 (O_163,N_2872,N_2595);
nor UO_164 (O_164,N_2794,N_2889);
nand UO_165 (O_165,N_2738,N_2970);
or UO_166 (O_166,N_2766,N_2726);
or UO_167 (O_167,N_2855,N_2736);
nand UO_168 (O_168,N_2873,N_2724);
nor UO_169 (O_169,N_2887,N_2618);
nor UO_170 (O_170,N_2741,N_2551);
xnor UO_171 (O_171,N_2871,N_2539);
nor UO_172 (O_172,N_2735,N_2479);
nand UO_173 (O_173,N_2617,N_2447);
nor UO_174 (O_174,N_2524,N_2899);
or UO_175 (O_175,N_2956,N_2497);
or UO_176 (O_176,N_2769,N_2754);
nor UO_177 (O_177,N_2665,N_2874);
nor UO_178 (O_178,N_2820,N_2652);
nand UO_179 (O_179,N_2506,N_2898);
and UO_180 (O_180,N_2681,N_2729);
nor UO_181 (O_181,N_2600,N_2817);
or UO_182 (O_182,N_2877,N_2961);
or UO_183 (O_183,N_2829,N_2585);
and UO_184 (O_184,N_2679,N_2456);
nor UO_185 (O_185,N_2471,N_2713);
and UO_186 (O_186,N_2634,N_2958);
and UO_187 (O_187,N_2707,N_2669);
or UO_188 (O_188,N_2628,N_2535);
and UO_189 (O_189,N_2990,N_2857);
nand UO_190 (O_190,N_2410,N_2435);
nand UO_191 (O_191,N_2528,N_2532);
nand UO_192 (O_192,N_2725,N_2799);
or UO_193 (O_193,N_2838,N_2733);
or UO_194 (O_194,N_2674,N_2716);
and UO_195 (O_195,N_2427,N_2534);
and UO_196 (O_196,N_2521,N_2921);
and UO_197 (O_197,N_2400,N_2537);
nand UO_198 (O_198,N_2888,N_2526);
nand UO_199 (O_199,N_2441,N_2826);
and UO_200 (O_200,N_2843,N_2784);
xnor UO_201 (O_201,N_2905,N_2703);
nor UO_202 (O_202,N_2656,N_2571);
and UO_203 (O_203,N_2591,N_2789);
nor UO_204 (O_204,N_2582,N_2814);
xnor UO_205 (O_205,N_2437,N_2854);
nand UO_206 (O_206,N_2602,N_2756);
xor UO_207 (O_207,N_2851,N_2971);
and UO_208 (O_208,N_2976,N_2746);
nand UO_209 (O_209,N_2630,N_2569);
or UO_210 (O_210,N_2987,N_2580);
nor UO_211 (O_211,N_2522,N_2866);
or UO_212 (O_212,N_2407,N_2616);
and UO_213 (O_213,N_2576,N_2476);
nor UO_214 (O_214,N_2706,N_2966);
and UO_215 (O_215,N_2657,N_2841);
nor UO_216 (O_216,N_2690,N_2403);
and UO_217 (O_217,N_2619,N_2751);
or UO_218 (O_218,N_2592,N_2806);
nor UO_219 (O_219,N_2902,N_2548);
or UO_220 (O_220,N_2730,N_2472);
and UO_221 (O_221,N_2765,N_2994);
and UO_222 (O_222,N_2952,N_2834);
and UO_223 (O_223,N_2803,N_2598);
nor UO_224 (O_224,N_2473,N_2529);
or UO_225 (O_225,N_2561,N_2546);
or UO_226 (O_226,N_2694,N_2696);
nor UO_227 (O_227,N_2536,N_2495);
and UO_228 (O_228,N_2631,N_2682);
nor UO_229 (O_229,N_2577,N_2944);
xor UO_230 (O_230,N_2935,N_2593);
nor UO_231 (O_231,N_2608,N_2648);
and UO_232 (O_232,N_2589,N_2708);
xnor UO_233 (O_233,N_2928,N_2554);
or UO_234 (O_234,N_2959,N_2862);
or UO_235 (O_235,N_2508,N_2663);
and UO_236 (O_236,N_2430,N_2929);
nor UO_237 (O_237,N_2808,N_2833);
nand UO_238 (O_238,N_2544,N_2438);
nor UO_239 (O_239,N_2622,N_2638);
and UO_240 (O_240,N_2777,N_2743);
nor UO_241 (O_241,N_2923,N_2590);
nand UO_242 (O_242,N_2500,N_2670);
or UO_243 (O_243,N_2566,N_2417);
xnor UO_244 (O_244,N_2893,N_2549);
or UO_245 (O_245,N_2700,N_2649);
nand UO_246 (O_246,N_2550,N_2836);
and UO_247 (O_247,N_2761,N_2768);
or UO_248 (O_248,N_2482,N_2431);
nand UO_249 (O_249,N_2543,N_2963);
and UO_250 (O_250,N_2953,N_2637);
nand UO_251 (O_251,N_2967,N_2687);
nor UO_252 (O_252,N_2507,N_2558);
or UO_253 (O_253,N_2718,N_2847);
nand UO_254 (O_254,N_2827,N_2463);
nand UO_255 (O_255,N_2936,N_2908);
and UO_256 (O_256,N_2573,N_2728);
nor UO_257 (O_257,N_2489,N_2641);
and UO_258 (O_258,N_2914,N_2611);
nand UO_259 (O_259,N_2781,N_2457);
nand UO_260 (O_260,N_2950,N_2643);
nor UO_261 (O_261,N_2454,N_2662);
nand UO_262 (O_262,N_2612,N_2969);
and UO_263 (O_263,N_2750,N_2557);
nor UO_264 (O_264,N_2692,N_2603);
or UO_265 (O_265,N_2749,N_2428);
and UO_266 (O_266,N_2486,N_2773);
or UO_267 (O_267,N_2623,N_2624);
nand UO_268 (O_268,N_2596,N_2699);
nand UO_269 (O_269,N_2422,N_2515);
or UO_270 (O_270,N_2962,N_2926);
or UO_271 (O_271,N_2740,N_2917);
and UO_272 (O_272,N_2465,N_2484);
or UO_273 (O_273,N_2940,N_2668);
xnor UO_274 (O_274,N_2485,N_2480);
nor UO_275 (O_275,N_2461,N_2869);
nand UO_276 (O_276,N_2892,N_2763);
and UO_277 (O_277,N_2837,N_2897);
xor UO_278 (O_278,N_2559,N_2661);
and UO_279 (O_279,N_2442,N_2890);
nand UO_280 (O_280,N_2709,N_2815);
and UO_281 (O_281,N_2745,N_2646);
or UO_282 (O_282,N_2891,N_2555);
and UO_283 (O_283,N_2805,N_2860);
nand UO_284 (O_284,N_2922,N_2737);
nand UO_285 (O_285,N_2494,N_2556);
or UO_286 (O_286,N_2802,N_2514);
xnor UO_287 (O_287,N_2459,N_2920);
or UO_288 (O_288,N_2449,N_2949);
or UO_289 (O_289,N_2527,N_2689);
nand UO_290 (O_290,N_2742,N_2770);
nand UO_291 (O_291,N_2989,N_2783);
xor UO_292 (O_292,N_2673,N_2667);
nand UO_293 (O_293,N_2695,N_2453);
xnor UO_294 (O_294,N_2883,N_2491);
and UO_295 (O_295,N_2509,N_2474);
xor UO_296 (O_296,N_2613,N_2530);
nor UO_297 (O_297,N_2983,N_2636);
nand UO_298 (O_298,N_2880,N_2776);
nor UO_299 (O_299,N_2977,N_2615);
nor UO_300 (O_300,N_2933,N_2414);
nor UO_301 (O_301,N_2648,N_2639);
and UO_302 (O_302,N_2449,N_2523);
nand UO_303 (O_303,N_2445,N_2795);
xnor UO_304 (O_304,N_2812,N_2809);
and UO_305 (O_305,N_2584,N_2651);
or UO_306 (O_306,N_2740,N_2919);
nor UO_307 (O_307,N_2910,N_2400);
nor UO_308 (O_308,N_2767,N_2919);
nand UO_309 (O_309,N_2981,N_2757);
nand UO_310 (O_310,N_2876,N_2668);
nor UO_311 (O_311,N_2817,N_2435);
nor UO_312 (O_312,N_2670,N_2469);
and UO_313 (O_313,N_2467,N_2984);
nor UO_314 (O_314,N_2888,N_2741);
nor UO_315 (O_315,N_2556,N_2944);
and UO_316 (O_316,N_2798,N_2507);
or UO_317 (O_317,N_2436,N_2753);
nand UO_318 (O_318,N_2402,N_2419);
nand UO_319 (O_319,N_2514,N_2540);
or UO_320 (O_320,N_2760,N_2586);
nor UO_321 (O_321,N_2952,N_2431);
or UO_322 (O_322,N_2766,N_2806);
xnor UO_323 (O_323,N_2514,N_2742);
xnor UO_324 (O_324,N_2996,N_2981);
nor UO_325 (O_325,N_2682,N_2799);
or UO_326 (O_326,N_2624,N_2449);
nor UO_327 (O_327,N_2506,N_2997);
and UO_328 (O_328,N_2453,N_2503);
nand UO_329 (O_329,N_2633,N_2741);
nor UO_330 (O_330,N_2604,N_2691);
and UO_331 (O_331,N_2778,N_2645);
nor UO_332 (O_332,N_2672,N_2553);
or UO_333 (O_333,N_2907,N_2966);
xor UO_334 (O_334,N_2655,N_2501);
and UO_335 (O_335,N_2624,N_2609);
nand UO_336 (O_336,N_2562,N_2775);
and UO_337 (O_337,N_2427,N_2410);
and UO_338 (O_338,N_2478,N_2658);
nor UO_339 (O_339,N_2455,N_2763);
or UO_340 (O_340,N_2607,N_2483);
nor UO_341 (O_341,N_2554,N_2625);
nor UO_342 (O_342,N_2617,N_2848);
nand UO_343 (O_343,N_2966,N_2543);
or UO_344 (O_344,N_2406,N_2985);
and UO_345 (O_345,N_2771,N_2438);
nor UO_346 (O_346,N_2662,N_2647);
nor UO_347 (O_347,N_2460,N_2635);
or UO_348 (O_348,N_2851,N_2417);
nand UO_349 (O_349,N_2622,N_2774);
and UO_350 (O_350,N_2695,N_2730);
and UO_351 (O_351,N_2587,N_2799);
nand UO_352 (O_352,N_2874,N_2918);
nor UO_353 (O_353,N_2417,N_2954);
nand UO_354 (O_354,N_2767,N_2893);
and UO_355 (O_355,N_2593,N_2740);
xor UO_356 (O_356,N_2444,N_2902);
or UO_357 (O_357,N_2917,N_2702);
and UO_358 (O_358,N_2633,N_2857);
and UO_359 (O_359,N_2932,N_2463);
or UO_360 (O_360,N_2603,N_2747);
nor UO_361 (O_361,N_2434,N_2494);
nand UO_362 (O_362,N_2865,N_2603);
or UO_363 (O_363,N_2409,N_2499);
xnor UO_364 (O_364,N_2612,N_2937);
nand UO_365 (O_365,N_2805,N_2722);
nor UO_366 (O_366,N_2804,N_2663);
and UO_367 (O_367,N_2703,N_2718);
or UO_368 (O_368,N_2862,N_2725);
and UO_369 (O_369,N_2591,N_2610);
nand UO_370 (O_370,N_2915,N_2965);
or UO_371 (O_371,N_2488,N_2444);
or UO_372 (O_372,N_2842,N_2684);
and UO_373 (O_373,N_2494,N_2461);
nand UO_374 (O_374,N_2682,N_2580);
and UO_375 (O_375,N_2933,N_2620);
or UO_376 (O_376,N_2873,N_2856);
nor UO_377 (O_377,N_2645,N_2437);
and UO_378 (O_378,N_2964,N_2936);
nand UO_379 (O_379,N_2997,N_2852);
and UO_380 (O_380,N_2805,N_2627);
nand UO_381 (O_381,N_2785,N_2816);
or UO_382 (O_382,N_2991,N_2705);
nand UO_383 (O_383,N_2438,N_2750);
nand UO_384 (O_384,N_2769,N_2840);
xnor UO_385 (O_385,N_2731,N_2774);
nand UO_386 (O_386,N_2413,N_2795);
and UO_387 (O_387,N_2843,N_2468);
nor UO_388 (O_388,N_2675,N_2409);
or UO_389 (O_389,N_2422,N_2882);
nor UO_390 (O_390,N_2784,N_2626);
nor UO_391 (O_391,N_2950,N_2663);
and UO_392 (O_392,N_2822,N_2994);
or UO_393 (O_393,N_2967,N_2521);
and UO_394 (O_394,N_2687,N_2878);
or UO_395 (O_395,N_2520,N_2729);
nor UO_396 (O_396,N_2747,N_2640);
nor UO_397 (O_397,N_2564,N_2514);
nor UO_398 (O_398,N_2704,N_2630);
or UO_399 (O_399,N_2694,N_2948);
nor UO_400 (O_400,N_2795,N_2934);
and UO_401 (O_401,N_2944,N_2840);
or UO_402 (O_402,N_2481,N_2873);
nor UO_403 (O_403,N_2853,N_2991);
and UO_404 (O_404,N_2609,N_2490);
or UO_405 (O_405,N_2745,N_2451);
and UO_406 (O_406,N_2839,N_2486);
nand UO_407 (O_407,N_2767,N_2638);
nand UO_408 (O_408,N_2617,N_2699);
and UO_409 (O_409,N_2545,N_2909);
or UO_410 (O_410,N_2842,N_2763);
or UO_411 (O_411,N_2511,N_2793);
nand UO_412 (O_412,N_2400,N_2606);
nor UO_413 (O_413,N_2456,N_2818);
and UO_414 (O_414,N_2591,N_2585);
and UO_415 (O_415,N_2507,N_2474);
nor UO_416 (O_416,N_2825,N_2926);
or UO_417 (O_417,N_2923,N_2973);
and UO_418 (O_418,N_2589,N_2881);
and UO_419 (O_419,N_2619,N_2674);
and UO_420 (O_420,N_2907,N_2854);
and UO_421 (O_421,N_2631,N_2728);
or UO_422 (O_422,N_2869,N_2619);
and UO_423 (O_423,N_2725,N_2491);
nand UO_424 (O_424,N_2798,N_2474);
and UO_425 (O_425,N_2526,N_2462);
nand UO_426 (O_426,N_2452,N_2536);
or UO_427 (O_427,N_2766,N_2513);
nor UO_428 (O_428,N_2926,N_2726);
or UO_429 (O_429,N_2485,N_2938);
and UO_430 (O_430,N_2670,N_2691);
xnor UO_431 (O_431,N_2666,N_2625);
nor UO_432 (O_432,N_2913,N_2405);
nand UO_433 (O_433,N_2444,N_2809);
or UO_434 (O_434,N_2902,N_2544);
nor UO_435 (O_435,N_2796,N_2901);
and UO_436 (O_436,N_2784,N_2663);
or UO_437 (O_437,N_2928,N_2871);
nor UO_438 (O_438,N_2490,N_2986);
nand UO_439 (O_439,N_2632,N_2760);
nor UO_440 (O_440,N_2662,N_2868);
or UO_441 (O_441,N_2753,N_2562);
and UO_442 (O_442,N_2779,N_2807);
xor UO_443 (O_443,N_2750,N_2790);
xor UO_444 (O_444,N_2658,N_2878);
nand UO_445 (O_445,N_2618,N_2739);
or UO_446 (O_446,N_2904,N_2788);
nor UO_447 (O_447,N_2498,N_2915);
and UO_448 (O_448,N_2531,N_2524);
nor UO_449 (O_449,N_2589,N_2537);
nor UO_450 (O_450,N_2610,N_2558);
or UO_451 (O_451,N_2804,N_2432);
and UO_452 (O_452,N_2651,N_2789);
xnor UO_453 (O_453,N_2794,N_2542);
nor UO_454 (O_454,N_2470,N_2768);
and UO_455 (O_455,N_2826,N_2436);
and UO_456 (O_456,N_2498,N_2648);
nor UO_457 (O_457,N_2728,N_2606);
nand UO_458 (O_458,N_2605,N_2787);
nand UO_459 (O_459,N_2691,N_2490);
or UO_460 (O_460,N_2747,N_2947);
nor UO_461 (O_461,N_2401,N_2517);
and UO_462 (O_462,N_2838,N_2677);
nor UO_463 (O_463,N_2686,N_2523);
or UO_464 (O_464,N_2517,N_2801);
or UO_465 (O_465,N_2970,N_2784);
xnor UO_466 (O_466,N_2647,N_2628);
nand UO_467 (O_467,N_2764,N_2859);
xnor UO_468 (O_468,N_2734,N_2952);
or UO_469 (O_469,N_2974,N_2853);
or UO_470 (O_470,N_2503,N_2983);
or UO_471 (O_471,N_2951,N_2436);
nand UO_472 (O_472,N_2574,N_2985);
nand UO_473 (O_473,N_2688,N_2610);
and UO_474 (O_474,N_2515,N_2792);
nor UO_475 (O_475,N_2677,N_2953);
nand UO_476 (O_476,N_2750,N_2505);
or UO_477 (O_477,N_2493,N_2533);
or UO_478 (O_478,N_2580,N_2623);
nor UO_479 (O_479,N_2845,N_2402);
and UO_480 (O_480,N_2554,N_2673);
nand UO_481 (O_481,N_2930,N_2698);
xnor UO_482 (O_482,N_2754,N_2986);
nor UO_483 (O_483,N_2512,N_2878);
or UO_484 (O_484,N_2599,N_2919);
nand UO_485 (O_485,N_2624,N_2792);
xnor UO_486 (O_486,N_2733,N_2607);
or UO_487 (O_487,N_2827,N_2401);
nor UO_488 (O_488,N_2716,N_2662);
or UO_489 (O_489,N_2859,N_2745);
nor UO_490 (O_490,N_2802,N_2754);
and UO_491 (O_491,N_2686,N_2638);
nand UO_492 (O_492,N_2670,N_2697);
nor UO_493 (O_493,N_2725,N_2817);
and UO_494 (O_494,N_2935,N_2723);
nand UO_495 (O_495,N_2719,N_2444);
or UO_496 (O_496,N_2926,N_2416);
nand UO_497 (O_497,N_2895,N_2441);
or UO_498 (O_498,N_2857,N_2957);
or UO_499 (O_499,N_2631,N_2861);
endmodule