module basic_500_3000_500_40_levels_2xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_432,In_184);
and U1 (N_1,In_332,In_171);
and U2 (N_2,In_422,In_223);
nor U3 (N_3,In_448,In_489);
or U4 (N_4,In_299,In_285);
nand U5 (N_5,In_58,In_36);
nand U6 (N_6,In_338,In_486);
nand U7 (N_7,In_412,In_301);
and U8 (N_8,In_323,In_267);
and U9 (N_9,In_304,In_399);
nand U10 (N_10,In_404,In_320);
and U11 (N_11,In_449,In_270);
nand U12 (N_12,In_316,In_75);
nor U13 (N_13,In_377,In_246);
nand U14 (N_14,In_344,In_112);
or U15 (N_15,In_196,In_149);
and U16 (N_16,In_30,In_67);
or U17 (N_17,In_341,In_427);
or U18 (N_18,In_5,In_212);
and U19 (N_19,In_497,In_366);
nor U20 (N_20,In_278,In_234);
nand U21 (N_21,In_87,In_494);
and U22 (N_22,In_18,In_292);
or U23 (N_23,In_307,In_124);
or U24 (N_24,In_115,In_90);
nand U25 (N_25,In_204,In_96);
xor U26 (N_26,In_379,In_159);
or U27 (N_27,In_403,In_82);
and U28 (N_28,In_41,In_227);
nand U29 (N_29,In_26,In_105);
and U30 (N_30,In_303,In_311);
or U31 (N_31,In_51,In_418);
nand U32 (N_32,In_407,In_150);
nor U33 (N_33,In_254,In_102);
nor U34 (N_34,In_91,In_376);
or U35 (N_35,In_268,In_77);
or U36 (N_36,In_321,In_243);
and U37 (N_37,In_62,In_45);
or U38 (N_38,In_187,In_161);
or U39 (N_39,In_257,In_261);
xor U40 (N_40,In_294,In_137);
nor U41 (N_41,In_471,In_310);
or U42 (N_42,In_460,In_176);
xnor U43 (N_43,In_76,In_308);
nor U44 (N_44,In_136,In_32);
nor U45 (N_45,In_312,In_279);
and U46 (N_46,In_461,In_283);
or U47 (N_47,In_358,In_386);
xor U48 (N_48,In_140,In_35);
nor U49 (N_49,In_499,In_64);
or U50 (N_50,In_206,In_1);
or U51 (N_51,In_492,In_194);
and U52 (N_52,In_333,In_127);
nor U53 (N_53,In_493,In_38);
xnor U54 (N_54,In_49,In_47);
or U55 (N_55,In_121,In_329);
nor U56 (N_56,In_396,In_479);
nand U57 (N_57,In_177,In_167);
nor U58 (N_58,In_473,In_475);
nor U59 (N_59,In_207,In_322);
xnor U60 (N_60,In_463,In_188);
nor U61 (N_61,In_384,In_220);
or U62 (N_62,In_264,In_317);
nor U63 (N_63,In_387,In_468);
nor U64 (N_64,In_394,In_346);
xor U65 (N_65,In_242,In_391);
nand U66 (N_66,In_309,In_371);
and U67 (N_67,In_426,In_6);
nor U68 (N_68,In_318,In_440);
or U69 (N_69,In_255,In_24);
nor U70 (N_70,In_129,In_455);
or U71 (N_71,In_89,In_147);
nand U72 (N_72,In_183,In_134);
nor U73 (N_73,In_495,In_469);
nand U74 (N_74,In_2,In_116);
or U75 (N_75,N_52,N_51);
nor U76 (N_76,N_5,In_375);
xnor U77 (N_77,In_25,In_233);
and U78 (N_78,In_466,In_98);
nand U79 (N_79,In_302,N_28);
or U80 (N_80,N_68,In_385);
xnor U81 (N_81,In_122,N_14);
nor U82 (N_82,In_101,In_153);
nor U83 (N_83,In_19,N_69);
nand U84 (N_84,In_256,In_88);
and U85 (N_85,In_238,In_457);
nor U86 (N_86,In_139,In_60);
or U87 (N_87,In_478,N_24);
or U88 (N_88,In_356,In_143);
nor U89 (N_89,In_453,In_109);
nor U90 (N_90,In_218,In_405);
or U91 (N_91,In_360,In_467);
and U92 (N_92,N_35,In_289);
nor U93 (N_93,N_23,In_288);
and U94 (N_94,N_63,In_23);
nand U95 (N_95,In_342,In_353);
and U96 (N_96,In_141,In_331);
or U97 (N_97,In_222,In_200);
nor U98 (N_98,In_182,In_78);
nand U99 (N_99,In_367,In_94);
and U100 (N_100,In_100,In_65);
nor U101 (N_101,In_185,In_232);
and U102 (N_102,In_85,In_205);
or U103 (N_103,In_144,In_382);
nand U104 (N_104,In_477,In_269);
and U105 (N_105,In_228,In_113);
or U106 (N_106,In_433,In_354);
and U107 (N_107,In_66,In_413);
or U108 (N_108,N_18,In_340);
nor U109 (N_109,In_476,In_214);
and U110 (N_110,In_458,In_103);
and U111 (N_111,In_210,N_34);
and U112 (N_112,In_21,In_199);
or U113 (N_113,In_31,In_50);
and U114 (N_114,In_348,In_290);
nand U115 (N_115,In_423,In_306);
nor U116 (N_116,In_68,N_19);
or U117 (N_117,In_408,In_249);
or U118 (N_118,In_111,N_62);
nand U119 (N_119,In_281,In_383);
nor U120 (N_120,N_66,In_215);
nor U121 (N_121,In_374,In_114);
nand U122 (N_122,In_8,In_451);
and U123 (N_123,In_328,In_158);
nor U124 (N_124,N_64,In_291);
and U125 (N_125,In_247,In_424);
nor U126 (N_126,In_484,In_296);
xor U127 (N_127,In_389,In_266);
or U128 (N_128,In_434,In_166);
and U129 (N_129,In_192,N_33);
and U130 (N_130,In_273,In_93);
or U131 (N_131,In_436,In_481);
nor U132 (N_132,In_414,In_14);
and U133 (N_133,In_431,N_49);
and U134 (N_134,In_104,In_216);
or U135 (N_135,In_39,In_482);
or U136 (N_136,In_397,N_16);
nand U137 (N_137,N_4,In_450);
and U138 (N_138,In_441,In_236);
xnor U139 (N_139,In_213,In_339);
nand U140 (N_140,In_401,In_483);
nand U141 (N_141,In_496,In_271);
and U142 (N_142,In_157,In_48);
nand U143 (N_143,In_409,In_175);
nor U144 (N_144,In_178,In_119);
nor U145 (N_145,In_92,In_364);
nand U146 (N_146,In_79,In_118);
nand U147 (N_147,In_170,In_355);
or U148 (N_148,In_370,In_231);
and U149 (N_149,In_319,N_42);
nand U150 (N_150,In_277,In_42);
nand U151 (N_151,In_430,In_84);
nor U152 (N_152,N_70,N_22);
and U153 (N_153,In_343,N_100);
and U154 (N_154,In_474,In_37);
and U155 (N_155,In_52,In_203);
nor U156 (N_156,In_193,In_126);
nand U157 (N_157,In_63,In_27);
and U158 (N_158,In_437,In_16);
nand U159 (N_159,N_106,N_2);
and U160 (N_160,N_74,In_191);
or U161 (N_161,N_75,In_416);
nand U162 (N_162,In_224,In_9);
or U163 (N_163,In_46,In_337);
or U164 (N_164,In_284,In_392);
nand U165 (N_165,In_145,In_73);
and U166 (N_166,N_109,In_260);
or U167 (N_167,In_373,N_83);
and U168 (N_168,In_417,In_240);
nor U169 (N_169,In_86,N_39);
and U170 (N_170,N_141,In_445);
or U171 (N_171,In_11,In_351);
and U172 (N_172,In_132,In_447);
or U173 (N_173,In_123,In_443);
and U174 (N_174,In_108,In_160);
nand U175 (N_175,N_80,N_147);
nor U176 (N_176,In_324,N_114);
xor U177 (N_177,N_58,N_84);
nor U178 (N_178,N_40,In_305);
nor U179 (N_179,In_29,In_189);
nand U180 (N_180,N_113,In_152);
and U181 (N_181,In_146,In_287);
and U182 (N_182,N_88,In_130);
nand U183 (N_183,N_7,In_7);
nand U184 (N_184,In_237,In_363);
or U185 (N_185,In_395,In_97);
and U186 (N_186,In_250,N_65);
and U187 (N_187,N_95,In_43);
nor U188 (N_188,In_61,In_327);
and U189 (N_189,N_140,In_345);
nor U190 (N_190,In_398,In_179);
nand U191 (N_191,In_258,In_55);
nor U192 (N_192,N_47,N_132);
nand U193 (N_193,In_280,In_465);
nor U194 (N_194,N_134,In_142);
nand U195 (N_195,N_73,N_136);
nand U196 (N_196,N_72,In_487);
nand U197 (N_197,N_21,N_93);
nor U198 (N_198,In_201,In_138);
or U199 (N_199,In_282,In_125);
and U200 (N_200,In_378,N_103);
nor U201 (N_201,N_123,In_421);
nand U202 (N_202,In_22,In_117);
or U203 (N_203,In_352,In_163);
or U204 (N_204,In_173,In_252);
nand U205 (N_205,N_3,In_110);
and U206 (N_206,In_198,In_272);
nand U207 (N_207,In_357,N_57);
or U208 (N_208,N_110,N_71);
nor U209 (N_209,N_139,In_393);
or U210 (N_210,In_133,In_53);
nand U211 (N_211,In_245,N_54);
nor U212 (N_212,In_181,N_121);
nand U213 (N_213,N_56,In_359);
nand U214 (N_214,In_253,In_13);
xnor U215 (N_215,N_9,N_25);
and U216 (N_216,N_146,In_350);
nor U217 (N_217,N_130,N_119);
nor U218 (N_218,N_116,N_11);
or U219 (N_219,In_297,In_44);
nand U220 (N_220,In_128,In_54);
and U221 (N_221,N_92,N_48);
or U222 (N_222,N_138,In_248);
nor U223 (N_223,In_300,In_444);
nand U224 (N_224,In_211,In_74);
nor U225 (N_225,N_115,N_145);
nand U226 (N_226,In_335,In_10);
nor U227 (N_227,N_212,In_368);
and U228 (N_228,In_454,In_326);
or U229 (N_229,In_406,N_32);
or U230 (N_230,N_161,N_144);
and U231 (N_231,N_13,In_20);
nand U232 (N_232,In_365,N_199);
and U233 (N_233,N_158,N_108);
or U234 (N_234,N_196,N_177);
nor U235 (N_235,N_164,N_91);
or U236 (N_236,In_411,In_313);
nand U237 (N_237,N_191,N_185);
nor U238 (N_238,In_219,In_251);
or U239 (N_239,In_380,In_154);
xnor U240 (N_240,N_150,In_286);
nand U241 (N_241,N_105,In_174);
nor U242 (N_242,In_168,N_220);
or U243 (N_243,In_71,In_470);
nand U244 (N_244,N_29,In_57);
nor U245 (N_245,In_388,In_107);
and U246 (N_246,N_135,N_15);
or U247 (N_247,In_259,In_40);
nand U248 (N_248,N_218,N_112);
or U249 (N_249,N_0,In_295);
or U250 (N_250,In_464,N_200);
or U251 (N_251,In_274,N_154);
nand U252 (N_252,N_107,In_400);
nand U253 (N_253,In_59,N_176);
or U254 (N_254,N_216,N_12);
and U255 (N_255,In_472,N_149);
nand U256 (N_256,N_203,N_90);
or U257 (N_257,N_1,N_202);
nor U258 (N_258,In_131,N_160);
nand U259 (N_259,In_80,In_244);
or U260 (N_260,In_81,In_235);
nor U261 (N_261,N_143,In_263);
and U262 (N_262,In_435,In_442);
nor U263 (N_263,In_265,N_209);
and U264 (N_264,N_97,In_241);
or U265 (N_265,N_208,In_390);
nor U266 (N_266,N_156,N_194);
or U267 (N_267,In_410,N_148);
nand U268 (N_268,In_459,N_94);
nand U269 (N_269,N_222,N_152);
nand U270 (N_270,N_221,In_491);
and U271 (N_271,In_425,N_38);
nor U272 (N_272,In_456,N_162);
and U273 (N_273,N_104,N_26);
nor U274 (N_274,In_275,N_167);
nor U275 (N_275,N_120,In_229);
or U276 (N_276,In_217,N_78);
nor U277 (N_277,In_56,N_102);
nand U278 (N_278,In_197,In_72);
nand U279 (N_279,N_125,In_169);
or U280 (N_280,In_148,N_201);
or U281 (N_281,N_169,N_53);
or U282 (N_282,N_213,N_81);
xor U283 (N_283,N_10,In_402);
nand U284 (N_284,In_164,In_162);
and U285 (N_285,In_314,N_60);
or U286 (N_286,N_184,In_276);
or U287 (N_287,N_43,In_420);
nor U288 (N_288,N_86,In_325);
and U289 (N_289,N_173,N_96);
nand U290 (N_290,In_262,In_330);
or U291 (N_291,N_190,N_101);
nor U292 (N_292,N_99,N_211);
or U293 (N_293,In_439,In_135);
nor U294 (N_294,N_183,In_480);
nor U295 (N_295,N_206,N_20);
or U296 (N_296,In_485,N_224);
or U297 (N_297,N_8,N_171);
nor U298 (N_298,In_180,In_34);
nor U299 (N_299,N_46,N_67);
nor U300 (N_300,N_284,In_209);
nand U301 (N_301,N_87,In_428);
nor U302 (N_302,N_189,N_117);
nand U303 (N_303,N_41,In_438);
nand U304 (N_304,N_188,N_234);
nand U305 (N_305,N_45,N_279);
and U306 (N_306,N_27,N_270);
nand U307 (N_307,N_288,In_230);
nor U308 (N_308,N_77,N_59);
nor U309 (N_309,N_259,In_165);
or U310 (N_310,In_369,N_280);
and U311 (N_311,In_462,N_268);
or U312 (N_312,N_241,N_111);
nor U313 (N_313,N_286,N_151);
and U314 (N_314,In_12,N_292);
and U315 (N_315,In_190,N_210);
or U316 (N_316,In_15,In_446);
nand U317 (N_317,In_347,In_225);
nor U318 (N_318,N_153,N_124);
or U319 (N_319,N_170,In_156);
nand U320 (N_320,In_195,N_207);
and U321 (N_321,In_336,In_0);
nor U322 (N_322,N_30,N_267);
and U323 (N_323,N_244,N_293);
nor U324 (N_324,N_255,N_232);
or U325 (N_325,N_258,N_192);
nor U326 (N_326,N_238,N_55);
or U327 (N_327,N_6,N_251);
or U328 (N_328,N_289,In_221);
or U329 (N_329,In_120,N_245);
nand U330 (N_330,N_295,N_248);
xnor U331 (N_331,In_70,N_242);
nor U332 (N_332,N_229,In_83);
nand U333 (N_333,N_253,N_198);
nor U334 (N_334,N_276,N_256);
and U335 (N_335,N_179,N_274);
and U336 (N_336,N_296,In_498);
nand U337 (N_337,N_275,In_488);
nor U338 (N_338,N_278,N_128);
and U339 (N_339,N_277,In_349);
nor U340 (N_340,N_282,N_85);
or U341 (N_341,N_298,N_215);
nand U342 (N_342,N_193,In_372);
or U343 (N_343,N_118,In_28);
nor U344 (N_344,N_37,N_17);
xor U345 (N_345,In_172,N_166);
and U346 (N_346,In_17,N_240);
or U347 (N_347,N_172,N_236);
nand U348 (N_348,N_142,N_165);
nand U349 (N_349,N_133,N_273);
and U350 (N_350,N_246,In_362);
nor U351 (N_351,N_257,N_131);
and U352 (N_352,N_195,N_182);
nor U353 (N_353,N_227,In_69);
and U354 (N_354,N_204,N_197);
and U355 (N_355,N_219,N_82);
nor U356 (N_356,N_163,In_298);
nand U357 (N_357,N_271,N_264);
nand U358 (N_358,N_243,In_99);
or U359 (N_359,N_79,N_89);
nor U360 (N_360,In_490,N_226);
nand U361 (N_361,In_95,N_231);
or U362 (N_362,In_293,N_235);
nor U363 (N_363,N_281,N_260);
nor U364 (N_364,In_452,In_202);
nand U365 (N_365,N_237,N_178);
or U366 (N_366,N_181,In_106);
nand U367 (N_367,N_98,N_230);
xnor U368 (N_368,In_361,N_223);
or U369 (N_369,In_33,N_187);
and U370 (N_370,N_265,In_4);
or U371 (N_371,N_291,In_3);
or U372 (N_372,N_175,N_129);
and U373 (N_373,N_168,In_315);
and U374 (N_374,N_217,N_254);
or U375 (N_375,In_239,N_249);
or U376 (N_376,N_155,N_359);
and U377 (N_377,N_180,N_310);
and U378 (N_378,N_364,N_344);
nand U379 (N_379,N_318,N_357);
or U380 (N_380,N_316,N_350);
nor U381 (N_381,N_362,N_300);
nand U382 (N_382,N_322,N_269);
or U383 (N_383,N_299,N_370);
and U384 (N_384,N_363,N_31);
nor U385 (N_385,N_337,N_354);
nor U386 (N_386,N_372,N_261);
nand U387 (N_387,N_283,N_250);
or U388 (N_388,N_321,N_368);
and U389 (N_389,In_186,N_327);
nor U390 (N_390,N_214,N_61);
and U391 (N_391,N_343,N_342);
and U392 (N_392,N_285,In_415);
xor U393 (N_393,N_332,N_306);
and U394 (N_394,N_294,N_367);
nor U395 (N_395,N_247,N_349);
nand U396 (N_396,N_347,N_309);
or U397 (N_397,N_228,N_317);
nor U398 (N_398,N_186,N_334);
or U399 (N_399,N_346,N_330);
nand U400 (N_400,N_159,In_334);
nor U401 (N_401,In_208,In_151);
and U402 (N_402,N_290,N_252);
nand U403 (N_403,N_311,N_373);
or U404 (N_404,N_329,N_352);
and U405 (N_405,N_297,N_358);
or U406 (N_406,N_326,N_239);
and U407 (N_407,N_301,N_314);
nor U408 (N_408,N_225,N_127);
or U409 (N_409,N_157,N_328);
nor U410 (N_410,N_339,N_351);
or U411 (N_411,N_319,N_371);
or U412 (N_412,N_355,N_336);
and U413 (N_413,N_307,N_305);
or U414 (N_414,N_356,N_323);
nand U415 (N_415,N_340,N_174);
nor U416 (N_416,In_429,N_369);
nand U417 (N_417,N_365,N_76);
and U418 (N_418,N_308,In_155);
nand U419 (N_419,N_335,N_338);
nand U420 (N_420,N_122,N_315);
nand U421 (N_421,N_366,N_361);
or U422 (N_422,N_313,N_345);
and U423 (N_423,N_312,N_320);
or U424 (N_424,N_348,N_50);
nand U425 (N_425,N_126,In_381);
or U426 (N_426,N_287,N_205);
or U427 (N_427,N_341,N_302);
and U428 (N_428,N_304,N_360);
or U429 (N_429,N_137,N_272);
nand U430 (N_430,N_36,N_303);
nand U431 (N_431,N_262,In_419);
or U432 (N_432,N_233,N_331);
and U433 (N_433,N_374,N_263);
and U434 (N_434,N_325,N_353);
and U435 (N_435,N_333,N_266);
or U436 (N_436,N_324,In_226);
or U437 (N_437,N_44,In_381);
nand U438 (N_438,N_338,N_283);
nand U439 (N_439,N_370,N_363);
and U440 (N_440,N_340,N_329);
nor U441 (N_441,N_299,N_225);
and U442 (N_442,N_369,N_342);
or U443 (N_443,N_50,N_326);
and U444 (N_444,N_301,N_44);
nor U445 (N_445,N_345,N_363);
xor U446 (N_446,N_366,N_320);
and U447 (N_447,N_297,N_340);
nand U448 (N_448,N_339,N_355);
nor U449 (N_449,N_335,N_250);
or U450 (N_450,N_408,N_410);
or U451 (N_451,N_386,N_400);
nor U452 (N_452,N_444,N_413);
or U453 (N_453,N_375,N_426);
or U454 (N_454,N_436,N_391);
nand U455 (N_455,N_420,N_381);
or U456 (N_456,N_378,N_405);
and U457 (N_457,N_385,N_445);
nor U458 (N_458,N_407,N_382);
and U459 (N_459,N_446,N_441);
nand U460 (N_460,N_425,N_409);
and U461 (N_461,N_398,N_417);
xnor U462 (N_462,N_387,N_437);
and U463 (N_463,N_412,N_394);
nor U464 (N_464,N_428,N_411);
or U465 (N_465,N_423,N_404);
nand U466 (N_466,N_395,N_438);
nor U467 (N_467,N_442,N_402);
and U468 (N_468,N_422,N_418);
xor U469 (N_469,N_392,N_434);
or U470 (N_470,N_447,N_435);
and U471 (N_471,N_377,N_376);
nand U472 (N_472,N_432,N_419);
nor U473 (N_473,N_439,N_440);
and U474 (N_474,N_429,N_430);
nand U475 (N_475,N_390,N_388);
nor U476 (N_476,N_379,N_421);
and U477 (N_477,N_427,N_384);
nor U478 (N_478,N_397,N_416);
nor U479 (N_479,N_449,N_431);
and U480 (N_480,N_415,N_403);
or U481 (N_481,N_389,N_433);
or U482 (N_482,N_401,N_448);
or U483 (N_483,N_414,N_380);
or U484 (N_484,N_383,N_443);
nor U485 (N_485,N_406,N_399);
nor U486 (N_486,N_396,N_393);
or U487 (N_487,N_424,N_401);
nand U488 (N_488,N_398,N_443);
nand U489 (N_489,N_388,N_442);
or U490 (N_490,N_380,N_421);
nand U491 (N_491,N_403,N_380);
nor U492 (N_492,N_413,N_393);
nor U493 (N_493,N_422,N_405);
nor U494 (N_494,N_422,N_440);
nand U495 (N_495,N_392,N_417);
nand U496 (N_496,N_424,N_446);
and U497 (N_497,N_397,N_378);
or U498 (N_498,N_409,N_392);
nand U499 (N_499,N_411,N_417);
xor U500 (N_500,N_417,N_441);
and U501 (N_501,N_380,N_448);
and U502 (N_502,N_391,N_399);
and U503 (N_503,N_409,N_385);
or U504 (N_504,N_427,N_412);
nor U505 (N_505,N_424,N_386);
or U506 (N_506,N_426,N_408);
or U507 (N_507,N_385,N_379);
nand U508 (N_508,N_381,N_426);
or U509 (N_509,N_402,N_446);
nand U510 (N_510,N_443,N_396);
and U511 (N_511,N_435,N_389);
and U512 (N_512,N_426,N_396);
or U513 (N_513,N_415,N_431);
or U514 (N_514,N_377,N_427);
nand U515 (N_515,N_436,N_412);
nand U516 (N_516,N_432,N_443);
or U517 (N_517,N_434,N_427);
and U518 (N_518,N_386,N_384);
and U519 (N_519,N_439,N_428);
nor U520 (N_520,N_431,N_425);
xnor U521 (N_521,N_400,N_380);
nor U522 (N_522,N_421,N_414);
or U523 (N_523,N_387,N_399);
nor U524 (N_524,N_423,N_395);
or U525 (N_525,N_488,N_464);
nand U526 (N_526,N_520,N_504);
or U527 (N_527,N_502,N_509);
nand U528 (N_528,N_487,N_483);
or U529 (N_529,N_450,N_501);
nor U530 (N_530,N_497,N_524);
or U531 (N_531,N_470,N_452);
nor U532 (N_532,N_473,N_481);
and U533 (N_533,N_479,N_451);
and U534 (N_534,N_466,N_522);
and U535 (N_535,N_508,N_462);
or U536 (N_536,N_468,N_453);
or U537 (N_537,N_475,N_496);
or U538 (N_538,N_480,N_458);
and U539 (N_539,N_516,N_490);
and U540 (N_540,N_505,N_506);
or U541 (N_541,N_486,N_484);
nand U542 (N_542,N_519,N_495);
and U543 (N_543,N_489,N_469);
nand U544 (N_544,N_491,N_500);
or U545 (N_545,N_511,N_471);
nand U546 (N_546,N_465,N_459);
or U547 (N_547,N_513,N_474);
xnor U548 (N_548,N_478,N_517);
and U549 (N_549,N_493,N_454);
or U550 (N_550,N_460,N_463);
or U551 (N_551,N_510,N_494);
and U552 (N_552,N_467,N_455);
nand U553 (N_553,N_492,N_518);
nand U554 (N_554,N_499,N_457);
and U555 (N_555,N_507,N_461);
xor U556 (N_556,N_456,N_515);
or U557 (N_557,N_482,N_472);
xor U558 (N_558,N_476,N_521);
and U559 (N_559,N_498,N_514);
nand U560 (N_560,N_523,N_477);
and U561 (N_561,N_512,N_503);
nor U562 (N_562,N_485,N_518);
nand U563 (N_563,N_469,N_516);
nand U564 (N_564,N_473,N_483);
and U565 (N_565,N_472,N_465);
and U566 (N_566,N_466,N_477);
and U567 (N_567,N_511,N_489);
nor U568 (N_568,N_492,N_460);
nand U569 (N_569,N_511,N_475);
nand U570 (N_570,N_467,N_492);
and U571 (N_571,N_474,N_517);
nor U572 (N_572,N_484,N_503);
and U573 (N_573,N_498,N_493);
and U574 (N_574,N_480,N_461);
xor U575 (N_575,N_458,N_453);
or U576 (N_576,N_515,N_507);
nand U577 (N_577,N_466,N_490);
nand U578 (N_578,N_475,N_498);
or U579 (N_579,N_479,N_506);
or U580 (N_580,N_463,N_489);
or U581 (N_581,N_459,N_510);
xnor U582 (N_582,N_491,N_484);
and U583 (N_583,N_500,N_464);
or U584 (N_584,N_456,N_468);
or U585 (N_585,N_463,N_478);
nand U586 (N_586,N_514,N_457);
nor U587 (N_587,N_521,N_460);
or U588 (N_588,N_478,N_458);
and U589 (N_589,N_457,N_477);
nand U590 (N_590,N_483,N_516);
nor U591 (N_591,N_458,N_505);
or U592 (N_592,N_524,N_472);
nand U593 (N_593,N_491,N_488);
and U594 (N_594,N_518,N_451);
or U595 (N_595,N_479,N_487);
nand U596 (N_596,N_482,N_477);
or U597 (N_597,N_516,N_515);
or U598 (N_598,N_510,N_468);
nor U599 (N_599,N_501,N_490);
nand U600 (N_600,N_557,N_576);
and U601 (N_601,N_541,N_554);
and U602 (N_602,N_568,N_569);
nand U603 (N_603,N_527,N_532);
nand U604 (N_604,N_563,N_595);
or U605 (N_605,N_581,N_533);
and U606 (N_606,N_579,N_571);
nor U607 (N_607,N_592,N_584);
and U608 (N_608,N_546,N_551);
or U609 (N_609,N_582,N_588);
nor U610 (N_610,N_570,N_531);
and U611 (N_611,N_564,N_580);
nand U612 (N_612,N_573,N_578);
nand U613 (N_613,N_548,N_577);
or U614 (N_614,N_590,N_542);
or U615 (N_615,N_550,N_583);
nand U616 (N_616,N_585,N_526);
nand U617 (N_617,N_549,N_566);
and U618 (N_618,N_556,N_597);
or U619 (N_619,N_591,N_540);
and U620 (N_620,N_598,N_565);
and U621 (N_621,N_562,N_536);
nand U622 (N_622,N_594,N_529);
nand U623 (N_623,N_530,N_534);
nand U624 (N_624,N_543,N_547);
and U625 (N_625,N_538,N_539);
or U626 (N_626,N_593,N_589);
nand U627 (N_627,N_596,N_599);
and U628 (N_628,N_586,N_587);
nor U629 (N_629,N_528,N_558);
and U630 (N_630,N_572,N_559);
xor U631 (N_631,N_545,N_555);
nand U632 (N_632,N_552,N_535);
nand U633 (N_633,N_525,N_575);
nand U634 (N_634,N_567,N_561);
nor U635 (N_635,N_553,N_537);
nor U636 (N_636,N_544,N_560);
and U637 (N_637,N_574,N_549);
and U638 (N_638,N_577,N_571);
or U639 (N_639,N_581,N_567);
and U640 (N_640,N_583,N_560);
nand U641 (N_641,N_546,N_557);
nand U642 (N_642,N_598,N_530);
nand U643 (N_643,N_541,N_586);
or U644 (N_644,N_575,N_542);
nor U645 (N_645,N_569,N_599);
or U646 (N_646,N_595,N_585);
nand U647 (N_647,N_570,N_592);
nand U648 (N_648,N_535,N_529);
nor U649 (N_649,N_575,N_541);
nor U650 (N_650,N_546,N_552);
or U651 (N_651,N_534,N_583);
nand U652 (N_652,N_559,N_575);
nor U653 (N_653,N_547,N_577);
nand U654 (N_654,N_528,N_579);
and U655 (N_655,N_564,N_525);
or U656 (N_656,N_578,N_544);
nand U657 (N_657,N_546,N_573);
or U658 (N_658,N_544,N_597);
nand U659 (N_659,N_544,N_576);
or U660 (N_660,N_581,N_566);
nor U661 (N_661,N_541,N_534);
or U662 (N_662,N_537,N_547);
nand U663 (N_663,N_578,N_579);
nand U664 (N_664,N_553,N_541);
nand U665 (N_665,N_534,N_557);
or U666 (N_666,N_543,N_525);
or U667 (N_667,N_526,N_527);
nor U668 (N_668,N_535,N_599);
xnor U669 (N_669,N_548,N_565);
and U670 (N_670,N_530,N_570);
xor U671 (N_671,N_561,N_543);
and U672 (N_672,N_561,N_550);
or U673 (N_673,N_590,N_551);
nand U674 (N_674,N_585,N_587);
nor U675 (N_675,N_633,N_617);
nor U676 (N_676,N_613,N_649);
or U677 (N_677,N_627,N_652);
or U678 (N_678,N_616,N_628);
and U679 (N_679,N_644,N_664);
nand U680 (N_680,N_630,N_665);
and U681 (N_681,N_629,N_648);
and U682 (N_682,N_622,N_673);
nand U683 (N_683,N_635,N_646);
or U684 (N_684,N_640,N_604);
nor U685 (N_685,N_618,N_638);
nor U686 (N_686,N_600,N_668);
nor U687 (N_687,N_657,N_631);
or U688 (N_688,N_653,N_607);
and U689 (N_689,N_660,N_658);
or U690 (N_690,N_670,N_669);
xnor U691 (N_691,N_634,N_656);
nand U692 (N_692,N_636,N_610);
nor U693 (N_693,N_615,N_672);
nand U694 (N_694,N_623,N_614);
and U695 (N_695,N_632,N_608);
or U696 (N_696,N_671,N_663);
nand U697 (N_697,N_621,N_654);
nand U698 (N_698,N_612,N_603);
xnor U699 (N_699,N_661,N_650);
nor U700 (N_700,N_666,N_620);
nor U701 (N_701,N_619,N_647);
or U702 (N_702,N_625,N_662);
nor U703 (N_703,N_605,N_626);
and U704 (N_704,N_601,N_655);
nor U705 (N_705,N_602,N_642);
nor U706 (N_706,N_659,N_606);
nor U707 (N_707,N_641,N_624);
nand U708 (N_708,N_643,N_674);
xnor U709 (N_709,N_645,N_637);
or U710 (N_710,N_639,N_611);
nand U711 (N_711,N_651,N_667);
nand U712 (N_712,N_609,N_671);
or U713 (N_713,N_630,N_612);
nand U714 (N_714,N_605,N_608);
or U715 (N_715,N_639,N_672);
and U716 (N_716,N_600,N_615);
and U717 (N_717,N_624,N_610);
and U718 (N_718,N_673,N_610);
and U719 (N_719,N_613,N_634);
or U720 (N_720,N_663,N_646);
nand U721 (N_721,N_619,N_663);
and U722 (N_722,N_668,N_667);
or U723 (N_723,N_612,N_653);
and U724 (N_724,N_670,N_625);
or U725 (N_725,N_618,N_651);
nor U726 (N_726,N_656,N_606);
nor U727 (N_727,N_640,N_629);
or U728 (N_728,N_633,N_613);
or U729 (N_729,N_624,N_670);
nor U730 (N_730,N_625,N_617);
and U731 (N_731,N_662,N_655);
nand U732 (N_732,N_647,N_664);
nand U733 (N_733,N_634,N_660);
nand U734 (N_734,N_639,N_646);
or U735 (N_735,N_635,N_655);
and U736 (N_736,N_665,N_622);
nand U737 (N_737,N_634,N_600);
and U738 (N_738,N_635,N_619);
nor U739 (N_739,N_638,N_620);
nor U740 (N_740,N_658,N_665);
nand U741 (N_741,N_650,N_642);
or U742 (N_742,N_640,N_608);
nor U743 (N_743,N_656,N_619);
and U744 (N_744,N_624,N_613);
xnor U745 (N_745,N_630,N_660);
and U746 (N_746,N_634,N_605);
or U747 (N_747,N_663,N_651);
nor U748 (N_748,N_600,N_638);
and U749 (N_749,N_630,N_602);
or U750 (N_750,N_695,N_693);
nor U751 (N_751,N_744,N_720);
nand U752 (N_752,N_742,N_694);
nor U753 (N_753,N_710,N_690);
or U754 (N_754,N_743,N_686);
or U755 (N_755,N_735,N_675);
and U756 (N_756,N_699,N_746);
and U757 (N_757,N_703,N_723);
nand U758 (N_758,N_677,N_713);
and U759 (N_759,N_700,N_680);
and U760 (N_760,N_738,N_717);
nand U761 (N_761,N_701,N_682);
or U762 (N_762,N_712,N_729);
and U763 (N_763,N_702,N_739);
or U764 (N_764,N_692,N_696);
xor U765 (N_765,N_725,N_741);
nor U766 (N_766,N_711,N_747);
nor U767 (N_767,N_709,N_683);
or U768 (N_768,N_724,N_687);
and U769 (N_769,N_726,N_740);
xnor U770 (N_770,N_721,N_748);
nor U771 (N_771,N_707,N_722);
nand U772 (N_772,N_678,N_714);
nor U773 (N_773,N_736,N_731);
or U774 (N_774,N_728,N_691);
and U775 (N_775,N_733,N_681);
nor U776 (N_776,N_715,N_734);
nand U777 (N_777,N_719,N_718);
or U778 (N_778,N_689,N_745);
xnor U779 (N_779,N_737,N_749);
or U780 (N_780,N_676,N_727);
and U781 (N_781,N_679,N_697);
nor U782 (N_782,N_708,N_688);
and U783 (N_783,N_704,N_684);
nand U784 (N_784,N_730,N_706);
nand U785 (N_785,N_732,N_705);
nand U786 (N_786,N_716,N_698);
and U787 (N_787,N_685,N_714);
nor U788 (N_788,N_702,N_711);
or U789 (N_789,N_699,N_733);
xnor U790 (N_790,N_721,N_689);
nand U791 (N_791,N_748,N_691);
or U792 (N_792,N_741,N_731);
nand U793 (N_793,N_742,N_702);
and U794 (N_794,N_693,N_707);
nor U795 (N_795,N_719,N_747);
and U796 (N_796,N_700,N_748);
nand U797 (N_797,N_724,N_725);
or U798 (N_798,N_697,N_694);
nand U799 (N_799,N_680,N_722);
or U800 (N_800,N_729,N_717);
and U801 (N_801,N_726,N_702);
nor U802 (N_802,N_706,N_712);
nor U803 (N_803,N_686,N_726);
nor U804 (N_804,N_712,N_741);
nand U805 (N_805,N_704,N_743);
nand U806 (N_806,N_703,N_683);
nor U807 (N_807,N_747,N_741);
nand U808 (N_808,N_681,N_687);
and U809 (N_809,N_700,N_710);
nand U810 (N_810,N_707,N_709);
nand U811 (N_811,N_679,N_689);
nand U812 (N_812,N_703,N_749);
or U813 (N_813,N_681,N_720);
nor U814 (N_814,N_676,N_686);
nor U815 (N_815,N_733,N_698);
and U816 (N_816,N_745,N_743);
or U817 (N_817,N_732,N_684);
nor U818 (N_818,N_698,N_721);
nand U819 (N_819,N_701,N_745);
or U820 (N_820,N_690,N_743);
nand U821 (N_821,N_698,N_730);
and U822 (N_822,N_730,N_748);
nand U823 (N_823,N_698,N_731);
and U824 (N_824,N_704,N_738);
or U825 (N_825,N_819,N_811);
or U826 (N_826,N_756,N_781);
nor U827 (N_827,N_752,N_798);
nand U828 (N_828,N_772,N_802);
nor U829 (N_829,N_821,N_779);
or U830 (N_830,N_786,N_790);
and U831 (N_831,N_767,N_784);
and U832 (N_832,N_796,N_783);
nand U833 (N_833,N_778,N_788);
nor U834 (N_834,N_758,N_753);
and U835 (N_835,N_801,N_813);
and U836 (N_836,N_824,N_780);
xnor U837 (N_837,N_766,N_805);
or U838 (N_838,N_791,N_760);
nor U839 (N_839,N_792,N_774);
nand U840 (N_840,N_750,N_800);
or U841 (N_841,N_794,N_757);
nor U842 (N_842,N_782,N_770);
nand U843 (N_843,N_806,N_817);
or U844 (N_844,N_759,N_765);
and U845 (N_845,N_804,N_814);
nand U846 (N_846,N_815,N_769);
and U847 (N_847,N_762,N_816);
or U848 (N_848,N_787,N_799);
or U849 (N_849,N_808,N_754);
and U850 (N_850,N_755,N_785);
nor U851 (N_851,N_803,N_773);
nor U852 (N_852,N_809,N_775);
nand U853 (N_853,N_812,N_768);
or U854 (N_854,N_797,N_795);
or U855 (N_855,N_807,N_810);
and U856 (N_856,N_789,N_823);
and U857 (N_857,N_761,N_764);
nand U858 (N_858,N_822,N_751);
nor U859 (N_859,N_793,N_777);
nand U860 (N_860,N_771,N_820);
nor U861 (N_861,N_763,N_818);
nand U862 (N_862,N_776,N_788);
and U863 (N_863,N_756,N_760);
nand U864 (N_864,N_763,N_815);
and U865 (N_865,N_813,N_804);
nand U866 (N_866,N_787,N_812);
nor U867 (N_867,N_824,N_794);
or U868 (N_868,N_811,N_804);
nand U869 (N_869,N_795,N_762);
nor U870 (N_870,N_815,N_800);
nor U871 (N_871,N_822,N_791);
nor U872 (N_872,N_753,N_793);
and U873 (N_873,N_762,N_820);
nor U874 (N_874,N_799,N_776);
or U875 (N_875,N_822,N_806);
or U876 (N_876,N_822,N_767);
nand U877 (N_877,N_761,N_766);
and U878 (N_878,N_780,N_785);
xnor U879 (N_879,N_780,N_776);
or U880 (N_880,N_813,N_760);
or U881 (N_881,N_765,N_772);
or U882 (N_882,N_795,N_788);
xor U883 (N_883,N_806,N_810);
nor U884 (N_884,N_791,N_797);
and U885 (N_885,N_812,N_753);
nand U886 (N_886,N_776,N_789);
or U887 (N_887,N_814,N_802);
or U888 (N_888,N_769,N_776);
nor U889 (N_889,N_761,N_788);
or U890 (N_890,N_824,N_769);
or U891 (N_891,N_762,N_798);
and U892 (N_892,N_779,N_754);
and U893 (N_893,N_820,N_763);
and U894 (N_894,N_785,N_805);
nor U895 (N_895,N_767,N_781);
nand U896 (N_896,N_811,N_767);
nand U897 (N_897,N_814,N_769);
and U898 (N_898,N_773,N_770);
and U899 (N_899,N_810,N_781);
or U900 (N_900,N_866,N_884);
nand U901 (N_901,N_838,N_868);
nor U902 (N_902,N_897,N_849);
nand U903 (N_903,N_886,N_891);
nor U904 (N_904,N_887,N_894);
and U905 (N_905,N_834,N_844);
nand U906 (N_906,N_839,N_864);
nor U907 (N_907,N_898,N_880);
and U908 (N_908,N_846,N_851);
and U909 (N_909,N_870,N_895);
nor U910 (N_910,N_859,N_873);
or U911 (N_911,N_865,N_833);
nor U912 (N_912,N_830,N_863);
nor U913 (N_913,N_843,N_856);
and U914 (N_914,N_829,N_871);
or U915 (N_915,N_862,N_879);
and U916 (N_916,N_867,N_882);
or U917 (N_917,N_848,N_857);
and U918 (N_918,N_854,N_853);
nor U919 (N_919,N_828,N_826);
nor U920 (N_920,N_861,N_872);
or U921 (N_921,N_878,N_835);
or U922 (N_922,N_836,N_881);
nand U923 (N_923,N_825,N_883);
nand U924 (N_924,N_876,N_832);
and U925 (N_925,N_899,N_841);
nand U926 (N_926,N_875,N_837);
and U927 (N_927,N_869,N_845);
or U928 (N_928,N_892,N_827);
xor U929 (N_929,N_896,N_860);
nand U930 (N_930,N_890,N_888);
and U931 (N_931,N_885,N_874);
or U932 (N_932,N_850,N_847);
nand U933 (N_933,N_889,N_858);
nand U934 (N_934,N_893,N_840);
and U935 (N_935,N_852,N_831);
nand U936 (N_936,N_855,N_842);
nand U937 (N_937,N_877,N_860);
nor U938 (N_938,N_880,N_843);
nand U939 (N_939,N_832,N_894);
and U940 (N_940,N_845,N_862);
nor U941 (N_941,N_898,N_890);
nand U942 (N_942,N_866,N_875);
and U943 (N_943,N_884,N_872);
and U944 (N_944,N_857,N_877);
nand U945 (N_945,N_848,N_825);
nand U946 (N_946,N_897,N_881);
nand U947 (N_947,N_848,N_859);
or U948 (N_948,N_851,N_856);
nand U949 (N_949,N_889,N_864);
and U950 (N_950,N_871,N_893);
nand U951 (N_951,N_855,N_886);
and U952 (N_952,N_880,N_834);
nor U953 (N_953,N_880,N_846);
or U954 (N_954,N_865,N_887);
nand U955 (N_955,N_834,N_898);
and U956 (N_956,N_842,N_838);
and U957 (N_957,N_894,N_848);
nand U958 (N_958,N_839,N_854);
nand U959 (N_959,N_856,N_868);
and U960 (N_960,N_874,N_852);
and U961 (N_961,N_868,N_887);
nand U962 (N_962,N_891,N_853);
or U963 (N_963,N_834,N_825);
or U964 (N_964,N_882,N_889);
or U965 (N_965,N_893,N_833);
nand U966 (N_966,N_867,N_861);
nand U967 (N_967,N_880,N_895);
and U968 (N_968,N_857,N_846);
nand U969 (N_969,N_845,N_898);
nand U970 (N_970,N_887,N_856);
or U971 (N_971,N_836,N_880);
nor U972 (N_972,N_875,N_867);
and U973 (N_973,N_857,N_854);
nor U974 (N_974,N_845,N_853);
and U975 (N_975,N_924,N_914);
or U976 (N_976,N_936,N_913);
or U977 (N_977,N_963,N_912);
and U978 (N_978,N_955,N_922);
or U979 (N_979,N_948,N_958);
and U980 (N_980,N_947,N_954);
and U981 (N_981,N_900,N_965);
nor U982 (N_982,N_961,N_923);
and U983 (N_983,N_919,N_939);
or U984 (N_984,N_915,N_974);
nor U985 (N_985,N_926,N_966);
and U986 (N_986,N_973,N_917);
or U987 (N_987,N_918,N_945);
and U988 (N_988,N_959,N_970);
nand U989 (N_989,N_967,N_907);
nor U990 (N_990,N_949,N_908);
or U991 (N_991,N_904,N_943);
nor U992 (N_992,N_933,N_931);
xnor U993 (N_993,N_957,N_901);
nor U994 (N_994,N_968,N_929);
or U995 (N_995,N_964,N_944);
nor U996 (N_996,N_911,N_934);
nand U997 (N_997,N_906,N_941);
xor U998 (N_998,N_972,N_909);
nor U999 (N_999,N_950,N_940);
or U1000 (N_1000,N_946,N_910);
and U1001 (N_1001,N_916,N_937);
nand U1002 (N_1002,N_942,N_925);
or U1003 (N_1003,N_903,N_938);
nor U1004 (N_1004,N_962,N_952);
and U1005 (N_1005,N_953,N_935);
nor U1006 (N_1006,N_905,N_902);
and U1007 (N_1007,N_930,N_928);
and U1008 (N_1008,N_956,N_969);
and U1009 (N_1009,N_951,N_932);
or U1010 (N_1010,N_927,N_971);
and U1011 (N_1011,N_920,N_921);
nor U1012 (N_1012,N_960,N_940);
or U1013 (N_1013,N_913,N_920);
nor U1014 (N_1014,N_924,N_931);
nor U1015 (N_1015,N_915,N_930);
or U1016 (N_1016,N_935,N_922);
or U1017 (N_1017,N_914,N_944);
and U1018 (N_1018,N_943,N_907);
nor U1019 (N_1019,N_972,N_948);
or U1020 (N_1020,N_914,N_960);
or U1021 (N_1021,N_962,N_972);
or U1022 (N_1022,N_916,N_926);
nor U1023 (N_1023,N_969,N_917);
and U1024 (N_1024,N_941,N_949);
nand U1025 (N_1025,N_912,N_941);
or U1026 (N_1026,N_969,N_934);
nand U1027 (N_1027,N_915,N_955);
and U1028 (N_1028,N_933,N_941);
nand U1029 (N_1029,N_917,N_930);
and U1030 (N_1030,N_969,N_923);
nand U1031 (N_1031,N_945,N_917);
nand U1032 (N_1032,N_954,N_904);
and U1033 (N_1033,N_970,N_946);
or U1034 (N_1034,N_961,N_966);
nand U1035 (N_1035,N_927,N_953);
or U1036 (N_1036,N_944,N_974);
nor U1037 (N_1037,N_956,N_931);
and U1038 (N_1038,N_930,N_911);
or U1039 (N_1039,N_949,N_923);
or U1040 (N_1040,N_942,N_945);
nor U1041 (N_1041,N_923,N_926);
and U1042 (N_1042,N_952,N_917);
nand U1043 (N_1043,N_932,N_935);
or U1044 (N_1044,N_911,N_903);
nor U1045 (N_1045,N_930,N_913);
nand U1046 (N_1046,N_963,N_925);
or U1047 (N_1047,N_906,N_972);
and U1048 (N_1048,N_952,N_915);
nor U1049 (N_1049,N_912,N_944);
or U1050 (N_1050,N_1023,N_1040);
or U1051 (N_1051,N_979,N_1041);
or U1052 (N_1052,N_995,N_1019);
or U1053 (N_1053,N_1035,N_1020);
or U1054 (N_1054,N_984,N_1031);
or U1055 (N_1055,N_1012,N_994);
or U1056 (N_1056,N_1032,N_999);
and U1057 (N_1057,N_987,N_989);
or U1058 (N_1058,N_1021,N_1014);
nor U1059 (N_1059,N_1022,N_1026);
nor U1060 (N_1060,N_1009,N_980);
nand U1061 (N_1061,N_991,N_1001);
and U1062 (N_1062,N_1010,N_1049);
or U1063 (N_1063,N_1013,N_1045);
or U1064 (N_1064,N_1029,N_1042);
nand U1065 (N_1065,N_1018,N_1024);
or U1066 (N_1066,N_981,N_1033);
nand U1067 (N_1067,N_992,N_1030);
nand U1068 (N_1068,N_1006,N_985);
nand U1069 (N_1069,N_1043,N_978);
nand U1070 (N_1070,N_1039,N_996);
or U1071 (N_1071,N_976,N_1004);
nor U1072 (N_1072,N_990,N_1011);
nor U1073 (N_1073,N_1047,N_986);
and U1074 (N_1074,N_975,N_982);
and U1075 (N_1075,N_1015,N_1036);
nor U1076 (N_1076,N_1037,N_997);
or U1077 (N_1077,N_1000,N_1028);
nor U1078 (N_1078,N_1002,N_1038);
nor U1079 (N_1079,N_1048,N_977);
nor U1080 (N_1080,N_1016,N_1007);
or U1081 (N_1081,N_1027,N_1046);
and U1082 (N_1082,N_1003,N_1005);
or U1083 (N_1083,N_983,N_988);
nor U1084 (N_1084,N_1008,N_1025);
nand U1085 (N_1085,N_998,N_1034);
and U1086 (N_1086,N_1044,N_993);
nor U1087 (N_1087,N_1017,N_981);
nand U1088 (N_1088,N_1016,N_1049);
and U1089 (N_1089,N_1028,N_1006);
or U1090 (N_1090,N_1040,N_1017);
nor U1091 (N_1091,N_1007,N_989);
or U1092 (N_1092,N_991,N_1011);
and U1093 (N_1093,N_1038,N_1040);
and U1094 (N_1094,N_1004,N_1015);
nor U1095 (N_1095,N_995,N_1046);
nor U1096 (N_1096,N_995,N_984);
nor U1097 (N_1097,N_992,N_1009);
and U1098 (N_1098,N_1012,N_1043);
nor U1099 (N_1099,N_984,N_1024);
nor U1100 (N_1100,N_988,N_1045);
nor U1101 (N_1101,N_1014,N_985);
or U1102 (N_1102,N_997,N_999);
or U1103 (N_1103,N_983,N_987);
nor U1104 (N_1104,N_1034,N_1035);
or U1105 (N_1105,N_989,N_1033);
nor U1106 (N_1106,N_1033,N_1036);
or U1107 (N_1107,N_1042,N_975);
nand U1108 (N_1108,N_985,N_1037);
nor U1109 (N_1109,N_1044,N_1017);
nor U1110 (N_1110,N_994,N_979);
nor U1111 (N_1111,N_1023,N_1019);
nand U1112 (N_1112,N_988,N_1046);
and U1113 (N_1113,N_1016,N_1035);
and U1114 (N_1114,N_1038,N_1014);
and U1115 (N_1115,N_1015,N_999);
nand U1116 (N_1116,N_989,N_1009);
or U1117 (N_1117,N_1048,N_992);
and U1118 (N_1118,N_1003,N_1012);
nor U1119 (N_1119,N_984,N_1009);
and U1120 (N_1120,N_1015,N_1047);
nand U1121 (N_1121,N_1036,N_1038);
nor U1122 (N_1122,N_992,N_980);
or U1123 (N_1123,N_989,N_1025);
nor U1124 (N_1124,N_983,N_1005);
and U1125 (N_1125,N_1088,N_1094);
and U1126 (N_1126,N_1110,N_1101);
nor U1127 (N_1127,N_1123,N_1120);
xor U1128 (N_1128,N_1121,N_1077);
nand U1129 (N_1129,N_1070,N_1107);
and U1130 (N_1130,N_1059,N_1063);
or U1131 (N_1131,N_1092,N_1052);
xnor U1132 (N_1132,N_1062,N_1082);
or U1133 (N_1133,N_1119,N_1074);
and U1134 (N_1134,N_1080,N_1087);
nor U1135 (N_1135,N_1068,N_1061);
nand U1136 (N_1136,N_1086,N_1089);
and U1137 (N_1137,N_1111,N_1085);
and U1138 (N_1138,N_1072,N_1060);
nand U1139 (N_1139,N_1096,N_1109);
nand U1140 (N_1140,N_1122,N_1073);
or U1141 (N_1141,N_1117,N_1075);
or U1142 (N_1142,N_1076,N_1053);
nor U1143 (N_1143,N_1055,N_1114);
nand U1144 (N_1144,N_1100,N_1115);
nand U1145 (N_1145,N_1103,N_1084);
or U1146 (N_1146,N_1054,N_1124);
and U1147 (N_1147,N_1065,N_1081);
or U1148 (N_1148,N_1057,N_1078);
or U1149 (N_1149,N_1051,N_1099);
or U1150 (N_1150,N_1050,N_1066);
nor U1151 (N_1151,N_1058,N_1093);
nand U1152 (N_1152,N_1102,N_1106);
and U1153 (N_1153,N_1091,N_1097);
and U1154 (N_1154,N_1067,N_1104);
nor U1155 (N_1155,N_1098,N_1113);
nor U1156 (N_1156,N_1064,N_1116);
nor U1157 (N_1157,N_1108,N_1112);
nor U1158 (N_1158,N_1118,N_1083);
nor U1159 (N_1159,N_1095,N_1079);
and U1160 (N_1160,N_1069,N_1090);
nand U1161 (N_1161,N_1105,N_1056);
or U1162 (N_1162,N_1071,N_1097);
and U1163 (N_1163,N_1103,N_1051);
and U1164 (N_1164,N_1076,N_1090);
and U1165 (N_1165,N_1121,N_1062);
nand U1166 (N_1166,N_1094,N_1072);
nand U1167 (N_1167,N_1107,N_1123);
nand U1168 (N_1168,N_1060,N_1116);
xnor U1169 (N_1169,N_1091,N_1089);
or U1170 (N_1170,N_1110,N_1094);
nand U1171 (N_1171,N_1117,N_1097);
and U1172 (N_1172,N_1066,N_1057);
nor U1173 (N_1173,N_1056,N_1109);
nor U1174 (N_1174,N_1086,N_1054);
or U1175 (N_1175,N_1103,N_1100);
or U1176 (N_1176,N_1114,N_1074);
or U1177 (N_1177,N_1107,N_1109);
nand U1178 (N_1178,N_1075,N_1121);
nor U1179 (N_1179,N_1078,N_1089);
and U1180 (N_1180,N_1097,N_1123);
or U1181 (N_1181,N_1121,N_1082);
nand U1182 (N_1182,N_1080,N_1091);
or U1183 (N_1183,N_1060,N_1066);
and U1184 (N_1184,N_1118,N_1107);
nand U1185 (N_1185,N_1107,N_1071);
and U1186 (N_1186,N_1059,N_1055);
nor U1187 (N_1187,N_1095,N_1121);
and U1188 (N_1188,N_1121,N_1055);
nand U1189 (N_1189,N_1060,N_1102);
nand U1190 (N_1190,N_1122,N_1068);
nand U1191 (N_1191,N_1053,N_1118);
and U1192 (N_1192,N_1123,N_1082);
or U1193 (N_1193,N_1078,N_1124);
xnor U1194 (N_1194,N_1103,N_1087);
or U1195 (N_1195,N_1075,N_1082);
nor U1196 (N_1196,N_1100,N_1058);
and U1197 (N_1197,N_1077,N_1124);
nor U1198 (N_1198,N_1115,N_1121);
nand U1199 (N_1199,N_1111,N_1061);
nand U1200 (N_1200,N_1198,N_1162);
xor U1201 (N_1201,N_1199,N_1188);
nor U1202 (N_1202,N_1158,N_1166);
nor U1203 (N_1203,N_1196,N_1126);
nor U1204 (N_1204,N_1159,N_1137);
xnor U1205 (N_1205,N_1174,N_1152);
nand U1206 (N_1206,N_1157,N_1147);
or U1207 (N_1207,N_1142,N_1143);
nor U1208 (N_1208,N_1192,N_1131);
nor U1209 (N_1209,N_1184,N_1177);
nor U1210 (N_1210,N_1130,N_1150);
nor U1211 (N_1211,N_1133,N_1181);
nor U1212 (N_1212,N_1136,N_1194);
nor U1213 (N_1213,N_1175,N_1151);
or U1214 (N_1214,N_1179,N_1160);
and U1215 (N_1215,N_1197,N_1168);
nand U1216 (N_1216,N_1189,N_1193);
and U1217 (N_1217,N_1171,N_1139);
or U1218 (N_1218,N_1190,N_1167);
and U1219 (N_1219,N_1173,N_1140);
and U1220 (N_1220,N_1172,N_1180);
and U1221 (N_1221,N_1170,N_1187);
nor U1222 (N_1222,N_1145,N_1148);
and U1223 (N_1223,N_1154,N_1178);
and U1224 (N_1224,N_1129,N_1169);
nor U1225 (N_1225,N_1191,N_1163);
nor U1226 (N_1226,N_1165,N_1141);
and U1227 (N_1227,N_1144,N_1183);
nand U1228 (N_1228,N_1176,N_1146);
or U1229 (N_1229,N_1185,N_1132);
and U1230 (N_1230,N_1164,N_1155);
nand U1231 (N_1231,N_1125,N_1128);
nand U1232 (N_1232,N_1135,N_1153);
nand U1233 (N_1233,N_1195,N_1156);
or U1234 (N_1234,N_1127,N_1134);
nand U1235 (N_1235,N_1182,N_1186);
nor U1236 (N_1236,N_1161,N_1149);
and U1237 (N_1237,N_1138,N_1170);
and U1238 (N_1238,N_1162,N_1134);
and U1239 (N_1239,N_1185,N_1187);
or U1240 (N_1240,N_1196,N_1185);
or U1241 (N_1241,N_1156,N_1140);
nor U1242 (N_1242,N_1126,N_1165);
nand U1243 (N_1243,N_1166,N_1134);
nor U1244 (N_1244,N_1159,N_1128);
and U1245 (N_1245,N_1149,N_1136);
and U1246 (N_1246,N_1148,N_1161);
or U1247 (N_1247,N_1154,N_1126);
or U1248 (N_1248,N_1156,N_1171);
nand U1249 (N_1249,N_1165,N_1189);
nor U1250 (N_1250,N_1184,N_1194);
nor U1251 (N_1251,N_1146,N_1133);
nor U1252 (N_1252,N_1130,N_1195);
and U1253 (N_1253,N_1157,N_1166);
nor U1254 (N_1254,N_1126,N_1146);
or U1255 (N_1255,N_1160,N_1168);
and U1256 (N_1256,N_1141,N_1136);
nand U1257 (N_1257,N_1183,N_1125);
nand U1258 (N_1258,N_1192,N_1135);
and U1259 (N_1259,N_1159,N_1182);
nor U1260 (N_1260,N_1164,N_1190);
and U1261 (N_1261,N_1143,N_1146);
xnor U1262 (N_1262,N_1185,N_1173);
or U1263 (N_1263,N_1199,N_1129);
nand U1264 (N_1264,N_1155,N_1185);
and U1265 (N_1265,N_1127,N_1135);
or U1266 (N_1266,N_1183,N_1178);
or U1267 (N_1267,N_1132,N_1175);
and U1268 (N_1268,N_1191,N_1185);
nor U1269 (N_1269,N_1155,N_1188);
and U1270 (N_1270,N_1152,N_1166);
and U1271 (N_1271,N_1165,N_1133);
or U1272 (N_1272,N_1167,N_1157);
or U1273 (N_1273,N_1164,N_1196);
and U1274 (N_1274,N_1191,N_1142);
nor U1275 (N_1275,N_1246,N_1213);
xnor U1276 (N_1276,N_1218,N_1222);
nand U1277 (N_1277,N_1220,N_1201);
nand U1278 (N_1278,N_1252,N_1257);
nand U1279 (N_1279,N_1219,N_1249);
or U1280 (N_1280,N_1248,N_1269);
xnor U1281 (N_1281,N_1216,N_1225);
and U1282 (N_1282,N_1260,N_1230);
xor U1283 (N_1283,N_1209,N_1244);
or U1284 (N_1284,N_1237,N_1243);
nand U1285 (N_1285,N_1235,N_1267);
nand U1286 (N_1286,N_1264,N_1223);
or U1287 (N_1287,N_1226,N_1261);
and U1288 (N_1288,N_1203,N_1229);
and U1289 (N_1289,N_1272,N_1265);
nand U1290 (N_1290,N_1206,N_1268);
and U1291 (N_1291,N_1263,N_1270);
nand U1292 (N_1292,N_1205,N_1236);
or U1293 (N_1293,N_1232,N_1241);
nand U1294 (N_1294,N_1271,N_1231);
and U1295 (N_1295,N_1274,N_1253);
nor U1296 (N_1296,N_1245,N_1273);
and U1297 (N_1297,N_1242,N_1224);
nand U1298 (N_1298,N_1259,N_1250);
xor U1299 (N_1299,N_1233,N_1221);
nor U1300 (N_1300,N_1251,N_1234);
or U1301 (N_1301,N_1238,N_1207);
nand U1302 (N_1302,N_1239,N_1212);
or U1303 (N_1303,N_1228,N_1256);
nor U1304 (N_1304,N_1204,N_1202);
and U1305 (N_1305,N_1214,N_1258);
nor U1306 (N_1306,N_1217,N_1210);
and U1307 (N_1307,N_1240,N_1247);
and U1308 (N_1308,N_1266,N_1200);
nand U1309 (N_1309,N_1254,N_1255);
nand U1310 (N_1310,N_1262,N_1215);
nand U1311 (N_1311,N_1211,N_1227);
nor U1312 (N_1312,N_1208,N_1266);
or U1313 (N_1313,N_1250,N_1241);
or U1314 (N_1314,N_1212,N_1222);
and U1315 (N_1315,N_1252,N_1234);
nand U1316 (N_1316,N_1227,N_1210);
or U1317 (N_1317,N_1265,N_1216);
nor U1318 (N_1318,N_1250,N_1231);
or U1319 (N_1319,N_1244,N_1231);
nand U1320 (N_1320,N_1235,N_1257);
nor U1321 (N_1321,N_1218,N_1227);
nand U1322 (N_1322,N_1230,N_1248);
and U1323 (N_1323,N_1207,N_1273);
nor U1324 (N_1324,N_1265,N_1252);
nand U1325 (N_1325,N_1211,N_1214);
nor U1326 (N_1326,N_1240,N_1249);
nand U1327 (N_1327,N_1224,N_1262);
nand U1328 (N_1328,N_1262,N_1250);
nand U1329 (N_1329,N_1225,N_1241);
or U1330 (N_1330,N_1200,N_1256);
nor U1331 (N_1331,N_1214,N_1271);
and U1332 (N_1332,N_1239,N_1224);
or U1333 (N_1333,N_1221,N_1240);
and U1334 (N_1334,N_1214,N_1244);
nor U1335 (N_1335,N_1229,N_1224);
nand U1336 (N_1336,N_1213,N_1259);
and U1337 (N_1337,N_1221,N_1252);
and U1338 (N_1338,N_1264,N_1271);
or U1339 (N_1339,N_1218,N_1270);
or U1340 (N_1340,N_1272,N_1231);
and U1341 (N_1341,N_1248,N_1242);
nand U1342 (N_1342,N_1269,N_1251);
or U1343 (N_1343,N_1266,N_1214);
or U1344 (N_1344,N_1249,N_1228);
and U1345 (N_1345,N_1224,N_1234);
and U1346 (N_1346,N_1265,N_1229);
or U1347 (N_1347,N_1257,N_1256);
nor U1348 (N_1348,N_1270,N_1242);
nand U1349 (N_1349,N_1268,N_1202);
nor U1350 (N_1350,N_1339,N_1313);
and U1351 (N_1351,N_1316,N_1320);
nor U1352 (N_1352,N_1318,N_1281);
nor U1353 (N_1353,N_1308,N_1332);
nand U1354 (N_1354,N_1275,N_1323);
and U1355 (N_1355,N_1346,N_1295);
nand U1356 (N_1356,N_1311,N_1335);
or U1357 (N_1357,N_1310,N_1278);
nor U1358 (N_1358,N_1343,N_1300);
nand U1359 (N_1359,N_1324,N_1317);
and U1360 (N_1360,N_1298,N_1342);
or U1361 (N_1361,N_1338,N_1327);
xor U1362 (N_1362,N_1277,N_1293);
or U1363 (N_1363,N_1289,N_1325);
and U1364 (N_1364,N_1345,N_1314);
and U1365 (N_1365,N_1330,N_1292);
nand U1366 (N_1366,N_1309,N_1328);
or U1367 (N_1367,N_1302,N_1287);
nand U1368 (N_1368,N_1334,N_1315);
nand U1369 (N_1369,N_1296,N_1299);
or U1370 (N_1370,N_1336,N_1285);
or U1371 (N_1371,N_1337,N_1344);
nor U1372 (N_1372,N_1301,N_1331);
and U1373 (N_1373,N_1341,N_1321);
nand U1374 (N_1374,N_1312,N_1306);
and U1375 (N_1375,N_1326,N_1282);
and U1376 (N_1376,N_1280,N_1294);
nor U1377 (N_1377,N_1284,N_1283);
and U1378 (N_1378,N_1347,N_1290);
or U1379 (N_1379,N_1286,N_1288);
nand U1380 (N_1380,N_1291,N_1333);
and U1381 (N_1381,N_1276,N_1340);
nor U1382 (N_1382,N_1322,N_1305);
nor U1383 (N_1383,N_1348,N_1329);
nor U1384 (N_1384,N_1307,N_1297);
nor U1385 (N_1385,N_1319,N_1279);
nand U1386 (N_1386,N_1304,N_1303);
and U1387 (N_1387,N_1349,N_1279);
or U1388 (N_1388,N_1302,N_1276);
or U1389 (N_1389,N_1289,N_1330);
and U1390 (N_1390,N_1300,N_1279);
nor U1391 (N_1391,N_1313,N_1333);
xnor U1392 (N_1392,N_1300,N_1325);
and U1393 (N_1393,N_1338,N_1339);
nand U1394 (N_1394,N_1319,N_1344);
xor U1395 (N_1395,N_1304,N_1344);
and U1396 (N_1396,N_1333,N_1324);
nand U1397 (N_1397,N_1309,N_1292);
and U1398 (N_1398,N_1324,N_1345);
nor U1399 (N_1399,N_1305,N_1275);
or U1400 (N_1400,N_1310,N_1329);
and U1401 (N_1401,N_1335,N_1325);
nand U1402 (N_1402,N_1347,N_1346);
nor U1403 (N_1403,N_1294,N_1338);
nand U1404 (N_1404,N_1342,N_1281);
nand U1405 (N_1405,N_1295,N_1344);
and U1406 (N_1406,N_1317,N_1330);
nor U1407 (N_1407,N_1279,N_1285);
nor U1408 (N_1408,N_1328,N_1343);
and U1409 (N_1409,N_1277,N_1321);
nor U1410 (N_1410,N_1328,N_1336);
nor U1411 (N_1411,N_1314,N_1348);
or U1412 (N_1412,N_1327,N_1333);
nand U1413 (N_1413,N_1345,N_1342);
nand U1414 (N_1414,N_1282,N_1345);
nor U1415 (N_1415,N_1278,N_1331);
and U1416 (N_1416,N_1330,N_1291);
or U1417 (N_1417,N_1311,N_1294);
nand U1418 (N_1418,N_1327,N_1320);
nand U1419 (N_1419,N_1296,N_1343);
or U1420 (N_1420,N_1319,N_1333);
xor U1421 (N_1421,N_1298,N_1339);
or U1422 (N_1422,N_1338,N_1315);
and U1423 (N_1423,N_1306,N_1333);
nor U1424 (N_1424,N_1330,N_1285);
or U1425 (N_1425,N_1374,N_1398);
nand U1426 (N_1426,N_1409,N_1360);
nor U1427 (N_1427,N_1389,N_1408);
nor U1428 (N_1428,N_1383,N_1402);
and U1429 (N_1429,N_1373,N_1406);
or U1430 (N_1430,N_1362,N_1416);
nor U1431 (N_1431,N_1407,N_1365);
nor U1432 (N_1432,N_1399,N_1417);
and U1433 (N_1433,N_1394,N_1414);
and U1434 (N_1434,N_1403,N_1397);
nand U1435 (N_1435,N_1387,N_1393);
nand U1436 (N_1436,N_1366,N_1367);
and U1437 (N_1437,N_1368,N_1378);
nand U1438 (N_1438,N_1391,N_1424);
nor U1439 (N_1439,N_1353,N_1359);
or U1440 (N_1440,N_1356,N_1355);
nor U1441 (N_1441,N_1363,N_1351);
xnor U1442 (N_1442,N_1396,N_1415);
xor U1443 (N_1443,N_1405,N_1412);
nor U1444 (N_1444,N_1420,N_1421);
nand U1445 (N_1445,N_1380,N_1375);
or U1446 (N_1446,N_1401,N_1404);
or U1447 (N_1447,N_1400,N_1376);
or U1448 (N_1448,N_1352,N_1390);
nor U1449 (N_1449,N_1370,N_1369);
and U1450 (N_1450,N_1357,N_1377);
and U1451 (N_1451,N_1423,N_1385);
nor U1452 (N_1452,N_1364,N_1379);
nor U1453 (N_1453,N_1410,N_1386);
nand U1454 (N_1454,N_1413,N_1372);
and U1455 (N_1455,N_1392,N_1358);
xnor U1456 (N_1456,N_1388,N_1361);
nor U1457 (N_1457,N_1418,N_1382);
nor U1458 (N_1458,N_1350,N_1411);
nor U1459 (N_1459,N_1395,N_1381);
nor U1460 (N_1460,N_1419,N_1371);
nor U1461 (N_1461,N_1422,N_1354);
and U1462 (N_1462,N_1384,N_1359);
and U1463 (N_1463,N_1419,N_1376);
and U1464 (N_1464,N_1416,N_1352);
or U1465 (N_1465,N_1393,N_1380);
or U1466 (N_1466,N_1370,N_1375);
nor U1467 (N_1467,N_1407,N_1398);
and U1468 (N_1468,N_1415,N_1424);
and U1469 (N_1469,N_1384,N_1365);
nand U1470 (N_1470,N_1382,N_1403);
and U1471 (N_1471,N_1403,N_1385);
nand U1472 (N_1472,N_1380,N_1358);
nand U1473 (N_1473,N_1382,N_1414);
nor U1474 (N_1474,N_1367,N_1361);
or U1475 (N_1475,N_1375,N_1389);
xnor U1476 (N_1476,N_1419,N_1410);
xnor U1477 (N_1477,N_1381,N_1415);
or U1478 (N_1478,N_1350,N_1373);
and U1479 (N_1479,N_1392,N_1356);
xnor U1480 (N_1480,N_1413,N_1362);
and U1481 (N_1481,N_1420,N_1354);
or U1482 (N_1482,N_1363,N_1411);
nand U1483 (N_1483,N_1387,N_1408);
and U1484 (N_1484,N_1392,N_1373);
nand U1485 (N_1485,N_1354,N_1380);
and U1486 (N_1486,N_1400,N_1410);
nor U1487 (N_1487,N_1416,N_1419);
or U1488 (N_1488,N_1376,N_1381);
and U1489 (N_1489,N_1369,N_1389);
nand U1490 (N_1490,N_1387,N_1412);
nand U1491 (N_1491,N_1412,N_1399);
nand U1492 (N_1492,N_1368,N_1383);
and U1493 (N_1493,N_1367,N_1393);
or U1494 (N_1494,N_1364,N_1377);
or U1495 (N_1495,N_1363,N_1417);
nand U1496 (N_1496,N_1407,N_1402);
nand U1497 (N_1497,N_1392,N_1420);
and U1498 (N_1498,N_1387,N_1389);
nor U1499 (N_1499,N_1356,N_1365);
or U1500 (N_1500,N_1483,N_1484);
nand U1501 (N_1501,N_1488,N_1495);
nand U1502 (N_1502,N_1438,N_1462);
xor U1503 (N_1503,N_1459,N_1498);
or U1504 (N_1504,N_1432,N_1426);
and U1505 (N_1505,N_1448,N_1429);
and U1506 (N_1506,N_1430,N_1463);
nand U1507 (N_1507,N_1489,N_1476);
and U1508 (N_1508,N_1445,N_1470);
nor U1509 (N_1509,N_1474,N_1431);
nand U1510 (N_1510,N_1425,N_1433);
nor U1511 (N_1511,N_1471,N_1443);
or U1512 (N_1512,N_1461,N_1475);
or U1513 (N_1513,N_1447,N_1439);
nor U1514 (N_1514,N_1456,N_1493);
or U1515 (N_1515,N_1464,N_1466);
nor U1516 (N_1516,N_1468,N_1444);
nand U1517 (N_1517,N_1460,N_1446);
nand U1518 (N_1518,N_1482,N_1490);
nor U1519 (N_1519,N_1472,N_1496);
nor U1520 (N_1520,N_1435,N_1457);
or U1521 (N_1521,N_1450,N_1497);
nand U1522 (N_1522,N_1458,N_1465);
and U1523 (N_1523,N_1480,N_1434);
nor U1524 (N_1524,N_1479,N_1427);
nor U1525 (N_1525,N_1437,N_1499);
and U1526 (N_1526,N_1494,N_1492);
or U1527 (N_1527,N_1449,N_1477);
or U1528 (N_1528,N_1436,N_1473);
and U1529 (N_1529,N_1491,N_1478);
nor U1530 (N_1530,N_1469,N_1441);
nor U1531 (N_1531,N_1428,N_1485);
or U1532 (N_1532,N_1440,N_1487);
or U1533 (N_1533,N_1486,N_1442);
nor U1534 (N_1534,N_1451,N_1481);
and U1535 (N_1535,N_1467,N_1454);
and U1536 (N_1536,N_1453,N_1452);
nor U1537 (N_1537,N_1455,N_1438);
nor U1538 (N_1538,N_1469,N_1495);
nor U1539 (N_1539,N_1438,N_1472);
nor U1540 (N_1540,N_1472,N_1482);
nand U1541 (N_1541,N_1429,N_1463);
nand U1542 (N_1542,N_1491,N_1475);
and U1543 (N_1543,N_1436,N_1491);
or U1544 (N_1544,N_1469,N_1462);
nor U1545 (N_1545,N_1451,N_1463);
and U1546 (N_1546,N_1425,N_1498);
nor U1547 (N_1547,N_1463,N_1475);
nand U1548 (N_1548,N_1458,N_1461);
nor U1549 (N_1549,N_1473,N_1499);
nand U1550 (N_1550,N_1451,N_1425);
and U1551 (N_1551,N_1443,N_1455);
nand U1552 (N_1552,N_1465,N_1474);
nand U1553 (N_1553,N_1454,N_1478);
nor U1554 (N_1554,N_1434,N_1464);
nor U1555 (N_1555,N_1427,N_1470);
nand U1556 (N_1556,N_1442,N_1452);
nand U1557 (N_1557,N_1465,N_1438);
nand U1558 (N_1558,N_1436,N_1454);
nor U1559 (N_1559,N_1441,N_1456);
nor U1560 (N_1560,N_1461,N_1447);
nand U1561 (N_1561,N_1472,N_1464);
and U1562 (N_1562,N_1481,N_1444);
or U1563 (N_1563,N_1498,N_1437);
xor U1564 (N_1564,N_1491,N_1442);
or U1565 (N_1565,N_1497,N_1449);
nor U1566 (N_1566,N_1431,N_1476);
nand U1567 (N_1567,N_1473,N_1480);
nor U1568 (N_1568,N_1474,N_1454);
or U1569 (N_1569,N_1456,N_1431);
and U1570 (N_1570,N_1474,N_1492);
or U1571 (N_1571,N_1426,N_1482);
xor U1572 (N_1572,N_1479,N_1446);
or U1573 (N_1573,N_1470,N_1431);
and U1574 (N_1574,N_1482,N_1477);
nor U1575 (N_1575,N_1545,N_1525);
or U1576 (N_1576,N_1540,N_1500);
and U1577 (N_1577,N_1538,N_1509);
nor U1578 (N_1578,N_1572,N_1565);
nor U1579 (N_1579,N_1523,N_1567);
or U1580 (N_1580,N_1534,N_1518);
or U1581 (N_1581,N_1529,N_1532);
and U1582 (N_1582,N_1530,N_1553);
and U1583 (N_1583,N_1546,N_1566);
or U1584 (N_1584,N_1558,N_1573);
nor U1585 (N_1585,N_1562,N_1542);
nand U1586 (N_1586,N_1516,N_1536);
nor U1587 (N_1587,N_1574,N_1514);
nand U1588 (N_1588,N_1549,N_1554);
nor U1589 (N_1589,N_1569,N_1510);
xnor U1590 (N_1590,N_1537,N_1543);
nor U1591 (N_1591,N_1519,N_1526);
nand U1592 (N_1592,N_1533,N_1535);
nor U1593 (N_1593,N_1571,N_1524);
and U1594 (N_1594,N_1520,N_1559);
and U1595 (N_1595,N_1561,N_1513);
and U1596 (N_1596,N_1527,N_1552);
and U1597 (N_1597,N_1570,N_1517);
nor U1598 (N_1598,N_1555,N_1557);
and U1599 (N_1599,N_1506,N_1563);
and U1600 (N_1600,N_1551,N_1564);
or U1601 (N_1601,N_1560,N_1539);
nor U1602 (N_1602,N_1502,N_1522);
and U1603 (N_1603,N_1507,N_1548);
nand U1604 (N_1604,N_1512,N_1550);
nand U1605 (N_1605,N_1528,N_1501);
nor U1606 (N_1606,N_1508,N_1515);
or U1607 (N_1607,N_1503,N_1541);
nand U1608 (N_1608,N_1568,N_1521);
and U1609 (N_1609,N_1547,N_1556);
nand U1610 (N_1610,N_1544,N_1511);
or U1611 (N_1611,N_1504,N_1505);
or U1612 (N_1612,N_1531,N_1500);
or U1613 (N_1613,N_1539,N_1534);
nand U1614 (N_1614,N_1562,N_1551);
and U1615 (N_1615,N_1520,N_1526);
nand U1616 (N_1616,N_1574,N_1508);
nor U1617 (N_1617,N_1571,N_1505);
or U1618 (N_1618,N_1532,N_1546);
and U1619 (N_1619,N_1502,N_1558);
nand U1620 (N_1620,N_1557,N_1507);
and U1621 (N_1621,N_1512,N_1532);
and U1622 (N_1622,N_1571,N_1539);
xor U1623 (N_1623,N_1555,N_1520);
nor U1624 (N_1624,N_1540,N_1521);
and U1625 (N_1625,N_1562,N_1529);
nand U1626 (N_1626,N_1532,N_1513);
nand U1627 (N_1627,N_1568,N_1544);
and U1628 (N_1628,N_1548,N_1512);
or U1629 (N_1629,N_1551,N_1571);
and U1630 (N_1630,N_1550,N_1567);
or U1631 (N_1631,N_1554,N_1500);
and U1632 (N_1632,N_1567,N_1514);
nand U1633 (N_1633,N_1535,N_1528);
and U1634 (N_1634,N_1546,N_1514);
xnor U1635 (N_1635,N_1536,N_1572);
nor U1636 (N_1636,N_1553,N_1505);
nor U1637 (N_1637,N_1568,N_1561);
and U1638 (N_1638,N_1500,N_1509);
nand U1639 (N_1639,N_1509,N_1543);
and U1640 (N_1640,N_1556,N_1565);
or U1641 (N_1641,N_1557,N_1566);
and U1642 (N_1642,N_1534,N_1510);
or U1643 (N_1643,N_1531,N_1528);
nor U1644 (N_1644,N_1526,N_1563);
and U1645 (N_1645,N_1513,N_1523);
or U1646 (N_1646,N_1511,N_1525);
or U1647 (N_1647,N_1537,N_1549);
or U1648 (N_1648,N_1569,N_1518);
xor U1649 (N_1649,N_1563,N_1510);
nand U1650 (N_1650,N_1595,N_1581);
nand U1651 (N_1651,N_1623,N_1615);
and U1652 (N_1652,N_1616,N_1629);
nand U1653 (N_1653,N_1618,N_1586);
and U1654 (N_1654,N_1599,N_1635);
and U1655 (N_1655,N_1631,N_1647);
nor U1656 (N_1656,N_1641,N_1626);
and U1657 (N_1657,N_1643,N_1646);
nor U1658 (N_1658,N_1576,N_1598);
nand U1659 (N_1659,N_1608,N_1597);
nor U1660 (N_1660,N_1648,N_1607);
nor U1661 (N_1661,N_1628,N_1632);
and U1662 (N_1662,N_1627,N_1589);
or U1663 (N_1663,N_1634,N_1606);
nor U1664 (N_1664,N_1590,N_1584);
or U1665 (N_1665,N_1620,N_1644);
nor U1666 (N_1666,N_1575,N_1630);
nand U1667 (N_1667,N_1610,N_1614);
or U1668 (N_1668,N_1594,N_1613);
nor U1669 (N_1669,N_1633,N_1611);
nor U1670 (N_1670,N_1621,N_1591);
or U1671 (N_1671,N_1582,N_1649);
and U1672 (N_1672,N_1602,N_1639);
nand U1673 (N_1673,N_1588,N_1624);
xnor U1674 (N_1674,N_1585,N_1580);
nor U1675 (N_1675,N_1600,N_1579);
or U1676 (N_1676,N_1619,N_1578);
nor U1677 (N_1677,N_1601,N_1596);
and U1678 (N_1678,N_1592,N_1642);
and U1679 (N_1679,N_1587,N_1625);
nor U1680 (N_1680,N_1605,N_1583);
nand U1681 (N_1681,N_1638,N_1609);
or U1682 (N_1682,N_1636,N_1603);
nand U1683 (N_1683,N_1640,N_1617);
nor U1684 (N_1684,N_1577,N_1593);
nor U1685 (N_1685,N_1637,N_1604);
and U1686 (N_1686,N_1612,N_1622);
nand U1687 (N_1687,N_1645,N_1594);
and U1688 (N_1688,N_1636,N_1601);
or U1689 (N_1689,N_1594,N_1644);
or U1690 (N_1690,N_1626,N_1599);
nor U1691 (N_1691,N_1613,N_1581);
or U1692 (N_1692,N_1648,N_1581);
and U1693 (N_1693,N_1633,N_1605);
nand U1694 (N_1694,N_1577,N_1640);
and U1695 (N_1695,N_1578,N_1614);
nor U1696 (N_1696,N_1600,N_1587);
nor U1697 (N_1697,N_1609,N_1588);
and U1698 (N_1698,N_1645,N_1609);
nor U1699 (N_1699,N_1606,N_1620);
or U1700 (N_1700,N_1588,N_1639);
xnor U1701 (N_1701,N_1617,N_1592);
or U1702 (N_1702,N_1623,N_1632);
nand U1703 (N_1703,N_1594,N_1636);
nor U1704 (N_1704,N_1592,N_1601);
nor U1705 (N_1705,N_1589,N_1649);
and U1706 (N_1706,N_1591,N_1627);
nor U1707 (N_1707,N_1584,N_1644);
xnor U1708 (N_1708,N_1645,N_1577);
and U1709 (N_1709,N_1642,N_1606);
and U1710 (N_1710,N_1576,N_1619);
nand U1711 (N_1711,N_1611,N_1598);
and U1712 (N_1712,N_1639,N_1587);
or U1713 (N_1713,N_1606,N_1598);
and U1714 (N_1714,N_1609,N_1627);
and U1715 (N_1715,N_1622,N_1644);
nor U1716 (N_1716,N_1615,N_1606);
and U1717 (N_1717,N_1626,N_1595);
or U1718 (N_1718,N_1622,N_1614);
xnor U1719 (N_1719,N_1575,N_1610);
or U1720 (N_1720,N_1608,N_1592);
and U1721 (N_1721,N_1629,N_1597);
or U1722 (N_1722,N_1611,N_1607);
and U1723 (N_1723,N_1642,N_1646);
and U1724 (N_1724,N_1616,N_1632);
and U1725 (N_1725,N_1684,N_1677);
and U1726 (N_1726,N_1718,N_1700);
and U1727 (N_1727,N_1679,N_1669);
and U1728 (N_1728,N_1690,N_1720);
and U1729 (N_1729,N_1656,N_1701);
nor U1730 (N_1730,N_1652,N_1672);
or U1731 (N_1731,N_1667,N_1710);
xor U1732 (N_1732,N_1716,N_1681);
or U1733 (N_1733,N_1658,N_1680);
or U1734 (N_1734,N_1707,N_1676);
nand U1735 (N_1735,N_1671,N_1685);
nand U1736 (N_1736,N_1703,N_1666);
nor U1737 (N_1737,N_1661,N_1668);
nand U1738 (N_1738,N_1651,N_1712);
nand U1739 (N_1739,N_1653,N_1663);
nor U1740 (N_1740,N_1691,N_1678);
xnor U1741 (N_1741,N_1713,N_1686);
nand U1742 (N_1742,N_1662,N_1655);
nand U1743 (N_1743,N_1705,N_1689);
nand U1744 (N_1744,N_1714,N_1660);
nor U1745 (N_1745,N_1715,N_1670);
or U1746 (N_1746,N_1650,N_1675);
and U1747 (N_1747,N_1708,N_1722);
nand U1748 (N_1748,N_1665,N_1699);
nand U1749 (N_1749,N_1706,N_1695);
xor U1750 (N_1750,N_1709,N_1674);
xor U1751 (N_1751,N_1654,N_1688);
or U1752 (N_1752,N_1693,N_1664);
nor U1753 (N_1753,N_1698,N_1719);
or U1754 (N_1754,N_1659,N_1702);
nand U1755 (N_1755,N_1711,N_1683);
or U1756 (N_1756,N_1721,N_1696);
or U1757 (N_1757,N_1657,N_1697);
nand U1758 (N_1758,N_1694,N_1682);
nor U1759 (N_1759,N_1673,N_1723);
or U1760 (N_1760,N_1704,N_1687);
or U1761 (N_1761,N_1692,N_1717);
nor U1762 (N_1762,N_1724,N_1705);
or U1763 (N_1763,N_1653,N_1691);
nand U1764 (N_1764,N_1711,N_1720);
or U1765 (N_1765,N_1692,N_1701);
nand U1766 (N_1766,N_1702,N_1719);
nand U1767 (N_1767,N_1710,N_1682);
nor U1768 (N_1768,N_1674,N_1664);
nand U1769 (N_1769,N_1675,N_1696);
and U1770 (N_1770,N_1701,N_1711);
or U1771 (N_1771,N_1684,N_1702);
or U1772 (N_1772,N_1713,N_1672);
nand U1773 (N_1773,N_1677,N_1708);
and U1774 (N_1774,N_1714,N_1683);
nor U1775 (N_1775,N_1720,N_1670);
and U1776 (N_1776,N_1720,N_1661);
nor U1777 (N_1777,N_1683,N_1687);
nand U1778 (N_1778,N_1672,N_1676);
nor U1779 (N_1779,N_1667,N_1658);
nor U1780 (N_1780,N_1688,N_1707);
nand U1781 (N_1781,N_1652,N_1702);
nand U1782 (N_1782,N_1663,N_1706);
or U1783 (N_1783,N_1655,N_1705);
or U1784 (N_1784,N_1687,N_1724);
nand U1785 (N_1785,N_1661,N_1667);
and U1786 (N_1786,N_1675,N_1667);
and U1787 (N_1787,N_1703,N_1655);
and U1788 (N_1788,N_1713,N_1699);
and U1789 (N_1789,N_1718,N_1659);
or U1790 (N_1790,N_1688,N_1650);
nand U1791 (N_1791,N_1678,N_1667);
or U1792 (N_1792,N_1659,N_1695);
or U1793 (N_1793,N_1652,N_1717);
nand U1794 (N_1794,N_1718,N_1672);
nand U1795 (N_1795,N_1704,N_1670);
nor U1796 (N_1796,N_1724,N_1654);
or U1797 (N_1797,N_1669,N_1694);
nor U1798 (N_1798,N_1658,N_1674);
and U1799 (N_1799,N_1677,N_1670);
nand U1800 (N_1800,N_1735,N_1763);
nand U1801 (N_1801,N_1755,N_1794);
and U1802 (N_1802,N_1761,N_1745);
nor U1803 (N_1803,N_1797,N_1758);
and U1804 (N_1804,N_1744,N_1726);
nand U1805 (N_1805,N_1736,N_1770);
nand U1806 (N_1806,N_1767,N_1799);
nand U1807 (N_1807,N_1731,N_1741);
or U1808 (N_1808,N_1789,N_1793);
or U1809 (N_1809,N_1787,N_1784);
xnor U1810 (N_1810,N_1768,N_1757);
and U1811 (N_1811,N_1746,N_1769);
nand U1812 (N_1812,N_1773,N_1747);
and U1813 (N_1813,N_1764,N_1756);
or U1814 (N_1814,N_1738,N_1730);
nor U1815 (N_1815,N_1743,N_1739);
nand U1816 (N_1816,N_1792,N_1729);
or U1817 (N_1817,N_1786,N_1725);
and U1818 (N_1818,N_1778,N_1788);
and U1819 (N_1819,N_1733,N_1762);
nand U1820 (N_1820,N_1765,N_1748);
or U1821 (N_1821,N_1790,N_1795);
and U1822 (N_1822,N_1752,N_1777);
nor U1823 (N_1823,N_1740,N_1782);
nor U1824 (N_1824,N_1732,N_1759);
nand U1825 (N_1825,N_1780,N_1781);
or U1826 (N_1826,N_1779,N_1742);
and U1827 (N_1827,N_1751,N_1774);
or U1828 (N_1828,N_1728,N_1771);
nor U1829 (N_1829,N_1785,N_1734);
nand U1830 (N_1830,N_1791,N_1727);
nand U1831 (N_1831,N_1783,N_1737);
and U1832 (N_1832,N_1749,N_1775);
nand U1833 (N_1833,N_1766,N_1772);
or U1834 (N_1834,N_1796,N_1753);
and U1835 (N_1835,N_1798,N_1760);
or U1836 (N_1836,N_1776,N_1750);
and U1837 (N_1837,N_1754,N_1741);
nor U1838 (N_1838,N_1764,N_1780);
nand U1839 (N_1839,N_1738,N_1791);
or U1840 (N_1840,N_1736,N_1756);
nor U1841 (N_1841,N_1775,N_1770);
nand U1842 (N_1842,N_1788,N_1755);
nand U1843 (N_1843,N_1797,N_1782);
and U1844 (N_1844,N_1771,N_1732);
nand U1845 (N_1845,N_1765,N_1750);
nor U1846 (N_1846,N_1731,N_1776);
and U1847 (N_1847,N_1798,N_1730);
and U1848 (N_1848,N_1727,N_1741);
nor U1849 (N_1849,N_1749,N_1781);
nor U1850 (N_1850,N_1738,N_1775);
and U1851 (N_1851,N_1750,N_1759);
and U1852 (N_1852,N_1751,N_1775);
nor U1853 (N_1853,N_1749,N_1798);
nor U1854 (N_1854,N_1789,N_1784);
nand U1855 (N_1855,N_1793,N_1754);
and U1856 (N_1856,N_1761,N_1740);
nor U1857 (N_1857,N_1730,N_1789);
or U1858 (N_1858,N_1726,N_1733);
nand U1859 (N_1859,N_1766,N_1785);
or U1860 (N_1860,N_1760,N_1792);
or U1861 (N_1861,N_1751,N_1770);
nand U1862 (N_1862,N_1737,N_1760);
and U1863 (N_1863,N_1775,N_1756);
or U1864 (N_1864,N_1797,N_1755);
and U1865 (N_1865,N_1739,N_1755);
and U1866 (N_1866,N_1757,N_1740);
xnor U1867 (N_1867,N_1754,N_1730);
and U1868 (N_1868,N_1771,N_1791);
nand U1869 (N_1869,N_1728,N_1798);
nand U1870 (N_1870,N_1726,N_1762);
nor U1871 (N_1871,N_1783,N_1763);
nor U1872 (N_1872,N_1759,N_1795);
nor U1873 (N_1873,N_1746,N_1760);
nand U1874 (N_1874,N_1727,N_1781);
and U1875 (N_1875,N_1835,N_1839);
or U1876 (N_1876,N_1873,N_1831);
and U1877 (N_1877,N_1820,N_1810);
or U1878 (N_1878,N_1809,N_1866);
or U1879 (N_1879,N_1857,N_1842);
nor U1880 (N_1880,N_1858,N_1836);
and U1881 (N_1881,N_1832,N_1814);
and U1882 (N_1882,N_1867,N_1871);
nand U1883 (N_1883,N_1843,N_1850);
nor U1884 (N_1884,N_1841,N_1860);
nor U1885 (N_1885,N_1816,N_1827);
and U1886 (N_1886,N_1854,N_1833);
or U1887 (N_1887,N_1869,N_1856);
and U1888 (N_1888,N_1802,N_1830);
nor U1889 (N_1889,N_1828,N_1864);
nor U1890 (N_1890,N_1812,N_1853);
nor U1891 (N_1891,N_1819,N_1824);
nor U1892 (N_1892,N_1818,N_1822);
or U1893 (N_1893,N_1817,N_1813);
or U1894 (N_1894,N_1805,N_1815);
and U1895 (N_1895,N_1862,N_1859);
or U1896 (N_1896,N_1825,N_1840);
or U1897 (N_1897,N_1870,N_1849);
nand U1898 (N_1898,N_1845,N_1811);
and U1899 (N_1899,N_1851,N_1838);
and U1900 (N_1900,N_1855,N_1801);
nand U1901 (N_1901,N_1861,N_1808);
nor U1902 (N_1902,N_1872,N_1803);
nor U1903 (N_1903,N_1834,N_1868);
or U1904 (N_1904,N_1821,N_1837);
or U1905 (N_1905,N_1852,N_1865);
nand U1906 (N_1906,N_1844,N_1846);
or U1907 (N_1907,N_1807,N_1806);
nor U1908 (N_1908,N_1823,N_1826);
or U1909 (N_1909,N_1804,N_1863);
nor U1910 (N_1910,N_1874,N_1829);
nand U1911 (N_1911,N_1848,N_1800);
nor U1912 (N_1912,N_1847,N_1819);
nor U1913 (N_1913,N_1846,N_1863);
nand U1914 (N_1914,N_1845,N_1860);
nor U1915 (N_1915,N_1871,N_1814);
and U1916 (N_1916,N_1832,N_1836);
nand U1917 (N_1917,N_1849,N_1847);
nor U1918 (N_1918,N_1817,N_1871);
and U1919 (N_1919,N_1840,N_1801);
nor U1920 (N_1920,N_1840,N_1871);
or U1921 (N_1921,N_1831,N_1825);
or U1922 (N_1922,N_1821,N_1835);
nand U1923 (N_1923,N_1850,N_1874);
or U1924 (N_1924,N_1851,N_1869);
or U1925 (N_1925,N_1833,N_1857);
nand U1926 (N_1926,N_1865,N_1851);
and U1927 (N_1927,N_1813,N_1810);
or U1928 (N_1928,N_1851,N_1846);
and U1929 (N_1929,N_1824,N_1800);
and U1930 (N_1930,N_1849,N_1865);
nand U1931 (N_1931,N_1850,N_1845);
nand U1932 (N_1932,N_1811,N_1865);
nand U1933 (N_1933,N_1822,N_1831);
nor U1934 (N_1934,N_1804,N_1842);
and U1935 (N_1935,N_1857,N_1829);
nor U1936 (N_1936,N_1864,N_1860);
and U1937 (N_1937,N_1822,N_1827);
nor U1938 (N_1938,N_1854,N_1864);
and U1939 (N_1939,N_1808,N_1832);
and U1940 (N_1940,N_1821,N_1866);
or U1941 (N_1941,N_1852,N_1862);
nor U1942 (N_1942,N_1862,N_1815);
nand U1943 (N_1943,N_1805,N_1830);
or U1944 (N_1944,N_1866,N_1865);
nand U1945 (N_1945,N_1850,N_1844);
and U1946 (N_1946,N_1831,N_1827);
or U1947 (N_1947,N_1819,N_1811);
or U1948 (N_1948,N_1846,N_1862);
nor U1949 (N_1949,N_1816,N_1841);
nand U1950 (N_1950,N_1942,N_1879);
nor U1951 (N_1951,N_1906,N_1930);
or U1952 (N_1952,N_1927,N_1903);
and U1953 (N_1953,N_1895,N_1911);
nand U1954 (N_1954,N_1889,N_1886);
nand U1955 (N_1955,N_1934,N_1890);
or U1956 (N_1956,N_1932,N_1929);
xor U1957 (N_1957,N_1936,N_1938);
and U1958 (N_1958,N_1905,N_1882);
nand U1959 (N_1959,N_1915,N_1909);
and U1960 (N_1960,N_1908,N_1902);
nor U1961 (N_1961,N_1896,N_1937);
and U1962 (N_1962,N_1875,N_1918);
nand U1963 (N_1963,N_1887,N_1926);
and U1964 (N_1964,N_1904,N_1913);
or U1965 (N_1965,N_1894,N_1898);
nor U1966 (N_1966,N_1924,N_1919);
or U1967 (N_1967,N_1912,N_1883);
xor U1968 (N_1968,N_1935,N_1893);
or U1969 (N_1969,N_1925,N_1910);
or U1970 (N_1970,N_1917,N_1897);
and U1971 (N_1971,N_1949,N_1914);
nand U1972 (N_1972,N_1944,N_1900);
nand U1973 (N_1973,N_1878,N_1939);
nor U1974 (N_1974,N_1943,N_1907);
nand U1975 (N_1975,N_1899,N_1877);
nand U1976 (N_1976,N_1941,N_1880);
nand U1977 (N_1977,N_1947,N_1920);
nand U1978 (N_1978,N_1916,N_1885);
and U1979 (N_1979,N_1923,N_1876);
nor U1980 (N_1980,N_1884,N_1891);
or U1981 (N_1981,N_1928,N_1922);
and U1982 (N_1982,N_1948,N_1892);
nor U1983 (N_1983,N_1933,N_1881);
nand U1984 (N_1984,N_1888,N_1946);
xnor U1985 (N_1985,N_1901,N_1945);
or U1986 (N_1986,N_1931,N_1940);
nand U1987 (N_1987,N_1921,N_1926);
nor U1988 (N_1988,N_1889,N_1890);
nor U1989 (N_1989,N_1876,N_1929);
nand U1990 (N_1990,N_1886,N_1906);
nand U1991 (N_1991,N_1888,N_1932);
or U1992 (N_1992,N_1946,N_1902);
or U1993 (N_1993,N_1938,N_1922);
nor U1994 (N_1994,N_1901,N_1895);
nor U1995 (N_1995,N_1926,N_1915);
nor U1996 (N_1996,N_1904,N_1934);
nor U1997 (N_1997,N_1934,N_1876);
nand U1998 (N_1998,N_1900,N_1887);
and U1999 (N_1999,N_1931,N_1893);
nor U2000 (N_2000,N_1909,N_1944);
nor U2001 (N_2001,N_1907,N_1938);
and U2002 (N_2002,N_1941,N_1921);
nor U2003 (N_2003,N_1928,N_1889);
and U2004 (N_2004,N_1898,N_1909);
nand U2005 (N_2005,N_1882,N_1902);
or U2006 (N_2006,N_1909,N_1928);
or U2007 (N_2007,N_1929,N_1885);
and U2008 (N_2008,N_1949,N_1925);
nand U2009 (N_2009,N_1933,N_1937);
or U2010 (N_2010,N_1880,N_1933);
or U2011 (N_2011,N_1934,N_1920);
nor U2012 (N_2012,N_1917,N_1924);
nand U2013 (N_2013,N_1915,N_1912);
nand U2014 (N_2014,N_1904,N_1917);
or U2015 (N_2015,N_1945,N_1898);
nor U2016 (N_2016,N_1884,N_1896);
nand U2017 (N_2017,N_1885,N_1948);
nor U2018 (N_2018,N_1914,N_1947);
nor U2019 (N_2019,N_1896,N_1883);
or U2020 (N_2020,N_1893,N_1911);
nor U2021 (N_2021,N_1904,N_1899);
nor U2022 (N_2022,N_1935,N_1934);
nand U2023 (N_2023,N_1889,N_1929);
nand U2024 (N_2024,N_1944,N_1885);
nor U2025 (N_2025,N_1992,N_2002);
nand U2026 (N_2026,N_2022,N_1981);
nand U2027 (N_2027,N_1965,N_1969);
and U2028 (N_2028,N_1971,N_1975);
or U2029 (N_2029,N_2015,N_2017);
nand U2030 (N_2030,N_2024,N_2009);
nor U2031 (N_2031,N_1991,N_2006);
or U2032 (N_2032,N_1976,N_1953);
nand U2033 (N_2033,N_1983,N_1951);
xor U2034 (N_2034,N_1968,N_2003);
or U2035 (N_2035,N_2000,N_2013);
and U2036 (N_2036,N_1986,N_2018);
nand U2037 (N_2037,N_2023,N_1972);
or U2038 (N_2038,N_2007,N_1978);
xnor U2039 (N_2039,N_1979,N_1954);
xnor U2040 (N_2040,N_1990,N_1985);
nand U2041 (N_2041,N_1955,N_1959);
nor U2042 (N_2042,N_1987,N_1996);
nor U2043 (N_2043,N_1950,N_1966);
and U2044 (N_2044,N_1970,N_1961);
and U2045 (N_2045,N_1974,N_2016);
or U2046 (N_2046,N_1962,N_2001);
nand U2047 (N_2047,N_2019,N_1999);
and U2048 (N_2048,N_1982,N_1956);
and U2049 (N_2049,N_2014,N_1967);
and U2050 (N_2050,N_2012,N_1952);
nand U2051 (N_2051,N_1963,N_1964);
xor U2052 (N_2052,N_1984,N_1980);
nand U2053 (N_2053,N_1993,N_1988);
nand U2054 (N_2054,N_2020,N_1957);
nor U2055 (N_2055,N_2021,N_1995);
nand U2056 (N_2056,N_1960,N_2004);
or U2057 (N_2057,N_1989,N_2008);
and U2058 (N_2058,N_2005,N_1998);
and U2059 (N_2059,N_1973,N_1994);
nand U2060 (N_2060,N_2011,N_2010);
and U2061 (N_2061,N_1958,N_1977);
nand U2062 (N_2062,N_1997,N_2001);
and U2063 (N_2063,N_1958,N_1999);
and U2064 (N_2064,N_1961,N_1962);
nor U2065 (N_2065,N_2020,N_2004);
or U2066 (N_2066,N_1981,N_1958);
nand U2067 (N_2067,N_1950,N_2018);
and U2068 (N_2068,N_1972,N_2005);
nand U2069 (N_2069,N_2008,N_1981);
nand U2070 (N_2070,N_1975,N_2017);
nor U2071 (N_2071,N_1984,N_1981);
xnor U2072 (N_2072,N_2024,N_2012);
nand U2073 (N_2073,N_2023,N_2004);
xnor U2074 (N_2074,N_1985,N_1974);
and U2075 (N_2075,N_1973,N_1998);
or U2076 (N_2076,N_2021,N_2019);
nor U2077 (N_2077,N_1988,N_1969);
or U2078 (N_2078,N_2000,N_1999);
and U2079 (N_2079,N_1997,N_2023);
and U2080 (N_2080,N_1982,N_1985);
or U2081 (N_2081,N_1950,N_1996);
and U2082 (N_2082,N_1969,N_2007);
or U2083 (N_2083,N_2012,N_1964);
and U2084 (N_2084,N_1971,N_2008);
nor U2085 (N_2085,N_2013,N_1964);
nor U2086 (N_2086,N_1974,N_1968);
xnor U2087 (N_2087,N_1967,N_1966);
nor U2088 (N_2088,N_2001,N_2003);
or U2089 (N_2089,N_2014,N_1964);
or U2090 (N_2090,N_1955,N_1996);
nand U2091 (N_2091,N_1952,N_1964);
or U2092 (N_2092,N_2024,N_2005);
or U2093 (N_2093,N_1976,N_1962);
nand U2094 (N_2094,N_1966,N_1983);
xnor U2095 (N_2095,N_2007,N_2017);
nand U2096 (N_2096,N_1997,N_2018);
and U2097 (N_2097,N_1963,N_1983);
and U2098 (N_2098,N_1970,N_1972);
nand U2099 (N_2099,N_1987,N_2018);
nor U2100 (N_2100,N_2077,N_2033);
and U2101 (N_2101,N_2095,N_2034);
and U2102 (N_2102,N_2087,N_2073);
nor U2103 (N_2103,N_2075,N_2091);
nor U2104 (N_2104,N_2064,N_2049);
nand U2105 (N_2105,N_2042,N_2030);
nor U2106 (N_2106,N_2084,N_2056);
nand U2107 (N_2107,N_2040,N_2089);
nor U2108 (N_2108,N_2031,N_2086);
or U2109 (N_2109,N_2041,N_2055);
nand U2110 (N_2110,N_2036,N_2026);
and U2111 (N_2111,N_2092,N_2079);
and U2112 (N_2112,N_2094,N_2047);
nand U2113 (N_2113,N_2076,N_2096);
nor U2114 (N_2114,N_2057,N_2070);
and U2115 (N_2115,N_2058,N_2062);
or U2116 (N_2116,N_2082,N_2068);
xor U2117 (N_2117,N_2078,N_2083);
nand U2118 (N_2118,N_2032,N_2061);
and U2119 (N_2119,N_2069,N_2037);
nand U2120 (N_2120,N_2098,N_2044);
or U2121 (N_2121,N_2090,N_2060);
nand U2122 (N_2122,N_2097,N_2045);
and U2123 (N_2123,N_2051,N_2099);
or U2124 (N_2124,N_2054,N_2067);
and U2125 (N_2125,N_2028,N_2072);
nand U2126 (N_2126,N_2039,N_2088);
nand U2127 (N_2127,N_2050,N_2066);
or U2128 (N_2128,N_2053,N_2080);
nor U2129 (N_2129,N_2093,N_2046);
nand U2130 (N_2130,N_2052,N_2074);
nor U2131 (N_2131,N_2063,N_2027);
nor U2132 (N_2132,N_2071,N_2025);
and U2133 (N_2133,N_2059,N_2048);
or U2134 (N_2134,N_2081,N_2038);
or U2135 (N_2135,N_2065,N_2029);
xor U2136 (N_2136,N_2035,N_2085);
nor U2137 (N_2137,N_2043,N_2045);
nor U2138 (N_2138,N_2094,N_2064);
nor U2139 (N_2139,N_2054,N_2029);
nor U2140 (N_2140,N_2026,N_2059);
or U2141 (N_2141,N_2056,N_2037);
nand U2142 (N_2142,N_2093,N_2076);
or U2143 (N_2143,N_2092,N_2058);
or U2144 (N_2144,N_2053,N_2042);
nand U2145 (N_2145,N_2094,N_2036);
nor U2146 (N_2146,N_2074,N_2094);
nand U2147 (N_2147,N_2029,N_2082);
and U2148 (N_2148,N_2083,N_2068);
nand U2149 (N_2149,N_2066,N_2095);
nor U2150 (N_2150,N_2088,N_2084);
nand U2151 (N_2151,N_2030,N_2038);
and U2152 (N_2152,N_2078,N_2080);
nor U2153 (N_2153,N_2049,N_2038);
and U2154 (N_2154,N_2075,N_2078);
and U2155 (N_2155,N_2070,N_2079);
nand U2156 (N_2156,N_2060,N_2026);
xor U2157 (N_2157,N_2065,N_2082);
nor U2158 (N_2158,N_2070,N_2041);
nand U2159 (N_2159,N_2097,N_2099);
and U2160 (N_2160,N_2084,N_2082);
and U2161 (N_2161,N_2035,N_2091);
and U2162 (N_2162,N_2058,N_2056);
or U2163 (N_2163,N_2091,N_2094);
or U2164 (N_2164,N_2069,N_2068);
or U2165 (N_2165,N_2057,N_2039);
and U2166 (N_2166,N_2025,N_2085);
or U2167 (N_2167,N_2033,N_2078);
or U2168 (N_2168,N_2042,N_2069);
and U2169 (N_2169,N_2072,N_2032);
and U2170 (N_2170,N_2093,N_2029);
nand U2171 (N_2171,N_2028,N_2048);
or U2172 (N_2172,N_2034,N_2086);
and U2173 (N_2173,N_2078,N_2067);
and U2174 (N_2174,N_2098,N_2072);
xor U2175 (N_2175,N_2121,N_2153);
nand U2176 (N_2176,N_2102,N_2145);
nor U2177 (N_2177,N_2113,N_2104);
nor U2178 (N_2178,N_2157,N_2118);
nor U2179 (N_2179,N_2106,N_2168);
and U2180 (N_2180,N_2125,N_2101);
nand U2181 (N_2181,N_2116,N_2149);
and U2182 (N_2182,N_2109,N_2172);
and U2183 (N_2183,N_2173,N_2117);
or U2184 (N_2184,N_2110,N_2140);
nand U2185 (N_2185,N_2166,N_2135);
nor U2186 (N_2186,N_2141,N_2114);
or U2187 (N_2187,N_2122,N_2151);
nand U2188 (N_2188,N_2128,N_2161);
and U2189 (N_2189,N_2138,N_2144);
or U2190 (N_2190,N_2164,N_2165);
and U2191 (N_2191,N_2124,N_2103);
or U2192 (N_2192,N_2156,N_2120);
nand U2193 (N_2193,N_2100,N_2171);
nand U2194 (N_2194,N_2148,N_2162);
nand U2195 (N_2195,N_2143,N_2142);
or U2196 (N_2196,N_2127,N_2158);
and U2197 (N_2197,N_2159,N_2137);
and U2198 (N_2198,N_2131,N_2150);
or U2199 (N_2199,N_2169,N_2152);
nand U2200 (N_2200,N_2107,N_2108);
or U2201 (N_2201,N_2126,N_2154);
and U2202 (N_2202,N_2147,N_2167);
nand U2203 (N_2203,N_2163,N_2132);
or U2204 (N_2204,N_2111,N_2160);
or U2205 (N_2205,N_2115,N_2130);
nor U2206 (N_2206,N_2129,N_2136);
nand U2207 (N_2207,N_2105,N_2133);
and U2208 (N_2208,N_2112,N_2123);
and U2209 (N_2209,N_2174,N_2119);
nor U2210 (N_2210,N_2146,N_2170);
and U2211 (N_2211,N_2134,N_2155);
nor U2212 (N_2212,N_2139,N_2155);
or U2213 (N_2213,N_2153,N_2168);
or U2214 (N_2214,N_2164,N_2103);
nand U2215 (N_2215,N_2166,N_2151);
nand U2216 (N_2216,N_2167,N_2104);
nand U2217 (N_2217,N_2107,N_2133);
nor U2218 (N_2218,N_2108,N_2127);
nor U2219 (N_2219,N_2118,N_2115);
nand U2220 (N_2220,N_2132,N_2169);
nand U2221 (N_2221,N_2124,N_2153);
and U2222 (N_2222,N_2127,N_2143);
or U2223 (N_2223,N_2117,N_2163);
nand U2224 (N_2224,N_2128,N_2158);
nand U2225 (N_2225,N_2148,N_2123);
and U2226 (N_2226,N_2130,N_2165);
nand U2227 (N_2227,N_2161,N_2143);
nand U2228 (N_2228,N_2105,N_2166);
nand U2229 (N_2229,N_2125,N_2104);
or U2230 (N_2230,N_2107,N_2137);
nor U2231 (N_2231,N_2107,N_2112);
nand U2232 (N_2232,N_2135,N_2170);
and U2233 (N_2233,N_2112,N_2173);
nand U2234 (N_2234,N_2163,N_2145);
and U2235 (N_2235,N_2162,N_2158);
and U2236 (N_2236,N_2112,N_2129);
nand U2237 (N_2237,N_2152,N_2162);
and U2238 (N_2238,N_2146,N_2112);
nand U2239 (N_2239,N_2103,N_2155);
nor U2240 (N_2240,N_2137,N_2134);
nor U2241 (N_2241,N_2113,N_2173);
and U2242 (N_2242,N_2174,N_2130);
and U2243 (N_2243,N_2133,N_2106);
nor U2244 (N_2244,N_2117,N_2165);
and U2245 (N_2245,N_2171,N_2173);
or U2246 (N_2246,N_2120,N_2141);
or U2247 (N_2247,N_2105,N_2159);
nand U2248 (N_2248,N_2106,N_2165);
nand U2249 (N_2249,N_2129,N_2111);
or U2250 (N_2250,N_2220,N_2206);
and U2251 (N_2251,N_2215,N_2186);
nor U2252 (N_2252,N_2241,N_2199);
or U2253 (N_2253,N_2222,N_2224);
nand U2254 (N_2254,N_2190,N_2242);
xnor U2255 (N_2255,N_2201,N_2209);
or U2256 (N_2256,N_2177,N_2179);
and U2257 (N_2257,N_2226,N_2195);
nor U2258 (N_2258,N_2188,N_2247);
or U2259 (N_2259,N_2248,N_2194);
and U2260 (N_2260,N_2211,N_2230);
or U2261 (N_2261,N_2185,N_2229);
nand U2262 (N_2262,N_2200,N_2181);
nor U2263 (N_2263,N_2180,N_2225);
nor U2264 (N_2264,N_2236,N_2193);
and U2265 (N_2265,N_2192,N_2249);
or U2266 (N_2266,N_2205,N_2234);
nor U2267 (N_2267,N_2191,N_2232);
and U2268 (N_2268,N_2237,N_2175);
or U2269 (N_2269,N_2184,N_2218);
and U2270 (N_2270,N_2228,N_2212);
or U2271 (N_2271,N_2223,N_2219);
nor U2272 (N_2272,N_2187,N_2214);
nor U2273 (N_2273,N_2235,N_2246);
and U2274 (N_2274,N_2208,N_2231);
nor U2275 (N_2275,N_2221,N_2217);
nor U2276 (N_2276,N_2197,N_2207);
nand U2277 (N_2277,N_2213,N_2198);
or U2278 (N_2278,N_2239,N_2240);
nand U2279 (N_2279,N_2202,N_2176);
and U2280 (N_2280,N_2196,N_2210);
nor U2281 (N_2281,N_2245,N_2244);
or U2282 (N_2282,N_2216,N_2233);
and U2283 (N_2283,N_2238,N_2178);
nor U2284 (N_2284,N_2189,N_2183);
nor U2285 (N_2285,N_2204,N_2227);
nand U2286 (N_2286,N_2203,N_2243);
nor U2287 (N_2287,N_2182,N_2190);
and U2288 (N_2288,N_2190,N_2206);
and U2289 (N_2289,N_2193,N_2175);
and U2290 (N_2290,N_2214,N_2194);
or U2291 (N_2291,N_2186,N_2197);
or U2292 (N_2292,N_2210,N_2204);
nand U2293 (N_2293,N_2232,N_2192);
xnor U2294 (N_2294,N_2213,N_2179);
or U2295 (N_2295,N_2205,N_2189);
and U2296 (N_2296,N_2175,N_2241);
and U2297 (N_2297,N_2180,N_2240);
and U2298 (N_2298,N_2214,N_2199);
nand U2299 (N_2299,N_2232,N_2180);
nor U2300 (N_2300,N_2223,N_2221);
nand U2301 (N_2301,N_2230,N_2218);
xor U2302 (N_2302,N_2182,N_2223);
or U2303 (N_2303,N_2244,N_2213);
nand U2304 (N_2304,N_2245,N_2228);
nor U2305 (N_2305,N_2214,N_2223);
nor U2306 (N_2306,N_2201,N_2240);
nand U2307 (N_2307,N_2183,N_2208);
or U2308 (N_2308,N_2187,N_2243);
nand U2309 (N_2309,N_2225,N_2188);
or U2310 (N_2310,N_2192,N_2245);
and U2311 (N_2311,N_2183,N_2232);
or U2312 (N_2312,N_2198,N_2200);
or U2313 (N_2313,N_2207,N_2249);
nand U2314 (N_2314,N_2199,N_2235);
xnor U2315 (N_2315,N_2219,N_2195);
nor U2316 (N_2316,N_2218,N_2219);
nor U2317 (N_2317,N_2240,N_2204);
xor U2318 (N_2318,N_2218,N_2217);
and U2319 (N_2319,N_2238,N_2235);
nand U2320 (N_2320,N_2210,N_2186);
nor U2321 (N_2321,N_2209,N_2211);
nand U2322 (N_2322,N_2223,N_2210);
nor U2323 (N_2323,N_2179,N_2239);
or U2324 (N_2324,N_2183,N_2202);
and U2325 (N_2325,N_2271,N_2254);
and U2326 (N_2326,N_2291,N_2288);
nor U2327 (N_2327,N_2262,N_2264);
nor U2328 (N_2328,N_2296,N_2306);
or U2329 (N_2329,N_2285,N_2284);
or U2330 (N_2330,N_2314,N_2268);
or U2331 (N_2331,N_2295,N_2280);
nand U2332 (N_2332,N_2265,N_2282);
or U2333 (N_2333,N_2298,N_2293);
and U2334 (N_2334,N_2260,N_2258);
and U2335 (N_2335,N_2252,N_2257);
nand U2336 (N_2336,N_2310,N_2292);
and U2337 (N_2337,N_2287,N_2319);
and U2338 (N_2338,N_2300,N_2315);
or U2339 (N_2339,N_2277,N_2261);
and U2340 (N_2340,N_2279,N_2308);
and U2341 (N_2341,N_2318,N_2301);
or U2342 (N_2342,N_2272,N_2259);
and U2343 (N_2343,N_2250,N_2304);
or U2344 (N_2344,N_2311,N_2269);
and U2345 (N_2345,N_2297,N_2303);
nor U2346 (N_2346,N_2305,N_2317);
or U2347 (N_2347,N_2255,N_2322);
nand U2348 (N_2348,N_2266,N_2273);
nand U2349 (N_2349,N_2307,N_2299);
and U2350 (N_2350,N_2278,N_2263);
nand U2351 (N_2351,N_2324,N_2286);
or U2352 (N_2352,N_2302,N_2316);
nor U2353 (N_2353,N_2256,N_2275);
nand U2354 (N_2354,N_2294,N_2253);
nand U2355 (N_2355,N_2289,N_2274);
and U2356 (N_2356,N_2320,N_2323);
and U2357 (N_2357,N_2283,N_2281);
nand U2358 (N_2358,N_2276,N_2321);
nand U2359 (N_2359,N_2309,N_2251);
and U2360 (N_2360,N_2312,N_2290);
or U2361 (N_2361,N_2267,N_2313);
or U2362 (N_2362,N_2270,N_2250);
or U2363 (N_2363,N_2299,N_2256);
nand U2364 (N_2364,N_2311,N_2279);
or U2365 (N_2365,N_2302,N_2281);
nand U2366 (N_2366,N_2320,N_2276);
nor U2367 (N_2367,N_2260,N_2280);
nor U2368 (N_2368,N_2250,N_2296);
nor U2369 (N_2369,N_2257,N_2250);
and U2370 (N_2370,N_2318,N_2255);
or U2371 (N_2371,N_2275,N_2269);
nand U2372 (N_2372,N_2290,N_2271);
and U2373 (N_2373,N_2262,N_2266);
or U2374 (N_2374,N_2262,N_2294);
and U2375 (N_2375,N_2290,N_2302);
or U2376 (N_2376,N_2255,N_2292);
nor U2377 (N_2377,N_2291,N_2322);
nor U2378 (N_2378,N_2274,N_2319);
and U2379 (N_2379,N_2296,N_2262);
or U2380 (N_2380,N_2255,N_2279);
nand U2381 (N_2381,N_2287,N_2300);
nor U2382 (N_2382,N_2267,N_2286);
nand U2383 (N_2383,N_2293,N_2311);
or U2384 (N_2384,N_2319,N_2317);
or U2385 (N_2385,N_2275,N_2260);
nand U2386 (N_2386,N_2320,N_2254);
nor U2387 (N_2387,N_2298,N_2272);
or U2388 (N_2388,N_2285,N_2309);
nor U2389 (N_2389,N_2298,N_2294);
nor U2390 (N_2390,N_2286,N_2259);
nor U2391 (N_2391,N_2270,N_2253);
nor U2392 (N_2392,N_2294,N_2272);
and U2393 (N_2393,N_2255,N_2256);
nor U2394 (N_2394,N_2253,N_2299);
or U2395 (N_2395,N_2264,N_2273);
and U2396 (N_2396,N_2320,N_2300);
or U2397 (N_2397,N_2314,N_2297);
nor U2398 (N_2398,N_2313,N_2301);
or U2399 (N_2399,N_2291,N_2324);
nor U2400 (N_2400,N_2338,N_2377);
and U2401 (N_2401,N_2359,N_2392);
or U2402 (N_2402,N_2367,N_2375);
nand U2403 (N_2403,N_2336,N_2364);
nand U2404 (N_2404,N_2357,N_2393);
nand U2405 (N_2405,N_2376,N_2396);
nor U2406 (N_2406,N_2390,N_2334);
nand U2407 (N_2407,N_2387,N_2339);
nor U2408 (N_2408,N_2383,N_2332);
nor U2409 (N_2409,N_2329,N_2354);
nand U2410 (N_2410,N_2347,N_2382);
nand U2411 (N_2411,N_2356,N_2388);
nor U2412 (N_2412,N_2343,N_2379);
and U2413 (N_2413,N_2325,N_2397);
or U2414 (N_2414,N_2361,N_2370);
nor U2415 (N_2415,N_2345,N_2351);
xnor U2416 (N_2416,N_2330,N_2389);
nand U2417 (N_2417,N_2381,N_2378);
nand U2418 (N_2418,N_2386,N_2327);
and U2419 (N_2419,N_2384,N_2337);
or U2420 (N_2420,N_2394,N_2353);
nor U2421 (N_2421,N_2366,N_2398);
nand U2422 (N_2422,N_2348,N_2342);
xor U2423 (N_2423,N_2346,N_2355);
or U2424 (N_2424,N_2380,N_2385);
and U2425 (N_2425,N_2373,N_2352);
or U2426 (N_2426,N_2360,N_2350);
and U2427 (N_2427,N_2368,N_2349);
nor U2428 (N_2428,N_2395,N_2363);
and U2429 (N_2429,N_2358,N_2335);
nor U2430 (N_2430,N_2369,N_2344);
nor U2431 (N_2431,N_2399,N_2340);
nor U2432 (N_2432,N_2331,N_2333);
nand U2433 (N_2433,N_2362,N_2391);
nor U2434 (N_2434,N_2372,N_2341);
or U2435 (N_2435,N_2365,N_2371);
nor U2436 (N_2436,N_2374,N_2326);
and U2437 (N_2437,N_2328,N_2381);
xor U2438 (N_2438,N_2388,N_2389);
and U2439 (N_2439,N_2326,N_2367);
and U2440 (N_2440,N_2384,N_2359);
xor U2441 (N_2441,N_2366,N_2385);
nor U2442 (N_2442,N_2395,N_2399);
nand U2443 (N_2443,N_2354,N_2333);
xor U2444 (N_2444,N_2381,N_2355);
nor U2445 (N_2445,N_2325,N_2394);
nand U2446 (N_2446,N_2339,N_2335);
and U2447 (N_2447,N_2395,N_2341);
nand U2448 (N_2448,N_2352,N_2357);
nand U2449 (N_2449,N_2325,N_2345);
nand U2450 (N_2450,N_2363,N_2340);
nand U2451 (N_2451,N_2392,N_2368);
nand U2452 (N_2452,N_2385,N_2367);
nor U2453 (N_2453,N_2338,N_2345);
nor U2454 (N_2454,N_2397,N_2328);
xnor U2455 (N_2455,N_2385,N_2379);
nor U2456 (N_2456,N_2375,N_2365);
and U2457 (N_2457,N_2393,N_2378);
nor U2458 (N_2458,N_2382,N_2364);
or U2459 (N_2459,N_2365,N_2393);
xor U2460 (N_2460,N_2346,N_2366);
or U2461 (N_2461,N_2333,N_2379);
xor U2462 (N_2462,N_2338,N_2375);
or U2463 (N_2463,N_2344,N_2385);
nand U2464 (N_2464,N_2350,N_2379);
or U2465 (N_2465,N_2397,N_2396);
nor U2466 (N_2466,N_2388,N_2327);
or U2467 (N_2467,N_2346,N_2374);
or U2468 (N_2468,N_2398,N_2329);
nand U2469 (N_2469,N_2362,N_2335);
and U2470 (N_2470,N_2356,N_2334);
and U2471 (N_2471,N_2338,N_2390);
and U2472 (N_2472,N_2333,N_2371);
and U2473 (N_2473,N_2363,N_2327);
or U2474 (N_2474,N_2326,N_2348);
nand U2475 (N_2475,N_2438,N_2439);
and U2476 (N_2476,N_2416,N_2407);
nand U2477 (N_2477,N_2408,N_2430);
or U2478 (N_2478,N_2414,N_2445);
nor U2479 (N_2479,N_2400,N_2453);
and U2480 (N_2480,N_2422,N_2410);
nand U2481 (N_2481,N_2423,N_2468);
nor U2482 (N_2482,N_2434,N_2461);
or U2483 (N_2483,N_2437,N_2465);
and U2484 (N_2484,N_2441,N_2442);
and U2485 (N_2485,N_2421,N_2425);
nand U2486 (N_2486,N_2454,N_2440);
or U2487 (N_2487,N_2449,N_2446);
or U2488 (N_2488,N_2463,N_2470);
nor U2489 (N_2489,N_2472,N_2459);
nor U2490 (N_2490,N_2436,N_2467);
nand U2491 (N_2491,N_2420,N_2415);
and U2492 (N_2492,N_2464,N_2409);
xor U2493 (N_2493,N_2458,N_2462);
or U2494 (N_2494,N_2435,N_2448);
nand U2495 (N_2495,N_2404,N_2431);
or U2496 (N_2496,N_2460,N_2419);
nand U2497 (N_2497,N_2457,N_2403);
nand U2498 (N_2498,N_2426,N_2469);
xor U2499 (N_2499,N_2466,N_2417);
nor U2500 (N_2500,N_2411,N_2432);
nand U2501 (N_2501,N_2451,N_2424);
nor U2502 (N_2502,N_2444,N_2413);
xor U2503 (N_2503,N_2418,N_2456);
and U2504 (N_2504,N_2474,N_2402);
and U2505 (N_2505,N_2401,N_2452);
nor U2506 (N_2506,N_2429,N_2428);
nand U2507 (N_2507,N_2405,N_2471);
nand U2508 (N_2508,N_2433,N_2412);
nor U2509 (N_2509,N_2427,N_2447);
or U2510 (N_2510,N_2473,N_2406);
nor U2511 (N_2511,N_2450,N_2443);
nor U2512 (N_2512,N_2455,N_2428);
nor U2513 (N_2513,N_2448,N_2412);
and U2514 (N_2514,N_2447,N_2402);
or U2515 (N_2515,N_2445,N_2439);
or U2516 (N_2516,N_2454,N_2474);
nand U2517 (N_2517,N_2427,N_2456);
or U2518 (N_2518,N_2432,N_2452);
or U2519 (N_2519,N_2457,N_2434);
and U2520 (N_2520,N_2443,N_2431);
and U2521 (N_2521,N_2417,N_2467);
nor U2522 (N_2522,N_2448,N_2414);
or U2523 (N_2523,N_2436,N_2408);
and U2524 (N_2524,N_2456,N_2423);
nor U2525 (N_2525,N_2442,N_2412);
and U2526 (N_2526,N_2420,N_2403);
nor U2527 (N_2527,N_2431,N_2437);
and U2528 (N_2528,N_2426,N_2461);
nand U2529 (N_2529,N_2430,N_2419);
and U2530 (N_2530,N_2445,N_2449);
or U2531 (N_2531,N_2464,N_2400);
or U2532 (N_2532,N_2432,N_2454);
or U2533 (N_2533,N_2458,N_2463);
or U2534 (N_2534,N_2432,N_2425);
nand U2535 (N_2535,N_2402,N_2462);
nor U2536 (N_2536,N_2451,N_2473);
xor U2537 (N_2537,N_2468,N_2421);
or U2538 (N_2538,N_2411,N_2446);
or U2539 (N_2539,N_2470,N_2425);
and U2540 (N_2540,N_2446,N_2462);
nor U2541 (N_2541,N_2414,N_2446);
nand U2542 (N_2542,N_2443,N_2417);
or U2543 (N_2543,N_2426,N_2401);
nor U2544 (N_2544,N_2424,N_2431);
and U2545 (N_2545,N_2446,N_2422);
and U2546 (N_2546,N_2448,N_2410);
and U2547 (N_2547,N_2469,N_2463);
nand U2548 (N_2548,N_2460,N_2469);
and U2549 (N_2549,N_2444,N_2441);
or U2550 (N_2550,N_2545,N_2511);
nand U2551 (N_2551,N_2515,N_2548);
nor U2552 (N_2552,N_2488,N_2491);
and U2553 (N_2553,N_2534,N_2538);
or U2554 (N_2554,N_2485,N_2547);
or U2555 (N_2555,N_2531,N_2527);
and U2556 (N_2556,N_2528,N_2493);
nand U2557 (N_2557,N_2524,N_2530);
or U2558 (N_2558,N_2475,N_2517);
nor U2559 (N_2559,N_2532,N_2501);
or U2560 (N_2560,N_2502,N_2525);
nand U2561 (N_2561,N_2522,N_2504);
nor U2562 (N_2562,N_2494,N_2498);
nor U2563 (N_2563,N_2549,N_2516);
and U2564 (N_2564,N_2539,N_2481);
nand U2565 (N_2565,N_2542,N_2512);
and U2566 (N_2566,N_2533,N_2500);
nand U2567 (N_2567,N_2489,N_2495);
nor U2568 (N_2568,N_2479,N_2476);
or U2569 (N_2569,N_2518,N_2477);
or U2570 (N_2570,N_2541,N_2507);
and U2571 (N_2571,N_2537,N_2496);
or U2572 (N_2572,N_2513,N_2544);
nor U2573 (N_2573,N_2520,N_2506);
xnor U2574 (N_2574,N_2536,N_2510);
and U2575 (N_2575,N_2514,N_2543);
nor U2576 (N_2576,N_2486,N_2546);
and U2577 (N_2577,N_2480,N_2503);
or U2578 (N_2578,N_2519,N_2482);
nand U2579 (N_2579,N_2521,N_2492);
nor U2580 (N_2580,N_2540,N_2508);
or U2581 (N_2581,N_2499,N_2483);
nor U2582 (N_2582,N_2497,N_2490);
nor U2583 (N_2583,N_2535,N_2484);
or U2584 (N_2584,N_2505,N_2529);
or U2585 (N_2585,N_2487,N_2509);
nand U2586 (N_2586,N_2478,N_2523);
nor U2587 (N_2587,N_2526,N_2506);
nor U2588 (N_2588,N_2537,N_2494);
or U2589 (N_2589,N_2515,N_2479);
and U2590 (N_2590,N_2478,N_2476);
nor U2591 (N_2591,N_2536,N_2521);
nand U2592 (N_2592,N_2541,N_2496);
nor U2593 (N_2593,N_2531,N_2538);
xor U2594 (N_2594,N_2507,N_2515);
nand U2595 (N_2595,N_2513,N_2517);
and U2596 (N_2596,N_2531,N_2483);
nand U2597 (N_2597,N_2497,N_2496);
and U2598 (N_2598,N_2488,N_2521);
or U2599 (N_2599,N_2480,N_2475);
nand U2600 (N_2600,N_2534,N_2483);
or U2601 (N_2601,N_2532,N_2543);
nor U2602 (N_2602,N_2503,N_2547);
or U2603 (N_2603,N_2496,N_2517);
nor U2604 (N_2604,N_2480,N_2537);
and U2605 (N_2605,N_2483,N_2479);
nor U2606 (N_2606,N_2536,N_2534);
and U2607 (N_2607,N_2545,N_2479);
nor U2608 (N_2608,N_2549,N_2522);
nor U2609 (N_2609,N_2500,N_2499);
nand U2610 (N_2610,N_2480,N_2499);
and U2611 (N_2611,N_2524,N_2509);
nand U2612 (N_2612,N_2497,N_2480);
xnor U2613 (N_2613,N_2527,N_2479);
and U2614 (N_2614,N_2519,N_2504);
and U2615 (N_2615,N_2484,N_2539);
or U2616 (N_2616,N_2516,N_2487);
or U2617 (N_2617,N_2516,N_2492);
nor U2618 (N_2618,N_2512,N_2534);
and U2619 (N_2619,N_2481,N_2520);
nand U2620 (N_2620,N_2516,N_2522);
or U2621 (N_2621,N_2510,N_2545);
or U2622 (N_2622,N_2508,N_2481);
and U2623 (N_2623,N_2507,N_2508);
xnor U2624 (N_2624,N_2497,N_2503);
nand U2625 (N_2625,N_2579,N_2618);
xnor U2626 (N_2626,N_2620,N_2597);
or U2627 (N_2627,N_2613,N_2595);
nor U2628 (N_2628,N_2558,N_2616);
nor U2629 (N_2629,N_2615,N_2576);
or U2630 (N_2630,N_2551,N_2607);
nand U2631 (N_2631,N_2568,N_2555);
or U2632 (N_2632,N_2572,N_2567);
nor U2633 (N_2633,N_2574,N_2566);
nor U2634 (N_2634,N_2575,N_2554);
and U2635 (N_2635,N_2577,N_2601);
or U2636 (N_2636,N_2561,N_2622);
nand U2637 (N_2637,N_2614,N_2588);
or U2638 (N_2638,N_2603,N_2617);
nand U2639 (N_2639,N_2593,N_2592);
and U2640 (N_2640,N_2606,N_2599);
nor U2641 (N_2641,N_2594,N_2587);
and U2642 (N_2642,N_2598,N_2557);
nor U2643 (N_2643,N_2583,N_2570);
or U2644 (N_2644,N_2582,N_2610);
and U2645 (N_2645,N_2609,N_2553);
nor U2646 (N_2646,N_2590,N_2578);
nand U2647 (N_2647,N_2621,N_2552);
nor U2648 (N_2648,N_2569,N_2605);
and U2649 (N_2649,N_2608,N_2596);
nor U2650 (N_2650,N_2602,N_2623);
nor U2651 (N_2651,N_2611,N_2580);
nand U2652 (N_2652,N_2562,N_2591);
nor U2653 (N_2653,N_2573,N_2586);
nor U2654 (N_2654,N_2556,N_2581);
or U2655 (N_2655,N_2624,N_2604);
and U2656 (N_2656,N_2585,N_2584);
nand U2657 (N_2657,N_2619,N_2565);
and U2658 (N_2658,N_2571,N_2564);
nand U2659 (N_2659,N_2563,N_2589);
and U2660 (N_2660,N_2600,N_2560);
and U2661 (N_2661,N_2559,N_2550);
nor U2662 (N_2662,N_2612,N_2553);
and U2663 (N_2663,N_2587,N_2606);
nand U2664 (N_2664,N_2608,N_2573);
or U2665 (N_2665,N_2593,N_2557);
or U2666 (N_2666,N_2555,N_2593);
nand U2667 (N_2667,N_2587,N_2619);
or U2668 (N_2668,N_2567,N_2574);
nand U2669 (N_2669,N_2587,N_2577);
or U2670 (N_2670,N_2609,N_2591);
nand U2671 (N_2671,N_2614,N_2560);
nor U2672 (N_2672,N_2617,N_2572);
nand U2673 (N_2673,N_2579,N_2552);
nor U2674 (N_2674,N_2621,N_2559);
nor U2675 (N_2675,N_2585,N_2597);
nand U2676 (N_2676,N_2578,N_2582);
nor U2677 (N_2677,N_2613,N_2576);
and U2678 (N_2678,N_2579,N_2619);
or U2679 (N_2679,N_2601,N_2617);
nand U2680 (N_2680,N_2562,N_2608);
nor U2681 (N_2681,N_2559,N_2599);
or U2682 (N_2682,N_2580,N_2559);
xnor U2683 (N_2683,N_2555,N_2582);
and U2684 (N_2684,N_2592,N_2615);
or U2685 (N_2685,N_2611,N_2573);
and U2686 (N_2686,N_2573,N_2554);
or U2687 (N_2687,N_2573,N_2605);
nand U2688 (N_2688,N_2559,N_2616);
or U2689 (N_2689,N_2607,N_2604);
and U2690 (N_2690,N_2558,N_2587);
and U2691 (N_2691,N_2588,N_2617);
or U2692 (N_2692,N_2581,N_2569);
nor U2693 (N_2693,N_2594,N_2609);
or U2694 (N_2694,N_2608,N_2601);
nand U2695 (N_2695,N_2566,N_2588);
nand U2696 (N_2696,N_2564,N_2568);
nor U2697 (N_2697,N_2610,N_2550);
and U2698 (N_2698,N_2590,N_2601);
or U2699 (N_2699,N_2560,N_2582);
nor U2700 (N_2700,N_2626,N_2680);
nand U2701 (N_2701,N_2662,N_2671);
and U2702 (N_2702,N_2636,N_2633);
or U2703 (N_2703,N_2690,N_2640);
and U2704 (N_2704,N_2639,N_2645);
nand U2705 (N_2705,N_2672,N_2637);
and U2706 (N_2706,N_2656,N_2689);
nand U2707 (N_2707,N_2635,N_2669);
nor U2708 (N_2708,N_2667,N_2697);
or U2709 (N_2709,N_2677,N_2684);
and U2710 (N_2710,N_2679,N_2657);
or U2711 (N_2711,N_2659,N_2681);
or U2712 (N_2712,N_2647,N_2699);
or U2713 (N_2713,N_2638,N_2666);
or U2714 (N_2714,N_2648,N_2695);
and U2715 (N_2715,N_2668,N_2664);
and U2716 (N_2716,N_2650,N_2674);
or U2717 (N_2717,N_2698,N_2642);
and U2718 (N_2718,N_2625,N_2655);
xnor U2719 (N_2719,N_2631,N_2661);
nor U2720 (N_2720,N_2665,N_2660);
and U2721 (N_2721,N_2653,N_2630);
nor U2722 (N_2722,N_2694,N_2627);
or U2723 (N_2723,N_2646,N_2675);
nand U2724 (N_2724,N_2685,N_2651);
and U2725 (N_2725,N_2658,N_2692);
nand U2726 (N_2726,N_2688,N_2634);
nand U2727 (N_2727,N_2643,N_2654);
or U2728 (N_2728,N_2652,N_2628);
and U2729 (N_2729,N_2682,N_2696);
nor U2730 (N_2730,N_2693,N_2644);
and U2731 (N_2731,N_2663,N_2686);
nand U2732 (N_2732,N_2687,N_2649);
and U2733 (N_2733,N_2629,N_2676);
xor U2734 (N_2734,N_2673,N_2632);
or U2735 (N_2735,N_2683,N_2691);
or U2736 (N_2736,N_2641,N_2670);
and U2737 (N_2737,N_2678,N_2682);
xor U2738 (N_2738,N_2636,N_2665);
and U2739 (N_2739,N_2670,N_2668);
nor U2740 (N_2740,N_2674,N_2627);
nor U2741 (N_2741,N_2689,N_2679);
nor U2742 (N_2742,N_2666,N_2692);
nand U2743 (N_2743,N_2684,N_2678);
and U2744 (N_2744,N_2663,N_2676);
or U2745 (N_2745,N_2674,N_2664);
and U2746 (N_2746,N_2651,N_2677);
nand U2747 (N_2747,N_2635,N_2647);
and U2748 (N_2748,N_2651,N_2673);
nor U2749 (N_2749,N_2665,N_2690);
nor U2750 (N_2750,N_2665,N_2633);
nand U2751 (N_2751,N_2664,N_2648);
nor U2752 (N_2752,N_2675,N_2631);
or U2753 (N_2753,N_2661,N_2682);
or U2754 (N_2754,N_2679,N_2626);
and U2755 (N_2755,N_2674,N_2662);
nand U2756 (N_2756,N_2665,N_2685);
nand U2757 (N_2757,N_2685,N_2642);
nor U2758 (N_2758,N_2670,N_2676);
nand U2759 (N_2759,N_2667,N_2647);
nand U2760 (N_2760,N_2675,N_2668);
nand U2761 (N_2761,N_2653,N_2688);
nor U2762 (N_2762,N_2641,N_2674);
or U2763 (N_2763,N_2678,N_2648);
and U2764 (N_2764,N_2686,N_2653);
or U2765 (N_2765,N_2631,N_2638);
or U2766 (N_2766,N_2643,N_2639);
and U2767 (N_2767,N_2644,N_2674);
or U2768 (N_2768,N_2694,N_2698);
nand U2769 (N_2769,N_2684,N_2627);
and U2770 (N_2770,N_2695,N_2659);
nand U2771 (N_2771,N_2651,N_2643);
or U2772 (N_2772,N_2636,N_2627);
xnor U2773 (N_2773,N_2658,N_2684);
and U2774 (N_2774,N_2633,N_2629);
xor U2775 (N_2775,N_2704,N_2742);
nand U2776 (N_2776,N_2715,N_2734);
nor U2777 (N_2777,N_2711,N_2762);
and U2778 (N_2778,N_2706,N_2739);
nand U2779 (N_2779,N_2707,N_2738);
xnor U2780 (N_2780,N_2746,N_2758);
nand U2781 (N_2781,N_2761,N_2732);
or U2782 (N_2782,N_2749,N_2769);
nand U2783 (N_2783,N_2759,N_2753);
or U2784 (N_2784,N_2747,N_2768);
or U2785 (N_2785,N_2720,N_2743);
nor U2786 (N_2786,N_2708,N_2702);
and U2787 (N_2787,N_2773,N_2745);
or U2788 (N_2788,N_2729,N_2719);
nor U2789 (N_2789,N_2752,N_2760);
nor U2790 (N_2790,N_2770,N_2744);
and U2791 (N_2791,N_2748,N_2757);
nor U2792 (N_2792,N_2767,N_2726);
nand U2793 (N_2793,N_2725,N_2733);
and U2794 (N_2794,N_2712,N_2735);
nor U2795 (N_2795,N_2771,N_2703);
or U2796 (N_2796,N_2740,N_2723);
and U2797 (N_2797,N_2730,N_2731);
and U2798 (N_2798,N_2772,N_2721);
nand U2799 (N_2799,N_2700,N_2722);
or U2800 (N_2800,N_2764,N_2736);
nor U2801 (N_2801,N_2705,N_2713);
nor U2802 (N_2802,N_2754,N_2714);
nand U2803 (N_2803,N_2755,N_2774);
xnor U2804 (N_2804,N_2716,N_2727);
and U2805 (N_2805,N_2701,N_2710);
xor U2806 (N_2806,N_2763,N_2750);
or U2807 (N_2807,N_2717,N_2718);
nand U2808 (N_2808,N_2709,N_2724);
and U2809 (N_2809,N_2765,N_2751);
nand U2810 (N_2810,N_2728,N_2737);
and U2811 (N_2811,N_2756,N_2741);
nand U2812 (N_2812,N_2766,N_2713);
and U2813 (N_2813,N_2726,N_2750);
nand U2814 (N_2814,N_2718,N_2764);
or U2815 (N_2815,N_2713,N_2706);
and U2816 (N_2816,N_2745,N_2761);
nand U2817 (N_2817,N_2705,N_2722);
nand U2818 (N_2818,N_2702,N_2763);
nor U2819 (N_2819,N_2717,N_2738);
or U2820 (N_2820,N_2719,N_2728);
or U2821 (N_2821,N_2729,N_2738);
nand U2822 (N_2822,N_2734,N_2736);
nand U2823 (N_2823,N_2770,N_2714);
nor U2824 (N_2824,N_2773,N_2759);
nor U2825 (N_2825,N_2722,N_2749);
or U2826 (N_2826,N_2757,N_2707);
or U2827 (N_2827,N_2763,N_2764);
nor U2828 (N_2828,N_2714,N_2750);
or U2829 (N_2829,N_2767,N_2748);
nand U2830 (N_2830,N_2729,N_2701);
nand U2831 (N_2831,N_2726,N_2764);
and U2832 (N_2832,N_2761,N_2704);
or U2833 (N_2833,N_2753,N_2700);
and U2834 (N_2834,N_2718,N_2714);
nor U2835 (N_2835,N_2709,N_2726);
nor U2836 (N_2836,N_2720,N_2755);
and U2837 (N_2837,N_2764,N_2760);
or U2838 (N_2838,N_2704,N_2770);
nand U2839 (N_2839,N_2709,N_2714);
nand U2840 (N_2840,N_2730,N_2758);
or U2841 (N_2841,N_2745,N_2729);
or U2842 (N_2842,N_2738,N_2747);
and U2843 (N_2843,N_2770,N_2700);
nor U2844 (N_2844,N_2761,N_2727);
nor U2845 (N_2845,N_2738,N_2764);
and U2846 (N_2846,N_2717,N_2711);
nor U2847 (N_2847,N_2752,N_2774);
or U2848 (N_2848,N_2739,N_2765);
and U2849 (N_2849,N_2731,N_2703);
nor U2850 (N_2850,N_2812,N_2813);
and U2851 (N_2851,N_2807,N_2814);
nor U2852 (N_2852,N_2805,N_2788);
nand U2853 (N_2853,N_2775,N_2816);
nor U2854 (N_2854,N_2849,N_2825);
and U2855 (N_2855,N_2784,N_2835);
or U2856 (N_2856,N_2776,N_2804);
and U2857 (N_2857,N_2777,N_2783);
nor U2858 (N_2858,N_2802,N_2789);
and U2859 (N_2859,N_2831,N_2824);
nand U2860 (N_2860,N_2842,N_2799);
nor U2861 (N_2861,N_2815,N_2790);
nor U2862 (N_2862,N_2827,N_2778);
and U2863 (N_2863,N_2846,N_2808);
or U2864 (N_2864,N_2823,N_2798);
and U2865 (N_2865,N_2803,N_2822);
nor U2866 (N_2866,N_2817,N_2793);
nor U2867 (N_2867,N_2832,N_2797);
nor U2868 (N_2868,N_2833,N_2826);
nor U2869 (N_2869,N_2806,N_2834);
or U2870 (N_2870,N_2836,N_2840);
nand U2871 (N_2871,N_2819,N_2818);
xor U2872 (N_2872,N_2786,N_2800);
and U2873 (N_2873,N_2779,N_2794);
nor U2874 (N_2874,N_2844,N_2785);
and U2875 (N_2875,N_2828,N_2810);
nand U2876 (N_2876,N_2829,N_2781);
and U2877 (N_2877,N_2820,N_2841);
or U2878 (N_2878,N_2848,N_2830);
nand U2879 (N_2879,N_2837,N_2782);
and U2880 (N_2880,N_2821,N_2811);
and U2881 (N_2881,N_2838,N_2795);
nand U2882 (N_2882,N_2809,N_2843);
nand U2883 (N_2883,N_2791,N_2839);
nor U2884 (N_2884,N_2787,N_2845);
and U2885 (N_2885,N_2792,N_2847);
and U2886 (N_2886,N_2780,N_2801);
nand U2887 (N_2887,N_2796,N_2789);
or U2888 (N_2888,N_2788,N_2779);
or U2889 (N_2889,N_2796,N_2811);
and U2890 (N_2890,N_2820,N_2778);
nor U2891 (N_2891,N_2827,N_2848);
and U2892 (N_2892,N_2822,N_2790);
xnor U2893 (N_2893,N_2807,N_2779);
nand U2894 (N_2894,N_2806,N_2847);
nand U2895 (N_2895,N_2799,N_2813);
and U2896 (N_2896,N_2833,N_2823);
xnor U2897 (N_2897,N_2798,N_2783);
or U2898 (N_2898,N_2825,N_2816);
nand U2899 (N_2899,N_2802,N_2787);
and U2900 (N_2900,N_2813,N_2839);
or U2901 (N_2901,N_2818,N_2834);
and U2902 (N_2902,N_2840,N_2783);
nor U2903 (N_2903,N_2793,N_2819);
and U2904 (N_2904,N_2824,N_2826);
nand U2905 (N_2905,N_2827,N_2836);
and U2906 (N_2906,N_2831,N_2804);
and U2907 (N_2907,N_2805,N_2804);
nor U2908 (N_2908,N_2818,N_2830);
nor U2909 (N_2909,N_2805,N_2779);
nor U2910 (N_2910,N_2846,N_2814);
xor U2911 (N_2911,N_2838,N_2836);
nor U2912 (N_2912,N_2784,N_2792);
nand U2913 (N_2913,N_2812,N_2779);
nand U2914 (N_2914,N_2792,N_2839);
or U2915 (N_2915,N_2818,N_2789);
nor U2916 (N_2916,N_2828,N_2799);
nor U2917 (N_2917,N_2836,N_2849);
and U2918 (N_2918,N_2783,N_2804);
or U2919 (N_2919,N_2837,N_2775);
xnor U2920 (N_2920,N_2784,N_2779);
and U2921 (N_2921,N_2825,N_2824);
and U2922 (N_2922,N_2776,N_2775);
nor U2923 (N_2923,N_2779,N_2801);
and U2924 (N_2924,N_2796,N_2820);
or U2925 (N_2925,N_2852,N_2920);
or U2926 (N_2926,N_2861,N_2859);
and U2927 (N_2927,N_2885,N_2880);
nor U2928 (N_2928,N_2882,N_2923);
nand U2929 (N_2929,N_2874,N_2899);
nor U2930 (N_2930,N_2879,N_2887);
or U2931 (N_2931,N_2918,N_2877);
nand U2932 (N_2932,N_2906,N_2904);
or U2933 (N_2933,N_2866,N_2868);
or U2934 (N_2934,N_2883,N_2863);
xnor U2935 (N_2935,N_2902,N_2855);
or U2936 (N_2936,N_2858,N_2865);
or U2937 (N_2937,N_2851,N_2854);
nand U2938 (N_2938,N_2875,N_2900);
nor U2939 (N_2939,N_2909,N_2924);
nand U2940 (N_2940,N_2895,N_2893);
or U2941 (N_2941,N_2889,N_2884);
or U2942 (N_2942,N_2891,N_2869);
nand U2943 (N_2943,N_2921,N_2894);
nand U2944 (N_2944,N_2915,N_2901);
nor U2945 (N_2945,N_2917,N_2898);
nor U2946 (N_2946,N_2857,N_2910);
and U2947 (N_2947,N_2916,N_2886);
nor U2948 (N_2948,N_2911,N_2919);
nor U2949 (N_2949,N_2907,N_2878);
and U2950 (N_2950,N_2864,N_2856);
nor U2951 (N_2951,N_2912,N_2873);
nand U2952 (N_2952,N_2871,N_2850);
or U2953 (N_2953,N_2896,N_2905);
nor U2954 (N_2954,N_2853,N_2897);
nor U2955 (N_2955,N_2922,N_2913);
or U2956 (N_2956,N_2872,N_2888);
and U2957 (N_2957,N_2903,N_2860);
or U2958 (N_2958,N_2908,N_2867);
nand U2959 (N_2959,N_2914,N_2881);
and U2960 (N_2960,N_2862,N_2870);
and U2961 (N_2961,N_2890,N_2876);
or U2962 (N_2962,N_2892,N_2869);
nor U2963 (N_2963,N_2902,N_2903);
or U2964 (N_2964,N_2892,N_2901);
nand U2965 (N_2965,N_2911,N_2892);
nor U2966 (N_2966,N_2920,N_2855);
xor U2967 (N_2967,N_2908,N_2886);
or U2968 (N_2968,N_2877,N_2883);
nor U2969 (N_2969,N_2912,N_2876);
nor U2970 (N_2970,N_2872,N_2896);
or U2971 (N_2971,N_2851,N_2887);
nor U2972 (N_2972,N_2918,N_2904);
nand U2973 (N_2973,N_2918,N_2854);
nor U2974 (N_2974,N_2919,N_2850);
nor U2975 (N_2975,N_2914,N_2850);
nand U2976 (N_2976,N_2907,N_2864);
or U2977 (N_2977,N_2903,N_2872);
or U2978 (N_2978,N_2860,N_2917);
and U2979 (N_2979,N_2853,N_2850);
nor U2980 (N_2980,N_2883,N_2902);
and U2981 (N_2981,N_2908,N_2866);
xnor U2982 (N_2982,N_2895,N_2870);
or U2983 (N_2983,N_2911,N_2884);
nand U2984 (N_2984,N_2879,N_2864);
and U2985 (N_2985,N_2913,N_2852);
nand U2986 (N_2986,N_2912,N_2859);
nand U2987 (N_2987,N_2884,N_2878);
and U2988 (N_2988,N_2900,N_2867);
or U2989 (N_2989,N_2865,N_2854);
and U2990 (N_2990,N_2885,N_2911);
or U2991 (N_2991,N_2898,N_2855);
or U2992 (N_2992,N_2878,N_2868);
nor U2993 (N_2993,N_2893,N_2888);
or U2994 (N_2994,N_2898,N_2921);
nand U2995 (N_2995,N_2865,N_2897);
and U2996 (N_2996,N_2907,N_2857);
nor U2997 (N_2997,N_2921,N_2856);
and U2998 (N_2998,N_2850,N_2924);
and U2999 (N_2999,N_2874,N_2892);
nand UO_0 (O_0,N_2968,N_2994);
xor UO_1 (O_1,N_2989,N_2983);
and UO_2 (O_2,N_2980,N_2974);
nand UO_3 (O_3,N_2955,N_2963);
nor UO_4 (O_4,N_2973,N_2965);
or UO_5 (O_5,N_2934,N_2954);
nor UO_6 (O_6,N_2982,N_2930);
nor UO_7 (O_7,N_2950,N_2978);
nor UO_8 (O_8,N_2999,N_2964);
nand UO_9 (O_9,N_2957,N_2969);
and UO_10 (O_10,N_2929,N_2940);
nor UO_11 (O_11,N_2971,N_2967);
or UO_12 (O_12,N_2938,N_2986);
and UO_13 (O_13,N_2952,N_2997);
and UO_14 (O_14,N_2979,N_2949);
or UO_15 (O_15,N_2945,N_2995);
or UO_16 (O_16,N_2946,N_2992);
nor UO_17 (O_17,N_2991,N_2942);
nand UO_18 (O_18,N_2987,N_2961);
or UO_19 (O_19,N_2948,N_2977);
nand UO_20 (O_20,N_2975,N_2993);
nor UO_21 (O_21,N_2990,N_2939);
or UO_22 (O_22,N_2931,N_2981);
or UO_23 (O_23,N_2976,N_2937);
or UO_24 (O_24,N_2972,N_2926);
and UO_25 (O_25,N_2984,N_2932);
nand UO_26 (O_26,N_2925,N_2959);
nor UO_27 (O_27,N_2998,N_2935);
or UO_28 (O_28,N_2951,N_2936);
nor UO_29 (O_29,N_2958,N_2985);
nand UO_30 (O_30,N_2947,N_2966);
and UO_31 (O_31,N_2962,N_2988);
or UO_32 (O_32,N_2933,N_2944);
and UO_33 (O_33,N_2956,N_2928);
and UO_34 (O_34,N_2941,N_2953);
nor UO_35 (O_35,N_2960,N_2996);
or UO_36 (O_36,N_2927,N_2943);
and UO_37 (O_37,N_2970,N_2994);
and UO_38 (O_38,N_2947,N_2965);
or UO_39 (O_39,N_2954,N_2943);
and UO_40 (O_40,N_2935,N_2997);
and UO_41 (O_41,N_2942,N_2943);
and UO_42 (O_42,N_2934,N_2963);
and UO_43 (O_43,N_2990,N_2938);
or UO_44 (O_44,N_2950,N_2955);
and UO_45 (O_45,N_2926,N_2986);
and UO_46 (O_46,N_2938,N_2972);
or UO_47 (O_47,N_2956,N_2979);
and UO_48 (O_48,N_2997,N_2994);
or UO_49 (O_49,N_2928,N_2998);
nand UO_50 (O_50,N_2954,N_2992);
or UO_51 (O_51,N_2939,N_2946);
and UO_52 (O_52,N_2980,N_2983);
nand UO_53 (O_53,N_2968,N_2982);
and UO_54 (O_54,N_2927,N_2958);
nand UO_55 (O_55,N_2994,N_2936);
or UO_56 (O_56,N_2928,N_2970);
nor UO_57 (O_57,N_2963,N_2993);
nand UO_58 (O_58,N_2972,N_2956);
nor UO_59 (O_59,N_2996,N_2938);
or UO_60 (O_60,N_2972,N_2950);
nor UO_61 (O_61,N_2947,N_2963);
or UO_62 (O_62,N_2925,N_2961);
or UO_63 (O_63,N_2931,N_2927);
or UO_64 (O_64,N_2948,N_2985);
nand UO_65 (O_65,N_2952,N_2943);
or UO_66 (O_66,N_2980,N_2984);
or UO_67 (O_67,N_2962,N_2937);
nand UO_68 (O_68,N_2955,N_2964);
or UO_69 (O_69,N_2987,N_2985);
or UO_70 (O_70,N_2938,N_2965);
or UO_71 (O_71,N_2940,N_2982);
or UO_72 (O_72,N_2984,N_2927);
or UO_73 (O_73,N_2985,N_2933);
nand UO_74 (O_74,N_2992,N_2938);
or UO_75 (O_75,N_2951,N_2997);
and UO_76 (O_76,N_2990,N_2980);
nand UO_77 (O_77,N_2932,N_2939);
and UO_78 (O_78,N_2979,N_2964);
nor UO_79 (O_79,N_2994,N_2971);
nor UO_80 (O_80,N_2999,N_2955);
nor UO_81 (O_81,N_2994,N_2965);
and UO_82 (O_82,N_2935,N_2991);
nor UO_83 (O_83,N_2983,N_2959);
nand UO_84 (O_84,N_2968,N_2938);
nor UO_85 (O_85,N_2934,N_2933);
or UO_86 (O_86,N_2974,N_2950);
nand UO_87 (O_87,N_2928,N_2984);
or UO_88 (O_88,N_2995,N_2976);
nor UO_89 (O_89,N_2931,N_2982);
or UO_90 (O_90,N_2984,N_2953);
or UO_91 (O_91,N_2962,N_2956);
or UO_92 (O_92,N_2969,N_2927);
and UO_93 (O_93,N_2949,N_2989);
or UO_94 (O_94,N_2984,N_2961);
and UO_95 (O_95,N_2980,N_2948);
nand UO_96 (O_96,N_2936,N_2990);
nand UO_97 (O_97,N_2985,N_2954);
nor UO_98 (O_98,N_2939,N_2929);
or UO_99 (O_99,N_2996,N_2941);
nor UO_100 (O_100,N_2944,N_2963);
xnor UO_101 (O_101,N_2952,N_2974);
nor UO_102 (O_102,N_2984,N_2930);
or UO_103 (O_103,N_2972,N_2969);
and UO_104 (O_104,N_2958,N_2946);
and UO_105 (O_105,N_2955,N_2994);
nor UO_106 (O_106,N_2984,N_2983);
nand UO_107 (O_107,N_2959,N_2933);
nand UO_108 (O_108,N_2976,N_2941);
nand UO_109 (O_109,N_2952,N_2989);
nor UO_110 (O_110,N_2977,N_2932);
nor UO_111 (O_111,N_2925,N_2940);
or UO_112 (O_112,N_2968,N_2957);
nor UO_113 (O_113,N_2968,N_2927);
and UO_114 (O_114,N_2928,N_2948);
nand UO_115 (O_115,N_2963,N_2949);
or UO_116 (O_116,N_2958,N_2993);
or UO_117 (O_117,N_2987,N_2941);
or UO_118 (O_118,N_2958,N_2929);
nand UO_119 (O_119,N_2970,N_2981);
xor UO_120 (O_120,N_2965,N_2995);
nand UO_121 (O_121,N_2988,N_2963);
or UO_122 (O_122,N_2975,N_2961);
xnor UO_123 (O_123,N_2974,N_2935);
or UO_124 (O_124,N_2937,N_2960);
and UO_125 (O_125,N_2961,N_2964);
and UO_126 (O_126,N_2927,N_2963);
nor UO_127 (O_127,N_2993,N_2959);
xor UO_128 (O_128,N_2963,N_2973);
and UO_129 (O_129,N_2975,N_2996);
nor UO_130 (O_130,N_2972,N_2935);
nor UO_131 (O_131,N_2955,N_2958);
or UO_132 (O_132,N_2964,N_2997);
or UO_133 (O_133,N_2956,N_2952);
or UO_134 (O_134,N_2953,N_2998);
or UO_135 (O_135,N_2990,N_2966);
nor UO_136 (O_136,N_2972,N_2963);
nor UO_137 (O_137,N_2980,N_2959);
and UO_138 (O_138,N_2980,N_2966);
nor UO_139 (O_139,N_2935,N_2976);
nand UO_140 (O_140,N_2960,N_2983);
or UO_141 (O_141,N_2929,N_2938);
or UO_142 (O_142,N_2940,N_2980);
nor UO_143 (O_143,N_2943,N_2975);
and UO_144 (O_144,N_2962,N_2975);
or UO_145 (O_145,N_2947,N_2949);
and UO_146 (O_146,N_2996,N_2951);
or UO_147 (O_147,N_2934,N_2986);
or UO_148 (O_148,N_2943,N_2973);
or UO_149 (O_149,N_2955,N_2962);
or UO_150 (O_150,N_2926,N_2970);
nand UO_151 (O_151,N_2956,N_2932);
or UO_152 (O_152,N_2997,N_2931);
nand UO_153 (O_153,N_2966,N_2965);
nand UO_154 (O_154,N_2958,N_2974);
nor UO_155 (O_155,N_2950,N_2991);
nor UO_156 (O_156,N_2985,N_2960);
or UO_157 (O_157,N_2933,N_2942);
or UO_158 (O_158,N_2976,N_2964);
and UO_159 (O_159,N_2944,N_2948);
nor UO_160 (O_160,N_2934,N_2937);
or UO_161 (O_161,N_2955,N_2995);
or UO_162 (O_162,N_2988,N_2957);
nor UO_163 (O_163,N_2982,N_2983);
or UO_164 (O_164,N_2975,N_2992);
and UO_165 (O_165,N_2990,N_2933);
nor UO_166 (O_166,N_2973,N_2944);
or UO_167 (O_167,N_2968,N_2984);
nand UO_168 (O_168,N_2936,N_2987);
and UO_169 (O_169,N_2934,N_2989);
or UO_170 (O_170,N_2950,N_2967);
nor UO_171 (O_171,N_2951,N_2993);
or UO_172 (O_172,N_2943,N_2960);
or UO_173 (O_173,N_2958,N_2995);
nor UO_174 (O_174,N_2960,N_2984);
or UO_175 (O_175,N_2947,N_2933);
or UO_176 (O_176,N_2960,N_2976);
xor UO_177 (O_177,N_2935,N_2990);
or UO_178 (O_178,N_2943,N_2987);
nor UO_179 (O_179,N_2927,N_2940);
nand UO_180 (O_180,N_2973,N_2983);
nand UO_181 (O_181,N_2976,N_2980);
or UO_182 (O_182,N_2977,N_2981);
or UO_183 (O_183,N_2970,N_2988);
xor UO_184 (O_184,N_2945,N_2929);
nand UO_185 (O_185,N_2965,N_2929);
nand UO_186 (O_186,N_2959,N_2981);
or UO_187 (O_187,N_2943,N_2957);
nor UO_188 (O_188,N_2972,N_2993);
nand UO_189 (O_189,N_2951,N_2937);
nor UO_190 (O_190,N_2998,N_2947);
or UO_191 (O_191,N_2971,N_2960);
nand UO_192 (O_192,N_2991,N_2989);
or UO_193 (O_193,N_2937,N_2931);
xnor UO_194 (O_194,N_2989,N_2959);
nand UO_195 (O_195,N_2955,N_2947);
and UO_196 (O_196,N_2974,N_2954);
nand UO_197 (O_197,N_2960,N_2986);
nand UO_198 (O_198,N_2960,N_2970);
nand UO_199 (O_199,N_2986,N_2971);
xor UO_200 (O_200,N_2943,N_2951);
nand UO_201 (O_201,N_2975,N_2966);
nor UO_202 (O_202,N_2997,N_2992);
and UO_203 (O_203,N_2943,N_2966);
nor UO_204 (O_204,N_2945,N_2956);
nor UO_205 (O_205,N_2927,N_2989);
and UO_206 (O_206,N_2925,N_2934);
nand UO_207 (O_207,N_2936,N_2928);
and UO_208 (O_208,N_2974,N_2994);
and UO_209 (O_209,N_2959,N_2973);
and UO_210 (O_210,N_2942,N_2954);
nand UO_211 (O_211,N_2951,N_2952);
or UO_212 (O_212,N_2946,N_2997);
or UO_213 (O_213,N_2964,N_2960);
or UO_214 (O_214,N_2939,N_2988);
nand UO_215 (O_215,N_2957,N_2966);
nor UO_216 (O_216,N_2926,N_2999);
nor UO_217 (O_217,N_2957,N_2931);
nand UO_218 (O_218,N_2944,N_2956);
nand UO_219 (O_219,N_2942,N_2951);
nand UO_220 (O_220,N_2999,N_2985);
nand UO_221 (O_221,N_2941,N_2966);
nor UO_222 (O_222,N_2968,N_2954);
nand UO_223 (O_223,N_2940,N_2987);
nor UO_224 (O_224,N_2969,N_2933);
nand UO_225 (O_225,N_2992,N_2931);
nor UO_226 (O_226,N_2994,N_2942);
nand UO_227 (O_227,N_2983,N_2966);
nor UO_228 (O_228,N_2951,N_2928);
and UO_229 (O_229,N_2975,N_2933);
nor UO_230 (O_230,N_2998,N_2965);
or UO_231 (O_231,N_2996,N_2962);
nor UO_232 (O_232,N_2976,N_2932);
nor UO_233 (O_233,N_2984,N_2934);
nand UO_234 (O_234,N_2973,N_2931);
or UO_235 (O_235,N_2987,N_2945);
or UO_236 (O_236,N_2942,N_2959);
or UO_237 (O_237,N_2929,N_2987);
or UO_238 (O_238,N_2995,N_2975);
or UO_239 (O_239,N_2946,N_2995);
nand UO_240 (O_240,N_2973,N_2995);
nor UO_241 (O_241,N_2973,N_2961);
nand UO_242 (O_242,N_2940,N_2981);
nor UO_243 (O_243,N_2959,N_2975);
and UO_244 (O_244,N_2972,N_2948);
and UO_245 (O_245,N_2965,N_2979);
nor UO_246 (O_246,N_2981,N_2978);
or UO_247 (O_247,N_2932,N_2971);
nand UO_248 (O_248,N_2953,N_2981);
nand UO_249 (O_249,N_2967,N_2972);
or UO_250 (O_250,N_2986,N_2997);
nand UO_251 (O_251,N_2961,N_2988);
nand UO_252 (O_252,N_2956,N_2954);
nor UO_253 (O_253,N_2975,N_2985);
nand UO_254 (O_254,N_2946,N_2976);
nand UO_255 (O_255,N_2956,N_2997);
or UO_256 (O_256,N_2966,N_2932);
nor UO_257 (O_257,N_2934,N_2950);
nor UO_258 (O_258,N_2952,N_2987);
and UO_259 (O_259,N_2979,N_2954);
nor UO_260 (O_260,N_2987,N_2976);
or UO_261 (O_261,N_2950,N_2977);
and UO_262 (O_262,N_2932,N_2941);
or UO_263 (O_263,N_2970,N_2969);
or UO_264 (O_264,N_2962,N_2938);
nand UO_265 (O_265,N_2954,N_2933);
and UO_266 (O_266,N_2970,N_2983);
and UO_267 (O_267,N_2926,N_2977);
or UO_268 (O_268,N_2982,N_2993);
and UO_269 (O_269,N_2992,N_2974);
or UO_270 (O_270,N_2997,N_2978);
and UO_271 (O_271,N_2942,N_2948);
or UO_272 (O_272,N_2960,N_2962);
nor UO_273 (O_273,N_2990,N_2957);
nand UO_274 (O_274,N_2974,N_2981);
nand UO_275 (O_275,N_2999,N_2973);
or UO_276 (O_276,N_2953,N_2994);
nor UO_277 (O_277,N_2996,N_2963);
nor UO_278 (O_278,N_2970,N_2963);
nand UO_279 (O_279,N_2932,N_2967);
nor UO_280 (O_280,N_2984,N_2933);
or UO_281 (O_281,N_2990,N_2977);
nand UO_282 (O_282,N_2956,N_2947);
nor UO_283 (O_283,N_2972,N_2958);
nor UO_284 (O_284,N_2927,N_2952);
nor UO_285 (O_285,N_2963,N_2999);
and UO_286 (O_286,N_2964,N_2972);
or UO_287 (O_287,N_2942,N_2936);
and UO_288 (O_288,N_2992,N_2957);
or UO_289 (O_289,N_2994,N_2950);
and UO_290 (O_290,N_2986,N_2940);
or UO_291 (O_291,N_2960,N_2968);
or UO_292 (O_292,N_2943,N_2994);
and UO_293 (O_293,N_2997,N_2991);
nand UO_294 (O_294,N_2967,N_2975);
xor UO_295 (O_295,N_2949,N_2935);
and UO_296 (O_296,N_2927,N_2957);
nand UO_297 (O_297,N_2993,N_2950);
and UO_298 (O_298,N_2963,N_2929);
nor UO_299 (O_299,N_2949,N_2969);
nor UO_300 (O_300,N_2992,N_2977);
and UO_301 (O_301,N_2957,N_2993);
nor UO_302 (O_302,N_2972,N_2946);
and UO_303 (O_303,N_2983,N_2957);
or UO_304 (O_304,N_2937,N_2965);
nor UO_305 (O_305,N_2960,N_2988);
nor UO_306 (O_306,N_2977,N_2976);
nand UO_307 (O_307,N_2966,N_2959);
and UO_308 (O_308,N_2930,N_2980);
and UO_309 (O_309,N_2943,N_2981);
and UO_310 (O_310,N_2989,N_2940);
and UO_311 (O_311,N_2944,N_2974);
and UO_312 (O_312,N_2940,N_2961);
nand UO_313 (O_313,N_2925,N_2944);
nor UO_314 (O_314,N_2983,N_2990);
nor UO_315 (O_315,N_2972,N_2996);
nand UO_316 (O_316,N_2972,N_2975);
or UO_317 (O_317,N_2957,N_2929);
nor UO_318 (O_318,N_2969,N_2998);
nor UO_319 (O_319,N_2926,N_2948);
nor UO_320 (O_320,N_2995,N_2951);
or UO_321 (O_321,N_2932,N_2944);
or UO_322 (O_322,N_2981,N_2990);
or UO_323 (O_323,N_2987,N_2995);
nand UO_324 (O_324,N_2951,N_2927);
nor UO_325 (O_325,N_2926,N_2941);
xnor UO_326 (O_326,N_2969,N_2954);
nand UO_327 (O_327,N_2960,N_2929);
nor UO_328 (O_328,N_2948,N_2965);
and UO_329 (O_329,N_2996,N_2945);
and UO_330 (O_330,N_2931,N_2993);
or UO_331 (O_331,N_2986,N_2949);
nand UO_332 (O_332,N_2960,N_2974);
nor UO_333 (O_333,N_2953,N_2938);
or UO_334 (O_334,N_2968,N_2947);
nand UO_335 (O_335,N_2962,N_2989);
nand UO_336 (O_336,N_2935,N_2982);
xnor UO_337 (O_337,N_2999,N_2967);
and UO_338 (O_338,N_2982,N_2976);
nor UO_339 (O_339,N_2955,N_2936);
nor UO_340 (O_340,N_2977,N_2979);
nor UO_341 (O_341,N_2989,N_2972);
and UO_342 (O_342,N_2979,N_2958);
or UO_343 (O_343,N_2970,N_2937);
and UO_344 (O_344,N_2966,N_2981);
nand UO_345 (O_345,N_2983,N_2992);
nand UO_346 (O_346,N_2982,N_2980);
or UO_347 (O_347,N_2965,N_2968);
or UO_348 (O_348,N_2970,N_2965);
or UO_349 (O_349,N_2966,N_2952);
or UO_350 (O_350,N_2953,N_2946);
and UO_351 (O_351,N_2954,N_2982);
and UO_352 (O_352,N_2934,N_2973);
nand UO_353 (O_353,N_2933,N_2950);
nor UO_354 (O_354,N_2938,N_2942);
and UO_355 (O_355,N_2929,N_2969);
and UO_356 (O_356,N_2999,N_2974);
nor UO_357 (O_357,N_2953,N_2951);
and UO_358 (O_358,N_2943,N_2965);
nor UO_359 (O_359,N_2947,N_2986);
nand UO_360 (O_360,N_2941,N_2950);
nor UO_361 (O_361,N_2955,N_2968);
nor UO_362 (O_362,N_2977,N_2984);
and UO_363 (O_363,N_2992,N_2944);
and UO_364 (O_364,N_2949,N_2953);
or UO_365 (O_365,N_2974,N_2971);
nor UO_366 (O_366,N_2941,N_2968);
or UO_367 (O_367,N_2998,N_2929);
and UO_368 (O_368,N_2934,N_2929);
nand UO_369 (O_369,N_2982,N_2986);
or UO_370 (O_370,N_2984,N_2957);
and UO_371 (O_371,N_2945,N_2989);
and UO_372 (O_372,N_2953,N_2929);
or UO_373 (O_373,N_2937,N_2947);
and UO_374 (O_374,N_2938,N_2984);
and UO_375 (O_375,N_2978,N_2931);
and UO_376 (O_376,N_2959,N_2969);
or UO_377 (O_377,N_2998,N_2983);
nor UO_378 (O_378,N_2945,N_2980);
or UO_379 (O_379,N_2964,N_2986);
or UO_380 (O_380,N_2989,N_2971);
nor UO_381 (O_381,N_2992,N_2961);
or UO_382 (O_382,N_2999,N_2933);
and UO_383 (O_383,N_2965,N_2993);
nor UO_384 (O_384,N_2951,N_2990);
xnor UO_385 (O_385,N_2972,N_2925);
or UO_386 (O_386,N_2972,N_2982);
nand UO_387 (O_387,N_2935,N_2932);
nor UO_388 (O_388,N_2941,N_2980);
nor UO_389 (O_389,N_2958,N_2926);
nand UO_390 (O_390,N_2994,N_2978);
or UO_391 (O_391,N_2925,N_2982);
and UO_392 (O_392,N_2959,N_2957);
nor UO_393 (O_393,N_2984,N_2956);
nand UO_394 (O_394,N_2996,N_2986);
nor UO_395 (O_395,N_2963,N_2928);
nand UO_396 (O_396,N_2990,N_2971);
or UO_397 (O_397,N_2931,N_2939);
nor UO_398 (O_398,N_2956,N_2959);
nor UO_399 (O_399,N_2948,N_2956);
nor UO_400 (O_400,N_2972,N_2928);
and UO_401 (O_401,N_2983,N_2995);
nand UO_402 (O_402,N_2974,N_2968);
or UO_403 (O_403,N_2990,N_2969);
and UO_404 (O_404,N_2942,N_2979);
or UO_405 (O_405,N_2961,N_2990);
nand UO_406 (O_406,N_2971,N_2930);
nor UO_407 (O_407,N_2945,N_2972);
or UO_408 (O_408,N_2933,N_2979);
or UO_409 (O_409,N_2981,N_2962);
nor UO_410 (O_410,N_2962,N_2950);
nor UO_411 (O_411,N_2935,N_2942);
nor UO_412 (O_412,N_2945,N_2932);
nor UO_413 (O_413,N_2953,N_2966);
nand UO_414 (O_414,N_2988,N_2965);
or UO_415 (O_415,N_2964,N_2956);
nand UO_416 (O_416,N_2975,N_2999);
and UO_417 (O_417,N_2945,N_2992);
or UO_418 (O_418,N_2976,N_2963);
nor UO_419 (O_419,N_2984,N_2971);
or UO_420 (O_420,N_2935,N_2927);
nand UO_421 (O_421,N_2999,N_2971);
and UO_422 (O_422,N_2989,N_2951);
nor UO_423 (O_423,N_2932,N_2985);
nor UO_424 (O_424,N_2953,N_2934);
and UO_425 (O_425,N_2933,N_2995);
nor UO_426 (O_426,N_2990,N_2931);
and UO_427 (O_427,N_2981,N_2984);
nand UO_428 (O_428,N_2967,N_2977);
or UO_429 (O_429,N_2928,N_2938);
xor UO_430 (O_430,N_2979,N_2971);
or UO_431 (O_431,N_2926,N_2955);
nand UO_432 (O_432,N_2999,N_2944);
xor UO_433 (O_433,N_2996,N_2952);
nand UO_434 (O_434,N_2926,N_2952);
xor UO_435 (O_435,N_2959,N_2944);
or UO_436 (O_436,N_2992,N_2995);
nand UO_437 (O_437,N_2977,N_2958);
nor UO_438 (O_438,N_2940,N_2958);
nor UO_439 (O_439,N_2926,N_2942);
nor UO_440 (O_440,N_2955,N_2976);
nand UO_441 (O_441,N_2949,N_2926);
or UO_442 (O_442,N_2996,N_2932);
nor UO_443 (O_443,N_2994,N_2934);
nor UO_444 (O_444,N_2987,N_2999);
and UO_445 (O_445,N_2935,N_2926);
and UO_446 (O_446,N_2955,N_2986);
nor UO_447 (O_447,N_2932,N_2940);
or UO_448 (O_448,N_2963,N_2936);
and UO_449 (O_449,N_2996,N_2939);
or UO_450 (O_450,N_2947,N_2989);
or UO_451 (O_451,N_2973,N_2962);
or UO_452 (O_452,N_2976,N_2975);
nand UO_453 (O_453,N_2968,N_2986);
or UO_454 (O_454,N_2992,N_2986);
nand UO_455 (O_455,N_2960,N_2980);
nor UO_456 (O_456,N_2988,N_2956);
nor UO_457 (O_457,N_2950,N_2939);
nand UO_458 (O_458,N_2932,N_2938);
or UO_459 (O_459,N_2980,N_2925);
or UO_460 (O_460,N_2983,N_2987);
nor UO_461 (O_461,N_2978,N_2925);
nand UO_462 (O_462,N_2960,N_2994);
or UO_463 (O_463,N_2968,N_2979);
nand UO_464 (O_464,N_2925,N_2931);
or UO_465 (O_465,N_2980,N_2986);
or UO_466 (O_466,N_2972,N_2973);
nand UO_467 (O_467,N_2946,N_2977);
nor UO_468 (O_468,N_2985,N_2996);
nand UO_469 (O_469,N_2986,N_2933);
nor UO_470 (O_470,N_2946,N_2984);
or UO_471 (O_471,N_2942,N_2955);
or UO_472 (O_472,N_2943,N_2979);
nand UO_473 (O_473,N_2977,N_2944);
and UO_474 (O_474,N_2962,N_2944);
nand UO_475 (O_475,N_2998,N_2925);
or UO_476 (O_476,N_2933,N_2926);
and UO_477 (O_477,N_2986,N_2967);
nand UO_478 (O_478,N_2961,N_2974);
nor UO_479 (O_479,N_2965,N_2928);
nor UO_480 (O_480,N_2967,N_2958);
nand UO_481 (O_481,N_2998,N_2942);
or UO_482 (O_482,N_2945,N_2991);
nand UO_483 (O_483,N_2943,N_2986);
or UO_484 (O_484,N_2988,N_2969);
nor UO_485 (O_485,N_2959,N_2977);
nor UO_486 (O_486,N_2933,N_2939);
nand UO_487 (O_487,N_2958,N_2968);
nor UO_488 (O_488,N_2988,N_2995);
nand UO_489 (O_489,N_2978,N_2951);
nor UO_490 (O_490,N_2929,N_2997);
nand UO_491 (O_491,N_2983,N_2941);
nand UO_492 (O_492,N_2932,N_2959);
nor UO_493 (O_493,N_2960,N_2947);
and UO_494 (O_494,N_2975,N_2930);
and UO_495 (O_495,N_2968,N_2937);
xnor UO_496 (O_496,N_2951,N_2972);
nand UO_497 (O_497,N_2977,N_2975);
nor UO_498 (O_498,N_2933,N_2972);
nor UO_499 (O_499,N_2964,N_2952);
endmodule