module basic_2000_20000_2500_4_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_344,In_379);
or U1 (N_1,In_517,In_1491);
and U2 (N_2,In_1554,In_571);
and U3 (N_3,In_194,In_1038);
and U4 (N_4,In_1634,In_1211);
nor U5 (N_5,In_1661,In_534);
nor U6 (N_6,In_1452,In_353);
nor U7 (N_7,In_953,In_1985);
and U8 (N_8,In_1997,In_1378);
xor U9 (N_9,In_1563,In_1672);
and U10 (N_10,In_1463,In_1006);
nor U11 (N_11,In_444,In_1181);
or U12 (N_12,In_1896,In_515);
xor U13 (N_13,In_640,In_36);
and U14 (N_14,In_1060,In_325);
xnor U15 (N_15,In_203,In_51);
and U16 (N_16,In_1961,In_1890);
nand U17 (N_17,In_18,In_700);
nand U18 (N_18,In_28,In_113);
and U19 (N_19,In_1779,In_8);
xnor U20 (N_20,In_1504,In_1995);
xor U21 (N_21,In_1965,In_1875);
nand U22 (N_22,In_1657,In_234);
nand U23 (N_23,In_1507,In_1146);
xnor U24 (N_24,In_1171,In_1560);
xnor U25 (N_25,In_797,In_24);
nand U26 (N_26,In_306,In_1544);
nand U27 (N_27,In_839,In_982);
xor U28 (N_28,In_473,In_1041);
nand U29 (N_29,In_259,In_462);
xnor U30 (N_30,In_1723,In_507);
and U31 (N_31,In_367,In_693);
nand U32 (N_32,In_1738,In_1577);
or U33 (N_33,In_209,In_1854);
and U34 (N_34,In_314,In_532);
or U35 (N_35,In_723,In_1673);
nor U36 (N_36,In_1832,In_315);
and U37 (N_37,In_552,In_1740);
or U38 (N_38,In_468,In_1201);
nand U39 (N_39,In_1527,In_1443);
nor U40 (N_40,In_1339,In_584);
nor U41 (N_41,In_1770,In_498);
nor U42 (N_42,In_1594,In_172);
xor U43 (N_43,In_124,In_1864);
xnor U44 (N_44,In_660,In_795);
and U45 (N_45,In_66,In_9);
xor U46 (N_46,In_486,In_1616);
or U47 (N_47,In_1222,In_1926);
nand U48 (N_48,In_728,In_1163);
and U49 (N_49,In_558,In_760);
or U50 (N_50,In_493,In_1731);
nand U51 (N_51,In_1477,In_228);
nand U52 (N_52,In_322,In_280);
and U53 (N_53,In_1863,In_218);
nor U54 (N_54,In_1903,In_1621);
nor U55 (N_55,In_765,In_1596);
nand U56 (N_56,In_451,In_1785);
nor U57 (N_57,In_1910,In_1606);
or U58 (N_58,In_427,In_26);
or U59 (N_59,In_1153,In_914);
nand U60 (N_60,In_964,In_1343);
xor U61 (N_61,In_184,In_852);
xor U62 (N_62,In_1633,In_505);
and U63 (N_63,In_1808,In_1022);
nor U64 (N_64,In_186,In_104);
nor U65 (N_65,In_230,In_565);
nand U66 (N_66,In_499,In_60);
nor U67 (N_67,In_1001,In_526);
and U68 (N_68,In_417,In_1963);
nand U69 (N_69,In_1775,In_93);
nor U70 (N_70,In_1458,In_889);
xor U71 (N_71,In_1059,In_118);
nor U72 (N_72,In_1879,In_1704);
or U73 (N_73,In_508,In_727);
nor U74 (N_74,In_879,In_549);
nor U75 (N_75,In_271,In_1356);
xor U76 (N_76,In_443,In_1278);
nor U77 (N_77,In_997,In_207);
nand U78 (N_78,In_109,In_869);
and U79 (N_79,In_1351,In_692);
or U80 (N_80,In_826,In_1043);
nor U81 (N_81,In_1391,In_158);
or U82 (N_82,In_1329,In_1856);
xnor U83 (N_83,In_1318,In_1630);
nand U84 (N_84,In_1931,In_1649);
and U85 (N_85,In_22,In_452);
nand U86 (N_86,In_89,In_17);
xor U87 (N_87,In_1906,In_685);
nand U88 (N_88,In_1110,In_1818);
and U89 (N_89,In_431,In_1459);
nand U90 (N_90,In_1279,In_482);
xor U91 (N_91,In_1091,In_1521);
nor U92 (N_92,In_1551,In_540);
or U93 (N_93,In_350,In_1710);
xor U94 (N_94,In_543,In_33);
nor U95 (N_95,In_1380,In_650);
nand U96 (N_96,In_136,In_1972);
and U97 (N_97,In_198,In_530);
or U98 (N_98,In_433,In_430);
nor U99 (N_99,In_1344,In_531);
xor U100 (N_100,In_324,In_423);
and U101 (N_101,In_1795,In_457);
nor U102 (N_102,In_1207,In_1976);
xnor U103 (N_103,In_305,In_667);
nand U104 (N_104,In_1028,In_1703);
and U105 (N_105,In_143,In_1450);
or U106 (N_106,In_616,In_695);
xor U107 (N_107,In_291,In_607);
or U108 (N_108,In_1453,In_1801);
or U109 (N_109,In_787,In_1117);
nand U110 (N_110,In_1918,In_1120);
and U111 (N_111,In_1601,In_1750);
and U112 (N_112,In_1708,In_1752);
nor U113 (N_113,In_436,In_72);
or U114 (N_114,In_1062,In_1923);
and U115 (N_115,In_1759,In_863);
nand U116 (N_116,In_276,In_1907);
and U117 (N_117,In_1855,In_220);
nor U118 (N_118,In_597,In_1846);
nor U119 (N_119,In_822,In_55);
nor U120 (N_120,In_1636,In_45);
nand U121 (N_121,In_166,In_311);
or U122 (N_122,In_1324,In_173);
and U123 (N_123,In_402,In_994);
nor U124 (N_124,In_1472,In_422);
and U125 (N_125,In_1783,In_1193);
nand U126 (N_126,In_469,In_358);
nand U127 (N_127,In_1036,In_490);
and U128 (N_128,In_320,In_1604);
and U129 (N_129,In_838,In_187);
nand U130 (N_130,In_1233,In_57);
nand U131 (N_131,In_546,In_1614);
and U132 (N_132,In_1899,In_248);
or U133 (N_133,In_1575,In_1248);
and U134 (N_134,In_1009,In_1470);
nor U135 (N_135,In_843,In_545);
or U136 (N_136,In_649,In_1953);
and U137 (N_137,In_1049,In_1056);
nand U138 (N_138,In_1415,In_1363);
and U139 (N_139,In_848,In_1786);
or U140 (N_140,In_567,In_1608);
or U141 (N_141,In_1300,In_290);
nor U142 (N_142,In_894,In_991);
or U143 (N_143,In_471,In_1951);
or U144 (N_144,In_524,In_909);
nor U145 (N_145,In_1115,In_1489);
nand U146 (N_146,In_939,In_1578);
nand U147 (N_147,In_195,In_1622);
nor U148 (N_148,In_1700,In_1683);
or U149 (N_149,In_1736,In_1256);
or U150 (N_150,In_731,In_213);
nor U151 (N_151,In_757,In_1400);
xor U152 (N_152,In_284,In_824);
nand U153 (N_153,In_1381,In_1707);
or U154 (N_154,In_1940,In_794);
nor U155 (N_155,In_1265,In_537);
xor U156 (N_156,In_1958,In_956);
nand U157 (N_157,In_1087,In_818);
or U158 (N_158,In_385,In_1188);
nor U159 (N_159,In_1333,In_1372);
or U160 (N_160,In_1493,In_192);
xnor U161 (N_161,In_1959,In_438);
and U162 (N_162,In_999,In_1682);
and U163 (N_163,In_935,In_340);
xnor U164 (N_164,In_1526,In_1600);
xnor U165 (N_165,In_189,In_758);
xnor U166 (N_166,In_1629,In_42);
nor U167 (N_167,In_608,In_352);
nand U168 (N_168,In_1639,In_535);
nor U169 (N_169,In_122,In_244);
xnor U170 (N_170,In_1199,In_153);
nor U171 (N_171,In_478,In_1019);
nand U172 (N_172,In_1418,In_132);
nor U173 (N_173,In_1177,In_197);
or U174 (N_174,In_674,In_83);
nand U175 (N_175,In_16,In_150);
xnor U176 (N_176,In_593,In_1154);
xor U177 (N_177,In_1838,In_1015);
nor U178 (N_178,In_1642,In_1371);
nand U179 (N_179,In_958,In_1756);
xnor U180 (N_180,In_561,In_729);
nor U181 (N_181,In_529,In_1425);
nor U182 (N_182,In_405,In_1238);
xor U183 (N_183,In_1320,In_1861);
and U184 (N_184,In_1688,In_116);
nand U185 (N_185,In_972,In_1132);
or U186 (N_186,In_1667,In_1429);
and U187 (N_187,In_1652,In_1074);
xor U188 (N_188,In_1294,In_1486);
and U189 (N_189,In_772,In_873);
or U190 (N_190,In_1155,In_544);
xnor U191 (N_191,In_210,In_1495);
or U192 (N_192,In_1757,In_1474);
or U193 (N_193,In_1658,In_1338);
or U194 (N_194,In_559,In_1749);
and U195 (N_195,In_790,In_653);
nor U196 (N_196,In_1471,In_1617);
nand U197 (N_197,In_955,In_1139);
and U198 (N_198,In_1308,In_390);
nor U199 (N_199,In_1124,In_1929);
xor U200 (N_200,In_1763,In_399);
xnor U201 (N_201,In_580,In_1190);
xnor U202 (N_202,In_809,In_1319);
nand U203 (N_203,In_1887,In_1274);
or U204 (N_204,In_648,In_27);
or U205 (N_205,In_1141,In_882);
and U206 (N_206,In_382,In_872);
or U207 (N_207,In_933,In_1802);
or U208 (N_208,In_348,In_121);
nor U209 (N_209,In_77,In_1911);
nand U210 (N_210,In_159,In_715);
nor U211 (N_211,In_1295,In_1179);
and U212 (N_212,In_1455,In_208);
nand U213 (N_213,In_1533,In_1721);
or U214 (N_214,In_1107,In_627);
nand U215 (N_215,In_1395,In_1747);
nand U216 (N_216,In_1946,In_1771);
nor U217 (N_217,In_1924,In_1392);
and U218 (N_218,In_298,In_883);
xor U219 (N_219,In_392,In_1241);
and U220 (N_220,In_823,In_878);
and U221 (N_221,In_375,In_1514);
or U222 (N_222,In_1925,In_988);
and U223 (N_223,In_181,In_223);
nor U224 (N_224,In_226,In_1086);
nor U225 (N_225,In_316,In_68);
xor U226 (N_226,In_447,In_412);
nand U227 (N_227,In_1886,In_1151);
nand U228 (N_228,In_1938,In_400);
and U229 (N_229,In_1824,In_1748);
nor U230 (N_230,In_1003,In_1511);
nor U231 (N_231,In_1244,In_773);
nand U232 (N_232,In_1535,In_48);
nor U233 (N_233,In_217,In_1121);
nand U234 (N_234,In_1161,In_1917);
or U235 (N_235,In_1335,In_762);
nand U236 (N_236,In_1494,In_1605);
nor U237 (N_237,In_286,In_1768);
or U238 (N_238,In_1585,In_793);
and U239 (N_239,In_71,In_485);
nor U240 (N_240,In_1525,In_455);
or U241 (N_241,In_1449,In_450);
or U242 (N_242,In_600,In_588);
and U243 (N_243,In_1815,In_0);
nand U244 (N_244,In_65,In_295);
nor U245 (N_245,In_1446,In_174);
xor U246 (N_246,In_1084,In_1964);
nor U247 (N_247,In_896,In_190);
nand U248 (N_248,In_1203,In_893);
nand U249 (N_249,In_706,In_1385);
nand U250 (N_250,In_59,In_233);
nor U251 (N_251,In_1692,In_1522);
nor U252 (N_252,In_1532,In_906);
nor U253 (N_253,In_1826,In_514);
and U254 (N_254,In_691,In_1568);
nand U255 (N_255,In_1461,In_100);
xnor U256 (N_256,In_1714,In_764);
and U257 (N_257,In_1042,In_969);
nand U258 (N_258,In_928,In_1993);
nand U259 (N_259,In_200,In_771);
xnor U260 (N_260,In_1099,In_1322);
nor U261 (N_261,In_458,In_1373);
and U262 (N_262,In_978,In_502);
and U263 (N_263,In_349,In_1696);
nand U264 (N_264,In_576,In_1083);
nand U265 (N_265,In_522,In_135);
xnor U266 (N_266,In_1383,In_1464);
or U267 (N_267,In_657,In_888);
and U268 (N_268,In_1957,In_1569);
xor U269 (N_269,In_837,In_779);
and U270 (N_270,In_364,In_743);
and U271 (N_271,In_983,In_215);
nand U272 (N_272,In_1726,In_2);
and U273 (N_273,In_652,In_819);
or U274 (N_274,In_374,In_1541);
and U275 (N_275,In_751,In_221);
nor U276 (N_276,In_1590,In_81);
nor U277 (N_277,In_1989,In_191);
and U278 (N_278,In_901,In_239);
nor U279 (N_279,In_841,In_719);
xnor U280 (N_280,In_1109,In_989);
nor U281 (N_281,In_912,In_354);
xor U282 (N_282,In_176,In_96);
nor U283 (N_283,In_708,In_753);
or U284 (N_284,In_1366,In_618);
nand U285 (N_285,In_911,In_378);
nand U286 (N_286,In_635,In_1516);
nand U287 (N_287,In_175,In_636);
nand U288 (N_288,In_1837,In_767);
nand U289 (N_289,In_668,In_1340);
xnor U290 (N_290,In_730,In_1209);
and U291 (N_291,In_256,In_1691);
and U292 (N_292,In_1979,In_363);
nor U293 (N_293,In_536,In_247);
nor U294 (N_294,In_97,In_1873);
nand U295 (N_295,In_1481,In_1693);
nor U296 (N_296,In_1921,In_1646);
xor U297 (N_297,In_756,In_1537);
xnor U298 (N_298,In_830,In_1713);
and U299 (N_299,In_1588,In_1390);
or U300 (N_300,In_1874,In_397);
and U301 (N_301,In_371,In_249);
nor U302 (N_302,In_778,In_1687);
xnor U303 (N_303,In_661,In_1719);
xor U304 (N_304,In_602,In_1160);
or U305 (N_305,In_1114,In_579);
nor U306 (N_306,In_1206,In_1102);
xor U307 (N_307,In_881,In_643);
nor U308 (N_308,In_804,In_1576);
or U309 (N_309,In_644,In_1579);
xor U310 (N_310,In_798,In_1014);
nor U311 (N_311,In_1296,In_995);
nor U312 (N_312,In_1411,In_235);
nand U313 (N_313,In_973,In_1310);
nand U314 (N_314,In_1572,In_44);
xnor U315 (N_315,In_1029,In_114);
or U316 (N_316,In_1829,In_961);
and U317 (N_317,In_1974,In_811);
or U318 (N_318,In_533,In_1305);
nor U319 (N_319,In_1349,In_3);
xnor U320 (N_320,In_1973,In_735);
or U321 (N_321,In_1169,In_1242);
or U322 (N_322,In_1651,In_1182);
nor U323 (N_323,In_733,In_1334);
nor U324 (N_324,In_624,In_1187);
xnor U325 (N_325,In_1799,In_717);
nand U326 (N_326,In_713,In_711);
or U327 (N_327,In_870,In_698);
or U328 (N_328,In_741,In_1135);
xnor U329 (N_329,In_1675,In_1625);
and U330 (N_330,In_1166,In_1094);
xnor U331 (N_331,In_1035,In_461);
xor U332 (N_332,In_1851,In_853);
nand U333 (N_333,In_1312,In_1325);
and U334 (N_334,In_1467,In_555);
nand U335 (N_335,In_931,In_918);
and U336 (N_336,In_628,In_1186);
and U337 (N_337,In_1880,In_321);
and U338 (N_338,In_501,In_130);
or U339 (N_339,In_394,In_747);
and U340 (N_340,In_1655,In_1663);
xor U341 (N_341,In_1313,In_877);
or U342 (N_342,In_1638,In_716);
xor U343 (N_343,In_1210,In_1828);
xor U344 (N_344,In_547,In_460);
and U345 (N_345,In_777,In_409);
nand U346 (N_346,In_871,In_1914);
xnor U347 (N_347,In_1599,In_1108);
and U348 (N_348,In_1219,In_222);
xor U349 (N_349,In_1417,In_1662);
and U350 (N_350,In_554,In_37);
nor U351 (N_351,In_1133,In_1192);
nand U352 (N_352,In_1399,In_898);
and U353 (N_353,In_370,In_1058);
nand U354 (N_354,In_921,In_376);
and U355 (N_355,In_278,In_1547);
xor U356 (N_356,In_1165,In_246);
nand U357 (N_357,In_1555,In_1127);
nand U358 (N_358,In_1023,In_1232);
or U359 (N_359,In_265,In_1212);
xor U360 (N_360,In_1326,In_539);
or U361 (N_361,In_996,In_915);
and U362 (N_362,In_404,In_488);
nor U363 (N_363,In_970,In_313);
nor U364 (N_364,In_125,In_832);
nor U365 (N_365,In_1040,In_516);
nand U366 (N_366,In_1462,In_86);
xnor U367 (N_367,In_850,In_411);
or U368 (N_368,In_211,In_151);
xor U369 (N_369,In_569,In_67);
nor U370 (N_370,In_710,In_1321);
xnor U371 (N_371,In_1438,In_1791);
or U372 (N_372,In_1044,In_846);
nor U373 (N_373,In_1552,In_1531);
nor U374 (N_374,In_1881,In_476);
nor U375 (N_375,In_1172,In_1309);
and U376 (N_376,In_19,In_445);
nand U377 (N_377,In_979,In_1920);
nand U378 (N_378,In_936,In_1919);
or U379 (N_379,In_631,In_948);
xor U380 (N_380,In_73,In_860);
or U381 (N_381,In_858,In_307);
and U382 (N_382,In_1792,In_336);
nand U383 (N_383,In_254,In_876);
nand U384 (N_384,In_1364,In_1517);
nand U385 (N_385,In_601,In_1408);
and U386 (N_386,In_1612,In_1705);
nand U387 (N_387,In_1912,In_1235);
and U388 (N_388,In_967,In_784);
or U389 (N_389,In_1697,In_959);
and U390 (N_390,In_1530,In_1559);
and U391 (N_391,In_1229,In_1025);
and U392 (N_392,In_312,In_1966);
xor U393 (N_393,In_416,In_1934);
xnor U394 (N_394,In_1287,In_1353);
xnor U395 (N_395,In_775,In_1034);
nor U396 (N_396,In_329,In_160);
nand U397 (N_397,In_1159,In_563);
and U398 (N_398,In_694,In_1039);
or U399 (N_399,In_1031,In_1227);
and U400 (N_400,In_1419,In_857);
xnor U401 (N_401,In_383,In_1285);
nand U402 (N_402,In_429,In_157);
nor U403 (N_403,In_261,In_1370);
nand U404 (N_404,In_1830,In_1476);
or U405 (N_405,In_806,In_739);
or U406 (N_406,In_296,In_1016);
nand U407 (N_407,In_1093,In_229);
and U408 (N_408,In_1473,In_1510);
and U409 (N_409,In_489,In_866);
nand U410 (N_410,In_1358,In_29);
xnor U411 (N_411,In_769,In_895);
xor U412 (N_412,In_268,In_1080);
and U413 (N_413,In_509,In_833);
and U414 (N_414,In_1998,In_677);
or U415 (N_415,In_1977,In_1733);
xor U416 (N_416,In_1478,In_1860);
or U417 (N_417,In_1928,In_709);
and U418 (N_418,In_842,In_987);
xnor U419 (N_419,In_52,In_908);
or U420 (N_420,In_162,In_74);
xnor U421 (N_421,In_323,In_591);
or U422 (N_422,In_1156,In_1746);
and U423 (N_423,In_1147,In_557);
or U424 (N_424,In_212,In_1125);
and U425 (N_425,In_1051,In_1627);
nor U426 (N_426,In_1788,In_1077);
nand U427 (N_427,In_389,In_1480);
nor U428 (N_428,In_224,In_718);
or U429 (N_429,In_1566,In_1286);
nand U430 (N_430,In_984,In_1952);
and U431 (N_431,In_1050,In_1345);
xor U432 (N_432,In_855,In_171);
or U433 (N_433,In_974,In_1072);
or U434 (N_434,In_1488,In_1061);
and U435 (N_435,In_1986,In_107);
nor U436 (N_436,In_1412,In_282);
or U437 (N_437,In_905,In_85);
or U438 (N_438,In_1943,In_1048);
and U439 (N_439,In_1987,In_1778);
nand U440 (N_440,In_1447,In_408);
or U441 (N_441,In_251,In_1571);
and U442 (N_442,In_814,In_1812);
xnor U443 (N_443,In_1005,In_696);
xor U444 (N_444,In_1076,In_164);
or U445 (N_445,In_69,In_1755);
and U446 (N_446,In_1671,In_614);
nor U447 (N_447,In_1439,In_670);
xor U448 (N_448,In_1969,In_886);
and U449 (N_449,In_41,In_847);
nor U450 (N_450,In_820,In_1362);
nand U451 (N_451,In_1445,In_1346);
xnor U452 (N_452,In_523,In_1002);
and U453 (N_453,In_237,In_862);
xor U454 (N_454,In_623,In_1119);
and U455 (N_455,In_464,In_289);
and U456 (N_456,In_892,In_672);
and U457 (N_457,In_138,In_1955);
nor U458 (N_458,In_1883,In_1970);
or U459 (N_459,In_477,In_334);
nor U460 (N_460,In_799,In_599);
nand U461 (N_461,In_1654,In_1845);
nand U462 (N_462,In_1950,In_1674);
nor U463 (N_463,In_446,In_87);
xnor U464 (N_464,In_1690,In_1584);
nand U465 (N_465,In_1536,In_518);
and U466 (N_466,In_1089,In_1609);
or U467 (N_467,In_1469,In_1456);
or U468 (N_468,In_35,In_317);
nand U469 (N_469,In_594,In_586);
and U470 (N_470,In_10,In_232);
and U471 (N_471,In_1574,In_1484);
nor U472 (N_472,In_1303,In_551);
nand U473 (N_473,In_737,In_475);
xor U474 (N_474,In_725,In_494);
and U475 (N_475,In_1680,In_834);
nand U476 (N_476,In_1284,In_1954);
and U477 (N_477,In_46,In_1404);
nor U478 (N_478,In_1431,In_1784);
xnor U479 (N_479,In_926,In_1999);
nor U480 (N_480,In_1460,In_550);
nor U481 (N_481,In_1433,In_142);
or U482 (N_482,In_418,In_345);
nor U483 (N_483,In_1067,In_407);
and U484 (N_484,In_658,In_528);
nand U485 (N_485,In_112,In_196);
nor U486 (N_486,In_5,In_1720);
or U487 (N_487,In_53,In_262);
nor U488 (N_488,In_467,In_605);
and U489 (N_489,In_1937,In_1162);
and U490 (N_490,In_1129,In_39);
nand U491 (N_491,In_1111,In_117);
xnor U492 (N_492,In_1401,In_582);
or U493 (N_493,In_742,In_632);
xor U494 (N_494,In_1564,In_442);
nand U495 (N_495,In_1501,In_342);
nor U496 (N_496,In_1503,In_637);
and U497 (N_497,In_1718,In_1289);
and U498 (N_498,In_1116,In_496);
xor U499 (N_499,In_459,In_1342);
and U500 (N_500,In_1293,In_856);
or U501 (N_501,In_788,In_681);
or U502 (N_502,In_625,In_58);
nand U503 (N_503,In_1138,In_219);
and U504 (N_504,In_1913,In_1732);
nor U505 (N_505,In_14,In_1558);
nor U506 (N_506,In_1157,In_1500);
nand U507 (N_507,In_1465,In_101);
or U508 (N_508,In_639,In_990);
and U509 (N_509,In_365,In_1306);
nand U510 (N_510,In_1774,In_1075);
and U511 (N_511,In_1332,In_1698);
or U512 (N_512,In_663,In_272);
nor U513 (N_513,In_553,In_170);
nor U514 (N_514,In_675,In_183);
xnor U515 (N_515,In_500,In_252);
nor U516 (N_516,In_1430,In_568);
or U517 (N_517,In_439,In_6);
nor U518 (N_518,In_1766,In_351);
nand U519 (N_519,In_1299,In_992);
nand U520 (N_520,In_527,In_1376);
and U521 (N_521,In_236,In_815);
nor U522 (N_522,In_1214,In_812);
nor U523 (N_523,In_1336,In_1282);
or U524 (N_524,In_264,In_1377);
xor U525 (N_525,In_1597,In_746);
and U526 (N_526,In_891,In_574);
nand U527 (N_527,In_770,In_1368);
or U528 (N_528,In_1947,In_1355);
nor U529 (N_529,In_1737,In_90);
nor U530 (N_530,In_620,In_1348);
nand U531 (N_531,In_904,In_642);
nand U532 (N_532,In_238,In_1106);
and U533 (N_533,In_1991,In_851);
xor U534 (N_534,In_1100,In_1835);
xor U535 (N_535,In_139,In_1055);
and U536 (N_536,In_373,In_705);
nand U537 (N_537,In_214,In_1839);
nand U538 (N_538,In_106,In_1528);
and U539 (N_539,In_1267,In_589);
xnor U540 (N_540,In_1302,In_1317);
nor U541 (N_541,In_369,In_1103);
xnor U542 (N_542,In_1885,In_310);
or U543 (N_543,In_1857,In_1379);
nand U544 (N_544,In_1648,In_1670);
nand U545 (N_545,In_1787,In_1717);
nand U546 (N_546,In_1226,In_301);
or U547 (N_547,In_1085,In_566);
xor U548 (N_548,In_168,In_748);
nor U549 (N_549,In_1772,In_401);
or U550 (N_550,In_1168,In_99);
nand U551 (N_551,In_1158,In_1669);
xor U552 (N_552,In_1330,In_319);
and U553 (N_553,In_581,In_656);
and U554 (N_554,In_1653,In_917);
xor U555 (N_555,In_366,In_867);
xor U556 (N_556,In_110,In_1297);
nand U557 (N_557,In_1534,In_1079);
nand U558 (N_558,In_1817,In_962);
xor U559 (N_559,In_585,In_188);
nand U560 (N_560,In_679,In_1565);
nand U561 (N_561,In_1247,In_932);
xnor U562 (N_562,In_103,In_277);
xnor U563 (N_563,In_966,In_492);
or U564 (N_564,In_1905,In_1741);
and U565 (N_565,In_428,In_398);
nand U566 (N_566,In_413,In_615);
nor U567 (N_567,In_626,In_1216);
nand U568 (N_568,In_548,In_333);
nand U569 (N_569,In_622,In_1220);
or U570 (N_570,In_929,In_1695);
nand U571 (N_571,In_724,In_1878);
and U572 (N_572,In_1386,In_1570);
or U573 (N_573,In_1760,In_61);
xnor U574 (N_574,In_1405,In_840);
and U575 (N_575,In_1679,In_140);
nor U576 (N_576,In_1867,In_808);
or U577 (N_577,In_796,In_937);
and U578 (N_578,In_1337,In_654);
nor U579 (N_579,In_487,In_592);
nand U580 (N_580,In_441,In_1643);
nor U581 (N_581,In_23,In_1548);
nand U582 (N_582,In_362,In_1017);
xor U583 (N_583,In_1258,In_360);
and U584 (N_584,In_12,In_1090);
or U585 (N_585,In_266,In_281);
or U586 (N_586,In_1607,In_1052);
xnor U587 (N_587,In_885,In_596);
nor U588 (N_588,In_1764,In_20);
and U589 (N_589,In_1257,In_1850);
nand U590 (N_590,In_155,In_1073);
nor U591 (N_591,In_269,In_1228);
or U592 (N_592,In_1699,In_1712);
or U593 (N_593,In_1483,In_1185);
xnor U594 (N_594,In_1805,In_1865);
nand U595 (N_595,In_123,In_1796);
or U596 (N_596,In_1234,In_242);
nor U597 (N_597,In_957,In_1497);
nor U598 (N_598,In_1422,In_732);
nand U599 (N_599,In_689,In_1853);
xnor U600 (N_600,In_1827,In_573);
and U601 (N_601,In_697,In_781);
or U602 (N_602,In_934,In_410);
nor U603 (N_603,In_1292,In_78);
nand U604 (N_604,In_119,In_396);
nand U605 (N_605,In_595,In_1866);
xor U606 (N_606,In_1403,In_1276);
nor U607 (N_607,In_513,In_137);
nor U608 (N_608,In_1095,In_1096);
nor U609 (N_609,In_1057,In_1432);
nand U610 (N_610,In_1112,In_1130);
nand U611 (N_611,In_802,In_1595);
nand U612 (N_612,In_1078,In_70);
nor U613 (N_613,In_25,In_275);
or U614 (N_614,In_621,In_1441);
and U615 (N_615,In_900,In_1859);
or U616 (N_616,In_30,In_332);
or U617 (N_617,In_34,In_335);
and U618 (N_618,In_257,In_1968);
or U619 (N_619,In_1620,In_1573);
xnor U620 (N_620,In_1762,In_300);
nand U621 (N_621,In_1420,In_149);
nand U622 (N_622,In_1252,In_1893);
and U623 (N_623,In_1217,In_165);
or U624 (N_624,In_1423,In_763);
and U625 (N_625,In_13,In_270);
and U626 (N_626,In_780,In_115);
and U627 (N_627,In_805,In_651);
or U628 (N_628,In_1933,In_177);
nand U629 (N_629,In_1515,In_1496);
xnor U630 (N_630,In_1421,In_1341);
and U631 (N_631,In_318,In_1394);
or U632 (N_632,In_1152,In_274);
nand U633 (N_633,In_1981,In_1935);
or U634 (N_634,In_1361,In_129);
xor U635 (N_635,In_598,In_664);
nand U636 (N_636,In_1064,In_676);
nand U637 (N_637,In_542,In_828);
and U638 (N_638,In_1328,In_1798);
or U639 (N_639,In_152,In_1069);
xnor U640 (N_640,In_1020,In_1140);
nor U641 (N_641,In_1561,In_403);
nand U642 (N_642,In_604,In_1382);
and U643 (N_643,In_180,In_1314);
nand U644 (N_644,In_1498,In_1123);
and U645 (N_645,In_1694,In_1686);
xnor U646 (N_646,In_414,In_47);
xor U647 (N_647,In_377,In_491);
nand U648 (N_648,In_577,In_1962);
nand U649 (N_649,In_1735,In_678);
nand U650 (N_650,In_1365,In_84);
or U651 (N_651,In_1045,In_1375);
nor U652 (N_652,In_845,In_1134);
nand U653 (N_653,In_4,In_126);
xnor U654 (N_654,In_1290,In_1941);
xor U655 (N_655,In_1945,In_913);
xor U656 (N_656,In_1761,In_722);
nand U657 (N_657,In_38,In_1980);
and U658 (N_658,In_1891,In_671);
xor U659 (N_659,In_1105,In_1844);
and U660 (N_660,In_1834,In_880);
or U661 (N_661,In_521,In_829);
nor U662 (N_662,In_484,In_1889);
nor U663 (N_663,In_1915,In_1066);
and U664 (N_664,In_1178,In_659);
nor U665 (N_665,In_346,In_1984);
and U666 (N_666,In_1685,In_907);
nand U667 (N_667,In_63,In_1706);
or U668 (N_668,In_1281,In_684);
xnor U669 (N_669,In_202,In_1825);
nand U670 (N_670,In_774,In_800);
nand U671 (N_671,In_381,In_1367);
and U672 (N_672,In_1032,In_1137);
and U673 (N_673,In_1689,In_94);
nor U674 (N_674,In_133,In_481);
nor U675 (N_675,In_1164,In_619);
or U676 (N_676,In_890,In_293);
nand U677 (N_677,In_1592,In_1803);
or U678 (N_678,In_924,In_1183);
and U679 (N_679,In_750,In_1518);
xnor U680 (N_680,In_1307,In_680);
and U681 (N_681,In_630,In_1262);
and U682 (N_682,In_279,In_1884);
or U683 (N_683,In_1315,In_421);
and U684 (N_684,In_1150,In_424);
nand U685 (N_685,In_1711,In_1268);
and U686 (N_686,In_167,In_1640);
xnor U687 (N_687,In_1702,In_241);
nand U688 (N_688,In_721,In_980);
nand U689 (N_689,In_641,In_1407);
nand U690 (N_690,In_1454,In_1782);
nor U691 (N_691,In_541,In_1148);
nand U692 (N_692,In_388,In_1716);
nor U693 (N_693,In_1451,In_1413);
xnor U694 (N_694,In_1191,In_1810);
and U695 (N_695,In_945,In_91);
or U696 (N_696,In_302,In_1819);
nor U697 (N_697,In_1174,In_304);
nand U698 (N_698,In_1092,In_712);
nand U699 (N_699,In_479,In_930);
or U700 (N_700,In_1868,In_1273);
or U701 (N_701,In_613,In_1288);
xnor U702 (N_702,In_645,In_288);
xnor U703 (N_703,In_1047,In_1468);
and U704 (N_704,In_570,In_134);
xnor U705 (N_705,In_1396,In_1442);
or U706 (N_706,In_1833,In_665);
nor U707 (N_707,In_1988,In_79);
or U708 (N_708,In_216,In_472);
or U709 (N_709,In_1623,In_1628);
or U710 (N_710,In_902,In_330);
nor U711 (N_711,In_783,In_273);
nor U712 (N_712,In_1224,In_1637);
nand U713 (N_713,In_1402,In_1013);
and U714 (N_714,In_328,In_425);
or U715 (N_715,In_1070,In_1466);
or U716 (N_716,In_1144,In_1457);
or U717 (N_717,In_1751,In_470);
and U718 (N_718,In_963,In_147);
or U719 (N_719,In_575,In_702);
xor U720 (N_720,In_1237,In_844);
xor U721 (N_721,In_1512,In_1251);
nand U722 (N_722,In_682,In_740);
and U723 (N_723,In_925,In_646);
or U724 (N_724,In_1524,In_1581);
and U725 (N_725,In_480,In_734);
or U726 (N_726,In_1249,In_835);
and U727 (N_727,In_327,In_525);
nand U728 (N_728,In_749,In_1054);
nand U729 (N_729,In_258,In_386);
nor U730 (N_730,In_1316,In_1167);
xnor U731 (N_731,In_285,In_1922);
or U732 (N_732,In_250,In_1769);
nand U733 (N_733,In_1208,In_56);
and U734 (N_734,In_789,In_1508);
or U735 (N_735,In_1836,In_243);
nand U736 (N_736,In_849,In_1804);
xor U737 (N_737,In_1448,In_395);
xor U738 (N_738,In_337,In_240);
and U739 (N_739,In_466,In_92);
xnor U740 (N_740,In_1843,In_634);
and U741 (N_741,In_1858,In_1589);
and U742 (N_742,In_1990,In_1033);
nand U743 (N_743,In_1888,In_1632);
xnor U744 (N_744,In_1357,In_813);
nand U745 (N_745,In_699,In_1221);
and U746 (N_746,In_1225,In_1820);
or U747 (N_747,In_1660,In_1149);
nor U748 (N_748,In_1068,In_148);
nor U749 (N_749,In_49,In_199);
and U750 (N_750,In_82,In_1932);
or U751 (N_751,In_1223,In_1631);
or U752 (N_752,In_497,In_1264);
xnor U753 (N_753,In_88,In_1656);
or U754 (N_754,In_1397,In_1082);
xor U755 (N_755,In_1189,In_1668);
and U756 (N_756,In_1104,In_292);
xnor U757 (N_757,In_1644,In_669);
xnor U758 (N_758,In_339,In_792);
xnor U759 (N_759,In_1807,In_1170);
and U760 (N_760,In_15,In_1739);
or U761 (N_761,In_1744,In_1352);
or U762 (N_762,In_255,In_1369);
nand U763 (N_763,In_406,In_920);
or U764 (N_764,In_263,In_1410);
or U765 (N_765,In_144,In_1350);
nor U766 (N_766,In_1666,In_453);
or U767 (N_767,In_701,In_1398);
nor U768 (N_768,In_899,In_583);
nor U769 (N_769,In_1198,In_294);
nor U770 (N_770,In_687,In_1814);
nand U771 (N_771,In_922,In_590);
nor U772 (N_772,In_1800,In_520);
nor U773 (N_773,In_985,In_1641);
and U774 (N_774,In_1916,In_511);
nor U775 (N_775,In_1546,In_1727);
xor U776 (N_776,In_1176,In_1291);
nor U777 (N_777,In_638,In_1505);
and U778 (N_778,In_861,In_1848);
and U779 (N_779,In_372,In_1246);
nand U780 (N_780,In_1902,In_440);
nand U781 (N_781,In_785,In_587);
nor U782 (N_782,In_1677,In_368);
nand U783 (N_783,In_432,In_1311);
nor U784 (N_784,In_1030,In_54);
xor U785 (N_785,In_1046,In_182);
and U786 (N_786,In_1586,In_1734);
nand U787 (N_787,In_1437,In_1260);
nand U788 (N_788,In_726,In_253);
and U789 (N_789,In_1948,In_1624);
xor U790 (N_790,In_759,In_720);
and U791 (N_791,In_1949,In_434);
xor U792 (N_792,In_976,In_1983);
or U793 (N_793,In_801,In_1619);
xnor U794 (N_794,In_606,In_1492);
xor U795 (N_795,In_1027,In_1231);
xor U796 (N_796,In_603,In_1485);
xor U797 (N_797,In_1610,In_1567);
nor U798 (N_798,In_1790,In_347);
or U799 (N_799,In_831,In_1583);
xor U800 (N_800,In_1475,In_1277);
xnor U801 (N_801,In_1427,In_946);
nand U802 (N_802,In_1841,In_1255);
or U803 (N_803,In_572,In_1197);
or U804 (N_804,In_504,In_1882);
and U805 (N_805,In_1414,In_95);
xnor U806 (N_806,In_1026,In_1971);
and U807 (N_807,In_1635,In_1101);
nand U808 (N_808,In_916,In_897);
nand U809 (N_809,In_556,In_1000);
nor U810 (N_810,In_1813,In_1113);
or U811 (N_811,In_1909,In_356);
nand U812 (N_812,In_874,In_1767);
nor U813 (N_813,In_1982,In_1545);
or U814 (N_814,In_361,In_951);
and U815 (N_815,In_1,In_1359);
or U816 (N_816,In_1960,In_111);
and U817 (N_817,In_178,In_1098);
nor U818 (N_818,In_1490,In_1862);
nand U819 (N_819,In_7,In_1809);
nor U820 (N_820,In_1012,In_1539);
xor U821 (N_821,In_1753,In_662);
nor U822 (N_822,In_141,In_688);
nand U823 (N_823,In_260,In_31);
nor U824 (N_824,In_1562,In_560);
and U825 (N_825,In_1550,In_968);
nand U826 (N_826,In_1822,In_1440);
and U827 (N_827,In_1200,In_807);
nand U828 (N_828,In_1996,In_32);
nor U829 (N_829,In_971,In_1849);
xnor U830 (N_830,In_128,In_1870);
or U831 (N_831,In_791,In_40);
nor U832 (N_832,In_1126,In_1010);
and U833 (N_833,In_1754,In_1259);
nand U834 (N_834,In_938,In_357);
or U835 (N_835,In_766,In_1847);
nor U836 (N_836,In_1743,In_1542);
and U837 (N_837,In_98,In_62);
or U838 (N_838,In_611,In_355);
nand U839 (N_839,In_1513,In_949);
and U840 (N_840,In_309,In_1967);
nor U841 (N_841,In_1816,In_297);
or U842 (N_842,In_1613,In_1011);
or U843 (N_843,In_562,In_704);
xnor U844 (N_844,In_506,In_1482);
nor U845 (N_845,In_512,In_1215);
or U846 (N_846,In_1136,In_1270);
nand U847 (N_847,In_975,In_1240);
xnor U848 (N_848,In_1553,In_1840);
nand U849 (N_849,In_1202,In_1908);
nand U850 (N_850,In_1776,In_1789);
nor U851 (N_851,In_380,In_1374);
xor U852 (N_852,In_947,In_993);
and U853 (N_853,In_1388,In_21);
or U854 (N_854,In_836,In_1598);
or U855 (N_855,In_1243,In_1239);
xnor U856 (N_856,In_738,In_1520);
and U857 (N_857,In_1898,In_1821);
nor U858 (N_858,In_903,In_1173);
nor U859 (N_859,In_1435,In_1901);
nand U860 (N_860,In_1806,In_503);
nand U861 (N_861,In_1876,In_1939);
and U862 (N_862,In_1645,In_1729);
xor U863 (N_863,In_1892,In_612);
and U864 (N_864,In_1354,In_308);
or U865 (N_865,In_1487,In_102);
xor U866 (N_866,In_647,In_1387);
xor U867 (N_867,In_755,In_1071);
or U868 (N_868,In_816,In_1709);
nor U869 (N_869,In_1436,In_1428);
xnor U870 (N_870,In_1143,In_1978);
nand U871 (N_871,In_201,In_1393);
and U872 (N_872,In_1894,In_1992);
xnor U873 (N_873,In_736,In_1024);
or U874 (N_874,In_1715,In_1852);
xnor U875 (N_875,In_454,In_782);
nand U876 (N_876,In_776,In_1773);
or U877 (N_877,In_120,In_1942);
or U878 (N_878,In_163,In_359);
nor U879 (N_879,In_64,In_1254);
and U880 (N_880,In_341,In_1499);
and U881 (N_881,In_283,In_1424);
and U882 (N_882,In_1543,In_1018);
nor U883 (N_883,In_923,In_950);
or U884 (N_884,In_225,In_1245);
and U885 (N_885,In_1323,In_435);
nor U886 (N_886,In_1626,In_875);
and U887 (N_887,In_1975,In_495);
xnor U888 (N_888,In_965,In_865);
or U889 (N_889,In_617,In_1529);
xnor U890 (N_890,In_943,In_683);
nor U891 (N_891,In_437,In_714);
and U892 (N_892,In_1831,In_338);
nand U893 (N_893,In_1384,In_146);
or U894 (N_894,In_131,In_127);
nand U895 (N_895,In_1416,In_1811);
nand U896 (N_896,In_1742,In_1204);
nand U897 (N_897,In_1280,In_1591);
nand U898 (N_898,In_927,In_1004);
and U899 (N_899,In_227,In_510);
xor U900 (N_900,In_1793,In_415);
and U901 (N_901,In_578,In_1593);
nor U902 (N_902,In_519,In_448);
nand U903 (N_903,In_1936,In_50);
xor U904 (N_904,In_1869,In_1184);
nor U905 (N_905,In_1272,In_1823);
nor U906 (N_906,In_483,In_1063);
and U907 (N_907,In_1266,In_1118);
xor U908 (N_908,In_1580,In_1081);
xor U909 (N_909,In_817,In_326);
and U910 (N_910,In_768,In_1389);
nor U911 (N_911,In_43,In_76);
and U912 (N_912,In_1681,In_387);
and U913 (N_913,In_954,In_1538);
or U914 (N_914,In_977,In_1298);
xnor U915 (N_915,In_1930,In_1895);
or U916 (N_916,In_1088,In_745);
xor U917 (N_917,In_1007,In_1283);
or U918 (N_918,In_1261,In_154);
and U919 (N_919,In_810,In_1780);
nor U920 (N_920,In_919,In_205);
nor U921 (N_921,In_1409,In_1180);
and U922 (N_922,In_231,In_474);
nand U923 (N_923,In_1523,In_1269);
nor U924 (N_924,In_1927,In_1263);
and U925 (N_925,In_1556,In_1509);
nor U926 (N_926,In_391,In_456);
and U927 (N_927,In_761,In_1195);
and U928 (N_928,In_1897,In_161);
and U929 (N_929,In_859,In_633);
or U930 (N_930,In_108,In_1615);
nand U931 (N_931,In_1360,In_1758);
nand U932 (N_932,In_206,In_1725);
xor U933 (N_933,In_1678,In_185);
or U934 (N_934,In_1994,In_1676);
nor U935 (N_935,In_803,In_1618);
and U936 (N_936,In_1797,In_1904);
xor U937 (N_937,In_941,In_1131);
and U938 (N_938,In_145,In_1765);
nor U939 (N_939,In_960,In_1956);
or U940 (N_940,In_752,In_419);
and U941 (N_941,In_1196,In_868);
nand U942 (N_942,In_80,In_1218);
or U943 (N_943,In_1730,In_986);
nor U944 (N_944,In_1250,In_1145);
nor U945 (N_945,In_1549,In_245);
and U946 (N_946,In_1722,In_463);
nor U947 (N_947,In_821,In_1275);
nor U948 (N_948,In_1213,In_105);
xnor U949 (N_949,In_11,In_1872);
or U950 (N_950,In_1582,In_1194);
or U951 (N_951,In_655,In_1603);
or U952 (N_952,In_610,In_998);
nor U953 (N_953,In_287,In_864);
and U954 (N_954,In_744,In_204);
or U955 (N_955,In_1122,In_666);
nand U956 (N_956,In_686,In_1444);
xnor U957 (N_957,In_1406,In_1944);
or U958 (N_958,In_1877,In_1426);
xnor U959 (N_959,In_1701,In_267);
and U960 (N_960,In_1236,In_1065);
and U961 (N_961,In_1230,In_564);
or U962 (N_962,In_673,In_1777);
nor U963 (N_963,In_910,In_1647);
or U964 (N_964,In_1175,In_169);
and U965 (N_965,In_981,In_1037);
nor U966 (N_966,In_538,In_384);
xnor U967 (N_967,In_887,In_1304);
and U968 (N_968,In_75,In_299);
nor U969 (N_969,In_193,In_465);
or U970 (N_970,In_690,In_703);
nand U971 (N_971,In_1842,In_1781);
and U972 (N_972,In_179,In_1900);
nand U973 (N_973,In_303,In_854);
or U974 (N_974,In_331,In_1008);
xor U975 (N_975,In_156,In_1434);
or U976 (N_976,In_1128,In_942);
nand U977 (N_977,In_1271,In_1053);
nand U978 (N_978,In_420,In_1659);
and U979 (N_979,In_1611,In_1301);
nand U980 (N_980,In_827,In_1745);
nor U981 (N_981,In_343,In_1519);
or U982 (N_982,In_393,In_1205);
nand U983 (N_983,In_609,In_1871);
or U984 (N_984,In_1479,In_1253);
and U985 (N_985,In_1327,In_1331);
nor U986 (N_986,In_629,In_1347);
and U987 (N_987,In_426,In_1557);
or U988 (N_988,In_944,In_1502);
xor U989 (N_989,In_707,In_940);
xnor U990 (N_990,In_1506,In_952);
and U991 (N_991,In_1724,In_1794);
xor U992 (N_992,In_1142,In_754);
nand U993 (N_993,In_1665,In_1728);
nand U994 (N_994,In_825,In_786);
xnor U995 (N_995,In_1664,In_1097);
nand U996 (N_996,In_1602,In_449);
and U997 (N_997,In_1021,In_1650);
xnor U998 (N_998,In_884,In_1684);
nand U999 (N_999,In_1540,In_1587);
xor U1000 (N_1000,In_234,In_1901);
xnor U1001 (N_1001,In_1656,In_1086);
xnor U1002 (N_1002,In_1012,In_1804);
and U1003 (N_1003,In_757,In_1620);
nor U1004 (N_1004,In_1083,In_216);
nor U1005 (N_1005,In_633,In_1813);
nor U1006 (N_1006,In_1063,In_719);
xor U1007 (N_1007,In_760,In_1441);
nor U1008 (N_1008,In_1221,In_1885);
xnor U1009 (N_1009,In_810,In_1599);
xor U1010 (N_1010,In_1485,In_1633);
xor U1011 (N_1011,In_1624,In_1734);
or U1012 (N_1012,In_1387,In_114);
nand U1013 (N_1013,In_957,In_874);
xor U1014 (N_1014,In_113,In_310);
xnor U1015 (N_1015,In_130,In_1031);
xor U1016 (N_1016,In_1277,In_1741);
nor U1017 (N_1017,In_1736,In_1463);
or U1018 (N_1018,In_243,In_331);
and U1019 (N_1019,In_1185,In_646);
or U1020 (N_1020,In_1854,In_698);
xor U1021 (N_1021,In_1018,In_1406);
or U1022 (N_1022,In_408,In_622);
or U1023 (N_1023,In_1488,In_1601);
xor U1024 (N_1024,In_381,In_1303);
nor U1025 (N_1025,In_197,In_1463);
or U1026 (N_1026,In_563,In_153);
nand U1027 (N_1027,In_378,In_473);
and U1028 (N_1028,In_721,In_589);
xnor U1029 (N_1029,In_1758,In_1673);
or U1030 (N_1030,In_415,In_1578);
and U1031 (N_1031,In_1782,In_1471);
nand U1032 (N_1032,In_913,In_1558);
and U1033 (N_1033,In_1303,In_1410);
nand U1034 (N_1034,In_340,In_1289);
xnor U1035 (N_1035,In_1098,In_1344);
xnor U1036 (N_1036,In_1196,In_1822);
xor U1037 (N_1037,In_1301,In_1828);
nor U1038 (N_1038,In_1036,In_266);
or U1039 (N_1039,In_1404,In_1793);
or U1040 (N_1040,In_514,In_1807);
xor U1041 (N_1041,In_1560,In_1572);
or U1042 (N_1042,In_1208,In_635);
or U1043 (N_1043,In_1457,In_1340);
or U1044 (N_1044,In_995,In_700);
and U1045 (N_1045,In_1277,In_1923);
nor U1046 (N_1046,In_1142,In_524);
nand U1047 (N_1047,In_817,In_496);
nand U1048 (N_1048,In_563,In_629);
or U1049 (N_1049,In_1311,In_84);
and U1050 (N_1050,In_51,In_939);
or U1051 (N_1051,In_162,In_1483);
and U1052 (N_1052,In_504,In_1644);
and U1053 (N_1053,In_1742,In_208);
nor U1054 (N_1054,In_140,In_1098);
nand U1055 (N_1055,In_904,In_902);
nor U1056 (N_1056,In_1361,In_255);
or U1057 (N_1057,In_230,In_93);
nor U1058 (N_1058,In_453,In_605);
or U1059 (N_1059,In_776,In_867);
and U1060 (N_1060,In_409,In_190);
nand U1061 (N_1061,In_935,In_1922);
and U1062 (N_1062,In_1289,In_1615);
and U1063 (N_1063,In_404,In_508);
nor U1064 (N_1064,In_1457,In_1490);
and U1065 (N_1065,In_3,In_1862);
nor U1066 (N_1066,In_1285,In_1476);
or U1067 (N_1067,In_1641,In_1416);
and U1068 (N_1068,In_1181,In_454);
and U1069 (N_1069,In_1996,In_1566);
or U1070 (N_1070,In_1940,In_1000);
nor U1071 (N_1071,In_91,In_908);
or U1072 (N_1072,In_1453,In_1048);
xor U1073 (N_1073,In_1491,In_1437);
xnor U1074 (N_1074,In_213,In_1724);
and U1075 (N_1075,In_768,In_1125);
or U1076 (N_1076,In_1145,In_308);
nand U1077 (N_1077,In_1322,In_1357);
and U1078 (N_1078,In_75,In_1663);
xor U1079 (N_1079,In_1002,In_1065);
nand U1080 (N_1080,In_81,In_1083);
nand U1081 (N_1081,In_77,In_1001);
and U1082 (N_1082,In_1913,In_1891);
nand U1083 (N_1083,In_1431,In_268);
and U1084 (N_1084,In_1732,In_617);
or U1085 (N_1085,In_331,In_67);
nand U1086 (N_1086,In_99,In_1905);
and U1087 (N_1087,In_971,In_1283);
nor U1088 (N_1088,In_824,In_1218);
xor U1089 (N_1089,In_983,In_1106);
xnor U1090 (N_1090,In_993,In_1828);
or U1091 (N_1091,In_84,In_830);
xor U1092 (N_1092,In_1440,In_656);
xnor U1093 (N_1093,In_1299,In_1256);
or U1094 (N_1094,In_1017,In_1029);
or U1095 (N_1095,In_1359,In_508);
nor U1096 (N_1096,In_1818,In_727);
or U1097 (N_1097,In_1320,In_1639);
nand U1098 (N_1098,In_929,In_1407);
or U1099 (N_1099,In_344,In_1887);
xnor U1100 (N_1100,In_1919,In_1399);
nand U1101 (N_1101,In_1605,In_1632);
nand U1102 (N_1102,In_1075,In_1525);
nor U1103 (N_1103,In_974,In_88);
nor U1104 (N_1104,In_572,In_264);
and U1105 (N_1105,In_1314,In_1927);
xnor U1106 (N_1106,In_197,In_1873);
and U1107 (N_1107,In_1346,In_1632);
and U1108 (N_1108,In_1416,In_60);
and U1109 (N_1109,In_1527,In_157);
and U1110 (N_1110,In_139,In_1301);
nor U1111 (N_1111,In_522,In_143);
or U1112 (N_1112,In_831,In_1223);
or U1113 (N_1113,In_532,In_1775);
and U1114 (N_1114,In_607,In_893);
nor U1115 (N_1115,In_1384,In_1338);
nor U1116 (N_1116,In_1278,In_1779);
or U1117 (N_1117,In_1437,In_968);
and U1118 (N_1118,In_880,In_155);
or U1119 (N_1119,In_1096,In_77);
nor U1120 (N_1120,In_256,In_1564);
or U1121 (N_1121,In_823,In_437);
nand U1122 (N_1122,In_244,In_643);
nand U1123 (N_1123,In_294,In_1370);
or U1124 (N_1124,In_1046,In_819);
nor U1125 (N_1125,In_397,In_1196);
nand U1126 (N_1126,In_1749,In_741);
or U1127 (N_1127,In_1546,In_1115);
nor U1128 (N_1128,In_1122,In_1685);
and U1129 (N_1129,In_1644,In_247);
nor U1130 (N_1130,In_361,In_37);
nor U1131 (N_1131,In_670,In_414);
and U1132 (N_1132,In_1173,In_264);
and U1133 (N_1133,In_1360,In_297);
nand U1134 (N_1134,In_1277,In_825);
xor U1135 (N_1135,In_175,In_770);
xor U1136 (N_1136,In_653,In_1824);
nor U1137 (N_1137,In_1422,In_1293);
or U1138 (N_1138,In_1249,In_602);
and U1139 (N_1139,In_612,In_769);
and U1140 (N_1140,In_1460,In_317);
xor U1141 (N_1141,In_1965,In_1790);
or U1142 (N_1142,In_441,In_1783);
nor U1143 (N_1143,In_1853,In_1319);
nand U1144 (N_1144,In_680,In_879);
nor U1145 (N_1145,In_1722,In_1149);
xor U1146 (N_1146,In_1299,In_1685);
or U1147 (N_1147,In_959,In_600);
nor U1148 (N_1148,In_1077,In_1651);
or U1149 (N_1149,In_1263,In_150);
xnor U1150 (N_1150,In_1985,In_901);
nor U1151 (N_1151,In_879,In_1121);
or U1152 (N_1152,In_621,In_1882);
nand U1153 (N_1153,In_964,In_394);
and U1154 (N_1154,In_1860,In_1410);
xnor U1155 (N_1155,In_801,In_1343);
nand U1156 (N_1156,In_619,In_1586);
or U1157 (N_1157,In_1167,In_930);
nand U1158 (N_1158,In_918,In_732);
and U1159 (N_1159,In_1085,In_994);
nor U1160 (N_1160,In_241,In_559);
or U1161 (N_1161,In_654,In_1401);
or U1162 (N_1162,In_1369,In_250);
or U1163 (N_1163,In_1390,In_1843);
xor U1164 (N_1164,In_64,In_1238);
xor U1165 (N_1165,In_1510,In_1871);
or U1166 (N_1166,In_1950,In_79);
or U1167 (N_1167,In_1779,In_823);
xor U1168 (N_1168,In_660,In_20);
xnor U1169 (N_1169,In_1700,In_1893);
nand U1170 (N_1170,In_495,In_724);
xor U1171 (N_1171,In_1318,In_1416);
nand U1172 (N_1172,In_1344,In_1652);
nand U1173 (N_1173,In_1257,In_1968);
nor U1174 (N_1174,In_408,In_1238);
nor U1175 (N_1175,In_1086,In_852);
nand U1176 (N_1176,In_1193,In_191);
or U1177 (N_1177,In_133,In_539);
xor U1178 (N_1178,In_1251,In_612);
nor U1179 (N_1179,In_1555,In_191);
and U1180 (N_1180,In_1922,In_1445);
nand U1181 (N_1181,In_1723,In_874);
or U1182 (N_1182,In_15,In_1523);
xnor U1183 (N_1183,In_673,In_1314);
and U1184 (N_1184,In_1343,In_970);
nand U1185 (N_1185,In_866,In_1797);
nand U1186 (N_1186,In_1102,In_974);
nand U1187 (N_1187,In_655,In_796);
nand U1188 (N_1188,In_140,In_1859);
or U1189 (N_1189,In_84,In_549);
nor U1190 (N_1190,In_1007,In_1286);
or U1191 (N_1191,In_244,In_1953);
xnor U1192 (N_1192,In_1740,In_38);
nand U1193 (N_1193,In_1103,In_850);
and U1194 (N_1194,In_804,In_462);
nand U1195 (N_1195,In_1583,In_439);
xor U1196 (N_1196,In_1580,In_1073);
nand U1197 (N_1197,In_1164,In_634);
nand U1198 (N_1198,In_1805,In_1560);
nor U1199 (N_1199,In_194,In_1919);
or U1200 (N_1200,In_1869,In_1828);
nor U1201 (N_1201,In_592,In_360);
or U1202 (N_1202,In_912,In_594);
nor U1203 (N_1203,In_1870,In_1421);
or U1204 (N_1204,In_590,In_888);
nor U1205 (N_1205,In_544,In_1548);
nand U1206 (N_1206,In_1452,In_447);
nor U1207 (N_1207,In_1600,In_1004);
nor U1208 (N_1208,In_1609,In_1479);
nor U1209 (N_1209,In_1933,In_280);
and U1210 (N_1210,In_232,In_1509);
or U1211 (N_1211,In_1913,In_1667);
and U1212 (N_1212,In_163,In_1017);
xor U1213 (N_1213,In_113,In_1340);
nand U1214 (N_1214,In_1741,In_1171);
and U1215 (N_1215,In_1643,In_1701);
xor U1216 (N_1216,In_555,In_1212);
and U1217 (N_1217,In_475,In_1529);
and U1218 (N_1218,In_546,In_138);
nor U1219 (N_1219,In_981,In_645);
nand U1220 (N_1220,In_176,In_1308);
or U1221 (N_1221,In_618,In_1947);
and U1222 (N_1222,In_1572,In_392);
nand U1223 (N_1223,In_376,In_272);
xnor U1224 (N_1224,In_800,In_47);
or U1225 (N_1225,In_1651,In_117);
nor U1226 (N_1226,In_309,In_178);
xor U1227 (N_1227,In_1072,In_1234);
or U1228 (N_1228,In_1334,In_1506);
nand U1229 (N_1229,In_781,In_519);
and U1230 (N_1230,In_1279,In_299);
nand U1231 (N_1231,In_895,In_1484);
or U1232 (N_1232,In_1756,In_676);
xor U1233 (N_1233,In_1322,In_1245);
xor U1234 (N_1234,In_71,In_1575);
or U1235 (N_1235,In_614,In_1988);
or U1236 (N_1236,In_127,In_1236);
xor U1237 (N_1237,In_793,In_839);
and U1238 (N_1238,In_825,In_1330);
nand U1239 (N_1239,In_961,In_1345);
and U1240 (N_1240,In_855,In_1998);
nand U1241 (N_1241,In_239,In_1488);
nor U1242 (N_1242,In_1178,In_1579);
and U1243 (N_1243,In_1685,In_1608);
nor U1244 (N_1244,In_1341,In_1269);
or U1245 (N_1245,In_543,In_1083);
xor U1246 (N_1246,In_598,In_970);
nor U1247 (N_1247,In_1178,In_674);
nor U1248 (N_1248,In_286,In_53);
and U1249 (N_1249,In_31,In_284);
nor U1250 (N_1250,In_312,In_956);
nand U1251 (N_1251,In_694,In_87);
nand U1252 (N_1252,In_1799,In_1060);
or U1253 (N_1253,In_1075,In_1524);
xnor U1254 (N_1254,In_1932,In_1039);
xor U1255 (N_1255,In_1209,In_1519);
nor U1256 (N_1256,In_1169,In_1017);
nand U1257 (N_1257,In_1492,In_1145);
or U1258 (N_1258,In_1,In_278);
or U1259 (N_1259,In_206,In_1142);
nor U1260 (N_1260,In_1016,In_21);
and U1261 (N_1261,In_1351,In_557);
xor U1262 (N_1262,In_818,In_1904);
and U1263 (N_1263,In_73,In_318);
nand U1264 (N_1264,In_67,In_1541);
and U1265 (N_1265,In_899,In_1642);
or U1266 (N_1266,In_1545,In_156);
and U1267 (N_1267,In_962,In_1850);
nand U1268 (N_1268,In_610,In_516);
xor U1269 (N_1269,In_1450,In_898);
nor U1270 (N_1270,In_1523,In_721);
or U1271 (N_1271,In_99,In_968);
and U1272 (N_1272,In_1857,In_1873);
nand U1273 (N_1273,In_622,In_478);
and U1274 (N_1274,In_1412,In_981);
and U1275 (N_1275,In_921,In_403);
and U1276 (N_1276,In_1020,In_837);
xnor U1277 (N_1277,In_85,In_1999);
and U1278 (N_1278,In_70,In_900);
nor U1279 (N_1279,In_1179,In_69);
nand U1280 (N_1280,In_1815,In_557);
and U1281 (N_1281,In_419,In_1778);
or U1282 (N_1282,In_1479,In_1906);
nor U1283 (N_1283,In_527,In_1235);
nand U1284 (N_1284,In_1219,In_1874);
nand U1285 (N_1285,In_136,In_1070);
and U1286 (N_1286,In_1896,In_28);
or U1287 (N_1287,In_1576,In_903);
nand U1288 (N_1288,In_735,In_1186);
nor U1289 (N_1289,In_1315,In_825);
xnor U1290 (N_1290,In_96,In_1168);
and U1291 (N_1291,In_1480,In_343);
and U1292 (N_1292,In_1052,In_612);
xor U1293 (N_1293,In_325,In_1870);
xor U1294 (N_1294,In_1197,In_589);
and U1295 (N_1295,In_1617,In_93);
nor U1296 (N_1296,In_745,In_1122);
or U1297 (N_1297,In_1052,In_797);
nand U1298 (N_1298,In_366,In_1388);
and U1299 (N_1299,In_378,In_400);
or U1300 (N_1300,In_982,In_738);
xor U1301 (N_1301,In_868,In_519);
nor U1302 (N_1302,In_320,In_4);
nand U1303 (N_1303,In_1128,In_1459);
nand U1304 (N_1304,In_1700,In_1912);
or U1305 (N_1305,In_151,In_1877);
nand U1306 (N_1306,In_1913,In_405);
nor U1307 (N_1307,In_1313,In_510);
and U1308 (N_1308,In_1127,In_147);
nand U1309 (N_1309,In_556,In_1202);
nand U1310 (N_1310,In_1209,In_551);
or U1311 (N_1311,In_1975,In_1482);
nand U1312 (N_1312,In_710,In_1465);
and U1313 (N_1313,In_148,In_690);
nand U1314 (N_1314,In_197,In_1793);
or U1315 (N_1315,In_1158,In_103);
or U1316 (N_1316,In_964,In_1161);
and U1317 (N_1317,In_464,In_481);
and U1318 (N_1318,In_1403,In_961);
or U1319 (N_1319,In_567,In_67);
xnor U1320 (N_1320,In_822,In_1599);
or U1321 (N_1321,In_1184,In_1421);
nor U1322 (N_1322,In_811,In_1410);
nor U1323 (N_1323,In_148,In_1756);
and U1324 (N_1324,In_1569,In_1442);
xor U1325 (N_1325,In_1050,In_937);
nand U1326 (N_1326,In_1122,In_398);
or U1327 (N_1327,In_1666,In_1855);
or U1328 (N_1328,In_202,In_380);
and U1329 (N_1329,In_1145,In_1092);
nor U1330 (N_1330,In_1571,In_1973);
nor U1331 (N_1331,In_1805,In_352);
nand U1332 (N_1332,In_1520,In_265);
nor U1333 (N_1333,In_546,In_195);
or U1334 (N_1334,In_1117,In_377);
nand U1335 (N_1335,In_795,In_957);
nand U1336 (N_1336,In_1753,In_1243);
nor U1337 (N_1337,In_190,In_206);
nand U1338 (N_1338,In_1155,In_952);
nand U1339 (N_1339,In_1441,In_1187);
and U1340 (N_1340,In_1947,In_1683);
and U1341 (N_1341,In_425,In_398);
nor U1342 (N_1342,In_1369,In_663);
and U1343 (N_1343,In_828,In_187);
xnor U1344 (N_1344,In_1048,In_1657);
nand U1345 (N_1345,In_1135,In_1214);
and U1346 (N_1346,In_269,In_1859);
and U1347 (N_1347,In_973,In_538);
nor U1348 (N_1348,In_1371,In_829);
and U1349 (N_1349,In_396,In_877);
and U1350 (N_1350,In_1238,In_1169);
and U1351 (N_1351,In_757,In_350);
nand U1352 (N_1352,In_908,In_1395);
nor U1353 (N_1353,In_149,In_387);
or U1354 (N_1354,In_130,In_1417);
and U1355 (N_1355,In_1573,In_730);
nand U1356 (N_1356,In_1124,In_740);
and U1357 (N_1357,In_138,In_159);
nand U1358 (N_1358,In_1701,In_1250);
xnor U1359 (N_1359,In_641,In_1218);
nor U1360 (N_1360,In_77,In_1688);
or U1361 (N_1361,In_154,In_1762);
nor U1362 (N_1362,In_1826,In_513);
nand U1363 (N_1363,In_1110,In_1735);
or U1364 (N_1364,In_1449,In_534);
nand U1365 (N_1365,In_967,In_1188);
xor U1366 (N_1366,In_1763,In_244);
nand U1367 (N_1367,In_646,In_1408);
nor U1368 (N_1368,In_1745,In_1546);
nand U1369 (N_1369,In_297,In_265);
and U1370 (N_1370,In_621,In_310);
nand U1371 (N_1371,In_458,In_71);
xnor U1372 (N_1372,In_1842,In_1471);
nand U1373 (N_1373,In_1626,In_9);
nand U1374 (N_1374,In_372,In_1712);
xnor U1375 (N_1375,In_80,In_1169);
nor U1376 (N_1376,In_488,In_389);
or U1377 (N_1377,In_537,In_1234);
or U1378 (N_1378,In_1525,In_1854);
xor U1379 (N_1379,In_728,In_644);
or U1380 (N_1380,In_1552,In_867);
nor U1381 (N_1381,In_1008,In_1356);
xor U1382 (N_1382,In_1280,In_1101);
or U1383 (N_1383,In_238,In_1512);
and U1384 (N_1384,In_1601,In_621);
nand U1385 (N_1385,In_1414,In_1411);
xor U1386 (N_1386,In_140,In_1744);
nor U1387 (N_1387,In_1269,In_329);
nand U1388 (N_1388,In_1314,In_1316);
and U1389 (N_1389,In_1047,In_1224);
or U1390 (N_1390,In_297,In_1639);
nand U1391 (N_1391,In_1112,In_1550);
nor U1392 (N_1392,In_1091,In_1375);
nand U1393 (N_1393,In_767,In_1997);
nor U1394 (N_1394,In_500,In_1360);
or U1395 (N_1395,In_1109,In_1707);
and U1396 (N_1396,In_856,In_1813);
xnor U1397 (N_1397,In_1784,In_1965);
nand U1398 (N_1398,In_569,In_948);
or U1399 (N_1399,In_1784,In_1779);
xnor U1400 (N_1400,In_307,In_1697);
xnor U1401 (N_1401,In_1862,In_1989);
and U1402 (N_1402,In_31,In_216);
nand U1403 (N_1403,In_1847,In_1587);
xnor U1404 (N_1404,In_1755,In_954);
xor U1405 (N_1405,In_1756,In_1252);
or U1406 (N_1406,In_850,In_938);
xor U1407 (N_1407,In_1729,In_423);
nand U1408 (N_1408,In_209,In_1560);
nand U1409 (N_1409,In_1505,In_1006);
and U1410 (N_1410,In_1560,In_778);
nand U1411 (N_1411,In_804,In_520);
xor U1412 (N_1412,In_684,In_1069);
or U1413 (N_1413,In_666,In_1029);
nand U1414 (N_1414,In_813,In_306);
xor U1415 (N_1415,In_1125,In_353);
xor U1416 (N_1416,In_572,In_1163);
xnor U1417 (N_1417,In_1766,In_1874);
nand U1418 (N_1418,In_1460,In_1733);
nor U1419 (N_1419,In_822,In_893);
xnor U1420 (N_1420,In_1702,In_474);
or U1421 (N_1421,In_1325,In_355);
nor U1422 (N_1422,In_1043,In_1304);
xor U1423 (N_1423,In_1990,In_1793);
xor U1424 (N_1424,In_496,In_912);
nor U1425 (N_1425,In_1477,In_1221);
nor U1426 (N_1426,In_1778,In_320);
and U1427 (N_1427,In_265,In_198);
nor U1428 (N_1428,In_919,In_1418);
and U1429 (N_1429,In_1599,In_994);
and U1430 (N_1430,In_336,In_1344);
or U1431 (N_1431,In_1385,In_1602);
nand U1432 (N_1432,In_1447,In_3);
nor U1433 (N_1433,In_1225,In_1680);
nor U1434 (N_1434,In_94,In_830);
or U1435 (N_1435,In_1633,In_1878);
or U1436 (N_1436,In_672,In_1107);
nor U1437 (N_1437,In_1746,In_1641);
or U1438 (N_1438,In_756,In_1955);
nand U1439 (N_1439,In_745,In_1275);
nor U1440 (N_1440,In_1237,In_336);
and U1441 (N_1441,In_1591,In_1460);
or U1442 (N_1442,In_250,In_950);
nor U1443 (N_1443,In_242,In_516);
and U1444 (N_1444,In_1480,In_1621);
or U1445 (N_1445,In_103,In_1121);
nand U1446 (N_1446,In_520,In_1426);
or U1447 (N_1447,In_1423,In_1116);
nand U1448 (N_1448,In_0,In_730);
and U1449 (N_1449,In_612,In_226);
and U1450 (N_1450,In_798,In_464);
nand U1451 (N_1451,In_1129,In_114);
xnor U1452 (N_1452,In_1370,In_341);
xnor U1453 (N_1453,In_739,In_443);
xor U1454 (N_1454,In_705,In_1248);
xor U1455 (N_1455,In_791,In_1073);
nor U1456 (N_1456,In_1102,In_1813);
nor U1457 (N_1457,In_1271,In_816);
or U1458 (N_1458,In_396,In_30);
nand U1459 (N_1459,In_1266,In_1546);
nand U1460 (N_1460,In_752,In_244);
nor U1461 (N_1461,In_1314,In_1586);
and U1462 (N_1462,In_1786,In_1823);
and U1463 (N_1463,In_444,In_1344);
nand U1464 (N_1464,In_836,In_1484);
xnor U1465 (N_1465,In_1266,In_1421);
or U1466 (N_1466,In_1115,In_1756);
nor U1467 (N_1467,In_1531,In_857);
or U1468 (N_1468,In_1385,In_1817);
xnor U1469 (N_1469,In_1347,In_343);
and U1470 (N_1470,In_1327,In_840);
and U1471 (N_1471,In_1424,In_1246);
xor U1472 (N_1472,In_1104,In_1123);
or U1473 (N_1473,In_151,In_962);
nand U1474 (N_1474,In_1783,In_1184);
or U1475 (N_1475,In_609,In_496);
and U1476 (N_1476,In_113,In_419);
and U1477 (N_1477,In_1681,In_1763);
nand U1478 (N_1478,In_1395,In_262);
and U1479 (N_1479,In_172,In_414);
nand U1480 (N_1480,In_1939,In_145);
xor U1481 (N_1481,In_1871,In_1385);
or U1482 (N_1482,In_660,In_1770);
nand U1483 (N_1483,In_222,In_223);
nand U1484 (N_1484,In_1613,In_299);
xor U1485 (N_1485,In_1543,In_811);
nand U1486 (N_1486,In_1531,In_1234);
nand U1487 (N_1487,In_979,In_907);
and U1488 (N_1488,In_292,In_1069);
nand U1489 (N_1489,In_1320,In_232);
or U1490 (N_1490,In_1420,In_1570);
nand U1491 (N_1491,In_1176,In_199);
or U1492 (N_1492,In_1312,In_822);
xor U1493 (N_1493,In_935,In_947);
xnor U1494 (N_1494,In_1205,In_903);
or U1495 (N_1495,In_1495,In_193);
or U1496 (N_1496,In_1833,In_1276);
and U1497 (N_1497,In_576,In_1942);
xor U1498 (N_1498,In_913,In_948);
nand U1499 (N_1499,In_643,In_364);
or U1500 (N_1500,In_782,In_1029);
or U1501 (N_1501,In_1885,In_1937);
and U1502 (N_1502,In_1335,In_1276);
nand U1503 (N_1503,In_868,In_417);
nor U1504 (N_1504,In_104,In_889);
nor U1505 (N_1505,In_381,In_1843);
nor U1506 (N_1506,In_57,In_610);
xor U1507 (N_1507,In_505,In_973);
or U1508 (N_1508,In_1877,In_1017);
nor U1509 (N_1509,In_907,In_1773);
xor U1510 (N_1510,In_642,In_411);
and U1511 (N_1511,In_1038,In_1843);
nor U1512 (N_1512,In_131,In_1694);
nand U1513 (N_1513,In_249,In_578);
nor U1514 (N_1514,In_531,In_1029);
or U1515 (N_1515,In_859,In_1720);
nand U1516 (N_1516,In_632,In_977);
xor U1517 (N_1517,In_448,In_1097);
xor U1518 (N_1518,In_164,In_760);
or U1519 (N_1519,In_1064,In_1952);
nand U1520 (N_1520,In_846,In_959);
nand U1521 (N_1521,In_346,In_114);
nor U1522 (N_1522,In_337,In_1213);
xnor U1523 (N_1523,In_1788,In_1269);
nor U1524 (N_1524,In_570,In_1791);
nand U1525 (N_1525,In_281,In_896);
nor U1526 (N_1526,In_207,In_274);
nor U1527 (N_1527,In_1824,In_174);
and U1528 (N_1528,In_363,In_1217);
nor U1529 (N_1529,In_51,In_23);
nand U1530 (N_1530,In_1556,In_238);
nand U1531 (N_1531,In_1876,In_629);
nor U1532 (N_1532,In_436,In_1210);
xor U1533 (N_1533,In_426,In_1578);
nand U1534 (N_1534,In_1523,In_114);
nand U1535 (N_1535,In_1303,In_31);
nor U1536 (N_1536,In_1940,In_774);
or U1537 (N_1537,In_1838,In_907);
nand U1538 (N_1538,In_1736,In_1958);
nand U1539 (N_1539,In_54,In_1278);
nor U1540 (N_1540,In_1782,In_1899);
nor U1541 (N_1541,In_1736,In_1532);
nor U1542 (N_1542,In_709,In_246);
or U1543 (N_1543,In_1070,In_254);
or U1544 (N_1544,In_1110,In_261);
and U1545 (N_1545,In_1752,In_392);
nor U1546 (N_1546,In_406,In_1085);
xor U1547 (N_1547,In_1997,In_431);
xnor U1548 (N_1548,In_1519,In_583);
nand U1549 (N_1549,In_358,In_776);
and U1550 (N_1550,In_1644,In_436);
xor U1551 (N_1551,In_216,In_508);
nand U1552 (N_1552,In_1089,In_1109);
nand U1553 (N_1553,In_1127,In_782);
or U1554 (N_1554,In_362,In_1588);
nor U1555 (N_1555,In_1947,In_58);
or U1556 (N_1556,In_837,In_1364);
nand U1557 (N_1557,In_775,In_1064);
and U1558 (N_1558,In_1751,In_1221);
and U1559 (N_1559,In_263,In_1239);
and U1560 (N_1560,In_476,In_675);
nor U1561 (N_1561,In_429,In_1214);
or U1562 (N_1562,In_363,In_544);
nor U1563 (N_1563,In_469,In_1586);
and U1564 (N_1564,In_1635,In_363);
nor U1565 (N_1565,In_14,In_736);
nand U1566 (N_1566,In_1278,In_136);
or U1567 (N_1567,In_1411,In_1617);
xnor U1568 (N_1568,In_41,In_1579);
nor U1569 (N_1569,In_1182,In_1785);
xnor U1570 (N_1570,In_416,In_863);
and U1571 (N_1571,In_1876,In_487);
xnor U1572 (N_1572,In_571,In_204);
xor U1573 (N_1573,In_667,In_7);
or U1574 (N_1574,In_534,In_1879);
and U1575 (N_1575,In_1650,In_703);
nand U1576 (N_1576,In_921,In_695);
nor U1577 (N_1577,In_466,In_166);
and U1578 (N_1578,In_229,In_1669);
and U1579 (N_1579,In_682,In_1037);
nor U1580 (N_1580,In_1965,In_238);
nor U1581 (N_1581,In_568,In_0);
or U1582 (N_1582,In_551,In_1111);
and U1583 (N_1583,In_970,In_1751);
nor U1584 (N_1584,In_721,In_1408);
nand U1585 (N_1585,In_79,In_1659);
or U1586 (N_1586,In_952,In_802);
nand U1587 (N_1587,In_1908,In_1670);
nand U1588 (N_1588,In_927,In_1310);
nor U1589 (N_1589,In_77,In_218);
xor U1590 (N_1590,In_810,In_1565);
nor U1591 (N_1591,In_1022,In_1279);
xnor U1592 (N_1592,In_67,In_122);
nand U1593 (N_1593,In_262,In_1672);
nand U1594 (N_1594,In_73,In_1339);
and U1595 (N_1595,In_1064,In_325);
xor U1596 (N_1596,In_202,In_796);
nand U1597 (N_1597,In_1829,In_60);
nor U1598 (N_1598,In_1954,In_107);
nand U1599 (N_1599,In_1613,In_594);
or U1600 (N_1600,In_1948,In_187);
xor U1601 (N_1601,In_1747,In_788);
nor U1602 (N_1602,In_299,In_1649);
or U1603 (N_1603,In_400,In_500);
nand U1604 (N_1604,In_1338,In_1884);
and U1605 (N_1605,In_1847,In_1694);
nand U1606 (N_1606,In_636,In_1349);
or U1607 (N_1607,In_462,In_906);
nand U1608 (N_1608,In_465,In_1549);
nand U1609 (N_1609,In_1837,In_944);
or U1610 (N_1610,In_790,In_95);
nor U1611 (N_1611,In_1809,In_1815);
and U1612 (N_1612,In_1320,In_403);
or U1613 (N_1613,In_1744,In_1308);
xnor U1614 (N_1614,In_1280,In_943);
nand U1615 (N_1615,In_331,In_545);
nor U1616 (N_1616,In_1903,In_946);
and U1617 (N_1617,In_319,In_1616);
or U1618 (N_1618,In_1638,In_676);
nor U1619 (N_1619,In_346,In_4);
or U1620 (N_1620,In_1831,In_47);
nand U1621 (N_1621,In_1412,In_397);
or U1622 (N_1622,In_515,In_131);
nand U1623 (N_1623,In_1596,In_933);
nor U1624 (N_1624,In_811,In_1126);
and U1625 (N_1625,In_74,In_702);
nand U1626 (N_1626,In_1348,In_1054);
or U1627 (N_1627,In_1679,In_1410);
nor U1628 (N_1628,In_1341,In_1660);
or U1629 (N_1629,In_1001,In_333);
and U1630 (N_1630,In_138,In_367);
xor U1631 (N_1631,In_983,In_1005);
xor U1632 (N_1632,In_1516,In_1799);
or U1633 (N_1633,In_187,In_636);
nor U1634 (N_1634,In_936,In_728);
xor U1635 (N_1635,In_781,In_610);
xnor U1636 (N_1636,In_210,In_490);
nand U1637 (N_1637,In_878,In_398);
and U1638 (N_1638,In_1306,In_1550);
xor U1639 (N_1639,In_1064,In_1945);
or U1640 (N_1640,In_595,In_870);
and U1641 (N_1641,In_2,In_1153);
and U1642 (N_1642,In_150,In_1109);
nand U1643 (N_1643,In_301,In_1728);
nor U1644 (N_1644,In_1243,In_848);
xnor U1645 (N_1645,In_1963,In_1185);
and U1646 (N_1646,In_972,In_1025);
nand U1647 (N_1647,In_352,In_1012);
nor U1648 (N_1648,In_926,In_397);
nand U1649 (N_1649,In_303,In_760);
and U1650 (N_1650,In_707,In_1957);
xnor U1651 (N_1651,In_860,In_1592);
nand U1652 (N_1652,In_1099,In_997);
and U1653 (N_1653,In_282,In_348);
xnor U1654 (N_1654,In_1405,In_475);
and U1655 (N_1655,In_1214,In_221);
xor U1656 (N_1656,In_666,In_769);
xor U1657 (N_1657,In_179,In_188);
nand U1658 (N_1658,In_1589,In_1360);
or U1659 (N_1659,In_430,In_211);
nand U1660 (N_1660,In_664,In_235);
xnor U1661 (N_1661,In_1845,In_997);
and U1662 (N_1662,In_1704,In_65);
or U1663 (N_1663,In_1225,In_1741);
nand U1664 (N_1664,In_1522,In_1715);
and U1665 (N_1665,In_463,In_730);
nand U1666 (N_1666,In_1725,In_1607);
nor U1667 (N_1667,In_1670,In_1192);
and U1668 (N_1668,In_1721,In_113);
nand U1669 (N_1669,In_831,In_1644);
or U1670 (N_1670,In_772,In_283);
nor U1671 (N_1671,In_1358,In_1447);
nand U1672 (N_1672,In_99,In_712);
or U1673 (N_1673,In_840,In_1679);
xnor U1674 (N_1674,In_155,In_1836);
xnor U1675 (N_1675,In_82,In_734);
nor U1676 (N_1676,In_522,In_207);
nor U1677 (N_1677,In_1242,In_438);
nor U1678 (N_1678,In_405,In_1454);
xor U1679 (N_1679,In_882,In_818);
nor U1680 (N_1680,In_323,In_862);
xnor U1681 (N_1681,In_1124,In_1406);
or U1682 (N_1682,In_845,In_1191);
xnor U1683 (N_1683,In_1313,In_654);
or U1684 (N_1684,In_1548,In_1022);
or U1685 (N_1685,In_1223,In_308);
or U1686 (N_1686,In_359,In_981);
or U1687 (N_1687,In_468,In_698);
xor U1688 (N_1688,In_134,In_514);
and U1689 (N_1689,In_1309,In_791);
nand U1690 (N_1690,In_8,In_499);
and U1691 (N_1691,In_349,In_1818);
xnor U1692 (N_1692,In_1920,In_69);
or U1693 (N_1693,In_777,In_1646);
xor U1694 (N_1694,In_353,In_321);
nor U1695 (N_1695,In_15,In_145);
nand U1696 (N_1696,In_640,In_1243);
and U1697 (N_1697,In_856,In_7);
nor U1698 (N_1698,In_1022,In_1795);
or U1699 (N_1699,In_673,In_1353);
and U1700 (N_1700,In_1474,In_272);
or U1701 (N_1701,In_782,In_897);
nor U1702 (N_1702,In_24,In_1280);
nand U1703 (N_1703,In_1734,In_337);
or U1704 (N_1704,In_87,In_337);
xor U1705 (N_1705,In_630,In_530);
or U1706 (N_1706,In_507,In_1165);
and U1707 (N_1707,In_829,In_1508);
and U1708 (N_1708,In_1542,In_1999);
nor U1709 (N_1709,In_1032,In_902);
nor U1710 (N_1710,In_947,In_1842);
xnor U1711 (N_1711,In_427,In_227);
nand U1712 (N_1712,In_168,In_328);
xnor U1713 (N_1713,In_145,In_815);
xor U1714 (N_1714,In_1739,In_1251);
nor U1715 (N_1715,In_865,In_1861);
or U1716 (N_1716,In_560,In_1046);
nor U1717 (N_1717,In_1887,In_761);
or U1718 (N_1718,In_443,In_1257);
or U1719 (N_1719,In_13,In_904);
or U1720 (N_1720,In_38,In_162);
xnor U1721 (N_1721,In_1900,In_1885);
xnor U1722 (N_1722,In_1558,In_800);
xnor U1723 (N_1723,In_1712,In_446);
nor U1724 (N_1724,In_678,In_1666);
and U1725 (N_1725,In_1203,In_1053);
nand U1726 (N_1726,In_365,In_1080);
nand U1727 (N_1727,In_737,In_1451);
xor U1728 (N_1728,In_406,In_1105);
nand U1729 (N_1729,In_316,In_499);
nand U1730 (N_1730,In_416,In_1193);
or U1731 (N_1731,In_419,In_1450);
or U1732 (N_1732,In_35,In_1895);
or U1733 (N_1733,In_811,In_316);
or U1734 (N_1734,In_766,In_132);
and U1735 (N_1735,In_1186,In_1712);
xnor U1736 (N_1736,In_48,In_912);
nand U1737 (N_1737,In_950,In_402);
nand U1738 (N_1738,In_1884,In_1297);
nand U1739 (N_1739,In_1417,In_1812);
and U1740 (N_1740,In_1119,In_106);
and U1741 (N_1741,In_1384,In_699);
nand U1742 (N_1742,In_180,In_1690);
nand U1743 (N_1743,In_665,In_707);
nor U1744 (N_1744,In_129,In_871);
and U1745 (N_1745,In_297,In_33);
and U1746 (N_1746,In_1402,In_1815);
nor U1747 (N_1747,In_1621,In_1612);
nand U1748 (N_1748,In_673,In_291);
and U1749 (N_1749,In_1965,In_999);
xor U1750 (N_1750,In_833,In_951);
or U1751 (N_1751,In_1171,In_1572);
and U1752 (N_1752,In_662,In_565);
and U1753 (N_1753,In_1426,In_1180);
or U1754 (N_1754,In_1250,In_1819);
nor U1755 (N_1755,In_1172,In_464);
or U1756 (N_1756,In_1380,In_376);
nand U1757 (N_1757,In_190,In_635);
xnor U1758 (N_1758,In_600,In_1808);
nor U1759 (N_1759,In_1249,In_432);
xor U1760 (N_1760,In_1936,In_594);
nand U1761 (N_1761,In_282,In_1678);
or U1762 (N_1762,In_1744,In_26);
and U1763 (N_1763,In_82,In_892);
nor U1764 (N_1764,In_472,In_1160);
nand U1765 (N_1765,In_1548,In_1336);
nor U1766 (N_1766,In_644,In_959);
and U1767 (N_1767,In_1372,In_1380);
or U1768 (N_1768,In_549,In_520);
nand U1769 (N_1769,In_1119,In_1533);
and U1770 (N_1770,In_678,In_441);
nand U1771 (N_1771,In_991,In_1289);
nor U1772 (N_1772,In_461,In_579);
nor U1773 (N_1773,In_1432,In_138);
and U1774 (N_1774,In_304,In_594);
xor U1775 (N_1775,In_1146,In_1593);
and U1776 (N_1776,In_928,In_1085);
xor U1777 (N_1777,In_1266,In_1855);
xnor U1778 (N_1778,In_708,In_404);
nand U1779 (N_1779,In_1834,In_1376);
and U1780 (N_1780,In_756,In_640);
xor U1781 (N_1781,In_1898,In_1869);
nor U1782 (N_1782,In_1846,In_36);
or U1783 (N_1783,In_544,In_118);
nor U1784 (N_1784,In_721,In_271);
and U1785 (N_1785,In_1090,In_652);
nand U1786 (N_1786,In_1380,In_1203);
or U1787 (N_1787,In_879,In_1902);
or U1788 (N_1788,In_418,In_1766);
nand U1789 (N_1789,In_301,In_922);
xor U1790 (N_1790,In_771,In_1992);
or U1791 (N_1791,In_618,In_1519);
nand U1792 (N_1792,In_536,In_412);
xnor U1793 (N_1793,In_1597,In_890);
nor U1794 (N_1794,In_1656,In_1774);
nor U1795 (N_1795,In_40,In_334);
xnor U1796 (N_1796,In_308,In_714);
and U1797 (N_1797,In_447,In_1518);
and U1798 (N_1798,In_700,In_86);
xor U1799 (N_1799,In_247,In_1881);
xnor U1800 (N_1800,In_788,In_1417);
xnor U1801 (N_1801,In_212,In_458);
and U1802 (N_1802,In_1645,In_1116);
nor U1803 (N_1803,In_1034,In_972);
nor U1804 (N_1804,In_374,In_718);
nor U1805 (N_1805,In_1202,In_1772);
xor U1806 (N_1806,In_1344,In_1220);
xnor U1807 (N_1807,In_397,In_604);
xor U1808 (N_1808,In_1707,In_1097);
nor U1809 (N_1809,In_1947,In_1230);
nand U1810 (N_1810,In_988,In_568);
xor U1811 (N_1811,In_1660,In_884);
and U1812 (N_1812,In_1510,In_1494);
or U1813 (N_1813,In_1828,In_289);
and U1814 (N_1814,In_1982,In_192);
and U1815 (N_1815,In_1825,In_89);
nor U1816 (N_1816,In_1550,In_898);
xnor U1817 (N_1817,In_311,In_220);
xnor U1818 (N_1818,In_1929,In_935);
or U1819 (N_1819,In_416,In_321);
or U1820 (N_1820,In_777,In_1747);
or U1821 (N_1821,In_250,In_998);
or U1822 (N_1822,In_1641,In_1706);
and U1823 (N_1823,In_1485,In_377);
nand U1824 (N_1824,In_1262,In_1537);
xnor U1825 (N_1825,In_1771,In_559);
or U1826 (N_1826,In_1074,In_312);
xnor U1827 (N_1827,In_1091,In_1995);
nand U1828 (N_1828,In_398,In_1808);
and U1829 (N_1829,In_1829,In_686);
or U1830 (N_1830,In_164,In_1410);
and U1831 (N_1831,In_1189,In_990);
xnor U1832 (N_1832,In_1075,In_1214);
xnor U1833 (N_1833,In_366,In_1737);
or U1834 (N_1834,In_863,In_1009);
nand U1835 (N_1835,In_1628,In_119);
nor U1836 (N_1836,In_1617,In_1719);
nor U1837 (N_1837,In_538,In_441);
xor U1838 (N_1838,In_1950,In_278);
xor U1839 (N_1839,In_1260,In_1307);
nand U1840 (N_1840,In_1269,In_1249);
nor U1841 (N_1841,In_171,In_1405);
xnor U1842 (N_1842,In_105,In_956);
or U1843 (N_1843,In_883,In_253);
nand U1844 (N_1844,In_832,In_1801);
nor U1845 (N_1845,In_391,In_184);
xor U1846 (N_1846,In_1060,In_925);
and U1847 (N_1847,In_35,In_1652);
nor U1848 (N_1848,In_1697,In_660);
or U1849 (N_1849,In_1956,In_801);
nor U1850 (N_1850,In_379,In_449);
xor U1851 (N_1851,In_1472,In_1895);
or U1852 (N_1852,In_614,In_1930);
nor U1853 (N_1853,In_1770,In_1570);
and U1854 (N_1854,In_1213,In_1750);
xor U1855 (N_1855,In_915,In_1743);
nor U1856 (N_1856,In_1665,In_150);
nor U1857 (N_1857,In_1360,In_188);
nand U1858 (N_1858,In_1358,In_1836);
nor U1859 (N_1859,In_1849,In_775);
nand U1860 (N_1860,In_1815,In_625);
nor U1861 (N_1861,In_1310,In_1064);
nand U1862 (N_1862,In_1489,In_1473);
nand U1863 (N_1863,In_1882,In_54);
or U1864 (N_1864,In_1890,In_1708);
nor U1865 (N_1865,In_1243,In_1540);
xnor U1866 (N_1866,In_1782,In_359);
or U1867 (N_1867,In_24,In_429);
nand U1868 (N_1868,In_1946,In_1261);
and U1869 (N_1869,In_725,In_1808);
nor U1870 (N_1870,In_843,In_702);
xnor U1871 (N_1871,In_707,In_215);
or U1872 (N_1872,In_756,In_1698);
or U1873 (N_1873,In_1724,In_1954);
nand U1874 (N_1874,In_589,In_1290);
nand U1875 (N_1875,In_478,In_987);
and U1876 (N_1876,In_889,In_1042);
nand U1877 (N_1877,In_1833,In_1772);
xor U1878 (N_1878,In_1967,In_1953);
and U1879 (N_1879,In_1245,In_307);
nor U1880 (N_1880,In_958,In_339);
nand U1881 (N_1881,In_372,In_1284);
and U1882 (N_1882,In_734,In_1519);
or U1883 (N_1883,In_689,In_814);
nor U1884 (N_1884,In_1894,In_658);
nand U1885 (N_1885,In_1877,In_747);
and U1886 (N_1886,In_696,In_1286);
or U1887 (N_1887,In_1822,In_1969);
and U1888 (N_1888,In_795,In_1725);
nand U1889 (N_1889,In_1205,In_686);
or U1890 (N_1890,In_972,In_463);
nand U1891 (N_1891,In_1754,In_980);
or U1892 (N_1892,In_252,In_574);
xnor U1893 (N_1893,In_416,In_230);
or U1894 (N_1894,In_408,In_1897);
or U1895 (N_1895,In_1588,In_1465);
nand U1896 (N_1896,In_1398,In_513);
or U1897 (N_1897,In_548,In_1290);
nor U1898 (N_1898,In_1990,In_724);
nor U1899 (N_1899,In_1010,In_1326);
nand U1900 (N_1900,In_395,In_102);
xor U1901 (N_1901,In_880,In_573);
or U1902 (N_1902,In_270,In_1200);
nor U1903 (N_1903,In_179,In_109);
nand U1904 (N_1904,In_1423,In_1679);
and U1905 (N_1905,In_600,In_1181);
or U1906 (N_1906,In_205,In_1958);
and U1907 (N_1907,In_510,In_1802);
nand U1908 (N_1908,In_1341,In_1834);
or U1909 (N_1909,In_965,In_1395);
nor U1910 (N_1910,In_1640,In_1634);
or U1911 (N_1911,In_240,In_1340);
xnor U1912 (N_1912,In_231,In_267);
nand U1913 (N_1913,In_1286,In_1616);
nor U1914 (N_1914,In_1959,In_89);
and U1915 (N_1915,In_88,In_446);
and U1916 (N_1916,In_1702,In_171);
or U1917 (N_1917,In_1144,In_714);
xor U1918 (N_1918,In_1432,In_87);
or U1919 (N_1919,In_524,In_1945);
nor U1920 (N_1920,In_888,In_18);
nand U1921 (N_1921,In_1208,In_381);
nand U1922 (N_1922,In_1306,In_1452);
xor U1923 (N_1923,In_178,In_1451);
nor U1924 (N_1924,In_479,In_97);
or U1925 (N_1925,In_1127,In_1777);
nor U1926 (N_1926,In_1461,In_1417);
or U1927 (N_1927,In_145,In_1424);
and U1928 (N_1928,In_1941,In_1408);
xor U1929 (N_1929,In_1075,In_1782);
or U1930 (N_1930,In_697,In_967);
nand U1931 (N_1931,In_1739,In_446);
and U1932 (N_1932,In_462,In_644);
and U1933 (N_1933,In_626,In_1189);
and U1934 (N_1934,In_749,In_1310);
or U1935 (N_1935,In_1398,In_306);
and U1936 (N_1936,In_235,In_1118);
nor U1937 (N_1937,In_1072,In_1451);
or U1938 (N_1938,In_1639,In_514);
nor U1939 (N_1939,In_702,In_348);
nor U1940 (N_1940,In_985,In_994);
or U1941 (N_1941,In_1994,In_978);
nor U1942 (N_1942,In_1210,In_978);
or U1943 (N_1943,In_134,In_322);
or U1944 (N_1944,In_1405,In_743);
or U1945 (N_1945,In_98,In_758);
or U1946 (N_1946,In_349,In_138);
nand U1947 (N_1947,In_759,In_185);
and U1948 (N_1948,In_515,In_110);
nor U1949 (N_1949,In_635,In_1356);
and U1950 (N_1950,In_939,In_321);
nand U1951 (N_1951,In_732,In_832);
xnor U1952 (N_1952,In_487,In_1593);
nor U1953 (N_1953,In_1346,In_371);
and U1954 (N_1954,In_1839,In_1478);
xor U1955 (N_1955,In_1187,In_843);
nand U1956 (N_1956,In_1162,In_1011);
xor U1957 (N_1957,In_1769,In_484);
and U1958 (N_1958,In_1590,In_1899);
xor U1959 (N_1959,In_1614,In_292);
and U1960 (N_1960,In_1434,In_1498);
or U1961 (N_1961,In_749,In_479);
nand U1962 (N_1962,In_267,In_852);
xnor U1963 (N_1963,In_1072,In_1667);
nor U1964 (N_1964,In_642,In_215);
nand U1965 (N_1965,In_1288,In_1567);
nor U1966 (N_1966,In_299,In_707);
nand U1967 (N_1967,In_1784,In_755);
or U1968 (N_1968,In_841,In_292);
or U1969 (N_1969,In_1484,In_1042);
and U1970 (N_1970,In_689,In_752);
nand U1971 (N_1971,In_1192,In_858);
and U1972 (N_1972,In_764,In_330);
nor U1973 (N_1973,In_538,In_342);
nor U1974 (N_1974,In_575,In_446);
and U1975 (N_1975,In_86,In_1995);
and U1976 (N_1976,In_498,In_1998);
nand U1977 (N_1977,In_1246,In_1464);
and U1978 (N_1978,In_1485,In_822);
and U1979 (N_1979,In_768,In_1272);
nor U1980 (N_1980,In_1288,In_1963);
or U1981 (N_1981,In_453,In_495);
xnor U1982 (N_1982,In_1778,In_699);
xor U1983 (N_1983,In_316,In_139);
xor U1984 (N_1984,In_984,In_1750);
xnor U1985 (N_1985,In_25,In_105);
and U1986 (N_1986,In_413,In_1811);
xnor U1987 (N_1987,In_490,In_189);
nand U1988 (N_1988,In_865,In_1011);
and U1989 (N_1989,In_332,In_935);
nand U1990 (N_1990,In_1937,In_1194);
nor U1991 (N_1991,In_1981,In_279);
xor U1992 (N_1992,In_1436,In_491);
nor U1993 (N_1993,In_898,In_1826);
or U1994 (N_1994,In_1524,In_452);
and U1995 (N_1995,In_593,In_919);
nand U1996 (N_1996,In_54,In_1899);
or U1997 (N_1997,In_1553,In_55);
nand U1998 (N_1998,In_1873,In_1915);
xnor U1999 (N_1999,In_467,In_1836);
and U2000 (N_2000,In_1972,In_433);
or U2001 (N_2001,In_1862,In_1441);
nand U2002 (N_2002,In_437,In_1809);
and U2003 (N_2003,In_1780,In_1069);
xor U2004 (N_2004,In_1405,In_1099);
xnor U2005 (N_2005,In_1239,In_1255);
xnor U2006 (N_2006,In_970,In_307);
nand U2007 (N_2007,In_1204,In_1568);
xnor U2008 (N_2008,In_923,In_1136);
nor U2009 (N_2009,In_1274,In_1218);
nand U2010 (N_2010,In_706,In_845);
and U2011 (N_2011,In_605,In_665);
and U2012 (N_2012,In_1310,In_564);
and U2013 (N_2013,In_925,In_221);
xor U2014 (N_2014,In_33,In_256);
and U2015 (N_2015,In_115,In_70);
and U2016 (N_2016,In_597,In_1042);
nor U2017 (N_2017,In_438,In_367);
or U2018 (N_2018,In_223,In_1701);
xnor U2019 (N_2019,In_339,In_1300);
and U2020 (N_2020,In_580,In_1701);
nor U2021 (N_2021,In_1238,In_637);
xnor U2022 (N_2022,In_1273,In_224);
nand U2023 (N_2023,In_260,In_142);
nor U2024 (N_2024,In_1154,In_68);
or U2025 (N_2025,In_1075,In_848);
nor U2026 (N_2026,In_1575,In_1196);
nand U2027 (N_2027,In_960,In_1763);
nor U2028 (N_2028,In_936,In_1619);
xor U2029 (N_2029,In_260,In_5);
or U2030 (N_2030,In_973,In_1005);
nor U2031 (N_2031,In_594,In_90);
or U2032 (N_2032,In_810,In_847);
xnor U2033 (N_2033,In_1857,In_1220);
or U2034 (N_2034,In_1327,In_1162);
xnor U2035 (N_2035,In_591,In_301);
xor U2036 (N_2036,In_0,In_1311);
xnor U2037 (N_2037,In_1894,In_504);
and U2038 (N_2038,In_680,In_389);
nor U2039 (N_2039,In_324,In_427);
and U2040 (N_2040,In_1838,In_1441);
and U2041 (N_2041,In_421,In_830);
xnor U2042 (N_2042,In_962,In_839);
nor U2043 (N_2043,In_1100,In_91);
nand U2044 (N_2044,In_266,In_702);
nor U2045 (N_2045,In_1233,In_618);
and U2046 (N_2046,In_1623,In_1810);
xor U2047 (N_2047,In_1103,In_577);
xnor U2048 (N_2048,In_146,In_1053);
nand U2049 (N_2049,In_46,In_1158);
and U2050 (N_2050,In_1993,In_1170);
and U2051 (N_2051,In_963,In_694);
or U2052 (N_2052,In_710,In_1860);
nand U2053 (N_2053,In_1684,In_358);
or U2054 (N_2054,In_405,In_680);
nand U2055 (N_2055,In_544,In_618);
or U2056 (N_2056,In_468,In_1046);
nor U2057 (N_2057,In_941,In_1100);
xnor U2058 (N_2058,In_1370,In_960);
and U2059 (N_2059,In_1705,In_424);
xor U2060 (N_2060,In_826,In_706);
and U2061 (N_2061,In_637,In_1837);
nand U2062 (N_2062,In_1550,In_1979);
nand U2063 (N_2063,In_1465,In_504);
xor U2064 (N_2064,In_1510,In_1079);
nor U2065 (N_2065,In_1831,In_111);
xor U2066 (N_2066,In_1194,In_1189);
nand U2067 (N_2067,In_1415,In_754);
and U2068 (N_2068,In_750,In_626);
nand U2069 (N_2069,In_796,In_1683);
xnor U2070 (N_2070,In_826,In_3);
or U2071 (N_2071,In_4,In_1214);
and U2072 (N_2072,In_891,In_335);
and U2073 (N_2073,In_712,In_1629);
nor U2074 (N_2074,In_811,In_535);
or U2075 (N_2075,In_1692,In_1292);
nand U2076 (N_2076,In_1431,In_1044);
nor U2077 (N_2077,In_1625,In_1308);
or U2078 (N_2078,In_1263,In_125);
nand U2079 (N_2079,In_683,In_1637);
xnor U2080 (N_2080,In_1884,In_1584);
nand U2081 (N_2081,In_770,In_1504);
xnor U2082 (N_2082,In_1472,In_177);
and U2083 (N_2083,In_806,In_35);
nand U2084 (N_2084,In_665,In_736);
nor U2085 (N_2085,In_734,In_72);
xnor U2086 (N_2086,In_603,In_253);
and U2087 (N_2087,In_755,In_1171);
or U2088 (N_2088,In_435,In_530);
or U2089 (N_2089,In_873,In_1580);
nor U2090 (N_2090,In_1705,In_1303);
nor U2091 (N_2091,In_820,In_678);
and U2092 (N_2092,In_1001,In_1439);
nor U2093 (N_2093,In_1913,In_1648);
xor U2094 (N_2094,In_97,In_1877);
xnor U2095 (N_2095,In_533,In_451);
xor U2096 (N_2096,In_1901,In_562);
nand U2097 (N_2097,In_198,In_1174);
xor U2098 (N_2098,In_193,In_903);
and U2099 (N_2099,In_1344,In_903);
and U2100 (N_2100,In_1723,In_1263);
or U2101 (N_2101,In_218,In_1319);
nor U2102 (N_2102,In_585,In_1004);
nand U2103 (N_2103,In_1005,In_299);
and U2104 (N_2104,In_876,In_1482);
nand U2105 (N_2105,In_632,In_1161);
nand U2106 (N_2106,In_1716,In_1341);
xnor U2107 (N_2107,In_1577,In_480);
xor U2108 (N_2108,In_258,In_1347);
xor U2109 (N_2109,In_1581,In_1258);
and U2110 (N_2110,In_578,In_874);
nor U2111 (N_2111,In_952,In_1562);
nand U2112 (N_2112,In_354,In_562);
nor U2113 (N_2113,In_1924,In_15);
nand U2114 (N_2114,In_1141,In_423);
nand U2115 (N_2115,In_845,In_622);
nand U2116 (N_2116,In_408,In_15);
nand U2117 (N_2117,In_730,In_437);
nand U2118 (N_2118,In_427,In_1480);
and U2119 (N_2119,In_211,In_311);
xnor U2120 (N_2120,In_505,In_185);
or U2121 (N_2121,In_1652,In_1169);
and U2122 (N_2122,In_1695,In_1836);
xnor U2123 (N_2123,In_514,In_1699);
nand U2124 (N_2124,In_1361,In_1589);
and U2125 (N_2125,In_309,In_684);
or U2126 (N_2126,In_1748,In_1689);
and U2127 (N_2127,In_942,In_274);
xnor U2128 (N_2128,In_1775,In_879);
xnor U2129 (N_2129,In_1242,In_526);
and U2130 (N_2130,In_746,In_875);
xor U2131 (N_2131,In_642,In_994);
xor U2132 (N_2132,In_1346,In_1208);
and U2133 (N_2133,In_148,In_1256);
xor U2134 (N_2134,In_648,In_179);
nand U2135 (N_2135,In_716,In_270);
xnor U2136 (N_2136,In_298,In_1105);
nor U2137 (N_2137,In_566,In_1019);
nand U2138 (N_2138,In_1106,In_1268);
nor U2139 (N_2139,In_23,In_1880);
or U2140 (N_2140,In_1708,In_547);
xnor U2141 (N_2141,In_210,In_1687);
xnor U2142 (N_2142,In_559,In_372);
nand U2143 (N_2143,In_329,In_1691);
nand U2144 (N_2144,In_314,In_1746);
nand U2145 (N_2145,In_1324,In_441);
nand U2146 (N_2146,In_1453,In_566);
or U2147 (N_2147,In_201,In_417);
xor U2148 (N_2148,In_1880,In_214);
or U2149 (N_2149,In_1818,In_1727);
or U2150 (N_2150,In_1647,In_1443);
or U2151 (N_2151,In_1912,In_579);
xnor U2152 (N_2152,In_177,In_1470);
xnor U2153 (N_2153,In_26,In_1425);
xnor U2154 (N_2154,In_782,In_469);
or U2155 (N_2155,In_73,In_934);
xnor U2156 (N_2156,In_334,In_1778);
nor U2157 (N_2157,In_20,In_788);
nand U2158 (N_2158,In_1010,In_1573);
or U2159 (N_2159,In_893,In_887);
or U2160 (N_2160,In_923,In_1770);
or U2161 (N_2161,In_691,In_1796);
nand U2162 (N_2162,In_911,In_591);
xnor U2163 (N_2163,In_307,In_897);
xnor U2164 (N_2164,In_979,In_1893);
nor U2165 (N_2165,In_764,In_124);
nand U2166 (N_2166,In_1594,In_287);
or U2167 (N_2167,In_747,In_1884);
and U2168 (N_2168,In_1848,In_765);
nand U2169 (N_2169,In_162,In_1450);
xnor U2170 (N_2170,In_417,In_625);
nand U2171 (N_2171,In_1466,In_413);
and U2172 (N_2172,In_296,In_1365);
xor U2173 (N_2173,In_918,In_243);
nor U2174 (N_2174,In_173,In_1595);
xnor U2175 (N_2175,In_1661,In_383);
and U2176 (N_2176,In_1154,In_1343);
xnor U2177 (N_2177,In_17,In_1814);
xnor U2178 (N_2178,In_1608,In_857);
nand U2179 (N_2179,In_1516,In_447);
and U2180 (N_2180,In_1869,In_336);
or U2181 (N_2181,In_266,In_1165);
xor U2182 (N_2182,In_841,In_1767);
xor U2183 (N_2183,In_249,In_1092);
nand U2184 (N_2184,In_158,In_1671);
nor U2185 (N_2185,In_104,In_1438);
or U2186 (N_2186,In_174,In_859);
nand U2187 (N_2187,In_1566,In_1129);
nand U2188 (N_2188,In_1214,In_1466);
or U2189 (N_2189,In_374,In_884);
or U2190 (N_2190,In_704,In_1138);
and U2191 (N_2191,In_1518,In_1031);
nand U2192 (N_2192,In_1422,In_565);
nor U2193 (N_2193,In_1569,In_1998);
nor U2194 (N_2194,In_1384,In_995);
xor U2195 (N_2195,In_1869,In_178);
and U2196 (N_2196,In_1884,In_117);
nand U2197 (N_2197,In_1157,In_1492);
and U2198 (N_2198,In_193,In_852);
nand U2199 (N_2199,In_1678,In_55);
or U2200 (N_2200,In_1317,In_1345);
xnor U2201 (N_2201,In_114,In_643);
nand U2202 (N_2202,In_788,In_495);
and U2203 (N_2203,In_997,In_538);
nand U2204 (N_2204,In_932,In_472);
nor U2205 (N_2205,In_484,In_1423);
and U2206 (N_2206,In_1409,In_714);
nand U2207 (N_2207,In_355,In_314);
or U2208 (N_2208,In_1929,In_1658);
nor U2209 (N_2209,In_1776,In_502);
and U2210 (N_2210,In_1975,In_691);
and U2211 (N_2211,In_1589,In_1532);
and U2212 (N_2212,In_864,In_897);
or U2213 (N_2213,In_828,In_1880);
or U2214 (N_2214,In_1277,In_1995);
nand U2215 (N_2215,In_236,In_489);
and U2216 (N_2216,In_1174,In_238);
nor U2217 (N_2217,In_1666,In_293);
or U2218 (N_2218,In_894,In_228);
nor U2219 (N_2219,In_1935,In_500);
nand U2220 (N_2220,In_1469,In_1414);
nor U2221 (N_2221,In_184,In_1512);
xnor U2222 (N_2222,In_1952,In_1209);
xor U2223 (N_2223,In_14,In_1424);
or U2224 (N_2224,In_1507,In_47);
xnor U2225 (N_2225,In_1589,In_558);
xor U2226 (N_2226,In_573,In_1886);
nand U2227 (N_2227,In_1565,In_1458);
nor U2228 (N_2228,In_1731,In_1065);
nand U2229 (N_2229,In_1952,In_245);
or U2230 (N_2230,In_1356,In_381);
or U2231 (N_2231,In_759,In_1381);
or U2232 (N_2232,In_467,In_942);
nand U2233 (N_2233,In_2,In_1332);
xor U2234 (N_2234,In_1863,In_683);
and U2235 (N_2235,In_1791,In_1221);
nor U2236 (N_2236,In_1160,In_989);
or U2237 (N_2237,In_933,In_968);
nor U2238 (N_2238,In_583,In_1277);
or U2239 (N_2239,In_55,In_609);
xor U2240 (N_2240,In_661,In_1961);
and U2241 (N_2241,In_1404,In_1876);
and U2242 (N_2242,In_1313,In_1815);
and U2243 (N_2243,In_457,In_1894);
and U2244 (N_2244,In_257,In_1248);
or U2245 (N_2245,In_299,In_856);
nor U2246 (N_2246,In_146,In_1715);
xnor U2247 (N_2247,In_1367,In_167);
nor U2248 (N_2248,In_455,In_166);
nand U2249 (N_2249,In_575,In_1175);
or U2250 (N_2250,In_128,In_269);
and U2251 (N_2251,In_52,In_207);
nand U2252 (N_2252,In_163,In_126);
nor U2253 (N_2253,In_263,In_869);
nor U2254 (N_2254,In_1085,In_1451);
and U2255 (N_2255,In_1502,In_1009);
xor U2256 (N_2256,In_1987,In_1353);
nand U2257 (N_2257,In_1928,In_1995);
nor U2258 (N_2258,In_934,In_1763);
nor U2259 (N_2259,In_1381,In_1471);
or U2260 (N_2260,In_988,In_1694);
xor U2261 (N_2261,In_189,In_1344);
nand U2262 (N_2262,In_870,In_1949);
or U2263 (N_2263,In_753,In_1345);
nor U2264 (N_2264,In_1388,In_130);
and U2265 (N_2265,In_1753,In_659);
or U2266 (N_2266,In_471,In_1867);
xnor U2267 (N_2267,In_785,In_797);
nor U2268 (N_2268,In_258,In_969);
and U2269 (N_2269,In_1818,In_1150);
nand U2270 (N_2270,In_1628,In_524);
nor U2271 (N_2271,In_1594,In_600);
nand U2272 (N_2272,In_837,In_1381);
nand U2273 (N_2273,In_1963,In_701);
and U2274 (N_2274,In_450,In_758);
or U2275 (N_2275,In_1122,In_735);
xnor U2276 (N_2276,In_272,In_1499);
nor U2277 (N_2277,In_1945,In_1853);
and U2278 (N_2278,In_1921,In_1183);
and U2279 (N_2279,In_554,In_1515);
or U2280 (N_2280,In_715,In_718);
nand U2281 (N_2281,In_1179,In_1398);
xor U2282 (N_2282,In_1705,In_762);
xnor U2283 (N_2283,In_1179,In_1127);
nand U2284 (N_2284,In_642,In_202);
or U2285 (N_2285,In_351,In_1794);
xnor U2286 (N_2286,In_315,In_1386);
and U2287 (N_2287,In_1575,In_1927);
nor U2288 (N_2288,In_537,In_110);
nor U2289 (N_2289,In_1378,In_1937);
xnor U2290 (N_2290,In_807,In_899);
and U2291 (N_2291,In_1715,In_94);
nor U2292 (N_2292,In_1618,In_1279);
and U2293 (N_2293,In_269,In_1617);
or U2294 (N_2294,In_1358,In_1314);
and U2295 (N_2295,In_458,In_1106);
xnor U2296 (N_2296,In_1481,In_993);
xor U2297 (N_2297,In_878,In_845);
nor U2298 (N_2298,In_1955,In_1051);
nor U2299 (N_2299,In_1709,In_1230);
xnor U2300 (N_2300,In_1249,In_739);
nor U2301 (N_2301,In_523,In_1909);
and U2302 (N_2302,In_620,In_1204);
and U2303 (N_2303,In_1824,In_1893);
xnor U2304 (N_2304,In_370,In_1278);
or U2305 (N_2305,In_1142,In_1058);
or U2306 (N_2306,In_1034,In_802);
nor U2307 (N_2307,In_142,In_1122);
xnor U2308 (N_2308,In_1415,In_1935);
or U2309 (N_2309,In_821,In_1005);
and U2310 (N_2310,In_118,In_1771);
nor U2311 (N_2311,In_608,In_1376);
nand U2312 (N_2312,In_1775,In_764);
or U2313 (N_2313,In_412,In_1396);
xnor U2314 (N_2314,In_392,In_954);
or U2315 (N_2315,In_1626,In_146);
and U2316 (N_2316,In_1347,In_1829);
nor U2317 (N_2317,In_938,In_236);
or U2318 (N_2318,In_1691,In_1666);
xor U2319 (N_2319,In_1233,In_1766);
nor U2320 (N_2320,In_544,In_838);
nand U2321 (N_2321,In_978,In_1934);
or U2322 (N_2322,In_536,In_1959);
xor U2323 (N_2323,In_1009,In_662);
nand U2324 (N_2324,In_206,In_1006);
nand U2325 (N_2325,In_1440,In_1463);
and U2326 (N_2326,In_122,In_933);
nor U2327 (N_2327,In_504,In_1414);
or U2328 (N_2328,In_1038,In_1755);
xnor U2329 (N_2329,In_1046,In_716);
nand U2330 (N_2330,In_1225,In_1840);
xor U2331 (N_2331,In_1776,In_1479);
xnor U2332 (N_2332,In_88,In_283);
nor U2333 (N_2333,In_1694,In_1441);
nand U2334 (N_2334,In_887,In_1759);
nor U2335 (N_2335,In_1372,In_1697);
or U2336 (N_2336,In_807,In_1000);
xnor U2337 (N_2337,In_1092,In_365);
nand U2338 (N_2338,In_718,In_397);
nor U2339 (N_2339,In_1243,In_376);
nand U2340 (N_2340,In_1874,In_478);
nor U2341 (N_2341,In_1189,In_1475);
or U2342 (N_2342,In_1832,In_219);
and U2343 (N_2343,In_1770,In_1815);
xnor U2344 (N_2344,In_1646,In_339);
nand U2345 (N_2345,In_885,In_533);
and U2346 (N_2346,In_817,In_995);
nand U2347 (N_2347,In_1052,In_822);
and U2348 (N_2348,In_1755,In_1118);
and U2349 (N_2349,In_1627,In_752);
xor U2350 (N_2350,In_1416,In_136);
nand U2351 (N_2351,In_1227,In_288);
or U2352 (N_2352,In_585,In_1653);
and U2353 (N_2353,In_429,In_27);
nor U2354 (N_2354,In_915,In_613);
nand U2355 (N_2355,In_724,In_1018);
nand U2356 (N_2356,In_443,In_1074);
nor U2357 (N_2357,In_1616,In_896);
nand U2358 (N_2358,In_1176,In_923);
nand U2359 (N_2359,In_981,In_1309);
nor U2360 (N_2360,In_1488,In_1792);
nor U2361 (N_2361,In_450,In_1402);
nand U2362 (N_2362,In_947,In_295);
and U2363 (N_2363,In_153,In_1886);
and U2364 (N_2364,In_1528,In_1080);
xor U2365 (N_2365,In_1412,In_994);
nand U2366 (N_2366,In_563,In_1036);
and U2367 (N_2367,In_1307,In_1450);
nand U2368 (N_2368,In_1990,In_40);
xor U2369 (N_2369,In_739,In_1857);
nor U2370 (N_2370,In_1729,In_806);
nor U2371 (N_2371,In_137,In_1822);
nand U2372 (N_2372,In_246,In_1911);
nor U2373 (N_2373,In_1663,In_1572);
and U2374 (N_2374,In_1754,In_1601);
nor U2375 (N_2375,In_311,In_361);
nor U2376 (N_2376,In_49,In_823);
and U2377 (N_2377,In_1290,In_1882);
nand U2378 (N_2378,In_717,In_1983);
or U2379 (N_2379,In_1149,In_999);
nand U2380 (N_2380,In_730,In_296);
nand U2381 (N_2381,In_864,In_518);
nand U2382 (N_2382,In_1924,In_274);
xnor U2383 (N_2383,In_138,In_1511);
and U2384 (N_2384,In_1466,In_914);
nand U2385 (N_2385,In_1601,In_1634);
or U2386 (N_2386,In_1515,In_1168);
nor U2387 (N_2387,In_1996,In_195);
nand U2388 (N_2388,In_10,In_160);
or U2389 (N_2389,In_259,In_1399);
xor U2390 (N_2390,In_1026,In_1181);
or U2391 (N_2391,In_1997,In_1563);
or U2392 (N_2392,In_1141,In_853);
nand U2393 (N_2393,In_555,In_212);
and U2394 (N_2394,In_714,In_1695);
xnor U2395 (N_2395,In_1368,In_1087);
or U2396 (N_2396,In_1295,In_1943);
nor U2397 (N_2397,In_542,In_1495);
xor U2398 (N_2398,In_1829,In_1109);
xnor U2399 (N_2399,In_518,In_146);
and U2400 (N_2400,In_1161,In_200);
nor U2401 (N_2401,In_1739,In_902);
or U2402 (N_2402,In_1198,In_608);
nand U2403 (N_2403,In_1955,In_1415);
nor U2404 (N_2404,In_769,In_746);
and U2405 (N_2405,In_1678,In_630);
nand U2406 (N_2406,In_1264,In_1059);
or U2407 (N_2407,In_1469,In_857);
xnor U2408 (N_2408,In_604,In_733);
and U2409 (N_2409,In_1998,In_1193);
nor U2410 (N_2410,In_1818,In_921);
xor U2411 (N_2411,In_1191,In_1996);
nor U2412 (N_2412,In_1406,In_1163);
and U2413 (N_2413,In_485,In_1262);
or U2414 (N_2414,In_243,In_747);
or U2415 (N_2415,In_1355,In_326);
nand U2416 (N_2416,In_101,In_1487);
nand U2417 (N_2417,In_1500,In_290);
nand U2418 (N_2418,In_1359,In_1401);
and U2419 (N_2419,In_337,In_1406);
nor U2420 (N_2420,In_1851,In_192);
and U2421 (N_2421,In_875,In_1194);
nor U2422 (N_2422,In_1910,In_1302);
nor U2423 (N_2423,In_314,In_53);
or U2424 (N_2424,In_1206,In_134);
xor U2425 (N_2425,In_1288,In_839);
nor U2426 (N_2426,In_31,In_345);
and U2427 (N_2427,In_97,In_1317);
nand U2428 (N_2428,In_1071,In_1207);
xor U2429 (N_2429,In_832,In_576);
nor U2430 (N_2430,In_317,In_1566);
nand U2431 (N_2431,In_1760,In_439);
nor U2432 (N_2432,In_700,In_1957);
and U2433 (N_2433,In_104,In_1195);
or U2434 (N_2434,In_1839,In_1179);
or U2435 (N_2435,In_533,In_1827);
nor U2436 (N_2436,In_723,In_1780);
and U2437 (N_2437,In_1344,In_934);
xor U2438 (N_2438,In_606,In_90);
nor U2439 (N_2439,In_931,In_983);
xor U2440 (N_2440,In_1718,In_789);
nor U2441 (N_2441,In_1688,In_1241);
nand U2442 (N_2442,In_1366,In_840);
or U2443 (N_2443,In_659,In_152);
and U2444 (N_2444,In_313,In_400);
and U2445 (N_2445,In_1104,In_953);
xnor U2446 (N_2446,In_190,In_102);
and U2447 (N_2447,In_1328,In_1935);
nor U2448 (N_2448,In_693,In_1606);
nor U2449 (N_2449,In_1316,In_1156);
xnor U2450 (N_2450,In_49,In_1674);
or U2451 (N_2451,In_1413,In_32);
nor U2452 (N_2452,In_1417,In_1458);
nor U2453 (N_2453,In_1853,In_1574);
nor U2454 (N_2454,In_1132,In_1571);
nand U2455 (N_2455,In_941,In_1530);
xnor U2456 (N_2456,In_920,In_849);
nor U2457 (N_2457,In_761,In_869);
xnor U2458 (N_2458,In_1478,In_204);
xor U2459 (N_2459,In_1278,In_979);
or U2460 (N_2460,In_118,In_619);
nand U2461 (N_2461,In_312,In_1188);
nor U2462 (N_2462,In_1664,In_1268);
nand U2463 (N_2463,In_1232,In_708);
nand U2464 (N_2464,In_190,In_1353);
nor U2465 (N_2465,In_1204,In_796);
and U2466 (N_2466,In_1932,In_1339);
nand U2467 (N_2467,In_1918,In_110);
or U2468 (N_2468,In_1041,In_1433);
and U2469 (N_2469,In_743,In_1852);
nand U2470 (N_2470,In_280,In_1662);
nand U2471 (N_2471,In_648,In_135);
or U2472 (N_2472,In_1298,In_522);
nor U2473 (N_2473,In_1716,In_509);
xnor U2474 (N_2474,In_1652,In_820);
or U2475 (N_2475,In_970,In_1557);
and U2476 (N_2476,In_1335,In_1234);
or U2477 (N_2477,In_44,In_556);
xnor U2478 (N_2478,In_1322,In_1986);
xor U2479 (N_2479,In_1545,In_1674);
nand U2480 (N_2480,In_1962,In_628);
nand U2481 (N_2481,In_371,In_1445);
or U2482 (N_2482,In_1747,In_273);
or U2483 (N_2483,In_120,In_787);
nor U2484 (N_2484,In_1820,In_1872);
nand U2485 (N_2485,In_1977,In_1141);
nor U2486 (N_2486,In_1934,In_1737);
or U2487 (N_2487,In_780,In_37);
nand U2488 (N_2488,In_698,In_158);
xor U2489 (N_2489,In_1635,In_1691);
and U2490 (N_2490,In_131,In_1587);
xnor U2491 (N_2491,In_1363,In_1236);
nor U2492 (N_2492,In_491,In_550);
nand U2493 (N_2493,In_576,In_404);
xnor U2494 (N_2494,In_332,In_231);
xnor U2495 (N_2495,In_647,In_1300);
xor U2496 (N_2496,In_1152,In_1605);
or U2497 (N_2497,In_1443,In_1613);
and U2498 (N_2498,In_1226,In_436);
or U2499 (N_2499,In_867,In_407);
nor U2500 (N_2500,In_545,In_345);
or U2501 (N_2501,In_32,In_1842);
xor U2502 (N_2502,In_807,In_1750);
or U2503 (N_2503,In_692,In_684);
or U2504 (N_2504,In_737,In_1784);
and U2505 (N_2505,In_4,In_270);
or U2506 (N_2506,In_1734,In_833);
or U2507 (N_2507,In_1163,In_968);
or U2508 (N_2508,In_620,In_1104);
nor U2509 (N_2509,In_1689,In_1090);
nand U2510 (N_2510,In_104,In_1056);
nor U2511 (N_2511,In_1001,In_1400);
xnor U2512 (N_2512,In_1643,In_1526);
and U2513 (N_2513,In_1224,In_1418);
nand U2514 (N_2514,In_137,In_1119);
or U2515 (N_2515,In_223,In_685);
xnor U2516 (N_2516,In_1157,In_1396);
xnor U2517 (N_2517,In_1432,In_493);
nand U2518 (N_2518,In_734,In_1268);
nand U2519 (N_2519,In_169,In_1998);
or U2520 (N_2520,In_1643,In_942);
xnor U2521 (N_2521,In_438,In_942);
xor U2522 (N_2522,In_604,In_725);
and U2523 (N_2523,In_422,In_192);
xnor U2524 (N_2524,In_535,In_1008);
nand U2525 (N_2525,In_1739,In_1181);
nand U2526 (N_2526,In_43,In_1756);
xor U2527 (N_2527,In_1628,In_449);
nor U2528 (N_2528,In_505,In_1839);
or U2529 (N_2529,In_0,In_1972);
nor U2530 (N_2530,In_1931,In_736);
xnor U2531 (N_2531,In_945,In_1376);
nor U2532 (N_2532,In_704,In_1152);
or U2533 (N_2533,In_301,In_51);
xor U2534 (N_2534,In_99,In_1559);
xor U2535 (N_2535,In_501,In_1556);
nand U2536 (N_2536,In_1492,In_7);
xor U2537 (N_2537,In_1272,In_362);
and U2538 (N_2538,In_160,In_59);
or U2539 (N_2539,In_1245,In_389);
and U2540 (N_2540,In_1986,In_1392);
xor U2541 (N_2541,In_1967,In_1706);
xnor U2542 (N_2542,In_914,In_7);
nand U2543 (N_2543,In_1812,In_809);
nand U2544 (N_2544,In_448,In_216);
nand U2545 (N_2545,In_21,In_1112);
xnor U2546 (N_2546,In_594,In_763);
xnor U2547 (N_2547,In_1155,In_1699);
and U2548 (N_2548,In_1046,In_1983);
nand U2549 (N_2549,In_1795,In_1234);
xnor U2550 (N_2550,In_1282,In_1266);
nor U2551 (N_2551,In_1480,In_738);
and U2552 (N_2552,In_1055,In_144);
xnor U2553 (N_2553,In_327,In_1786);
nor U2554 (N_2554,In_1081,In_1697);
and U2555 (N_2555,In_885,In_646);
or U2556 (N_2556,In_1129,In_1511);
or U2557 (N_2557,In_1195,In_1091);
nor U2558 (N_2558,In_1369,In_1539);
or U2559 (N_2559,In_218,In_624);
or U2560 (N_2560,In_1739,In_1918);
nor U2561 (N_2561,In_712,In_44);
xnor U2562 (N_2562,In_708,In_586);
nor U2563 (N_2563,In_1482,In_1723);
nor U2564 (N_2564,In_1727,In_1895);
nand U2565 (N_2565,In_1978,In_719);
and U2566 (N_2566,In_1880,In_979);
xnor U2567 (N_2567,In_815,In_431);
xor U2568 (N_2568,In_807,In_1533);
or U2569 (N_2569,In_426,In_1320);
xor U2570 (N_2570,In_999,In_411);
or U2571 (N_2571,In_1953,In_1843);
xnor U2572 (N_2572,In_1767,In_858);
xnor U2573 (N_2573,In_1532,In_1533);
or U2574 (N_2574,In_672,In_1864);
or U2575 (N_2575,In_1879,In_57);
nand U2576 (N_2576,In_1861,In_570);
nand U2577 (N_2577,In_525,In_1543);
nand U2578 (N_2578,In_1879,In_853);
xnor U2579 (N_2579,In_438,In_1398);
nor U2580 (N_2580,In_1612,In_1133);
xor U2581 (N_2581,In_529,In_1031);
or U2582 (N_2582,In_858,In_570);
or U2583 (N_2583,In_1281,In_779);
nor U2584 (N_2584,In_1382,In_917);
xnor U2585 (N_2585,In_818,In_1334);
nand U2586 (N_2586,In_941,In_313);
and U2587 (N_2587,In_1038,In_53);
nand U2588 (N_2588,In_1290,In_1827);
nor U2589 (N_2589,In_1191,In_1865);
nor U2590 (N_2590,In_1254,In_1977);
or U2591 (N_2591,In_657,In_570);
xnor U2592 (N_2592,In_667,In_1054);
and U2593 (N_2593,In_241,In_445);
nor U2594 (N_2594,In_1441,In_456);
nor U2595 (N_2595,In_1253,In_717);
and U2596 (N_2596,In_1790,In_1364);
nor U2597 (N_2597,In_1520,In_1788);
xor U2598 (N_2598,In_1382,In_1844);
nor U2599 (N_2599,In_1604,In_737);
or U2600 (N_2600,In_1016,In_1815);
nand U2601 (N_2601,In_1909,In_1587);
nor U2602 (N_2602,In_183,In_1175);
nor U2603 (N_2603,In_1592,In_183);
and U2604 (N_2604,In_223,In_916);
nand U2605 (N_2605,In_495,In_1455);
or U2606 (N_2606,In_1135,In_1865);
nor U2607 (N_2607,In_367,In_257);
nand U2608 (N_2608,In_811,In_1073);
xnor U2609 (N_2609,In_345,In_1780);
nand U2610 (N_2610,In_494,In_700);
xnor U2611 (N_2611,In_786,In_415);
nand U2612 (N_2612,In_310,In_752);
xnor U2613 (N_2613,In_899,In_523);
nor U2614 (N_2614,In_163,In_1107);
and U2615 (N_2615,In_1632,In_26);
nand U2616 (N_2616,In_1662,In_352);
xnor U2617 (N_2617,In_1507,In_159);
xnor U2618 (N_2618,In_1678,In_1452);
nand U2619 (N_2619,In_873,In_1278);
or U2620 (N_2620,In_1478,In_728);
nand U2621 (N_2621,In_1955,In_788);
and U2622 (N_2622,In_1472,In_1411);
or U2623 (N_2623,In_941,In_817);
nor U2624 (N_2624,In_500,In_1581);
xnor U2625 (N_2625,In_210,In_477);
nand U2626 (N_2626,In_1654,In_1257);
xnor U2627 (N_2627,In_1069,In_1387);
nor U2628 (N_2628,In_620,In_609);
nand U2629 (N_2629,In_922,In_570);
and U2630 (N_2630,In_1679,In_374);
or U2631 (N_2631,In_1506,In_493);
and U2632 (N_2632,In_2,In_1208);
or U2633 (N_2633,In_948,In_612);
nand U2634 (N_2634,In_1992,In_6);
and U2635 (N_2635,In_1032,In_592);
and U2636 (N_2636,In_814,In_112);
xor U2637 (N_2637,In_1528,In_1340);
xor U2638 (N_2638,In_1796,In_523);
nor U2639 (N_2639,In_1387,In_77);
nor U2640 (N_2640,In_479,In_220);
or U2641 (N_2641,In_1596,In_33);
nand U2642 (N_2642,In_1999,In_458);
nand U2643 (N_2643,In_1757,In_803);
and U2644 (N_2644,In_1377,In_1989);
nor U2645 (N_2645,In_886,In_1442);
nor U2646 (N_2646,In_885,In_537);
and U2647 (N_2647,In_936,In_1522);
or U2648 (N_2648,In_52,In_606);
and U2649 (N_2649,In_1092,In_214);
nand U2650 (N_2650,In_1587,In_1820);
nor U2651 (N_2651,In_1508,In_1472);
nor U2652 (N_2652,In_934,In_1256);
xor U2653 (N_2653,In_950,In_1315);
and U2654 (N_2654,In_1395,In_1459);
nand U2655 (N_2655,In_1862,In_1077);
and U2656 (N_2656,In_1065,In_786);
nor U2657 (N_2657,In_126,In_923);
xor U2658 (N_2658,In_840,In_160);
or U2659 (N_2659,In_290,In_1780);
and U2660 (N_2660,In_1255,In_1582);
or U2661 (N_2661,In_1509,In_1981);
nor U2662 (N_2662,In_1435,In_513);
nor U2663 (N_2663,In_695,In_1002);
and U2664 (N_2664,In_1940,In_1636);
nor U2665 (N_2665,In_1984,In_1188);
or U2666 (N_2666,In_1659,In_753);
nand U2667 (N_2667,In_222,In_821);
xnor U2668 (N_2668,In_1061,In_1500);
and U2669 (N_2669,In_379,In_1560);
and U2670 (N_2670,In_175,In_1614);
xor U2671 (N_2671,In_548,In_643);
or U2672 (N_2672,In_454,In_1503);
nor U2673 (N_2673,In_1651,In_329);
nand U2674 (N_2674,In_733,In_1789);
nand U2675 (N_2675,In_1606,In_415);
xnor U2676 (N_2676,In_1427,In_1213);
nor U2677 (N_2677,In_82,In_1414);
xnor U2678 (N_2678,In_1024,In_1705);
and U2679 (N_2679,In_644,In_927);
and U2680 (N_2680,In_1934,In_911);
xnor U2681 (N_2681,In_701,In_1205);
xor U2682 (N_2682,In_543,In_296);
xor U2683 (N_2683,In_215,In_1779);
nand U2684 (N_2684,In_902,In_1257);
nand U2685 (N_2685,In_1160,In_1547);
or U2686 (N_2686,In_92,In_178);
and U2687 (N_2687,In_20,In_30);
or U2688 (N_2688,In_325,In_1944);
nand U2689 (N_2689,In_673,In_519);
and U2690 (N_2690,In_1591,In_392);
and U2691 (N_2691,In_435,In_1414);
or U2692 (N_2692,In_1790,In_498);
and U2693 (N_2693,In_1714,In_1309);
or U2694 (N_2694,In_99,In_1043);
xor U2695 (N_2695,In_1704,In_1460);
or U2696 (N_2696,In_1389,In_256);
nor U2697 (N_2697,In_1862,In_864);
xnor U2698 (N_2698,In_1033,In_535);
or U2699 (N_2699,In_1119,In_482);
or U2700 (N_2700,In_1316,In_288);
xnor U2701 (N_2701,In_1281,In_1391);
or U2702 (N_2702,In_1999,In_227);
xor U2703 (N_2703,In_1025,In_1239);
nand U2704 (N_2704,In_1754,In_1437);
xor U2705 (N_2705,In_1441,In_878);
and U2706 (N_2706,In_392,In_1200);
nor U2707 (N_2707,In_1654,In_51);
or U2708 (N_2708,In_1026,In_517);
or U2709 (N_2709,In_1177,In_1957);
xor U2710 (N_2710,In_1234,In_1619);
nor U2711 (N_2711,In_1438,In_1498);
and U2712 (N_2712,In_1295,In_81);
xor U2713 (N_2713,In_1853,In_1457);
or U2714 (N_2714,In_776,In_1819);
xnor U2715 (N_2715,In_842,In_283);
nor U2716 (N_2716,In_1814,In_1537);
or U2717 (N_2717,In_1268,In_871);
nand U2718 (N_2718,In_583,In_199);
or U2719 (N_2719,In_1729,In_1002);
and U2720 (N_2720,In_810,In_1792);
nand U2721 (N_2721,In_1946,In_1856);
nor U2722 (N_2722,In_1761,In_472);
and U2723 (N_2723,In_1919,In_1050);
xnor U2724 (N_2724,In_1942,In_1473);
and U2725 (N_2725,In_634,In_127);
xnor U2726 (N_2726,In_1858,In_1998);
nand U2727 (N_2727,In_14,In_391);
or U2728 (N_2728,In_162,In_427);
or U2729 (N_2729,In_1755,In_1036);
xor U2730 (N_2730,In_1865,In_568);
nor U2731 (N_2731,In_1339,In_1248);
xnor U2732 (N_2732,In_1152,In_768);
nor U2733 (N_2733,In_1148,In_982);
xnor U2734 (N_2734,In_1757,In_1384);
or U2735 (N_2735,In_174,In_1462);
nand U2736 (N_2736,In_1081,In_737);
nor U2737 (N_2737,In_1114,In_750);
nand U2738 (N_2738,In_188,In_402);
xnor U2739 (N_2739,In_481,In_276);
nand U2740 (N_2740,In_1280,In_732);
nor U2741 (N_2741,In_217,In_507);
nor U2742 (N_2742,In_1474,In_1885);
xor U2743 (N_2743,In_1507,In_1604);
and U2744 (N_2744,In_622,In_438);
and U2745 (N_2745,In_65,In_803);
or U2746 (N_2746,In_629,In_1404);
xnor U2747 (N_2747,In_1396,In_1569);
and U2748 (N_2748,In_199,In_1734);
and U2749 (N_2749,In_1402,In_795);
nor U2750 (N_2750,In_1208,In_1475);
xor U2751 (N_2751,In_1650,In_1324);
xnor U2752 (N_2752,In_1708,In_1743);
or U2753 (N_2753,In_268,In_1143);
and U2754 (N_2754,In_1389,In_1250);
xnor U2755 (N_2755,In_677,In_967);
nor U2756 (N_2756,In_800,In_491);
nand U2757 (N_2757,In_1774,In_1296);
and U2758 (N_2758,In_700,In_1958);
or U2759 (N_2759,In_292,In_1439);
xor U2760 (N_2760,In_1819,In_1939);
nand U2761 (N_2761,In_218,In_577);
xnor U2762 (N_2762,In_119,In_1089);
nor U2763 (N_2763,In_575,In_1405);
nand U2764 (N_2764,In_1590,In_911);
nand U2765 (N_2765,In_1334,In_240);
or U2766 (N_2766,In_1233,In_1618);
and U2767 (N_2767,In_11,In_707);
and U2768 (N_2768,In_125,In_697);
and U2769 (N_2769,In_177,In_955);
xnor U2770 (N_2770,In_309,In_1167);
nand U2771 (N_2771,In_1213,In_1974);
or U2772 (N_2772,In_144,In_878);
xor U2773 (N_2773,In_506,In_322);
nor U2774 (N_2774,In_1844,In_729);
xnor U2775 (N_2775,In_1167,In_438);
and U2776 (N_2776,In_542,In_163);
nand U2777 (N_2777,In_1650,In_1971);
xor U2778 (N_2778,In_1699,In_248);
or U2779 (N_2779,In_1562,In_668);
nand U2780 (N_2780,In_625,In_1157);
and U2781 (N_2781,In_650,In_1630);
xnor U2782 (N_2782,In_711,In_264);
or U2783 (N_2783,In_224,In_1298);
nor U2784 (N_2784,In_1303,In_669);
nor U2785 (N_2785,In_1629,In_1702);
or U2786 (N_2786,In_1187,In_583);
or U2787 (N_2787,In_1390,In_352);
xor U2788 (N_2788,In_818,In_1635);
nand U2789 (N_2789,In_1429,In_1954);
nand U2790 (N_2790,In_1480,In_785);
and U2791 (N_2791,In_894,In_1074);
and U2792 (N_2792,In_1692,In_703);
xnor U2793 (N_2793,In_1057,In_1423);
and U2794 (N_2794,In_1536,In_916);
and U2795 (N_2795,In_211,In_1848);
nand U2796 (N_2796,In_1051,In_992);
nor U2797 (N_2797,In_1622,In_1859);
and U2798 (N_2798,In_438,In_1385);
xor U2799 (N_2799,In_217,In_1443);
and U2800 (N_2800,In_1561,In_951);
and U2801 (N_2801,In_772,In_1683);
nand U2802 (N_2802,In_1418,In_1046);
and U2803 (N_2803,In_1,In_20);
or U2804 (N_2804,In_1331,In_1177);
or U2805 (N_2805,In_157,In_129);
and U2806 (N_2806,In_319,In_1417);
or U2807 (N_2807,In_1755,In_138);
nand U2808 (N_2808,In_1325,In_853);
or U2809 (N_2809,In_760,In_166);
nand U2810 (N_2810,In_1960,In_748);
and U2811 (N_2811,In_435,In_1796);
and U2812 (N_2812,In_1057,In_1137);
nand U2813 (N_2813,In_1339,In_1645);
nand U2814 (N_2814,In_1490,In_1189);
and U2815 (N_2815,In_78,In_623);
and U2816 (N_2816,In_1047,In_1);
xor U2817 (N_2817,In_134,In_1951);
nor U2818 (N_2818,In_1128,In_718);
nor U2819 (N_2819,In_1759,In_214);
xnor U2820 (N_2820,In_1038,In_1415);
nor U2821 (N_2821,In_1987,In_20);
nor U2822 (N_2822,In_515,In_1647);
or U2823 (N_2823,In_154,In_1757);
nor U2824 (N_2824,In_604,In_1476);
nand U2825 (N_2825,In_1693,In_182);
nor U2826 (N_2826,In_1136,In_139);
nand U2827 (N_2827,In_1433,In_65);
and U2828 (N_2828,In_1798,In_1987);
xor U2829 (N_2829,In_1040,In_1662);
nand U2830 (N_2830,In_475,In_1838);
nand U2831 (N_2831,In_31,In_488);
nand U2832 (N_2832,In_1901,In_286);
and U2833 (N_2833,In_1091,In_527);
xor U2834 (N_2834,In_125,In_216);
xor U2835 (N_2835,In_1849,In_1404);
or U2836 (N_2836,In_794,In_600);
nand U2837 (N_2837,In_1770,In_22);
nor U2838 (N_2838,In_901,In_1865);
and U2839 (N_2839,In_147,In_380);
and U2840 (N_2840,In_38,In_1391);
nand U2841 (N_2841,In_251,In_172);
nand U2842 (N_2842,In_1606,In_543);
nor U2843 (N_2843,In_70,In_1024);
or U2844 (N_2844,In_1217,In_297);
or U2845 (N_2845,In_1717,In_1163);
or U2846 (N_2846,In_1216,In_1863);
nor U2847 (N_2847,In_1274,In_473);
and U2848 (N_2848,In_1958,In_128);
or U2849 (N_2849,In_1562,In_1817);
nor U2850 (N_2850,In_1403,In_1320);
xnor U2851 (N_2851,In_1102,In_1720);
or U2852 (N_2852,In_176,In_155);
nand U2853 (N_2853,In_161,In_1024);
and U2854 (N_2854,In_1667,In_857);
xor U2855 (N_2855,In_182,In_479);
and U2856 (N_2856,In_1117,In_1371);
nand U2857 (N_2857,In_1574,In_925);
nand U2858 (N_2858,In_656,In_231);
and U2859 (N_2859,In_714,In_205);
and U2860 (N_2860,In_1181,In_574);
and U2861 (N_2861,In_1450,In_582);
nor U2862 (N_2862,In_826,In_284);
xnor U2863 (N_2863,In_1813,In_1710);
xor U2864 (N_2864,In_1613,In_1435);
nand U2865 (N_2865,In_523,In_1515);
xor U2866 (N_2866,In_885,In_241);
nor U2867 (N_2867,In_196,In_1748);
or U2868 (N_2868,In_1710,In_1353);
nor U2869 (N_2869,In_1748,In_1012);
xor U2870 (N_2870,In_1258,In_120);
nand U2871 (N_2871,In_44,In_168);
or U2872 (N_2872,In_950,In_1288);
nand U2873 (N_2873,In_33,In_1182);
xor U2874 (N_2874,In_289,In_1209);
nor U2875 (N_2875,In_794,In_1833);
nand U2876 (N_2876,In_877,In_683);
and U2877 (N_2877,In_255,In_1092);
or U2878 (N_2878,In_1864,In_1678);
xnor U2879 (N_2879,In_1548,In_1158);
nor U2880 (N_2880,In_316,In_1441);
and U2881 (N_2881,In_1897,In_886);
and U2882 (N_2882,In_1433,In_1478);
or U2883 (N_2883,In_1056,In_803);
or U2884 (N_2884,In_1989,In_1532);
nand U2885 (N_2885,In_1898,In_1287);
and U2886 (N_2886,In_568,In_1591);
nor U2887 (N_2887,In_1198,In_1388);
nor U2888 (N_2888,In_179,In_1495);
nor U2889 (N_2889,In_1418,In_478);
xor U2890 (N_2890,In_1070,In_1590);
xnor U2891 (N_2891,In_676,In_1273);
nor U2892 (N_2892,In_41,In_1729);
and U2893 (N_2893,In_40,In_598);
nand U2894 (N_2894,In_839,In_831);
or U2895 (N_2895,In_371,In_1669);
and U2896 (N_2896,In_1781,In_635);
nand U2897 (N_2897,In_1194,In_1080);
or U2898 (N_2898,In_508,In_1462);
xor U2899 (N_2899,In_749,In_370);
and U2900 (N_2900,In_837,In_1740);
nand U2901 (N_2901,In_1908,In_1398);
nand U2902 (N_2902,In_1523,In_89);
or U2903 (N_2903,In_1935,In_1712);
xor U2904 (N_2904,In_251,In_354);
or U2905 (N_2905,In_1963,In_652);
nand U2906 (N_2906,In_412,In_1674);
and U2907 (N_2907,In_145,In_1104);
or U2908 (N_2908,In_1681,In_1255);
nand U2909 (N_2909,In_1505,In_1678);
and U2910 (N_2910,In_41,In_1504);
and U2911 (N_2911,In_1310,In_579);
and U2912 (N_2912,In_251,In_1590);
nand U2913 (N_2913,In_285,In_1536);
xnor U2914 (N_2914,In_1921,In_1949);
and U2915 (N_2915,In_1344,In_1768);
nand U2916 (N_2916,In_612,In_443);
and U2917 (N_2917,In_958,In_940);
or U2918 (N_2918,In_958,In_714);
nand U2919 (N_2919,In_1651,In_822);
nand U2920 (N_2920,In_939,In_1408);
and U2921 (N_2921,In_957,In_1380);
nor U2922 (N_2922,In_1305,In_171);
nand U2923 (N_2923,In_1909,In_1681);
nand U2924 (N_2924,In_1688,In_1538);
nor U2925 (N_2925,In_1952,In_591);
nor U2926 (N_2926,In_1133,In_760);
and U2927 (N_2927,In_1871,In_171);
and U2928 (N_2928,In_540,In_494);
or U2929 (N_2929,In_198,In_904);
and U2930 (N_2930,In_881,In_1291);
nand U2931 (N_2931,In_1178,In_574);
xnor U2932 (N_2932,In_467,In_187);
nand U2933 (N_2933,In_281,In_1776);
or U2934 (N_2934,In_1899,In_1934);
or U2935 (N_2935,In_589,In_197);
nand U2936 (N_2936,In_1621,In_1074);
xor U2937 (N_2937,In_1271,In_527);
and U2938 (N_2938,In_245,In_231);
or U2939 (N_2939,In_83,In_1174);
and U2940 (N_2940,In_1294,In_0);
or U2941 (N_2941,In_574,In_628);
and U2942 (N_2942,In_623,In_1363);
xor U2943 (N_2943,In_539,In_1580);
xnor U2944 (N_2944,In_23,In_1886);
xor U2945 (N_2945,In_269,In_634);
nand U2946 (N_2946,In_1359,In_138);
or U2947 (N_2947,In_1782,In_1159);
and U2948 (N_2948,In_664,In_1489);
nand U2949 (N_2949,In_1037,In_1650);
xor U2950 (N_2950,In_286,In_218);
nand U2951 (N_2951,In_1754,In_10);
xnor U2952 (N_2952,In_1958,In_329);
xor U2953 (N_2953,In_893,In_1780);
xor U2954 (N_2954,In_220,In_1661);
xnor U2955 (N_2955,In_1235,In_570);
or U2956 (N_2956,In_87,In_222);
nor U2957 (N_2957,In_310,In_1265);
and U2958 (N_2958,In_1932,In_1255);
or U2959 (N_2959,In_1284,In_964);
and U2960 (N_2960,In_1713,In_441);
or U2961 (N_2961,In_1234,In_1597);
nand U2962 (N_2962,In_642,In_881);
and U2963 (N_2963,In_978,In_444);
xnor U2964 (N_2964,In_1746,In_1855);
or U2965 (N_2965,In_1807,In_1509);
xnor U2966 (N_2966,In_460,In_757);
xnor U2967 (N_2967,In_132,In_852);
nand U2968 (N_2968,In_1118,In_1097);
nand U2969 (N_2969,In_1774,In_1005);
xor U2970 (N_2970,In_1395,In_1114);
nand U2971 (N_2971,In_680,In_454);
xor U2972 (N_2972,In_1198,In_100);
or U2973 (N_2973,In_51,In_766);
nand U2974 (N_2974,In_1466,In_540);
or U2975 (N_2975,In_199,In_1990);
nor U2976 (N_2976,In_1956,In_87);
or U2977 (N_2977,In_851,In_1813);
xor U2978 (N_2978,In_145,In_1701);
nand U2979 (N_2979,In_1707,In_610);
xor U2980 (N_2980,In_658,In_682);
xor U2981 (N_2981,In_727,In_1407);
nand U2982 (N_2982,In_762,In_220);
or U2983 (N_2983,In_1139,In_291);
and U2984 (N_2984,In_1625,In_947);
or U2985 (N_2985,In_1818,In_5);
xnor U2986 (N_2986,In_181,In_317);
nor U2987 (N_2987,In_988,In_1577);
nand U2988 (N_2988,In_1979,In_655);
or U2989 (N_2989,In_1122,In_644);
xor U2990 (N_2990,In_1486,In_976);
or U2991 (N_2991,In_755,In_1541);
or U2992 (N_2992,In_1553,In_1715);
nor U2993 (N_2993,In_468,In_1877);
nor U2994 (N_2994,In_1137,In_1823);
nand U2995 (N_2995,In_1218,In_1401);
or U2996 (N_2996,In_884,In_1294);
and U2997 (N_2997,In_1310,In_1143);
nand U2998 (N_2998,In_1208,In_1077);
nand U2999 (N_2999,In_618,In_790);
or U3000 (N_3000,In_836,In_1807);
and U3001 (N_3001,In_1840,In_836);
or U3002 (N_3002,In_103,In_1620);
nand U3003 (N_3003,In_974,In_964);
nor U3004 (N_3004,In_1341,In_1317);
xnor U3005 (N_3005,In_1530,In_1873);
nand U3006 (N_3006,In_1287,In_1475);
nor U3007 (N_3007,In_1720,In_772);
and U3008 (N_3008,In_1409,In_691);
and U3009 (N_3009,In_346,In_1360);
and U3010 (N_3010,In_1564,In_109);
or U3011 (N_3011,In_924,In_1884);
xor U3012 (N_3012,In_559,In_237);
nor U3013 (N_3013,In_201,In_1903);
xor U3014 (N_3014,In_140,In_552);
and U3015 (N_3015,In_1831,In_1737);
and U3016 (N_3016,In_385,In_701);
or U3017 (N_3017,In_1672,In_1392);
nor U3018 (N_3018,In_1501,In_1062);
nand U3019 (N_3019,In_1665,In_666);
xor U3020 (N_3020,In_942,In_373);
nor U3021 (N_3021,In_1591,In_1377);
and U3022 (N_3022,In_1794,In_456);
nand U3023 (N_3023,In_1951,In_755);
nand U3024 (N_3024,In_95,In_1339);
nand U3025 (N_3025,In_1328,In_295);
or U3026 (N_3026,In_822,In_1020);
nor U3027 (N_3027,In_1632,In_496);
nand U3028 (N_3028,In_735,In_840);
nand U3029 (N_3029,In_1969,In_359);
and U3030 (N_3030,In_1073,In_1134);
nor U3031 (N_3031,In_111,In_1563);
or U3032 (N_3032,In_69,In_1857);
xor U3033 (N_3033,In_494,In_1920);
or U3034 (N_3034,In_573,In_1728);
and U3035 (N_3035,In_532,In_383);
nand U3036 (N_3036,In_1917,In_1444);
or U3037 (N_3037,In_79,In_1362);
nand U3038 (N_3038,In_1591,In_1755);
nor U3039 (N_3039,In_1800,In_418);
or U3040 (N_3040,In_425,In_39);
nand U3041 (N_3041,In_1472,In_125);
or U3042 (N_3042,In_1426,In_843);
and U3043 (N_3043,In_1788,In_1096);
and U3044 (N_3044,In_1356,In_779);
xor U3045 (N_3045,In_1540,In_917);
and U3046 (N_3046,In_171,In_1598);
or U3047 (N_3047,In_1275,In_476);
nand U3048 (N_3048,In_429,In_1496);
nor U3049 (N_3049,In_1394,In_1672);
xor U3050 (N_3050,In_307,In_147);
or U3051 (N_3051,In_23,In_1632);
and U3052 (N_3052,In_791,In_180);
nor U3053 (N_3053,In_1013,In_1086);
nor U3054 (N_3054,In_1023,In_67);
and U3055 (N_3055,In_1258,In_1172);
xnor U3056 (N_3056,In_740,In_483);
xor U3057 (N_3057,In_1191,In_1336);
nand U3058 (N_3058,In_1792,In_1210);
or U3059 (N_3059,In_1283,In_137);
xor U3060 (N_3060,In_11,In_1780);
xor U3061 (N_3061,In_1087,In_174);
nor U3062 (N_3062,In_1962,In_990);
and U3063 (N_3063,In_1957,In_145);
nand U3064 (N_3064,In_1811,In_1225);
or U3065 (N_3065,In_462,In_753);
nand U3066 (N_3066,In_220,In_72);
nand U3067 (N_3067,In_1408,In_450);
nand U3068 (N_3068,In_308,In_896);
and U3069 (N_3069,In_1300,In_1163);
nor U3070 (N_3070,In_1842,In_1767);
nand U3071 (N_3071,In_1852,In_669);
and U3072 (N_3072,In_392,In_1725);
xor U3073 (N_3073,In_1932,In_107);
xnor U3074 (N_3074,In_260,In_450);
nand U3075 (N_3075,In_132,In_1258);
nand U3076 (N_3076,In_913,In_1716);
xnor U3077 (N_3077,In_1053,In_1442);
nor U3078 (N_3078,In_1930,In_1392);
nand U3079 (N_3079,In_1417,In_1528);
nand U3080 (N_3080,In_850,In_1441);
or U3081 (N_3081,In_1135,In_780);
nor U3082 (N_3082,In_1079,In_614);
or U3083 (N_3083,In_487,In_1521);
nand U3084 (N_3084,In_163,In_1449);
nand U3085 (N_3085,In_1830,In_449);
xor U3086 (N_3086,In_698,In_538);
nand U3087 (N_3087,In_858,In_1386);
or U3088 (N_3088,In_1144,In_1580);
nor U3089 (N_3089,In_10,In_1784);
xor U3090 (N_3090,In_1726,In_1743);
nor U3091 (N_3091,In_803,In_465);
nand U3092 (N_3092,In_206,In_228);
xnor U3093 (N_3093,In_1714,In_264);
or U3094 (N_3094,In_138,In_756);
and U3095 (N_3095,In_136,In_300);
or U3096 (N_3096,In_1380,In_1831);
xnor U3097 (N_3097,In_1754,In_1782);
nor U3098 (N_3098,In_153,In_1646);
xor U3099 (N_3099,In_583,In_1961);
nand U3100 (N_3100,In_543,In_1663);
nor U3101 (N_3101,In_975,In_1028);
nor U3102 (N_3102,In_1643,In_1519);
and U3103 (N_3103,In_203,In_814);
nor U3104 (N_3104,In_741,In_140);
nor U3105 (N_3105,In_961,In_204);
xor U3106 (N_3106,In_1905,In_1260);
nand U3107 (N_3107,In_118,In_1495);
or U3108 (N_3108,In_1332,In_1102);
nor U3109 (N_3109,In_1505,In_1869);
and U3110 (N_3110,In_390,In_1130);
nor U3111 (N_3111,In_880,In_691);
or U3112 (N_3112,In_1816,In_992);
nor U3113 (N_3113,In_1114,In_1625);
or U3114 (N_3114,In_846,In_726);
or U3115 (N_3115,In_1099,In_1460);
xnor U3116 (N_3116,In_1716,In_925);
nand U3117 (N_3117,In_1890,In_1358);
and U3118 (N_3118,In_1790,In_1796);
and U3119 (N_3119,In_1749,In_1877);
xnor U3120 (N_3120,In_33,In_661);
or U3121 (N_3121,In_1395,In_1051);
or U3122 (N_3122,In_274,In_743);
or U3123 (N_3123,In_1341,In_496);
or U3124 (N_3124,In_1335,In_800);
nand U3125 (N_3125,In_1730,In_1159);
nor U3126 (N_3126,In_581,In_1384);
and U3127 (N_3127,In_1763,In_860);
or U3128 (N_3128,In_1474,In_168);
nor U3129 (N_3129,In_776,In_227);
xor U3130 (N_3130,In_1170,In_1772);
nor U3131 (N_3131,In_696,In_33);
and U3132 (N_3132,In_1232,In_1547);
and U3133 (N_3133,In_1530,In_1624);
or U3134 (N_3134,In_1187,In_1392);
nor U3135 (N_3135,In_586,In_1268);
nor U3136 (N_3136,In_1648,In_802);
and U3137 (N_3137,In_812,In_1034);
nor U3138 (N_3138,In_973,In_588);
and U3139 (N_3139,In_1540,In_79);
nor U3140 (N_3140,In_453,In_1317);
and U3141 (N_3141,In_1317,In_1667);
and U3142 (N_3142,In_599,In_717);
or U3143 (N_3143,In_1973,In_849);
or U3144 (N_3144,In_96,In_326);
nor U3145 (N_3145,In_1588,In_1314);
nor U3146 (N_3146,In_1047,In_1011);
or U3147 (N_3147,In_164,In_1090);
xnor U3148 (N_3148,In_531,In_308);
or U3149 (N_3149,In_1866,In_254);
nor U3150 (N_3150,In_63,In_708);
nor U3151 (N_3151,In_1366,In_501);
or U3152 (N_3152,In_1948,In_51);
xor U3153 (N_3153,In_1106,In_1812);
and U3154 (N_3154,In_1631,In_1136);
xor U3155 (N_3155,In_891,In_1557);
xor U3156 (N_3156,In_1190,In_1276);
xnor U3157 (N_3157,In_1171,In_1146);
or U3158 (N_3158,In_390,In_13);
nand U3159 (N_3159,In_462,In_1494);
or U3160 (N_3160,In_1617,In_54);
nor U3161 (N_3161,In_1954,In_429);
nand U3162 (N_3162,In_1370,In_665);
nor U3163 (N_3163,In_1663,In_1407);
nor U3164 (N_3164,In_369,In_1217);
and U3165 (N_3165,In_726,In_1950);
or U3166 (N_3166,In_1585,In_776);
nor U3167 (N_3167,In_5,In_1992);
and U3168 (N_3168,In_1177,In_1910);
nand U3169 (N_3169,In_1452,In_115);
or U3170 (N_3170,In_994,In_1031);
nand U3171 (N_3171,In_366,In_1599);
or U3172 (N_3172,In_210,In_1245);
or U3173 (N_3173,In_1930,In_31);
or U3174 (N_3174,In_193,In_1308);
and U3175 (N_3175,In_1851,In_538);
nand U3176 (N_3176,In_674,In_648);
nor U3177 (N_3177,In_221,In_25);
xor U3178 (N_3178,In_755,In_386);
nand U3179 (N_3179,In_1978,In_1867);
and U3180 (N_3180,In_1048,In_626);
xor U3181 (N_3181,In_964,In_202);
nor U3182 (N_3182,In_493,In_51);
and U3183 (N_3183,In_163,In_55);
or U3184 (N_3184,In_1073,In_399);
nor U3185 (N_3185,In_1799,In_481);
or U3186 (N_3186,In_1066,In_1244);
or U3187 (N_3187,In_1726,In_159);
nand U3188 (N_3188,In_774,In_757);
nor U3189 (N_3189,In_1281,In_310);
or U3190 (N_3190,In_1503,In_129);
and U3191 (N_3191,In_1442,In_1592);
or U3192 (N_3192,In_1237,In_583);
nand U3193 (N_3193,In_1036,In_938);
and U3194 (N_3194,In_1271,In_329);
xor U3195 (N_3195,In_1991,In_1524);
or U3196 (N_3196,In_1764,In_946);
and U3197 (N_3197,In_353,In_1249);
nor U3198 (N_3198,In_1577,In_964);
nor U3199 (N_3199,In_70,In_629);
xor U3200 (N_3200,In_771,In_559);
nand U3201 (N_3201,In_510,In_1741);
or U3202 (N_3202,In_1324,In_1365);
nor U3203 (N_3203,In_916,In_1306);
xnor U3204 (N_3204,In_1199,In_189);
nor U3205 (N_3205,In_1987,In_892);
and U3206 (N_3206,In_1252,In_87);
or U3207 (N_3207,In_1398,In_1572);
nand U3208 (N_3208,In_1545,In_71);
nand U3209 (N_3209,In_1508,In_255);
xor U3210 (N_3210,In_1914,In_1857);
xnor U3211 (N_3211,In_554,In_695);
and U3212 (N_3212,In_403,In_932);
or U3213 (N_3213,In_681,In_1649);
xor U3214 (N_3214,In_1813,In_1299);
and U3215 (N_3215,In_698,In_1859);
or U3216 (N_3216,In_1266,In_1648);
xor U3217 (N_3217,In_28,In_370);
and U3218 (N_3218,In_1711,In_1570);
xnor U3219 (N_3219,In_1468,In_1344);
xnor U3220 (N_3220,In_1893,In_90);
xor U3221 (N_3221,In_1371,In_1276);
nor U3222 (N_3222,In_164,In_1980);
nor U3223 (N_3223,In_99,In_1621);
or U3224 (N_3224,In_320,In_192);
nor U3225 (N_3225,In_264,In_547);
nor U3226 (N_3226,In_1585,In_487);
nand U3227 (N_3227,In_1561,In_530);
nand U3228 (N_3228,In_55,In_1635);
nor U3229 (N_3229,In_1616,In_1060);
xor U3230 (N_3230,In_1580,In_1115);
and U3231 (N_3231,In_720,In_1660);
or U3232 (N_3232,In_1999,In_855);
nand U3233 (N_3233,In_477,In_721);
and U3234 (N_3234,In_888,In_330);
and U3235 (N_3235,In_736,In_1392);
and U3236 (N_3236,In_1539,In_1707);
or U3237 (N_3237,In_1343,In_255);
xor U3238 (N_3238,In_216,In_141);
xnor U3239 (N_3239,In_1627,In_1982);
nor U3240 (N_3240,In_1430,In_1011);
nand U3241 (N_3241,In_1969,In_1553);
and U3242 (N_3242,In_382,In_587);
or U3243 (N_3243,In_1978,In_1716);
nor U3244 (N_3244,In_1541,In_1515);
nor U3245 (N_3245,In_149,In_897);
and U3246 (N_3246,In_118,In_1903);
nor U3247 (N_3247,In_1852,In_1724);
nor U3248 (N_3248,In_174,In_734);
or U3249 (N_3249,In_67,In_1624);
or U3250 (N_3250,In_1657,In_1982);
xnor U3251 (N_3251,In_559,In_614);
and U3252 (N_3252,In_1096,In_1468);
xor U3253 (N_3253,In_1795,In_625);
nor U3254 (N_3254,In_894,In_463);
nor U3255 (N_3255,In_910,In_87);
or U3256 (N_3256,In_880,In_1889);
nor U3257 (N_3257,In_1540,In_1475);
nor U3258 (N_3258,In_438,In_1777);
nand U3259 (N_3259,In_1588,In_1030);
and U3260 (N_3260,In_984,In_134);
or U3261 (N_3261,In_1852,In_623);
nor U3262 (N_3262,In_1263,In_1640);
nor U3263 (N_3263,In_1328,In_1189);
or U3264 (N_3264,In_511,In_1240);
or U3265 (N_3265,In_1121,In_1819);
and U3266 (N_3266,In_1378,In_1538);
xor U3267 (N_3267,In_1117,In_93);
and U3268 (N_3268,In_1433,In_128);
xnor U3269 (N_3269,In_279,In_1950);
nor U3270 (N_3270,In_543,In_1566);
or U3271 (N_3271,In_962,In_1359);
and U3272 (N_3272,In_801,In_383);
xnor U3273 (N_3273,In_497,In_1298);
nand U3274 (N_3274,In_730,In_201);
xor U3275 (N_3275,In_1931,In_1136);
xnor U3276 (N_3276,In_879,In_1236);
xor U3277 (N_3277,In_1733,In_1310);
xor U3278 (N_3278,In_1745,In_958);
and U3279 (N_3279,In_1932,In_570);
nor U3280 (N_3280,In_1976,In_1126);
nand U3281 (N_3281,In_909,In_670);
xnor U3282 (N_3282,In_745,In_1141);
xnor U3283 (N_3283,In_821,In_903);
and U3284 (N_3284,In_96,In_1781);
nor U3285 (N_3285,In_640,In_366);
xor U3286 (N_3286,In_1196,In_444);
or U3287 (N_3287,In_1511,In_249);
nor U3288 (N_3288,In_1534,In_1617);
xor U3289 (N_3289,In_1442,In_956);
xor U3290 (N_3290,In_614,In_1856);
or U3291 (N_3291,In_988,In_1031);
nand U3292 (N_3292,In_1351,In_772);
and U3293 (N_3293,In_1136,In_1756);
and U3294 (N_3294,In_634,In_1799);
nor U3295 (N_3295,In_42,In_1388);
and U3296 (N_3296,In_1050,In_1425);
or U3297 (N_3297,In_1580,In_17);
nor U3298 (N_3298,In_1716,In_1120);
nor U3299 (N_3299,In_1661,In_1864);
nor U3300 (N_3300,In_1634,In_1727);
or U3301 (N_3301,In_1550,In_1630);
and U3302 (N_3302,In_690,In_1274);
nor U3303 (N_3303,In_97,In_1548);
and U3304 (N_3304,In_174,In_878);
nand U3305 (N_3305,In_746,In_88);
or U3306 (N_3306,In_423,In_1688);
or U3307 (N_3307,In_317,In_610);
or U3308 (N_3308,In_160,In_1545);
xor U3309 (N_3309,In_381,In_1898);
and U3310 (N_3310,In_1374,In_1906);
and U3311 (N_3311,In_669,In_968);
nor U3312 (N_3312,In_421,In_1083);
or U3313 (N_3313,In_1937,In_1748);
and U3314 (N_3314,In_1826,In_665);
nand U3315 (N_3315,In_1333,In_436);
or U3316 (N_3316,In_192,In_1317);
xor U3317 (N_3317,In_1439,In_406);
nand U3318 (N_3318,In_482,In_1613);
nor U3319 (N_3319,In_511,In_678);
or U3320 (N_3320,In_1367,In_524);
nor U3321 (N_3321,In_1299,In_152);
nand U3322 (N_3322,In_122,In_1244);
xor U3323 (N_3323,In_1996,In_892);
and U3324 (N_3324,In_1708,In_977);
and U3325 (N_3325,In_1906,In_1647);
nand U3326 (N_3326,In_608,In_1615);
and U3327 (N_3327,In_1773,In_317);
or U3328 (N_3328,In_1808,In_885);
nand U3329 (N_3329,In_559,In_1670);
nand U3330 (N_3330,In_923,In_1077);
nor U3331 (N_3331,In_1024,In_31);
nor U3332 (N_3332,In_87,In_240);
nand U3333 (N_3333,In_491,In_1617);
xor U3334 (N_3334,In_1042,In_1808);
and U3335 (N_3335,In_46,In_1983);
nand U3336 (N_3336,In_913,In_1665);
xnor U3337 (N_3337,In_1351,In_1498);
xor U3338 (N_3338,In_1520,In_1038);
and U3339 (N_3339,In_1725,In_1559);
nand U3340 (N_3340,In_625,In_1949);
nand U3341 (N_3341,In_458,In_699);
nand U3342 (N_3342,In_770,In_1381);
and U3343 (N_3343,In_1032,In_521);
nand U3344 (N_3344,In_1095,In_1405);
nand U3345 (N_3345,In_1027,In_437);
and U3346 (N_3346,In_1957,In_1631);
nor U3347 (N_3347,In_293,In_1001);
or U3348 (N_3348,In_746,In_1574);
xnor U3349 (N_3349,In_12,In_1893);
nor U3350 (N_3350,In_691,In_557);
or U3351 (N_3351,In_661,In_1064);
nor U3352 (N_3352,In_1027,In_1404);
nor U3353 (N_3353,In_1202,In_166);
and U3354 (N_3354,In_290,In_1700);
nor U3355 (N_3355,In_1440,In_1252);
nand U3356 (N_3356,In_408,In_56);
xnor U3357 (N_3357,In_1973,In_917);
nor U3358 (N_3358,In_509,In_1957);
or U3359 (N_3359,In_865,In_616);
xnor U3360 (N_3360,In_570,In_593);
and U3361 (N_3361,In_1361,In_917);
or U3362 (N_3362,In_705,In_1747);
xnor U3363 (N_3363,In_1917,In_1136);
nand U3364 (N_3364,In_1810,In_212);
nor U3365 (N_3365,In_1093,In_1424);
nor U3366 (N_3366,In_961,In_726);
nand U3367 (N_3367,In_496,In_32);
and U3368 (N_3368,In_1003,In_1989);
nand U3369 (N_3369,In_552,In_1895);
nand U3370 (N_3370,In_113,In_1604);
nor U3371 (N_3371,In_337,In_664);
or U3372 (N_3372,In_783,In_697);
and U3373 (N_3373,In_1599,In_1207);
nand U3374 (N_3374,In_869,In_1987);
or U3375 (N_3375,In_424,In_1794);
and U3376 (N_3376,In_910,In_834);
nand U3377 (N_3377,In_1406,In_1620);
and U3378 (N_3378,In_245,In_969);
nand U3379 (N_3379,In_466,In_474);
nand U3380 (N_3380,In_5,In_1003);
nand U3381 (N_3381,In_377,In_593);
or U3382 (N_3382,In_623,In_1492);
and U3383 (N_3383,In_1570,In_624);
xnor U3384 (N_3384,In_152,In_233);
nand U3385 (N_3385,In_1812,In_1699);
or U3386 (N_3386,In_661,In_821);
xnor U3387 (N_3387,In_686,In_726);
or U3388 (N_3388,In_827,In_1025);
and U3389 (N_3389,In_170,In_381);
xor U3390 (N_3390,In_1496,In_1575);
or U3391 (N_3391,In_591,In_397);
or U3392 (N_3392,In_1154,In_1939);
and U3393 (N_3393,In_375,In_1460);
and U3394 (N_3394,In_1179,In_612);
xnor U3395 (N_3395,In_488,In_1070);
nor U3396 (N_3396,In_976,In_764);
nand U3397 (N_3397,In_1106,In_1014);
nor U3398 (N_3398,In_1252,In_1210);
nor U3399 (N_3399,In_1156,In_432);
nor U3400 (N_3400,In_991,In_1998);
xnor U3401 (N_3401,In_1412,In_541);
nand U3402 (N_3402,In_1332,In_148);
or U3403 (N_3403,In_1134,In_1854);
and U3404 (N_3404,In_261,In_631);
xor U3405 (N_3405,In_1971,In_91);
nand U3406 (N_3406,In_150,In_1182);
or U3407 (N_3407,In_1721,In_1001);
or U3408 (N_3408,In_155,In_355);
nand U3409 (N_3409,In_93,In_1410);
xnor U3410 (N_3410,In_33,In_452);
xnor U3411 (N_3411,In_949,In_369);
and U3412 (N_3412,In_357,In_229);
nor U3413 (N_3413,In_342,In_1059);
or U3414 (N_3414,In_536,In_1155);
nor U3415 (N_3415,In_1784,In_1375);
xor U3416 (N_3416,In_1757,In_1037);
nand U3417 (N_3417,In_1200,In_542);
nand U3418 (N_3418,In_1933,In_68);
nor U3419 (N_3419,In_756,In_974);
nand U3420 (N_3420,In_1641,In_679);
xnor U3421 (N_3421,In_1909,In_1442);
xor U3422 (N_3422,In_601,In_908);
nand U3423 (N_3423,In_25,In_1266);
nor U3424 (N_3424,In_401,In_282);
or U3425 (N_3425,In_1312,In_479);
and U3426 (N_3426,In_1473,In_680);
xnor U3427 (N_3427,In_1113,In_331);
nor U3428 (N_3428,In_1303,In_1167);
and U3429 (N_3429,In_1587,In_1768);
nand U3430 (N_3430,In_143,In_126);
or U3431 (N_3431,In_1007,In_829);
or U3432 (N_3432,In_597,In_624);
or U3433 (N_3433,In_1610,In_964);
xnor U3434 (N_3434,In_1725,In_1951);
or U3435 (N_3435,In_1566,In_1015);
and U3436 (N_3436,In_128,In_1055);
nor U3437 (N_3437,In_280,In_488);
nand U3438 (N_3438,In_478,In_1153);
or U3439 (N_3439,In_747,In_1408);
and U3440 (N_3440,In_410,In_519);
or U3441 (N_3441,In_1694,In_201);
nor U3442 (N_3442,In_754,In_1771);
xor U3443 (N_3443,In_857,In_1117);
and U3444 (N_3444,In_1008,In_1407);
or U3445 (N_3445,In_184,In_781);
nor U3446 (N_3446,In_1926,In_584);
nand U3447 (N_3447,In_424,In_1359);
or U3448 (N_3448,In_1474,In_397);
and U3449 (N_3449,In_325,In_323);
nor U3450 (N_3450,In_1307,In_1908);
and U3451 (N_3451,In_9,In_569);
nand U3452 (N_3452,In_35,In_1074);
nor U3453 (N_3453,In_38,In_59);
nand U3454 (N_3454,In_1293,In_1287);
and U3455 (N_3455,In_69,In_1189);
nor U3456 (N_3456,In_508,In_46);
or U3457 (N_3457,In_836,In_283);
or U3458 (N_3458,In_334,In_1373);
and U3459 (N_3459,In_277,In_1026);
nor U3460 (N_3460,In_154,In_295);
nor U3461 (N_3461,In_1244,In_13);
and U3462 (N_3462,In_1997,In_1241);
nand U3463 (N_3463,In_684,In_777);
and U3464 (N_3464,In_226,In_678);
nor U3465 (N_3465,In_1641,In_1220);
nor U3466 (N_3466,In_1455,In_737);
or U3467 (N_3467,In_1330,In_1772);
nor U3468 (N_3468,In_344,In_912);
and U3469 (N_3469,In_1569,In_1593);
or U3470 (N_3470,In_617,In_142);
nor U3471 (N_3471,In_479,In_860);
and U3472 (N_3472,In_386,In_964);
xnor U3473 (N_3473,In_612,In_1434);
xnor U3474 (N_3474,In_1181,In_1701);
nand U3475 (N_3475,In_804,In_1724);
and U3476 (N_3476,In_68,In_1805);
and U3477 (N_3477,In_143,In_547);
xnor U3478 (N_3478,In_1968,In_352);
or U3479 (N_3479,In_1792,In_245);
or U3480 (N_3480,In_77,In_1907);
nand U3481 (N_3481,In_1820,In_941);
nand U3482 (N_3482,In_1548,In_773);
or U3483 (N_3483,In_1508,In_1462);
nand U3484 (N_3484,In_166,In_941);
nor U3485 (N_3485,In_1520,In_1565);
xor U3486 (N_3486,In_169,In_1128);
nor U3487 (N_3487,In_1737,In_1765);
or U3488 (N_3488,In_114,In_964);
xnor U3489 (N_3489,In_490,In_269);
nand U3490 (N_3490,In_1644,In_914);
and U3491 (N_3491,In_269,In_805);
and U3492 (N_3492,In_609,In_290);
nand U3493 (N_3493,In_1052,In_982);
nand U3494 (N_3494,In_391,In_1499);
or U3495 (N_3495,In_1821,In_967);
or U3496 (N_3496,In_1672,In_110);
and U3497 (N_3497,In_578,In_97);
nor U3498 (N_3498,In_465,In_1434);
and U3499 (N_3499,In_1409,In_196);
and U3500 (N_3500,In_1702,In_1675);
xnor U3501 (N_3501,In_1851,In_205);
and U3502 (N_3502,In_119,In_1733);
or U3503 (N_3503,In_948,In_1315);
nand U3504 (N_3504,In_1060,In_915);
and U3505 (N_3505,In_942,In_1843);
and U3506 (N_3506,In_604,In_1305);
nand U3507 (N_3507,In_1988,In_65);
or U3508 (N_3508,In_783,In_972);
or U3509 (N_3509,In_1864,In_407);
nand U3510 (N_3510,In_35,In_812);
nand U3511 (N_3511,In_504,In_931);
and U3512 (N_3512,In_1196,In_1991);
and U3513 (N_3513,In_1034,In_724);
nor U3514 (N_3514,In_910,In_1307);
or U3515 (N_3515,In_1285,In_1143);
xnor U3516 (N_3516,In_181,In_1286);
or U3517 (N_3517,In_180,In_1377);
and U3518 (N_3518,In_1714,In_1397);
nand U3519 (N_3519,In_329,In_1116);
xor U3520 (N_3520,In_208,In_528);
nand U3521 (N_3521,In_1843,In_798);
nand U3522 (N_3522,In_1508,In_1570);
nand U3523 (N_3523,In_699,In_1801);
or U3524 (N_3524,In_1683,In_1747);
nor U3525 (N_3525,In_1416,In_645);
nor U3526 (N_3526,In_1111,In_1996);
nor U3527 (N_3527,In_1500,In_1021);
or U3528 (N_3528,In_965,In_195);
or U3529 (N_3529,In_609,In_986);
xnor U3530 (N_3530,In_1984,In_1190);
and U3531 (N_3531,In_1734,In_244);
and U3532 (N_3532,In_122,In_1464);
nand U3533 (N_3533,In_751,In_1247);
xnor U3534 (N_3534,In_1319,In_342);
nand U3535 (N_3535,In_519,In_1708);
nand U3536 (N_3536,In_1889,In_827);
or U3537 (N_3537,In_637,In_916);
xnor U3538 (N_3538,In_1097,In_447);
xor U3539 (N_3539,In_185,In_178);
xnor U3540 (N_3540,In_1476,In_1881);
or U3541 (N_3541,In_1816,In_538);
and U3542 (N_3542,In_1745,In_642);
nor U3543 (N_3543,In_1222,In_873);
and U3544 (N_3544,In_1923,In_477);
and U3545 (N_3545,In_1286,In_555);
nand U3546 (N_3546,In_1990,In_117);
nor U3547 (N_3547,In_1417,In_219);
nand U3548 (N_3548,In_767,In_1205);
nor U3549 (N_3549,In_1137,In_1406);
nand U3550 (N_3550,In_1387,In_988);
xnor U3551 (N_3551,In_988,In_219);
and U3552 (N_3552,In_1111,In_187);
nand U3553 (N_3553,In_1281,In_306);
and U3554 (N_3554,In_1352,In_1902);
xor U3555 (N_3555,In_571,In_1788);
or U3556 (N_3556,In_258,In_1632);
nor U3557 (N_3557,In_1923,In_1082);
xor U3558 (N_3558,In_212,In_1702);
nor U3559 (N_3559,In_1790,In_815);
xnor U3560 (N_3560,In_1251,In_70);
xor U3561 (N_3561,In_819,In_1827);
xor U3562 (N_3562,In_1546,In_739);
or U3563 (N_3563,In_275,In_1778);
nand U3564 (N_3564,In_674,In_1592);
and U3565 (N_3565,In_1194,In_1122);
xnor U3566 (N_3566,In_1707,In_1372);
or U3567 (N_3567,In_1707,In_1466);
or U3568 (N_3568,In_1643,In_1946);
xor U3569 (N_3569,In_1388,In_846);
or U3570 (N_3570,In_941,In_1213);
and U3571 (N_3571,In_332,In_106);
nand U3572 (N_3572,In_37,In_382);
nand U3573 (N_3573,In_368,In_210);
nor U3574 (N_3574,In_879,In_584);
nand U3575 (N_3575,In_1534,In_647);
xnor U3576 (N_3576,In_56,In_476);
or U3577 (N_3577,In_24,In_691);
xnor U3578 (N_3578,In_296,In_1362);
xnor U3579 (N_3579,In_1524,In_873);
xor U3580 (N_3580,In_1565,In_1491);
xnor U3581 (N_3581,In_1273,In_624);
or U3582 (N_3582,In_1606,In_1608);
and U3583 (N_3583,In_241,In_1067);
nor U3584 (N_3584,In_967,In_1945);
and U3585 (N_3585,In_1789,In_841);
nand U3586 (N_3586,In_472,In_1210);
xnor U3587 (N_3587,In_1994,In_828);
nand U3588 (N_3588,In_1092,In_112);
nor U3589 (N_3589,In_1045,In_1448);
and U3590 (N_3590,In_1054,In_1585);
and U3591 (N_3591,In_439,In_579);
and U3592 (N_3592,In_87,In_235);
or U3593 (N_3593,In_1519,In_145);
xnor U3594 (N_3594,In_1084,In_487);
nand U3595 (N_3595,In_730,In_609);
or U3596 (N_3596,In_390,In_1406);
nand U3597 (N_3597,In_1525,In_1724);
xnor U3598 (N_3598,In_1490,In_445);
and U3599 (N_3599,In_40,In_1396);
or U3600 (N_3600,In_1376,In_1330);
or U3601 (N_3601,In_1536,In_293);
xnor U3602 (N_3602,In_1942,In_1799);
nand U3603 (N_3603,In_956,In_1638);
or U3604 (N_3604,In_7,In_443);
and U3605 (N_3605,In_1607,In_489);
nand U3606 (N_3606,In_1537,In_1109);
xor U3607 (N_3607,In_1063,In_233);
nand U3608 (N_3608,In_1885,In_1104);
nor U3609 (N_3609,In_1919,In_1786);
xnor U3610 (N_3610,In_732,In_1132);
xnor U3611 (N_3611,In_1162,In_1505);
nand U3612 (N_3612,In_1806,In_1675);
xnor U3613 (N_3613,In_1071,In_480);
or U3614 (N_3614,In_1292,In_215);
nor U3615 (N_3615,In_1923,In_1100);
xor U3616 (N_3616,In_887,In_728);
nor U3617 (N_3617,In_177,In_632);
xnor U3618 (N_3618,In_1360,In_684);
and U3619 (N_3619,In_825,In_1741);
nor U3620 (N_3620,In_845,In_1479);
nor U3621 (N_3621,In_965,In_261);
or U3622 (N_3622,In_1009,In_1697);
nor U3623 (N_3623,In_999,In_336);
nand U3624 (N_3624,In_62,In_1790);
nor U3625 (N_3625,In_1480,In_191);
xor U3626 (N_3626,In_1574,In_811);
xor U3627 (N_3627,In_1092,In_567);
or U3628 (N_3628,In_996,In_2);
or U3629 (N_3629,In_542,In_1226);
nor U3630 (N_3630,In_759,In_58);
nand U3631 (N_3631,In_1518,In_1109);
xor U3632 (N_3632,In_1218,In_991);
and U3633 (N_3633,In_1162,In_712);
xor U3634 (N_3634,In_1249,In_77);
nand U3635 (N_3635,In_1870,In_922);
or U3636 (N_3636,In_1021,In_1864);
nand U3637 (N_3637,In_1140,In_137);
and U3638 (N_3638,In_1150,In_656);
nand U3639 (N_3639,In_1434,In_37);
nand U3640 (N_3640,In_1494,In_1914);
nand U3641 (N_3641,In_905,In_749);
nand U3642 (N_3642,In_872,In_1573);
nor U3643 (N_3643,In_1208,In_46);
and U3644 (N_3644,In_151,In_1911);
and U3645 (N_3645,In_1868,In_123);
or U3646 (N_3646,In_1450,In_1989);
or U3647 (N_3647,In_1574,In_943);
nor U3648 (N_3648,In_494,In_1548);
xor U3649 (N_3649,In_144,In_1544);
or U3650 (N_3650,In_576,In_1263);
or U3651 (N_3651,In_1468,In_1900);
or U3652 (N_3652,In_64,In_1603);
and U3653 (N_3653,In_948,In_1687);
and U3654 (N_3654,In_591,In_535);
nand U3655 (N_3655,In_688,In_349);
nor U3656 (N_3656,In_1603,In_681);
nand U3657 (N_3657,In_1292,In_1654);
nand U3658 (N_3658,In_57,In_1672);
nand U3659 (N_3659,In_1974,In_546);
xnor U3660 (N_3660,In_1101,In_661);
nand U3661 (N_3661,In_802,In_323);
or U3662 (N_3662,In_879,In_369);
or U3663 (N_3663,In_1439,In_531);
or U3664 (N_3664,In_658,In_304);
or U3665 (N_3665,In_1426,In_516);
xnor U3666 (N_3666,In_949,In_1533);
xor U3667 (N_3667,In_1250,In_221);
or U3668 (N_3668,In_421,In_1643);
nor U3669 (N_3669,In_1938,In_364);
or U3670 (N_3670,In_1849,In_757);
nor U3671 (N_3671,In_401,In_1241);
or U3672 (N_3672,In_964,In_40);
xnor U3673 (N_3673,In_1336,In_1613);
xnor U3674 (N_3674,In_1494,In_1402);
xnor U3675 (N_3675,In_449,In_1382);
nor U3676 (N_3676,In_240,In_372);
nand U3677 (N_3677,In_1986,In_957);
xnor U3678 (N_3678,In_1221,In_289);
xnor U3679 (N_3679,In_164,In_476);
and U3680 (N_3680,In_1889,In_884);
nand U3681 (N_3681,In_836,In_1024);
and U3682 (N_3682,In_1657,In_1862);
nor U3683 (N_3683,In_1645,In_284);
or U3684 (N_3684,In_82,In_324);
nand U3685 (N_3685,In_689,In_1665);
and U3686 (N_3686,In_128,In_1549);
and U3687 (N_3687,In_1581,In_1177);
nor U3688 (N_3688,In_1832,In_255);
and U3689 (N_3689,In_245,In_964);
or U3690 (N_3690,In_1605,In_768);
or U3691 (N_3691,In_71,In_219);
nand U3692 (N_3692,In_1056,In_587);
xor U3693 (N_3693,In_62,In_756);
and U3694 (N_3694,In_848,In_1821);
nand U3695 (N_3695,In_13,In_628);
and U3696 (N_3696,In_426,In_1706);
or U3697 (N_3697,In_198,In_1772);
nand U3698 (N_3698,In_489,In_1042);
xnor U3699 (N_3699,In_45,In_605);
or U3700 (N_3700,In_145,In_1370);
nor U3701 (N_3701,In_855,In_1129);
nor U3702 (N_3702,In_103,In_1809);
nand U3703 (N_3703,In_1634,In_170);
and U3704 (N_3704,In_938,In_332);
nand U3705 (N_3705,In_55,In_1047);
xnor U3706 (N_3706,In_599,In_440);
nand U3707 (N_3707,In_1883,In_176);
nand U3708 (N_3708,In_636,In_1122);
xnor U3709 (N_3709,In_99,In_191);
nand U3710 (N_3710,In_793,In_1481);
nor U3711 (N_3711,In_523,In_104);
xnor U3712 (N_3712,In_1669,In_1099);
or U3713 (N_3713,In_524,In_789);
nand U3714 (N_3714,In_1763,In_1982);
nor U3715 (N_3715,In_1914,In_1396);
nor U3716 (N_3716,In_1918,In_1253);
and U3717 (N_3717,In_1896,In_1498);
and U3718 (N_3718,In_1781,In_1002);
nand U3719 (N_3719,In_1411,In_1608);
xnor U3720 (N_3720,In_1861,In_478);
and U3721 (N_3721,In_926,In_1317);
nor U3722 (N_3722,In_1882,In_1256);
nand U3723 (N_3723,In_1273,In_1010);
nor U3724 (N_3724,In_1601,In_1728);
and U3725 (N_3725,In_288,In_990);
xnor U3726 (N_3726,In_226,In_655);
or U3727 (N_3727,In_874,In_745);
and U3728 (N_3728,In_628,In_1791);
and U3729 (N_3729,In_1586,In_118);
nor U3730 (N_3730,In_964,In_1650);
and U3731 (N_3731,In_629,In_749);
nor U3732 (N_3732,In_17,In_207);
xnor U3733 (N_3733,In_1133,In_1395);
nand U3734 (N_3734,In_1896,In_72);
or U3735 (N_3735,In_396,In_1994);
nor U3736 (N_3736,In_1861,In_543);
or U3737 (N_3737,In_1452,In_1032);
xnor U3738 (N_3738,In_67,In_788);
nand U3739 (N_3739,In_687,In_593);
or U3740 (N_3740,In_995,In_648);
and U3741 (N_3741,In_158,In_1864);
nor U3742 (N_3742,In_341,In_813);
or U3743 (N_3743,In_1926,In_1339);
or U3744 (N_3744,In_1722,In_224);
nand U3745 (N_3745,In_486,In_169);
and U3746 (N_3746,In_1797,In_1956);
xor U3747 (N_3747,In_744,In_1534);
nand U3748 (N_3748,In_1702,In_1150);
or U3749 (N_3749,In_1608,In_1328);
and U3750 (N_3750,In_1891,In_493);
or U3751 (N_3751,In_529,In_1665);
nor U3752 (N_3752,In_487,In_806);
and U3753 (N_3753,In_1116,In_794);
nor U3754 (N_3754,In_1061,In_497);
nor U3755 (N_3755,In_721,In_1517);
and U3756 (N_3756,In_1177,In_671);
nor U3757 (N_3757,In_311,In_1705);
xor U3758 (N_3758,In_825,In_1508);
and U3759 (N_3759,In_420,In_1003);
nor U3760 (N_3760,In_860,In_1782);
and U3761 (N_3761,In_1574,In_408);
nand U3762 (N_3762,In_166,In_1413);
nor U3763 (N_3763,In_259,In_1157);
and U3764 (N_3764,In_1030,In_1488);
nand U3765 (N_3765,In_950,In_215);
and U3766 (N_3766,In_658,In_1604);
nand U3767 (N_3767,In_1442,In_1527);
or U3768 (N_3768,In_1234,In_706);
xor U3769 (N_3769,In_1079,In_1491);
and U3770 (N_3770,In_778,In_1350);
and U3771 (N_3771,In_752,In_464);
nand U3772 (N_3772,In_321,In_1643);
nor U3773 (N_3773,In_467,In_1865);
or U3774 (N_3774,In_360,In_16);
xor U3775 (N_3775,In_425,In_633);
or U3776 (N_3776,In_1335,In_1286);
or U3777 (N_3777,In_1767,In_183);
nand U3778 (N_3778,In_1941,In_1263);
or U3779 (N_3779,In_277,In_864);
nand U3780 (N_3780,In_478,In_1207);
nand U3781 (N_3781,In_1093,In_579);
and U3782 (N_3782,In_562,In_1021);
and U3783 (N_3783,In_77,In_796);
nand U3784 (N_3784,In_1156,In_1350);
xor U3785 (N_3785,In_970,In_667);
nand U3786 (N_3786,In_521,In_716);
nand U3787 (N_3787,In_295,In_814);
or U3788 (N_3788,In_1381,In_1009);
nand U3789 (N_3789,In_1325,In_611);
nand U3790 (N_3790,In_118,In_1006);
nor U3791 (N_3791,In_539,In_1635);
or U3792 (N_3792,In_110,In_1180);
and U3793 (N_3793,In_1887,In_306);
or U3794 (N_3794,In_121,In_1379);
or U3795 (N_3795,In_662,In_571);
and U3796 (N_3796,In_1485,In_728);
nand U3797 (N_3797,In_322,In_171);
nand U3798 (N_3798,In_1771,In_975);
xor U3799 (N_3799,In_1685,In_785);
nor U3800 (N_3800,In_31,In_1264);
nand U3801 (N_3801,In_1735,In_1710);
xnor U3802 (N_3802,In_495,In_1180);
and U3803 (N_3803,In_472,In_1953);
or U3804 (N_3804,In_157,In_868);
nor U3805 (N_3805,In_1736,In_176);
or U3806 (N_3806,In_1929,In_268);
or U3807 (N_3807,In_454,In_822);
and U3808 (N_3808,In_179,In_1977);
or U3809 (N_3809,In_1853,In_1912);
nor U3810 (N_3810,In_1335,In_11);
xnor U3811 (N_3811,In_995,In_1896);
xnor U3812 (N_3812,In_237,In_1290);
or U3813 (N_3813,In_1476,In_1303);
and U3814 (N_3814,In_949,In_1174);
nor U3815 (N_3815,In_1252,In_337);
nor U3816 (N_3816,In_1275,In_654);
and U3817 (N_3817,In_822,In_1156);
nand U3818 (N_3818,In_488,In_1192);
nand U3819 (N_3819,In_770,In_1458);
and U3820 (N_3820,In_1705,In_114);
and U3821 (N_3821,In_232,In_1093);
nor U3822 (N_3822,In_1298,In_1702);
nor U3823 (N_3823,In_934,In_1204);
or U3824 (N_3824,In_18,In_831);
or U3825 (N_3825,In_1694,In_1426);
or U3826 (N_3826,In_332,In_1585);
and U3827 (N_3827,In_606,In_211);
xnor U3828 (N_3828,In_1835,In_1747);
nand U3829 (N_3829,In_1304,In_294);
nor U3830 (N_3830,In_34,In_475);
xor U3831 (N_3831,In_1126,In_1859);
xor U3832 (N_3832,In_597,In_554);
and U3833 (N_3833,In_809,In_1653);
nor U3834 (N_3834,In_1494,In_1100);
nor U3835 (N_3835,In_295,In_1);
xor U3836 (N_3836,In_1104,In_1278);
nand U3837 (N_3837,In_1717,In_1824);
xor U3838 (N_3838,In_826,In_1102);
nand U3839 (N_3839,In_1918,In_1457);
or U3840 (N_3840,In_1075,In_1083);
nand U3841 (N_3841,In_1255,In_399);
and U3842 (N_3842,In_1297,In_1435);
xnor U3843 (N_3843,In_32,In_203);
or U3844 (N_3844,In_1405,In_631);
or U3845 (N_3845,In_1926,In_17);
or U3846 (N_3846,In_78,In_880);
xnor U3847 (N_3847,In_716,In_1352);
nand U3848 (N_3848,In_639,In_738);
xnor U3849 (N_3849,In_1598,In_1193);
and U3850 (N_3850,In_346,In_1824);
nand U3851 (N_3851,In_595,In_520);
nand U3852 (N_3852,In_1132,In_206);
and U3853 (N_3853,In_1757,In_482);
nor U3854 (N_3854,In_1118,In_654);
nor U3855 (N_3855,In_1455,In_164);
and U3856 (N_3856,In_1387,In_589);
or U3857 (N_3857,In_1224,In_207);
and U3858 (N_3858,In_272,In_472);
nor U3859 (N_3859,In_417,In_66);
nor U3860 (N_3860,In_1764,In_1001);
or U3861 (N_3861,In_1878,In_1215);
xor U3862 (N_3862,In_867,In_946);
xor U3863 (N_3863,In_298,In_961);
xnor U3864 (N_3864,In_880,In_263);
and U3865 (N_3865,In_929,In_234);
nand U3866 (N_3866,In_595,In_5);
or U3867 (N_3867,In_1785,In_915);
xnor U3868 (N_3868,In_1942,In_1079);
and U3869 (N_3869,In_1004,In_1811);
nor U3870 (N_3870,In_1090,In_541);
and U3871 (N_3871,In_516,In_295);
xor U3872 (N_3872,In_1319,In_1183);
nand U3873 (N_3873,In_78,In_1668);
nand U3874 (N_3874,In_1641,In_501);
nand U3875 (N_3875,In_534,In_932);
and U3876 (N_3876,In_1306,In_328);
and U3877 (N_3877,In_1043,In_1704);
xor U3878 (N_3878,In_74,In_1397);
nor U3879 (N_3879,In_474,In_650);
and U3880 (N_3880,In_1142,In_1910);
or U3881 (N_3881,In_1800,In_1156);
xnor U3882 (N_3882,In_1864,In_1244);
nor U3883 (N_3883,In_1708,In_328);
and U3884 (N_3884,In_488,In_743);
nor U3885 (N_3885,In_436,In_957);
and U3886 (N_3886,In_29,In_465);
xor U3887 (N_3887,In_468,In_1431);
nand U3888 (N_3888,In_52,In_1415);
xor U3889 (N_3889,In_653,In_869);
xnor U3890 (N_3890,In_453,In_689);
or U3891 (N_3891,In_504,In_1511);
or U3892 (N_3892,In_1025,In_128);
nor U3893 (N_3893,In_1330,In_872);
nor U3894 (N_3894,In_849,In_1597);
nand U3895 (N_3895,In_1845,In_895);
nor U3896 (N_3896,In_629,In_1863);
or U3897 (N_3897,In_177,In_1454);
xor U3898 (N_3898,In_1223,In_1024);
xnor U3899 (N_3899,In_1781,In_1293);
nor U3900 (N_3900,In_1181,In_355);
and U3901 (N_3901,In_1082,In_346);
and U3902 (N_3902,In_1766,In_733);
or U3903 (N_3903,In_1111,In_1905);
nand U3904 (N_3904,In_602,In_1920);
xnor U3905 (N_3905,In_1978,In_10);
nor U3906 (N_3906,In_898,In_220);
or U3907 (N_3907,In_1653,In_1945);
or U3908 (N_3908,In_330,In_1838);
or U3909 (N_3909,In_460,In_252);
nand U3910 (N_3910,In_940,In_1616);
and U3911 (N_3911,In_1836,In_640);
nand U3912 (N_3912,In_1201,In_471);
nand U3913 (N_3913,In_1158,In_390);
or U3914 (N_3914,In_1020,In_248);
and U3915 (N_3915,In_1796,In_200);
nand U3916 (N_3916,In_1267,In_31);
or U3917 (N_3917,In_1141,In_739);
and U3918 (N_3918,In_949,In_1822);
or U3919 (N_3919,In_411,In_998);
and U3920 (N_3920,In_508,In_671);
nand U3921 (N_3921,In_1255,In_376);
xnor U3922 (N_3922,In_1695,In_704);
nor U3923 (N_3923,In_1716,In_514);
and U3924 (N_3924,In_1609,In_662);
nor U3925 (N_3925,In_1051,In_1215);
and U3926 (N_3926,In_939,In_1732);
nor U3927 (N_3927,In_470,In_1998);
xor U3928 (N_3928,In_1626,In_316);
and U3929 (N_3929,In_1234,In_533);
or U3930 (N_3930,In_872,In_1458);
nand U3931 (N_3931,In_439,In_681);
xor U3932 (N_3932,In_635,In_855);
or U3933 (N_3933,In_1420,In_1660);
xor U3934 (N_3934,In_580,In_794);
xnor U3935 (N_3935,In_702,In_1544);
nand U3936 (N_3936,In_1152,In_1858);
xor U3937 (N_3937,In_533,In_1430);
or U3938 (N_3938,In_967,In_1711);
or U3939 (N_3939,In_917,In_648);
xnor U3940 (N_3940,In_415,In_973);
or U3941 (N_3941,In_1546,In_326);
xor U3942 (N_3942,In_580,In_449);
or U3943 (N_3943,In_1236,In_1563);
and U3944 (N_3944,In_312,In_532);
or U3945 (N_3945,In_1201,In_1812);
nor U3946 (N_3946,In_996,In_1934);
or U3947 (N_3947,In_1707,In_476);
or U3948 (N_3948,In_943,In_1677);
and U3949 (N_3949,In_694,In_1389);
or U3950 (N_3950,In_636,In_1901);
nand U3951 (N_3951,In_1788,In_1159);
nand U3952 (N_3952,In_128,In_716);
xor U3953 (N_3953,In_1628,In_1787);
xor U3954 (N_3954,In_1806,In_1955);
and U3955 (N_3955,In_1866,In_1670);
nor U3956 (N_3956,In_1156,In_1003);
and U3957 (N_3957,In_1967,In_583);
and U3958 (N_3958,In_1618,In_376);
xor U3959 (N_3959,In_157,In_1072);
or U3960 (N_3960,In_1702,In_959);
nor U3961 (N_3961,In_1740,In_296);
xor U3962 (N_3962,In_1131,In_1225);
nand U3963 (N_3963,In_1861,In_123);
xor U3964 (N_3964,In_1494,In_48);
or U3965 (N_3965,In_634,In_653);
nor U3966 (N_3966,In_1020,In_116);
or U3967 (N_3967,In_1682,In_1469);
or U3968 (N_3968,In_41,In_1);
and U3969 (N_3969,In_601,In_817);
xnor U3970 (N_3970,In_734,In_569);
nand U3971 (N_3971,In_474,In_960);
xor U3972 (N_3972,In_320,In_569);
nand U3973 (N_3973,In_798,In_728);
and U3974 (N_3974,In_655,In_1005);
or U3975 (N_3975,In_862,In_1798);
nand U3976 (N_3976,In_1951,In_1651);
nor U3977 (N_3977,In_708,In_867);
or U3978 (N_3978,In_221,In_141);
nor U3979 (N_3979,In_1650,In_1444);
and U3980 (N_3980,In_1791,In_699);
or U3981 (N_3981,In_649,In_108);
nand U3982 (N_3982,In_1644,In_1005);
nor U3983 (N_3983,In_1270,In_502);
or U3984 (N_3984,In_1723,In_9);
or U3985 (N_3985,In_248,In_792);
xor U3986 (N_3986,In_1927,In_1864);
nand U3987 (N_3987,In_753,In_1756);
nand U3988 (N_3988,In_1716,In_896);
or U3989 (N_3989,In_1758,In_1919);
xnor U3990 (N_3990,In_795,In_936);
nand U3991 (N_3991,In_40,In_956);
nand U3992 (N_3992,In_226,In_1790);
nand U3993 (N_3993,In_795,In_961);
xnor U3994 (N_3994,In_1535,In_545);
nor U3995 (N_3995,In_159,In_697);
or U3996 (N_3996,In_1371,In_1145);
nor U3997 (N_3997,In_1021,In_756);
xor U3998 (N_3998,In_1542,In_1807);
nor U3999 (N_3999,In_937,In_1243);
nand U4000 (N_4000,In_1026,In_243);
and U4001 (N_4001,In_0,In_1418);
or U4002 (N_4002,In_587,In_615);
or U4003 (N_4003,In_1730,In_937);
xnor U4004 (N_4004,In_764,In_1111);
xnor U4005 (N_4005,In_1636,In_538);
or U4006 (N_4006,In_1002,In_1719);
nand U4007 (N_4007,In_187,In_1594);
or U4008 (N_4008,In_1955,In_1838);
xor U4009 (N_4009,In_1732,In_827);
nand U4010 (N_4010,In_727,In_739);
or U4011 (N_4011,In_335,In_927);
nor U4012 (N_4012,In_359,In_454);
xor U4013 (N_4013,In_1821,In_1555);
xnor U4014 (N_4014,In_1488,In_1908);
or U4015 (N_4015,In_1867,In_900);
nor U4016 (N_4016,In_815,In_461);
nor U4017 (N_4017,In_1265,In_1991);
nand U4018 (N_4018,In_1,In_665);
or U4019 (N_4019,In_930,In_1089);
or U4020 (N_4020,In_1641,In_1659);
nand U4021 (N_4021,In_888,In_953);
nand U4022 (N_4022,In_590,In_1096);
and U4023 (N_4023,In_1498,In_1253);
nor U4024 (N_4024,In_1171,In_1677);
xnor U4025 (N_4025,In_1252,In_1542);
xor U4026 (N_4026,In_1326,In_1041);
nor U4027 (N_4027,In_1187,In_43);
and U4028 (N_4028,In_539,In_1604);
xor U4029 (N_4029,In_1453,In_946);
and U4030 (N_4030,In_913,In_725);
or U4031 (N_4031,In_67,In_915);
or U4032 (N_4032,In_728,In_374);
or U4033 (N_4033,In_671,In_656);
and U4034 (N_4034,In_1715,In_730);
and U4035 (N_4035,In_583,In_216);
nor U4036 (N_4036,In_1770,In_745);
nor U4037 (N_4037,In_850,In_394);
nor U4038 (N_4038,In_1736,In_772);
nor U4039 (N_4039,In_98,In_661);
and U4040 (N_4040,In_217,In_1788);
or U4041 (N_4041,In_1294,In_707);
or U4042 (N_4042,In_183,In_9);
nor U4043 (N_4043,In_362,In_1286);
or U4044 (N_4044,In_119,In_1977);
nand U4045 (N_4045,In_1419,In_1245);
and U4046 (N_4046,In_1580,In_222);
and U4047 (N_4047,In_1390,In_1431);
or U4048 (N_4048,In_8,In_1916);
or U4049 (N_4049,In_178,In_1343);
or U4050 (N_4050,In_1289,In_1744);
and U4051 (N_4051,In_996,In_1263);
or U4052 (N_4052,In_748,In_357);
or U4053 (N_4053,In_58,In_1110);
or U4054 (N_4054,In_1553,In_1913);
xor U4055 (N_4055,In_100,In_393);
or U4056 (N_4056,In_787,In_1997);
nor U4057 (N_4057,In_470,In_991);
and U4058 (N_4058,In_1372,In_1069);
nand U4059 (N_4059,In_711,In_1534);
xor U4060 (N_4060,In_1127,In_1173);
or U4061 (N_4061,In_37,In_319);
nand U4062 (N_4062,In_1244,In_822);
nor U4063 (N_4063,In_1925,In_1187);
and U4064 (N_4064,In_1025,In_1114);
and U4065 (N_4065,In_954,In_589);
xor U4066 (N_4066,In_291,In_1004);
xnor U4067 (N_4067,In_64,In_1658);
or U4068 (N_4068,In_188,In_407);
and U4069 (N_4069,In_412,In_1933);
xnor U4070 (N_4070,In_1384,In_171);
and U4071 (N_4071,In_487,In_1000);
nand U4072 (N_4072,In_1021,In_1597);
nor U4073 (N_4073,In_1121,In_148);
nand U4074 (N_4074,In_1728,In_1619);
nand U4075 (N_4075,In_466,In_1400);
nor U4076 (N_4076,In_1179,In_1665);
nor U4077 (N_4077,In_874,In_1504);
and U4078 (N_4078,In_543,In_1947);
and U4079 (N_4079,In_1551,In_1056);
xnor U4080 (N_4080,In_1297,In_1325);
and U4081 (N_4081,In_63,In_224);
nand U4082 (N_4082,In_373,In_424);
nor U4083 (N_4083,In_1375,In_1043);
nand U4084 (N_4084,In_139,In_1054);
nor U4085 (N_4085,In_159,In_265);
nand U4086 (N_4086,In_1533,In_735);
and U4087 (N_4087,In_966,In_1134);
xor U4088 (N_4088,In_1774,In_670);
xor U4089 (N_4089,In_706,In_751);
nand U4090 (N_4090,In_1531,In_1422);
and U4091 (N_4091,In_1746,In_1356);
nor U4092 (N_4092,In_401,In_1345);
nor U4093 (N_4093,In_566,In_498);
nand U4094 (N_4094,In_1967,In_540);
xnor U4095 (N_4095,In_64,In_277);
or U4096 (N_4096,In_1958,In_210);
or U4097 (N_4097,In_693,In_1900);
and U4098 (N_4098,In_196,In_1645);
xor U4099 (N_4099,In_375,In_943);
and U4100 (N_4100,In_244,In_265);
xor U4101 (N_4101,In_118,In_772);
or U4102 (N_4102,In_652,In_1463);
nor U4103 (N_4103,In_1630,In_1418);
and U4104 (N_4104,In_990,In_1183);
nand U4105 (N_4105,In_1666,In_398);
nor U4106 (N_4106,In_599,In_82);
nor U4107 (N_4107,In_807,In_920);
nand U4108 (N_4108,In_1747,In_807);
xor U4109 (N_4109,In_1641,In_1388);
xor U4110 (N_4110,In_1512,In_412);
xor U4111 (N_4111,In_178,In_336);
or U4112 (N_4112,In_976,In_38);
nand U4113 (N_4113,In_1928,In_1277);
xor U4114 (N_4114,In_1507,In_1761);
nand U4115 (N_4115,In_712,In_1523);
and U4116 (N_4116,In_1287,In_1993);
xor U4117 (N_4117,In_1385,In_1634);
or U4118 (N_4118,In_1607,In_244);
nor U4119 (N_4119,In_606,In_250);
xnor U4120 (N_4120,In_97,In_1374);
and U4121 (N_4121,In_1916,In_742);
and U4122 (N_4122,In_747,In_1158);
or U4123 (N_4123,In_34,In_1045);
or U4124 (N_4124,In_329,In_1105);
or U4125 (N_4125,In_1824,In_921);
nor U4126 (N_4126,In_1412,In_370);
and U4127 (N_4127,In_858,In_163);
xnor U4128 (N_4128,In_975,In_725);
nor U4129 (N_4129,In_851,In_1489);
xnor U4130 (N_4130,In_1023,In_234);
and U4131 (N_4131,In_1476,In_1694);
or U4132 (N_4132,In_1768,In_408);
nand U4133 (N_4133,In_76,In_1469);
xor U4134 (N_4134,In_452,In_967);
xnor U4135 (N_4135,In_924,In_1843);
xnor U4136 (N_4136,In_905,In_268);
or U4137 (N_4137,In_1772,In_169);
or U4138 (N_4138,In_1690,In_1050);
nand U4139 (N_4139,In_346,In_639);
nor U4140 (N_4140,In_1489,In_526);
nor U4141 (N_4141,In_668,In_1225);
xor U4142 (N_4142,In_1317,In_1894);
or U4143 (N_4143,In_1725,In_1296);
nor U4144 (N_4144,In_1178,In_728);
or U4145 (N_4145,In_1917,In_1075);
xnor U4146 (N_4146,In_922,In_46);
nor U4147 (N_4147,In_1649,In_1672);
and U4148 (N_4148,In_253,In_840);
xnor U4149 (N_4149,In_700,In_844);
and U4150 (N_4150,In_1878,In_499);
or U4151 (N_4151,In_1914,In_1296);
nand U4152 (N_4152,In_1057,In_1308);
nand U4153 (N_4153,In_1644,In_617);
nor U4154 (N_4154,In_1419,In_1539);
nand U4155 (N_4155,In_1277,In_1504);
nor U4156 (N_4156,In_1796,In_300);
and U4157 (N_4157,In_1471,In_1225);
xnor U4158 (N_4158,In_1147,In_926);
nor U4159 (N_4159,In_224,In_30);
or U4160 (N_4160,In_8,In_755);
nand U4161 (N_4161,In_858,In_653);
and U4162 (N_4162,In_596,In_816);
or U4163 (N_4163,In_1209,In_879);
nand U4164 (N_4164,In_1144,In_1305);
xnor U4165 (N_4165,In_1798,In_1057);
nand U4166 (N_4166,In_1713,In_545);
or U4167 (N_4167,In_29,In_1792);
and U4168 (N_4168,In_461,In_408);
nor U4169 (N_4169,In_1671,In_961);
xor U4170 (N_4170,In_425,In_1368);
xnor U4171 (N_4171,In_1286,In_197);
nor U4172 (N_4172,In_800,In_359);
xnor U4173 (N_4173,In_1345,In_540);
and U4174 (N_4174,In_1906,In_543);
and U4175 (N_4175,In_625,In_1297);
or U4176 (N_4176,In_617,In_1776);
nor U4177 (N_4177,In_1014,In_101);
or U4178 (N_4178,In_985,In_236);
and U4179 (N_4179,In_1986,In_1015);
xor U4180 (N_4180,In_828,In_1692);
and U4181 (N_4181,In_1503,In_898);
or U4182 (N_4182,In_989,In_1164);
nor U4183 (N_4183,In_1226,In_842);
or U4184 (N_4184,In_140,In_484);
or U4185 (N_4185,In_2,In_183);
nor U4186 (N_4186,In_943,In_1828);
xor U4187 (N_4187,In_120,In_464);
nand U4188 (N_4188,In_1753,In_362);
xor U4189 (N_4189,In_1665,In_199);
nand U4190 (N_4190,In_1177,In_916);
xor U4191 (N_4191,In_1827,In_1426);
xnor U4192 (N_4192,In_1318,In_326);
nor U4193 (N_4193,In_105,In_1761);
or U4194 (N_4194,In_426,In_994);
nor U4195 (N_4195,In_130,In_871);
xnor U4196 (N_4196,In_1768,In_1821);
and U4197 (N_4197,In_1391,In_1318);
xor U4198 (N_4198,In_1838,In_1163);
and U4199 (N_4199,In_1322,In_1809);
or U4200 (N_4200,In_1576,In_771);
nor U4201 (N_4201,In_1032,In_813);
nor U4202 (N_4202,In_593,In_1644);
nor U4203 (N_4203,In_938,In_114);
or U4204 (N_4204,In_1004,In_1775);
and U4205 (N_4205,In_1,In_667);
nand U4206 (N_4206,In_1781,In_20);
and U4207 (N_4207,In_1650,In_1567);
nor U4208 (N_4208,In_354,In_69);
nor U4209 (N_4209,In_185,In_686);
xor U4210 (N_4210,In_610,In_1686);
xor U4211 (N_4211,In_992,In_491);
xor U4212 (N_4212,In_1147,In_917);
nor U4213 (N_4213,In_306,In_1960);
and U4214 (N_4214,In_16,In_225);
and U4215 (N_4215,In_1785,In_455);
nand U4216 (N_4216,In_1688,In_1127);
or U4217 (N_4217,In_926,In_1901);
and U4218 (N_4218,In_1452,In_649);
nand U4219 (N_4219,In_1539,In_1869);
or U4220 (N_4220,In_215,In_730);
nand U4221 (N_4221,In_794,In_1792);
xnor U4222 (N_4222,In_1685,In_335);
nor U4223 (N_4223,In_731,In_626);
nand U4224 (N_4224,In_1414,In_1569);
xnor U4225 (N_4225,In_618,In_765);
and U4226 (N_4226,In_93,In_1099);
and U4227 (N_4227,In_1649,In_35);
nor U4228 (N_4228,In_861,In_1650);
or U4229 (N_4229,In_822,In_314);
and U4230 (N_4230,In_1175,In_1539);
nand U4231 (N_4231,In_1176,In_1876);
xor U4232 (N_4232,In_1528,In_1608);
nand U4233 (N_4233,In_1691,In_1270);
and U4234 (N_4234,In_764,In_1783);
nor U4235 (N_4235,In_1040,In_1740);
xor U4236 (N_4236,In_150,In_919);
or U4237 (N_4237,In_1139,In_467);
xor U4238 (N_4238,In_789,In_848);
nor U4239 (N_4239,In_1183,In_1889);
xnor U4240 (N_4240,In_215,In_478);
and U4241 (N_4241,In_1113,In_1294);
nor U4242 (N_4242,In_370,In_103);
nand U4243 (N_4243,In_1681,In_1862);
and U4244 (N_4244,In_1507,In_1803);
xor U4245 (N_4245,In_135,In_1547);
nor U4246 (N_4246,In_575,In_232);
xnor U4247 (N_4247,In_1023,In_1225);
nand U4248 (N_4248,In_992,In_1562);
nor U4249 (N_4249,In_169,In_1047);
nor U4250 (N_4250,In_1520,In_665);
nand U4251 (N_4251,In_1333,In_1093);
nand U4252 (N_4252,In_1922,In_1113);
and U4253 (N_4253,In_201,In_304);
and U4254 (N_4254,In_492,In_1304);
nor U4255 (N_4255,In_1680,In_1810);
or U4256 (N_4256,In_78,In_1256);
nor U4257 (N_4257,In_1510,In_873);
or U4258 (N_4258,In_882,In_1265);
or U4259 (N_4259,In_1343,In_1591);
xnor U4260 (N_4260,In_1407,In_1977);
and U4261 (N_4261,In_1972,In_460);
nand U4262 (N_4262,In_955,In_1074);
nand U4263 (N_4263,In_119,In_823);
nor U4264 (N_4264,In_177,In_527);
or U4265 (N_4265,In_927,In_1739);
or U4266 (N_4266,In_555,In_862);
nand U4267 (N_4267,In_250,In_752);
nand U4268 (N_4268,In_666,In_1740);
nand U4269 (N_4269,In_1174,In_1340);
and U4270 (N_4270,In_827,In_578);
nand U4271 (N_4271,In_915,In_1102);
and U4272 (N_4272,In_439,In_834);
and U4273 (N_4273,In_1299,In_1744);
or U4274 (N_4274,In_1034,In_185);
nor U4275 (N_4275,In_138,In_1663);
or U4276 (N_4276,In_351,In_1329);
xor U4277 (N_4277,In_471,In_84);
and U4278 (N_4278,In_447,In_1688);
and U4279 (N_4279,In_868,In_340);
nor U4280 (N_4280,In_751,In_884);
and U4281 (N_4281,In_1213,In_525);
and U4282 (N_4282,In_1523,In_125);
and U4283 (N_4283,In_1593,In_17);
or U4284 (N_4284,In_1242,In_138);
or U4285 (N_4285,In_626,In_1591);
nor U4286 (N_4286,In_536,In_1592);
nor U4287 (N_4287,In_428,In_1631);
nor U4288 (N_4288,In_79,In_769);
xor U4289 (N_4289,In_1002,In_149);
xnor U4290 (N_4290,In_1237,In_1446);
and U4291 (N_4291,In_828,In_1301);
and U4292 (N_4292,In_1832,In_107);
or U4293 (N_4293,In_1707,In_1324);
and U4294 (N_4294,In_825,In_1617);
nand U4295 (N_4295,In_709,In_804);
nor U4296 (N_4296,In_605,In_996);
xor U4297 (N_4297,In_508,In_1925);
or U4298 (N_4298,In_19,In_1545);
or U4299 (N_4299,In_1732,In_719);
nor U4300 (N_4300,In_1860,In_239);
nand U4301 (N_4301,In_620,In_824);
nor U4302 (N_4302,In_1449,In_1301);
nor U4303 (N_4303,In_628,In_1070);
or U4304 (N_4304,In_313,In_643);
or U4305 (N_4305,In_686,In_504);
nor U4306 (N_4306,In_1612,In_502);
nand U4307 (N_4307,In_784,In_995);
and U4308 (N_4308,In_1781,In_516);
and U4309 (N_4309,In_1908,In_637);
or U4310 (N_4310,In_1616,In_1039);
nand U4311 (N_4311,In_247,In_1307);
xor U4312 (N_4312,In_1449,In_573);
nor U4313 (N_4313,In_1097,In_418);
nand U4314 (N_4314,In_1142,In_763);
and U4315 (N_4315,In_289,In_460);
and U4316 (N_4316,In_1710,In_228);
nand U4317 (N_4317,In_772,In_237);
and U4318 (N_4318,In_1202,In_88);
xor U4319 (N_4319,In_1230,In_1321);
and U4320 (N_4320,In_510,In_497);
xor U4321 (N_4321,In_1420,In_800);
and U4322 (N_4322,In_1587,In_319);
or U4323 (N_4323,In_1901,In_917);
or U4324 (N_4324,In_826,In_1352);
nand U4325 (N_4325,In_1733,In_414);
or U4326 (N_4326,In_1130,In_1548);
xnor U4327 (N_4327,In_1949,In_1163);
nand U4328 (N_4328,In_73,In_949);
xor U4329 (N_4329,In_1531,In_485);
nand U4330 (N_4330,In_66,In_1825);
or U4331 (N_4331,In_1853,In_354);
and U4332 (N_4332,In_1246,In_273);
nand U4333 (N_4333,In_438,In_247);
or U4334 (N_4334,In_580,In_635);
and U4335 (N_4335,In_950,In_408);
or U4336 (N_4336,In_729,In_418);
and U4337 (N_4337,In_1847,In_1268);
or U4338 (N_4338,In_981,In_843);
nor U4339 (N_4339,In_440,In_1715);
nand U4340 (N_4340,In_811,In_1239);
nand U4341 (N_4341,In_1365,In_1635);
or U4342 (N_4342,In_1411,In_1526);
xnor U4343 (N_4343,In_584,In_1602);
and U4344 (N_4344,In_1177,In_1566);
nand U4345 (N_4345,In_1946,In_788);
or U4346 (N_4346,In_859,In_1743);
xnor U4347 (N_4347,In_506,In_1446);
or U4348 (N_4348,In_1479,In_704);
nor U4349 (N_4349,In_1683,In_356);
or U4350 (N_4350,In_810,In_734);
and U4351 (N_4351,In_608,In_266);
and U4352 (N_4352,In_40,In_142);
or U4353 (N_4353,In_1847,In_807);
and U4354 (N_4354,In_1749,In_760);
and U4355 (N_4355,In_1547,In_1289);
or U4356 (N_4356,In_1377,In_1163);
nor U4357 (N_4357,In_1827,In_1126);
nand U4358 (N_4358,In_1602,In_1658);
xnor U4359 (N_4359,In_10,In_840);
or U4360 (N_4360,In_1289,In_1876);
nor U4361 (N_4361,In_1357,In_1661);
xnor U4362 (N_4362,In_1104,In_1715);
nand U4363 (N_4363,In_722,In_947);
nor U4364 (N_4364,In_1181,In_1856);
nor U4365 (N_4365,In_1329,In_539);
or U4366 (N_4366,In_1984,In_1630);
or U4367 (N_4367,In_87,In_1336);
nor U4368 (N_4368,In_289,In_1142);
nor U4369 (N_4369,In_732,In_809);
and U4370 (N_4370,In_1429,In_37);
and U4371 (N_4371,In_1659,In_1445);
xnor U4372 (N_4372,In_622,In_1020);
nor U4373 (N_4373,In_111,In_379);
xor U4374 (N_4374,In_1201,In_1688);
or U4375 (N_4375,In_1268,In_1936);
xor U4376 (N_4376,In_958,In_624);
and U4377 (N_4377,In_1504,In_1357);
nor U4378 (N_4378,In_1671,In_1947);
xnor U4379 (N_4379,In_994,In_1187);
or U4380 (N_4380,In_1642,In_1782);
or U4381 (N_4381,In_1046,In_948);
nand U4382 (N_4382,In_1365,In_549);
or U4383 (N_4383,In_1062,In_276);
xor U4384 (N_4384,In_1267,In_332);
nand U4385 (N_4385,In_402,In_300);
and U4386 (N_4386,In_1752,In_1825);
nand U4387 (N_4387,In_82,In_974);
and U4388 (N_4388,In_1759,In_1855);
or U4389 (N_4389,In_618,In_695);
and U4390 (N_4390,In_202,In_1074);
xnor U4391 (N_4391,In_1735,In_1625);
nor U4392 (N_4392,In_12,In_357);
xor U4393 (N_4393,In_973,In_1212);
nand U4394 (N_4394,In_907,In_805);
and U4395 (N_4395,In_148,In_1281);
nand U4396 (N_4396,In_304,In_1978);
and U4397 (N_4397,In_1015,In_816);
nor U4398 (N_4398,In_1601,In_1522);
or U4399 (N_4399,In_500,In_116);
and U4400 (N_4400,In_1285,In_981);
and U4401 (N_4401,In_723,In_468);
xor U4402 (N_4402,In_1137,In_693);
xor U4403 (N_4403,In_114,In_465);
and U4404 (N_4404,In_1006,In_166);
nand U4405 (N_4405,In_89,In_1511);
xnor U4406 (N_4406,In_5,In_677);
nand U4407 (N_4407,In_861,In_651);
xnor U4408 (N_4408,In_625,In_1426);
or U4409 (N_4409,In_1479,In_732);
or U4410 (N_4410,In_1777,In_1096);
nor U4411 (N_4411,In_1120,In_1141);
and U4412 (N_4412,In_1844,In_934);
xor U4413 (N_4413,In_118,In_1910);
and U4414 (N_4414,In_1696,In_1785);
xor U4415 (N_4415,In_1892,In_893);
xnor U4416 (N_4416,In_1739,In_911);
nand U4417 (N_4417,In_1782,In_52);
nor U4418 (N_4418,In_87,In_1530);
or U4419 (N_4419,In_1185,In_691);
and U4420 (N_4420,In_652,In_1275);
nor U4421 (N_4421,In_707,In_396);
nand U4422 (N_4422,In_779,In_1348);
nor U4423 (N_4423,In_1237,In_779);
or U4424 (N_4424,In_242,In_1460);
nor U4425 (N_4425,In_462,In_821);
nor U4426 (N_4426,In_238,In_690);
nand U4427 (N_4427,In_114,In_1391);
nor U4428 (N_4428,In_430,In_1995);
and U4429 (N_4429,In_664,In_224);
nand U4430 (N_4430,In_1832,In_587);
and U4431 (N_4431,In_248,In_804);
and U4432 (N_4432,In_1648,In_1828);
xor U4433 (N_4433,In_1740,In_1816);
xor U4434 (N_4434,In_1779,In_419);
or U4435 (N_4435,In_1431,In_1701);
nand U4436 (N_4436,In_15,In_1371);
nor U4437 (N_4437,In_44,In_1610);
and U4438 (N_4438,In_907,In_540);
nand U4439 (N_4439,In_999,In_1276);
xnor U4440 (N_4440,In_1744,In_1543);
xor U4441 (N_4441,In_599,In_632);
xnor U4442 (N_4442,In_1864,In_1356);
nor U4443 (N_4443,In_312,In_123);
nor U4444 (N_4444,In_591,In_1321);
nor U4445 (N_4445,In_482,In_1863);
xor U4446 (N_4446,In_604,In_877);
xor U4447 (N_4447,In_1153,In_660);
or U4448 (N_4448,In_1530,In_1320);
or U4449 (N_4449,In_771,In_97);
nand U4450 (N_4450,In_1519,In_1664);
nor U4451 (N_4451,In_1548,In_1831);
nor U4452 (N_4452,In_248,In_1771);
and U4453 (N_4453,In_905,In_1474);
nor U4454 (N_4454,In_931,In_1347);
xor U4455 (N_4455,In_1886,In_259);
nand U4456 (N_4456,In_1951,In_1338);
nand U4457 (N_4457,In_1808,In_1727);
and U4458 (N_4458,In_1690,In_1125);
or U4459 (N_4459,In_1787,In_1827);
and U4460 (N_4460,In_1656,In_456);
or U4461 (N_4461,In_1471,In_1886);
nor U4462 (N_4462,In_917,In_1206);
nand U4463 (N_4463,In_945,In_418);
xnor U4464 (N_4464,In_1426,In_871);
nor U4465 (N_4465,In_1917,In_1863);
nand U4466 (N_4466,In_510,In_881);
xor U4467 (N_4467,In_1270,In_808);
xnor U4468 (N_4468,In_564,In_152);
nand U4469 (N_4469,In_595,In_1286);
xnor U4470 (N_4470,In_1907,In_1123);
and U4471 (N_4471,In_1722,In_891);
nand U4472 (N_4472,In_1767,In_673);
or U4473 (N_4473,In_599,In_1849);
xor U4474 (N_4474,In_458,In_827);
xor U4475 (N_4475,In_1156,In_278);
nand U4476 (N_4476,In_1953,In_1948);
xnor U4477 (N_4477,In_101,In_184);
nor U4478 (N_4478,In_248,In_151);
nand U4479 (N_4479,In_212,In_564);
or U4480 (N_4480,In_1729,In_24);
xor U4481 (N_4481,In_1032,In_1022);
nand U4482 (N_4482,In_68,In_520);
nor U4483 (N_4483,In_1097,In_1282);
nor U4484 (N_4484,In_1420,In_1722);
nor U4485 (N_4485,In_1233,In_1137);
xor U4486 (N_4486,In_1078,In_732);
or U4487 (N_4487,In_636,In_1838);
xor U4488 (N_4488,In_1892,In_827);
or U4489 (N_4489,In_771,In_94);
nor U4490 (N_4490,In_139,In_1087);
nor U4491 (N_4491,In_1640,In_964);
and U4492 (N_4492,In_1603,In_1631);
nor U4493 (N_4493,In_909,In_338);
and U4494 (N_4494,In_1558,In_1583);
nand U4495 (N_4495,In_239,In_559);
nor U4496 (N_4496,In_1759,In_1847);
and U4497 (N_4497,In_1214,In_1743);
nand U4498 (N_4498,In_1111,In_224);
nand U4499 (N_4499,In_1404,In_1960);
nor U4500 (N_4500,In_1468,In_1476);
nand U4501 (N_4501,In_1491,In_1126);
and U4502 (N_4502,In_246,In_1908);
nor U4503 (N_4503,In_399,In_1469);
nor U4504 (N_4504,In_1650,In_61);
and U4505 (N_4505,In_1193,In_322);
xnor U4506 (N_4506,In_1556,In_271);
xnor U4507 (N_4507,In_1728,In_1898);
xor U4508 (N_4508,In_492,In_199);
xnor U4509 (N_4509,In_525,In_387);
or U4510 (N_4510,In_1718,In_634);
xor U4511 (N_4511,In_1856,In_303);
xnor U4512 (N_4512,In_1296,In_1352);
or U4513 (N_4513,In_93,In_1979);
nand U4514 (N_4514,In_243,In_1378);
nor U4515 (N_4515,In_300,In_1427);
and U4516 (N_4516,In_1753,In_1119);
nor U4517 (N_4517,In_76,In_1818);
nand U4518 (N_4518,In_289,In_73);
nor U4519 (N_4519,In_58,In_1024);
nor U4520 (N_4520,In_696,In_517);
and U4521 (N_4521,In_1433,In_948);
nor U4522 (N_4522,In_39,In_488);
and U4523 (N_4523,In_874,In_813);
nand U4524 (N_4524,In_1311,In_619);
nor U4525 (N_4525,In_1692,In_381);
and U4526 (N_4526,In_481,In_236);
xor U4527 (N_4527,In_479,In_781);
xor U4528 (N_4528,In_1652,In_1080);
xnor U4529 (N_4529,In_421,In_1043);
nand U4530 (N_4530,In_1520,In_125);
and U4531 (N_4531,In_1790,In_1988);
or U4532 (N_4532,In_1404,In_435);
nor U4533 (N_4533,In_1394,In_819);
or U4534 (N_4534,In_1981,In_1574);
nor U4535 (N_4535,In_629,In_1370);
and U4536 (N_4536,In_461,In_386);
nand U4537 (N_4537,In_1018,In_1380);
and U4538 (N_4538,In_1529,In_788);
and U4539 (N_4539,In_1062,In_1010);
xor U4540 (N_4540,In_142,In_1632);
and U4541 (N_4541,In_187,In_1861);
or U4542 (N_4542,In_1426,In_290);
or U4543 (N_4543,In_1012,In_52);
and U4544 (N_4544,In_1086,In_1364);
nor U4545 (N_4545,In_1240,In_1939);
nor U4546 (N_4546,In_1676,In_358);
and U4547 (N_4547,In_970,In_1450);
xor U4548 (N_4548,In_1289,In_354);
nand U4549 (N_4549,In_1495,In_713);
and U4550 (N_4550,In_1681,In_1563);
nor U4551 (N_4551,In_1670,In_1238);
or U4552 (N_4552,In_40,In_624);
nor U4553 (N_4553,In_167,In_1205);
nand U4554 (N_4554,In_135,In_1928);
nor U4555 (N_4555,In_781,In_414);
nor U4556 (N_4556,In_1501,In_209);
or U4557 (N_4557,In_904,In_1204);
or U4558 (N_4558,In_1039,In_1802);
or U4559 (N_4559,In_1591,In_733);
or U4560 (N_4560,In_1100,In_444);
or U4561 (N_4561,In_142,In_559);
nor U4562 (N_4562,In_772,In_1839);
xor U4563 (N_4563,In_1453,In_747);
or U4564 (N_4564,In_628,In_916);
or U4565 (N_4565,In_1629,In_1478);
xor U4566 (N_4566,In_455,In_279);
or U4567 (N_4567,In_177,In_1385);
xor U4568 (N_4568,In_1152,In_396);
or U4569 (N_4569,In_1647,In_35);
and U4570 (N_4570,In_358,In_369);
xor U4571 (N_4571,In_1712,In_563);
nand U4572 (N_4572,In_1998,In_921);
nand U4573 (N_4573,In_1138,In_1518);
nand U4574 (N_4574,In_1779,In_278);
nor U4575 (N_4575,In_1855,In_281);
and U4576 (N_4576,In_1509,In_322);
nand U4577 (N_4577,In_1731,In_1983);
nor U4578 (N_4578,In_1783,In_352);
nand U4579 (N_4579,In_1546,In_1849);
nor U4580 (N_4580,In_779,In_674);
and U4581 (N_4581,In_1208,In_1089);
xor U4582 (N_4582,In_1544,In_553);
or U4583 (N_4583,In_700,In_486);
nand U4584 (N_4584,In_872,In_1350);
or U4585 (N_4585,In_1587,In_862);
and U4586 (N_4586,In_162,In_849);
xor U4587 (N_4587,In_971,In_716);
xor U4588 (N_4588,In_983,In_684);
xnor U4589 (N_4589,In_0,In_142);
nor U4590 (N_4590,In_934,In_1359);
nand U4591 (N_4591,In_1488,In_1544);
nand U4592 (N_4592,In_677,In_941);
or U4593 (N_4593,In_1691,In_1609);
nor U4594 (N_4594,In_67,In_233);
xnor U4595 (N_4595,In_1691,In_1340);
nor U4596 (N_4596,In_1687,In_916);
xor U4597 (N_4597,In_1753,In_1663);
nand U4598 (N_4598,In_411,In_469);
and U4599 (N_4599,In_41,In_401);
nand U4600 (N_4600,In_1914,In_1285);
and U4601 (N_4601,In_110,In_1945);
nand U4602 (N_4602,In_21,In_168);
xor U4603 (N_4603,In_1492,In_1896);
and U4604 (N_4604,In_978,In_694);
or U4605 (N_4605,In_490,In_1788);
xnor U4606 (N_4606,In_1053,In_1346);
nand U4607 (N_4607,In_371,In_1184);
and U4608 (N_4608,In_335,In_1722);
nand U4609 (N_4609,In_1515,In_1239);
xor U4610 (N_4610,In_318,In_1894);
xor U4611 (N_4611,In_1267,In_241);
nand U4612 (N_4612,In_329,In_1654);
nand U4613 (N_4613,In_936,In_302);
or U4614 (N_4614,In_1311,In_57);
and U4615 (N_4615,In_328,In_1019);
and U4616 (N_4616,In_427,In_65);
nor U4617 (N_4617,In_788,In_318);
nor U4618 (N_4618,In_1940,In_216);
and U4619 (N_4619,In_1627,In_528);
xnor U4620 (N_4620,In_316,In_1678);
nand U4621 (N_4621,In_404,In_586);
xor U4622 (N_4622,In_793,In_486);
xnor U4623 (N_4623,In_576,In_244);
nand U4624 (N_4624,In_1864,In_1619);
nand U4625 (N_4625,In_476,In_1640);
nor U4626 (N_4626,In_152,In_966);
nand U4627 (N_4627,In_1844,In_1204);
nor U4628 (N_4628,In_1629,In_27);
or U4629 (N_4629,In_1526,In_305);
xnor U4630 (N_4630,In_1534,In_1927);
xnor U4631 (N_4631,In_161,In_296);
nand U4632 (N_4632,In_655,In_1619);
xnor U4633 (N_4633,In_444,In_1747);
or U4634 (N_4634,In_110,In_58);
and U4635 (N_4635,In_1856,In_234);
nand U4636 (N_4636,In_11,In_1005);
nand U4637 (N_4637,In_1564,In_1277);
or U4638 (N_4638,In_1554,In_1588);
or U4639 (N_4639,In_1317,In_520);
nor U4640 (N_4640,In_297,In_675);
xor U4641 (N_4641,In_1900,In_1924);
xnor U4642 (N_4642,In_1221,In_1382);
and U4643 (N_4643,In_917,In_743);
and U4644 (N_4644,In_237,In_83);
nand U4645 (N_4645,In_1852,In_1831);
nor U4646 (N_4646,In_1906,In_1736);
or U4647 (N_4647,In_1526,In_666);
nor U4648 (N_4648,In_717,In_1708);
and U4649 (N_4649,In_1121,In_1028);
xor U4650 (N_4650,In_641,In_594);
and U4651 (N_4651,In_353,In_1594);
or U4652 (N_4652,In_17,In_1946);
xnor U4653 (N_4653,In_722,In_1940);
xnor U4654 (N_4654,In_1955,In_526);
or U4655 (N_4655,In_451,In_1960);
or U4656 (N_4656,In_494,In_1541);
and U4657 (N_4657,In_418,In_1910);
nand U4658 (N_4658,In_1730,In_1578);
or U4659 (N_4659,In_1770,In_1197);
xnor U4660 (N_4660,In_1562,In_35);
xnor U4661 (N_4661,In_938,In_1043);
nand U4662 (N_4662,In_1496,In_1000);
nand U4663 (N_4663,In_1413,In_1627);
xnor U4664 (N_4664,In_705,In_1192);
nand U4665 (N_4665,In_753,In_1159);
xor U4666 (N_4666,In_231,In_1412);
and U4667 (N_4667,In_1931,In_538);
xnor U4668 (N_4668,In_1177,In_1456);
and U4669 (N_4669,In_281,In_491);
and U4670 (N_4670,In_1001,In_1188);
and U4671 (N_4671,In_202,In_414);
and U4672 (N_4672,In_1454,In_392);
xor U4673 (N_4673,In_1507,In_1832);
nand U4674 (N_4674,In_1623,In_1601);
nor U4675 (N_4675,In_944,In_1792);
xnor U4676 (N_4676,In_186,In_787);
nand U4677 (N_4677,In_260,In_1632);
nor U4678 (N_4678,In_570,In_766);
and U4679 (N_4679,In_1290,In_1646);
nand U4680 (N_4680,In_1515,In_1499);
or U4681 (N_4681,In_1800,In_408);
nor U4682 (N_4682,In_805,In_1810);
or U4683 (N_4683,In_1925,In_1104);
or U4684 (N_4684,In_660,In_1532);
or U4685 (N_4685,In_527,In_1720);
or U4686 (N_4686,In_423,In_856);
nor U4687 (N_4687,In_1857,In_720);
nand U4688 (N_4688,In_1141,In_485);
xor U4689 (N_4689,In_351,In_1306);
nor U4690 (N_4690,In_1654,In_1451);
nor U4691 (N_4691,In_323,In_1388);
or U4692 (N_4692,In_558,In_549);
xnor U4693 (N_4693,In_427,In_1540);
xor U4694 (N_4694,In_852,In_718);
xnor U4695 (N_4695,In_1673,In_1298);
or U4696 (N_4696,In_80,In_1037);
nand U4697 (N_4697,In_1523,In_924);
or U4698 (N_4698,In_1258,In_426);
nor U4699 (N_4699,In_310,In_134);
xnor U4700 (N_4700,In_1657,In_1878);
nand U4701 (N_4701,In_1869,In_356);
nand U4702 (N_4702,In_45,In_1201);
nor U4703 (N_4703,In_489,In_2);
or U4704 (N_4704,In_1567,In_918);
and U4705 (N_4705,In_950,In_183);
or U4706 (N_4706,In_1622,In_133);
nand U4707 (N_4707,In_155,In_493);
and U4708 (N_4708,In_237,In_336);
nor U4709 (N_4709,In_258,In_497);
xor U4710 (N_4710,In_550,In_1188);
and U4711 (N_4711,In_7,In_1258);
xor U4712 (N_4712,In_1133,In_577);
or U4713 (N_4713,In_1428,In_1456);
xnor U4714 (N_4714,In_300,In_1188);
xnor U4715 (N_4715,In_1339,In_569);
nor U4716 (N_4716,In_136,In_776);
and U4717 (N_4717,In_1050,In_823);
nand U4718 (N_4718,In_11,In_1620);
or U4719 (N_4719,In_437,In_1375);
xor U4720 (N_4720,In_1789,In_1617);
nand U4721 (N_4721,In_531,In_1430);
and U4722 (N_4722,In_476,In_274);
nand U4723 (N_4723,In_92,In_1948);
nor U4724 (N_4724,In_291,In_130);
nand U4725 (N_4725,In_10,In_125);
nor U4726 (N_4726,In_1764,In_408);
or U4727 (N_4727,In_1307,In_5);
nand U4728 (N_4728,In_1164,In_1633);
and U4729 (N_4729,In_662,In_1236);
nor U4730 (N_4730,In_701,In_745);
nand U4731 (N_4731,In_742,In_675);
xnor U4732 (N_4732,In_954,In_811);
nor U4733 (N_4733,In_1658,In_767);
xor U4734 (N_4734,In_34,In_783);
or U4735 (N_4735,In_1278,In_1542);
or U4736 (N_4736,In_469,In_523);
nor U4737 (N_4737,In_172,In_1674);
and U4738 (N_4738,In_1097,In_199);
or U4739 (N_4739,In_1833,In_1464);
xor U4740 (N_4740,In_446,In_1580);
and U4741 (N_4741,In_1584,In_1053);
nor U4742 (N_4742,In_898,In_1604);
and U4743 (N_4743,In_1752,In_1894);
xnor U4744 (N_4744,In_0,In_1935);
nor U4745 (N_4745,In_206,In_440);
xnor U4746 (N_4746,In_1511,In_536);
and U4747 (N_4747,In_1411,In_1974);
and U4748 (N_4748,In_1636,In_66);
and U4749 (N_4749,In_102,In_90);
xor U4750 (N_4750,In_548,In_1882);
xnor U4751 (N_4751,In_283,In_1604);
and U4752 (N_4752,In_459,In_1984);
nand U4753 (N_4753,In_777,In_1448);
nand U4754 (N_4754,In_132,In_96);
and U4755 (N_4755,In_705,In_232);
nor U4756 (N_4756,In_456,In_1165);
nand U4757 (N_4757,In_972,In_1490);
and U4758 (N_4758,In_1539,In_64);
and U4759 (N_4759,In_1329,In_1335);
or U4760 (N_4760,In_1160,In_1210);
xnor U4761 (N_4761,In_1214,In_565);
xnor U4762 (N_4762,In_74,In_56);
nand U4763 (N_4763,In_1252,In_342);
nor U4764 (N_4764,In_1463,In_346);
nor U4765 (N_4765,In_550,In_135);
nand U4766 (N_4766,In_867,In_1946);
xor U4767 (N_4767,In_298,In_1029);
nor U4768 (N_4768,In_218,In_1920);
nand U4769 (N_4769,In_102,In_1737);
xnor U4770 (N_4770,In_514,In_1652);
nand U4771 (N_4771,In_994,In_1731);
nor U4772 (N_4772,In_1823,In_1931);
or U4773 (N_4773,In_1378,In_199);
and U4774 (N_4774,In_611,In_683);
nor U4775 (N_4775,In_1602,In_1612);
nand U4776 (N_4776,In_1609,In_1981);
or U4777 (N_4777,In_1621,In_998);
nor U4778 (N_4778,In_1849,In_924);
or U4779 (N_4779,In_1120,In_1022);
nor U4780 (N_4780,In_1772,In_877);
xor U4781 (N_4781,In_1902,In_762);
nand U4782 (N_4782,In_976,In_532);
nand U4783 (N_4783,In_285,In_1466);
nor U4784 (N_4784,In_320,In_1616);
xnor U4785 (N_4785,In_679,In_1322);
nor U4786 (N_4786,In_1421,In_1123);
and U4787 (N_4787,In_306,In_663);
xnor U4788 (N_4788,In_1875,In_1146);
xor U4789 (N_4789,In_1196,In_1153);
xor U4790 (N_4790,In_172,In_637);
and U4791 (N_4791,In_791,In_364);
xnor U4792 (N_4792,In_748,In_1187);
or U4793 (N_4793,In_558,In_1356);
nor U4794 (N_4794,In_1439,In_1016);
nand U4795 (N_4795,In_888,In_411);
nor U4796 (N_4796,In_1439,In_25);
and U4797 (N_4797,In_1732,In_1833);
nand U4798 (N_4798,In_1794,In_1924);
xor U4799 (N_4799,In_517,In_1249);
and U4800 (N_4800,In_132,In_23);
and U4801 (N_4801,In_1645,In_730);
nor U4802 (N_4802,In_254,In_1271);
xor U4803 (N_4803,In_133,In_625);
nand U4804 (N_4804,In_935,In_937);
and U4805 (N_4805,In_1863,In_545);
nand U4806 (N_4806,In_734,In_1782);
xor U4807 (N_4807,In_1492,In_1295);
nand U4808 (N_4808,In_1174,In_562);
and U4809 (N_4809,In_284,In_1938);
or U4810 (N_4810,In_1083,In_346);
nor U4811 (N_4811,In_750,In_1558);
or U4812 (N_4812,In_1958,In_662);
or U4813 (N_4813,In_1803,In_118);
nor U4814 (N_4814,In_1887,In_1038);
or U4815 (N_4815,In_335,In_1076);
and U4816 (N_4816,In_1702,In_1606);
and U4817 (N_4817,In_170,In_1384);
nor U4818 (N_4818,In_885,In_1162);
nand U4819 (N_4819,In_952,In_181);
nor U4820 (N_4820,In_826,In_173);
xor U4821 (N_4821,In_16,In_295);
nand U4822 (N_4822,In_1803,In_1008);
xnor U4823 (N_4823,In_448,In_1348);
xnor U4824 (N_4824,In_1517,In_645);
xnor U4825 (N_4825,In_1427,In_1488);
nor U4826 (N_4826,In_99,In_501);
nand U4827 (N_4827,In_1276,In_1456);
nor U4828 (N_4828,In_1260,In_1601);
xor U4829 (N_4829,In_911,In_1670);
or U4830 (N_4830,In_191,In_1020);
nor U4831 (N_4831,In_669,In_166);
and U4832 (N_4832,In_1186,In_1500);
nor U4833 (N_4833,In_1396,In_1495);
nand U4834 (N_4834,In_37,In_1964);
or U4835 (N_4835,In_961,In_518);
nor U4836 (N_4836,In_607,In_178);
or U4837 (N_4837,In_1087,In_1693);
and U4838 (N_4838,In_374,In_1742);
nor U4839 (N_4839,In_458,In_1811);
xor U4840 (N_4840,In_1652,In_703);
nor U4841 (N_4841,In_473,In_550);
or U4842 (N_4842,In_1959,In_1854);
nand U4843 (N_4843,In_1698,In_1760);
nand U4844 (N_4844,In_1575,In_735);
and U4845 (N_4845,In_672,In_582);
and U4846 (N_4846,In_1201,In_612);
xnor U4847 (N_4847,In_858,In_888);
nor U4848 (N_4848,In_1213,In_223);
or U4849 (N_4849,In_1460,In_951);
nand U4850 (N_4850,In_1655,In_1594);
nand U4851 (N_4851,In_159,In_195);
nand U4852 (N_4852,In_1956,In_1724);
and U4853 (N_4853,In_1472,In_1380);
nor U4854 (N_4854,In_1943,In_1635);
nand U4855 (N_4855,In_1328,In_90);
xnor U4856 (N_4856,In_1117,In_1394);
and U4857 (N_4857,In_97,In_714);
or U4858 (N_4858,In_310,In_1979);
or U4859 (N_4859,In_1584,In_1668);
xor U4860 (N_4860,In_331,In_1272);
or U4861 (N_4861,In_1060,In_333);
or U4862 (N_4862,In_271,In_1997);
nor U4863 (N_4863,In_1886,In_1138);
nor U4864 (N_4864,In_1191,In_732);
and U4865 (N_4865,In_247,In_1335);
and U4866 (N_4866,In_1662,In_1265);
and U4867 (N_4867,In_1971,In_432);
and U4868 (N_4868,In_488,In_1178);
or U4869 (N_4869,In_1080,In_1352);
or U4870 (N_4870,In_1891,In_1898);
or U4871 (N_4871,In_306,In_949);
xnor U4872 (N_4872,In_1270,In_9);
or U4873 (N_4873,In_334,In_1004);
and U4874 (N_4874,In_696,In_1124);
nor U4875 (N_4875,In_1091,In_1038);
and U4876 (N_4876,In_1512,In_905);
nand U4877 (N_4877,In_1427,In_22);
or U4878 (N_4878,In_1064,In_642);
nand U4879 (N_4879,In_141,In_1026);
or U4880 (N_4880,In_1301,In_469);
xnor U4881 (N_4881,In_535,In_764);
and U4882 (N_4882,In_470,In_1551);
and U4883 (N_4883,In_527,In_1070);
nand U4884 (N_4884,In_1433,In_501);
nor U4885 (N_4885,In_808,In_417);
nand U4886 (N_4886,In_185,In_1152);
xor U4887 (N_4887,In_1160,In_423);
or U4888 (N_4888,In_242,In_1741);
xnor U4889 (N_4889,In_904,In_670);
nand U4890 (N_4890,In_1421,In_12);
nor U4891 (N_4891,In_247,In_515);
nand U4892 (N_4892,In_298,In_1646);
xnor U4893 (N_4893,In_38,In_35);
nand U4894 (N_4894,In_229,In_1654);
nor U4895 (N_4895,In_375,In_1978);
nor U4896 (N_4896,In_859,In_1633);
and U4897 (N_4897,In_624,In_1630);
nand U4898 (N_4898,In_580,In_1432);
nand U4899 (N_4899,In_146,In_907);
xnor U4900 (N_4900,In_459,In_288);
or U4901 (N_4901,In_905,In_1468);
nor U4902 (N_4902,In_518,In_1468);
nor U4903 (N_4903,In_1805,In_678);
nand U4904 (N_4904,In_1566,In_1288);
nand U4905 (N_4905,In_29,In_725);
nand U4906 (N_4906,In_1307,In_1014);
nor U4907 (N_4907,In_804,In_315);
nand U4908 (N_4908,In_1687,In_1125);
nor U4909 (N_4909,In_343,In_1004);
nor U4910 (N_4910,In_845,In_1932);
or U4911 (N_4911,In_1252,In_1944);
or U4912 (N_4912,In_375,In_685);
xnor U4913 (N_4913,In_836,In_1883);
or U4914 (N_4914,In_1664,In_1611);
and U4915 (N_4915,In_341,In_512);
and U4916 (N_4916,In_1907,In_772);
nor U4917 (N_4917,In_1094,In_997);
or U4918 (N_4918,In_726,In_145);
xnor U4919 (N_4919,In_853,In_406);
nor U4920 (N_4920,In_692,In_378);
and U4921 (N_4921,In_579,In_1506);
or U4922 (N_4922,In_125,In_57);
nor U4923 (N_4923,In_180,In_241);
xnor U4924 (N_4924,In_206,In_1376);
or U4925 (N_4925,In_1047,In_136);
or U4926 (N_4926,In_652,In_60);
nor U4927 (N_4927,In_699,In_578);
and U4928 (N_4928,In_954,In_1393);
or U4929 (N_4929,In_1308,In_314);
xor U4930 (N_4930,In_1515,In_873);
and U4931 (N_4931,In_503,In_1382);
xor U4932 (N_4932,In_792,In_1216);
xor U4933 (N_4933,In_1287,In_403);
or U4934 (N_4934,In_1331,In_1963);
and U4935 (N_4935,In_1764,In_1144);
nand U4936 (N_4936,In_274,In_1018);
nor U4937 (N_4937,In_1513,In_102);
xor U4938 (N_4938,In_404,In_1853);
or U4939 (N_4939,In_959,In_986);
nor U4940 (N_4940,In_1661,In_635);
or U4941 (N_4941,In_663,In_1962);
or U4942 (N_4942,In_763,In_982);
nand U4943 (N_4943,In_1489,In_279);
and U4944 (N_4944,In_1581,In_140);
and U4945 (N_4945,In_959,In_480);
nor U4946 (N_4946,In_1008,In_309);
nor U4947 (N_4947,In_1408,In_1367);
nor U4948 (N_4948,In_360,In_847);
nand U4949 (N_4949,In_1628,In_40);
nor U4950 (N_4950,In_101,In_1613);
or U4951 (N_4951,In_454,In_1701);
nand U4952 (N_4952,In_356,In_343);
or U4953 (N_4953,In_392,In_956);
or U4954 (N_4954,In_1207,In_30);
and U4955 (N_4955,In_1559,In_1243);
nor U4956 (N_4956,In_1442,In_1982);
nor U4957 (N_4957,In_672,In_1255);
and U4958 (N_4958,In_434,In_558);
nor U4959 (N_4959,In_1057,In_846);
and U4960 (N_4960,In_896,In_1058);
and U4961 (N_4961,In_1301,In_775);
and U4962 (N_4962,In_564,In_1426);
xnor U4963 (N_4963,In_1846,In_1362);
xnor U4964 (N_4964,In_307,In_1928);
nand U4965 (N_4965,In_427,In_398);
xor U4966 (N_4966,In_361,In_540);
nor U4967 (N_4967,In_1723,In_683);
nor U4968 (N_4968,In_265,In_47);
nor U4969 (N_4969,In_1424,In_1599);
nor U4970 (N_4970,In_1583,In_769);
or U4971 (N_4971,In_44,In_749);
xor U4972 (N_4972,In_847,In_181);
xnor U4973 (N_4973,In_380,In_1307);
nand U4974 (N_4974,In_224,In_1562);
and U4975 (N_4975,In_889,In_914);
and U4976 (N_4976,In_1588,In_762);
xor U4977 (N_4977,In_670,In_1393);
or U4978 (N_4978,In_265,In_1079);
and U4979 (N_4979,In_99,In_373);
nand U4980 (N_4980,In_1652,In_1077);
xor U4981 (N_4981,In_604,In_123);
or U4982 (N_4982,In_1978,In_97);
and U4983 (N_4983,In_1776,In_118);
and U4984 (N_4984,In_1239,In_1200);
nor U4985 (N_4985,In_486,In_495);
xnor U4986 (N_4986,In_160,In_283);
nor U4987 (N_4987,In_1466,In_1489);
nand U4988 (N_4988,In_1340,In_311);
nand U4989 (N_4989,In_1463,In_1400);
xnor U4990 (N_4990,In_1702,In_1744);
nor U4991 (N_4991,In_209,In_269);
or U4992 (N_4992,In_628,In_1327);
and U4993 (N_4993,In_302,In_538);
xor U4994 (N_4994,In_1151,In_285);
nand U4995 (N_4995,In_360,In_854);
and U4996 (N_4996,In_503,In_1756);
and U4997 (N_4997,In_1842,In_1582);
and U4998 (N_4998,In_1364,In_421);
and U4999 (N_4999,In_1958,In_403);
and U5000 (N_5000,N_2379,N_3226);
or U5001 (N_5001,N_1460,N_3286);
and U5002 (N_5002,N_1874,N_1248);
or U5003 (N_5003,N_25,N_1892);
or U5004 (N_5004,N_965,N_2137);
xnor U5005 (N_5005,N_3296,N_3657);
nand U5006 (N_5006,N_120,N_3891);
xor U5007 (N_5007,N_4099,N_4833);
and U5008 (N_5008,N_542,N_521);
nand U5009 (N_5009,N_969,N_4827);
and U5010 (N_5010,N_3275,N_2670);
xor U5011 (N_5011,N_1616,N_391);
and U5012 (N_5012,N_4314,N_3335);
xnor U5013 (N_5013,N_1280,N_2496);
xor U5014 (N_5014,N_1314,N_3260);
and U5015 (N_5015,N_3503,N_1072);
nor U5016 (N_5016,N_3633,N_1338);
nor U5017 (N_5017,N_4257,N_3549);
xor U5018 (N_5018,N_4641,N_1962);
nand U5019 (N_5019,N_2764,N_4916);
or U5020 (N_5020,N_2781,N_4326);
nand U5021 (N_5021,N_2629,N_456);
or U5022 (N_5022,N_3636,N_2297);
xor U5023 (N_5023,N_4535,N_180);
nor U5024 (N_5024,N_4419,N_4788);
and U5025 (N_5025,N_1080,N_2085);
nor U5026 (N_5026,N_4799,N_400);
nand U5027 (N_5027,N_1190,N_3515);
xnor U5028 (N_5028,N_3300,N_1744);
nand U5029 (N_5029,N_1995,N_892);
and U5030 (N_5030,N_914,N_1233);
xor U5031 (N_5031,N_1556,N_2836);
or U5032 (N_5032,N_4136,N_4014);
nand U5033 (N_5033,N_3783,N_4117);
nand U5034 (N_5034,N_3931,N_1804);
or U5035 (N_5035,N_1160,N_2959);
or U5036 (N_5036,N_3736,N_3211);
xor U5037 (N_5037,N_1590,N_2437);
nor U5038 (N_5038,N_4220,N_4829);
xnor U5039 (N_5039,N_3488,N_440);
nor U5040 (N_5040,N_1014,N_28);
or U5041 (N_5041,N_2156,N_4696);
nor U5042 (N_5042,N_2061,N_3537);
or U5043 (N_5043,N_3060,N_382);
or U5044 (N_5044,N_1776,N_2325);
or U5045 (N_5045,N_436,N_4366);
or U5046 (N_5046,N_48,N_3778);
nand U5047 (N_5047,N_4906,N_1917);
nand U5048 (N_5048,N_4560,N_2722);
and U5049 (N_5049,N_4589,N_1857);
nor U5050 (N_5050,N_3903,N_1216);
nor U5051 (N_5051,N_3767,N_3444);
nor U5052 (N_5052,N_477,N_1468);
xnor U5053 (N_5053,N_4893,N_1279);
nand U5054 (N_5054,N_4819,N_1195);
or U5055 (N_5055,N_2433,N_4236);
or U5056 (N_5056,N_747,N_3340);
and U5057 (N_5057,N_366,N_3996);
or U5058 (N_5058,N_2253,N_1512);
or U5059 (N_5059,N_1258,N_4736);
nand U5060 (N_5060,N_2912,N_4785);
or U5061 (N_5061,N_2470,N_666);
and U5062 (N_5062,N_3617,N_4392);
or U5063 (N_5063,N_2802,N_870);
xor U5064 (N_5064,N_1900,N_3268);
and U5065 (N_5065,N_4017,N_1820);
xor U5066 (N_5066,N_4184,N_4395);
and U5067 (N_5067,N_1440,N_4700);
nand U5068 (N_5068,N_1656,N_514);
or U5069 (N_5069,N_72,N_1806);
xor U5070 (N_5070,N_2858,N_3811);
xor U5071 (N_5071,N_2189,N_4515);
nand U5072 (N_5072,N_4120,N_93);
and U5073 (N_5073,N_2949,N_3535);
nand U5074 (N_5074,N_1403,N_523);
nor U5075 (N_5075,N_81,N_1681);
nand U5076 (N_5076,N_3435,N_3545);
or U5077 (N_5077,N_3789,N_579);
nand U5078 (N_5078,N_2247,N_3177);
nor U5079 (N_5079,N_2821,N_460);
and U5080 (N_5080,N_1538,N_3803);
nand U5081 (N_5081,N_2035,N_3153);
and U5082 (N_5082,N_2195,N_4559);
nor U5083 (N_5083,N_3396,N_2312);
xor U5084 (N_5084,N_1424,N_3733);
and U5085 (N_5085,N_322,N_1124);
nor U5086 (N_5086,N_794,N_4600);
or U5087 (N_5087,N_2684,N_3639);
nand U5088 (N_5088,N_2720,N_3283);
nor U5089 (N_5089,N_1557,N_4263);
xnor U5090 (N_5090,N_2546,N_4424);
and U5091 (N_5091,N_3566,N_264);
nor U5092 (N_5092,N_2425,N_3320);
and U5093 (N_5093,N_3788,N_479);
xor U5094 (N_5094,N_1396,N_3460);
and U5095 (N_5095,N_3748,N_4754);
nor U5096 (N_5096,N_3229,N_3579);
or U5097 (N_5097,N_800,N_4606);
nor U5098 (N_5098,N_2105,N_2032);
nand U5099 (N_5099,N_3687,N_4382);
and U5100 (N_5100,N_511,N_118);
and U5101 (N_5101,N_2748,N_3560);
or U5102 (N_5102,N_3380,N_4423);
or U5103 (N_5103,N_2547,N_3563);
nor U5104 (N_5104,N_3495,N_3347);
nand U5105 (N_5105,N_1311,N_2905);
and U5106 (N_5106,N_749,N_504);
or U5107 (N_5107,N_3117,N_1691);
xnor U5108 (N_5108,N_3987,N_2552);
or U5109 (N_5109,N_4988,N_4210);
or U5110 (N_5110,N_2669,N_2401);
and U5111 (N_5111,N_2309,N_2889);
and U5112 (N_5112,N_2106,N_503);
and U5113 (N_5113,N_1435,N_3136);
xor U5114 (N_5114,N_3955,N_3288);
and U5115 (N_5115,N_4155,N_549);
or U5116 (N_5116,N_3934,N_2757);
nand U5117 (N_5117,N_1352,N_291);
or U5118 (N_5118,N_110,N_3963);
nor U5119 (N_5119,N_4965,N_4302);
and U5120 (N_5120,N_1650,N_2682);
nor U5121 (N_5121,N_1020,N_1098);
and U5122 (N_5122,N_4996,N_4024);
and U5123 (N_5123,N_3466,N_4585);
and U5124 (N_5124,N_2279,N_4027);
or U5125 (N_5125,N_792,N_1096);
and U5126 (N_5126,N_774,N_3302);
and U5127 (N_5127,N_709,N_2770);
nand U5128 (N_5128,N_750,N_2248);
or U5129 (N_5129,N_4753,N_4898);
xor U5130 (N_5130,N_3475,N_4088);
and U5131 (N_5131,N_1724,N_2639);
and U5132 (N_5132,N_4828,N_3050);
nand U5133 (N_5133,N_3632,N_3561);
or U5134 (N_5134,N_3386,N_3345);
nand U5135 (N_5135,N_3081,N_4957);
nand U5136 (N_5136,N_4948,N_1492);
nor U5137 (N_5137,N_114,N_1772);
or U5138 (N_5138,N_3543,N_128);
xor U5139 (N_5139,N_1012,N_1399);
and U5140 (N_5140,N_2302,N_4476);
and U5141 (N_5141,N_2488,N_4687);
nor U5142 (N_5142,N_1376,N_1182);
or U5143 (N_5143,N_4322,N_2625);
xor U5144 (N_5144,N_153,N_813);
and U5145 (N_5145,N_4640,N_1618);
nor U5146 (N_5146,N_4356,N_2579);
xor U5147 (N_5147,N_4531,N_1977);
and U5148 (N_5148,N_2469,N_4285);
nand U5149 (N_5149,N_4016,N_2915);
and U5150 (N_5150,N_222,N_3509);
and U5151 (N_5151,N_4746,N_2212);
nor U5152 (N_5152,N_2107,N_1447);
and U5153 (N_5153,N_1059,N_340);
xor U5154 (N_5154,N_199,N_746);
nand U5155 (N_5155,N_814,N_1620);
and U5156 (N_5156,N_4518,N_4271);
nor U5157 (N_5157,N_2218,N_2752);
or U5158 (N_5158,N_986,N_1277);
nand U5159 (N_5159,N_304,N_2603);
nand U5160 (N_5160,N_1763,N_2076);
or U5161 (N_5161,N_3672,N_4351);
or U5162 (N_5162,N_2719,N_2004);
xnor U5163 (N_5163,N_3763,N_1034);
nand U5164 (N_5164,N_3093,N_1676);
or U5165 (N_5165,N_4260,N_4547);
nor U5166 (N_5166,N_4976,N_2311);
or U5167 (N_5167,N_148,N_748);
xnor U5168 (N_5168,N_1646,N_2755);
and U5169 (N_5169,N_3354,N_4170);
nand U5170 (N_5170,N_2332,N_2323);
nand U5171 (N_5171,N_33,N_4660);
and U5172 (N_5172,N_4508,N_1095);
and U5173 (N_5173,N_1973,N_2987);
nor U5174 (N_5174,N_4764,N_2376);
nand U5175 (N_5175,N_4722,N_589);
xor U5176 (N_5176,N_1450,N_3508);
nor U5177 (N_5177,N_14,N_879);
or U5178 (N_5178,N_3562,N_1601);
nor U5179 (N_5179,N_899,N_4288);
xnor U5180 (N_5180,N_4379,N_1050);
xor U5181 (N_5181,N_2850,N_1120);
and U5182 (N_5182,N_2732,N_1048);
or U5183 (N_5183,N_1436,N_2175);
and U5184 (N_5184,N_189,N_374);
or U5185 (N_5185,N_2344,N_3336);
or U5186 (N_5186,N_3063,N_192);
or U5187 (N_5187,N_1079,N_4448);
or U5188 (N_5188,N_334,N_1149);
or U5189 (N_5189,N_1934,N_3362);
or U5190 (N_5190,N_2319,N_1322);
nand U5191 (N_5191,N_1923,N_4738);
or U5192 (N_5192,N_2204,N_4406);
and U5193 (N_5193,N_3200,N_1673);
nand U5194 (N_5194,N_587,N_2466);
or U5195 (N_5195,N_4704,N_3127);
xnor U5196 (N_5196,N_1654,N_4383);
or U5197 (N_5197,N_2266,N_1877);
nor U5198 (N_5198,N_2733,N_2068);
and U5199 (N_5199,N_4331,N_1209);
xnor U5200 (N_5200,N_3062,N_2951);
or U5201 (N_5201,N_3254,N_386);
and U5202 (N_5202,N_4609,N_163);
and U5203 (N_5203,N_2818,N_1637);
xor U5204 (N_5204,N_3355,N_2996);
nand U5205 (N_5205,N_2555,N_1334);
and U5206 (N_5206,N_2386,N_1888);
nor U5207 (N_5207,N_4457,N_2591);
and U5208 (N_5208,N_4525,N_2994);
nand U5209 (N_5209,N_3526,N_2898);
and U5210 (N_5210,N_586,N_1915);
and U5211 (N_5211,N_2119,N_3680);
nand U5212 (N_5212,N_3592,N_2589);
or U5213 (N_5213,N_1873,N_946);
nand U5214 (N_5214,N_3197,N_4035);
or U5215 (N_5215,N_1169,N_2853);
xor U5216 (N_5216,N_1064,N_3252);
nor U5217 (N_5217,N_936,N_1348);
xnor U5218 (N_5218,N_2354,N_2141);
and U5219 (N_5219,N_2007,N_1087);
nand U5220 (N_5220,N_3860,N_4173);
or U5221 (N_5221,N_286,N_4144);
or U5222 (N_5222,N_2054,N_1342);
or U5223 (N_5223,N_3168,N_562);
nor U5224 (N_5224,N_883,N_3970);
nor U5225 (N_5225,N_3284,N_2094);
or U5226 (N_5226,N_232,N_4388);
nand U5227 (N_5227,N_1069,N_381);
and U5228 (N_5228,N_4370,N_780);
xnor U5229 (N_5229,N_1743,N_990);
and U5230 (N_5230,N_1379,N_2772);
nand U5231 (N_5231,N_4223,N_3704);
xnor U5232 (N_5232,N_1102,N_3096);
nand U5233 (N_5233,N_3149,N_3879);
xnor U5234 (N_5234,N_2811,N_851);
or U5235 (N_5235,N_2228,N_2863);
xor U5236 (N_5236,N_3175,N_301);
nor U5237 (N_5237,N_2055,N_882);
xor U5238 (N_5238,N_1949,N_1307);
xor U5239 (N_5239,N_2396,N_658);
or U5240 (N_5240,N_842,N_2717);
or U5241 (N_5241,N_2161,N_1373);
and U5242 (N_5242,N_4172,N_4509);
xnor U5243 (N_5243,N_3641,N_3843);
nand U5244 (N_5244,N_4488,N_3519);
or U5245 (N_5245,N_445,N_4338);
nand U5246 (N_5246,N_4368,N_2262);
xnor U5247 (N_5247,N_4743,N_2940);
and U5248 (N_5248,N_2724,N_2436);
and U5249 (N_5249,N_3462,N_1648);
and U5250 (N_5250,N_1276,N_463);
or U5251 (N_5251,N_2118,N_3115);
or U5252 (N_5252,N_1000,N_1525);
nand U5253 (N_5253,N_464,N_170);
xor U5254 (N_5254,N_1391,N_1769);
xnor U5255 (N_5255,N_3206,N_3741);
xnor U5256 (N_5256,N_3679,N_531);
nor U5257 (N_5257,N_3458,N_3204);
nand U5258 (N_5258,N_4817,N_3323);
and U5259 (N_5259,N_1895,N_1813);
nor U5260 (N_5260,N_4041,N_804);
nor U5261 (N_5261,N_2519,N_890);
xor U5262 (N_5262,N_3699,N_1253);
xnor U5263 (N_5263,N_1153,N_3586);
nand U5264 (N_5264,N_2807,N_2533);
and U5265 (N_5265,N_10,N_619);
and U5266 (N_5266,N_4871,N_4689);
xnor U5267 (N_5267,N_3010,N_1051);
xor U5268 (N_5268,N_2340,N_341);
or U5269 (N_5269,N_2271,N_1572);
and U5270 (N_5270,N_3048,N_2730);
xnor U5271 (N_5271,N_938,N_2986);
and U5272 (N_5272,N_1210,N_2593);
nor U5273 (N_5273,N_1380,N_3321);
nor U5274 (N_5274,N_4294,N_635);
nor U5275 (N_5275,N_519,N_2924);
nand U5276 (N_5276,N_98,N_3399);
and U5277 (N_5277,N_297,N_2147);
and U5278 (N_5278,N_3027,N_3674);
nor U5279 (N_5279,N_4066,N_785);
nor U5280 (N_5280,N_4514,N_730);
nor U5281 (N_5281,N_2485,N_644);
nand U5282 (N_5282,N_4800,N_2024);
and U5283 (N_5283,N_3079,N_3933);
or U5284 (N_5284,N_1966,N_3766);
xnor U5285 (N_5285,N_1581,N_3465);
nor U5286 (N_5286,N_3293,N_3802);
or U5287 (N_5287,N_2272,N_2193);
and U5288 (N_5288,N_2171,N_2217);
nor U5289 (N_5289,N_1996,N_2345);
xnor U5290 (N_5290,N_2492,N_3607);
nor U5291 (N_5291,N_1768,N_1818);
or U5292 (N_5292,N_2245,N_2065);
nand U5293 (N_5293,N_3266,N_3518);
xor U5294 (N_5294,N_843,N_3496);
xnor U5295 (N_5295,N_3927,N_845);
xnor U5296 (N_5296,N_91,N_2442);
xor U5297 (N_5297,N_4007,N_1497);
or U5298 (N_5298,N_1249,N_2962);
or U5299 (N_5299,N_4771,N_1580);
and U5300 (N_5300,N_4458,N_1699);
nand U5301 (N_5301,N_4078,N_4082);
nand U5302 (N_5302,N_1453,N_1786);
nor U5303 (N_5303,N_1615,N_3107);
and U5304 (N_5304,N_411,N_471);
nand U5305 (N_5305,N_97,N_4029);
nand U5306 (N_5306,N_1163,N_3898);
xnor U5307 (N_5307,N_1871,N_1922);
nor U5308 (N_5308,N_1863,N_3764);
or U5309 (N_5309,N_691,N_2185);
nor U5310 (N_5310,N_3279,N_1562);
nand U5311 (N_5311,N_1055,N_2698);
and U5312 (N_5312,N_3734,N_2);
and U5313 (N_5313,N_3270,N_4634);
xnor U5314 (N_5314,N_2444,N_1952);
or U5315 (N_5315,N_3393,N_639);
nor U5316 (N_5316,N_3609,N_3038);
or U5317 (N_5317,N_4346,N_3546);
or U5318 (N_5318,N_4287,N_1803);
nand U5319 (N_5319,N_1008,N_3326);
and U5320 (N_5320,N_3624,N_1510);
xor U5321 (N_5321,N_3012,N_1033);
and U5322 (N_5322,N_2851,N_2683);
xor U5323 (N_5323,N_1552,N_4079);
and U5324 (N_5324,N_442,N_3572);
nand U5325 (N_5325,N_345,N_3423);
nor U5326 (N_5326,N_3962,N_540);
or U5327 (N_5327,N_4101,N_3779);
or U5328 (N_5328,N_169,N_4703);
nand U5329 (N_5329,N_4218,N_3652);
and U5330 (N_5330,N_4032,N_3431);
xnor U5331 (N_5331,N_3352,N_3249);
xor U5332 (N_5332,N_4189,N_3398);
nand U5333 (N_5333,N_904,N_3377);
nor U5334 (N_5334,N_4554,N_1545);
or U5335 (N_5335,N_2315,N_1729);
and U5336 (N_5336,N_2398,N_1198);
nand U5337 (N_5337,N_1047,N_4021);
nand U5338 (N_5338,N_2829,N_4723);
nand U5339 (N_5339,N_1765,N_795);
and U5340 (N_5340,N_3432,N_4915);
nor U5341 (N_5341,N_3816,N_1641);
nor U5342 (N_5342,N_3900,N_3565);
and U5343 (N_5343,N_4334,N_3080);
nand U5344 (N_5344,N_4197,N_856);
xor U5345 (N_5345,N_3799,N_3813);
nand U5346 (N_5346,N_4921,N_3282);
or U5347 (N_5347,N_2461,N_1106);
and U5348 (N_5348,N_4434,N_3961);
nor U5349 (N_5349,N_3071,N_887);
nand U5350 (N_5350,N_2567,N_2139);
and U5351 (N_5351,N_4286,N_4697);
nor U5352 (N_5352,N_3676,N_4216);
and U5353 (N_5353,N_1548,N_2935);
and U5354 (N_5354,N_3188,N_2009);
and U5355 (N_5355,N_4654,N_4283);
or U5356 (N_5356,N_307,N_623);
nor U5357 (N_5357,N_3649,N_2739);
and U5358 (N_5358,N_538,N_4137);
nand U5359 (N_5359,N_1173,N_1009);
or U5360 (N_5360,N_4802,N_4883);
nor U5361 (N_5361,N_4923,N_3928);
and U5362 (N_5362,N_4087,N_615);
nor U5363 (N_5363,N_557,N_4427);
and U5364 (N_5364,N_4147,N_3866);
or U5365 (N_5365,N_3400,N_2120);
and U5366 (N_5366,N_4768,N_4524);
xor U5367 (N_5367,N_1706,N_3276);
xnor U5368 (N_5368,N_4450,N_1415);
nand U5369 (N_5369,N_117,N_3945);
xnor U5370 (N_5370,N_1591,N_3628);
nor U5371 (N_5371,N_2928,N_3512);
nand U5372 (N_5372,N_1986,N_1134);
or U5373 (N_5373,N_2943,N_182);
nor U5374 (N_5374,N_3610,N_337);
and U5375 (N_5375,N_1491,N_4623);
nor U5376 (N_5376,N_3539,N_2092);
or U5377 (N_5377,N_2746,N_2978);
xor U5378 (N_5378,N_3247,N_2524);
or U5379 (N_5379,N_2016,N_403);
nand U5380 (N_5380,N_4719,N_4683);
and U5381 (N_5381,N_4964,N_3787);
nand U5382 (N_5382,N_3479,N_1375);
or U5383 (N_5383,N_4157,N_2048);
nor U5384 (N_5384,N_292,N_3834);
and U5385 (N_5385,N_4232,N_3376);
and U5386 (N_5386,N_3494,N_1068);
nand U5387 (N_5387,N_3534,N_2144);
or U5388 (N_5388,N_2981,N_778);
nand U5389 (N_5389,N_2630,N_1371);
nand U5390 (N_5390,N_3710,N_1222);
and U5391 (N_5391,N_962,N_2244);
nand U5392 (N_5392,N_2516,N_4038);
or U5393 (N_5393,N_465,N_1550);
xnor U5394 (N_5394,N_1636,N_909);
xnor U5395 (N_5395,N_4487,N_3890);
xor U5396 (N_5396,N_4501,N_2693);
nand U5397 (N_5397,N_1519,N_2631);
xor U5398 (N_5398,N_4061,N_2690);
or U5399 (N_5399,N_2930,N_1695);
nand U5400 (N_5400,N_2718,N_683);
xor U5401 (N_5401,N_4397,N_3424);
nor U5402 (N_5402,N_1145,N_3749);
and U5403 (N_5403,N_4786,N_1758);
and U5404 (N_5404,N_2080,N_2356);
nor U5405 (N_5405,N_3611,N_4414);
xnor U5406 (N_5406,N_1549,N_4646);
nor U5407 (N_5407,N_1669,N_581);
nand U5408 (N_5408,N_1383,N_3068);
or U5409 (N_5409,N_4505,N_347);
xnor U5410 (N_5410,N_520,N_4954);
nor U5411 (N_5411,N_3404,N_484);
xor U5412 (N_5412,N_2481,N_41);
or U5413 (N_5413,N_1728,N_1031);
or U5414 (N_5414,N_1180,N_3058);
or U5415 (N_5415,N_434,N_410);
nand U5416 (N_5416,N_420,N_246);
xnor U5417 (N_5417,N_4244,N_283);
or U5418 (N_5418,N_2849,N_4238);
and U5419 (N_5419,N_2077,N_377);
nand U5420 (N_5420,N_3123,N_1869);
or U5421 (N_5421,N_1975,N_2153);
or U5422 (N_5422,N_1679,N_1740);
nand U5423 (N_5423,N_2478,N_2737);
nand U5424 (N_5424,N_437,N_3274);
nor U5425 (N_5425,N_409,N_1146);
nand U5426 (N_5426,N_744,N_1594);
nand U5427 (N_5427,N_3645,N_2167);
nand U5428 (N_5428,N_116,N_931);
xor U5429 (N_5429,N_2365,N_4549);
nor U5430 (N_5430,N_3194,N_3199);
nand U5431 (N_5431,N_578,N_2740);
nand U5432 (N_5432,N_1269,N_3057);
nor U5433 (N_5433,N_4064,N_1807);
or U5434 (N_5434,N_2942,N_3634);
xor U5435 (N_5435,N_4122,N_2441);
and U5436 (N_5436,N_1746,N_4649);
and U5437 (N_5437,N_2251,N_1866);
xnor U5438 (N_5438,N_4308,N_629);
nor U5439 (N_5439,N_4201,N_4469);
nor U5440 (N_5440,N_2238,N_1619);
and U5441 (N_5441,N_1236,N_2677);
nand U5442 (N_5442,N_4116,N_4046);
nand U5443 (N_5443,N_996,N_1386);
nor U5444 (N_5444,N_4112,N_2400);
nand U5445 (N_5445,N_601,N_90);
nor U5446 (N_5446,N_3725,N_862);
xor U5447 (N_5447,N_1896,N_3133);
or U5448 (N_5448,N_3869,N_4729);
nand U5449 (N_5449,N_1870,N_4164);
and U5450 (N_5450,N_2665,N_1238);
and U5451 (N_5451,N_1805,N_3339);
nor U5452 (N_5452,N_4720,N_2627);
xnor U5453 (N_5453,N_547,N_782);
or U5454 (N_5454,N_3456,N_3904);
or U5455 (N_5455,N_1286,N_4203);
and U5456 (N_5456,N_4854,N_4413);
nand U5457 (N_5457,N_1795,N_1239);
xnor U5458 (N_5458,N_3712,N_4999);
xnor U5459 (N_5459,N_1514,N_1762);
nand U5460 (N_5460,N_3908,N_1467);
xnor U5461 (N_5461,N_1644,N_1204);
or U5462 (N_5462,N_819,N_4199);
xnor U5463 (N_5463,N_4669,N_976);
and U5464 (N_5464,N_1285,N_4674);
xor U5465 (N_5465,N_496,N_4822);
xnor U5466 (N_5466,N_3831,N_1148);
nand U5467 (N_5467,N_3969,N_3420);
or U5468 (N_5468,N_2965,N_2176);
and U5469 (N_5469,N_1496,N_2574);
nand U5470 (N_5470,N_584,N_622);
xor U5471 (N_5471,N_852,N_2150);
or U5472 (N_5472,N_4482,N_3896);
xnor U5473 (N_5473,N_65,N_3245);
nand U5474 (N_5474,N_759,N_3443);
and U5475 (N_5475,N_4150,N_2155);
nand U5476 (N_5476,N_2929,N_1416);
and U5477 (N_5477,N_2227,N_530);
nor U5478 (N_5478,N_2003,N_330);
nor U5479 (N_5479,N_1540,N_1321);
and U5480 (N_5480,N_4275,N_103);
nand U5481 (N_5481,N_3008,N_3716);
or U5482 (N_5482,N_417,N_375);
nor U5483 (N_5483,N_1187,N_2636);
or U5484 (N_5484,N_392,N_3568);
and U5485 (N_5485,N_684,N_3433);
nor U5486 (N_5486,N_111,N_11);
or U5487 (N_5487,N_4242,N_1702);
nor U5488 (N_5488,N_2694,N_2310);
and U5489 (N_5489,N_4912,N_4569);
xor U5490 (N_5490,N_2439,N_2357);
nand U5491 (N_5491,N_4058,N_388);
nand U5492 (N_5492,N_3744,N_82);
nor U5493 (N_5493,N_2179,N_4337);
nor U5494 (N_5494,N_3,N_122);
nand U5495 (N_5495,N_4566,N_4750);
xor U5496 (N_5496,N_2729,N_803);
or U5497 (N_5497,N_3836,N_2371);
nor U5498 (N_5498,N_4068,N_157);
nand U5499 (N_5499,N_3997,N_929);
nand U5500 (N_5500,N_1796,N_4779);
nor U5501 (N_5501,N_2526,N_3406);
and U5502 (N_5502,N_78,N_1211);
and U5503 (N_5503,N_2038,N_2184);
nand U5504 (N_5504,N_2809,N_1651);
xor U5505 (N_5505,N_2070,N_3478);
xnor U5506 (N_5506,N_2369,N_3122);
nor U5507 (N_5507,N_4810,N_3812);
xnor U5508 (N_5508,N_1939,N_3576);
nor U5509 (N_5509,N_3793,N_4707);
nor U5510 (N_5510,N_4726,N_218);
or U5511 (N_5511,N_2261,N_3223);
xor U5512 (N_5512,N_3281,N_1404);
nor U5513 (N_5513,N_3210,N_1060);
nand U5514 (N_5514,N_4929,N_1183);
or U5515 (N_5515,N_4130,N_4090);
nor U5516 (N_5516,N_2662,N_1355);
xor U5517 (N_5517,N_265,N_947);
nor U5518 (N_5518,N_3654,N_1791);
and U5519 (N_5519,N_4798,N_1049);
nor U5520 (N_5520,N_1797,N_4666);
nor U5521 (N_5521,N_2078,N_993);
or U5522 (N_5522,N_4229,N_1684);
nor U5523 (N_5523,N_4299,N_4284);
or U5524 (N_5524,N_2545,N_4);
and U5525 (N_5525,N_4960,N_3824);
nand U5526 (N_5526,N_2170,N_543);
nor U5527 (N_5527,N_4962,N_2633);
xor U5528 (N_5528,N_2933,N_2890);
or U5529 (N_5529,N_3378,N_1584);
nand U5530 (N_5530,N_4652,N_1369);
and U5531 (N_5531,N_3312,N_3191);
xnor U5532 (N_5532,N_877,N_2919);
or U5533 (N_5533,N_1135,N_802);
or U5534 (N_5534,N_4598,N_1897);
and U5535 (N_5535,N_4303,N_2979);
and U5536 (N_5536,N_1612,N_3360);
and U5537 (N_5537,N_4715,N_4234);
and U5538 (N_5538,N_3762,N_119);
or U5539 (N_5539,N_3761,N_3946);
nand U5540 (N_5540,N_2765,N_475);
nor U5541 (N_5541,N_3309,N_290);
xor U5542 (N_5542,N_1954,N_1388);
or U5543 (N_5543,N_1988,N_494);
or U5544 (N_5544,N_1046,N_1174);
and U5545 (N_5545,N_1751,N_3440);
or U5546 (N_5546,N_1118,N_2964);
or U5547 (N_5547,N_2801,N_3520);
nand U5548 (N_5548,N_43,N_3089);
and U5549 (N_5549,N_3977,N_2455);
nor U5550 (N_5550,N_4769,N_3614);
and U5551 (N_5551,N_1189,N_4040);
or U5552 (N_5552,N_967,N_378);
nand U5553 (N_5553,N_317,N_419);
and U5554 (N_5554,N_3294,N_9);
xor U5555 (N_5555,N_1518,N_2337);
xor U5556 (N_5556,N_772,N_4572);
or U5557 (N_5557,N_1766,N_3132);
xnor U5558 (N_5558,N_3959,N_630);
xnor U5559 (N_5559,N_4995,N_3979);
nor U5560 (N_5560,N_4865,N_1030);
and U5561 (N_5561,N_742,N_1508);
nor U5562 (N_5562,N_2592,N_3161);
or U5563 (N_5563,N_2602,N_1945);
xnor U5564 (N_5564,N_3324,N_2957);
nand U5565 (N_5565,N_3669,N_701);
xnor U5566 (N_5566,N_3501,N_3740);
nand U5567 (N_5567,N_2329,N_1052);
xnor U5568 (N_5568,N_522,N_3041);
and U5569 (N_5569,N_4783,N_96);
nand U5570 (N_5570,N_2215,N_2913);
and U5571 (N_5571,N_3852,N_4429);
and U5572 (N_5572,N_2681,N_529);
or U5573 (N_5573,N_3411,N_2330);
and U5574 (N_5574,N_3061,N_3616);
xnor U5575 (N_5575,N_3837,N_806);
or U5576 (N_5576,N_3299,N_4421);
xnor U5577 (N_5577,N_3165,N_1465);
and U5578 (N_5578,N_606,N_4836);
nand U5579 (N_5579,N_1574,N_561);
nand U5580 (N_5580,N_4862,N_2234);
nor U5581 (N_5581,N_2278,N_4451);
and U5582 (N_5582,N_4168,N_4702);
and U5583 (N_5583,N_4952,N_3818);
or U5584 (N_5584,N_3434,N_3973);
nor U5585 (N_5585,N_2463,N_4968);
xnor U5586 (N_5586,N_2879,N_1504);
and U5587 (N_5587,N_4228,N_4327);
or U5588 (N_5588,N_1177,N_603);
or U5589 (N_5589,N_3148,N_3729);
and U5590 (N_5590,N_3702,N_4853);
or U5591 (N_5591,N_4857,N_761);
nor U5592 (N_5592,N_1607,N_389);
and U5593 (N_5593,N_1073,N_3113);
or U5594 (N_5594,N_4823,N_1745);
and U5595 (N_5595,N_512,N_508);
or U5596 (N_5596,N_1312,N_613);
nor U5597 (N_5597,N_469,N_4162);
nand U5598 (N_5598,N_608,N_160);
nand U5599 (N_5599,N_324,N_517);
nor U5600 (N_5600,N_3999,N_3544);
nand U5601 (N_5601,N_3248,N_3559);
and U5602 (N_5602,N_220,N_2842);
xnor U5603 (N_5603,N_3361,N_50);
nand U5604 (N_5604,N_835,N_1812);
and U5605 (N_5605,N_1576,N_313);
or U5606 (N_5606,N_2026,N_942);
and U5607 (N_5607,N_4766,N_2199);
or U5608 (N_5608,N_4156,N_4790);
nand U5609 (N_5609,N_3510,N_3912);
or U5610 (N_5610,N_4249,N_745);
and U5611 (N_5611,N_399,N_3310);
nand U5612 (N_5612,N_4489,N_4985);
xnor U5613 (N_5613,N_4807,N_1502);
or U5614 (N_5614,N_3451,N_211);
nor U5615 (N_5615,N_4742,N_4447);
xnor U5616 (N_5616,N_4716,N_1275);
and U5617 (N_5617,N_4477,N_2535);
or U5618 (N_5618,N_3730,N_4980);
xnor U5619 (N_5619,N_4553,N_3727);
nor U5620 (N_5620,N_2422,N_4565);
or U5621 (N_5621,N_3455,N_2250);
nor U5622 (N_5622,N_705,N_4591);
or U5623 (N_5623,N_2382,N_3626);
and U5624 (N_5624,N_672,N_3792);
and U5625 (N_5625,N_1726,N_136);
and U5626 (N_5626,N_4721,N_2623);
nor U5627 (N_5627,N_4042,N_2663);
xnor U5628 (N_5628,N_3615,N_1879);
or U5629 (N_5629,N_326,N_1251);
xor U5630 (N_5630,N_2892,N_686);
xnor U5631 (N_5631,N_4814,N_1981);
xor U5632 (N_5632,N_438,N_1592);
xor U5633 (N_5633,N_212,N_3950);
xnor U5634 (N_5634,N_4935,N_1319);
or U5635 (N_5635,N_2880,N_412);
nor U5636 (N_5636,N_766,N_3913);
xor U5637 (N_5637,N_1992,N_2900);
nand U5638 (N_5638,N_1625,N_1446);
nand U5639 (N_5639,N_826,N_2872);
and U5640 (N_5640,N_4272,N_2927);
nand U5641 (N_5641,N_4939,N_1527);
and U5642 (N_5642,N_3909,N_739);
xnor U5643 (N_5643,N_2571,N_3438);
or U5644 (N_5644,N_2109,N_2281);
nor U5645 (N_5645,N_1881,N_2213);
and U5646 (N_5646,N_1074,N_1214);
nor U5647 (N_5647,N_2826,N_4930);
and U5648 (N_5648,N_27,N_4376);
or U5649 (N_5649,N_4381,N_1696);
nor U5650 (N_5650,N_4387,N_3665);
and U5651 (N_5651,N_811,N_2468);
xnor U5652 (N_5652,N_2317,N_1315);
nand U5653 (N_5653,N_1710,N_4097);
xor U5654 (N_5654,N_1473,N_3746);
and U5655 (N_5655,N_61,N_483);
and U5656 (N_5656,N_4363,N_1);
or U5657 (N_5657,N_4604,N_2058);
or U5658 (N_5658,N_4324,N_4731);
or U5659 (N_5659,N_1774,N_2785);
nand U5660 (N_5660,N_1964,N_3745);
nor U5661 (N_5661,N_2936,N_4903);
nand U5662 (N_5662,N_1571,N_4163);
xnor U5663 (N_5663,N_2710,N_1741);
nand U5664 (N_5664,N_3753,N_2243);
or U5665 (N_5665,N_1292,N_3150);
nand U5666 (N_5666,N_676,N_2859);
and U5667 (N_5667,N_4552,N_3506);
xnor U5668 (N_5668,N_4842,N_1910);
nor U5669 (N_5669,N_4103,N_1536);
nor U5670 (N_5670,N_3826,N_2703);
and U5671 (N_5671,N_1221,N_2615);
xnor U5672 (N_5672,N_4362,N_791);
nand U5673 (N_5673,N_4770,N_1856);
nand U5674 (N_5674,N_2728,N_3608);
nor U5675 (N_5675,N_3118,N_3292);
or U5676 (N_5676,N_2619,N_1853);
and U5677 (N_5677,N_3646,N_202);
and U5678 (N_5678,N_1335,N_274);
nand U5679 (N_5679,N_241,N_2705);
or U5680 (N_5680,N_4310,N_2168);
xnor U5681 (N_5681,N_628,N_2128);
or U5682 (N_5682,N_2052,N_2438);
and U5683 (N_5683,N_1240,N_2559);
xor U5684 (N_5684,N_945,N_3228);
nor U5685 (N_5685,N_3937,N_2203);
and U5686 (N_5686,N_2887,N_4459);
nand U5687 (N_5687,N_2335,N_3956);
nand U5688 (N_5688,N_2449,N_263);
and U5689 (N_5689,N_754,N_2404);
and U5690 (N_5690,N_3042,N_3358);
nand U5691 (N_5691,N_2146,N_1894);
xor U5692 (N_5692,N_3577,N_4400);
or U5693 (N_5693,N_3667,N_3325);
nor U5694 (N_5694,N_3034,N_210);
or U5695 (N_5695,N_1200,N_335);
and U5696 (N_5696,N_911,N_4613);
nor U5697 (N_5697,N_4139,N_4013);
xor U5698 (N_5698,N_38,N_1953);
nor U5699 (N_5699,N_1674,N_446);
nor U5700 (N_5700,N_3169,N_3124);
nand U5701 (N_5701,N_2820,N_3907);
xor U5702 (N_5702,N_3151,N_269);
nand U5703 (N_5703,N_450,N_898);
or U5704 (N_5704,N_4767,N_991);
or U5705 (N_5705,N_2706,N_1529);
nor U5706 (N_5706,N_4364,N_4153);
nand U5707 (N_5707,N_2843,N_889);
or U5708 (N_5708,N_332,N_2419);
xnor U5709 (N_5709,N_509,N_567);
nand U5710 (N_5710,N_3500,N_2513);
nor U5711 (N_5711,N_626,N_4063);
and U5712 (N_5712,N_2225,N_1771);
and U5713 (N_5713,N_4837,N_2847);
or U5714 (N_5714,N_1463,N_3743);
or U5715 (N_5715,N_4936,N_2368);
xor U5716 (N_5716,N_956,N_3975);
nand U5717 (N_5717,N_1814,N_4404);
nand U5718 (N_5718,N_689,N_2808);
or U5719 (N_5719,N_4864,N_3986);
or U5720 (N_5720,N_855,N_4268);
xnor U5721 (N_5721,N_674,N_1043);
and U5722 (N_5722,N_3187,N_861);
nor U5723 (N_5723,N_2017,N_1076);
and U5724 (N_5724,N_2945,N_3137);
nor U5725 (N_5725,N_84,N_4787);
nand U5726 (N_5726,N_1722,N_3643);
and U5727 (N_5727,N_3297,N_1867);
or U5728 (N_5728,N_1501,N_3648);
nor U5729 (N_5729,N_4863,N_1105);
nand U5730 (N_5730,N_4737,N_4624);
nand U5731 (N_5731,N_2129,N_156);
or U5732 (N_5732,N_4192,N_4775);
and U5733 (N_5733,N_3967,N_3230);
xnor U5734 (N_5734,N_2828,N_2394);
xnor U5735 (N_5735,N_2590,N_3035);
nand U5736 (N_5736,N_1883,N_645);
and U5737 (N_5737,N_205,N_4293);
nor U5738 (N_5738,N_1622,N_2861);
xnor U5739 (N_5739,N_1513,N_3660);
or U5740 (N_5740,N_2968,N_837);
xor U5741 (N_5741,N_1841,N_3043);
or U5742 (N_5742,N_2283,N_2429);
nand U5743 (N_5743,N_1242,N_594);
nand U5744 (N_5744,N_1831,N_662);
xor U5745 (N_5745,N_4280,N_4152);
xnor U5746 (N_5746,N_67,N_1439);
nor U5747 (N_5747,N_656,N_2410);
xnor U5748 (N_5748,N_3938,N_4874);
and U5749 (N_5749,N_1166,N_4597);
or U5750 (N_5750,N_526,N_2108);
or U5751 (N_5751,N_1787,N_2066);
and U5752 (N_5752,N_3120,N_255);
or U5753 (N_5753,N_2654,N_3939);
nand U5754 (N_5754,N_944,N_1101);
and U5755 (N_5755,N_499,N_3445);
nand U5756 (N_5756,N_498,N_755);
nand U5757 (N_5757,N_2164,N_4852);
nor U5758 (N_5758,N_2423,N_2166);
or U5759 (N_5759,N_1868,N_2715);
nor U5760 (N_5760,N_849,N_2268);
or U5761 (N_5761,N_354,N_3715);
or U5762 (N_5762,N_83,N_2896);
nor U5763 (N_5763,N_805,N_2503);
nand U5764 (N_5764,N_3265,N_1125);
xor U5765 (N_5765,N_2643,N_3739);
and U5766 (N_5766,N_597,N_3231);
or U5767 (N_5767,N_1357,N_1932);
and U5768 (N_5768,N_3430,N_1734);
or U5769 (N_5769,N_1756,N_2561);
nand U5770 (N_5770,N_1567,N_2350);
and U5771 (N_5771,N_1539,N_654);
and U5772 (N_5772,N_384,N_4258);
nor U5773 (N_5773,N_4071,N_4091);
or U5774 (N_5774,N_4276,N_367);
nor U5775 (N_5775,N_4676,N_3873);
and U5776 (N_5776,N_1389,N_858);
xor U5777 (N_5777,N_3517,N_1793);
and U5778 (N_5778,N_3718,N_3521);
nor U5779 (N_5779,N_1230,N_4384);
or U5780 (N_5780,N_4815,N_1639);
nor U5781 (N_5781,N_2641,N_532);
or U5782 (N_5782,N_2673,N_233);
nand U5783 (N_5783,N_1485,N_124);
xnor U5784 (N_5784,N_2445,N_4592);
nand U5785 (N_5785,N_428,N_1162);
nor U5786 (N_5786,N_4067,N_4507);
nand U5787 (N_5787,N_866,N_2486);
nor U5788 (N_5788,N_3542,N_312);
nand U5789 (N_5789,N_46,N_2505);
nor U5790 (N_5790,N_2906,N_978);
or U5791 (N_5791,N_1299,N_3403);
xor U5792 (N_5792,N_3178,N_700);
and U5793 (N_5793,N_3516,N_4650);
nor U5794 (N_5794,N_308,N_2308);
or U5795 (N_5795,N_2125,N_3548);
or U5796 (N_5796,N_492,N_187);
or U5797 (N_5797,N_196,N_3083);
nand U5798 (N_5798,N_323,N_544);
or U5799 (N_5799,N_2680,N_4845);
nand U5800 (N_5800,N_2992,N_4497);
or U5801 (N_5801,N_651,N_3601);
nand U5802 (N_5802,N_1717,N_1495);
nor U5803 (N_5803,N_2908,N_430);
xor U5804 (N_5804,N_1126,N_3287);
nor U5805 (N_5805,N_271,N_294);
nor U5806 (N_5806,N_1547,N_1689);
or U5807 (N_5807,N_2214,N_1579);
or U5808 (N_5808,N_4213,N_2282);
nor U5809 (N_5809,N_770,N_4587);
xnor U5810 (N_5810,N_2659,N_448);
nor U5811 (N_5811,N_3209,N_1950);
and U5812 (N_5812,N_1506,N_2824);
nor U5813 (N_5813,N_1889,N_1003);
and U5814 (N_5814,N_2183,N_1919);
nor U5815 (N_5815,N_1021,N_4107);
nor U5816 (N_5816,N_2464,N_1642);
nand U5817 (N_5817,N_3181,N_3876);
xor U5818 (N_5818,N_4300,N_1372);
nand U5819 (N_5819,N_1621,N_1767);
nand U5820 (N_5820,N_175,N_1032);
and U5821 (N_5821,N_3830,N_2657);
nor U5822 (N_5822,N_2576,N_4686);
or U5823 (N_5823,N_2355,N_237);
xnor U5824 (N_5824,N_1731,N_2408);
nor U5825 (N_5825,N_810,N_3606);
nor U5826 (N_5826,N_179,N_4655);
xor U5827 (N_5827,N_2976,N_1585);
or U5828 (N_5828,N_1693,N_3246);
xnor U5829 (N_5829,N_4776,N_556);
and U5830 (N_5830,N_569,N_3864);
nor U5831 (N_5831,N_3272,N_3694);
xnor U5832 (N_5832,N_1212,N_4596);
xnor U5833 (N_5833,N_4006,N_4306);
and U5834 (N_5834,N_1980,N_1711);
or U5835 (N_5835,N_4782,N_3306);
nand U5836 (N_5836,N_3155,N_3951);
and U5837 (N_5837,N_3032,N_2426);
nand U5838 (N_5838,N_395,N_2381);
xor U5839 (N_5839,N_2377,N_2769);
nand U5840 (N_5840,N_3708,N_1564);
or U5841 (N_5841,N_80,N_4291);
xnor U5842 (N_5842,N_4019,N_4727);
and U5843 (N_5843,N_3737,N_66);
xor U5844 (N_5844,N_3037,N_4437);
nand U5845 (N_5845,N_4323,N_2046);
or U5846 (N_5846,N_2257,N_1246);
nand U5847 (N_5847,N_3110,N_3116);
or U5848 (N_5848,N_2235,N_661);
or U5849 (N_5849,N_2926,N_4896);
xnor U5850 (N_5850,N_3439,N_200);
nand U5851 (N_5851,N_4274,N_4733);
xnor U5852 (N_5852,N_45,N_4281);
nor U5853 (N_5853,N_528,N_1354);
xor U5854 (N_5854,N_4160,N_1176);
nand U5855 (N_5855,N_1738,N_2766);
nand U5856 (N_5856,N_3220,N_2029);
and U5857 (N_5857,N_4973,N_4359);
nor U5858 (N_5858,N_3541,N_872);
xor U5859 (N_5859,N_4125,N_4399);
xor U5860 (N_5860,N_359,N_2294);
xor U5861 (N_5861,N_4262,N_2787);
nand U5862 (N_5862,N_2595,N_4876);
or U5863 (N_5863,N_2044,N_3142);
and U5864 (N_5864,N_2884,N_3205);
nor U5865 (N_5865,N_534,N_3207);
xnor U5866 (N_5866,N_4678,N_58);
or U5867 (N_5867,N_1438,N_507);
nor U5868 (N_5868,N_4927,N_536);
nor U5869 (N_5869,N_4377,N_3487);
nor U5870 (N_5870,N_3459,N_2130);
or U5871 (N_5871,N_2521,N_1344);
nor U5872 (N_5872,N_1154,N_421);
nand U5873 (N_5873,N_3700,N_1083);
or U5874 (N_5874,N_1847,N_4290);
nor U5875 (N_5875,N_3045,N_2789);
nand U5876 (N_5876,N_568,N_1172);
xor U5877 (N_5877,N_3828,N_2606);
xor U5878 (N_5878,N_3463,N_4086);
nand U5879 (N_5879,N_168,N_4060);
nand U5880 (N_5880,N_70,N_596);
or U5881 (N_5881,N_1703,N_847);
nor U5882 (N_5882,N_1957,N_4023);
or U5883 (N_5883,N_1281,N_3504);
and U5884 (N_5884,N_1516,N_4994);
nor U5885 (N_5885,N_4221,N_4297);
or U5886 (N_5886,N_4914,N_4897);
nor U5887 (N_5887,N_231,N_2483);
nand U5888 (N_5888,N_3681,N_1822);
nor U5889 (N_5889,N_1810,N_671);
nor U5890 (N_5890,N_3768,N_681);
or U5891 (N_5891,N_2512,N_4418);
xnor U5892 (N_5892,N_4253,N_1901);
or U5893 (N_5893,N_958,N_2726);
nand U5894 (N_5894,N_2901,N_3750);
and U5895 (N_5895,N_2661,N_3261);
or U5896 (N_5896,N_444,N_2020);
and U5897 (N_5897,N_3388,N_1596);
nand U5898 (N_5898,N_1927,N_1066);
nand U5899 (N_5899,N_3942,N_1918);
or U5900 (N_5900,N_2971,N_1413);
nand U5901 (N_5901,N_3002,N_287);
nand U5902 (N_5902,N_3815,N_183);
nor U5903 (N_5903,N_257,N_3499);
and U5904 (N_5904,N_225,N_2554);
nor U5905 (N_5905,N_1569,N_753);
and U5906 (N_5906,N_4403,N_921);
and U5907 (N_5907,N_1359,N_2773);
or U5908 (N_5908,N_2779,N_559);
nand U5909 (N_5909,N_3344,N_4576);
or U5910 (N_5910,N_2321,N_361);
xnor U5911 (N_5911,N_2079,N_3469);
nand U5912 (N_5912,N_4454,N_2451);
and U5913 (N_5913,N_2753,N_2136);
and U5914 (N_5914,N_4811,N_406);
xor U5915 (N_5915,N_145,N_4398);
xor U5916 (N_5916,N_1511,N_3391);
xor U5917 (N_5917,N_951,N_1997);
or U5918 (N_5918,N_524,N_2346);
nor U5919 (N_5919,N_3854,N_1882);
and U5920 (N_5920,N_217,N_3221);
nor U5921 (N_5921,N_1400,N_2938);
xnor U5922 (N_5922,N_2497,N_533);
nor U5923 (N_5923,N_1428,N_2490);
nor U5924 (N_5924,N_1001,N_2053);
and U5925 (N_5925,N_2001,N_998);
xnor U5926 (N_5926,N_2974,N_3806);
and U5927 (N_5927,N_3253,N_3203);
nor U5928 (N_5928,N_3732,N_833);
and U5929 (N_5929,N_123,N_478);
xnor U5930 (N_5930,N_4127,N_4922);
xnor U5931 (N_5931,N_3492,N_4892);
or U5932 (N_5932,N_4296,N_1156);
nor U5933 (N_5933,N_2612,N_4673);
nand U5934 (N_5934,N_4026,N_3551);
nor U5935 (N_5935,N_1994,N_850);
and U5936 (N_5936,N_3557,N_633);
nand U5937 (N_5937,N_3735,N_338);
nor U5938 (N_5938,N_4261,N_1799);
or U5939 (N_5939,N_3794,N_3104);
xor U5940 (N_5940,N_4452,N_2034);
xor U5941 (N_5941,N_1666,N_4273);
and U5942 (N_5942,N_47,N_268);
and U5943 (N_5943,N_288,N_907);
or U5944 (N_5944,N_1317,N_3130);
and U5945 (N_5945,N_1332,N_4224);
xor U5946 (N_5946,N_2018,N_2778);
and U5947 (N_5947,N_2868,N_4093);
nor U5948 (N_5948,N_1405,N_3785);
nand U5949 (N_5949,N_2888,N_4512);
and U5950 (N_5950,N_1989,N_4529);
nand U5951 (N_5951,N_2714,N_4159);
nor U5952 (N_5952,N_919,N_4135);
nor U5953 (N_5953,N_73,N_3232);
and U5954 (N_5954,N_2482,N_1137);
and U5955 (N_5955,N_4219,N_4390);
nand U5956 (N_5956,N_1067,N_3840);
xnor U5957 (N_5957,N_839,N_3280);
or U5958 (N_5958,N_2822,N_4834);
nor U5959 (N_5959,N_3706,N_1770);
nand U5960 (N_5960,N_1522,N_2101);
nor U5961 (N_5961,N_229,N_2431);
or U5962 (N_5962,N_1951,N_4031);
xnor U5963 (N_5963,N_2723,N_4661);
and U5964 (N_5964,N_3871,N_4098);
nand U5965 (N_5965,N_2169,N_266);
xor U5966 (N_5966,N_2293,N_132);
nand U5967 (N_5967,N_2267,N_4832);
nor U5968 (N_5968,N_2022,N_4571);
and U5969 (N_5969,N_2254,N_2196);
and U5970 (N_5970,N_2841,N_306);
or U5971 (N_5971,N_3771,N_1271);
nand U5972 (N_5972,N_1611,N_4431);
nor U5973 (N_5973,N_979,N_1266);
xor U5974 (N_5974,N_955,N_716);
and U5975 (N_5975,N_4352,N_4420);
xor U5976 (N_5976,N_2230,N_53);
or U5977 (N_5977,N_4708,N_4904);
nand U5978 (N_5978,N_1107,N_1103);
nor U5979 (N_5979,N_272,N_1623);
xor U5980 (N_5980,N_1010,N_2688);
nand U5981 (N_5981,N_2701,N_4690);
or U5982 (N_5982,N_2062,N_4885);
nor U5983 (N_5983,N_155,N_3684);
or U5984 (N_5984,N_372,N_4638);
nor U5985 (N_5985,N_4859,N_4902);
xor U5986 (N_5986,N_71,N_1205);
or U5987 (N_5987,N_4498,N_1170);
or U5988 (N_5988,N_4668,N_1481);
or U5989 (N_5989,N_2743,N_1168);
and U5990 (N_5990,N_3867,N_2735);
and U5991 (N_5991,N_2240,N_2624);
or U5992 (N_5992,N_1065,N_2734);
nor U5993 (N_5993,N_1542,N_1418);
or U5994 (N_5994,N_610,N_3738);
or U5995 (N_5995,N_4481,N_2259);
xor U5996 (N_5996,N_2982,N_1613);
and U5997 (N_5997,N_2832,N_467);
and U5998 (N_5998,N_652,N_2786);
and U5999 (N_5999,N_3851,N_801);
nand U6000 (N_6000,N_4567,N_314);
nand U6001 (N_6001,N_4012,N_415);
and U6002 (N_6002,N_3003,N_1909);
or U6003 (N_6003,N_248,N_429);
nand U6004 (N_6004,N_4756,N_3327);
or U6005 (N_6005,N_4499,N_1298);
xnor U6006 (N_6006,N_927,N_3952);
nand U6007 (N_6007,N_4958,N_2206);
and U6008 (N_6008,N_4900,N_4179);
or U6009 (N_6009,N_4496,N_60);
nor U6010 (N_6010,N_3289,N_1267);
nand U6011 (N_6011,N_4556,N_3677);
xor U6012 (N_6012,N_3372,N_832);
xnor U6013 (N_6013,N_1129,N_688);
or U6014 (N_6014,N_823,N_3285);
or U6015 (N_6015,N_194,N_3857);
nand U6016 (N_6016,N_727,N_1115);
xor U6017 (N_6017,N_455,N_3357);
nand U6018 (N_6018,N_4520,N_443);
nor U6019 (N_6019,N_4528,N_3918);
nand U6020 (N_6020,N_4405,N_3429);
nand U6021 (N_6021,N_3759,N_985);
nor U6022 (N_6022,N_4480,N_668);
and U6023 (N_6023,N_690,N_2608);
nor U6024 (N_6024,N_1903,N_838);
nand U6025 (N_6025,N_4020,N_869);
xnor U6026 (N_6026,N_89,N_1875);
nand U6027 (N_6027,N_1968,N_2796);
or U6028 (N_6028,N_2110,N_2852);
xor U6029 (N_6029,N_1053,N_4115);
nand U6030 (N_6030,N_2952,N_4433);
nand U6031 (N_6031,N_298,N_2761);
nand U6032 (N_6032,N_4563,N_4206);
nor U6033 (N_6033,N_2745,N_4781);
nor U6034 (N_6034,N_3949,N_2833);
or U6035 (N_6035,N_3072,N_3419);
nor U6036 (N_6036,N_2409,N_740);
nor U6037 (N_6037,N_250,N_1301);
or U6038 (N_6038,N_2618,N_2027);
nor U6039 (N_6039,N_4003,N_2806);
and U6040 (N_6040,N_4430,N_1110);
nand U6041 (N_6041,N_2881,N_427);
nor U6042 (N_6042,N_3427,N_824);
nor U6043 (N_6043,N_1353,N_4096);
xor U6044 (N_6044,N_4267,N_2095);
nor U6045 (N_6045,N_1350,N_2047);
xor U6046 (N_6046,N_1458,N_2180);
nand U6047 (N_6047,N_2160,N_2658);
nand U6048 (N_6048,N_3587,N_3394);
xnor U6049 (N_6049,N_2328,N_2983);
nand U6050 (N_6050,N_4313,N_997);
nand U6051 (N_6051,N_1848,N_527);
or U6052 (N_6052,N_2923,N_3442);
xnor U6053 (N_6053,N_3091,N_457);
or U6054 (N_6054,N_4034,N_206);
or U6055 (N_6055,N_4626,N_2604);
and U6056 (N_6056,N_1565,N_1955);
and U6057 (N_6057,N_2907,N_1531);
xor U6058 (N_6058,N_1259,N_2993);
nor U6059 (N_6059,N_1943,N_4795);
xnor U6060 (N_6060,N_3100,N_3006);
xor U6061 (N_6061,N_402,N_765);
xnor U6062 (N_6062,N_2370,N_2675);
or U6063 (N_6063,N_4278,N_3588);
nand U6064 (N_6064,N_3101,N_4590);
and U6065 (N_6065,N_2074,N_2019);
nor U6066 (N_6066,N_950,N_2830);
nor U6067 (N_6067,N_4207,N_1245);
xor U6068 (N_6068,N_4851,N_4350);
xor U6069 (N_6069,N_4369,N_3437);
xor U6070 (N_6070,N_4517,N_891);
xor U6071 (N_6071,N_2021,N_2088);
nor U6072 (N_6072,N_370,N_4386);
nand U6073 (N_6073,N_1862,N_1184);
or U6074 (N_6074,N_3822,N_2116);
or U6075 (N_6075,N_2343,N_571);
or U6076 (N_6076,N_779,N_1282);
nor U6077 (N_6077,N_4580,N_422);
and U6078 (N_6078,N_3472,N_4671);
or U6079 (N_6079,N_2301,N_4672);
nand U6080 (N_6080,N_353,N_667);
and U6081 (N_6081,N_1027,N_2508);
nand U6082 (N_6082,N_2560,N_728);
nand U6083 (N_6083,N_30,N_1780);
nand U6084 (N_6084,N_4523,N_462);
xor U6085 (N_6085,N_488,N_2415);
or U6086 (N_6086,N_768,N_2738);
and U6087 (N_6087,N_502,N_2333);
nor U6088 (N_6088,N_141,N_751);
nand U6089 (N_6089,N_2632,N_1257);
nand U6090 (N_6090,N_431,N_432);
or U6091 (N_6091,N_3982,N_3018);
nand U6092 (N_6092,N_2233,N_4466);
xnor U6093 (N_6093,N_1306,N_1698);
and U6094 (N_6094,N_2380,N_2197);
nor U6095 (N_6095,N_1227,N_2132);
nor U6096 (N_6096,N_1058,N_3921);
xnor U6097 (N_6097,N_1202,N_2866);
xnor U6098 (N_6098,N_151,N_158);
nor U6099 (N_6099,N_1963,N_2477);
and U6100 (N_6100,N_3872,N_893);
or U6101 (N_6101,N_2543,N_1560);
or U6102 (N_6102,N_4618,N_1985);
and U6103 (N_6103,N_230,N_3166);
xor U6104 (N_6104,N_1893,N_2403);
xnor U6105 (N_6105,N_2831,N_1629);
and U6106 (N_6106,N_975,N_1785);
xor U6107 (N_6107,N_79,N_3242);
nor U6108 (N_6108,N_3893,N_15);
and U6109 (N_6109,N_1855,N_439);
or U6110 (N_6110,N_1004,N_1331);
xor U6111 (N_6111,N_4548,N_830);
nor U6112 (N_6112,N_4472,N_293);
nor U6113 (N_6113,N_2932,N_1111);
xnor U6114 (N_6114,N_1819,N_3070);
and U6115 (N_6115,N_1499,N_4951);
nor U6116 (N_6116,N_4025,N_3167);
or U6117 (N_6117,N_197,N_4343);
and U6118 (N_6118,N_3192,N_865);
nand U6119 (N_6119,N_853,N_2316);
xnor U6120 (N_6120,N_3989,N_2096);
nor U6121 (N_6121,N_3602,N_4380);
and U6122 (N_6122,N_1672,N_1690);
nor U6123 (N_6123,N_4051,N_1305);
or U6124 (N_6124,N_960,N_2867);
xor U6125 (N_6125,N_776,N_2548);
nor U6126 (N_6126,N_1196,N_3695);
nor U6127 (N_6127,N_2792,N_3525);
and U6128 (N_6128,N_3383,N_356);
nand U6129 (N_6129,N_4409,N_1523);
nand U6130 (N_6130,N_64,N_3583);
xnor U6131 (N_6131,N_1147,N_3784);
xor U6132 (N_6132,N_459,N_207);
nor U6133 (N_6133,N_1029,N_2742);
nor U6134 (N_6134,N_4573,N_3941);
or U6135 (N_6135,N_4953,N_2008);
nor U6136 (N_6136,N_3882,N_4111);
or U6137 (N_6137,N_3098,N_2277);
nand U6138 (N_6138,N_4663,N_4375);
or U6139 (N_6139,N_1825,N_1061);
nor U6140 (N_6140,N_4320,N_362);
nand U6141 (N_6141,N_901,N_4986);
nand U6142 (N_6142,N_1735,N_1688);
nand U6143 (N_6143,N_3555,N_165);
or U6144 (N_6144,N_2413,N_1062);
and U6145 (N_6145,N_2500,N_3795);
xor U6146 (N_6146,N_546,N_548);
nor U6147 (N_6147,N_4621,N_4462);
or U6148 (N_6148,N_1303,N_3464);
xnor U6149 (N_6149,N_2848,N_2069);
nor U6150 (N_6150,N_1337,N_1165);
xnor U6151 (N_6151,N_1351,N_797);
nand U6152 (N_6152,N_4247,N_2869);
xnor U6153 (N_6153,N_333,N_1026);
nand U6154 (N_6154,N_4891,N_980);
nand U6155 (N_6155,N_857,N_3255);
and U6156 (N_6156,N_2385,N_1777);
xnor U6157 (N_6157,N_1617,N_710);
nor U6158 (N_6158,N_4701,N_1217);
xor U6159 (N_6159,N_3497,N_1864);
xor U6160 (N_6160,N_1606,N_4446);
or U6161 (N_6161,N_4972,N_8);
xor U6162 (N_6162,N_2124,N_1956);
or U6163 (N_6163,N_3030,N_3407);
and U6164 (N_6164,N_2607,N_4245);
nand U6165 (N_6165,N_551,N_3685);
and U6166 (N_6166,N_2989,N_3111);
xnor U6167 (N_6167,N_3020,N_1898);
nor U6168 (N_6168,N_1039,N_1832);
nor U6169 (N_6169,N_3625,N_4158);
xor U6170 (N_6170,N_3629,N_1990);
or U6171 (N_6171,N_3696,N_1364);
nand U6172 (N_6172,N_4574,N_2475);
or U6173 (N_6173,N_4056,N_4166);
or U6174 (N_6174,N_1140,N_767);
xnor U6175 (N_6175,N_1323,N_3146);
xor U6176 (N_6176,N_234,N_1982);
xnor U6177 (N_6177,N_1037,N_106);
nand U6178 (N_6178,N_4901,N_2904);
and U6179 (N_6179,N_4104,N_4118);
or U6180 (N_6180,N_4974,N_614);
nand U6181 (N_6181,N_2300,N_2692);
nand U6182 (N_6182,N_3023,N_706);
xor U6183 (N_6183,N_4358,N_3827);
nand U6184 (N_6184,N_3454,N_4527);
nand U6185 (N_6185,N_917,N_1775);
nand U6186 (N_6186,N_3065,N_4975);
nor U6187 (N_6187,N_2006,N_1075);
and U6188 (N_6188,N_4109,N_35);
nor U6189 (N_6189,N_4205,N_107);
or U6190 (N_6190,N_3369,N_713);
or U6191 (N_6191,N_4165,N_2651);
xor U6192 (N_6192,N_2650,N_238);
nor U6193 (N_6193,N_1042,N_2660);
nand U6194 (N_6194,N_468,N_4619);
or U6195 (N_6195,N_3705,N_1947);
or U6196 (N_6196,N_695,N_3028);
xor U6197 (N_6197,N_4910,N_4270);
xnor U6198 (N_6198,N_1941,N_3498);
xnor U6199 (N_6199,N_3888,N_1430);
nor U6200 (N_6200,N_611,N_1374);
xor U6201 (N_6201,N_2051,N_2997);
xnor U6202 (N_6202,N_149,N_1089);
and U6203 (N_6203,N_13,N_2598);
xnor U6204 (N_6204,N_1599,N_2721);
and U6205 (N_6205,N_2111,N_2876);
xnor U6206 (N_6206,N_493,N_2882);
and U6207 (N_6207,N_4611,N_2656);
or U6208 (N_6208,N_3258,N_3661);
and U6209 (N_6209,N_4265,N_941);
or U6210 (N_6210,N_4226,N_387);
xor U6211 (N_6211,N_2564,N_4918);
nor U6212 (N_6212,N_3102,N_3703);
nand U6213 (N_6213,N_3305,N_4984);
xnor U6214 (N_6214,N_62,N_4730);
or U6215 (N_6215,N_4941,N_2495);
nand U6216 (N_6216,N_4759,N_3040);
and U6217 (N_6217,N_3064,N_1408);
or U6218 (N_6218,N_4808,N_3446);
nand U6219 (N_6219,N_1390,N_4667);
xnor U6220 (N_6220,N_3972,N_1608);
xnor U6221 (N_6221,N_783,N_2331);
xnor U6222 (N_6222,N_4200,N_769);
nor U6223 (N_6223,N_2373,N_4861);
xnor U6224 (N_6224,N_4124,N_4616);
and U6225 (N_6225,N_786,N_4653);
or U6226 (N_6226,N_3530,N_1077);
nand U6227 (N_6227,N_276,N_2784);
nand U6228 (N_6228,N_3313,N_2351);
nand U6229 (N_6229,N_4677,N_4342);
xor U6230 (N_6230,N_682,N_2783);
nor U6231 (N_6231,N_3605,N_1604);
nand U6232 (N_6232,N_2397,N_3395);
xnor U6233 (N_6233,N_2702,N_2040);
or U6234 (N_6234,N_408,N_239);
and U6235 (N_6235,N_2322,N_1678);
nand U6236 (N_6236,N_1310,N_2953);
xnor U6237 (N_6237,N_2402,N_665);
nor U6238 (N_6238,N_2528,N_1843);
xor U6239 (N_6239,N_1692,N_1427);
nor U6240 (N_6240,N_1343,N_2303);
or U6241 (N_6241,N_4188,N_57);
xor U6242 (N_6242,N_582,N_4575);
nand U6243 (N_6243,N_1131,N_964);
nor U6244 (N_6244,N_2775,N_4083);
and U6245 (N_6245,N_1117,N_129);
and U6246 (N_6246,N_193,N_4950);
and U6247 (N_6247,N_1630,N_2501);
nand U6248 (N_6248,N_3392,N_1175);
nand U6249 (N_6249,N_3692,N_680);
xor U6250 (N_6250,N_34,N_4998);
xor U6251 (N_6251,N_423,N_4643);
xor U6252 (N_6252,N_4069,N_4463);
or U6253 (N_6253,N_458,N_4339);
or U6254 (N_6254,N_3889,N_2479);
or U6255 (N_6255,N_3484,N_1452);
nor U6256 (N_6256,N_2348,N_781);
xor U6257 (N_6257,N_3954,N_1116);
or U6258 (N_6258,N_5,N_1660);
and U6259 (N_6259,N_4680,N_1671);
xor U6260 (N_6260,N_1749,N_999);
and U6261 (N_6261,N_2291,N_3914);
nor U6262 (N_6262,N_2450,N_703);
or U6263 (N_6263,N_4539,N_3301);
or U6264 (N_6264,N_1781,N_1800);
or U6265 (N_6265,N_894,N_3841);
nor U6266 (N_6266,N_1318,N_1121);
xnor U6267 (N_6267,N_1093,N_2041);
xnor U6268 (N_6268,N_4411,N_2515);
xnor U6269 (N_6269,N_4855,N_4981);
nor U6270 (N_6270,N_474,N_572);
nand U6271 (N_6271,N_4755,N_2148);
or U6272 (N_6272,N_3171,N_2803);
xor U6273 (N_6273,N_1657,N_1589);
xnor U6274 (N_6274,N_4631,N_4277);
nand U6275 (N_6275,N_598,N_4625);
nand U6276 (N_6276,N_1097,N_1263);
nor U6277 (N_6277,N_204,N_4692);
nor U6278 (N_6278,N_4180,N_959);
and U6279 (N_6279,N_4739,N_3862);
xnor U6280 (N_6280,N_101,N_2762);
xnor U6281 (N_6281,N_476,N_3656);
nand U6282 (N_6282,N_284,N_1108);
and U6283 (N_6283,N_2473,N_1635);
or U6284 (N_6284,N_1002,N_653);
nand U6285 (N_6285,N_675,N_4309);
nand U6286 (N_6286,N_1568,N_1090);
nand U6287 (N_6287,N_2865,N_974);
and U6288 (N_6288,N_555,N_49);
nor U6289 (N_6289,N_171,N_2428);
nand U6290 (N_6290,N_4441,N_4825);
or U6291 (N_6291,N_4550,N_2712);
and U6292 (N_6292,N_22,N_1779);
and U6293 (N_6293,N_4856,N_1455);
and U6294 (N_6294,N_3031,N_2159);
xnor U6295 (N_6295,N_2995,N_1891);
and U6296 (N_6296,N_2489,N_94);
xor U6297 (N_6297,N_4632,N_4835);
and U6298 (N_6298,N_553,N_203);
or U6299 (N_6299,N_4292,N_1397);
xor U6300 (N_6300,N_407,N_3129);
nand U6301 (N_6301,N_1270,N_1448);
nand U6302 (N_6302,N_2446,N_3604);
and U6303 (N_6303,N_1426,N_4304);
nor U6304 (N_6304,N_4131,N_4717);
nand U6305 (N_6305,N_3723,N_3832);
or U6306 (N_6306,N_600,N_2966);
and U6307 (N_6307,N_1546,N_4455);
or U6308 (N_6308,N_4983,N_2950);
xor U6309 (N_6309,N_793,N_2306);
nand U6310 (N_6310,N_19,N_4956);
or U6311 (N_6311,N_718,N_4415);
nand U6312 (N_6312,N_181,N_2642);
nand U6313 (N_6313,N_1677,N_2914);
xnor U6314 (N_6314,N_1459,N_995);
and U6315 (N_6315,N_4167,N_3381);
nand U6316 (N_6316,N_3760,N_2793);
xnor U6317 (N_6317,N_3690,N_2097);
and U6318 (N_6318,N_1420,N_2036);
xor U6319 (N_6319,N_1649,N_3371);
nor U6320 (N_6320,N_4562,N_2452);
nor U6321 (N_6321,N_4340,N_2819);
nand U6322 (N_6322,N_1171,N_1959);
xnor U6323 (N_6323,N_2324,N_1846);
and U6324 (N_6324,N_1754,N_2522);
and U6325 (N_6325,N_516,N_4635);
nand U6326 (N_6326,N_3202,N_4000);
and U6327 (N_6327,N_4432,N_3635);
or U6328 (N_6328,N_878,N_2071);
xor U6329 (N_6329,N_2687,N_2158);
xor U6330 (N_6330,N_3662,N_1850);
xnor U6331 (N_6331,N_2091,N_4830);
nor U6332 (N_6332,N_1475,N_670);
xor U6333 (N_6333,N_4955,N_1667);
xnor U6334 (N_6334,N_3698,N_1225);
nand U6335 (N_6335,N_4407,N_1194);
nor U6336 (N_6336,N_3885,N_3798);
or U6337 (N_6337,N_2102,N_4533);
xnor U6338 (N_6338,N_228,N_1653);
nand U6339 (N_6339,N_2025,N_4502);
nand U6340 (N_6340,N_1339,N_971);
or U6341 (N_6341,N_164,N_1707);
xor U6342 (N_6342,N_1748,N_39);
nand U6343 (N_6343,N_1363,N_3775);
nand U6344 (N_6344,N_2931,N_1433);
nand U6345 (N_6345,N_2573,N_2903);
nor U6346 (N_6346,N_2558,N_2172);
or U6347 (N_6347,N_251,N_1284);
and U6348 (N_6348,N_4943,N_4561);
nor U6349 (N_6349,N_3436,N_3256);
xor U6350 (N_6350,N_1421,N_2750);
xor U6351 (N_6351,N_3263,N_515);
and U6352 (N_6352,N_4251,N_1398);
nor U6353 (N_6353,N_1509,N_2587);
nand U6354 (N_6354,N_1057,N_441);
xnor U6355 (N_6355,N_2173,N_930);
xnor U6356 (N_6356,N_4094,N_1329);
xnor U6357 (N_6357,N_2620,N_2856);
and U6358 (N_6358,N_2999,N_3078);
nor U6359 (N_6359,N_3971,N_1304);
nor U6360 (N_6360,N_1878,N_2367);
or U6361 (N_6361,N_4534,N_3574);
or U6362 (N_6362,N_1708,N_3239);
xnor U6363 (N_6363,N_1808,N_1948);
xnor U6364 (N_6364,N_3627,N_4979);
xnor U6365 (N_6365,N_1197,N_3839);
xor U6366 (N_6366,N_4875,N_4839);
xor U6367 (N_6367,N_1361,N_1811);
and U6368 (N_6368,N_188,N_4728);
and U6369 (N_6369,N_2563,N_3051);
and U6370 (N_6370,N_4259,N_948);
nand U6371 (N_6371,N_4797,N_2958);
and U6372 (N_6372,N_3630,N_3250);
nor U6373 (N_6373,N_2190,N_2628);
nand U6374 (N_6374,N_2383,N_133);
xnor U6375 (N_6375,N_2406,N_4648);
nand U6376 (N_6376,N_1360,N_1466);
nand U6377 (N_6377,N_2610,N_4558);
nand U6378 (N_6378,N_3786,N_3158);
nor U6379 (N_6379,N_4329,N_3138);
nor U6380 (N_6380,N_1826,N_2364);
xnor U6381 (N_6381,N_2674,N_3097);
or U6382 (N_6382,N_1727,N_2117);
nor U6383 (N_6383,N_3315,N_1188);
or U6384 (N_6384,N_2782,N_694);
xor U6385 (N_6385,N_3001,N_719);
nor U6386 (N_6386,N_2777,N_2638);
nor U6387 (N_6387,N_2840,N_2947);
xor U6388 (N_6388,N_539,N_1834);
and U6389 (N_6389,N_1704,N_2014);
or U6390 (N_6390,N_3894,N_4204);
nor U6391 (N_6391,N_4917,N_1289);
nand U6392 (N_6392,N_2458,N_788);
and U6393 (N_6393,N_227,N_4467);
nand U6394 (N_6394,N_698,N_2216);
and U6395 (N_6395,N_4473,N_1979);
or U6396 (N_6396,N_1283,N_52);
nand U6397 (N_6397,N_860,N_4394);
or U6398 (N_6398,N_1633,N_4444);
and U6399 (N_6399,N_2873,N_4176);
or U6400 (N_6400,N_1999,N_2617);
or U6401 (N_6401,N_32,N_4129);
xor U6402 (N_6402,N_4146,N_1543);
xor U6403 (N_6403,N_3801,N_4991);
or U6404 (N_6404,N_4778,N_3126);
and U6405 (N_6405,N_3780,N_1626);
and U6406 (N_6406,N_2374,N_2874);
and U6407 (N_6407,N_3338,N_1931);
nand U6408 (N_6408,N_820,N_1394);
nand U6409 (N_6409,N_1241,N_3756);
nand U6410 (N_6410,N_631,N_2780);
or U6411 (N_6411,N_1794,N_3331);
nand U6412 (N_6412,N_4630,N_3095);
nand U6413 (N_6413,N_4211,N_105);
nor U6414 (N_6414,N_4620,N_258);
and U6415 (N_6415,N_4408,N_3640);
or U6416 (N_6416,N_4777,N_916);
xor U6417 (N_6417,N_2917,N_2000);
or U6418 (N_6418,N_3856,N_4584);
and U6419 (N_6419,N_3193,N_4142);
or U6420 (N_6420,N_4357,N_343);
or U6421 (N_6421,N_495,N_1782);
nand U6422 (N_6422,N_2453,N_3415);
xnor U6423 (N_6423,N_2208,N_4538);
nor U6424 (N_6424,N_1845,N_1384);
or U6425 (N_6425,N_3821,N_3054);
nor U6426 (N_6426,N_1274,N_1505);
nand U6427 (N_6427,N_4089,N_3968);
and U6428 (N_6428,N_1938,N_405);
nand U6429 (N_6429,N_3183,N_3529);
xor U6430 (N_6430,N_4780,N_4393);
or U6431 (N_6431,N_1839,N_161);
or U6432 (N_6432,N_1432,N_3491);
nand U6433 (N_6433,N_2075,N_2749);
nor U6434 (N_6434,N_4500,N_3540);
or U6435 (N_6435,N_2122,N_4445);
or U6436 (N_6436,N_796,N_815);
and U6437 (N_6437,N_4557,N_4212);
and U6438 (N_6438,N_3447,N_1493);
nand U6439 (N_6439,N_2362,N_2857);
nand U6440 (N_6440,N_2652,N_2562);
nor U6441 (N_6441,N_393,N_2577);
nand U6442 (N_6442,N_583,N_2596);
or U6443 (N_6443,N_2336,N_3215);
nor U6444 (N_6444,N_4886,N_1185);
nand U6445 (N_6445,N_4456,N_4484);
or U6446 (N_6446,N_401,N_3059);
and U6447 (N_6447,N_773,N_487);
and U6448 (N_6448,N_4752,N_2256);
nor U6449 (N_6449,N_1840,N_1783);
and U6450 (N_6450,N_1451,N_2621);
and U6451 (N_6451,N_4033,N_3237);
and U6452 (N_6452,N_743,N_2725);
xnor U6453 (N_6453,N_2191,N_2509);
xor U6454 (N_6454,N_1167,N_4997);
nor U6455 (N_6455,N_1827,N_20);
nor U6456 (N_6456,N_2265,N_4977);
nor U6457 (N_6457,N_369,N_2427);
or U6458 (N_6458,N_472,N_953);
or U6459 (N_6459,N_2844,N_3121);
and U6460 (N_6460,N_640,N_4073);
nand U6461 (N_6461,N_712,N_325);
or U6462 (N_6462,N_4493,N_4568);
nand U6463 (N_6463,N_2113,N_2440);
nor U6464 (N_6464,N_663,N_12);
xnor U6465 (N_6465,N_881,N_2030);
or U6466 (N_6466,N_2534,N_943);
or U6467 (N_6467,N_913,N_4231);
or U6468 (N_6468,N_3007,N_1725);
nand U6469 (N_6469,N_3022,N_4938);
nand U6470 (N_6470,N_3330,N_4070);
nor U6471 (N_6471,N_2549,N_1852);
or U6472 (N_6472,N_2646,N_2626);
and U6473 (N_6473,N_2540,N_3139);
and U6474 (N_6474,N_3319,N_1159);
nor U6475 (N_6475,N_3620,N_1349);
xnor U6476 (N_6476,N_510,N_1605);
and U6477 (N_6477,N_738,N_4662);
nand U6478 (N_6478,N_758,N_2855);
or U6479 (N_6479,N_1181,N_2815);
and U6480 (N_6480,N_1113,N_1880);
nand U6481 (N_6481,N_4878,N_3156);
xor U6482 (N_6482,N_2581,N_537);
xor U6483 (N_6483,N_37,N_2570);
and U6484 (N_6484,N_1441,N_550);
xor U6485 (N_6485,N_3029,N_3618);
nor U6486 (N_6486,N_4801,N_1886);
nor U6487 (N_6487,N_21,N_513);
or U6488 (N_6488,N_2493,N_678);
xor U6489 (N_6489,N_848,N_1697);
nand U6490 (N_6490,N_4813,N_617);
xnor U6491 (N_6491,N_2393,N_1192);
or U6492 (N_6492,N_176,N_1011);
xnor U6493 (N_6493,N_3807,N_2797);
xnor U6494 (N_6494,N_3796,N_1345);
xor U6495 (N_6495,N_3853,N_4426);
nor U6496 (N_6496,N_1327,N_799);
xnor U6497 (N_6497,N_4048,N_3009);
xnor U6498 (N_6498,N_2121,N_4468);
xnor U6499 (N_6499,N_3134,N_373);
nor U6500 (N_6500,N_2093,N_2498);
nor U6501 (N_6501,N_1643,N_3238);
and U6502 (N_6502,N_2585,N_2264);
xnor U6503 (N_6503,N_1392,N_4241);
xor U6504 (N_6504,N_1362,N_1254);
nand U6505 (N_6505,N_2644,N_2223);
nand U6506 (N_6506,N_1682,N_576);
nand U6507 (N_6507,N_1730,N_970);
and U6508 (N_6508,N_1750,N_3994);
nor U6509 (N_6509,N_4349,N_296);
nor U6510 (N_6510,N_3752,N_1598);
and U6511 (N_6511,N_2599,N_4821);
or U6512 (N_6512,N_4018,N_2280);
or U6513 (N_6513,N_1675,N_4494);
or U6514 (N_6514,N_295,N_3244);
nand U6515 (N_6515,N_552,N_1476);
or U6516 (N_6516,N_992,N_2395);
or U6517 (N_6517,N_4932,N_3663);
nand U6518 (N_6518,N_3052,N_1469);
nand U6519 (N_6519,N_723,N_4607);
and U6520 (N_6520,N_4838,N_2823);
nor U6521 (N_6521,N_2566,N_4311);
xnor U6522 (N_6522,N_2467,N_4812);
and U6523 (N_6523,N_580,N_2274);
nor U6524 (N_6524,N_1028,N_4659);
xnor U6525 (N_6525,N_1752,N_1328);
nor U6526 (N_6526,N_1340,N_4001);
nand U6527 (N_6527,N_4820,N_1155);
nor U6528 (N_6528,N_2314,N_447);
xor U6529 (N_6529,N_1566,N_4791);
xor U6530 (N_6530,N_2788,N_983);
xor U6531 (N_6531,N_4470,N_3719);
nand U6532 (N_6532,N_2580,N_2307);
nor U6533 (N_6533,N_775,N_2707);
nor U6534 (N_6534,N_1201,N_642);
xnor U6535 (N_6535,N_4461,N_3790);
nor U6536 (N_6536,N_2635,N_4435);
or U6537 (N_6537,N_139,N_69);
xor U6538 (N_6538,N_873,N_3776);
nor U6539 (N_6539,N_135,N_126);
xnor U6540 (N_6540,N_2236,N_4601);
or U6541 (N_6541,N_154,N_4513);
nor U6542 (N_6542,N_3467,N_4062);
nand U6543 (N_6543,N_1570,N_3642);
xnor U6544 (N_6544,N_1296,N_2487);
and U6545 (N_6545,N_1151,N_2709);
xnor U6546 (N_6546,N_4546,N_4940);
nor U6547 (N_6547,N_591,N_3418);
or U6548 (N_6548,N_3714,N_1885);
xor U6549 (N_6549,N_1256,N_3172);
xor U6550 (N_6550,N_1215,N_3726);
nand U6551 (N_6551,N_3878,N_3859);
nor U6552 (N_6552,N_3644,N_2241);
xor U6553 (N_6553,N_1790,N_2287);
nor U6554 (N_6554,N_4872,N_1300);
or U6555 (N_6555,N_115,N_1417);
nor U6556 (N_6556,N_2057,N_2825);
nand U6557 (N_6557,N_3631,N_4134);
and U6558 (N_6558,N_2285,N_490);
xnor U6559 (N_6559,N_3351,N_4422);
or U6560 (N_6560,N_3013,N_4353);
and U6561 (N_6561,N_3208,N_121);
and U6562 (N_6562,N_3916,N_1287);
and U6563 (N_6563,N_3364,N_4009);
or U6564 (N_6564,N_75,N_3958);
xor U6565 (N_6565,N_4905,N_1640);
nor U6566 (N_6566,N_2956,N_2207);
or U6567 (N_6567,N_3957,N_2060);
nand U6568 (N_6568,N_3049,N_363);
nand U6569 (N_6569,N_6,N_2711);
nand U6570 (N_6570,N_2648,N_1070);
nand U6571 (N_6571,N_535,N_2010);
and U6572 (N_6572,N_1715,N_2435);
nand U6573 (N_6573,N_282,N_4289);
nand U6574 (N_6574,N_593,N_3317);
xnor U6575 (N_6575,N_109,N_1228);
xnor U6576 (N_6576,N_1946,N_1407);
and U6577 (N_6577,N_1138,N_1207);
nand U6578 (N_6578,N_4105,N_2460);
and U6579 (N_6579,N_3868,N_2768);
xnor U6580 (N_6580,N_637,N_554);
or U6581 (N_6581,N_679,N_3835);
nor U6582 (N_6582,N_1933,N_3597);
or U6583 (N_6583,N_3217,N_1631);
nand U6584 (N_6584,N_2289,N_249);
or U6585 (N_6585,N_1178,N_563);
nor U6586 (N_6586,N_1920,N_3384);
and U6587 (N_6587,N_327,N_4004);
xnor U6588 (N_6588,N_3005,N_2162);
xnor U6589 (N_6589,N_3844,N_2200);
and U6590 (N_6590,N_2089,N_864);
xnor U6591 (N_6591,N_558,N_3304);
and U6592 (N_6592,N_3373,N_4198);
or U6593 (N_6593,N_1663,N_2814);
nor U6594 (N_6594,N_4578,N_4081);
xor U6595 (N_6595,N_3984,N_885);
xnor U6596 (N_6596,N_4333,N_2776);
xor U6597 (N_6597,N_3346,N_1788);
or U6598 (N_6598,N_687,N_1486);
and U6599 (N_6599,N_1086,N_708);
or U6600 (N_6600,N_3322,N_2805);
xnor U6601 (N_6601,N_3905,N_4602);
nor U6602 (N_6602,N_2028,N_4214);
nand U6603 (N_6603,N_125,N_2462);
or U6604 (N_6604,N_1532,N_1809);
nand U6605 (N_6605,N_2465,N_3033);
nor U6606 (N_6606,N_4075,N_2099);
xnor U6607 (N_6607,N_3055,N_4804);
xor U6608 (N_6608,N_2835,N_1930);
and U6609 (N_6609,N_912,N_1534);
nand U6610 (N_6610,N_3948,N_2114);
nor U6611 (N_6611,N_3099,N_1732);
xor U6612 (N_6612,N_609,N_235);
and U6613 (N_6613,N_3162,N_3709);
or U6614 (N_6614,N_4714,N_1701);
and U6615 (N_6615,N_1445,N_95);
nor U6616 (N_6616,N_3547,N_1712);
nor U6617 (N_6617,N_4269,N_3507);
xor U6618 (N_6618,N_1733,N_426);
xnor U6619 (N_6619,N_4335,N_2471);
and U6620 (N_6620,N_1844,N_2963);
nand U6621 (N_6621,N_2517,N_3046);
xor U6622 (N_6622,N_240,N_3262);
or U6623 (N_6623,N_4831,N_1412);
and U6624 (N_6624,N_3810,N_2174);
nand U6625 (N_6625,N_2229,N_112);
or U6626 (N_6626,N_3990,N_1040);
and U6627 (N_6627,N_3514,N_219);
xor U6628 (N_6628,N_816,N_2605);
and U6629 (N_6629,N_4092,N_433);
or U6630 (N_6630,N_2286,N_1261);
and U6631 (N_6631,N_352,N_4603);
xor U6632 (N_6632,N_44,N_40);
nand U6633 (N_6633,N_3757,N_840);
xnor U6634 (N_6634,N_3011,N_4140);
and U6635 (N_6635,N_2708,N_3953);
or U6636 (N_6636,N_3410,N_741);
or U6637 (N_6637,N_1193,N_2023);
nand U6638 (N_6638,N_669,N_3385);
nor U6639 (N_6639,N_4315,N_4844);
and U6640 (N_6640,N_4633,N_3140);
and U6641 (N_6641,N_602,N_1652);
nand U6642 (N_6642,N_1223,N_1588);
or U6643 (N_6643,N_1661,N_1600);
nand U6644 (N_6644,N_2326,N_2804);
xnor U6645 (N_6645,N_1132,N_2550);
or U6646 (N_6646,N_1109,N_2794);
xnor U6647 (N_6647,N_394,N_722);
nand U6648 (N_6648,N_518,N_726);
and U6649 (N_6649,N_2578,N_564);
and U6650 (N_6650,N_4043,N_2392);
xor U6651 (N_6651,N_1036,N_3090);
nor U6652 (N_6652,N_3817,N_4510);
nand U6653 (N_6653,N_4990,N_3552);
nor U6654 (N_6654,N_3457,N_1487);
xor U6655 (N_6655,N_634,N_2420);
nand U6656 (N_6656,N_2664,N_4647);
nand U6657 (N_6657,N_3585,N_3235);
or U6658 (N_6658,N_2275,N_3594);
or U6659 (N_6659,N_3944,N_1899);
and U6660 (N_6660,N_1764,N_3570);
xnor U6661 (N_6661,N_2198,N_4911);
or U6662 (N_6662,N_2961,N_3670);
nand U6663 (N_6663,N_3886,N_3349);
and U6664 (N_6664,N_3774,N_3452);
nor U6665 (N_6665,N_2050,N_1444);
or U6666 (N_6666,N_4321,N_3569);
and U6667 (N_6667,N_3343,N_473);
xnor U6668 (N_6668,N_590,N_871);
and U6669 (N_6669,N_4438,N_4174);
or U6670 (N_6670,N_896,N_270);
nor U6671 (N_6671,N_2799,N_186);
or U6672 (N_6672,N_1887,N_1984);
xor U6673 (N_6673,N_4054,N_2430);
nand U6674 (N_6674,N_3147,N_104);
nor U6675 (N_6675,N_4762,N_4506);
and U6676 (N_6676,N_51,N_4372);
xor U6677 (N_6677,N_1429,N_3688);
and U6678 (N_6678,N_2457,N_1603);
and U6679 (N_6679,N_1158,N_4132);
nand U6680 (N_6680,N_4149,N_380);
or U6681 (N_6681,N_3858,N_714);
nor U6682 (N_6682,N_1302,N_4947);
nor U6683 (N_6683,N_2954,N_771);
xnor U6684 (N_6684,N_1902,N_350);
nor U6685 (N_6685,N_3985,N_2276);
xor U6686 (N_6686,N_2891,N_605);
nand U6687 (N_6687,N_3316,N_3892);
and U6688 (N_6688,N_3341,N_3578);
and U6689 (N_6689,N_1833,N_1308);
nand U6690 (N_6690,N_3829,N_150);
and U6691 (N_6691,N_3490,N_846);
or U6692 (N_6692,N_177,N_1025);
nor U6693 (N_6693,N_3241,N_4050);
xnor U6694 (N_6694,N_1716,N_2011);
xnor U6695 (N_6695,N_1961,N_3428);
or U6696 (N_6696,N_2937,N_737);
or U6697 (N_6697,N_4028,N_625);
xnor U6698 (N_6698,N_1320,N_4449);
nand U6699 (N_6699,N_4100,N_1017);
and U6700 (N_6700,N_2270,N_2541);
xor U6701 (N_6701,N_1136,N_886);
nand U6702 (N_6702,N_4011,N_3880);
nand U6703 (N_6703,N_244,N_54);
nand U6704 (N_6704,N_144,N_1680);
nor U6705 (N_6705,N_3314,N_3522);
xnor U6706 (N_6706,N_2948,N_336);
and U6707 (N_6707,N_2043,N_2899);
xor U6708 (N_6708,N_2854,N_3701);
and U6709 (N_6709,N_1970,N_1586);
xor U6710 (N_6710,N_1295,N_3865);
nand U6711 (N_6711,N_3267,N_2756);
and U6712 (N_6712,N_790,N_305);
xor U6713 (N_6713,N_4264,N_4145);
xnor U6714 (N_6714,N_925,N_2480);
nor U6715 (N_6715,N_711,N_3356);
nor U6716 (N_6716,N_2916,N_4039);
xnor U6717 (N_6717,N_3612,N_2298);
or U6718 (N_6718,N_254,N_451);
nand U6719 (N_6719,N_3359,N_2897);
and U6720 (N_6720,N_4884,N_371);
nor U6721 (N_6721,N_131,N_3846);
nor U6722 (N_6722,N_1936,N_3584);
and U6723 (N_6723,N_4784,N_2600);
or U6724 (N_6724,N_664,N_1798);
and U6725 (N_6725,N_1913,N_4378);
or U6726 (N_6726,N_968,N_1907);
or U6727 (N_6727,N_1018,N_2520);
and U6728 (N_6728,N_660,N_355);
or U6729 (N_6729,N_3930,N_3332);
or U6730 (N_6730,N_2292,N_2491);
nand U6731 (N_6731,N_4907,N_1865);
nor U6732 (N_6732,N_2700,N_3236);
xnor U6733 (N_6733,N_453,N_4987);
nor U6734 (N_6734,N_1431,N_4588);
nand U6735 (N_6735,N_2893,N_2145);
xor U6736 (N_6736,N_2967,N_1739);
or U6737 (N_6737,N_4185,N_2103);
and U6738 (N_6738,N_4254,N_4301);
and U6739 (N_6739,N_3943,N_4371);
or U6740 (N_6740,N_1226,N_130);
or U6741 (N_6741,N_191,N_525);
and U6742 (N_6742,N_1099,N_2895);
xor U6743 (N_6743,N_1150,N_928);
nor U6744 (N_6744,N_3881,N_2647);
and U6745 (N_6745,N_2813,N_18);
xor U6746 (N_6746,N_585,N_2339);
nor U6747 (N_6747,N_2542,N_501);
nand U6748 (N_6748,N_1395,N_3966);
and U6749 (N_6749,N_1670,N_3988);
and U6750 (N_6750,N_641,N_1082);
or U6751 (N_6751,N_1213,N_253);
or U6752 (N_6752,N_2985,N_3925);
nor U6753 (N_6753,N_1714,N_1755);
and U6754 (N_6754,N_1747,N_3056);
xor U6755 (N_6755,N_1742,N_26);
or U6756 (N_6756,N_398,N_648);
nor U6757 (N_6757,N_2839,N_1632);
and U6758 (N_6758,N_365,N_3453);
or U6759 (N_6759,N_1152,N_4072);
nand U6760 (N_6760,N_4465,N_184);
or U6761 (N_6761,N_2258,N_3758);
xor U6762 (N_6762,N_1161,N_3004);
and U6763 (N_6763,N_3571,N_1500);
nor U6764 (N_6764,N_3145,N_4316);
xor U6765 (N_6765,N_1563,N_828);
nor U6766 (N_6766,N_4530,N_1141);
nand U6767 (N_6767,N_1718,N_1944);
and U6768 (N_6768,N_1597,N_1479);
or U6769 (N_6769,N_4908,N_616);
xor U6770 (N_6770,N_3613,N_2151);
nand U6771 (N_6771,N_4688,N_2837);
or U6772 (N_6772,N_303,N_3233);
or U6773 (N_6773,N_4961,N_3647);
xnor U6774 (N_6774,N_3408,N_4057);
and U6775 (N_6775,N_4536,N_573);
xor U6776 (N_6776,N_4037,N_2201);
nor U6777 (N_6777,N_390,N_1022);
and U6778 (N_6778,N_2411,N_1232);
or U6779 (N_6779,N_2232,N_1925);
nor U6780 (N_6780,N_3461,N_2375);
nand U6781 (N_6781,N_1143,N_4361);
xor U6782 (N_6782,N_2536,N_4840);
nor U6783 (N_6783,N_867,N_2713);
and U6784 (N_6784,N_497,N_1081);
nor U6785 (N_6785,N_2002,N_2634);
xor U6786 (N_6786,N_4796,N_1528);
nand U6787 (N_6787,N_4516,N_3935);
xnor U6788 (N_6788,N_2991,N_1470);
and U6789 (N_6789,N_3668,N_4765);
xor U6790 (N_6790,N_173,N_29);
xnor U6791 (N_6791,N_915,N_4196);
and U6792 (N_6792,N_1573,N_4126);
and U6793 (N_6793,N_236,N_1023);
nor U6794 (N_6794,N_4202,N_1244);
nand U6795 (N_6795,N_3653,N_4629);
nor U6796 (N_6796,N_2031,N_2072);
and U6797 (N_6797,N_541,N_4555);
nand U6798 (N_6798,N_252,N_279);
and U6799 (N_6799,N_565,N_818);
or U6800 (N_6800,N_659,N_3850);
or U6801 (N_6801,N_500,N_68);
or U6802 (N_6802,N_1358,N_3747);
xnor U6803 (N_6803,N_2443,N_588);
nand U6804 (N_6804,N_646,N_1220);
xor U6805 (N_6805,N_808,N_1998);
or U6806 (N_6806,N_1045,N_1019);
or U6807 (N_6807,N_3144,N_1713);
or U6808 (N_6808,N_4030,N_3087);
xnor U6809 (N_6809,N_3533,N_3974);
nand U6810 (N_6810,N_3502,N_3105);
xor U6811 (N_6811,N_3489,N_4645);
nand U6812 (N_6812,N_3899,N_3922);
and U6813 (N_6813,N_1367,N_1462);
xor U6814 (N_6814,N_545,N_2424);
xnor U6815 (N_6815,N_1993,N_2378);
and U6816 (N_6816,N_3227,N_152);
nor U6817 (N_6817,N_127,N_385);
nor U6818 (N_6818,N_4705,N_2582);
or U6819 (N_6819,N_1628,N_3940);
xor U6820 (N_6820,N_3074,N_4982);
and U6821 (N_6821,N_1273,N_4102);
or U6822 (N_6822,N_4595,N_2067);
nand U6823 (N_6823,N_3000,N_1940);
xor U6824 (N_6824,N_4055,N_4471);
xnor U6825 (N_6825,N_577,N_4605);
and U6826 (N_6826,N_185,N_4944);
xnor U6827 (N_6827,N_4504,N_172);
xnor U6828 (N_6828,N_4937,N_3527);
or U6829 (N_6829,N_647,N_4240);
xnor U6830 (N_6830,N_1247,N_449);
and U6831 (N_6831,N_3025,N_4193);
xnor U6832 (N_6832,N_4846,N_3251);
xnor U6833 (N_6833,N_2514,N_3713);
or U6834 (N_6834,N_2583,N_4761);
xnor U6835 (N_6835,N_319,N_1368);
nand U6836 (N_6836,N_994,N_3021);
and U6837 (N_6837,N_4015,N_1044);
xor U6838 (N_6838,N_4282,N_4485);
nand U6839 (N_6839,N_2763,N_2320);
nand U6840 (N_6840,N_4230,N_575);
nand U6841 (N_6841,N_3755,N_2601);
and U6842 (N_6842,N_1761,N_3599);
or U6843 (N_6843,N_2231,N_2902);
or U6844 (N_6844,N_310,N_3141);
and U6845 (N_6845,N_4933,N_3993);
or U6846 (N_6846,N_1942,N_4867);
and U6847 (N_6847,N_3073,N_1503);
xor U6848 (N_6848,N_138,N_4138);
nor U6849 (N_6849,N_875,N_595);
and U6850 (N_6850,N_4691,N_42);
and U6851 (N_6851,N_146,N_4712);
nor U6852 (N_6852,N_1723,N_4849);
xor U6853 (N_6853,N_3820,N_2133);
nor U6854 (N_6854,N_1142,N_2939);
xnor U6855 (N_6855,N_2655,N_2187);
nand U6856 (N_6856,N_1823,N_4266);
xor U6857 (N_6857,N_454,N_2747);
nor U6858 (N_6858,N_349,N_3528);
and U6859 (N_6859,N_4080,N_2305);
nand U6860 (N_6860,N_2352,N_2182);
nor U6861 (N_6861,N_2810,N_895);
nor U6862 (N_6862,N_3143,N_1914);
nand U6863 (N_6863,N_1935,N_277);
and U6864 (N_6864,N_86,N_3877);
xnor U6865 (N_6865,N_1524,N_3731);
or U6866 (N_6866,N_638,N_4410);
xor U6867 (N_6867,N_1419,N_2741);
xor U6868 (N_6868,N_2551,N_1206);
nor U6869 (N_6869,N_4235,N_4227);
xnor U6870 (N_6870,N_2827,N_2506);
xnor U6871 (N_6871,N_2081,N_2296);
xnor U6872 (N_6872,N_4684,N_1582);
nor U6873 (N_6873,N_2588,N_2391);
xnor U6874 (N_6874,N_3426,N_1559);
xor U6875 (N_6875,N_221,N_4491);
and U6876 (N_6876,N_2134,N_1521);
nand U6877 (N_6877,N_4582,N_63);
nand U6878 (N_6878,N_3978,N_2249);
nor U6879 (N_6879,N_1119,N_2875);
xnor U6880 (N_6880,N_1330,N_3353);
nand U6881 (N_6881,N_3397,N_3186);
and U6882 (N_6882,N_2142,N_2263);
or U6883 (N_6883,N_3742,N_4969);
nand U6884 (N_6884,N_732,N_4970);
nor U6885 (N_6885,N_2817,N_2616);
xor U6886 (N_6886,N_1759,N_2816);
xor U6887 (N_6887,N_4741,N_841);
or U6888 (N_6888,N_2143,N_2290);
or U6889 (N_6889,N_3190,N_243);
and U6890 (N_6890,N_3082,N_278);
nor U6891 (N_6891,N_4608,N_4967);
nand U6892 (N_6892,N_4773,N_3219);
nand U6893 (N_6893,N_1860,N_2530);
or U6894 (N_6894,N_4866,N_1294);
nand U6895 (N_6895,N_3754,N_1229);
and U6896 (N_6896,N_4881,N_2502);
xnor U6897 (N_6897,N_3673,N_4190);
nor U6898 (N_6898,N_3412,N_677);
nand U6899 (N_6899,N_981,N_949);
nor U6900 (N_6900,N_1838,N_245);
nand U6901 (N_6901,N_2640,N_1130);
or U6902 (N_6902,N_208,N_2363);
and U6903 (N_6903,N_3363,N_2744);
and U6904 (N_6904,N_1423,N_2800);
xnor U6905 (N_6905,N_55,N_1366);
and U6906 (N_6906,N_1760,N_1578);
and U6907 (N_6907,N_3804,N_3947);
and U6908 (N_6908,N_2565,N_3485);
or U6909 (N_6909,N_982,N_3915);
nand U6910 (N_6910,N_1665,N_2911);
or U6911 (N_6911,N_1309,N_3416);
or U6912 (N_6912,N_1179,N_379);
and U6913 (N_6913,N_632,N_1687);
nor U6914 (N_6914,N_2100,N_1088);
xnor U6915 (N_6915,N_1474,N_299);
and U6916 (N_6916,N_3777,N_2611);
nor U6917 (N_6917,N_2342,N_1464);
nor U6918 (N_6918,N_1614,N_1517);
and U6919 (N_6919,N_618,N_4239);
and U6920 (N_6920,N_2894,N_1393);
xnor U6921 (N_6921,N_267,N_2671);
xnor U6922 (N_6922,N_3109,N_1231);
nand U6923 (N_6923,N_1816,N_798);
nor U6924 (N_6924,N_4869,N_3717);
or U6925 (N_6925,N_4949,N_1250);
xor U6926 (N_6926,N_900,N_3185);
xnor U6927 (N_6927,N_4312,N_300);
or U6928 (N_6928,N_2649,N_4679);
nand U6929 (N_6929,N_3782,N_763);
nand U6930 (N_6930,N_3379,N_2955);
or U6931 (N_6931,N_3689,N_854);
xnor U6932 (N_6932,N_4706,N_1526);
and U6933 (N_6933,N_3596,N_1553);
nand U6934 (N_6934,N_4128,N_1849);
xnor U6935 (N_6935,N_4718,N_1854);
nor U6936 (N_6936,N_2448,N_2421);
or U6937 (N_6937,N_3531,N_685);
and U6938 (N_6938,N_725,N_56);
nor U6939 (N_6939,N_489,N_1541);
nand U6940 (N_6940,N_2846,N_461);
or U6941 (N_6941,N_4486,N_4725);
and U6942 (N_6942,N_3298,N_4541);
nor U6943 (N_6943,N_2529,N_2353);
or U6944 (N_6944,N_4579,N_4763);
nor U6945 (N_6945,N_2553,N_2798);
xnor U6946 (N_6946,N_4593,N_2531);
nand U6947 (N_6947,N_4735,N_1144);
or U6948 (N_6948,N_3014,N_3066);
or U6949 (N_6949,N_821,N_1721);
or U6950 (N_6950,N_3076,N_4332);
nor U6951 (N_6951,N_1757,N_905);
and U6952 (N_6952,N_1784,N_1555);
and U6953 (N_6953,N_1208,N_4385);
nand U6954 (N_6954,N_2584,N_2205);
or U6955 (N_6955,N_397,N_3991);
xor U6956 (N_6956,N_2246,N_2812);
xor U6957 (N_6957,N_1449,N_3389);
and U6958 (N_6958,N_1041,N_3271);
nor U6959 (N_6959,N_910,N_3348);
or U6960 (N_6960,N_696,N_1402);
nor U6961 (N_6961,N_4699,N_4169);
nand U6962 (N_6962,N_2417,N_4246);
nor U6963 (N_6963,N_3417,N_4945);
xor U6964 (N_6964,N_3159,N_4803);
or U6965 (N_6965,N_2090,N_2864);
nand U6966 (N_6966,N_3382,N_3923);
nand U6967 (N_6967,N_4045,N_2838);
or U6968 (N_6968,N_3693,N_3189);
and U6969 (N_6969,N_3573,N_4114);
or U6970 (N_6970,N_560,N_2568);
or U6971 (N_6971,N_74,N_1802);
nand U6972 (N_6972,N_1575,N_4143);
or U6973 (N_6973,N_2609,N_825);
nor U6974 (N_6974,N_4298,N_2418);
xor U6975 (N_6975,N_3932,N_4396);
xnor U6976 (N_6976,N_920,N_4760);
nor U6977 (N_6977,N_3365,N_4920);
xor U6978 (N_6978,N_1792,N_1218);
nand U6979 (N_6979,N_3483,N_4402);
nor U6980 (N_6980,N_4347,N_922);
and U6981 (N_6981,N_1127,N_4794);
nor U6982 (N_6982,N_3441,N_3409);
xor U6983 (N_6983,N_3902,N_884);
xnor U6984 (N_6984,N_3170,N_1461);
xnor U6985 (N_6985,N_3825,N_3201);
xnor U6986 (N_6986,N_1252,N_3838);
or U6987 (N_6987,N_2921,N_4182);
and U6988 (N_6988,N_4354,N_4711);
nand U6989 (N_6989,N_4963,N_3675);
xor U6990 (N_6990,N_789,N_1969);
nand U6991 (N_6991,N_592,N_1054);
nor U6992 (N_6992,N_1454,N_2679);
xnor U6993 (N_6993,N_1324,N_1664);
nor U6994 (N_6994,N_4657,N_4888);
and U6995 (N_6995,N_1700,N_1015);
nand U6996 (N_6996,N_174,N_1291);
or U6997 (N_6997,N_3088,N_100);
nor U6998 (N_6998,N_3556,N_4401);
and U6999 (N_6999,N_3213,N_1736);
or U7000 (N_7000,N_3370,N_908);
nand U7001 (N_7001,N_2042,N_2459);
and U7002 (N_7002,N_1520,N_3897);
xor U7003 (N_7003,N_1078,N_4341);
nor U7004 (N_7004,N_2988,N_1325);
xor U7005 (N_7005,N_2037,N_733);
nand U7006 (N_7006,N_2073,N_23);
nor U7007 (N_7007,N_2791,N_2990);
nor U7008 (N_7008,N_3114,N_3621);
nor U7009 (N_7009,N_4751,N_4710);
xnor U7010 (N_7010,N_368,N_3845);
or U7011 (N_7011,N_1016,N_4675);
or U7012 (N_7012,N_315,N_351);
nor U7013 (N_7013,N_88,N_3450);
or U7014 (N_7014,N_4084,N_3603);
and U7015 (N_7015,N_3290,N_159);
nor U7016 (N_7016,N_316,N_2086);
xnor U7017 (N_7017,N_259,N_2327);
or U7018 (N_7018,N_4416,N_977);
nor U7019 (N_7019,N_242,N_1262);
nand U7020 (N_7020,N_4959,N_3240);
or U7021 (N_7021,N_720,N_3651);
nand U7022 (N_7022,N_4841,N_3505);
nand U7023 (N_7023,N_2098,N_1890);
nor U7024 (N_7024,N_933,N_3024);
nand U7025 (N_7025,N_3964,N_1005);
or U7026 (N_7026,N_1411,N_4279);
nor U7027 (N_7027,N_1272,N_906);
or U7028 (N_7028,N_863,N_3600);
xor U7029 (N_7029,N_416,N_2523);
xnor U7030 (N_7030,N_470,N_932);
and U7031 (N_7031,N_2572,N_3180);
nand U7032 (N_7032,N_1987,N_1164);
xor U7033 (N_7033,N_1929,N_4913);
nand U7034 (N_7034,N_4233,N_2318);
or U7035 (N_7035,N_3277,N_4889);
xnor U7036 (N_7036,N_4847,N_414);
and U7037 (N_7037,N_2112,N_4307);
xor U7038 (N_7038,N_3983,N_4793);
or U7039 (N_7039,N_2177,N_1801);
xor U7040 (N_7040,N_1498,N_3295);
xnor U7041 (N_7041,N_2622,N_92);
or U7042 (N_7042,N_1378,N_413);
nor U7043 (N_7043,N_3765,N_4428);
nor U7044 (N_7044,N_4121,N_4809);
or U7045 (N_7045,N_4526,N_3773);
nand U7046 (N_7046,N_3819,N_3911);
xnor U7047 (N_7047,N_717,N_2984);
and U7048 (N_7048,N_3553,N_4740);
or U7049 (N_7049,N_4665,N_1507);
or U7050 (N_7050,N_963,N_4848);
nor U7051 (N_7051,N_735,N_2135);
or U7052 (N_7052,N_4325,N_2637);
nand U7053 (N_7053,N_4919,N_2689);
xor U7054 (N_7054,N_4076,N_3039);
nor U7055 (N_7055,N_4490,N_2883);
or U7056 (N_7056,N_2760,N_1114);
nand U7057 (N_7057,N_2059,N_3671);
nand U7058 (N_7058,N_166,N_4545);
xor U7059 (N_7059,N_4171,N_4095);
or U7060 (N_7060,N_4644,N_1958);
nor U7061 (N_7061,N_3849,N_2575);
nand U7062 (N_7062,N_924,N_4154);
or U7063 (N_7063,N_223,N_3920);
xor U7064 (N_7064,N_2224,N_4732);
nand U7065 (N_7065,N_4077,N_4022);
nand U7066 (N_7066,N_1084,N_2569);
nand U7067 (N_7067,N_4583,N_2252);
xnor U7068 (N_7068,N_1537,N_140);
nor U7069 (N_7069,N_1456,N_1662);
nand U7070 (N_7070,N_620,N_3992);
xnor U7071 (N_7071,N_621,N_1268);
or U7072 (N_7072,N_4877,N_3401);
and U7073 (N_7073,N_1457,N_1442);
nor U7074 (N_7074,N_4178,N_1385);
xnor U7075 (N_7075,N_3781,N_4928);
or U7076 (N_7076,N_3195,N_3333);
nand U7077 (N_7077,N_4544,N_2126);
and U7078 (N_7078,N_566,N_24);
and U7079 (N_7079,N_2556,N_4966);
nand U7080 (N_7080,N_3337,N_1471);
nand U7081 (N_7081,N_4305,N_3580);
xnor U7082 (N_7082,N_715,N_3135);
or U7083 (N_7083,N_1290,N_4537);
xor U7084 (N_7084,N_3157,N_4693);
xor U7085 (N_7085,N_1830,N_3448);
or U7086 (N_7086,N_4106,N_3390);
nor U7087 (N_7087,N_2980,N_1237);
and U7088 (N_7088,N_655,N_4993);
nand U7089 (N_7089,N_4373,N_4148);
or U7090 (N_7090,N_2083,N_1234);
and U7091 (N_7091,N_4570,N_4237);
nor U7092 (N_7092,N_3291,N_570);
and U7093 (N_7093,N_247,N_2973);
and U7094 (N_7094,N_3481,N_3308);
xor U7095 (N_7095,N_1414,N_1906);
nand U7096 (N_7096,N_3711,N_3884);
or U7097 (N_7097,N_4191,N_2157);
xor U7098 (N_7098,N_3015,N_3473);
nand U7099 (N_7099,N_3106,N_3414);
xnor U7100 (N_7100,N_1370,N_4391);
or U7101 (N_7101,N_2975,N_1260);
and U7102 (N_7102,N_2389,N_3225);
and U7103 (N_7103,N_2557,N_4425);
and U7104 (N_7104,N_3218,N_2284);
nand U7105 (N_7105,N_2860,N_1928);
xor U7106 (N_7106,N_4503,N_3591);
xnor U7107 (N_7107,N_903,N_2934);
and U7108 (N_7108,N_2012,N_1063);
nor U7109 (N_7109,N_702,N_2716);
or U7110 (N_7110,N_4713,N_4594);
nor U7111 (N_7111,N_1488,N_787);
and U7112 (N_7112,N_2871,N_1422);
nand U7113 (N_7113,N_3847,N_3196);
nand U7114 (N_7114,N_3154,N_4860);
nor U7115 (N_7115,N_1092,N_134);
xnor U7116 (N_7116,N_692,N_4044);
and U7117 (N_7117,N_3328,N_4682);
nand U7118 (N_7118,N_1377,N_704);
and U7119 (N_7119,N_1265,N_764);
nor U7120 (N_7120,N_4792,N_1971);
and U7121 (N_7121,N_2476,N_2063);
xnor U7122 (N_7122,N_4256,N_3883);
or U7123 (N_7123,N_1645,N_4610);
nand U7124 (N_7124,N_4581,N_76);
or U7125 (N_7125,N_4328,N_1243);
and U7126 (N_7126,N_273,N_876);
nand U7127 (N_7127,N_2474,N_1387);
nor U7128 (N_7128,N_4685,N_1884);
xor U7129 (N_7129,N_2127,N_822);
or U7130 (N_7130,N_486,N_3329);
and U7131 (N_7131,N_3558,N_2597);
or U7132 (N_7132,N_829,N_1595);
nand U7133 (N_7133,N_339,N_4442);
and U7134 (N_7134,N_1911,N_1842);
and U7135 (N_7135,N_2795,N_4052);
or U7136 (N_7136,N_3581,N_2149);
or U7137 (N_7137,N_3536,N_3791);
nor U7138 (N_7138,N_1858,N_4252);
nand U7139 (N_7139,N_2834,N_4586);
nor U7140 (N_7140,N_4374,N_4695);
nand U7141 (N_7141,N_4639,N_1912);
xor U7142 (N_7142,N_1647,N_1991);
nor U7143 (N_7143,N_3047,N_1071);
or U7144 (N_7144,N_4564,N_988);
nor U7145 (N_7145,N_1773,N_4348);
or U7146 (N_7146,N_1978,N_902);
or U7147 (N_7147,N_3164,N_4747);
and U7148 (N_7148,N_918,N_1326);
or U7149 (N_7149,N_4336,N_2202);
nor U7150 (N_7150,N_137,N_1753);
nor U7151 (N_7151,N_3375,N_162);
nand U7152 (N_7152,N_3017,N_1443);
and U7153 (N_7153,N_3311,N_2909);
xor U7154 (N_7154,N_85,N_2239);
xor U7155 (N_7155,N_3805,N_844);
and U7156 (N_7156,N_1341,N_3523);
xnor U7157 (N_7157,N_3924,N_4899);
and U7158 (N_7158,N_3470,N_1686);
xnor U7159 (N_7159,N_4617,N_3084);
nand U7160 (N_7160,N_2242,N_3318);
or U7161 (N_7161,N_3808,N_2922);
xnor U7162 (N_7162,N_987,N_4843);
xor U7163 (N_7163,N_4119,N_1297);
nand U7164 (N_7164,N_2699,N_3212);
xnor U7165 (N_7165,N_4978,N_2472);
and U7166 (N_7166,N_2774,N_2507);
xnor U7167 (N_7167,N_2082,N_4627);
or U7168 (N_7168,N_1705,N_1609);
and U7169 (N_7169,N_736,N_3917);
nand U7170 (N_7170,N_481,N_1544);
and U7171 (N_7171,N_2359,N_1483);
and U7172 (N_7172,N_880,N_142);
and U7173 (N_7173,N_215,N_3119);
xnor U7174 (N_7174,N_346,N_3769);
nand U7175 (N_7175,N_3131,N_4181);
nand U7176 (N_7176,N_2056,N_3198);
xnor U7177 (N_7177,N_4651,N_3224);
xor U7178 (N_7178,N_4412,N_348);
xnor U7179 (N_7179,N_827,N_4521);
or U7180 (N_7180,N_4670,N_404);
nor U7181 (N_7181,N_3421,N_4658);
xnor U7182 (N_7182,N_1905,N_2504);
nor U7183 (N_7183,N_4008,N_3582);
xnor U7184 (N_7184,N_1085,N_2862);
and U7185 (N_7185,N_3664,N_4879);
nand U7186 (N_7186,N_2972,N_1577);
and U7187 (N_7187,N_2696,N_4318);
xor U7188 (N_7188,N_4195,N_2977);
or U7189 (N_7189,N_2544,N_3173);
xnor U7190 (N_7190,N_36,N_937);
or U7191 (N_7191,N_167,N_3697);
nand U7192 (N_7192,N_2594,N_4177);
and U7193 (N_7193,N_2432,N_2454);
nand U7194 (N_7194,N_4248,N_1558);
nand U7195 (N_7195,N_1976,N_3575);
nor U7196 (N_7196,N_4946,N_1484);
and U7197 (N_7197,N_328,N_643);
xor U7198 (N_7198,N_649,N_3044);
xnor U7199 (N_7199,N_506,N_178);
nand U7200 (N_7200,N_4243,N_3524);
or U7201 (N_7201,N_1425,N_957);
xor U7202 (N_7202,N_3176,N_3863);
nor U7203 (N_7203,N_424,N_4436);
or U7204 (N_7204,N_2920,N_1694);
or U7205 (N_7205,N_2334,N_3686);
or U7206 (N_7206,N_3532,N_2255);
and U7207 (N_7207,N_2510,N_4522);
xor U7208 (N_7208,N_4926,N_364);
or U7209 (N_7209,N_3182,N_3476);
or U7210 (N_7210,N_3638,N_4389);
nand U7211 (N_7211,N_3538,N_302);
nand U7212 (N_7212,N_4209,N_657);
and U7213 (N_7213,N_17,N_4217);
and U7214 (N_7214,N_16,N_4141);
or U7215 (N_7215,N_2653,N_4511);
nand U7216 (N_7216,N_2405,N_77);
and U7217 (N_7217,N_376,N_2226);
nand U7218 (N_7218,N_4010,N_318);
nor U7219 (N_7219,N_1123,N_3422);
and U7220 (N_7220,N_2537,N_3367);
or U7221 (N_7221,N_1638,N_4805);
nor U7222 (N_7222,N_3682,N_262);
nor U7223 (N_7223,N_4417,N_190);
and U7224 (N_7224,N_3179,N_807);
and U7225 (N_7225,N_574,N_1851);
xnor U7226 (N_7226,N_2407,N_2525);
nor U7227 (N_7227,N_2645,N_3077);
or U7228 (N_7228,N_3637,N_612);
nand U7229 (N_7229,N_3770,N_3721);
nand U7230 (N_7230,N_4478,N_1965);
or U7231 (N_7231,N_4047,N_201);
nor U7232 (N_7232,N_1489,N_260);
or U7233 (N_7233,N_2910,N_2123);
nand U7234 (N_7234,N_1409,N_2273);
nor U7235 (N_7235,N_4758,N_831);
nand U7236 (N_7236,N_2946,N_2288);
and U7237 (N_7237,N_4295,N_834);
xor U7238 (N_7238,N_4222,N_4890);
or U7239 (N_7239,N_1333,N_1219);
nor U7240 (N_7240,N_1561,N_4345);
and U7241 (N_7241,N_3075,N_4108);
and U7242 (N_7242,N_2666,N_1593);
or U7243 (N_7243,N_4183,N_2188);
xnor U7244 (N_7244,N_2154,N_817);
or U7245 (N_7245,N_731,N_3797);
nand U7246 (N_7246,N_289,N_2222);
nor U7247 (N_7247,N_1038,N_4483);
xnor U7248 (N_7248,N_4208,N_1835);
nand U7249 (N_7249,N_3998,N_1472);
and U7250 (N_7250,N_2759,N_2538);
or U7251 (N_7251,N_874,N_809);
nand U7252 (N_7252,N_4858,N_3995);
nor U7253 (N_7253,N_329,N_729);
or U7254 (N_7254,N_2304,N_3402);
and U7255 (N_7255,N_3619,N_4826);
and U7256 (N_7256,N_224,N_2181);
or U7257 (N_7257,N_4709,N_1406);
nor U7258 (N_7258,N_4894,N_1817);
nand U7259 (N_7259,N_4532,N_2237);
nor U7260 (N_7260,N_99,N_3425);
and U7261 (N_7261,N_3666,N_3598);
nand U7262 (N_7262,N_3678,N_4059);
nand U7263 (N_7263,N_4005,N_2165);
nor U7264 (N_7264,N_2049,N_3342);
nor U7265 (N_7265,N_2969,N_4870);
and U7266 (N_7266,N_3482,N_3724);
or U7267 (N_7267,N_2152,N_926);
or U7268 (N_7268,N_2697,N_1658);
xor U7269 (N_7269,N_2691,N_1924);
xnor U7270 (N_7270,N_2527,N_3259);
and U7271 (N_7271,N_3350,N_1255);
or U7272 (N_7272,N_3257,N_4749);
xnor U7273 (N_7273,N_311,N_604);
nand U7274 (N_7274,N_1916,N_4065);
and U7275 (N_7275,N_4698,N_4255);
and U7276 (N_7276,N_1482,N_1908);
xnor U7277 (N_7277,N_2384,N_309);
nand U7278 (N_7278,N_2295,N_2886);
nor U7279 (N_7279,N_1494,N_2686);
nand U7280 (N_7280,N_760,N_1815);
or U7281 (N_7281,N_2754,N_1336);
or U7282 (N_7282,N_3981,N_1490);
nor U7283 (N_7283,N_1610,N_1937);
xnor U7284 (N_7284,N_3222,N_972);
nor U7285 (N_7285,N_2727,N_1139);
nand U7286 (N_7286,N_756,N_954);
nor U7287 (N_7287,N_3234,N_485);
xnor U7288 (N_7288,N_4475,N_4355);
or U7289 (N_7289,N_2790,N_2013);
nand U7290 (N_7290,N_2349,N_3833);
nor U7291 (N_7291,N_2372,N_2751);
nor U7292 (N_7292,N_868,N_2416);
or U7293 (N_7293,N_1035,N_2532);
or U7294 (N_7294,N_3163,N_1583);
xor U7295 (N_7295,N_3086,N_1264);
nand U7296 (N_7296,N_4474,N_3901);
nand U7297 (N_7297,N_4744,N_2194);
nand U7298 (N_7298,N_777,N_3589);
and U7299 (N_7299,N_1382,N_724);
or U7300 (N_7300,N_1316,N_3374);
nand U7301 (N_7301,N_4636,N_607);
nor U7302 (N_7302,N_1401,N_1602);
nand U7303 (N_7303,N_1685,N_3814);
and U7304 (N_7304,N_1530,N_320);
and U7305 (N_7305,N_3128,N_3069);
or U7306 (N_7306,N_2668,N_4367);
nand U7307 (N_7307,N_2104,N_2358);
and U7308 (N_7308,N_3085,N_4133);
nor U7309 (N_7309,N_4989,N_1203);
or U7310 (N_7310,N_1437,N_836);
nor U7311 (N_7311,N_3184,N_4931);
xor U7312 (N_7312,N_3895,N_3307);
nand U7313 (N_7313,N_1836,N_2131);
nand U7314 (N_7314,N_3019,N_1824);
or U7315 (N_7315,N_3593,N_1720);
or U7316 (N_7316,N_331,N_3728);
xor U7317 (N_7317,N_4360,N_4440);
xnor U7318 (N_7318,N_3919,N_87);
xnor U7319 (N_7319,N_599,N_1278);
nor U7320 (N_7320,N_2260,N_4895);
nor U7321 (N_7321,N_2613,N_1112);
or U7322 (N_7322,N_4319,N_3094);
nor U7323 (N_7323,N_2511,N_4443);
nor U7324 (N_7324,N_2925,N_2087);
and U7325 (N_7325,N_466,N_1876);
xor U7326 (N_7326,N_4085,N_2138);
xor U7327 (N_7327,N_4330,N_4495);
nand U7328 (N_7328,N_4599,N_1627);
or U7329 (N_7329,N_935,N_1186);
nor U7330 (N_7330,N_2870,N_636);
xnor U7331 (N_7331,N_697,N_59);
nor U7332 (N_7332,N_216,N_3053);
xnor U7333 (N_7333,N_4880,N_627);
nor U7334 (N_7334,N_1478,N_4942);
nor U7335 (N_7335,N_2045,N_281);
and U7336 (N_7336,N_3480,N_2685);
and U7337 (N_7337,N_4925,N_213);
and U7338 (N_7338,N_102,N_721);
nor U7339 (N_7339,N_3067,N_940);
and U7340 (N_7340,N_1967,N_4724);
or U7341 (N_7341,N_989,N_650);
or U7342 (N_7342,N_1410,N_923);
nor U7343 (N_7343,N_1122,N_1365);
nand U7344 (N_7344,N_4873,N_3554);
xor U7345 (N_7345,N_3264,N_4664);
nor U7346 (N_7346,N_2518,N_2269);
xor U7347 (N_7347,N_3405,N_3160);
nand U7348 (N_7348,N_2221,N_4806);
nand U7349 (N_7349,N_2614,N_784);
or U7350 (N_7350,N_2960,N_4250);
xnor U7351 (N_7351,N_418,N_214);
nor U7352 (N_7352,N_3334,N_3855);
xor U7353 (N_7353,N_3468,N_699);
and U7354 (N_7354,N_1007,N_1133);
nor U7355 (N_7355,N_285,N_1104);
nor U7356 (N_7356,N_4774,N_2338);
or U7357 (N_7357,N_3874,N_2209);
nand U7358 (N_7358,N_4215,N_3809);
xnor U7359 (N_7359,N_4615,N_3842);
xnor U7360 (N_7360,N_2064,N_2015);
and U7361 (N_7361,N_3174,N_4110);
nand U7362 (N_7362,N_3622,N_4816);
and U7363 (N_7363,N_3112,N_452);
and U7364 (N_7364,N_1554,N_888);
and U7365 (N_7365,N_4194,N_4519);
or U7366 (N_7366,N_425,N_2039);
or U7367 (N_7367,N_2313,N_4053);
xnor U7368 (N_7368,N_480,N_1056);
xnor U7369 (N_7369,N_4992,N_3875);
nand U7370 (N_7370,N_4175,N_4479);
and U7371 (N_7371,N_0,N_3929);
or U7372 (N_7372,N_1157,N_3493);
nor U7373 (N_7373,N_4681,N_321);
xnor U7374 (N_7374,N_2299,N_1100);
and U7375 (N_7375,N_3036,N_3707);
or U7376 (N_7376,N_3691,N_1828);
nor U7377 (N_7377,N_3108,N_3477);
and U7378 (N_7378,N_3303,N_2676);
nor U7379 (N_7379,N_897,N_812);
nor U7380 (N_7380,N_4614,N_4049);
nor U7381 (N_7381,N_4887,N_4460);
nand U7382 (N_7382,N_1224,N_1477);
or U7383 (N_7383,N_1859,N_4757);
nor U7384 (N_7384,N_1655,N_2220);
or U7385 (N_7385,N_280,N_2758);
nand U7386 (N_7386,N_344,N_3659);
or U7387 (N_7387,N_195,N_3861);
xnor U7388 (N_7388,N_3366,N_966);
or U7389 (N_7389,N_383,N_1006);
nor U7390 (N_7390,N_4542,N_1535);
or U7391 (N_7391,N_1974,N_3887);
nor U7392 (N_7392,N_3368,N_2387);
nand U7393 (N_7393,N_624,N_3278);
or U7394 (N_7394,N_1288,N_2178);
and U7395 (N_7395,N_2412,N_4612);
nand U7396 (N_7396,N_1829,N_3486);
xor U7397 (N_7397,N_3658,N_3772);
or U7398 (N_7398,N_4772,N_984);
nor U7399 (N_7399,N_2767,N_2941);
nor U7400 (N_7400,N_435,N_2140);
nand U7401 (N_7401,N_3926,N_3910);
and U7402 (N_7402,N_3513,N_2499);
or U7403 (N_7403,N_2186,N_2845);
and U7404 (N_7404,N_2771,N_1719);
xor U7405 (N_7405,N_4924,N_3595);
or U7406 (N_7406,N_4868,N_4492);
nor U7407 (N_7407,N_147,N_4818);
and U7408 (N_7408,N_2341,N_4850);
nor U7409 (N_7409,N_2033,N_1837);
or U7410 (N_7410,N_2484,N_4971);
xor U7411 (N_7411,N_673,N_4464);
and U7412 (N_7412,N_2005,N_3650);
and U7413 (N_7413,N_1480,N_4745);
xnor U7414 (N_7414,N_1921,N_1683);
and U7415 (N_7415,N_1904,N_3567);
nand U7416 (N_7416,N_4637,N_4543);
and U7417 (N_7417,N_4694,N_2456);
or U7418 (N_7418,N_2414,N_198);
nor U7419 (N_7419,N_1356,N_2667);
nor U7420 (N_7420,N_2361,N_1821);
and U7421 (N_7421,N_1293,N_2434);
nand U7422 (N_7422,N_1515,N_1235);
nand U7423 (N_7423,N_4789,N_2672);
nor U7424 (N_7424,N_2360,N_357);
and U7425 (N_7425,N_2366,N_360);
and U7426 (N_7426,N_209,N_143);
and U7427 (N_7427,N_4036,N_4748);
and U7428 (N_7428,N_2736,N_3214);
or U7429 (N_7429,N_2539,N_762);
or U7430 (N_7430,N_3870,N_1199);
nand U7431 (N_7431,N_3474,N_2998);
nor U7432 (N_7432,N_3103,N_1191);
nand U7433 (N_7433,N_1861,N_108);
nand U7434 (N_7434,N_491,N_3511);
xnor U7435 (N_7435,N_3016,N_1972);
or U7436 (N_7436,N_1668,N_2163);
xor U7437 (N_7437,N_1737,N_1659);
nand U7438 (N_7438,N_4540,N_3960);
or U7439 (N_7439,N_2210,N_4656);
and U7440 (N_7440,N_2219,N_4577);
nor U7441 (N_7441,N_256,N_2447);
or U7442 (N_7442,N_734,N_482);
nand U7443 (N_7443,N_7,N_505);
and U7444 (N_7444,N_2678,N_3655);
nor U7445 (N_7445,N_2192,N_693);
xor U7446 (N_7446,N_1434,N_2211);
nand U7447 (N_7447,N_3980,N_3623);
and U7448 (N_7448,N_396,N_2944);
nor U7449 (N_7449,N_2084,N_2388);
or U7450 (N_7450,N_1709,N_2877);
nand U7451 (N_7451,N_4622,N_1778);
xor U7452 (N_7452,N_1024,N_3092);
and U7453 (N_7453,N_3026,N_3936);
nor U7454 (N_7454,N_4123,N_1587);
xor U7455 (N_7455,N_2731,N_3823);
nand U7456 (N_7456,N_2115,N_973);
and U7457 (N_7457,N_1624,N_1313);
nand U7458 (N_7458,N_3800,N_113);
nor U7459 (N_7459,N_3471,N_4002);
and U7460 (N_7460,N_4551,N_4344);
xnor U7461 (N_7461,N_261,N_4628);
nand U7462 (N_7462,N_1983,N_3243);
nor U7463 (N_7463,N_1128,N_2695);
nor U7464 (N_7464,N_1926,N_275);
xnor U7465 (N_7465,N_226,N_1960);
or U7466 (N_7466,N_1551,N_2885);
or U7467 (N_7467,N_3683,N_2878);
xor U7468 (N_7468,N_3720,N_342);
xor U7469 (N_7469,N_4734,N_2970);
or U7470 (N_7470,N_3273,N_4113);
or U7471 (N_7471,N_3965,N_3216);
or U7472 (N_7472,N_1346,N_4909);
or U7473 (N_7473,N_1789,N_31);
and U7474 (N_7474,N_1533,N_1634);
or U7475 (N_7475,N_3125,N_3152);
or U7476 (N_7476,N_2586,N_3269);
nor U7477 (N_7477,N_4186,N_4074);
or U7478 (N_7478,N_4225,N_4642);
nor U7479 (N_7479,N_4317,N_2390);
nor U7480 (N_7480,N_1347,N_3449);
nand U7481 (N_7481,N_757,N_4365);
nand U7482 (N_7482,N_3848,N_4161);
nor U7483 (N_7483,N_3751,N_4453);
xor U7484 (N_7484,N_4934,N_4439);
nand U7485 (N_7485,N_4882,N_3722);
nand U7486 (N_7486,N_934,N_1091);
xnor U7487 (N_7487,N_961,N_4151);
or U7488 (N_7488,N_4187,N_2494);
and U7489 (N_7489,N_939,N_3413);
xnor U7490 (N_7490,N_3976,N_358);
nor U7491 (N_7491,N_859,N_1381);
xor U7492 (N_7492,N_952,N_3906);
nor U7493 (N_7493,N_2704,N_4824);
or U7494 (N_7494,N_1094,N_3387);
nor U7495 (N_7495,N_3550,N_707);
xor U7496 (N_7496,N_2399,N_752);
xnor U7497 (N_7497,N_2918,N_3564);
and U7498 (N_7498,N_2347,N_3590);
nor U7499 (N_7499,N_1872,N_1013);
xnor U7500 (N_7500,N_4017,N_30);
nand U7501 (N_7501,N_2566,N_3857);
or U7502 (N_7502,N_180,N_4161);
and U7503 (N_7503,N_3781,N_2861);
and U7504 (N_7504,N_552,N_1455);
or U7505 (N_7505,N_3594,N_2531);
and U7506 (N_7506,N_230,N_4493);
xor U7507 (N_7507,N_1876,N_3406);
nor U7508 (N_7508,N_1609,N_366);
nand U7509 (N_7509,N_2653,N_679);
and U7510 (N_7510,N_2778,N_1994);
xnor U7511 (N_7511,N_4105,N_2873);
xnor U7512 (N_7512,N_2815,N_2621);
or U7513 (N_7513,N_649,N_580);
xnor U7514 (N_7514,N_3981,N_4127);
and U7515 (N_7515,N_1555,N_154);
or U7516 (N_7516,N_578,N_2470);
nand U7517 (N_7517,N_2392,N_2944);
or U7518 (N_7518,N_4995,N_184);
xnor U7519 (N_7519,N_2853,N_1775);
and U7520 (N_7520,N_4441,N_1518);
xor U7521 (N_7521,N_1860,N_3517);
xor U7522 (N_7522,N_3870,N_684);
or U7523 (N_7523,N_1811,N_4753);
xor U7524 (N_7524,N_2842,N_4091);
or U7525 (N_7525,N_3728,N_4420);
nand U7526 (N_7526,N_1499,N_2279);
or U7527 (N_7527,N_1565,N_4005);
xnor U7528 (N_7528,N_1562,N_851);
nand U7529 (N_7529,N_2037,N_3477);
or U7530 (N_7530,N_1927,N_1169);
nand U7531 (N_7531,N_1310,N_4183);
xnor U7532 (N_7532,N_3631,N_2337);
xor U7533 (N_7533,N_4627,N_4526);
nor U7534 (N_7534,N_364,N_4320);
xnor U7535 (N_7535,N_447,N_1440);
nor U7536 (N_7536,N_4767,N_1267);
xor U7537 (N_7537,N_1257,N_2837);
or U7538 (N_7538,N_1465,N_3344);
nor U7539 (N_7539,N_4871,N_2016);
nor U7540 (N_7540,N_73,N_2964);
or U7541 (N_7541,N_2211,N_1602);
and U7542 (N_7542,N_1609,N_1315);
or U7543 (N_7543,N_1392,N_1825);
nand U7544 (N_7544,N_547,N_731);
nand U7545 (N_7545,N_3102,N_1504);
or U7546 (N_7546,N_2466,N_4053);
nor U7547 (N_7547,N_2014,N_3125);
nand U7548 (N_7548,N_4706,N_741);
or U7549 (N_7549,N_4721,N_1071);
or U7550 (N_7550,N_1777,N_2798);
nor U7551 (N_7551,N_607,N_4816);
nor U7552 (N_7552,N_3822,N_3407);
xor U7553 (N_7553,N_643,N_1434);
nor U7554 (N_7554,N_4502,N_3943);
and U7555 (N_7555,N_1817,N_2821);
xor U7556 (N_7556,N_3054,N_799);
xor U7557 (N_7557,N_4750,N_2267);
or U7558 (N_7558,N_1595,N_2810);
nand U7559 (N_7559,N_3626,N_3579);
nand U7560 (N_7560,N_404,N_4216);
and U7561 (N_7561,N_1563,N_1628);
xor U7562 (N_7562,N_4644,N_4769);
nor U7563 (N_7563,N_4178,N_4785);
nor U7564 (N_7564,N_3930,N_4112);
xor U7565 (N_7565,N_2717,N_2697);
nand U7566 (N_7566,N_1690,N_2281);
nor U7567 (N_7567,N_1851,N_4200);
and U7568 (N_7568,N_4185,N_2341);
xnor U7569 (N_7569,N_403,N_0);
nor U7570 (N_7570,N_3491,N_363);
and U7571 (N_7571,N_351,N_2962);
or U7572 (N_7572,N_4586,N_3895);
nand U7573 (N_7573,N_1682,N_1048);
or U7574 (N_7574,N_1227,N_2314);
or U7575 (N_7575,N_4575,N_2749);
nand U7576 (N_7576,N_4400,N_3525);
nand U7577 (N_7577,N_2303,N_1272);
xnor U7578 (N_7578,N_1064,N_690);
and U7579 (N_7579,N_2477,N_2533);
and U7580 (N_7580,N_1880,N_1340);
xor U7581 (N_7581,N_2128,N_3144);
xnor U7582 (N_7582,N_695,N_4161);
or U7583 (N_7583,N_3999,N_2187);
and U7584 (N_7584,N_3948,N_726);
or U7585 (N_7585,N_4451,N_3672);
nor U7586 (N_7586,N_3973,N_848);
or U7587 (N_7587,N_2574,N_3081);
xor U7588 (N_7588,N_909,N_3304);
or U7589 (N_7589,N_4156,N_3784);
nand U7590 (N_7590,N_3159,N_2767);
nand U7591 (N_7591,N_3423,N_1497);
and U7592 (N_7592,N_1299,N_136);
nor U7593 (N_7593,N_1320,N_2841);
xnor U7594 (N_7594,N_2540,N_592);
nand U7595 (N_7595,N_3804,N_3096);
nor U7596 (N_7596,N_2083,N_4835);
and U7597 (N_7597,N_1542,N_3573);
xor U7598 (N_7598,N_518,N_4137);
nor U7599 (N_7599,N_1432,N_3089);
xor U7600 (N_7600,N_1076,N_1660);
xor U7601 (N_7601,N_1683,N_1117);
or U7602 (N_7602,N_2397,N_2523);
and U7603 (N_7603,N_560,N_513);
xor U7604 (N_7604,N_2508,N_4451);
nor U7605 (N_7605,N_1202,N_2016);
nor U7606 (N_7606,N_3248,N_1854);
nor U7607 (N_7607,N_1592,N_4414);
nor U7608 (N_7608,N_4698,N_3508);
nand U7609 (N_7609,N_1116,N_2908);
nand U7610 (N_7610,N_479,N_3933);
xor U7611 (N_7611,N_3773,N_1492);
xnor U7612 (N_7612,N_2251,N_1520);
or U7613 (N_7613,N_3647,N_34);
and U7614 (N_7614,N_1210,N_513);
and U7615 (N_7615,N_4056,N_96);
nor U7616 (N_7616,N_1834,N_3009);
or U7617 (N_7617,N_446,N_3027);
or U7618 (N_7618,N_2899,N_3163);
or U7619 (N_7619,N_215,N_3839);
xnor U7620 (N_7620,N_4030,N_1627);
nand U7621 (N_7621,N_4727,N_2335);
nor U7622 (N_7622,N_1665,N_4482);
xnor U7623 (N_7623,N_1426,N_3274);
nand U7624 (N_7624,N_4886,N_3871);
or U7625 (N_7625,N_2330,N_4807);
nor U7626 (N_7626,N_519,N_1915);
or U7627 (N_7627,N_546,N_2311);
xor U7628 (N_7628,N_4223,N_1542);
and U7629 (N_7629,N_4753,N_1972);
and U7630 (N_7630,N_1528,N_2254);
xor U7631 (N_7631,N_2124,N_3344);
xnor U7632 (N_7632,N_2777,N_4859);
and U7633 (N_7633,N_1756,N_4791);
xnor U7634 (N_7634,N_3126,N_3098);
nand U7635 (N_7635,N_2757,N_3681);
xor U7636 (N_7636,N_1945,N_3214);
nand U7637 (N_7637,N_4022,N_3272);
xor U7638 (N_7638,N_2746,N_1008);
nand U7639 (N_7639,N_701,N_2201);
nand U7640 (N_7640,N_3804,N_4105);
or U7641 (N_7641,N_3942,N_784);
nand U7642 (N_7642,N_303,N_990);
and U7643 (N_7643,N_4934,N_3787);
xor U7644 (N_7644,N_4934,N_2578);
or U7645 (N_7645,N_626,N_314);
nor U7646 (N_7646,N_856,N_2174);
and U7647 (N_7647,N_1687,N_2472);
and U7648 (N_7648,N_3146,N_4644);
nor U7649 (N_7649,N_1121,N_1539);
xnor U7650 (N_7650,N_4487,N_3046);
nand U7651 (N_7651,N_251,N_2569);
and U7652 (N_7652,N_451,N_991);
and U7653 (N_7653,N_2017,N_3096);
and U7654 (N_7654,N_3956,N_1569);
and U7655 (N_7655,N_3641,N_1014);
xnor U7656 (N_7656,N_857,N_525);
nor U7657 (N_7657,N_2165,N_215);
nand U7658 (N_7658,N_4218,N_1398);
and U7659 (N_7659,N_488,N_1234);
or U7660 (N_7660,N_4546,N_123);
or U7661 (N_7661,N_165,N_2925);
or U7662 (N_7662,N_189,N_277);
nor U7663 (N_7663,N_1781,N_2047);
xnor U7664 (N_7664,N_4214,N_1292);
and U7665 (N_7665,N_1193,N_4575);
nor U7666 (N_7666,N_2828,N_1993);
and U7667 (N_7667,N_1720,N_3786);
nor U7668 (N_7668,N_853,N_1474);
or U7669 (N_7669,N_4377,N_107);
nor U7670 (N_7670,N_2914,N_3245);
xor U7671 (N_7671,N_4812,N_2943);
xor U7672 (N_7672,N_862,N_1071);
nor U7673 (N_7673,N_4091,N_1781);
or U7674 (N_7674,N_4281,N_2951);
nor U7675 (N_7675,N_4458,N_2161);
xor U7676 (N_7676,N_4539,N_34);
xor U7677 (N_7677,N_654,N_4348);
nand U7678 (N_7678,N_70,N_2615);
or U7679 (N_7679,N_4264,N_2601);
nand U7680 (N_7680,N_3732,N_1887);
nor U7681 (N_7681,N_3291,N_855);
nor U7682 (N_7682,N_3498,N_1189);
nor U7683 (N_7683,N_502,N_759);
or U7684 (N_7684,N_1829,N_1329);
nand U7685 (N_7685,N_4798,N_2276);
xnor U7686 (N_7686,N_4301,N_2627);
or U7687 (N_7687,N_792,N_181);
xnor U7688 (N_7688,N_148,N_2642);
nand U7689 (N_7689,N_134,N_2116);
or U7690 (N_7690,N_3783,N_4040);
nand U7691 (N_7691,N_3475,N_4834);
or U7692 (N_7692,N_1001,N_816);
nor U7693 (N_7693,N_4869,N_921);
xor U7694 (N_7694,N_3976,N_2286);
nand U7695 (N_7695,N_3522,N_3294);
nand U7696 (N_7696,N_1707,N_4619);
nor U7697 (N_7697,N_498,N_913);
nand U7698 (N_7698,N_959,N_576);
and U7699 (N_7699,N_845,N_3827);
nand U7700 (N_7700,N_276,N_979);
nand U7701 (N_7701,N_2373,N_2969);
or U7702 (N_7702,N_4909,N_3006);
or U7703 (N_7703,N_3602,N_523);
or U7704 (N_7704,N_4939,N_2871);
nor U7705 (N_7705,N_1615,N_1430);
xnor U7706 (N_7706,N_657,N_2460);
xor U7707 (N_7707,N_3280,N_4133);
nand U7708 (N_7708,N_4226,N_1409);
nor U7709 (N_7709,N_2854,N_4166);
nand U7710 (N_7710,N_2590,N_3290);
or U7711 (N_7711,N_1871,N_2408);
or U7712 (N_7712,N_3748,N_4735);
and U7713 (N_7713,N_1248,N_415);
and U7714 (N_7714,N_3055,N_3153);
and U7715 (N_7715,N_4231,N_2058);
nand U7716 (N_7716,N_4080,N_4600);
or U7717 (N_7717,N_1218,N_1224);
or U7718 (N_7718,N_2221,N_2770);
nand U7719 (N_7719,N_2640,N_690);
or U7720 (N_7720,N_4377,N_4830);
or U7721 (N_7721,N_1396,N_1649);
and U7722 (N_7722,N_4471,N_57);
nand U7723 (N_7723,N_2170,N_3414);
nor U7724 (N_7724,N_899,N_4575);
or U7725 (N_7725,N_537,N_2330);
xor U7726 (N_7726,N_3344,N_1951);
nor U7727 (N_7727,N_2561,N_2182);
nand U7728 (N_7728,N_878,N_3857);
or U7729 (N_7729,N_1023,N_2334);
nor U7730 (N_7730,N_1351,N_1759);
nor U7731 (N_7731,N_400,N_3823);
or U7732 (N_7732,N_3410,N_4905);
nand U7733 (N_7733,N_1409,N_1810);
nor U7734 (N_7734,N_2521,N_1395);
or U7735 (N_7735,N_4436,N_1401);
nand U7736 (N_7736,N_3386,N_2432);
and U7737 (N_7737,N_3098,N_2046);
or U7738 (N_7738,N_987,N_4031);
nand U7739 (N_7739,N_4378,N_539);
nor U7740 (N_7740,N_2462,N_3695);
nand U7741 (N_7741,N_3651,N_3891);
nand U7742 (N_7742,N_719,N_3437);
xor U7743 (N_7743,N_1276,N_2549);
and U7744 (N_7744,N_1300,N_2186);
nand U7745 (N_7745,N_4617,N_1688);
and U7746 (N_7746,N_1980,N_723);
nor U7747 (N_7747,N_1852,N_4518);
and U7748 (N_7748,N_3223,N_4557);
nor U7749 (N_7749,N_523,N_4239);
and U7750 (N_7750,N_2324,N_1100);
or U7751 (N_7751,N_2441,N_1098);
and U7752 (N_7752,N_1317,N_13);
nand U7753 (N_7753,N_1040,N_3163);
xor U7754 (N_7754,N_4942,N_332);
nor U7755 (N_7755,N_4476,N_1932);
xor U7756 (N_7756,N_178,N_121);
and U7757 (N_7757,N_1307,N_670);
and U7758 (N_7758,N_421,N_245);
xnor U7759 (N_7759,N_1278,N_1173);
nand U7760 (N_7760,N_2271,N_529);
and U7761 (N_7761,N_1613,N_633);
nand U7762 (N_7762,N_683,N_647);
xnor U7763 (N_7763,N_275,N_2989);
and U7764 (N_7764,N_1812,N_2909);
nand U7765 (N_7765,N_2552,N_1959);
nor U7766 (N_7766,N_2586,N_1530);
and U7767 (N_7767,N_1355,N_2834);
or U7768 (N_7768,N_1500,N_128);
or U7769 (N_7769,N_4291,N_4540);
nor U7770 (N_7770,N_869,N_3429);
nand U7771 (N_7771,N_2173,N_2541);
or U7772 (N_7772,N_1412,N_4804);
or U7773 (N_7773,N_4553,N_4112);
xnor U7774 (N_7774,N_4797,N_3009);
or U7775 (N_7775,N_4703,N_3642);
or U7776 (N_7776,N_1534,N_2095);
or U7777 (N_7777,N_1696,N_3313);
nand U7778 (N_7778,N_1722,N_1079);
or U7779 (N_7779,N_1549,N_890);
nand U7780 (N_7780,N_3717,N_3849);
xor U7781 (N_7781,N_3623,N_2981);
xnor U7782 (N_7782,N_2975,N_3345);
xor U7783 (N_7783,N_3036,N_1967);
and U7784 (N_7784,N_4991,N_4116);
nor U7785 (N_7785,N_4795,N_4870);
and U7786 (N_7786,N_945,N_4370);
nand U7787 (N_7787,N_264,N_2920);
xor U7788 (N_7788,N_711,N_4221);
nor U7789 (N_7789,N_1228,N_4119);
or U7790 (N_7790,N_2249,N_4385);
nor U7791 (N_7791,N_244,N_3587);
and U7792 (N_7792,N_1744,N_2857);
xnor U7793 (N_7793,N_2756,N_4306);
nor U7794 (N_7794,N_4449,N_3550);
or U7795 (N_7795,N_374,N_3385);
nor U7796 (N_7796,N_2657,N_862);
nor U7797 (N_7797,N_260,N_119);
or U7798 (N_7798,N_4534,N_2667);
nand U7799 (N_7799,N_2835,N_3226);
xnor U7800 (N_7800,N_3826,N_4835);
nand U7801 (N_7801,N_1676,N_3789);
nor U7802 (N_7802,N_157,N_2768);
and U7803 (N_7803,N_2087,N_2509);
nor U7804 (N_7804,N_2609,N_1529);
and U7805 (N_7805,N_1510,N_4744);
or U7806 (N_7806,N_2778,N_1099);
nand U7807 (N_7807,N_1757,N_4446);
nor U7808 (N_7808,N_4268,N_3722);
or U7809 (N_7809,N_2439,N_200);
xor U7810 (N_7810,N_383,N_3226);
nor U7811 (N_7811,N_3816,N_2639);
and U7812 (N_7812,N_3903,N_1357);
or U7813 (N_7813,N_4764,N_4752);
xor U7814 (N_7814,N_4005,N_1749);
and U7815 (N_7815,N_766,N_1310);
and U7816 (N_7816,N_4913,N_1992);
or U7817 (N_7817,N_1349,N_2097);
nor U7818 (N_7818,N_4966,N_1857);
or U7819 (N_7819,N_4429,N_1412);
nor U7820 (N_7820,N_1704,N_3278);
and U7821 (N_7821,N_4118,N_358);
or U7822 (N_7822,N_538,N_1694);
nand U7823 (N_7823,N_4815,N_1779);
or U7824 (N_7824,N_2922,N_2158);
nand U7825 (N_7825,N_4666,N_4245);
xnor U7826 (N_7826,N_2420,N_4457);
and U7827 (N_7827,N_2928,N_1670);
and U7828 (N_7828,N_1213,N_1067);
or U7829 (N_7829,N_2188,N_1644);
or U7830 (N_7830,N_3227,N_1676);
nor U7831 (N_7831,N_381,N_1906);
nor U7832 (N_7832,N_775,N_2593);
or U7833 (N_7833,N_107,N_1540);
xnor U7834 (N_7834,N_1272,N_1804);
nand U7835 (N_7835,N_1377,N_2875);
nand U7836 (N_7836,N_4356,N_2336);
or U7837 (N_7837,N_2305,N_72);
or U7838 (N_7838,N_2064,N_3169);
nand U7839 (N_7839,N_419,N_1508);
nand U7840 (N_7840,N_2831,N_2810);
or U7841 (N_7841,N_3700,N_2836);
or U7842 (N_7842,N_4278,N_3097);
xnor U7843 (N_7843,N_1114,N_2619);
nor U7844 (N_7844,N_2480,N_1705);
nand U7845 (N_7845,N_108,N_1034);
xnor U7846 (N_7846,N_675,N_2497);
nor U7847 (N_7847,N_1571,N_2129);
nor U7848 (N_7848,N_1494,N_3771);
and U7849 (N_7849,N_252,N_2266);
and U7850 (N_7850,N_2982,N_3658);
or U7851 (N_7851,N_2497,N_325);
nor U7852 (N_7852,N_2063,N_3159);
and U7853 (N_7853,N_1098,N_4662);
and U7854 (N_7854,N_3777,N_1358);
and U7855 (N_7855,N_3444,N_2201);
xnor U7856 (N_7856,N_4954,N_3848);
nor U7857 (N_7857,N_2176,N_2622);
nand U7858 (N_7858,N_2951,N_39);
and U7859 (N_7859,N_1173,N_3616);
and U7860 (N_7860,N_893,N_4771);
nor U7861 (N_7861,N_4938,N_615);
xor U7862 (N_7862,N_149,N_1347);
nor U7863 (N_7863,N_222,N_1288);
xnor U7864 (N_7864,N_3245,N_2854);
nor U7865 (N_7865,N_1492,N_2743);
and U7866 (N_7866,N_4056,N_2038);
or U7867 (N_7867,N_479,N_1019);
or U7868 (N_7868,N_3788,N_2552);
or U7869 (N_7869,N_3938,N_3148);
or U7870 (N_7870,N_4511,N_592);
xor U7871 (N_7871,N_2060,N_4630);
and U7872 (N_7872,N_4036,N_3621);
and U7873 (N_7873,N_1547,N_3943);
and U7874 (N_7874,N_1791,N_1189);
nor U7875 (N_7875,N_3013,N_4900);
and U7876 (N_7876,N_4869,N_3024);
and U7877 (N_7877,N_801,N_3483);
or U7878 (N_7878,N_4293,N_162);
or U7879 (N_7879,N_990,N_2053);
nand U7880 (N_7880,N_3055,N_3388);
nor U7881 (N_7881,N_2606,N_3195);
xor U7882 (N_7882,N_1130,N_1810);
and U7883 (N_7883,N_1286,N_4013);
and U7884 (N_7884,N_4252,N_4007);
xnor U7885 (N_7885,N_1986,N_598);
nor U7886 (N_7886,N_595,N_2106);
xor U7887 (N_7887,N_2531,N_354);
and U7888 (N_7888,N_3923,N_1171);
or U7889 (N_7889,N_3712,N_4140);
and U7890 (N_7890,N_1306,N_3112);
nand U7891 (N_7891,N_4909,N_2969);
nand U7892 (N_7892,N_3179,N_2148);
and U7893 (N_7893,N_1135,N_4223);
nand U7894 (N_7894,N_2518,N_1705);
nor U7895 (N_7895,N_541,N_1110);
xnor U7896 (N_7896,N_1601,N_242);
or U7897 (N_7897,N_1616,N_2063);
or U7898 (N_7898,N_140,N_3388);
nand U7899 (N_7899,N_3075,N_3178);
and U7900 (N_7900,N_90,N_810);
xor U7901 (N_7901,N_4999,N_865);
xor U7902 (N_7902,N_1471,N_1062);
or U7903 (N_7903,N_568,N_332);
and U7904 (N_7904,N_3390,N_953);
xnor U7905 (N_7905,N_1190,N_316);
xor U7906 (N_7906,N_999,N_4453);
and U7907 (N_7907,N_4153,N_654);
or U7908 (N_7908,N_1004,N_3345);
nand U7909 (N_7909,N_1406,N_2031);
or U7910 (N_7910,N_2129,N_2489);
nand U7911 (N_7911,N_547,N_3235);
or U7912 (N_7912,N_4700,N_1641);
nor U7913 (N_7913,N_3196,N_2834);
and U7914 (N_7914,N_526,N_4226);
xor U7915 (N_7915,N_3186,N_2141);
and U7916 (N_7916,N_2783,N_4373);
or U7917 (N_7917,N_2355,N_3675);
nor U7918 (N_7918,N_1623,N_3643);
or U7919 (N_7919,N_1952,N_4273);
nand U7920 (N_7920,N_598,N_2426);
or U7921 (N_7921,N_165,N_3873);
or U7922 (N_7922,N_1990,N_1059);
xor U7923 (N_7923,N_3257,N_4450);
xnor U7924 (N_7924,N_232,N_1349);
xnor U7925 (N_7925,N_3723,N_4485);
nor U7926 (N_7926,N_4638,N_763);
nor U7927 (N_7927,N_38,N_4345);
xnor U7928 (N_7928,N_2227,N_2066);
nor U7929 (N_7929,N_92,N_4940);
nor U7930 (N_7930,N_1379,N_3205);
or U7931 (N_7931,N_4452,N_2385);
or U7932 (N_7932,N_4853,N_4314);
xnor U7933 (N_7933,N_3220,N_420);
or U7934 (N_7934,N_2423,N_3522);
and U7935 (N_7935,N_795,N_264);
and U7936 (N_7936,N_3089,N_2603);
or U7937 (N_7937,N_4091,N_3352);
nand U7938 (N_7938,N_1880,N_2240);
nand U7939 (N_7939,N_3375,N_3345);
nand U7940 (N_7940,N_4278,N_810);
or U7941 (N_7941,N_3938,N_3329);
and U7942 (N_7942,N_111,N_721);
xnor U7943 (N_7943,N_206,N_215);
xor U7944 (N_7944,N_2322,N_4148);
nand U7945 (N_7945,N_3102,N_1393);
or U7946 (N_7946,N_2072,N_4593);
or U7947 (N_7947,N_3368,N_3067);
nand U7948 (N_7948,N_144,N_676);
nand U7949 (N_7949,N_2590,N_1949);
or U7950 (N_7950,N_1908,N_2477);
or U7951 (N_7951,N_277,N_3094);
xnor U7952 (N_7952,N_2007,N_3628);
nor U7953 (N_7953,N_3466,N_3795);
or U7954 (N_7954,N_2913,N_3515);
or U7955 (N_7955,N_3490,N_3613);
and U7956 (N_7956,N_2203,N_554);
nor U7957 (N_7957,N_53,N_2825);
xor U7958 (N_7958,N_18,N_3286);
nand U7959 (N_7959,N_4365,N_1422);
xor U7960 (N_7960,N_410,N_2883);
nand U7961 (N_7961,N_1145,N_1260);
xor U7962 (N_7962,N_1511,N_1029);
xnor U7963 (N_7963,N_3371,N_4083);
and U7964 (N_7964,N_816,N_4852);
xor U7965 (N_7965,N_2578,N_4381);
nand U7966 (N_7966,N_3657,N_1500);
nand U7967 (N_7967,N_3113,N_3975);
and U7968 (N_7968,N_1100,N_2335);
nand U7969 (N_7969,N_4408,N_1305);
nor U7970 (N_7970,N_1972,N_3297);
xnor U7971 (N_7971,N_1841,N_2948);
and U7972 (N_7972,N_44,N_4046);
and U7973 (N_7973,N_1093,N_1389);
nor U7974 (N_7974,N_1502,N_59);
or U7975 (N_7975,N_1644,N_2687);
nor U7976 (N_7976,N_2092,N_3484);
nand U7977 (N_7977,N_2872,N_391);
or U7978 (N_7978,N_4045,N_3867);
xnor U7979 (N_7979,N_3554,N_904);
or U7980 (N_7980,N_4954,N_2544);
nor U7981 (N_7981,N_2198,N_3836);
nor U7982 (N_7982,N_2814,N_2799);
and U7983 (N_7983,N_3707,N_2978);
nor U7984 (N_7984,N_4759,N_1720);
xnor U7985 (N_7985,N_3520,N_4596);
and U7986 (N_7986,N_1430,N_2703);
and U7987 (N_7987,N_2635,N_949);
and U7988 (N_7988,N_2965,N_2871);
nand U7989 (N_7989,N_1455,N_2885);
nand U7990 (N_7990,N_3130,N_1954);
and U7991 (N_7991,N_3624,N_121);
and U7992 (N_7992,N_2038,N_3334);
xor U7993 (N_7993,N_3557,N_1486);
nand U7994 (N_7994,N_1965,N_4723);
nor U7995 (N_7995,N_1523,N_4210);
nor U7996 (N_7996,N_3033,N_4644);
and U7997 (N_7997,N_4924,N_1127);
xor U7998 (N_7998,N_421,N_2716);
or U7999 (N_7999,N_938,N_3600);
or U8000 (N_8000,N_540,N_1302);
nand U8001 (N_8001,N_2282,N_574);
nor U8002 (N_8002,N_4355,N_471);
and U8003 (N_8003,N_1255,N_4818);
nand U8004 (N_8004,N_4833,N_540);
nor U8005 (N_8005,N_252,N_2242);
or U8006 (N_8006,N_1040,N_1318);
or U8007 (N_8007,N_294,N_1335);
nand U8008 (N_8008,N_4205,N_142);
xnor U8009 (N_8009,N_2214,N_1938);
nand U8010 (N_8010,N_4053,N_4718);
nor U8011 (N_8011,N_2281,N_1075);
and U8012 (N_8012,N_4472,N_274);
and U8013 (N_8013,N_1075,N_4455);
nand U8014 (N_8014,N_4382,N_4732);
nand U8015 (N_8015,N_2986,N_1462);
and U8016 (N_8016,N_713,N_2091);
or U8017 (N_8017,N_3267,N_719);
nand U8018 (N_8018,N_1883,N_1683);
nor U8019 (N_8019,N_2617,N_3416);
nand U8020 (N_8020,N_2699,N_4357);
and U8021 (N_8021,N_3974,N_794);
nand U8022 (N_8022,N_1483,N_682);
or U8023 (N_8023,N_4165,N_3309);
xnor U8024 (N_8024,N_2900,N_1143);
nor U8025 (N_8025,N_2137,N_3675);
xor U8026 (N_8026,N_4604,N_725);
nand U8027 (N_8027,N_3150,N_2640);
or U8028 (N_8028,N_1437,N_2459);
nand U8029 (N_8029,N_1177,N_2931);
xnor U8030 (N_8030,N_1883,N_4497);
nand U8031 (N_8031,N_3066,N_3710);
and U8032 (N_8032,N_87,N_3679);
or U8033 (N_8033,N_198,N_730);
and U8034 (N_8034,N_818,N_4750);
and U8035 (N_8035,N_480,N_1986);
nand U8036 (N_8036,N_455,N_3722);
and U8037 (N_8037,N_3670,N_4547);
nor U8038 (N_8038,N_1110,N_1663);
or U8039 (N_8039,N_2348,N_3595);
xnor U8040 (N_8040,N_1576,N_2605);
xor U8041 (N_8041,N_3916,N_2091);
and U8042 (N_8042,N_3861,N_852);
or U8043 (N_8043,N_4455,N_2180);
and U8044 (N_8044,N_69,N_3360);
nor U8045 (N_8045,N_2553,N_4013);
nand U8046 (N_8046,N_2535,N_2964);
and U8047 (N_8047,N_209,N_1711);
nor U8048 (N_8048,N_4702,N_4017);
or U8049 (N_8049,N_3203,N_247);
and U8050 (N_8050,N_2975,N_4594);
xor U8051 (N_8051,N_3327,N_3139);
xnor U8052 (N_8052,N_1973,N_4459);
nor U8053 (N_8053,N_206,N_1645);
and U8054 (N_8054,N_21,N_4031);
xnor U8055 (N_8055,N_3988,N_4590);
nand U8056 (N_8056,N_4696,N_852);
nand U8057 (N_8057,N_2648,N_338);
and U8058 (N_8058,N_1436,N_2561);
nand U8059 (N_8059,N_398,N_2993);
xor U8060 (N_8060,N_3127,N_3658);
or U8061 (N_8061,N_1464,N_4833);
and U8062 (N_8062,N_1268,N_960);
xor U8063 (N_8063,N_2484,N_2888);
nand U8064 (N_8064,N_100,N_2658);
and U8065 (N_8065,N_1078,N_1256);
nor U8066 (N_8066,N_4285,N_1207);
nor U8067 (N_8067,N_3848,N_3349);
or U8068 (N_8068,N_2626,N_1075);
nor U8069 (N_8069,N_4709,N_1556);
nor U8070 (N_8070,N_72,N_1517);
nor U8071 (N_8071,N_4607,N_3103);
nor U8072 (N_8072,N_1664,N_2632);
xor U8073 (N_8073,N_1909,N_4055);
or U8074 (N_8074,N_4863,N_1553);
or U8075 (N_8075,N_2243,N_1904);
xnor U8076 (N_8076,N_546,N_292);
or U8077 (N_8077,N_3895,N_2102);
nand U8078 (N_8078,N_148,N_3070);
nor U8079 (N_8079,N_3786,N_269);
xnor U8080 (N_8080,N_1813,N_2245);
xor U8081 (N_8081,N_1202,N_4787);
xor U8082 (N_8082,N_3683,N_779);
nor U8083 (N_8083,N_515,N_399);
xor U8084 (N_8084,N_2349,N_2635);
and U8085 (N_8085,N_4602,N_1540);
nand U8086 (N_8086,N_1727,N_3574);
or U8087 (N_8087,N_4899,N_276);
and U8088 (N_8088,N_2501,N_3441);
or U8089 (N_8089,N_923,N_3247);
or U8090 (N_8090,N_2616,N_785);
or U8091 (N_8091,N_4744,N_4065);
and U8092 (N_8092,N_3296,N_4193);
xnor U8093 (N_8093,N_2821,N_3512);
and U8094 (N_8094,N_2185,N_3786);
or U8095 (N_8095,N_730,N_529);
nand U8096 (N_8096,N_4824,N_2782);
nand U8097 (N_8097,N_2403,N_164);
and U8098 (N_8098,N_223,N_4397);
xor U8099 (N_8099,N_2588,N_3395);
nor U8100 (N_8100,N_3526,N_2431);
and U8101 (N_8101,N_4336,N_4449);
and U8102 (N_8102,N_2937,N_407);
nor U8103 (N_8103,N_1364,N_3698);
and U8104 (N_8104,N_159,N_569);
or U8105 (N_8105,N_2683,N_4648);
or U8106 (N_8106,N_3237,N_1966);
and U8107 (N_8107,N_1045,N_4957);
and U8108 (N_8108,N_1606,N_2630);
nand U8109 (N_8109,N_1824,N_716);
nor U8110 (N_8110,N_3549,N_3534);
and U8111 (N_8111,N_2860,N_300);
or U8112 (N_8112,N_4696,N_3859);
and U8113 (N_8113,N_3840,N_2150);
nand U8114 (N_8114,N_3754,N_32);
xor U8115 (N_8115,N_4986,N_1603);
xnor U8116 (N_8116,N_4024,N_2701);
and U8117 (N_8117,N_2164,N_404);
nor U8118 (N_8118,N_1049,N_1159);
nor U8119 (N_8119,N_3672,N_4295);
nand U8120 (N_8120,N_4368,N_77);
and U8121 (N_8121,N_886,N_3531);
nor U8122 (N_8122,N_301,N_1233);
xnor U8123 (N_8123,N_2106,N_3011);
nor U8124 (N_8124,N_2044,N_4666);
or U8125 (N_8125,N_1951,N_2407);
nor U8126 (N_8126,N_4661,N_2472);
or U8127 (N_8127,N_1300,N_2686);
xnor U8128 (N_8128,N_2128,N_2618);
xor U8129 (N_8129,N_607,N_436);
nand U8130 (N_8130,N_2903,N_3015);
or U8131 (N_8131,N_3852,N_2304);
and U8132 (N_8132,N_811,N_1886);
or U8133 (N_8133,N_3546,N_755);
nor U8134 (N_8134,N_2524,N_4564);
nand U8135 (N_8135,N_162,N_342);
xor U8136 (N_8136,N_3375,N_3219);
nand U8137 (N_8137,N_3252,N_194);
nand U8138 (N_8138,N_4370,N_2672);
nand U8139 (N_8139,N_383,N_4190);
or U8140 (N_8140,N_2836,N_4498);
or U8141 (N_8141,N_2853,N_4711);
nand U8142 (N_8142,N_2434,N_4781);
nand U8143 (N_8143,N_1107,N_2109);
nand U8144 (N_8144,N_142,N_3958);
nand U8145 (N_8145,N_2436,N_3224);
and U8146 (N_8146,N_2493,N_436);
nor U8147 (N_8147,N_1611,N_1962);
or U8148 (N_8148,N_3605,N_3859);
and U8149 (N_8149,N_1203,N_746);
or U8150 (N_8150,N_4983,N_1016);
or U8151 (N_8151,N_4279,N_2525);
nand U8152 (N_8152,N_2486,N_1431);
nor U8153 (N_8153,N_1049,N_2381);
nand U8154 (N_8154,N_666,N_1496);
and U8155 (N_8155,N_1432,N_2917);
xnor U8156 (N_8156,N_822,N_2237);
nor U8157 (N_8157,N_122,N_3797);
or U8158 (N_8158,N_1919,N_998);
and U8159 (N_8159,N_2626,N_2240);
xnor U8160 (N_8160,N_2278,N_2743);
and U8161 (N_8161,N_1934,N_2280);
xnor U8162 (N_8162,N_1115,N_1490);
and U8163 (N_8163,N_3534,N_658);
nand U8164 (N_8164,N_227,N_1652);
and U8165 (N_8165,N_1452,N_3426);
nor U8166 (N_8166,N_581,N_4410);
xnor U8167 (N_8167,N_3384,N_2577);
xor U8168 (N_8168,N_683,N_4071);
nand U8169 (N_8169,N_4314,N_3887);
nand U8170 (N_8170,N_1230,N_4441);
and U8171 (N_8171,N_4032,N_1569);
and U8172 (N_8172,N_2346,N_1569);
nand U8173 (N_8173,N_2751,N_1295);
xnor U8174 (N_8174,N_4857,N_3797);
or U8175 (N_8175,N_4019,N_3598);
nor U8176 (N_8176,N_393,N_0);
nor U8177 (N_8177,N_2426,N_4773);
or U8178 (N_8178,N_3784,N_968);
nand U8179 (N_8179,N_1077,N_1598);
or U8180 (N_8180,N_1609,N_2740);
nor U8181 (N_8181,N_4576,N_1380);
or U8182 (N_8182,N_4725,N_3117);
xnor U8183 (N_8183,N_156,N_3362);
nand U8184 (N_8184,N_821,N_3604);
nand U8185 (N_8185,N_3497,N_2555);
and U8186 (N_8186,N_2383,N_4648);
and U8187 (N_8187,N_573,N_1577);
nand U8188 (N_8188,N_118,N_1342);
nor U8189 (N_8189,N_4896,N_140);
nor U8190 (N_8190,N_2726,N_2913);
nand U8191 (N_8191,N_2668,N_183);
xnor U8192 (N_8192,N_3415,N_4273);
or U8193 (N_8193,N_2389,N_2563);
and U8194 (N_8194,N_4282,N_1188);
xor U8195 (N_8195,N_4598,N_4167);
nand U8196 (N_8196,N_147,N_3145);
xor U8197 (N_8197,N_39,N_651);
nand U8198 (N_8198,N_852,N_3186);
nor U8199 (N_8199,N_3171,N_1234);
nand U8200 (N_8200,N_3492,N_1806);
and U8201 (N_8201,N_3522,N_2251);
and U8202 (N_8202,N_3837,N_2832);
nor U8203 (N_8203,N_2463,N_3788);
and U8204 (N_8204,N_1928,N_220);
or U8205 (N_8205,N_3030,N_4612);
nand U8206 (N_8206,N_3400,N_3232);
nand U8207 (N_8207,N_57,N_3989);
or U8208 (N_8208,N_968,N_4482);
and U8209 (N_8209,N_2612,N_2599);
and U8210 (N_8210,N_663,N_1004);
or U8211 (N_8211,N_1290,N_4856);
and U8212 (N_8212,N_4522,N_3134);
or U8213 (N_8213,N_3920,N_1116);
or U8214 (N_8214,N_1197,N_117);
and U8215 (N_8215,N_2096,N_1023);
nand U8216 (N_8216,N_2484,N_3683);
xor U8217 (N_8217,N_2864,N_1319);
and U8218 (N_8218,N_2120,N_3334);
nand U8219 (N_8219,N_3178,N_1220);
xor U8220 (N_8220,N_1462,N_318);
or U8221 (N_8221,N_4534,N_1477);
nand U8222 (N_8222,N_3942,N_3297);
nor U8223 (N_8223,N_2056,N_1701);
and U8224 (N_8224,N_1628,N_460);
and U8225 (N_8225,N_4501,N_4391);
or U8226 (N_8226,N_1288,N_4161);
nand U8227 (N_8227,N_2618,N_3162);
nand U8228 (N_8228,N_260,N_4010);
xor U8229 (N_8229,N_2240,N_4988);
nand U8230 (N_8230,N_1128,N_485);
xor U8231 (N_8231,N_2100,N_62);
nand U8232 (N_8232,N_3276,N_2436);
nand U8233 (N_8233,N_4722,N_3360);
xnor U8234 (N_8234,N_1775,N_1763);
or U8235 (N_8235,N_1673,N_2085);
and U8236 (N_8236,N_3540,N_731);
and U8237 (N_8237,N_4609,N_4729);
nand U8238 (N_8238,N_4609,N_2918);
or U8239 (N_8239,N_4976,N_3491);
xor U8240 (N_8240,N_536,N_3252);
or U8241 (N_8241,N_2679,N_3616);
or U8242 (N_8242,N_3255,N_4706);
nand U8243 (N_8243,N_1051,N_482);
and U8244 (N_8244,N_427,N_2911);
and U8245 (N_8245,N_4477,N_4992);
nor U8246 (N_8246,N_1069,N_1832);
xnor U8247 (N_8247,N_1857,N_324);
nor U8248 (N_8248,N_1873,N_525);
nand U8249 (N_8249,N_602,N_13);
nor U8250 (N_8250,N_4738,N_2950);
nor U8251 (N_8251,N_1635,N_1297);
and U8252 (N_8252,N_3787,N_4728);
xnor U8253 (N_8253,N_762,N_3883);
nand U8254 (N_8254,N_4565,N_3245);
nor U8255 (N_8255,N_567,N_4237);
xor U8256 (N_8256,N_4274,N_1805);
nand U8257 (N_8257,N_2949,N_4993);
nor U8258 (N_8258,N_1863,N_623);
or U8259 (N_8259,N_451,N_1299);
xnor U8260 (N_8260,N_1362,N_348);
or U8261 (N_8261,N_886,N_176);
nor U8262 (N_8262,N_2370,N_2575);
or U8263 (N_8263,N_4834,N_1558);
xnor U8264 (N_8264,N_2486,N_2746);
xor U8265 (N_8265,N_3288,N_4246);
xor U8266 (N_8266,N_4264,N_2852);
xnor U8267 (N_8267,N_1318,N_1152);
and U8268 (N_8268,N_3029,N_2951);
or U8269 (N_8269,N_3038,N_1100);
xor U8270 (N_8270,N_4064,N_917);
nor U8271 (N_8271,N_1620,N_4574);
nand U8272 (N_8272,N_3940,N_4412);
or U8273 (N_8273,N_1894,N_2624);
or U8274 (N_8274,N_3082,N_4555);
and U8275 (N_8275,N_58,N_2856);
and U8276 (N_8276,N_4366,N_2930);
or U8277 (N_8277,N_903,N_439);
xor U8278 (N_8278,N_4414,N_4385);
xor U8279 (N_8279,N_2264,N_730);
xnor U8280 (N_8280,N_1007,N_2492);
nand U8281 (N_8281,N_497,N_2082);
nand U8282 (N_8282,N_4033,N_4811);
xnor U8283 (N_8283,N_3346,N_3067);
xor U8284 (N_8284,N_4524,N_3067);
xnor U8285 (N_8285,N_756,N_1295);
nand U8286 (N_8286,N_756,N_4561);
nor U8287 (N_8287,N_1282,N_3153);
and U8288 (N_8288,N_2145,N_835);
nor U8289 (N_8289,N_160,N_1639);
xnor U8290 (N_8290,N_862,N_1792);
or U8291 (N_8291,N_488,N_1691);
and U8292 (N_8292,N_4101,N_3602);
and U8293 (N_8293,N_3722,N_1724);
nand U8294 (N_8294,N_2785,N_1572);
nand U8295 (N_8295,N_4476,N_3666);
nor U8296 (N_8296,N_1076,N_4361);
nor U8297 (N_8297,N_4123,N_3687);
nor U8298 (N_8298,N_1060,N_2359);
xnor U8299 (N_8299,N_4423,N_1488);
nand U8300 (N_8300,N_944,N_1503);
nor U8301 (N_8301,N_221,N_2945);
and U8302 (N_8302,N_143,N_67);
and U8303 (N_8303,N_1947,N_329);
xnor U8304 (N_8304,N_2414,N_3399);
and U8305 (N_8305,N_1178,N_4165);
or U8306 (N_8306,N_3306,N_1564);
nand U8307 (N_8307,N_2974,N_3751);
xor U8308 (N_8308,N_4973,N_4267);
xor U8309 (N_8309,N_3157,N_1009);
nand U8310 (N_8310,N_2750,N_3289);
and U8311 (N_8311,N_1947,N_534);
and U8312 (N_8312,N_4864,N_4849);
and U8313 (N_8313,N_3691,N_1129);
and U8314 (N_8314,N_2905,N_640);
xor U8315 (N_8315,N_1617,N_2763);
nor U8316 (N_8316,N_552,N_1883);
nand U8317 (N_8317,N_3015,N_3858);
xnor U8318 (N_8318,N_4791,N_4986);
or U8319 (N_8319,N_1890,N_2042);
and U8320 (N_8320,N_4421,N_1414);
xnor U8321 (N_8321,N_4757,N_1685);
nand U8322 (N_8322,N_2346,N_3385);
nand U8323 (N_8323,N_2652,N_3659);
xor U8324 (N_8324,N_3362,N_4492);
and U8325 (N_8325,N_2029,N_1846);
xnor U8326 (N_8326,N_1856,N_407);
or U8327 (N_8327,N_363,N_4709);
or U8328 (N_8328,N_2327,N_407);
and U8329 (N_8329,N_699,N_2593);
and U8330 (N_8330,N_710,N_2753);
nand U8331 (N_8331,N_283,N_720);
or U8332 (N_8332,N_2766,N_593);
or U8333 (N_8333,N_557,N_335);
nand U8334 (N_8334,N_364,N_4011);
or U8335 (N_8335,N_1178,N_1480);
and U8336 (N_8336,N_2584,N_172);
or U8337 (N_8337,N_913,N_4853);
nor U8338 (N_8338,N_2577,N_711);
or U8339 (N_8339,N_981,N_91);
and U8340 (N_8340,N_4064,N_164);
xor U8341 (N_8341,N_1073,N_1907);
nor U8342 (N_8342,N_2367,N_1044);
or U8343 (N_8343,N_1519,N_1969);
nor U8344 (N_8344,N_3299,N_4448);
nor U8345 (N_8345,N_2925,N_4710);
and U8346 (N_8346,N_2946,N_1292);
or U8347 (N_8347,N_4936,N_2997);
nand U8348 (N_8348,N_1360,N_1529);
and U8349 (N_8349,N_1833,N_1775);
nor U8350 (N_8350,N_663,N_815);
or U8351 (N_8351,N_3279,N_4399);
or U8352 (N_8352,N_3485,N_3924);
xnor U8353 (N_8353,N_3494,N_4048);
or U8354 (N_8354,N_2068,N_2652);
or U8355 (N_8355,N_3729,N_2226);
and U8356 (N_8356,N_2034,N_4266);
or U8357 (N_8357,N_53,N_1742);
nor U8358 (N_8358,N_3580,N_1126);
nor U8359 (N_8359,N_1996,N_2039);
and U8360 (N_8360,N_1784,N_2029);
or U8361 (N_8361,N_1503,N_2989);
nand U8362 (N_8362,N_4598,N_4998);
or U8363 (N_8363,N_2329,N_4320);
nor U8364 (N_8364,N_4306,N_319);
and U8365 (N_8365,N_943,N_2349);
nor U8366 (N_8366,N_228,N_1693);
xor U8367 (N_8367,N_2724,N_3615);
nor U8368 (N_8368,N_846,N_4483);
nand U8369 (N_8369,N_2290,N_2721);
xor U8370 (N_8370,N_4973,N_2058);
and U8371 (N_8371,N_2995,N_2603);
and U8372 (N_8372,N_382,N_819);
or U8373 (N_8373,N_2819,N_1155);
and U8374 (N_8374,N_3161,N_903);
xor U8375 (N_8375,N_3214,N_2802);
and U8376 (N_8376,N_208,N_3250);
nor U8377 (N_8377,N_1937,N_2586);
nand U8378 (N_8378,N_1562,N_1819);
and U8379 (N_8379,N_2237,N_840);
and U8380 (N_8380,N_4095,N_649);
nor U8381 (N_8381,N_521,N_986);
xor U8382 (N_8382,N_4408,N_4961);
or U8383 (N_8383,N_2508,N_3066);
or U8384 (N_8384,N_4836,N_4502);
or U8385 (N_8385,N_841,N_2145);
xnor U8386 (N_8386,N_4277,N_3460);
nor U8387 (N_8387,N_3134,N_4173);
and U8388 (N_8388,N_3149,N_1781);
xnor U8389 (N_8389,N_544,N_4903);
xor U8390 (N_8390,N_1077,N_1211);
nand U8391 (N_8391,N_4095,N_4900);
xnor U8392 (N_8392,N_1315,N_4010);
or U8393 (N_8393,N_1395,N_4622);
nand U8394 (N_8394,N_4628,N_1059);
nor U8395 (N_8395,N_3449,N_4025);
and U8396 (N_8396,N_1740,N_3620);
nor U8397 (N_8397,N_1386,N_409);
or U8398 (N_8398,N_1492,N_4261);
nand U8399 (N_8399,N_1894,N_2220);
nand U8400 (N_8400,N_3990,N_4705);
or U8401 (N_8401,N_1055,N_12);
nor U8402 (N_8402,N_1027,N_2923);
or U8403 (N_8403,N_684,N_1043);
xor U8404 (N_8404,N_4931,N_3082);
xor U8405 (N_8405,N_1472,N_4628);
xor U8406 (N_8406,N_2345,N_4861);
and U8407 (N_8407,N_2448,N_1988);
or U8408 (N_8408,N_1988,N_267);
and U8409 (N_8409,N_4861,N_1517);
or U8410 (N_8410,N_351,N_4778);
and U8411 (N_8411,N_952,N_4865);
or U8412 (N_8412,N_1875,N_3215);
nor U8413 (N_8413,N_4529,N_1277);
nand U8414 (N_8414,N_1148,N_4589);
nor U8415 (N_8415,N_166,N_3441);
and U8416 (N_8416,N_3387,N_164);
nor U8417 (N_8417,N_4044,N_1345);
and U8418 (N_8418,N_1251,N_450);
xor U8419 (N_8419,N_1634,N_3107);
xor U8420 (N_8420,N_4852,N_891);
nand U8421 (N_8421,N_3691,N_881);
nand U8422 (N_8422,N_3615,N_3623);
xor U8423 (N_8423,N_2988,N_3867);
xor U8424 (N_8424,N_3063,N_1765);
and U8425 (N_8425,N_2942,N_1263);
nor U8426 (N_8426,N_196,N_2663);
or U8427 (N_8427,N_1046,N_651);
and U8428 (N_8428,N_740,N_4637);
and U8429 (N_8429,N_1693,N_3683);
nand U8430 (N_8430,N_1597,N_1809);
xnor U8431 (N_8431,N_3656,N_2448);
nor U8432 (N_8432,N_623,N_1540);
nand U8433 (N_8433,N_3018,N_2554);
nor U8434 (N_8434,N_3544,N_947);
xnor U8435 (N_8435,N_4438,N_2303);
xor U8436 (N_8436,N_4600,N_2133);
nand U8437 (N_8437,N_3177,N_681);
xor U8438 (N_8438,N_762,N_3966);
and U8439 (N_8439,N_397,N_119);
and U8440 (N_8440,N_3810,N_886);
xnor U8441 (N_8441,N_3832,N_2610);
or U8442 (N_8442,N_320,N_2565);
or U8443 (N_8443,N_813,N_4935);
or U8444 (N_8444,N_1625,N_1172);
nor U8445 (N_8445,N_2338,N_2776);
nor U8446 (N_8446,N_523,N_4650);
nand U8447 (N_8447,N_3815,N_951);
or U8448 (N_8448,N_4410,N_4872);
xnor U8449 (N_8449,N_2034,N_3608);
nand U8450 (N_8450,N_511,N_4470);
and U8451 (N_8451,N_2941,N_4076);
or U8452 (N_8452,N_3238,N_4066);
nand U8453 (N_8453,N_2652,N_4996);
and U8454 (N_8454,N_3664,N_4930);
or U8455 (N_8455,N_3018,N_4064);
or U8456 (N_8456,N_4720,N_2248);
and U8457 (N_8457,N_174,N_777);
or U8458 (N_8458,N_4211,N_4218);
xor U8459 (N_8459,N_3710,N_4860);
nand U8460 (N_8460,N_1446,N_170);
nor U8461 (N_8461,N_1438,N_3671);
or U8462 (N_8462,N_1880,N_322);
or U8463 (N_8463,N_1058,N_1072);
and U8464 (N_8464,N_1717,N_3654);
and U8465 (N_8465,N_3069,N_341);
and U8466 (N_8466,N_872,N_2897);
xnor U8467 (N_8467,N_3046,N_3825);
nand U8468 (N_8468,N_1255,N_2800);
and U8469 (N_8469,N_2921,N_3074);
nand U8470 (N_8470,N_2745,N_1788);
nand U8471 (N_8471,N_960,N_785);
or U8472 (N_8472,N_1444,N_4025);
nand U8473 (N_8473,N_227,N_2938);
nand U8474 (N_8474,N_1876,N_3060);
or U8475 (N_8475,N_4424,N_1532);
xor U8476 (N_8476,N_1304,N_4082);
and U8477 (N_8477,N_635,N_1479);
nand U8478 (N_8478,N_1094,N_4321);
nand U8479 (N_8479,N_3251,N_4032);
xnor U8480 (N_8480,N_4292,N_2498);
xor U8481 (N_8481,N_798,N_659);
nand U8482 (N_8482,N_1386,N_4435);
nand U8483 (N_8483,N_478,N_3902);
xnor U8484 (N_8484,N_2640,N_986);
nor U8485 (N_8485,N_2878,N_488);
or U8486 (N_8486,N_4511,N_116);
and U8487 (N_8487,N_1766,N_3548);
xor U8488 (N_8488,N_1703,N_3733);
xnor U8489 (N_8489,N_3231,N_1853);
nand U8490 (N_8490,N_4426,N_1874);
or U8491 (N_8491,N_4842,N_1824);
nor U8492 (N_8492,N_3210,N_2838);
xor U8493 (N_8493,N_2563,N_4401);
nand U8494 (N_8494,N_806,N_1873);
xnor U8495 (N_8495,N_3443,N_3278);
and U8496 (N_8496,N_867,N_396);
xor U8497 (N_8497,N_3427,N_723);
nor U8498 (N_8498,N_1565,N_1309);
nor U8499 (N_8499,N_657,N_4605);
nor U8500 (N_8500,N_1851,N_3815);
xor U8501 (N_8501,N_1614,N_734);
and U8502 (N_8502,N_3424,N_2292);
xor U8503 (N_8503,N_2338,N_252);
nand U8504 (N_8504,N_3713,N_4448);
nand U8505 (N_8505,N_4908,N_1248);
and U8506 (N_8506,N_4485,N_276);
or U8507 (N_8507,N_1808,N_2325);
nor U8508 (N_8508,N_3347,N_1804);
and U8509 (N_8509,N_4464,N_4264);
and U8510 (N_8510,N_3379,N_4510);
xor U8511 (N_8511,N_1038,N_4631);
or U8512 (N_8512,N_3500,N_3170);
or U8513 (N_8513,N_4416,N_1471);
nor U8514 (N_8514,N_804,N_2437);
xnor U8515 (N_8515,N_4926,N_1762);
and U8516 (N_8516,N_2979,N_1334);
and U8517 (N_8517,N_1485,N_4454);
or U8518 (N_8518,N_4368,N_667);
or U8519 (N_8519,N_2842,N_119);
nor U8520 (N_8520,N_4346,N_1759);
nor U8521 (N_8521,N_2315,N_3586);
and U8522 (N_8522,N_3419,N_760);
xnor U8523 (N_8523,N_2922,N_399);
xnor U8524 (N_8524,N_3884,N_3188);
nor U8525 (N_8525,N_106,N_2996);
xnor U8526 (N_8526,N_1370,N_1091);
and U8527 (N_8527,N_3633,N_2413);
nor U8528 (N_8528,N_702,N_1051);
or U8529 (N_8529,N_2652,N_3306);
xnor U8530 (N_8530,N_784,N_2861);
nand U8531 (N_8531,N_3697,N_4346);
or U8532 (N_8532,N_3520,N_1778);
nor U8533 (N_8533,N_4324,N_129);
nand U8534 (N_8534,N_301,N_4257);
or U8535 (N_8535,N_3425,N_14);
nor U8536 (N_8536,N_2511,N_716);
or U8537 (N_8537,N_358,N_3636);
or U8538 (N_8538,N_4265,N_1929);
or U8539 (N_8539,N_4891,N_727);
and U8540 (N_8540,N_2006,N_1648);
nand U8541 (N_8541,N_131,N_1552);
nand U8542 (N_8542,N_3738,N_751);
xnor U8543 (N_8543,N_3937,N_1851);
or U8544 (N_8544,N_3852,N_1906);
nor U8545 (N_8545,N_3742,N_2709);
nand U8546 (N_8546,N_3468,N_681);
and U8547 (N_8547,N_2472,N_1175);
or U8548 (N_8548,N_4542,N_1960);
and U8549 (N_8549,N_998,N_3591);
xor U8550 (N_8550,N_4955,N_4761);
nor U8551 (N_8551,N_3201,N_4749);
nand U8552 (N_8552,N_3951,N_4432);
nor U8553 (N_8553,N_4790,N_2155);
xnor U8554 (N_8554,N_2129,N_3213);
and U8555 (N_8555,N_4128,N_169);
xor U8556 (N_8556,N_1942,N_4572);
and U8557 (N_8557,N_4026,N_399);
and U8558 (N_8558,N_3813,N_586);
or U8559 (N_8559,N_4317,N_212);
nand U8560 (N_8560,N_1466,N_4277);
and U8561 (N_8561,N_3296,N_4985);
or U8562 (N_8562,N_2045,N_883);
nor U8563 (N_8563,N_2969,N_2446);
nor U8564 (N_8564,N_3763,N_827);
xor U8565 (N_8565,N_4983,N_2143);
nor U8566 (N_8566,N_742,N_2498);
or U8567 (N_8567,N_169,N_1282);
and U8568 (N_8568,N_4258,N_4278);
nor U8569 (N_8569,N_2726,N_548);
nor U8570 (N_8570,N_4088,N_2652);
xnor U8571 (N_8571,N_4313,N_1944);
nor U8572 (N_8572,N_1965,N_4253);
nand U8573 (N_8573,N_972,N_868);
xor U8574 (N_8574,N_2608,N_3734);
and U8575 (N_8575,N_4400,N_1768);
and U8576 (N_8576,N_3666,N_834);
xnor U8577 (N_8577,N_3533,N_3066);
or U8578 (N_8578,N_3106,N_825);
nand U8579 (N_8579,N_1795,N_2412);
nand U8580 (N_8580,N_2286,N_105);
or U8581 (N_8581,N_1505,N_2512);
nor U8582 (N_8582,N_4082,N_3185);
and U8583 (N_8583,N_3833,N_299);
xnor U8584 (N_8584,N_3642,N_849);
or U8585 (N_8585,N_3691,N_4200);
xor U8586 (N_8586,N_1211,N_680);
nor U8587 (N_8587,N_229,N_2228);
nor U8588 (N_8588,N_1113,N_3778);
nand U8589 (N_8589,N_3913,N_2623);
nand U8590 (N_8590,N_4329,N_441);
xor U8591 (N_8591,N_458,N_361);
nor U8592 (N_8592,N_88,N_4179);
xor U8593 (N_8593,N_4723,N_1051);
xnor U8594 (N_8594,N_2273,N_1891);
nand U8595 (N_8595,N_3112,N_2273);
xnor U8596 (N_8596,N_1558,N_2013);
xor U8597 (N_8597,N_3415,N_2871);
and U8598 (N_8598,N_1429,N_4551);
or U8599 (N_8599,N_3835,N_783);
and U8600 (N_8600,N_4243,N_2565);
or U8601 (N_8601,N_357,N_789);
nand U8602 (N_8602,N_3602,N_4221);
xnor U8603 (N_8603,N_1861,N_3392);
nand U8604 (N_8604,N_591,N_3364);
nand U8605 (N_8605,N_680,N_4425);
nand U8606 (N_8606,N_4920,N_3105);
nand U8607 (N_8607,N_4067,N_948);
nor U8608 (N_8608,N_434,N_4524);
nand U8609 (N_8609,N_3364,N_4349);
or U8610 (N_8610,N_3181,N_3437);
nor U8611 (N_8611,N_3165,N_1475);
nor U8612 (N_8612,N_4887,N_2165);
xnor U8613 (N_8613,N_782,N_2258);
xor U8614 (N_8614,N_2132,N_4319);
nand U8615 (N_8615,N_4843,N_3195);
nor U8616 (N_8616,N_629,N_1263);
and U8617 (N_8617,N_1633,N_3227);
nor U8618 (N_8618,N_4799,N_2421);
or U8619 (N_8619,N_2677,N_1911);
or U8620 (N_8620,N_2646,N_3620);
nor U8621 (N_8621,N_1540,N_3318);
or U8622 (N_8622,N_1415,N_4611);
or U8623 (N_8623,N_4140,N_4596);
or U8624 (N_8624,N_1157,N_775);
and U8625 (N_8625,N_3367,N_3049);
nand U8626 (N_8626,N_1171,N_2569);
nor U8627 (N_8627,N_1122,N_323);
xor U8628 (N_8628,N_1990,N_4260);
nand U8629 (N_8629,N_4264,N_687);
nand U8630 (N_8630,N_2061,N_3096);
and U8631 (N_8631,N_2657,N_1277);
and U8632 (N_8632,N_690,N_4203);
nor U8633 (N_8633,N_2134,N_4803);
and U8634 (N_8634,N_2878,N_1165);
and U8635 (N_8635,N_4493,N_257);
xnor U8636 (N_8636,N_4577,N_4406);
and U8637 (N_8637,N_874,N_4555);
xnor U8638 (N_8638,N_1864,N_3482);
and U8639 (N_8639,N_1346,N_1673);
xnor U8640 (N_8640,N_4924,N_2274);
or U8641 (N_8641,N_248,N_2800);
nand U8642 (N_8642,N_3478,N_4745);
nor U8643 (N_8643,N_4892,N_3979);
and U8644 (N_8644,N_140,N_372);
nor U8645 (N_8645,N_3999,N_4337);
and U8646 (N_8646,N_291,N_1512);
nand U8647 (N_8647,N_2347,N_2771);
and U8648 (N_8648,N_1695,N_2967);
nand U8649 (N_8649,N_2058,N_3256);
or U8650 (N_8650,N_924,N_2574);
nand U8651 (N_8651,N_2916,N_4588);
xnor U8652 (N_8652,N_761,N_3177);
or U8653 (N_8653,N_4414,N_4361);
nand U8654 (N_8654,N_4159,N_1048);
or U8655 (N_8655,N_582,N_2707);
and U8656 (N_8656,N_4913,N_3892);
nand U8657 (N_8657,N_4107,N_3242);
xor U8658 (N_8658,N_489,N_2803);
nand U8659 (N_8659,N_2631,N_42);
and U8660 (N_8660,N_2946,N_4737);
and U8661 (N_8661,N_2333,N_794);
nor U8662 (N_8662,N_233,N_4885);
nor U8663 (N_8663,N_963,N_1364);
or U8664 (N_8664,N_2652,N_2617);
nand U8665 (N_8665,N_3963,N_252);
nor U8666 (N_8666,N_506,N_4962);
nand U8667 (N_8667,N_3944,N_1520);
or U8668 (N_8668,N_3274,N_4092);
and U8669 (N_8669,N_156,N_413);
or U8670 (N_8670,N_3677,N_1927);
nand U8671 (N_8671,N_1544,N_363);
nand U8672 (N_8672,N_3978,N_2552);
and U8673 (N_8673,N_1791,N_3252);
nor U8674 (N_8674,N_2802,N_3693);
xnor U8675 (N_8675,N_4421,N_4692);
nor U8676 (N_8676,N_1550,N_2207);
nand U8677 (N_8677,N_2983,N_349);
nand U8678 (N_8678,N_777,N_1147);
nand U8679 (N_8679,N_4597,N_573);
or U8680 (N_8680,N_2536,N_2775);
nor U8681 (N_8681,N_2548,N_3922);
or U8682 (N_8682,N_3417,N_4563);
nand U8683 (N_8683,N_4611,N_2613);
xnor U8684 (N_8684,N_2283,N_3455);
nand U8685 (N_8685,N_1857,N_1866);
and U8686 (N_8686,N_1830,N_1958);
xnor U8687 (N_8687,N_3178,N_3406);
nand U8688 (N_8688,N_2448,N_1399);
or U8689 (N_8689,N_3349,N_2439);
xor U8690 (N_8690,N_562,N_4828);
and U8691 (N_8691,N_4485,N_3787);
or U8692 (N_8692,N_1232,N_4426);
and U8693 (N_8693,N_4833,N_2674);
or U8694 (N_8694,N_4184,N_4775);
nor U8695 (N_8695,N_1818,N_3905);
nand U8696 (N_8696,N_1938,N_3734);
nor U8697 (N_8697,N_4153,N_438);
or U8698 (N_8698,N_976,N_2553);
and U8699 (N_8699,N_152,N_3163);
nor U8700 (N_8700,N_1495,N_2641);
xnor U8701 (N_8701,N_3247,N_509);
nor U8702 (N_8702,N_1534,N_1851);
and U8703 (N_8703,N_1392,N_401);
nand U8704 (N_8704,N_2524,N_2402);
xor U8705 (N_8705,N_1914,N_376);
nand U8706 (N_8706,N_3496,N_3584);
nor U8707 (N_8707,N_522,N_3231);
and U8708 (N_8708,N_4571,N_2177);
xnor U8709 (N_8709,N_2609,N_2581);
xnor U8710 (N_8710,N_2663,N_267);
xor U8711 (N_8711,N_1697,N_2140);
or U8712 (N_8712,N_3681,N_2737);
xor U8713 (N_8713,N_2028,N_2176);
or U8714 (N_8714,N_3401,N_1176);
or U8715 (N_8715,N_4410,N_3546);
nor U8716 (N_8716,N_3946,N_859);
nor U8717 (N_8717,N_742,N_2876);
or U8718 (N_8718,N_2975,N_2588);
or U8719 (N_8719,N_1510,N_4166);
or U8720 (N_8720,N_518,N_744);
xnor U8721 (N_8721,N_4154,N_1656);
and U8722 (N_8722,N_693,N_748);
or U8723 (N_8723,N_421,N_2651);
and U8724 (N_8724,N_896,N_828);
nor U8725 (N_8725,N_2267,N_3741);
or U8726 (N_8726,N_2212,N_2809);
xor U8727 (N_8727,N_2839,N_839);
nand U8728 (N_8728,N_3693,N_501);
xor U8729 (N_8729,N_2816,N_1506);
nor U8730 (N_8730,N_125,N_1850);
nor U8731 (N_8731,N_3205,N_4774);
or U8732 (N_8732,N_4422,N_792);
nor U8733 (N_8733,N_3343,N_4114);
or U8734 (N_8734,N_2006,N_4073);
nand U8735 (N_8735,N_419,N_416);
nand U8736 (N_8736,N_267,N_2200);
and U8737 (N_8737,N_482,N_656);
xor U8738 (N_8738,N_442,N_673);
nand U8739 (N_8739,N_2586,N_3668);
nor U8740 (N_8740,N_1806,N_180);
nor U8741 (N_8741,N_3987,N_2781);
xor U8742 (N_8742,N_4681,N_4028);
nor U8743 (N_8743,N_3876,N_4980);
nor U8744 (N_8744,N_2218,N_880);
and U8745 (N_8745,N_1331,N_2797);
xor U8746 (N_8746,N_4529,N_1234);
nor U8747 (N_8747,N_4109,N_1087);
nor U8748 (N_8748,N_4256,N_4217);
nand U8749 (N_8749,N_3442,N_1295);
and U8750 (N_8750,N_1661,N_4023);
nand U8751 (N_8751,N_4960,N_4996);
or U8752 (N_8752,N_1274,N_179);
xor U8753 (N_8753,N_979,N_3652);
xnor U8754 (N_8754,N_4442,N_326);
or U8755 (N_8755,N_635,N_3057);
xor U8756 (N_8756,N_542,N_2807);
xnor U8757 (N_8757,N_1207,N_1186);
nand U8758 (N_8758,N_3409,N_3958);
xnor U8759 (N_8759,N_1568,N_251);
nand U8760 (N_8760,N_1938,N_3494);
nor U8761 (N_8761,N_4169,N_3979);
nand U8762 (N_8762,N_140,N_1843);
nand U8763 (N_8763,N_1555,N_3525);
nand U8764 (N_8764,N_3026,N_1388);
nand U8765 (N_8765,N_733,N_1072);
and U8766 (N_8766,N_69,N_4753);
nand U8767 (N_8767,N_2582,N_117);
and U8768 (N_8768,N_1566,N_101);
nor U8769 (N_8769,N_1747,N_780);
nor U8770 (N_8770,N_1332,N_4051);
nor U8771 (N_8771,N_2820,N_4150);
nand U8772 (N_8772,N_1629,N_3815);
and U8773 (N_8773,N_4859,N_1861);
or U8774 (N_8774,N_4580,N_3701);
and U8775 (N_8775,N_4089,N_1991);
and U8776 (N_8776,N_2803,N_2722);
and U8777 (N_8777,N_4873,N_1234);
and U8778 (N_8778,N_2813,N_3856);
nand U8779 (N_8779,N_3783,N_419);
nor U8780 (N_8780,N_2632,N_167);
nand U8781 (N_8781,N_2458,N_1056);
and U8782 (N_8782,N_21,N_4122);
nor U8783 (N_8783,N_1316,N_4738);
and U8784 (N_8784,N_1622,N_4704);
xnor U8785 (N_8785,N_1448,N_4035);
or U8786 (N_8786,N_1443,N_2782);
and U8787 (N_8787,N_3287,N_4709);
or U8788 (N_8788,N_2680,N_664);
nor U8789 (N_8789,N_3801,N_3737);
xor U8790 (N_8790,N_39,N_2718);
or U8791 (N_8791,N_1818,N_2528);
and U8792 (N_8792,N_1624,N_2002);
xnor U8793 (N_8793,N_2167,N_4390);
or U8794 (N_8794,N_335,N_2065);
xor U8795 (N_8795,N_2240,N_4385);
xnor U8796 (N_8796,N_1218,N_3519);
or U8797 (N_8797,N_2770,N_3247);
nand U8798 (N_8798,N_2189,N_386);
nand U8799 (N_8799,N_2106,N_1460);
nand U8800 (N_8800,N_534,N_3752);
nand U8801 (N_8801,N_3263,N_3232);
nand U8802 (N_8802,N_3857,N_2551);
or U8803 (N_8803,N_389,N_450);
xnor U8804 (N_8804,N_4175,N_4067);
nand U8805 (N_8805,N_4148,N_2303);
nand U8806 (N_8806,N_4333,N_3808);
and U8807 (N_8807,N_3705,N_3156);
or U8808 (N_8808,N_19,N_1716);
or U8809 (N_8809,N_4738,N_834);
nand U8810 (N_8810,N_4898,N_233);
xnor U8811 (N_8811,N_835,N_1033);
nor U8812 (N_8812,N_2347,N_3695);
nor U8813 (N_8813,N_95,N_559);
nor U8814 (N_8814,N_716,N_1553);
nand U8815 (N_8815,N_3495,N_4234);
or U8816 (N_8816,N_3429,N_4062);
or U8817 (N_8817,N_4052,N_25);
nand U8818 (N_8818,N_2023,N_4856);
nand U8819 (N_8819,N_4281,N_4710);
or U8820 (N_8820,N_999,N_1305);
nand U8821 (N_8821,N_4580,N_2976);
or U8822 (N_8822,N_2592,N_3767);
nand U8823 (N_8823,N_3100,N_2741);
or U8824 (N_8824,N_179,N_2725);
and U8825 (N_8825,N_4171,N_3160);
or U8826 (N_8826,N_498,N_4489);
and U8827 (N_8827,N_2641,N_3633);
xor U8828 (N_8828,N_335,N_3241);
nor U8829 (N_8829,N_1020,N_4743);
nand U8830 (N_8830,N_2133,N_1502);
or U8831 (N_8831,N_1661,N_4760);
or U8832 (N_8832,N_2884,N_4096);
and U8833 (N_8833,N_4529,N_3840);
nand U8834 (N_8834,N_2405,N_3154);
nor U8835 (N_8835,N_212,N_256);
xor U8836 (N_8836,N_1654,N_1308);
and U8837 (N_8837,N_1837,N_2741);
xnor U8838 (N_8838,N_1105,N_1527);
xor U8839 (N_8839,N_4012,N_1745);
nor U8840 (N_8840,N_1059,N_2964);
or U8841 (N_8841,N_3408,N_4266);
nand U8842 (N_8842,N_4598,N_1110);
and U8843 (N_8843,N_3556,N_2829);
or U8844 (N_8844,N_2970,N_1495);
nor U8845 (N_8845,N_3118,N_4826);
and U8846 (N_8846,N_261,N_1601);
nand U8847 (N_8847,N_303,N_1138);
nor U8848 (N_8848,N_334,N_1260);
and U8849 (N_8849,N_3153,N_1332);
and U8850 (N_8850,N_4348,N_2809);
nand U8851 (N_8851,N_2510,N_3557);
nand U8852 (N_8852,N_712,N_3221);
nand U8853 (N_8853,N_367,N_3672);
or U8854 (N_8854,N_2392,N_2698);
or U8855 (N_8855,N_2578,N_1805);
and U8856 (N_8856,N_566,N_2717);
nor U8857 (N_8857,N_4652,N_2609);
and U8858 (N_8858,N_2316,N_1635);
and U8859 (N_8859,N_2717,N_448);
or U8860 (N_8860,N_436,N_2648);
and U8861 (N_8861,N_1997,N_4224);
xnor U8862 (N_8862,N_2479,N_2050);
xnor U8863 (N_8863,N_439,N_3466);
nor U8864 (N_8864,N_3633,N_2127);
nor U8865 (N_8865,N_3837,N_4065);
xor U8866 (N_8866,N_2408,N_1988);
and U8867 (N_8867,N_767,N_1535);
xor U8868 (N_8868,N_1569,N_1404);
xor U8869 (N_8869,N_525,N_4157);
xor U8870 (N_8870,N_4338,N_2866);
nand U8871 (N_8871,N_3180,N_3462);
xor U8872 (N_8872,N_3909,N_4693);
nor U8873 (N_8873,N_1180,N_1072);
and U8874 (N_8874,N_4053,N_227);
or U8875 (N_8875,N_3528,N_2642);
nor U8876 (N_8876,N_352,N_3986);
nor U8877 (N_8877,N_3736,N_2508);
and U8878 (N_8878,N_2698,N_1043);
nand U8879 (N_8879,N_464,N_534);
nor U8880 (N_8880,N_1874,N_615);
nor U8881 (N_8881,N_1185,N_4922);
and U8882 (N_8882,N_3262,N_557);
xnor U8883 (N_8883,N_394,N_1907);
or U8884 (N_8884,N_4908,N_4237);
or U8885 (N_8885,N_1201,N_2511);
nor U8886 (N_8886,N_1994,N_3116);
and U8887 (N_8887,N_514,N_3857);
and U8888 (N_8888,N_1607,N_1935);
nand U8889 (N_8889,N_432,N_2484);
nor U8890 (N_8890,N_1257,N_3009);
xor U8891 (N_8891,N_2406,N_3677);
nand U8892 (N_8892,N_179,N_278);
nor U8893 (N_8893,N_2307,N_1600);
and U8894 (N_8894,N_4996,N_4973);
xor U8895 (N_8895,N_1338,N_4095);
nor U8896 (N_8896,N_4386,N_4174);
or U8897 (N_8897,N_2002,N_1900);
nor U8898 (N_8898,N_1657,N_1432);
or U8899 (N_8899,N_288,N_4728);
or U8900 (N_8900,N_1065,N_1746);
xor U8901 (N_8901,N_3658,N_4405);
nand U8902 (N_8902,N_3680,N_2162);
xor U8903 (N_8903,N_2123,N_3952);
nor U8904 (N_8904,N_350,N_218);
xor U8905 (N_8905,N_4839,N_1641);
xor U8906 (N_8906,N_3670,N_1363);
nor U8907 (N_8907,N_3347,N_717);
xor U8908 (N_8908,N_1456,N_306);
nand U8909 (N_8909,N_2016,N_2791);
and U8910 (N_8910,N_1868,N_2812);
or U8911 (N_8911,N_4156,N_3657);
or U8912 (N_8912,N_1300,N_3482);
nand U8913 (N_8913,N_2968,N_464);
nand U8914 (N_8914,N_4326,N_200);
nor U8915 (N_8915,N_939,N_2107);
xnor U8916 (N_8916,N_4222,N_1747);
nor U8917 (N_8917,N_1745,N_3985);
nor U8918 (N_8918,N_2142,N_2285);
nand U8919 (N_8919,N_3329,N_1074);
or U8920 (N_8920,N_2961,N_830);
xor U8921 (N_8921,N_4800,N_1977);
nor U8922 (N_8922,N_4845,N_1018);
or U8923 (N_8923,N_3275,N_4385);
nand U8924 (N_8924,N_18,N_4574);
nor U8925 (N_8925,N_4051,N_1520);
nor U8926 (N_8926,N_3499,N_406);
or U8927 (N_8927,N_1821,N_74);
nor U8928 (N_8928,N_2667,N_260);
nor U8929 (N_8929,N_771,N_2157);
xnor U8930 (N_8930,N_399,N_1546);
xnor U8931 (N_8931,N_3434,N_1970);
nor U8932 (N_8932,N_4916,N_1043);
xor U8933 (N_8933,N_4215,N_744);
and U8934 (N_8934,N_3717,N_235);
xor U8935 (N_8935,N_4371,N_241);
nand U8936 (N_8936,N_4082,N_3615);
nand U8937 (N_8937,N_4799,N_4626);
nor U8938 (N_8938,N_3790,N_541);
nand U8939 (N_8939,N_893,N_2028);
or U8940 (N_8940,N_1442,N_3547);
and U8941 (N_8941,N_3306,N_1809);
or U8942 (N_8942,N_3175,N_1707);
nand U8943 (N_8943,N_4083,N_4283);
nor U8944 (N_8944,N_1758,N_4694);
nand U8945 (N_8945,N_1139,N_4362);
and U8946 (N_8946,N_4656,N_1283);
and U8947 (N_8947,N_2323,N_2929);
and U8948 (N_8948,N_869,N_3425);
nor U8949 (N_8949,N_3642,N_4692);
nor U8950 (N_8950,N_3136,N_4598);
xnor U8951 (N_8951,N_3515,N_3159);
xnor U8952 (N_8952,N_1833,N_2430);
and U8953 (N_8953,N_4234,N_3122);
nor U8954 (N_8954,N_3257,N_3862);
or U8955 (N_8955,N_2864,N_908);
and U8956 (N_8956,N_1951,N_2969);
and U8957 (N_8957,N_2391,N_4716);
nor U8958 (N_8958,N_631,N_2456);
and U8959 (N_8959,N_1465,N_75);
or U8960 (N_8960,N_111,N_1385);
xor U8961 (N_8961,N_2523,N_1910);
and U8962 (N_8962,N_3500,N_3295);
nand U8963 (N_8963,N_3157,N_3457);
xor U8964 (N_8964,N_1112,N_1360);
or U8965 (N_8965,N_1580,N_1785);
or U8966 (N_8966,N_1266,N_2335);
xnor U8967 (N_8967,N_466,N_1635);
nor U8968 (N_8968,N_2841,N_2704);
xor U8969 (N_8969,N_3880,N_3849);
and U8970 (N_8970,N_2273,N_326);
nand U8971 (N_8971,N_2468,N_3866);
nor U8972 (N_8972,N_4628,N_3511);
xnor U8973 (N_8973,N_4741,N_4260);
nand U8974 (N_8974,N_3702,N_2515);
or U8975 (N_8975,N_4377,N_3353);
nor U8976 (N_8976,N_1643,N_4783);
xnor U8977 (N_8977,N_2125,N_4275);
nor U8978 (N_8978,N_4676,N_3630);
nand U8979 (N_8979,N_960,N_2767);
or U8980 (N_8980,N_4675,N_223);
nand U8981 (N_8981,N_793,N_3228);
or U8982 (N_8982,N_804,N_1388);
nand U8983 (N_8983,N_2538,N_3667);
or U8984 (N_8984,N_3499,N_2808);
and U8985 (N_8985,N_3769,N_3921);
and U8986 (N_8986,N_1022,N_2929);
xnor U8987 (N_8987,N_933,N_3188);
and U8988 (N_8988,N_4842,N_1767);
xnor U8989 (N_8989,N_3097,N_2845);
or U8990 (N_8990,N_1619,N_4305);
xnor U8991 (N_8991,N_2886,N_2435);
or U8992 (N_8992,N_4077,N_3171);
xnor U8993 (N_8993,N_417,N_2366);
nand U8994 (N_8994,N_688,N_3902);
or U8995 (N_8995,N_3958,N_3446);
nor U8996 (N_8996,N_3959,N_3916);
nand U8997 (N_8997,N_604,N_3838);
xor U8998 (N_8998,N_1743,N_2847);
and U8999 (N_8999,N_1552,N_3417);
and U9000 (N_9000,N_4706,N_3994);
and U9001 (N_9001,N_1135,N_4479);
and U9002 (N_9002,N_742,N_782);
nor U9003 (N_9003,N_755,N_2878);
or U9004 (N_9004,N_4750,N_4140);
nand U9005 (N_9005,N_634,N_1960);
and U9006 (N_9006,N_895,N_4751);
or U9007 (N_9007,N_4906,N_4648);
and U9008 (N_9008,N_844,N_2649);
nand U9009 (N_9009,N_4008,N_3792);
nor U9010 (N_9010,N_4866,N_1613);
nor U9011 (N_9011,N_1348,N_774);
or U9012 (N_9012,N_1282,N_2963);
or U9013 (N_9013,N_884,N_3922);
nand U9014 (N_9014,N_723,N_374);
nor U9015 (N_9015,N_2583,N_4754);
nand U9016 (N_9016,N_2616,N_3747);
nand U9017 (N_9017,N_3573,N_4160);
nand U9018 (N_9018,N_1277,N_4419);
or U9019 (N_9019,N_1763,N_4458);
or U9020 (N_9020,N_4368,N_1039);
or U9021 (N_9021,N_3594,N_906);
xor U9022 (N_9022,N_4821,N_2894);
xnor U9023 (N_9023,N_2837,N_3546);
nand U9024 (N_9024,N_609,N_2304);
or U9025 (N_9025,N_1275,N_3238);
nand U9026 (N_9026,N_2458,N_1241);
and U9027 (N_9027,N_2105,N_4252);
and U9028 (N_9028,N_1835,N_4374);
nor U9029 (N_9029,N_4575,N_3538);
nand U9030 (N_9030,N_2578,N_4704);
nand U9031 (N_9031,N_4214,N_4671);
nand U9032 (N_9032,N_756,N_848);
and U9033 (N_9033,N_2809,N_2774);
nand U9034 (N_9034,N_1705,N_3947);
or U9035 (N_9035,N_1196,N_2005);
nor U9036 (N_9036,N_1165,N_1675);
nand U9037 (N_9037,N_2198,N_2478);
nor U9038 (N_9038,N_3499,N_4514);
nor U9039 (N_9039,N_2701,N_1781);
and U9040 (N_9040,N_343,N_1221);
or U9041 (N_9041,N_40,N_1002);
nand U9042 (N_9042,N_2567,N_4512);
or U9043 (N_9043,N_2622,N_1170);
and U9044 (N_9044,N_3792,N_610);
nand U9045 (N_9045,N_4572,N_2196);
or U9046 (N_9046,N_510,N_2294);
nor U9047 (N_9047,N_3885,N_666);
xor U9048 (N_9048,N_4836,N_4283);
or U9049 (N_9049,N_4897,N_3939);
or U9050 (N_9050,N_4954,N_817);
nor U9051 (N_9051,N_1397,N_959);
and U9052 (N_9052,N_619,N_469);
and U9053 (N_9053,N_4137,N_3435);
or U9054 (N_9054,N_789,N_3013);
xnor U9055 (N_9055,N_809,N_4507);
nand U9056 (N_9056,N_4643,N_4767);
nor U9057 (N_9057,N_1863,N_1004);
nor U9058 (N_9058,N_1693,N_4441);
xnor U9059 (N_9059,N_4528,N_4019);
nand U9060 (N_9060,N_1049,N_1806);
or U9061 (N_9061,N_4146,N_2500);
nor U9062 (N_9062,N_1036,N_471);
nor U9063 (N_9063,N_4952,N_1012);
or U9064 (N_9064,N_1536,N_314);
or U9065 (N_9065,N_1713,N_3754);
and U9066 (N_9066,N_4671,N_2118);
or U9067 (N_9067,N_4945,N_1904);
nand U9068 (N_9068,N_1630,N_758);
nor U9069 (N_9069,N_4163,N_3483);
nor U9070 (N_9070,N_582,N_522);
nor U9071 (N_9071,N_1641,N_4717);
nor U9072 (N_9072,N_445,N_3236);
nand U9073 (N_9073,N_2830,N_3091);
and U9074 (N_9074,N_1188,N_2262);
and U9075 (N_9075,N_677,N_987);
nand U9076 (N_9076,N_3117,N_1647);
xor U9077 (N_9077,N_1182,N_1690);
and U9078 (N_9078,N_4639,N_1809);
and U9079 (N_9079,N_1728,N_4786);
or U9080 (N_9080,N_4135,N_46);
or U9081 (N_9081,N_4141,N_3977);
and U9082 (N_9082,N_478,N_2366);
or U9083 (N_9083,N_4469,N_3928);
or U9084 (N_9084,N_4649,N_1857);
nand U9085 (N_9085,N_2953,N_4285);
nor U9086 (N_9086,N_2166,N_4150);
xor U9087 (N_9087,N_587,N_4416);
nor U9088 (N_9088,N_4952,N_2813);
xor U9089 (N_9089,N_4355,N_4335);
nand U9090 (N_9090,N_307,N_2927);
and U9091 (N_9091,N_959,N_3995);
nor U9092 (N_9092,N_1186,N_50);
or U9093 (N_9093,N_2550,N_4939);
or U9094 (N_9094,N_1777,N_3621);
nand U9095 (N_9095,N_560,N_1160);
and U9096 (N_9096,N_3211,N_3219);
and U9097 (N_9097,N_4775,N_3957);
nand U9098 (N_9098,N_3374,N_3186);
and U9099 (N_9099,N_715,N_3212);
or U9100 (N_9100,N_1021,N_3281);
nor U9101 (N_9101,N_4262,N_4246);
nor U9102 (N_9102,N_1749,N_740);
nor U9103 (N_9103,N_2526,N_4645);
or U9104 (N_9104,N_4464,N_1588);
or U9105 (N_9105,N_3993,N_2089);
or U9106 (N_9106,N_4774,N_4924);
nor U9107 (N_9107,N_3297,N_4588);
xor U9108 (N_9108,N_1847,N_431);
nor U9109 (N_9109,N_829,N_493);
nand U9110 (N_9110,N_1125,N_3984);
nor U9111 (N_9111,N_3237,N_418);
nand U9112 (N_9112,N_2856,N_4496);
nor U9113 (N_9113,N_1595,N_3249);
nor U9114 (N_9114,N_4774,N_2122);
and U9115 (N_9115,N_911,N_517);
or U9116 (N_9116,N_4745,N_2598);
nand U9117 (N_9117,N_418,N_3167);
and U9118 (N_9118,N_872,N_1195);
or U9119 (N_9119,N_351,N_4070);
nor U9120 (N_9120,N_2625,N_331);
xor U9121 (N_9121,N_2644,N_4256);
nand U9122 (N_9122,N_4610,N_4597);
nor U9123 (N_9123,N_84,N_640);
xor U9124 (N_9124,N_3012,N_3941);
nand U9125 (N_9125,N_1534,N_4074);
xnor U9126 (N_9126,N_1096,N_3088);
or U9127 (N_9127,N_2825,N_918);
and U9128 (N_9128,N_2872,N_3295);
nor U9129 (N_9129,N_4957,N_1673);
nand U9130 (N_9130,N_2782,N_2547);
xnor U9131 (N_9131,N_1307,N_2518);
and U9132 (N_9132,N_2224,N_3526);
nor U9133 (N_9133,N_3462,N_2680);
xor U9134 (N_9134,N_1816,N_1886);
nor U9135 (N_9135,N_3733,N_2570);
nand U9136 (N_9136,N_3980,N_428);
or U9137 (N_9137,N_1042,N_1860);
nand U9138 (N_9138,N_986,N_3899);
nand U9139 (N_9139,N_734,N_2011);
or U9140 (N_9140,N_2090,N_3912);
or U9141 (N_9141,N_1568,N_1993);
xor U9142 (N_9142,N_4628,N_613);
xnor U9143 (N_9143,N_2025,N_1767);
xor U9144 (N_9144,N_1600,N_540);
nand U9145 (N_9145,N_1447,N_1513);
or U9146 (N_9146,N_3786,N_2082);
nor U9147 (N_9147,N_1949,N_4075);
nor U9148 (N_9148,N_2642,N_314);
or U9149 (N_9149,N_4728,N_721);
or U9150 (N_9150,N_2261,N_509);
nor U9151 (N_9151,N_1309,N_4678);
nand U9152 (N_9152,N_2864,N_4877);
and U9153 (N_9153,N_3654,N_199);
xor U9154 (N_9154,N_577,N_86);
and U9155 (N_9155,N_691,N_917);
xnor U9156 (N_9156,N_4218,N_495);
nand U9157 (N_9157,N_961,N_3996);
xor U9158 (N_9158,N_3352,N_1713);
nand U9159 (N_9159,N_4589,N_1213);
and U9160 (N_9160,N_1778,N_808);
or U9161 (N_9161,N_2825,N_3086);
nand U9162 (N_9162,N_2235,N_2009);
and U9163 (N_9163,N_3928,N_2202);
and U9164 (N_9164,N_254,N_3053);
and U9165 (N_9165,N_422,N_1596);
and U9166 (N_9166,N_2858,N_4052);
nand U9167 (N_9167,N_450,N_1316);
and U9168 (N_9168,N_171,N_1329);
or U9169 (N_9169,N_1769,N_2240);
nor U9170 (N_9170,N_409,N_3123);
or U9171 (N_9171,N_2169,N_3520);
nor U9172 (N_9172,N_948,N_86);
nand U9173 (N_9173,N_574,N_4644);
xor U9174 (N_9174,N_1618,N_322);
xor U9175 (N_9175,N_4993,N_1190);
nor U9176 (N_9176,N_1203,N_599);
and U9177 (N_9177,N_4910,N_81);
xnor U9178 (N_9178,N_4501,N_1830);
nand U9179 (N_9179,N_4861,N_2297);
xor U9180 (N_9180,N_3361,N_4225);
and U9181 (N_9181,N_1074,N_2173);
and U9182 (N_9182,N_4585,N_517);
nor U9183 (N_9183,N_4555,N_2742);
xnor U9184 (N_9184,N_3188,N_3392);
or U9185 (N_9185,N_2922,N_1789);
and U9186 (N_9186,N_1158,N_59);
nor U9187 (N_9187,N_2099,N_4337);
nor U9188 (N_9188,N_1898,N_2503);
and U9189 (N_9189,N_3669,N_2047);
nor U9190 (N_9190,N_1735,N_2833);
xnor U9191 (N_9191,N_1053,N_2535);
or U9192 (N_9192,N_2841,N_2753);
xnor U9193 (N_9193,N_1324,N_2000);
xor U9194 (N_9194,N_4773,N_912);
xor U9195 (N_9195,N_3826,N_1371);
nor U9196 (N_9196,N_4932,N_1537);
xnor U9197 (N_9197,N_4567,N_4436);
and U9198 (N_9198,N_2475,N_1137);
xnor U9199 (N_9199,N_3035,N_4848);
nor U9200 (N_9200,N_1116,N_4729);
or U9201 (N_9201,N_2366,N_4973);
nand U9202 (N_9202,N_1444,N_3358);
xnor U9203 (N_9203,N_274,N_4965);
and U9204 (N_9204,N_4553,N_4261);
and U9205 (N_9205,N_1752,N_1035);
xnor U9206 (N_9206,N_1103,N_1431);
nand U9207 (N_9207,N_3088,N_3238);
nand U9208 (N_9208,N_3490,N_2253);
nor U9209 (N_9209,N_3981,N_4499);
nand U9210 (N_9210,N_3133,N_626);
and U9211 (N_9211,N_778,N_4267);
and U9212 (N_9212,N_1729,N_4558);
and U9213 (N_9213,N_4667,N_4016);
nand U9214 (N_9214,N_476,N_4081);
xor U9215 (N_9215,N_3928,N_4707);
nor U9216 (N_9216,N_895,N_2975);
nor U9217 (N_9217,N_1744,N_948);
nand U9218 (N_9218,N_2885,N_2966);
or U9219 (N_9219,N_3482,N_2565);
nor U9220 (N_9220,N_2151,N_724);
xor U9221 (N_9221,N_3619,N_329);
xnor U9222 (N_9222,N_1711,N_4065);
xnor U9223 (N_9223,N_2094,N_3902);
nor U9224 (N_9224,N_3767,N_1803);
nand U9225 (N_9225,N_1804,N_2569);
and U9226 (N_9226,N_4532,N_4980);
and U9227 (N_9227,N_3736,N_4993);
nand U9228 (N_9228,N_3738,N_3972);
nand U9229 (N_9229,N_4882,N_672);
nor U9230 (N_9230,N_3434,N_2528);
and U9231 (N_9231,N_330,N_4789);
nor U9232 (N_9232,N_539,N_356);
nor U9233 (N_9233,N_3170,N_298);
or U9234 (N_9234,N_3324,N_242);
nand U9235 (N_9235,N_972,N_2271);
nor U9236 (N_9236,N_1619,N_4730);
xnor U9237 (N_9237,N_425,N_2915);
nor U9238 (N_9238,N_1476,N_95);
and U9239 (N_9239,N_653,N_4023);
nand U9240 (N_9240,N_1629,N_3771);
nor U9241 (N_9241,N_4831,N_1108);
xnor U9242 (N_9242,N_2162,N_1947);
nand U9243 (N_9243,N_3797,N_1906);
xor U9244 (N_9244,N_4923,N_3551);
xor U9245 (N_9245,N_1297,N_4255);
nor U9246 (N_9246,N_4955,N_2989);
and U9247 (N_9247,N_3158,N_4431);
or U9248 (N_9248,N_522,N_4807);
or U9249 (N_9249,N_1103,N_2188);
and U9250 (N_9250,N_42,N_124);
xor U9251 (N_9251,N_2474,N_2413);
and U9252 (N_9252,N_3287,N_2118);
xor U9253 (N_9253,N_1933,N_1782);
xor U9254 (N_9254,N_3331,N_4232);
nor U9255 (N_9255,N_3790,N_2905);
nand U9256 (N_9256,N_1459,N_2529);
xnor U9257 (N_9257,N_3897,N_965);
and U9258 (N_9258,N_4154,N_1248);
or U9259 (N_9259,N_3434,N_3230);
or U9260 (N_9260,N_3428,N_4111);
nand U9261 (N_9261,N_1605,N_4457);
nor U9262 (N_9262,N_5,N_2501);
or U9263 (N_9263,N_1403,N_4339);
nor U9264 (N_9264,N_2458,N_671);
nand U9265 (N_9265,N_2850,N_3822);
and U9266 (N_9266,N_2617,N_3290);
nand U9267 (N_9267,N_1612,N_1879);
and U9268 (N_9268,N_1005,N_37);
nand U9269 (N_9269,N_74,N_2928);
nand U9270 (N_9270,N_317,N_1231);
nand U9271 (N_9271,N_3314,N_559);
and U9272 (N_9272,N_1530,N_1330);
nor U9273 (N_9273,N_2507,N_3063);
or U9274 (N_9274,N_4618,N_1307);
nand U9275 (N_9275,N_3610,N_483);
xor U9276 (N_9276,N_3093,N_627);
nand U9277 (N_9277,N_3712,N_3072);
and U9278 (N_9278,N_2945,N_3243);
xor U9279 (N_9279,N_4518,N_3316);
nand U9280 (N_9280,N_1354,N_2386);
and U9281 (N_9281,N_4478,N_4933);
nor U9282 (N_9282,N_838,N_589);
xnor U9283 (N_9283,N_3344,N_482);
and U9284 (N_9284,N_4477,N_2853);
nor U9285 (N_9285,N_2424,N_3074);
xor U9286 (N_9286,N_4608,N_4820);
nor U9287 (N_9287,N_2051,N_4395);
nor U9288 (N_9288,N_1177,N_4005);
xnor U9289 (N_9289,N_342,N_4435);
nand U9290 (N_9290,N_613,N_2177);
and U9291 (N_9291,N_2820,N_4524);
nand U9292 (N_9292,N_504,N_3274);
nor U9293 (N_9293,N_2955,N_4770);
and U9294 (N_9294,N_1967,N_1786);
nor U9295 (N_9295,N_4420,N_1016);
and U9296 (N_9296,N_1150,N_3712);
xnor U9297 (N_9297,N_1300,N_1697);
nand U9298 (N_9298,N_1551,N_3663);
xnor U9299 (N_9299,N_4531,N_1680);
and U9300 (N_9300,N_3753,N_1254);
nor U9301 (N_9301,N_4316,N_3076);
nand U9302 (N_9302,N_4878,N_4403);
xnor U9303 (N_9303,N_1385,N_3627);
nor U9304 (N_9304,N_3474,N_4792);
nor U9305 (N_9305,N_3455,N_693);
and U9306 (N_9306,N_3685,N_4778);
nor U9307 (N_9307,N_3832,N_1769);
xnor U9308 (N_9308,N_64,N_565);
nor U9309 (N_9309,N_643,N_4689);
xnor U9310 (N_9310,N_2972,N_2283);
and U9311 (N_9311,N_384,N_3997);
or U9312 (N_9312,N_4486,N_3429);
or U9313 (N_9313,N_4562,N_3479);
nand U9314 (N_9314,N_1812,N_4519);
or U9315 (N_9315,N_1728,N_3386);
nor U9316 (N_9316,N_1076,N_1483);
xor U9317 (N_9317,N_4399,N_3573);
and U9318 (N_9318,N_239,N_4243);
and U9319 (N_9319,N_1342,N_2734);
nand U9320 (N_9320,N_4449,N_2437);
nand U9321 (N_9321,N_3490,N_233);
nand U9322 (N_9322,N_4089,N_668);
or U9323 (N_9323,N_4093,N_1816);
or U9324 (N_9324,N_1054,N_619);
nor U9325 (N_9325,N_1481,N_419);
nand U9326 (N_9326,N_4438,N_4753);
nand U9327 (N_9327,N_1454,N_4628);
or U9328 (N_9328,N_4613,N_3694);
and U9329 (N_9329,N_1348,N_2314);
nand U9330 (N_9330,N_4210,N_4777);
nor U9331 (N_9331,N_1939,N_2478);
xnor U9332 (N_9332,N_4710,N_2879);
and U9333 (N_9333,N_2537,N_3135);
xnor U9334 (N_9334,N_1684,N_4201);
nor U9335 (N_9335,N_4550,N_261);
xor U9336 (N_9336,N_2577,N_2421);
nor U9337 (N_9337,N_4970,N_913);
xor U9338 (N_9338,N_1429,N_1515);
and U9339 (N_9339,N_1530,N_2376);
or U9340 (N_9340,N_2040,N_4951);
nand U9341 (N_9341,N_3976,N_2073);
nand U9342 (N_9342,N_4869,N_3068);
nand U9343 (N_9343,N_927,N_4322);
nand U9344 (N_9344,N_4153,N_809);
nand U9345 (N_9345,N_572,N_4990);
and U9346 (N_9346,N_1101,N_3382);
xor U9347 (N_9347,N_379,N_237);
nand U9348 (N_9348,N_1494,N_3514);
or U9349 (N_9349,N_631,N_1346);
xor U9350 (N_9350,N_3373,N_3949);
nor U9351 (N_9351,N_3336,N_218);
nand U9352 (N_9352,N_4329,N_660);
and U9353 (N_9353,N_661,N_3002);
and U9354 (N_9354,N_1483,N_2486);
nand U9355 (N_9355,N_4444,N_4872);
and U9356 (N_9356,N_4280,N_4367);
or U9357 (N_9357,N_587,N_3045);
nor U9358 (N_9358,N_4736,N_927);
nand U9359 (N_9359,N_733,N_3263);
or U9360 (N_9360,N_4526,N_2765);
or U9361 (N_9361,N_3701,N_3338);
nor U9362 (N_9362,N_778,N_4152);
nand U9363 (N_9363,N_1842,N_1458);
nand U9364 (N_9364,N_921,N_188);
nor U9365 (N_9365,N_2628,N_1004);
or U9366 (N_9366,N_362,N_2848);
nor U9367 (N_9367,N_126,N_4244);
or U9368 (N_9368,N_4944,N_4593);
nor U9369 (N_9369,N_3941,N_2942);
nor U9370 (N_9370,N_2139,N_4408);
or U9371 (N_9371,N_2149,N_4042);
nand U9372 (N_9372,N_3466,N_2576);
nor U9373 (N_9373,N_3588,N_3348);
or U9374 (N_9374,N_694,N_1709);
or U9375 (N_9375,N_1633,N_4659);
nor U9376 (N_9376,N_2411,N_220);
nor U9377 (N_9377,N_275,N_2950);
nor U9378 (N_9378,N_1460,N_4963);
or U9379 (N_9379,N_1968,N_3255);
xnor U9380 (N_9380,N_1230,N_2909);
nand U9381 (N_9381,N_3747,N_4409);
or U9382 (N_9382,N_4890,N_2907);
nor U9383 (N_9383,N_486,N_4899);
or U9384 (N_9384,N_3409,N_1601);
xnor U9385 (N_9385,N_3052,N_2451);
nor U9386 (N_9386,N_2766,N_3046);
xnor U9387 (N_9387,N_3858,N_1594);
or U9388 (N_9388,N_1121,N_692);
nand U9389 (N_9389,N_3628,N_3810);
or U9390 (N_9390,N_1588,N_3692);
and U9391 (N_9391,N_3755,N_1155);
nor U9392 (N_9392,N_127,N_1254);
nand U9393 (N_9393,N_3711,N_1214);
nand U9394 (N_9394,N_4487,N_1187);
xor U9395 (N_9395,N_966,N_987);
nor U9396 (N_9396,N_116,N_2025);
nand U9397 (N_9397,N_4118,N_1507);
nor U9398 (N_9398,N_4457,N_143);
and U9399 (N_9399,N_942,N_4188);
or U9400 (N_9400,N_4337,N_4963);
xnor U9401 (N_9401,N_4635,N_1216);
nor U9402 (N_9402,N_3159,N_2852);
nor U9403 (N_9403,N_3919,N_3182);
xnor U9404 (N_9404,N_3254,N_4498);
xor U9405 (N_9405,N_2323,N_742);
nor U9406 (N_9406,N_2168,N_4081);
or U9407 (N_9407,N_3823,N_1085);
nand U9408 (N_9408,N_1606,N_1841);
nor U9409 (N_9409,N_4482,N_3887);
nor U9410 (N_9410,N_3236,N_3419);
and U9411 (N_9411,N_2485,N_4368);
or U9412 (N_9412,N_2068,N_4198);
nand U9413 (N_9413,N_2382,N_4492);
nand U9414 (N_9414,N_4470,N_575);
nand U9415 (N_9415,N_3199,N_4284);
nor U9416 (N_9416,N_2965,N_1672);
or U9417 (N_9417,N_2263,N_4523);
and U9418 (N_9418,N_4156,N_1545);
nand U9419 (N_9419,N_3153,N_2932);
or U9420 (N_9420,N_4630,N_2103);
xor U9421 (N_9421,N_624,N_887);
or U9422 (N_9422,N_2271,N_3361);
nor U9423 (N_9423,N_1991,N_3744);
nand U9424 (N_9424,N_1598,N_1429);
and U9425 (N_9425,N_201,N_3375);
nor U9426 (N_9426,N_1238,N_494);
xnor U9427 (N_9427,N_4044,N_379);
nor U9428 (N_9428,N_2595,N_956);
nor U9429 (N_9429,N_3796,N_1976);
nand U9430 (N_9430,N_1017,N_2463);
nand U9431 (N_9431,N_2688,N_574);
or U9432 (N_9432,N_3616,N_2582);
nor U9433 (N_9433,N_1717,N_4967);
or U9434 (N_9434,N_614,N_4282);
and U9435 (N_9435,N_628,N_4178);
nand U9436 (N_9436,N_1917,N_1674);
xor U9437 (N_9437,N_544,N_4797);
nor U9438 (N_9438,N_3348,N_2627);
nand U9439 (N_9439,N_3497,N_4533);
nand U9440 (N_9440,N_3961,N_2480);
xnor U9441 (N_9441,N_4598,N_4211);
nand U9442 (N_9442,N_3615,N_962);
and U9443 (N_9443,N_3670,N_1732);
xor U9444 (N_9444,N_1132,N_1874);
or U9445 (N_9445,N_4715,N_3826);
and U9446 (N_9446,N_2944,N_2788);
and U9447 (N_9447,N_2554,N_4879);
or U9448 (N_9448,N_4285,N_3068);
and U9449 (N_9449,N_3120,N_1122);
or U9450 (N_9450,N_2596,N_3588);
or U9451 (N_9451,N_536,N_2217);
nand U9452 (N_9452,N_1781,N_2062);
or U9453 (N_9453,N_1789,N_2887);
or U9454 (N_9454,N_661,N_4008);
and U9455 (N_9455,N_3207,N_2734);
and U9456 (N_9456,N_103,N_697);
xor U9457 (N_9457,N_1891,N_3407);
or U9458 (N_9458,N_4071,N_3765);
and U9459 (N_9459,N_2979,N_1696);
xor U9460 (N_9460,N_4992,N_2863);
or U9461 (N_9461,N_2049,N_1651);
nand U9462 (N_9462,N_3086,N_3151);
xnor U9463 (N_9463,N_975,N_2632);
nand U9464 (N_9464,N_4404,N_133);
and U9465 (N_9465,N_1476,N_2458);
or U9466 (N_9466,N_3734,N_2671);
xnor U9467 (N_9467,N_1925,N_774);
and U9468 (N_9468,N_4889,N_4992);
and U9469 (N_9469,N_2541,N_4921);
xnor U9470 (N_9470,N_2091,N_4981);
nor U9471 (N_9471,N_3391,N_4153);
nor U9472 (N_9472,N_3615,N_4020);
xnor U9473 (N_9473,N_2927,N_4440);
nor U9474 (N_9474,N_794,N_188);
and U9475 (N_9475,N_1795,N_949);
or U9476 (N_9476,N_3121,N_921);
and U9477 (N_9477,N_3417,N_3505);
and U9478 (N_9478,N_4474,N_882);
xor U9479 (N_9479,N_3046,N_2212);
nand U9480 (N_9480,N_4339,N_3207);
nand U9481 (N_9481,N_3343,N_1783);
nor U9482 (N_9482,N_4816,N_3373);
nand U9483 (N_9483,N_629,N_1190);
or U9484 (N_9484,N_827,N_51);
xnor U9485 (N_9485,N_1819,N_4868);
or U9486 (N_9486,N_3128,N_3763);
and U9487 (N_9487,N_2323,N_1713);
and U9488 (N_9488,N_3356,N_879);
nor U9489 (N_9489,N_4888,N_1521);
nand U9490 (N_9490,N_998,N_4753);
and U9491 (N_9491,N_1660,N_2184);
and U9492 (N_9492,N_4259,N_4666);
and U9493 (N_9493,N_389,N_2797);
nand U9494 (N_9494,N_4711,N_690);
nand U9495 (N_9495,N_807,N_3324);
or U9496 (N_9496,N_2548,N_4988);
or U9497 (N_9497,N_1784,N_3733);
nand U9498 (N_9498,N_1048,N_3228);
and U9499 (N_9499,N_1126,N_2825);
xnor U9500 (N_9500,N_696,N_4380);
nor U9501 (N_9501,N_2824,N_1844);
and U9502 (N_9502,N_1206,N_423);
and U9503 (N_9503,N_768,N_3836);
xor U9504 (N_9504,N_2397,N_1766);
or U9505 (N_9505,N_3928,N_1891);
nand U9506 (N_9506,N_369,N_2735);
nor U9507 (N_9507,N_1228,N_1168);
xor U9508 (N_9508,N_4811,N_3238);
xnor U9509 (N_9509,N_3975,N_1430);
nor U9510 (N_9510,N_2937,N_4480);
xnor U9511 (N_9511,N_1545,N_2627);
nor U9512 (N_9512,N_4390,N_4243);
nor U9513 (N_9513,N_1026,N_4104);
and U9514 (N_9514,N_4281,N_174);
xor U9515 (N_9515,N_1130,N_1056);
xor U9516 (N_9516,N_768,N_3990);
or U9517 (N_9517,N_2257,N_6);
or U9518 (N_9518,N_1062,N_1744);
nand U9519 (N_9519,N_1664,N_4847);
nor U9520 (N_9520,N_2401,N_1466);
and U9521 (N_9521,N_2443,N_4385);
xor U9522 (N_9522,N_4495,N_3987);
xnor U9523 (N_9523,N_2731,N_874);
nor U9524 (N_9524,N_1809,N_1897);
nand U9525 (N_9525,N_4757,N_1312);
and U9526 (N_9526,N_2220,N_1943);
xnor U9527 (N_9527,N_324,N_3962);
nor U9528 (N_9528,N_3405,N_627);
xor U9529 (N_9529,N_1917,N_4443);
nor U9530 (N_9530,N_2951,N_4168);
nor U9531 (N_9531,N_350,N_4095);
xnor U9532 (N_9532,N_52,N_2401);
nand U9533 (N_9533,N_4084,N_160);
nand U9534 (N_9534,N_2403,N_4914);
or U9535 (N_9535,N_104,N_1045);
nand U9536 (N_9536,N_1821,N_4058);
nand U9537 (N_9537,N_2765,N_2992);
xor U9538 (N_9538,N_483,N_535);
or U9539 (N_9539,N_799,N_4766);
nand U9540 (N_9540,N_571,N_4509);
nor U9541 (N_9541,N_4544,N_3955);
nor U9542 (N_9542,N_1046,N_1951);
and U9543 (N_9543,N_1377,N_4959);
nand U9544 (N_9544,N_1371,N_696);
xnor U9545 (N_9545,N_2452,N_4766);
nand U9546 (N_9546,N_3624,N_1537);
nand U9547 (N_9547,N_4272,N_2588);
and U9548 (N_9548,N_3794,N_3352);
nand U9549 (N_9549,N_2177,N_4593);
xnor U9550 (N_9550,N_2932,N_2642);
xor U9551 (N_9551,N_3398,N_4485);
and U9552 (N_9552,N_1592,N_3623);
or U9553 (N_9553,N_3295,N_1927);
and U9554 (N_9554,N_437,N_3872);
xnor U9555 (N_9555,N_51,N_4117);
or U9556 (N_9556,N_1533,N_4610);
or U9557 (N_9557,N_119,N_4206);
nor U9558 (N_9558,N_2825,N_4526);
xnor U9559 (N_9559,N_1499,N_258);
nor U9560 (N_9560,N_1102,N_4821);
xnor U9561 (N_9561,N_2377,N_1407);
nand U9562 (N_9562,N_602,N_4061);
nor U9563 (N_9563,N_1452,N_3472);
and U9564 (N_9564,N_1924,N_1516);
or U9565 (N_9565,N_3010,N_2652);
xor U9566 (N_9566,N_2055,N_3410);
or U9567 (N_9567,N_1337,N_3194);
and U9568 (N_9568,N_3349,N_4383);
nor U9569 (N_9569,N_561,N_4090);
xor U9570 (N_9570,N_989,N_3445);
nand U9571 (N_9571,N_788,N_2504);
and U9572 (N_9572,N_2852,N_993);
nor U9573 (N_9573,N_3927,N_2612);
or U9574 (N_9574,N_3953,N_165);
and U9575 (N_9575,N_2992,N_856);
and U9576 (N_9576,N_2397,N_2820);
xnor U9577 (N_9577,N_1911,N_4394);
nand U9578 (N_9578,N_20,N_4279);
or U9579 (N_9579,N_1013,N_928);
or U9580 (N_9580,N_3409,N_2553);
nand U9581 (N_9581,N_1197,N_1573);
nor U9582 (N_9582,N_1420,N_2865);
xnor U9583 (N_9583,N_2757,N_1132);
nor U9584 (N_9584,N_2036,N_828);
nand U9585 (N_9585,N_437,N_2945);
nand U9586 (N_9586,N_755,N_790);
nor U9587 (N_9587,N_592,N_31);
and U9588 (N_9588,N_1242,N_4973);
xnor U9589 (N_9589,N_2976,N_2096);
or U9590 (N_9590,N_3667,N_1792);
nor U9591 (N_9591,N_4914,N_2946);
xor U9592 (N_9592,N_2721,N_443);
and U9593 (N_9593,N_4997,N_3112);
nand U9594 (N_9594,N_3095,N_2836);
or U9595 (N_9595,N_3999,N_361);
xnor U9596 (N_9596,N_3122,N_2961);
xnor U9597 (N_9597,N_701,N_3085);
xnor U9598 (N_9598,N_1894,N_2040);
xnor U9599 (N_9599,N_3125,N_3291);
nor U9600 (N_9600,N_4605,N_3258);
nand U9601 (N_9601,N_3164,N_2617);
or U9602 (N_9602,N_3605,N_652);
and U9603 (N_9603,N_2489,N_2973);
or U9604 (N_9604,N_4127,N_2782);
xnor U9605 (N_9605,N_759,N_2226);
nand U9606 (N_9606,N_3886,N_3398);
nand U9607 (N_9607,N_2843,N_309);
or U9608 (N_9608,N_325,N_820);
xnor U9609 (N_9609,N_3497,N_39);
xor U9610 (N_9610,N_2586,N_82);
xnor U9611 (N_9611,N_910,N_3949);
nor U9612 (N_9612,N_3865,N_1615);
nor U9613 (N_9613,N_3889,N_1421);
xnor U9614 (N_9614,N_3813,N_2006);
nand U9615 (N_9615,N_3109,N_3);
xnor U9616 (N_9616,N_2356,N_2748);
and U9617 (N_9617,N_3166,N_341);
and U9618 (N_9618,N_911,N_790);
nor U9619 (N_9619,N_794,N_1515);
and U9620 (N_9620,N_835,N_2087);
nand U9621 (N_9621,N_4537,N_2796);
xor U9622 (N_9622,N_4424,N_2018);
and U9623 (N_9623,N_4700,N_56);
nor U9624 (N_9624,N_1629,N_3241);
xnor U9625 (N_9625,N_350,N_2060);
or U9626 (N_9626,N_2081,N_4884);
and U9627 (N_9627,N_2328,N_746);
or U9628 (N_9628,N_3405,N_3831);
or U9629 (N_9629,N_1100,N_4887);
and U9630 (N_9630,N_3265,N_1903);
nand U9631 (N_9631,N_1630,N_3);
nand U9632 (N_9632,N_1709,N_2757);
nor U9633 (N_9633,N_214,N_2358);
or U9634 (N_9634,N_2451,N_2264);
and U9635 (N_9635,N_3511,N_1674);
nor U9636 (N_9636,N_643,N_4930);
nand U9637 (N_9637,N_3408,N_1737);
and U9638 (N_9638,N_341,N_501);
nand U9639 (N_9639,N_624,N_4549);
xnor U9640 (N_9640,N_1826,N_259);
nor U9641 (N_9641,N_1861,N_1892);
xnor U9642 (N_9642,N_2115,N_3472);
or U9643 (N_9643,N_2167,N_4540);
xnor U9644 (N_9644,N_3245,N_2899);
and U9645 (N_9645,N_1235,N_3612);
nor U9646 (N_9646,N_4717,N_1073);
and U9647 (N_9647,N_3867,N_1193);
or U9648 (N_9648,N_1916,N_3359);
or U9649 (N_9649,N_1049,N_3792);
nor U9650 (N_9650,N_2948,N_1394);
xor U9651 (N_9651,N_1312,N_2126);
nand U9652 (N_9652,N_1363,N_3357);
nand U9653 (N_9653,N_741,N_713);
nor U9654 (N_9654,N_1826,N_2667);
nor U9655 (N_9655,N_4361,N_2440);
xnor U9656 (N_9656,N_300,N_3382);
xor U9657 (N_9657,N_686,N_1011);
or U9658 (N_9658,N_75,N_3909);
or U9659 (N_9659,N_4938,N_3903);
or U9660 (N_9660,N_2847,N_3670);
xnor U9661 (N_9661,N_3387,N_1167);
or U9662 (N_9662,N_345,N_4721);
nor U9663 (N_9663,N_364,N_4219);
nand U9664 (N_9664,N_1913,N_1189);
and U9665 (N_9665,N_1589,N_108);
nand U9666 (N_9666,N_3548,N_3593);
xnor U9667 (N_9667,N_4106,N_1466);
and U9668 (N_9668,N_2522,N_1000);
and U9669 (N_9669,N_1270,N_3624);
and U9670 (N_9670,N_1817,N_1811);
and U9671 (N_9671,N_3342,N_220);
and U9672 (N_9672,N_3875,N_1387);
nor U9673 (N_9673,N_1582,N_4748);
nand U9674 (N_9674,N_1130,N_826);
or U9675 (N_9675,N_1469,N_633);
xor U9676 (N_9676,N_3225,N_1923);
nor U9677 (N_9677,N_1890,N_3327);
nor U9678 (N_9678,N_1705,N_755);
xnor U9679 (N_9679,N_913,N_1216);
xor U9680 (N_9680,N_2475,N_1558);
or U9681 (N_9681,N_3876,N_493);
and U9682 (N_9682,N_1166,N_7);
nor U9683 (N_9683,N_4335,N_2131);
and U9684 (N_9684,N_764,N_4012);
nor U9685 (N_9685,N_687,N_1918);
xnor U9686 (N_9686,N_4747,N_1835);
and U9687 (N_9687,N_2033,N_2352);
nand U9688 (N_9688,N_588,N_2534);
nor U9689 (N_9689,N_2477,N_4136);
nand U9690 (N_9690,N_4151,N_1470);
or U9691 (N_9691,N_3558,N_2683);
nor U9692 (N_9692,N_2975,N_2459);
nand U9693 (N_9693,N_3529,N_2675);
xor U9694 (N_9694,N_4173,N_4059);
or U9695 (N_9695,N_4348,N_3790);
and U9696 (N_9696,N_4299,N_821);
or U9697 (N_9697,N_2420,N_121);
xnor U9698 (N_9698,N_4539,N_3826);
xnor U9699 (N_9699,N_2799,N_4151);
or U9700 (N_9700,N_3789,N_4094);
nand U9701 (N_9701,N_3598,N_543);
and U9702 (N_9702,N_1444,N_4033);
nor U9703 (N_9703,N_2456,N_4816);
or U9704 (N_9704,N_3984,N_178);
or U9705 (N_9705,N_477,N_453);
xor U9706 (N_9706,N_2037,N_78);
and U9707 (N_9707,N_3013,N_746);
or U9708 (N_9708,N_2269,N_3800);
or U9709 (N_9709,N_1317,N_4732);
nor U9710 (N_9710,N_1480,N_4224);
nand U9711 (N_9711,N_1909,N_1223);
nand U9712 (N_9712,N_3313,N_4491);
nand U9713 (N_9713,N_1885,N_1766);
or U9714 (N_9714,N_1691,N_693);
nand U9715 (N_9715,N_3483,N_1442);
xor U9716 (N_9716,N_4774,N_2151);
and U9717 (N_9717,N_2088,N_1612);
xor U9718 (N_9718,N_2163,N_4300);
or U9719 (N_9719,N_2019,N_3527);
xor U9720 (N_9720,N_3356,N_91);
nor U9721 (N_9721,N_711,N_2722);
nor U9722 (N_9722,N_2424,N_1226);
xor U9723 (N_9723,N_3930,N_2257);
or U9724 (N_9724,N_4040,N_4190);
xnor U9725 (N_9725,N_3153,N_473);
nor U9726 (N_9726,N_2191,N_1120);
nor U9727 (N_9727,N_4825,N_3778);
nand U9728 (N_9728,N_4764,N_3138);
or U9729 (N_9729,N_1860,N_2790);
nor U9730 (N_9730,N_3461,N_4048);
nor U9731 (N_9731,N_126,N_1578);
or U9732 (N_9732,N_800,N_2008);
nand U9733 (N_9733,N_3849,N_1239);
nor U9734 (N_9734,N_616,N_4682);
xor U9735 (N_9735,N_4967,N_3068);
nand U9736 (N_9736,N_1937,N_2375);
or U9737 (N_9737,N_250,N_937);
or U9738 (N_9738,N_2506,N_1596);
and U9739 (N_9739,N_2288,N_2045);
xor U9740 (N_9740,N_607,N_3474);
nand U9741 (N_9741,N_2806,N_4227);
xnor U9742 (N_9742,N_2036,N_1837);
xnor U9743 (N_9743,N_2183,N_3001);
or U9744 (N_9744,N_3780,N_2573);
nor U9745 (N_9745,N_4121,N_4086);
xor U9746 (N_9746,N_3067,N_67);
nand U9747 (N_9747,N_4338,N_4752);
nor U9748 (N_9748,N_614,N_2120);
and U9749 (N_9749,N_2174,N_2115);
nand U9750 (N_9750,N_3248,N_4934);
and U9751 (N_9751,N_2829,N_295);
nand U9752 (N_9752,N_2926,N_1815);
or U9753 (N_9753,N_2072,N_4964);
nand U9754 (N_9754,N_3019,N_1757);
xor U9755 (N_9755,N_3238,N_826);
nand U9756 (N_9756,N_2603,N_3051);
nor U9757 (N_9757,N_1184,N_1590);
or U9758 (N_9758,N_2551,N_2251);
xnor U9759 (N_9759,N_1368,N_0);
xnor U9760 (N_9760,N_4,N_4375);
nor U9761 (N_9761,N_168,N_246);
or U9762 (N_9762,N_2943,N_4503);
nand U9763 (N_9763,N_1226,N_3018);
and U9764 (N_9764,N_1197,N_1928);
xor U9765 (N_9765,N_3490,N_2862);
xor U9766 (N_9766,N_4761,N_2015);
or U9767 (N_9767,N_4207,N_1678);
nor U9768 (N_9768,N_452,N_1690);
nor U9769 (N_9769,N_654,N_1619);
or U9770 (N_9770,N_3799,N_4173);
and U9771 (N_9771,N_3355,N_2546);
or U9772 (N_9772,N_1443,N_1523);
nand U9773 (N_9773,N_2280,N_2457);
and U9774 (N_9774,N_2100,N_4522);
or U9775 (N_9775,N_2962,N_3545);
xnor U9776 (N_9776,N_1192,N_3695);
and U9777 (N_9777,N_176,N_1585);
and U9778 (N_9778,N_908,N_4661);
nor U9779 (N_9779,N_1246,N_2607);
xor U9780 (N_9780,N_4730,N_2764);
nor U9781 (N_9781,N_4252,N_1896);
nand U9782 (N_9782,N_1840,N_1237);
nor U9783 (N_9783,N_1954,N_3349);
xnor U9784 (N_9784,N_2307,N_2422);
xnor U9785 (N_9785,N_4611,N_4780);
nor U9786 (N_9786,N_1663,N_3254);
and U9787 (N_9787,N_4001,N_3127);
nor U9788 (N_9788,N_194,N_79);
nor U9789 (N_9789,N_568,N_1800);
or U9790 (N_9790,N_503,N_1279);
or U9791 (N_9791,N_4719,N_3889);
xor U9792 (N_9792,N_1487,N_3924);
and U9793 (N_9793,N_472,N_4136);
and U9794 (N_9794,N_2548,N_4543);
nand U9795 (N_9795,N_3198,N_3782);
xor U9796 (N_9796,N_912,N_159);
and U9797 (N_9797,N_3201,N_2702);
nand U9798 (N_9798,N_2070,N_3749);
nand U9799 (N_9799,N_1693,N_839);
nor U9800 (N_9800,N_1336,N_3163);
xnor U9801 (N_9801,N_1524,N_1684);
xor U9802 (N_9802,N_1111,N_3296);
nor U9803 (N_9803,N_1394,N_2871);
nand U9804 (N_9804,N_4807,N_4556);
and U9805 (N_9805,N_2309,N_3004);
and U9806 (N_9806,N_3564,N_3708);
or U9807 (N_9807,N_2810,N_3793);
nor U9808 (N_9808,N_1683,N_4194);
and U9809 (N_9809,N_3216,N_447);
and U9810 (N_9810,N_3967,N_4650);
nor U9811 (N_9811,N_3350,N_1434);
or U9812 (N_9812,N_4164,N_3203);
xnor U9813 (N_9813,N_2094,N_4444);
nand U9814 (N_9814,N_233,N_4060);
or U9815 (N_9815,N_2495,N_1851);
nor U9816 (N_9816,N_731,N_1460);
nor U9817 (N_9817,N_1254,N_3280);
xnor U9818 (N_9818,N_435,N_1090);
xnor U9819 (N_9819,N_729,N_3866);
nand U9820 (N_9820,N_1947,N_4697);
xnor U9821 (N_9821,N_945,N_2193);
nand U9822 (N_9822,N_3635,N_261);
xnor U9823 (N_9823,N_3766,N_3616);
xnor U9824 (N_9824,N_4273,N_966);
xnor U9825 (N_9825,N_557,N_4145);
xnor U9826 (N_9826,N_91,N_1722);
nor U9827 (N_9827,N_1307,N_1563);
xor U9828 (N_9828,N_3845,N_1227);
and U9829 (N_9829,N_1378,N_705);
xor U9830 (N_9830,N_3383,N_3454);
and U9831 (N_9831,N_2567,N_2892);
nand U9832 (N_9832,N_4641,N_1310);
or U9833 (N_9833,N_386,N_3963);
nor U9834 (N_9834,N_2167,N_3249);
xor U9835 (N_9835,N_4769,N_232);
and U9836 (N_9836,N_2769,N_4571);
or U9837 (N_9837,N_400,N_1654);
nor U9838 (N_9838,N_3352,N_2760);
and U9839 (N_9839,N_848,N_1909);
nor U9840 (N_9840,N_3954,N_4123);
and U9841 (N_9841,N_496,N_1436);
nor U9842 (N_9842,N_164,N_2181);
and U9843 (N_9843,N_2474,N_3091);
and U9844 (N_9844,N_1065,N_4235);
and U9845 (N_9845,N_4642,N_498);
and U9846 (N_9846,N_460,N_1823);
and U9847 (N_9847,N_1194,N_4475);
xnor U9848 (N_9848,N_393,N_1731);
and U9849 (N_9849,N_1252,N_1579);
xor U9850 (N_9850,N_3018,N_2466);
nor U9851 (N_9851,N_2116,N_3652);
nor U9852 (N_9852,N_2047,N_2566);
xnor U9853 (N_9853,N_2037,N_2425);
or U9854 (N_9854,N_3466,N_3700);
nand U9855 (N_9855,N_680,N_2760);
or U9856 (N_9856,N_4471,N_359);
nor U9857 (N_9857,N_3370,N_4998);
and U9858 (N_9858,N_177,N_4776);
and U9859 (N_9859,N_2677,N_3384);
nor U9860 (N_9860,N_971,N_1420);
xnor U9861 (N_9861,N_3053,N_4043);
and U9862 (N_9862,N_2161,N_929);
nor U9863 (N_9863,N_4149,N_4763);
and U9864 (N_9864,N_3575,N_2918);
xnor U9865 (N_9865,N_399,N_4537);
xnor U9866 (N_9866,N_957,N_2200);
and U9867 (N_9867,N_110,N_1840);
nor U9868 (N_9868,N_1699,N_3552);
or U9869 (N_9869,N_2421,N_3184);
nand U9870 (N_9870,N_3267,N_3836);
and U9871 (N_9871,N_2617,N_1010);
or U9872 (N_9872,N_2475,N_178);
nand U9873 (N_9873,N_2372,N_2808);
nand U9874 (N_9874,N_4253,N_1244);
nand U9875 (N_9875,N_4627,N_4728);
nand U9876 (N_9876,N_4011,N_4852);
nand U9877 (N_9877,N_3133,N_4017);
xnor U9878 (N_9878,N_1772,N_256);
nor U9879 (N_9879,N_655,N_1760);
nand U9880 (N_9880,N_739,N_4054);
or U9881 (N_9881,N_4363,N_4828);
nand U9882 (N_9882,N_983,N_2544);
and U9883 (N_9883,N_2676,N_1120);
nand U9884 (N_9884,N_2122,N_121);
and U9885 (N_9885,N_3878,N_3502);
or U9886 (N_9886,N_2719,N_473);
nor U9887 (N_9887,N_426,N_2428);
or U9888 (N_9888,N_138,N_196);
xor U9889 (N_9889,N_4034,N_1308);
or U9890 (N_9890,N_1064,N_1307);
nor U9891 (N_9891,N_1731,N_738);
xnor U9892 (N_9892,N_3597,N_447);
xor U9893 (N_9893,N_1615,N_1216);
nand U9894 (N_9894,N_2372,N_2441);
and U9895 (N_9895,N_502,N_2150);
and U9896 (N_9896,N_2314,N_1956);
and U9897 (N_9897,N_3422,N_1481);
nand U9898 (N_9898,N_3926,N_1162);
nand U9899 (N_9899,N_2738,N_3579);
and U9900 (N_9900,N_1859,N_4308);
or U9901 (N_9901,N_1916,N_4779);
nand U9902 (N_9902,N_1760,N_4957);
xor U9903 (N_9903,N_2819,N_1109);
nand U9904 (N_9904,N_4622,N_249);
or U9905 (N_9905,N_3642,N_4211);
xnor U9906 (N_9906,N_1911,N_4574);
or U9907 (N_9907,N_2377,N_4846);
nor U9908 (N_9908,N_1792,N_4098);
xor U9909 (N_9909,N_419,N_983);
and U9910 (N_9910,N_4320,N_2547);
xnor U9911 (N_9911,N_3694,N_1843);
xor U9912 (N_9912,N_3514,N_2520);
and U9913 (N_9913,N_2878,N_939);
xnor U9914 (N_9914,N_1221,N_488);
and U9915 (N_9915,N_342,N_3698);
or U9916 (N_9916,N_495,N_243);
and U9917 (N_9917,N_4,N_2443);
xor U9918 (N_9918,N_3151,N_904);
nor U9919 (N_9919,N_4714,N_2043);
and U9920 (N_9920,N_1566,N_3143);
and U9921 (N_9921,N_3921,N_1868);
nand U9922 (N_9922,N_1192,N_4232);
and U9923 (N_9923,N_720,N_655);
and U9924 (N_9924,N_4692,N_1443);
nand U9925 (N_9925,N_2550,N_4762);
nand U9926 (N_9926,N_868,N_4777);
or U9927 (N_9927,N_3704,N_2956);
or U9928 (N_9928,N_970,N_650);
xnor U9929 (N_9929,N_662,N_264);
nand U9930 (N_9930,N_608,N_2423);
or U9931 (N_9931,N_3028,N_2567);
xor U9932 (N_9932,N_1938,N_4185);
nand U9933 (N_9933,N_4247,N_367);
xnor U9934 (N_9934,N_1655,N_4392);
and U9935 (N_9935,N_4572,N_2674);
nand U9936 (N_9936,N_381,N_2032);
or U9937 (N_9937,N_1675,N_1480);
or U9938 (N_9938,N_1769,N_546);
nor U9939 (N_9939,N_4797,N_1031);
and U9940 (N_9940,N_877,N_1962);
and U9941 (N_9941,N_3761,N_2611);
nand U9942 (N_9942,N_4918,N_1623);
nand U9943 (N_9943,N_2072,N_4451);
nand U9944 (N_9944,N_41,N_1782);
nor U9945 (N_9945,N_1657,N_2291);
and U9946 (N_9946,N_1607,N_4110);
nand U9947 (N_9947,N_2193,N_1871);
or U9948 (N_9948,N_1419,N_4329);
and U9949 (N_9949,N_3224,N_821);
or U9950 (N_9950,N_1492,N_3756);
and U9951 (N_9951,N_446,N_3502);
nand U9952 (N_9952,N_385,N_3801);
nand U9953 (N_9953,N_2131,N_2279);
nand U9954 (N_9954,N_3079,N_3254);
and U9955 (N_9955,N_1054,N_1270);
xor U9956 (N_9956,N_4098,N_4472);
or U9957 (N_9957,N_1237,N_2906);
xnor U9958 (N_9958,N_4233,N_4147);
nor U9959 (N_9959,N_568,N_2733);
xnor U9960 (N_9960,N_3084,N_4541);
and U9961 (N_9961,N_144,N_2321);
and U9962 (N_9962,N_1464,N_1037);
nor U9963 (N_9963,N_965,N_2111);
or U9964 (N_9964,N_2679,N_2307);
and U9965 (N_9965,N_4181,N_1709);
nor U9966 (N_9966,N_1180,N_1867);
or U9967 (N_9967,N_3805,N_4950);
and U9968 (N_9968,N_3535,N_1671);
or U9969 (N_9969,N_4865,N_332);
nor U9970 (N_9970,N_233,N_1509);
nand U9971 (N_9971,N_4489,N_3980);
xnor U9972 (N_9972,N_3963,N_764);
nand U9973 (N_9973,N_2360,N_3663);
or U9974 (N_9974,N_3217,N_1465);
or U9975 (N_9975,N_4237,N_4435);
nor U9976 (N_9976,N_2809,N_4116);
and U9977 (N_9977,N_1039,N_4148);
xnor U9978 (N_9978,N_2677,N_1289);
and U9979 (N_9979,N_1618,N_272);
nand U9980 (N_9980,N_1506,N_427);
nand U9981 (N_9981,N_4832,N_2594);
or U9982 (N_9982,N_56,N_2762);
and U9983 (N_9983,N_3695,N_4911);
nand U9984 (N_9984,N_2025,N_1854);
nor U9985 (N_9985,N_2897,N_239);
and U9986 (N_9986,N_3664,N_629);
xor U9987 (N_9987,N_1407,N_3189);
or U9988 (N_9988,N_2986,N_3435);
nand U9989 (N_9989,N_1397,N_1628);
and U9990 (N_9990,N_1504,N_3246);
or U9991 (N_9991,N_109,N_4497);
nand U9992 (N_9992,N_3823,N_1562);
or U9993 (N_9993,N_3043,N_3163);
or U9994 (N_9994,N_261,N_209);
nand U9995 (N_9995,N_4477,N_1636);
nor U9996 (N_9996,N_2786,N_4225);
or U9997 (N_9997,N_1621,N_564);
nand U9998 (N_9998,N_2735,N_4643);
and U9999 (N_9999,N_3234,N_3062);
nand U10000 (N_10000,N_6189,N_5140);
nand U10001 (N_10001,N_6096,N_5375);
nand U10002 (N_10002,N_5447,N_9263);
nor U10003 (N_10003,N_7222,N_5281);
nor U10004 (N_10004,N_7982,N_5847);
and U10005 (N_10005,N_7703,N_8051);
xnor U10006 (N_10006,N_7950,N_9051);
nand U10007 (N_10007,N_5323,N_8883);
and U10008 (N_10008,N_6834,N_7103);
and U10009 (N_10009,N_7123,N_8748);
and U10010 (N_10010,N_7642,N_8287);
xnor U10011 (N_10011,N_9898,N_7890);
xor U10012 (N_10012,N_8201,N_9466);
and U10013 (N_10013,N_7005,N_7754);
and U10014 (N_10014,N_9628,N_8858);
and U10015 (N_10015,N_7900,N_6922);
or U10016 (N_10016,N_5940,N_6888);
and U10017 (N_10017,N_8388,N_6958);
or U10018 (N_10018,N_8677,N_5324);
or U10019 (N_10019,N_5529,N_7092);
xor U10020 (N_10020,N_5124,N_7139);
and U10021 (N_10021,N_6463,N_9750);
xor U10022 (N_10022,N_5951,N_6711);
or U10023 (N_10023,N_7290,N_9804);
xnor U10024 (N_10024,N_5679,N_7779);
nor U10025 (N_10025,N_5607,N_6854);
nor U10026 (N_10026,N_5631,N_7370);
or U10027 (N_10027,N_5967,N_5247);
nand U10028 (N_10028,N_6311,N_9534);
nand U10029 (N_10029,N_9245,N_8273);
xnor U10030 (N_10030,N_7111,N_8231);
and U10031 (N_10031,N_7035,N_7940);
and U10032 (N_10032,N_7130,N_5546);
or U10033 (N_10033,N_6914,N_7063);
xnor U10034 (N_10034,N_8684,N_5822);
or U10035 (N_10035,N_7125,N_5682);
xnor U10036 (N_10036,N_5540,N_8136);
or U10037 (N_10037,N_7456,N_5509);
and U10038 (N_10038,N_9574,N_9447);
or U10039 (N_10039,N_7104,N_8354);
and U10040 (N_10040,N_9114,N_9984);
and U10041 (N_10041,N_9860,N_7712);
or U10042 (N_10042,N_6484,N_9770);
nand U10043 (N_10043,N_7183,N_5470);
nand U10044 (N_10044,N_5922,N_6064);
and U10045 (N_10045,N_8185,N_9444);
nor U10046 (N_10046,N_9886,N_7659);
or U10047 (N_10047,N_9474,N_7473);
nand U10048 (N_10048,N_7804,N_7869);
and U10049 (N_10049,N_8798,N_8838);
and U10050 (N_10050,N_8847,N_7674);
nand U10051 (N_10051,N_7540,N_5126);
and U10052 (N_10052,N_7307,N_9838);
nand U10053 (N_10053,N_7590,N_6299);
and U10054 (N_10054,N_6348,N_6763);
and U10055 (N_10055,N_8471,N_7671);
and U10056 (N_10056,N_9455,N_9772);
xnor U10057 (N_10057,N_9739,N_5480);
nor U10058 (N_10058,N_7425,N_8258);
nand U10059 (N_10059,N_7335,N_7911);
xor U10060 (N_10060,N_7833,N_7858);
xnor U10061 (N_10061,N_8779,N_9759);
or U10062 (N_10062,N_8164,N_5634);
xnor U10063 (N_10063,N_8633,N_8813);
or U10064 (N_10064,N_9260,N_8652);
and U10065 (N_10065,N_9837,N_7166);
nor U10066 (N_10066,N_6894,N_7876);
xor U10067 (N_10067,N_6966,N_7587);
nor U10068 (N_10068,N_6669,N_8766);
nand U10069 (N_10069,N_5612,N_5418);
nor U10070 (N_10070,N_8458,N_9340);
nand U10071 (N_10071,N_6611,N_7791);
nand U10072 (N_10072,N_5037,N_5226);
xnor U10073 (N_10073,N_7354,N_6037);
and U10074 (N_10074,N_7592,N_7664);
nor U10075 (N_10075,N_8356,N_9244);
or U10076 (N_10076,N_5970,N_8674);
or U10077 (N_10077,N_5718,N_5563);
nand U10078 (N_10078,N_9951,N_6618);
nor U10079 (N_10079,N_7661,N_7666);
xor U10080 (N_10080,N_9981,N_5672);
and U10081 (N_10081,N_5830,N_8315);
or U10082 (N_10082,N_5639,N_9994);
xor U10083 (N_10083,N_9350,N_6731);
or U10084 (N_10084,N_7356,N_6367);
nor U10085 (N_10085,N_6572,N_6694);
or U10086 (N_10086,N_5963,N_9955);
nand U10087 (N_10087,N_5659,N_5971);
nand U10088 (N_10088,N_7640,N_9880);
nor U10089 (N_10089,N_5044,N_8196);
xor U10090 (N_10090,N_7541,N_6857);
xnor U10091 (N_10091,N_5255,N_9891);
xnor U10092 (N_10092,N_5845,N_7505);
xor U10093 (N_10093,N_9809,N_5163);
and U10094 (N_10094,N_9449,N_9776);
xnor U10095 (N_10095,N_5860,N_5493);
and U10096 (N_10096,N_5176,N_7156);
xor U10097 (N_10097,N_6068,N_7693);
nor U10098 (N_10098,N_7514,N_8954);
and U10099 (N_10099,N_6291,N_7377);
xnor U10100 (N_10100,N_8984,N_7714);
nor U10101 (N_10101,N_7716,N_8704);
nand U10102 (N_10102,N_8861,N_7360);
and U10103 (N_10103,N_8931,N_9013);
and U10104 (N_10104,N_9131,N_6858);
and U10105 (N_10105,N_7147,N_6401);
nor U10106 (N_10106,N_9042,N_8447);
xnor U10107 (N_10107,N_7470,N_7096);
xor U10108 (N_10108,N_9728,N_8599);
nor U10109 (N_10109,N_6636,N_7722);
xor U10110 (N_10110,N_6635,N_5249);
xor U10111 (N_10111,N_5646,N_5203);
and U10112 (N_10112,N_9366,N_6289);
xnor U10113 (N_10113,N_5614,N_8452);
nor U10114 (N_10114,N_9354,N_7174);
nor U10115 (N_10115,N_6728,N_9718);
and U10116 (N_10116,N_5537,N_8139);
xor U10117 (N_10117,N_6103,N_5328);
or U10118 (N_10118,N_7965,N_8152);
xnor U10119 (N_10119,N_5991,N_7769);
or U10120 (N_10120,N_8832,N_6087);
or U10121 (N_10121,N_5776,N_8419);
and U10122 (N_10122,N_8735,N_8805);
or U10123 (N_10123,N_7079,N_7095);
xnor U10124 (N_10124,N_8113,N_9963);
xor U10125 (N_10125,N_8584,N_9765);
nor U10126 (N_10126,N_5005,N_9351);
nor U10127 (N_10127,N_5178,N_8513);
xnor U10128 (N_10128,N_6327,N_6126);
or U10129 (N_10129,N_8585,N_5744);
and U10130 (N_10130,N_9814,N_9287);
nor U10131 (N_10131,N_9106,N_6623);
and U10132 (N_10132,N_5969,N_7195);
xor U10133 (N_10133,N_8836,N_6890);
or U10134 (N_10134,N_8294,N_9735);
nor U10135 (N_10135,N_9296,N_5851);
nor U10136 (N_10136,N_7181,N_7741);
xnor U10137 (N_10137,N_9933,N_5390);
and U10138 (N_10138,N_5012,N_8071);
nor U10139 (N_10139,N_6021,N_5272);
or U10140 (N_10140,N_7549,N_5087);
and U10141 (N_10141,N_8439,N_5371);
or U10142 (N_10142,N_5266,N_7022);
nand U10143 (N_10143,N_6417,N_8162);
and U10144 (N_10144,N_7085,N_8223);
xor U10145 (N_10145,N_7158,N_8739);
nand U10146 (N_10146,N_9241,N_9868);
and U10147 (N_10147,N_8877,N_6477);
and U10148 (N_10148,N_6221,N_8111);
nor U10149 (N_10149,N_8026,N_8450);
and U10150 (N_10150,N_8500,N_8322);
and U10151 (N_10151,N_8569,N_9542);
and U10152 (N_10152,N_7772,N_5974);
nor U10153 (N_10153,N_5652,N_5750);
xnor U10154 (N_10154,N_6673,N_8588);
and U10155 (N_10155,N_9655,N_9831);
xor U10156 (N_10156,N_8332,N_5849);
nand U10157 (N_10157,N_8522,N_9871);
nor U10158 (N_10158,N_5960,N_5271);
and U10159 (N_10159,N_6491,N_9974);
or U10160 (N_10160,N_6138,N_6295);
nor U10161 (N_10161,N_9352,N_9294);
xor U10162 (N_10162,N_7177,N_8644);
nand U10163 (N_10163,N_5472,N_9907);
nand U10164 (N_10164,N_9285,N_7534);
nor U10165 (N_10165,N_9635,N_8107);
nor U10166 (N_10166,N_9614,N_9458);
xnor U10167 (N_10167,N_7263,N_7961);
xnor U10168 (N_10168,N_8761,N_8446);
xor U10169 (N_10169,N_8243,N_5709);
nor U10170 (N_10170,N_5702,N_8815);
or U10171 (N_10171,N_7270,N_7586);
and U10172 (N_10172,N_8819,N_6577);
and U10173 (N_10173,N_9341,N_7972);
nand U10174 (N_10174,N_9423,N_7065);
or U10175 (N_10175,N_7831,N_7764);
and U10176 (N_10176,N_7854,N_6274);
and U10177 (N_10177,N_7364,N_8755);
or U10178 (N_10178,N_6581,N_9324);
xor U10179 (N_10179,N_9806,N_8765);
or U10180 (N_10180,N_8590,N_8023);
and U10181 (N_10181,N_6895,N_7271);
or U10182 (N_10182,N_6841,N_8080);
xor U10183 (N_10183,N_5107,N_6811);
nand U10184 (N_10184,N_9227,N_9038);
or U10185 (N_10185,N_7516,N_6789);
and U10186 (N_10186,N_5216,N_7896);
nor U10187 (N_10187,N_9870,N_8905);
and U10188 (N_10188,N_7999,N_6778);
nand U10189 (N_10189,N_6826,N_9566);
and U10190 (N_10190,N_6710,N_8002);
and U10191 (N_10191,N_7365,N_9248);
or U10192 (N_10192,N_9454,N_9191);
nor U10193 (N_10193,N_5399,N_7368);
nand U10194 (N_10194,N_6297,N_5411);
and U10195 (N_10195,N_5731,N_8682);
xor U10196 (N_10196,N_8799,N_5597);
and U10197 (N_10197,N_5593,N_5681);
or U10198 (N_10198,N_8508,N_5932);
xor U10199 (N_10199,N_9118,N_9727);
nor U10200 (N_10200,N_9151,N_7559);
nor U10201 (N_10201,N_6564,N_7188);
and U10202 (N_10202,N_9893,N_6959);
xor U10203 (N_10203,N_9987,N_7403);
nand U10204 (N_10204,N_9210,N_7287);
nand U10205 (N_10205,N_5078,N_9308);
xnor U10206 (N_10206,N_8632,N_5384);
nor U10207 (N_10207,N_6093,N_7702);
nand U10208 (N_10208,N_5200,N_9314);
xnor U10209 (N_10209,N_7259,N_7939);
nand U10210 (N_10210,N_7609,N_7112);
nor U10211 (N_10211,N_5992,N_5142);
and U10212 (N_10212,N_6988,N_7224);
xnor U10213 (N_10213,N_7927,N_5143);
xor U10214 (N_10214,N_5567,N_5250);
and U10215 (N_10215,N_6012,N_5613);
and U10216 (N_10216,N_8147,N_8475);
xnor U10217 (N_10217,N_7719,N_8497);
nor U10218 (N_10218,N_5476,N_9839);
nor U10219 (N_10219,N_5899,N_7450);
nor U10220 (N_10220,N_5393,N_5721);
nand U10221 (N_10221,N_8562,N_5090);
xnor U10222 (N_10222,N_8964,N_7128);
xnor U10223 (N_10223,N_8340,N_5400);
nor U10224 (N_10224,N_8169,N_8323);
nor U10225 (N_10225,N_6163,N_9374);
nand U10226 (N_10226,N_5968,N_9148);
or U10227 (N_10227,N_5474,N_6300);
and U10228 (N_10228,N_6115,N_7021);
nor U10229 (N_10229,N_5108,N_8846);
nand U10230 (N_10230,N_9903,N_8227);
and U10231 (N_10231,N_9368,N_8790);
xnor U10232 (N_10232,N_8369,N_7350);
or U10233 (N_10233,N_8993,N_7020);
nor U10234 (N_10234,N_9373,N_9767);
nor U10235 (N_10235,N_6361,N_8156);
nand U10236 (N_10236,N_7688,N_9762);
xor U10237 (N_10237,N_7875,N_6753);
xnor U10238 (N_10238,N_8372,N_5915);
nor U10239 (N_10239,N_7878,N_7004);
or U10240 (N_10240,N_9045,N_9208);
xor U10241 (N_10241,N_7543,N_6089);
and U10242 (N_10242,N_9818,N_8728);
or U10243 (N_10243,N_9766,N_7373);
and U10244 (N_10244,N_8863,N_6624);
xor U10245 (N_10245,N_6146,N_7978);
or U10246 (N_10246,N_9559,N_6492);
nand U10247 (N_10247,N_8721,N_6500);
nor U10248 (N_10248,N_7881,N_6457);
nor U10249 (N_10249,N_6503,N_7109);
or U10250 (N_10250,N_8854,N_9026);
xor U10251 (N_10251,N_7126,N_6815);
and U10252 (N_10252,N_6397,N_8628);
and U10253 (N_10253,N_6133,N_6533);
or U10254 (N_10254,N_6252,N_9471);
nor U10255 (N_10255,N_8699,N_7518);
nor U10256 (N_10256,N_5436,N_5088);
nand U10257 (N_10257,N_5585,N_5064);
xnor U10258 (N_10258,N_7283,N_8787);
and U10259 (N_10259,N_9292,N_5928);
nand U10260 (N_10260,N_5385,N_9769);
nand U10261 (N_10261,N_9424,N_7605);
nand U10262 (N_10262,N_6985,N_8134);
and U10263 (N_10263,N_6324,N_7249);
or U10264 (N_10264,N_9078,N_6706);
nor U10265 (N_10265,N_8958,N_5347);
nand U10266 (N_10266,N_7062,N_6601);
nor U10267 (N_10267,N_5780,N_7553);
xor U10268 (N_10268,N_5818,N_8039);
nand U10269 (N_10269,N_7221,N_5554);
nand U10270 (N_10270,N_7846,N_8128);
and U10271 (N_10271,N_6856,N_8896);
or U10272 (N_10272,N_7208,N_7561);
nor U10273 (N_10273,N_5769,N_8664);
nor U10274 (N_10274,N_9153,N_9799);
and U10275 (N_10275,N_6145,N_7494);
or U10276 (N_10276,N_5318,N_7775);
nor U10277 (N_10277,N_8274,N_5890);
nand U10278 (N_10278,N_9719,N_5020);
and U10279 (N_10279,N_5715,N_9509);
xnor U10280 (N_10280,N_6201,N_6810);
nor U10281 (N_10281,N_6363,N_8347);
and U10282 (N_10282,N_6742,N_9108);
and U10283 (N_10283,N_5207,N_6812);
xor U10284 (N_10284,N_6264,N_5265);
nand U10285 (N_10285,N_5295,N_6045);
and U10286 (N_10286,N_5764,N_6376);
nor U10287 (N_10287,N_9920,N_7254);
and U10288 (N_10288,N_6308,N_7870);
nor U10289 (N_10289,N_9006,N_9518);
and U10290 (N_10290,N_9124,N_8501);
nor U10291 (N_10291,N_9001,N_7520);
xnor U10292 (N_10292,N_9333,N_8921);
nor U10293 (N_10293,N_9076,N_6210);
xnor U10294 (N_10294,N_6035,N_5130);
and U10295 (N_10295,N_5965,N_8224);
xor U10296 (N_10296,N_5988,N_8624);
xnor U10297 (N_10297,N_5542,N_8215);
nor U10298 (N_10298,N_7479,N_9475);
nor U10299 (N_10299,N_5927,N_9515);
or U10300 (N_10300,N_9710,N_6285);
or U10301 (N_10301,N_8641,N_9005);
xnor U10302 (N_10302,N_5367,N_5030);
xnor U10303 (N_10303,N_6479,N_7720);
xnor U10304 (N_10304,N_8404,N_8157);
or U10305 (N_10305,N_5536,N_6650);
or U10306 (N_10306,N_6509,N_6388);
or U10307 (N_10307,N_7839,N_8962);
or U10308 (N_10308,N_9089,N_7967);
nand U10309 (N_10309,N_8495,N_9028);
nand U10310 (N_10310,N_9500,N_8065);
nor U10311 (N_10311,N_5417,N_5051);
and U10312 (N_10312,N_7436,N_9327);
nor U10313 (N_10313,N_9395,N_6796);
or U10314 (N_10314,N_5598,N_8472);
xor U10315 (N_10315,N_8010,N_5722);
and U10316 (N_10316,N_7813,N_8410);
and U10317 (N_10317,N_9486,N_6256);
xor U10318 (N_10318,N_6545,N_6597);
or U10319 (N_10319,N_5670,N_8432);
or U10320 (N_10320,N_5955,N_9178);
or U10321 (N_10321,N_5221,N_5684);
nor U10322 (N_10322,N_5264,N_8353);
xnor U10323 (N_10323,N_7261,N_9582);
nor U10324 (N_10324,N_9999,N_5017);
nand U10325 (N_10325,N_5716,N_9971);
and U10326 (N_10326,N_8100,N_7376);
nand U10327 (N_10327,N_9978,N_6434);
and U10328 (N_10328,N_9309,N_5194);
and U10329 (N_10329,N_6424,N_6560);
and U10330 (N_10330,N_5491,N_9499);
nand U10331 (N_10331,N_5309,N_9567);
and U10332 (N_10332,N_6884,N_9157);
nor U10333 (N_10333,N_5177,N_6233);
nand U10334 (N_10334,N_9494,N_5768);
nand U10335 (N_10335,N_8277,N_7851);
nand U10336 (N_10336,N_7342,N_8578);
and U10337 (N_10337,N_7031,N_5014);
nand U10338 (N_10338,N_9495,N_8745);
nor U10339 (N_10339,N_7616,N_5519);
or U10340 (N_10340,N_6192,N_7765);
nor U10341 (N_10341,N_8346,N_9683);
nor U10342 (N_10342,N_8932,N_6693);
nor U10343 (N_10343,N_7116,N_9253);
xor U10344 (N_10344,N_6516,N_8672);
and U10345 (N_10345,N_9697,N_9502);
nor U10346 (N_10346,N_8556,N_9996);
nand U10347 (N_10347,N_9177,N_5408);
nand U10348 (N_10348,N_9159,N_5161);
xor U10349 (N_10349,N_9513,N_8831);
or U10350 (N_10350,N_8498,N_5827);
nor U10351 (N_10351,N_8592,N_7901);
xnor U10352 (N_10352,N_8987,N_9830);
nand U10353 (N_10353,N_5321,N_9144);
and U10354 (N_10354,N_5495,N_9347);
or U10355 (N_10355,N_9460,N_9859);
xor U10356 (N_10356,N_8526,N_7766);
and U10357 (N_10357,N_7424,N_9729);
or U10358 (N_10358,N_8923,N_7212);
or U10359 (N_10359,N_8373,N_7347);
and U10360 (N_10360,N_5713,N_9132);
nor U10361 (N_10361,N_5944,N_5676);
or U10362 (N_10362,N_5914,N_6406);
and U10363 (N_10363,N_8749,N_6475);
xnor U10364 (N_10364,N_6391,N_6371);
nor U10365 (N_10365,N_6108,N_8236);
and U10366 (N_10366,N_9861,N_5002);
or U10367 (N_10367,N_8757,N_5215);
xor U10368 (N_10368,N_9319,N_5821);
xor U10369 (N_10369,N_9597,N_7193);
xor U10370 (N_10370,N_8520,N_5869);
and U10371 (N_10371,N_9717,N_8310);
nand U10372 (N_10372,N_5139,N_8537);
nand U10373 (N_10373,N_7284,N_8967);
nor U10374 (N_10374,N_9700,N_8423);
xnor U10375 (N_10375,N_7301,N_9036);
xnor U10376 (N_10376,N_9320,N_9977);
xnor U10377 (N_10377,N_7988,N_6842);
nand U10378 (N_10378,N_5609,N_9875);
or U10379 (N_10379,N_5084,N_6752);
xnor U10380 (N_10380,N_9563,N_7289);
and U10381 (N_10381,N_9685,N_7977);
nor U10382 (N_10382,N_8217,N_8013);
or U10383 (N_10383,N_7189,N_6634);
and U10384 (N_10384,N_6850,N_7244);
xnor U10385 (N_10385,N_7574,N_5867);
nor U10386 (N_10386,N_5277,N_6058);
and U10387 (N_10387,N_7902,N_6521);
nor U10388 (N_10388,N_7969,N_6798);
xnor U10389 (N_10389,N_7461,N_6907);
nand U10390 (N_10390,N_7708,N_8853);
nor U10391 (N_10391,N_8237,N_9535);
xor U10392 (N_10392,N_8581,N_8160);
xor U10393 (N_10393,N_9295,N_8737);
nor U10394 (N_10394,N_9232,N_8770);
nor U10395 (N_10395,N_6255,N_9321);
or U10396 (N_10396,N_7155,N_6909);
nand U10397 (N_10397,N_6121,N_5949);
or U10398 (N_10398,N_5106,N_8148);
nand U10399 (N_10399,N_6134,N_9317);
nor U10400 (N_10400,N_8078,N_6226);
and U10401 (N_10401,N_5326,N_5437);
or U10402 (N_10402,N_7957,N_8575);
or U10403 (N_10403,N_9015,N_8397);
or U10404 (N_10404,N_7608,N_7197);
nor U10405 (N_10405,N_5578,N_8087);
nand U10406 (N_10406,N_6237,N_9081);
and U10407 (N_10407,N_7532,N_9443);
nand U10408 (N_10408,N_8239,N_9749);
and U10409 (N_10409,N_9902,N_5314);
xnor U10410 (N_10410,N_7084,N_7142);
and U10411 (N_10411,N_5748,N_6975);
and U10412 (N_10412,N_5343,N_8339);
nor U10413 (N_10413,N_9438,N_6681);
or U10414 (N_10414,N_5198,N_5462);
nand U10415 (N_10415,N_6809,N_5784);
and U10416 (N_10416,N_8132,N_8099);
nor U10417 (N_10417,N_9023,N_9464);
xnor U10418 (N_10418,N_6433,N_7325);
and U10419 (N_10419,N_6236,N_5414);
and U10420 (N_10420,N_7599,N_9901);
and U10421 (N_10421,N_8260,N_8555);
nor U10422 (N_10422,N_5816,N_8491);
nor U10423 (N_10423,N_8117,N_8341);
nand U10424 (N_10424,N_5972,N_8792);
nand U10425 (N_10425,N_6523,N_6642);
or U10426 (N_10426,N_9916,N_5705);
or U10427 (N_10427,N_9425,N_5558);
and U10428 (N_10428,N_7119,N_7997);
nor U10429 (N_10429,N_5370,N_9097);
nor U10430 (N_10430,N_7229,N_6281);
nand U10431 (N_10431,N_7898,N_8859);
nor U10432 (N_10432,N_8681,N_6531);
nor U10433 (N_10433,N_7986,N_9297);
nand U10434 (N_10434,N_9704,N_6334);
nor U10435 (N_10435,N_9249,N_7288);
nand U10436 (N_10436,N_8504,N_5921);
nor U10437 (N_10437,N_5649,N_9848);
or U10438 (N_10438,N_7487,N_5859);
nor U10439 (N_10439,N_8464,N_5870);
or U10440 (N_10440,N_5782,N_7865);
or U10441 (N_10441,N_6620,N_7275);
and U10442 (N_10442,N_5154,N_8158);
nand U10443 (N_10443,N_9549,N_8240);
or U10444 (N_10444,N_9399,N_7526);
or U10445 (N_10445,N_9586,N_6213);
and U10446 (N_10446,N_5683,N_8691);
xor U10447 (N_10447,N_7246,N_5092);
nor U10448 (N_10448,N_6898,N_9259);
xnor U10449 (N_10449,N_6766,N_5792);
and U10450 (N_10450,N_5937,N_7462);
and U10451 (N_10451,N_5892,N_8208);
nand U10452 (N_10452,N_9541,N_7899);
nand U10453 (N_10453,N_6048,N_6645);
nand U10454 (N_10454,N_9034,N_6558);
xnor U10455 (N_10455,N_6891,N_6976);
nand U10456 (N_10456,N_7161,N_5605);
xor U10457 (N_10457,N_8803,N_9270);
or U10458 (N_10458,N_9666,N_9103);
and U10459 (N_10459,N_5112,N_5357);
nand U10460 (N_10460,N_8259,N_8095);
nor U10461 (N_10461,N_9525,N_7515);
xnor U10462 (N_10462,N_5018,N_5538);
and U10463 (N_10463,N_5745,N_8700);
nand U10464 (N_10464,N_7756,N_8058);
nor U10465 (N_10465,N_5785,N_5740);
or U10466 (N_10466,N_8285,N_5588);
nor U10467 (N_10467,N_9083,N_9128);
and U10468 (N_10468,N_6218,N_7832);
nor U10469 (N_10469,N_8695,N_9018);
or U10470 (N_10470,N_9622,N_9119);
or U10471 (N_10471,N_7299,N_6055);
or U10472 (N_10472,N_8143,N_6392);
or U10473 (N_10473,N_9516,N_5455);
nand U10474 (N_10474,N_7575,N_5043);
nand U10475 (N_10475,N_8084,N_8380);
or U10476 (N_10476,N_8789,N_6339);
nand U10477 (N_10477,N_6395,N_6360);
nand U10478 (N_10478,N_9141,N_7476);
nand U10479 (N_10479,N_7660,N_8591);
nand U10480 (N_10480,N_5527,N_6724);
xor U10481 (N_10481,N_6172,N_5435);
xor U10482 (N_10482,N_8431,N_9215);
and U10483 (N_10483,N_9928,N_5879);
nor U10484 (N_10484,N_8338,N_7573);
or U10485 (N_10485,N_9998,N_6946);
or U10486 (N_10486,N_9049,N_6587);
xnor U10487 (N_10487,N_7625,N_7538);
nor U10488 (N_10488,N_9853,N_5736);
nor U10489 (N_10489,N_7032,N_9162);
or U10490 (N_10490,N_8956,N_7859);
or U10491 (N_10491,N_5443,N_8370);
nand U10492 (N_10492,N_8783,N_7781);
nor U10493 (N_10493,N_8509,N_5283);
and U10494 (N_10494,N_5333,N_9310);
or U10495 (N_10495,N_8206,N_7941);
and U10496 (N_10496,N_7430,N_5048);
xor U10497 (N_10497,N_5286,N_5783);
nand U10498 (N_10498,N_6905,N_8389);
nand U10499 (N_10499,N_7747,N_7406);
nor U10500 (N_10500,N_7524,N_8873);
nor U10501 (N_10501,N_7621,N_8383);
and U10502 (N_10502,N_5948,N_6876);
xnor U10503 (N_10503,N_5072,N_7519);
xnor U10504 (N_10504,N_7809,N_6819);
nand U10505 (N_10505,N_8442,N_7340);
nor U10506 (N_10506,N_6132,N_7968);
xnor U10507 (N_10507,N_5421,N_5961);
or U10508 (N_10508,N_5381,N_9279);
nand U10509 (N_10509,N_6969,N_5186);
xor U10510 (N_10510,N_5813,N_5619);
nand U10511 (N_10511,N_7334,N_7956);
and U10512 (N_10512,N_9620,N_5185);
nor U10513 (N_10513,N_9179,N_7278);
nor U10514 (N_10514,N_7071,N_8769);
nand U10515 (N_10515,N_7670,N_5604);
and U10516 (N_10516,N_9139,N_6152);
nor U10517 (N_10517,N_8225,N_5906);
xnor U10518 (N_10518,N_8382,N_9820);
nor U10519 (N_10519,N_6384,N_7404);
and U10520 (N_10520,N_8516,N_9676);
or U10521 (N_10521,N_5981,N_9615);
and U10522 (N_10522,N_5982,N_7190);
xnor U10523 (N_10523,N_5823,N_9504);
or U10524 (N_10524,N_9069,N_7607);
nand U10525 (N_10525,N_6862,N_8563);
nand U10526 (N_10526,N_8616,N_6278);
xnor U10527 (N_10527,N_5853,N_8546);
nor U10528 (N_10528,N_6268,N_6426);
and U10529 (N_10529,N_8436,N_6124);
xnor U10530 (N_10530,N_5373,N_7011);
nor U10531 (N_10531,N_8096,N_6117);
nand U10532 (N_10532,N_5205,N_6202);
nor U10533 (N_10533,N_9812,N_7752);
and U10534 (N_10534,N_8933,N_9883);
nor U10535 (N_10535,N_7316,N_5640);
and U10536 (N_10536,N_9573,N_9756);
and U10537 (N_10537,N_8909,N_6610);
nand U10538 (N_10538,N_5548,N_6331);
and U10539 (N_10539,N_9680,N_9432);
nand U10540 (N_10540,N_8210,N_9422);
nand U10541 (N_10541,N_8673,N_7646);
and U10542 (N_10542,N_9572,N_6465);
nor U10543 (N_10543,N_6594,N_9732);
nor U10544 (N_10544,N_9370,N_7952);
nand U10545 (N_10545,N_5446,N_6079);
xnor U10546 (N_10546,N_6276,N_7245);
nor U10547 (N_10547,N_5913,N_6524);
nor U10548 (N_10548,N_7755,N_6232);
nor U10549 (N_10549,N_6649,N_8955);
nor U10550 (N_10550,N_9950,N_6818);
and U10551 (N_10551,N_5695,N_7564);
xnor U10552 (N_10552,N_9129,N_7086);
and U10553 (N_10553,N_6925,N_9712);
nand U10554 (N_10554,N_7160,N_9599);
or U10555 (N_10555,N_6284,N_6801);
and U10556 (N_10556,N_7576,N_6389);
xor U10557 (N_10557,N_6217,N_5448);
nor U10558 (N_10558,N_8758,N_6670);
nand U10559 (N_10559,N_8828,N_7731);
or U10560 (N_10560,N_9705,N_8189);
nor U10561 (N_10561,N_6788,N_8936);
and U10562 (N_10562,N_5902,N_9689);
xor U10563 (N_10563,N_8503,N_5268);
nor U10564 (N_10564,N_6086,N_5338);
and U10565 (N_10565,N_5195,N_9944);
and U10566 (N_10566,N_6051,N_5855);
nor U10567 (N_10567,N_6193,N_7821);
nor U10568 (N_10568,N_5799,N_9277);
nand U10569 (N_10569,N_9064,N_9536);
or U10570 (N_10570,N_9918,N_7555);
nor U10571 (N_10571,N_9736,N_5581);
and U10572 (N_10572,N_6143,N_5365);
xor U10573 (N_10573,N_9854,N_7321);
or U10574 (N_10574,N_9892,N_8890);
nand U10575 (N_10575,N_7184,N_7954);
nand U10576 (N_10576,N_7971,N_9477);
nor U10577 (N_10577,N_9810,N_8401);
or U10578 (N_10578,N_9647,N_8917);
and U10579 (N_10579,N_9329,N_5865);
nor U10580 (N_10580,N_6080,N_8199);
xor U10581 (N_10581,N_6190,N_5594);
xor U10582 (N_10582,N_8659,N_8103);
nor U10583 (N_10583,N_6609,N_5524);
and U10584 (N_10584,N_9929,N_7921);
nor U10585 (N_10585,N_6077,N_9577);
xor U10586 (N_10586,N_7595,N_5405);
nor U10587 (N_10587,N_5663,N_9470);
xnor U10588 (N_10588,N_6345,N_9059);
nand U10589 (N_10589,N_9364,N_5643);
nand U10590 (N_10590,N_6957,N_5717);
nand U10591 (N_10591,N_7219,N_8793);
xnor U10592 (N_10592,N_9665,N_6544);
xnor U10593 (N_10593,N_8056,N_7199);
and U10594 (N_10594,N_7394,N_6916);
nor U10595 (N_10595,N_9166,N_9053);
xor U10596 (N_10596,N_6427,N_6663);
or U10597 (N_10597,N_5582,N_5229);
or U10598 (N_10598,N_7148,N_6541);
and U10599 (N_10599,N_9927,N_8319);
and U10600 (N_10600,N_6203,N_8415);
xor U10601 (N_10601,N_9757,N_9501);
or U10602 (N_10602,N_5817,N_8881);
xnor U10603 (N_10603,N_8427,N_6404);
or U10604 (N_10604,N_7087,N_7154);
and U10605 (N_10605,N_8408,N_8183);
nand U10606 (N_10606,N_7281,N_9488);
xnor U10607 (N_10607,N_9008,N_9337);
nand U10608 (N_10608,N_9205,N_9238);
xnor U10609 (N_10609,N_6254,N_8988);
and U10610 (N_10610,N_7606,N_9307);
nand U10611 (N_10611,N_9881,N_8075);
and U10612 (N_10612,N_6748,N_9925);
nand U10613 (N_10613,N_7276,N_8387);
nand U10614 (N_10614,N_5747,N_5611);
nor U10615 (N_10615,N_9539,N_9446);
xor U10616 (N_10616,N_8586,N_7723);
nand U10617 (N_10617,N_6407,N_5260);
or U10618 (N_10618,N_6902,N_5127);
nand U10619 (N_10619,N_8732,N_6241);
and U10620 (N_10620,N_6656,N_6795);
or U10621 (N_10621,N_7651,N_8015);
and U10622 (N_10622,N_8646,N_7628);
nand U10623 (N_10623,N_6896,N_8292);
xnor U10624 (N_10624,N_7850,N_6150);
xnor U10625 (N_10625,N_5403,N_5341);
nor U10626 (N_10626,N_9593,N_5151);
and U10627 (N_10627,N_8214,N_9585);
nor U10628 (N_10628,N_7074,N_6159);
and U10629 (N_10629,N_7114,N_7678);
nand U10630 (N_10630,N_5997,N_7243);
nor U10631 (N_10631,N_6118,N_5591);
nor U10632 (N_10632,N_5415,N_9519);
nor U10633 (N_10633,N_8906,N_9899);
xor U10634 (N_10634,N_6437,N_6599);
nand U10635 (N_10635,N_5905,N_6813);
nand U10636 (N_10636,N_5526,N_9764);
nor U10637 (N_10637,N_8037,N_5039);
nand U10638 (N_10638,N_8251,N_9796);
xor U10639 (N_10639,N_8451,N_7268);
or U10640 (N_10640,N_8266,N_8035);
or U10641 (N_10641,N_9027,N_6675);
and U10642 (N_10642,N_9592,N_6928);
nor U10643 (N_10643,N_6488,N_5241);
and U10644 (N_10644,N_6992,N_9560);
xor U10645 (N_10645,N_9019,N_5395);
nand U10646 (N_10646,N_9428,N_9581);
and U10647 (N_10647,N_8879,N_9196);
and U10648 (N_10648,N_6141,N_8488);
or U10649 (N_10649,N_7295,N_6183);
or U10650 (N_10650,N_6009,N_6915);
or U10651 (N_10651,N_9117,N_9113);
or U10652 (N_10652,N_5871,N_6296);
xor U10653 (N_10653,N_8647,N_7689);
nand U10654 (N_10654,N_5391,N_7203);
xor U10655 (N_10655,N_5293,N_7959);
nand U10656 (N_10656,N_5958,N_6554);
or U10657 (N_10657,N_8193,N_8760);
nor U10658 (N_10658,N_7408,N_7571);
or U10659 (N_10659,N_6350,N_7010);
and U10660 (N_10660,N_9138,N_8360);
and U10661 (N_10661,N_9442,N_5202);
or U10662 (N_10662,N_6478,N_8109);
or U10663 (N_10663,N_8621,N_8460);
and U10664 (N_10664,N_8384,N_7691);
or U10665 (N_10665,N_5144,N_9913);
and U10666 (N_10666,N_8742,N_7568);
xor U10667 (N_10667,N_8860,N_7964);
nor U10668 (N_10668,N_8663,N_5406);
or U10669 (N_10669,N_5819,N_6069);
nand U10670 (N_10670,N_7162,N_9773);
nand U10671 (N_10671,N_6804,N_7987);
nand U10672 (N_10672,N_8309,N_5298);
and U10673 (N_10673,N_5361,N_6563);
xor U10674 (N_10674,N_9361,N_5118);
and U10675 (N_10675,N_8200,N_6725);
nor U10676 (N_10676,N_9720,N_5145);
xor U10677 (N_10677,N_7787,N_7294);
nand U10678 (N_10678,N_9983,N_9220);
xnor U10679 (N_10679,N_5085,N_9823);
nand U10680 (N_10680,N_5532,N_6184);
nand U10681 (N_10681,N_6621,N_5477);
nor U10682 (N_10682,N_5995,N_8538);
and U10683 (N_10683,N_5042,N_9404);
and U10684 (N_10684,N_9211,N_6897);
or U10685 (N_10685,N_6738,N_8335);
nor U10686 (N_10686,N_7547,N_9264);
xnor U10687 (N_10687,N_8949,N_9052);
nand U10688 (N_10688,N_7319,N_5539);
nor U10689 (N_10689,N_8651,N_7483);
and U10690 (N_10690,N_8097,N_8784);
nor U10691 (N_10691,N_5552,N_5113);
and U10692 (N_10692,N_5730,N_7700);
nand U10693 (N_10693,N_9529,N_8031);
or U10694 (N_10694,N_8175,N_5376);
nor U10695 (N_10695,N_6655,N_9239);
nor U10696 (N_10696,N_8864,N_8568);
nand U10697 (N_10697,N_5320,N_9163);
or U10698 (N_10698,N_5401,N_9561);
nor U10699 (N_10699,N_5006,N_9418);
or U10700 (N_10700,N_9497,N_7603);
nor U10701 (N_10701,N_6831,N_9072);
nor U10702 (N_10702,N_7466,N_6761);
or U10703 (N_10703,N_5452,N_9885);
or U10704 (N_10704,N_7758,N_7655);
nor U10705 (N_10705,N_5848,N_6783);
nor U10706 (N_10706,N_9686,N_6030);
xor U10707 (N_10707,N_9631,N_5978);
nor U10708 (N_10708,N_7579,N_6440);
or U10709 (N_10709,N_5273,N_6793);
xnor U10710 (N_10710,N_5525,N_9578);
or U10711 (N_10711,N_9652,N_8337);
and U10712 (N_10712,N_7434,N_7551);
nor U10713 (N_10713,N_9387,N_7435);
nor U10714 (N_10714,N_8907,N_5121);
or U10715 (N_10715,N_6158,N_9485);
nor U10716 (N_10716,N_5544,N_9047);
xnor U10717 (N_10717,N_6510,N_5334);
and U10718 (N_10718,N_7849,N_9247);
or U10719 (N_10719,N_7297,N_5975);
nand U10720 (N_10720,N_9669,N_9594);
nand U10721 (N_10721,N_5111,N_7282);
nor U10722 (N_10722,N_9734,N_5924);
nor U10723 (N_10723,N_7310,N_5274);
or U10724 (N_10724,N_5930,N_7273);
nand U10725 (N_10725,N_5840,N_8634);
nand U10726 (N_10726,N_6338,N_9234);
or U10727 (N_10727,N_5576,N_8714);
nor U10728 (N_10728,N_9445,N_5698);
and U10729 (N_10729,N_6851,N_8692);
nor U10730 (N_10730,N_8868,N_5101);
nor U10731 (N_10731,N_8247,N_9068);
xnor U10732 (N_10732,N_9679,N_6882);
nor U10733 (N_10733,N_8852,N_6169);
or U10734 (N_10734,N_7492,N_6374);
or U10735 (N_10735,N_6947,N_6864);
nor U10736 (N_10736,N_5592,N_8751);
and U10737 (N_10737,N_9115,N_8059);
nor U10738 (N_10738,N_8965,N_9240);
and U10739 (N_10739,N_6066,N_8235);
nor U10740 (N_10740,N_8957,N_5315);
xnor U10741 (N_10741,N_7973,N_5966);
nand U10742 (N_10742,N_8939,N_9506);
nor U10743 (N_10743,N_5657,N_5079);
nand U10744 (N_10744,N_8006,N_7405);
or U10745 (N_10745,N_8990,N_8130);
or U10746 (N_10746,N_9057,N_5918);
or U10747 (N_10747,N_9376,N_5864);
nand U10748 (N_10748,N_8474,N_6668);
nor U10749 (N_10749,N_9909,N_7118);
and U10750 (N_10750,N_7737,N_8938);
xor U10751 (N_10751,N_8257,N_5999);
or U10752 (N_10752,N_6180,N_7721);
xor U10753 (N_10753,N_5132,N_9396);
xnor U10754 (N_10754,N_9698,N_5956);
nand U10755 (N_10755,N_7734,N_7175);
nor U10756 (N_10756,N_8226,N_6722);
or U10757 (N_10757,N_9643,N_6176);
xnor U10758 (N_10758,N_7008,N_5175);
nor U10759 (N_10759,N_7653,N_9988);
nor U10760 (N_10760,N_6325,N_8234);
or U10761 (N_10761,N_5601,N_9617);
and U10762 (N_10762,N_7361,N_9298);
nand U10763 (N_10763,N_7788,N_6442);
nand U10764 (N_10764,N_9725,N_6718);
nor U10765 (N_10765,N_6964,N_7317);
nor U10766 (N_10766,N_6847,N_6084);
or U10767 (N_10767,N_8839,N_7996);
nor U10768 (N_10768,N_6050,N_5873);
and U10769 (N_10769,N_6240,N_7391);
nor U10770 (N_10770,N_6449,N_5711);
nand U10771 (N_10771,N_7449,N_6242);
xor U10772 (N_10772,N_5431,N_5310);
or U10773 (N_10773,N_6480,N_5678);
nor U10774 (N_10774,N_9283,N_6918);
nor U10775 (N_10775,N_9203,N_5117);
and U10776 (N_10776,N_6416,N_6157);
nand U10777 (N_10777,N_9480,N_6848);
nor U10778 (N_10778,N_8612,N_8043);
nor U10779 (N_10779,N_6933,N_5296);
or U10780 (N_10780,N_7277,N_8178);
and U10781 (N_10781,N_7773,N_5487);
or U10782 (N_10782,N_8166,N_8593);
nor U10783 (N_10783,N_7043,N_8090);
nand U10784 (N_10784,N_9741,N_5521);
or U10785 (N_10785,N_8280,N_9199);
nor U10786 (N_10786,N_8348,N_8551);
or U10787 (N_10787,N_6177,N_7643);
or U10788 (N_10788,N_8899,N_9692);
nand U10789 (N_10789,N_6776,N_5157);
and U10790 (N_10790,N_6341,N_8637);
or U10791 (N_10791,N_9408,N_6173);
nor U10792 (N_10792,N_8232,N_5095);
nand U10793 (N_10793,N_5882,N_6455);
xor U10794 (N_10794,N_7830,N_9575);
or U10795 (N_10795,N_8118,N_5047);
and U10796 (N_10796,N_6661,N_7742);
nor U10797 (N_10797,N_8848,N_7381);
and U10798 (N_10798,N_8393,N_7304);
nor U10799 (N_10799,N_5007,N_5618);
and U10800 (N_10800,N_7038,N_8565);
nor U10801 (N_10801,N_6487,N_7654);
nand U10802 (N_10802,N_6073,N_5647);
xor U10803 (N_10803,N_9623,N_6310);
nand U10804 (N_10804,N_7622,N_8082);
nand U10805 (N_10805,N_6489,N_5138);
nand U10806 (N_10806,N_8151,N_6097);
nand U10807 (N_10807,N_6188,N_6153);
nand U10808 (N_10808,N_5565,N_7920);
nand U10809 (N_10809,N_8445,N_6092);
xor U10810 (N_10810,N_8477,N_9947);
or U10811 (N_10811,N_8468,N_5919);
xnor U10812 (N_10812,N_7728,N_8493);
and U10813 (N_10813,N_9569,N_7054);
xor U10814 (N_10814,N_9849,N_6777);
xor U10815 (N_10815,N_5858,N_6627);
xor U10816 (N_10816,N_6987,N_8916);
xnor U10817 (N_10817,N_6405,N_9032);
and U10818 (N_10818,N_8448,N_9570);
and U10819 (N_10819,N_8676,N_8482);
or U10820 (N_10820,N_9372,N_7615);
nand U10821 (N_10821,N_7771,N_7783);
or U10822 (N_10822,N_8252,N_6782);
and U10823 (N_10823,N_6393,N_5248);
or U10824 (N_10824,N_9478,N_6608);
or U10825 (N_10825,N_9325,N_9212);
or U10826 (N_10826,N_7762,N_9579);
or U10827 (N_10827,N_8499,N_6013);
or U10828 (N_10828,N_5786,N_5471);
nand U10829 (N_10829,N_6282,N_7928);
or U10830 (N_10830,N_6730,N_7588);
xnor U10831 (N_10831,N_6504,N_7422);
and U10832 (N_10832,N_5189,N_7751);
nor U10833 (N_10833,N_8576,N_8326);
nand U10834 (N_10834,N_8441,N_9224);
and U10835 (N_10835,N_6020,N_9548);
nand U10836 (N_10836,N_5522,N_5288);
nor U10837 (N_10837,N_6468,N_8307);
or U10838 (N_10838,N_5697,N_9798);
xor U10839 (N_10839,N_5622,N_5779);
nor U10840 (N_10840,N_9044,N_5206);
nor U10841 (N_10841,N_5056,N_9538);
nand U10842 (N_10842,N_8689,N_6027);
and U10843 (N_10843,N_8920,N_9523);
nand U10844 (N_10844,N_6007,N_6682);
nand U10845 (N_10845,N_9152,N_7320);
nand U10846 (N_10846,N_9807,N_7872);
nor U10847 (N_10847,N_8595,N_8487);
or U10848 (N_10848,N_8736,N_7490);
and U10849 (N_10849,N_7232,N_5772);
and U10850 (N_10850,N_5872,N_7624);
or U10851 (N_10851,N_8069,N_6780);
nor U10852 (N_10852,N_7915,N_5426);
or U10853 (N_10853,N_6151,N_5809);
or U10854 (N_10854,N_6496,N_8284);
nor U10855 (N_10855,N_5854,N_8057);
xor U10856 (N_10856,N_7336,N_8211);
and U10857 (N_10857,N_8461,N_6983);
nand U10858 (N_10858,N_6733,N_8668);
nand U10859 (N_10859,N_5074,N_7465);
and U10860 (N_10860,N_5900,N_7026);
nand U10861 (N_10861,N_9462,N_5236);
xnor U10862 (N_10862,N_7383,N_9348);
and U10863 (N_10863,N_7395,N_8722);
nand U10864 (N_10864,N_9774,N_8998);
xor U10865 (N_10865,N_8731,N_7763);
or U10866 (N_10866,N_8855,N_9322);
nor U10867 (N_10867,N_8534,N_6859);
and U10868 (N_10868,N_6322,N_7631);
xnor U10869 (N_10869,N_7799,N_6836);
or U10870 (N_10870,N_8979,N_9972);
nor U10871 (N_10871,N_8897,N_5029);
and U10872 (N_10872,N_7049,N_5410);
and U10873 (N_10873,N_5896,N_7338);
nor U10874 (N_10874,N_9980,N_8145);
or U10875 (N_10875,N_8768,N_9430);
nand U10876 (N_10876,N_6756,N_5383);
and U10877 (N_10877,N_8081,N_6336);
and U10878 (N_10878,N_5661,N_9255);
and U10879 (N_10879,N_5123,N_5833);
or U10880 (N_10880,N_9745,N_9982);
and U10881 (N_10881,N_6977,N_5019);
or U10882 (N_10882,N_5881,N_6059);
nor U10883 (N_10883,N_9167,N_9884);
and U10884 (N_10884,N_6337,N_5034);
nand U10885 (N_10885,N_8729,N_8288);
or U10886 (N_10886,N_7152,N_6744);
nor U10887 (N_10887,N_5351,N_8544);
nor U10888 (N_10888,N_6955,N_7372);
or U10889 (N_10889,N_8449,N_9855);
nor U10890 (N_10890,N_8030,N_5492);
nor U10891 (N_10891,N_8900,N_9863);
or U10892 (N_10892,N_6368,N_9276);
nor U10893 (N_10893,N_5758,N_5091);
nand U10894 (N_10894,N_7895,N_6835);
nand U10895 (N_10895,N_6832,N_9805);
or U10896 (N_10896,N_7274,N_8696);
or U10897 (N_10897,N_8466,N_8602);
or U10898 (N_10898,N_7472,N_7879);
nor U10899 (N_10899,N_5430,N_6411);
and U10900 (N_10900,N_8876,N_8951);
xnor U10901 (N_10901,N_6366,N_8375);
nand U10902 (N_10902,N_7318,N_7414);
nand U10903 (N_10903,N_7604,N_9416);
xnor U10904 (N_10904,N_5081,N_5170);
or U10905 (N_10905,N_8527,N_8114);
and U10906 (N_10906,N_5237,N_6961);
nor U10907 (N_10907,N_7840,N_8934);
or U10908 (N_10908,N_6113,N_9121);
and U10909 (N_10909,N_6754,N_6306);
nor U10910 (N_10910,N_6220,N_6743);
or U10911 (N_10911,N_6569,N_9328);
nor U10912 (N_10912,N_6094,N_9637);
nand U10913 (N_10913,N_8597,N_6960);
xnor U10914 (N_10914,N_9949,N_6104);
nor U10915 (N_10915,N_6617,N_6616);
xor U10916 (N_10916,N_6447,N_6559);
and U10917 (N_10917,N_8741,N_7384);
nor U10918 (N_10918,N_9304,N_7669);
and U10919 (N_10919,N_7623,N_7352);
or U10920 (N_10920,N_9420,N_7542);
or U10921 (N_10921,N_9826,N_6063);
xor U10922 (N_10922,N_7556,N_7746);
nor U10923 (N_10923,N_5933,N_9751);
and U10924 (N_10924,N_5734,N_8044);
nand U10925 (N_10925,N_6290,N_8066);
and U10926 (N_10926,N_6592,N_6340);
nor U10927 (N_10927,N_5423,N_5908);
nor U10928 (N_10928,N_6049,N_9101);
xor U10929 (N_10929,N_6807,N_7570);
nor U10930 (N_10930,N_5600,N_7293);
nor U10931 (N_10931,N_9701,N_9457);
or U10932 (N_10932,N_5196,N_9230);
xnor U10933 (N_10933,N_6528,N_5337);
nand U10934 (N_10934,N_7083,N_8922);
and U10935 (N_10935,N_5790,N_7835);
or U10936 (N_10936,N_7429,N_6527);
or U10937 (N_10937,N_6344,N_9369);
nand U10938 (N_10938,N_6514,N_8480);
nand U10939 (N_10939,N_6615,N_9965);
nor U10940 (N_10940,N_7205,N_8774);
xnor U10941 (N_10941,N_6485,N_6603);
and U10942 (N_10942,N_9024,N_6652);
nor U10943 (N_10943,N_8912,N_8141);
nor U10944 (N_10944,N_6588,N_5562);
nor U10945 (N_10945,N_8822,N_5572);
and U10946 (N_10946,N_5159,N_7217);
xnor U10947 (N_10947,N_9964,N_7565);
or U10948 (N_10948,N_8983,N_6292);
or U10949 (N_10949,N_6224,N_7066);
nand U10950 (N_10950,N_6840,N_7907);
and U10951 (N_10951,N_9181,N_5916);
nor U10952 (N_10952,N_5841,N_9312);
nor U10953 (N_10953,N_8708,N_8106);
and U10954 (N_10954,N_7739,N_8834);
nand U10955 (N_10955,N_6702,N_7369);
xor U10956 (N_10956,N_5584,N_9435);
nor U10957 (N_10957,N_7572,N_9721);
nor U10958 (N_10958,N_5387,N_5319);
nand U10959 (N_10959,N_7844,N_9930);
or U10960 (N_10960,N_8469,N_6515);
nand U10961 (N_10961,N_6482,N_5699);
or U10962 (N_10962,N_6827,N_7124);
nor U10963 (N_10963,N_5829,N_6768);
nor U10964 (N_10964,N_9379,N_5685);
nand U10965 (N_10965,N_6140,N_8888);
nand U10966 (N_10966,N_9986,N_7852);
xor U10967 (N_10967,N_6265,N_5671);
nor U10968 (N_10968,N_7585,N_6529);
nor U10969 (N_10969,N_8413,N_5146);
and U10970 (N_10970,N_8666,N_9145);
nand U10971 (N_10971,N_5861,N_9703);
nand U10972 (N_10972,N_9194,N_6472);
and U10973 (N_10973,N_9236,N_5287);
and U10974 (N_10974,N_8119,N_5067);
xor U10975 (N_10975,N_9846,N_8935);
xnor U10976 (N_10976,N_8992,N_9954);
and U10977 (N_10977,N_8943,N_9781);
or U10978 (N_10978,N_7485,N_6923);
xnor U10979 (N_10979,N_7251,N_5061);
or U10980 (N_10980,N_6130,N_9095);
xor U10981 (N_10981,N_6390,N_6333);
nand U10982 (N_10982,N_9588,N_7888);
nand U10983 (N_10983,N_6474,N_6223);
xnor U10984 (N_10984,N_7469,N_5004);
xor U10985 (N_10985,N_7767,N_8173);
and U10986 (N_10986,N_9524,N_9706);
nand U10987 (N_10987,N_6708,N_8281);
nor U10988 (N_10988,N_5602,N_8759);
and U10989 (N_10989,N_6273,N_5468);
nand U10990 (N_10990,N_5703,N_9932);
and U10991 (N_10991,N_6358,N_8658);
xnor U10992 (N_10992,N_7842,N_8571);
or U10993 (N_10993,N_9218,N_6934);
xnor U10994 (N_10994,N_7311,N_9790);
and U10995 (N_10995,N_5330,N_7019);
nand U10996 (N_10996,N_9109,N_7962);
nor U10997 (N_10997,N_6346,N_8963);
or U10998 (N_10998,N_6316,N_8600);
nor U10999 (N_10999,N_5093,N_6222);
or U11000 (N_11000,N_9168,N_8541);
or U11001 (N_11001,N_5313,N_8980);
or U11002 (N_11002,N_7632,N_6209);
xor U11003 (N_11003,N_5925,N_6070);
nor U11004 (N_11004,N_8098,N_7167);
and U11005 (N_11005,N_9605,N_7909);
and U11006 (N_11006,N_8776,N_7242);
and U11007 (N_11007,N_7502,N_5439);
nor U11008 (N_11008,N_6135,N_9591);
or U11009 (N_11009,N_8355,N_7171);
xor U11010 (N_11010,N_8627,N_8414);
nor U11011 (N_11011,N_8007,N_5725);
and U11012 (N_11012,N_5125,N_7501);
or U11013 (N_11013,N_5016,N_5197);
nand U11014 (N_11014,N_5339,N_9970);
or U11015 (N_11015,N_7300,N_5304);
and U11016 (N_11016,N_8762,N_9228);
nor U11017 (N_11017,N_7214,N_5355);
nor U11018 (N_11018,N_9037,N_7009);
and U11019 (N_11019,N_7444,N_5946);
xor U11020 (N_11020,N_8465,N_6654);
and U11021 (N_11021,N_9493,N_5141);
nand U11022 (N_11022,N_7495,N_8456);
nor U11023 (N_11023,N_6863,N_7847);
and U11024 (N_11024,N_7057,N_7701);
and U11025 (N_11025,N_5561,N_9087);
or U11026 (N_11026,N_9726,N_8778);
nand U11027 (N_11027,N_5520,N_7816);
nor U11028 (N_11028,N_7007,N_9134);
nand U11029 (N_11029,N_7508,N_7894);
nor U11030 (N_11030,N_9331,N_9343);
nor U11031 (N_11031,N_8086,N_7706);
and U11032 (N_11032,N_9007,N_5291);
nor U11033 (N_11033,N_6741,N_9624);
xor U11034 (N_11034,N_8928,N_9537);
or U11035 (N_11035,N_6467,N_7150);
xor U11036 (N_11036,N_8314,N_6944);
and U11037 (N_11037,N_5233,N_8910);
nand U11038 (N_11038,N_9252,N_9071);
xnor U11039 (N_11039,N_7201,N_6382);
nand U11040 (N_11040,N_6996,N_6525);
nand U11041 (N_11041,N_6552,N_6567);
or U11042 (N_11042,N_6512,N_9063);
and U11043 (N_11043,N_6838,N_7705);
or U11044 (N_11044,N_5227,N_6206);
nor U11045 (N_11045,N_7530,N_9459);
nand U11046 (N_11046,N_8278,N_8690);
nand U11047 (N_11047,N_9360,N_8654);
nand U11048 (N_11048,N_7808,N_8807);
xor U11049 (N_11049,N_5432,N_5050);
nor U11050 (N_11050,N_6506,N_7877);
nand U11051 (N_11051,N_7090,N_8064);
xnor U11052 (N_11052,N_5497,N_5316);
and U11053 (N_11053,N_9663,N_6110);
nor U11054 (N_11054,N_6526,N_8519);
nor U11055 (N_11055,N_6805,N_6362);
nand U11056 (N_11056,N_6638,N_8424);
xnor U11057 (N_11057,N_9936,N_9758);
and U11058 (N_11058,N_7002,N_8352);
xor U11059 (N_11059,N_9800,N_7818);
xnor U11060 (N_11060,N_9150,N_6486);
nor U11061 (N_11061,N_5606,N_8865);
xor U11062 (N_11062,N_6573,N_8567);
xnor U11063 (N_11063,N_9229,N_9123);
and U11064 (N_11064,N_5038,N_5033);
or U11065 (N_11065,N_9125,N_8648);
nor U11066 (N_11066,N_9862,N_7528);
nand U11067 (N_11067,N_9066,N_9958);
nor U11068 (N_11068,N_6227,N_6546);
or U11069 (N_11069,N_5834,N_6727);
and U11070 (N_11070,N_6041,N_8560);
or U11071 (N_11071,N_7437,N_8428);
nand U11072 (N_11072,N_9890,N_8688);
nor U11073 (N_11073,N_7337,N_6874);
and U11074 (N_11074,N_5743,N_5800);
nand U11075 (N_11075,N_5179,N_6033);
and U11076 (N_11076,N_5184,N_5270);
nand U11077 (N_11077,N_5089,N_9183);
nor U11078 (N_11078,N_5077,N_7068);
xnor U11079 (N_11079,N_9336,N_8874);
and U11080 (N_11080,N_5626,N_5156);
xnor U11081 (N_11081,N_8198,N_9431);
nor U11082 (N_11082,N_9213,N_8242);
and U11083 (N_11083,N_8312,N_9997);
or U11084 (N_11084,N_5115,N_7749);
nand U11085 (N_11085,N_7477,N_6814);
nand U11086 (N_11086,N_5502,N_9256);
nor U11087 (N_11087,N_5535,N_9911);
nor U11088 (N_11088,N_8635,N_8574);
nand U11089 (N_11089,N_9896,N_7247);
xnor U11090 (N_11090,N_5027,N_7861);
nor U11091 (N_11091,N_8182,N_8045);
nor U11092 (N_11092,N_7697,N_6230);
xor U11093 (N_11093,N_9484,N_7919);
or U11094 (N_11094,N_7510,N_8330);
or U11095 (N_11095,N_6982,N_9110);
xor U11096 (N_11096,N_9388,N_8364);
xor U11097 (N_11097,N_6820,N_5832);
xor U11098 (N_11098,N_8542,N_9910);
nand U11099 (N_11099,N_6373,N_5015);
xnor U11100 (N_11100,N_7963,N_6317);
xnor U11101 (N_11101,N_9250,N_9565);
and U11102 (N_11102,N_9254,N_6448);
nor U11103 (N_11103,N_5810,N_6978);
or U11104 (N_11104,N_5889,N_6539);
or U11105 (N_11105,N_5364,N_6721);
and U11106 (N_11106,N_9702,N_6762);
or U11107 (N_11107,N_8622,N_5754);
nand U11108 (N_11108,N_5041,N_8351);
and U11109 (N_11109,N_8530,N_5893);
nor U11110 (N_11110,N_6576,N_5063);
nor U11111 (N_11111,N_7690,N_5878);
nor U11112 (N_11112,N_5556,N_7991);
xnor U11113 (N_11113,N_9606,N_7042);
or U11114 (N_11114,N_6123,N_6394);
and U11115 (N_11115,N_8609,N_7078);
or U11116 (N_11116,N_6354,N_7499);
xor U11117 (N_11117,N_9054,N_8212);
or U11118 (N_11118,N_8400,N_7108);
or U11119 (N_11119,N_5648,N_7048);
xnor U11120 (N_11120,N_6800,N_5311);
and U11121 (N_11121,N_6412,N_6464);
xor U11122 (N_11122,N_6139,N_7211);
nand U11123 (N_11123,N_6785,N_8074);
nand U11124 (N_11124,N_5422,N_5305);
and U11125 (N_11125,N_9349,N_8794);
nand U11126 (N_11126,N_6910,N_9461);
nor U11127 (N_11127,N_7272,N_7136);
nand U11128 (N_11128,N_9187,N_6430);
and U11129 (N_11129,N_9724,N_6309);
xor U11130 (N_11130,N_7885,N_6746);
nand U11131 (N_11131,N_7034,N_7339);
or U11132 (N_11132,N_9632,N_9362);
nand U11133 (N_11133,N_9650,N_7252);
nor U11134 (N_11134,N_6100,N_6963);
nor U11135 (N_11135,N_6343,N_6830);
or U11136 (N_11136,N_9100,N_9571);
xor U11137 (N_11137,N_6414,N_8875);
nor U11138 (N_11138,N_6698,N_7481);
nor U11139 (N_11139,N_5603,N_7302);
or U11140 (N_11140,N_6870,N_8733);
nor U11141 (N_11141,N_6402,N_8893);
nand U11142 (N_11142,N_8545,N_9707);
and U11143 (N_11143,N_8286,N_5760);
nor U11144 (N_11144,N_8582,N_8061);
nor U11145 (N_11145,N_7562,N_9962);
nand U11146 (N_11146,N_5909,N_6769);
xor U11147 (N_11147,N_7024,N_5620);
and U11148 (N_11148,N_9828,N_6740);
or U11149 (N_11149,N_6453,N_5920);
nor U11150 (N_11150,N_9985,N_5765);
nor U11151 (N_11151,N_9483,N_9888);
xor U11152 (N_11152,N_5465,N_9904);
nor U11153 (N_11153,N_8886,N_7829);
xnor U11154 (N_11154,N_9681,N_8521);
and U11155 (N_11155,N_9576,N_8720);
nor U11156 (N_11156,N_8753,N_8902);
or U11157 (N_11157,N_9912,N_9690);
xor U11158 (N_11158,N_5852,N_8025);
and U11159 (N_11159,N_5345,N_7097);
nand U11160 (N_11160,N_9785,N_9742);
nand U11161 (N_11161,N_5850,N_8422);
nand U11162 (N_11162,N_6758,N_8561);
and U11163 (N_11163,N_7210,N_8344);
xor U11164 (N_11164,N_8919,N_6330);
xor U11165 (N_11165,N_8250,N_5806);
and U11166 (N_11166,N_6250,N_7966);
or U11167 (N_11167,N_7411,N_6799);
nor U11168 (N_11168,N_9434,N_6182);
or U11169 (N_11169,N_7323,N_5973);
nor U11170 (N_11170,N_8268,N_5583);
xnor U11171 (N_11171,N_9243,N_7385);
or U11172 (N_11172,N_7220,N_6685);
xor U11173 (N_11173,N_6720,N_5500);
or U11174 (N_11174,N_6156,N_6245);
nand U11175 (N_11175,N_9231,N_8892);
or U11176 (N_11176,N_7134,N_6379);
nand U11177 (N_11177,N_8041,N_7315);
xor U11178 (N_11178,N_6532,N_5342);
nor U11179 (N_11179,N_7550,N_8036);
nand U11180 (N_11180,N_6469,N_8034);
and U11181 (N_11181,N_5441,N_7464);
nand U11182 (N_11182,N_5505,N_9274);
nor U11183 (N_11183,N_5162,N_8618);
nor U11184 (N_11184,N_9301,N_5989);
xor U11185 (N_11185,N_9345,N_7231);
nor U11186 (N_11186,N_8153,N_5224);
nor U11187 (N_11187,N_8611,N_6990);
nor U11188 (N_11188,N_8564,N_5787);
xnor U11189 (N_11189,N_9778,N_6128);
nand U11190 (N_11190,N_7017,N_9269);
or U11191 (N_11191,N_9410,N_7416);
nand U11192 (N_11192,N_9801,N_8165);
and U11193 (N_11193,N_5488,N_8462);
or U11194 (N_11194,N_6637,N_7380);
and U11195 (N_11195,N_7786,N_7955);
or U11196 (N_11196,N_9695,N_5059);
or U11197 (N_11197,N_9546,N_6972);
and U11198 (N_11198,N_6772,N_9439);
or U11199 (N_11199,N_6833,N_5712);
or U11200 (N_11200,N_9667,N_8914);
and U11201 (N_11201,N_7792,N_5083);
nand U11202 (N_11202,N_5008,N_7094);
xnor U11203 (N_11203,N_9922,N_8771);
or U11204 (N_11204,N_8180,N_9225);
nand U11205 (N_11205,N_8818,N_9039);
nor U11206 (N_11206,N_9339,N_9598);
nor U11207 (N_11207,N_9363,N_7386);
xor U11208 (N_11208,N_7745,N_6712);
nand U11209 (N_11209,N_5183,N_7713);
xor U11210 (N_11210,N_5547,N_8290);
or U11211 (N_11211,N_5805,N_5035);
nand U11212 (N_11212,N_5245,N_6550);
xor U11213 (N_11213,N_7525,N_6879);
or U11214 (N_11214,N_5329,N_5891);
and U11215 (N_11215,N_5404,N_8438);
and U11216 (N_11216,N_7291,N_7375);
and U11217 (N_11217,N_9046,N_5706);
or U11218 (N_11218,N_9289,N_8850);
or U11219 (N_11219,N_7537,N_5182);
and U11220 (N_11220,N_6797,N_8172);
xor U11221 (N_11221,N_6014,N_7458);
or U11222 (N_11222,N_6660,N_8945);
nor U11223 (N_11223,N_6967,N_8554);
xnor U11224 (N_11224,N_8068,N_8052);
xor U11225 (N_11225,N_8655,N_8042);
nand U11226 (N_11226,N_5494,N_7729);
and U11227 (N_11227,N_6570,N_6991);
or U11228 (N_11228,N_8746,N_7306);
nor U11229 (N_11229,N_6646,N_6889);
xor U11230 (N_11230,N_7539,N_6431);
or U11231 (N_11231,N_5269,N_9744);
nor U11232 (N_11232,N_5874,N_9678);
nand U11233 (N_11233,N_9311,N_5011);
nor U11234 (N_11234,N_7234,N_8358);
and U11235 (N_11235,N_9190,N_9473);
xnor U11236 (N_11236,N_7827,N_7324);
xor U11237 (N_11237,N_7186,N_5942);
and U11238 (N_11238,N_8171,N_6709);
xor U11239 (N_11239,N_5894,N_5923);
nand U11240 (N_11240,N_6053,N_6631);
and U11241 (N_11241,N_5994,N_8374);
xor U11242 (N_11242,N_8872,N_5666);
xor U11243 (N_11243,N_8548,N_9452);
or U11244 (N_11244,N_7563,N_5506);
and U11245 (N_11245,N_5746,N_5453);
nand U11246 (N_11246,N_5243,N_8885);
nand U11247 (N_11247,N_5009,N_5463);
nor U11248 (N_11248,N_6403,N_8617);
or U11249 (N_11249,N_8587,N_5511);
and U11250 (N_11250,N_6950,N_9041);
nor U11251 (N_11251,N_5010,N_7279);
nor U11252 (N_11252,N_6680,N_7938);
nand U11253 (N_11253,N_9530,N_7358);
or U11254 (N_11254,N_5642,N_9604);
or U11255 (N_11255,N_8149,N_7419);
nor U11256 (N_11256,N_7934,N_5755);
nand U11257 (N_11257,N_5428,N_5363);
or U11258 (N_11258,N_9222,N_9968);
nor U11259 (N_11259,N_9380,N_8952);
and U11260 (N_11260,N_7129,N_9096);
nor U11261 (N_11261,N_5550,N_7453);
or U11262 (N_11262,N_7455,N_6399);
and U11263 (N_11263,N_9143,N_9429);
and U11264 (N_11264,N_7730,N_6239);
xnor U11265 (N_11265,N_6119,N_7627);
or U11266 (N_11266,N_9664,N_5073);
nor U11267 (N_11267,N_9346,N_5263);
nand U11268 (N_11268,N_8202,N_5420);
and U11269 (N_11269,N_5001,N_7743);
nand U11270 (N_11270,N_5637,N_9386);
nand U11271 (N_11271,N_8079,N_8221);
or U11272 (N_11272,N_6628,N_9894);
xor U11273 (N_11273,N_5586,N_6258);
nor U11274 (N_11274,N_6704,N_5013);
or U11275 (N_11275,N_5109,N_7351);
nor U11276 (N_11276,N_6719,N_9136);
xor U11277 (N_11277,N_8418,N_8392);
xor U11278 (N_11278,N_7794,N_6369);
nand U11279 (N_11279,N_9334,N_9815);
and U11280 (N_11280,N_9779,N_5350);
and U11281 (N_11281,N_6703,N_7016);
nor U11282 (N_11282,N_5577,N_7484);
xor U11283 (N_11283,N_9554,N_5427);
and U11284 (N_11284,N_8181,N_5075);
nand U11285 (N_11285,N_5060,N_6520);
xnor U11286 (N_11286,N_9512,N_5979);
and U11287 (N_11287,N_7138,N_8638);
nand U11288 (N_11288,N_5590,N_8233);
xor U11289 (N_11289,N_8801,N_7636);
nor U11290 (N_11290,N_8845,N_6678);
and U11291 (N_11291,N_8835,N_8391);
nand U11292 (N_11292,N_8867,N_6319);
nand U11293 (N_11293,N_8155,N_5412);
xnor U11294 (N_11294,N_6196,N_9527);
nand U11295 (N_11295,N_9367,N_9302);
and U11296 (N_11296,N_7760,N_5442);
xor U11297 (N_11297,N_7349,N_6713);
nand U11298 (N_11298,N_5568,N_8126);
nand U11299 (N_11299,N_9867,N_7353);
nand U11300 (N_11300,N_5457,N_5773);
or U11301 (N_11301,N_7522,N_5508);
and U11302 (N_11302,N_9383,N_9931);
nor U11303 (N_11303,N_9866,N_7474);
or U11304 (N_11304,N_8636,N_9029);
and U11305 (N_11305,N_6205,N_8911);
xor U11306 (N_11306,N_5798,N_6266);
xor U11307 (N_11307,N_9638,N_9286);
or U11308 (N_11308,N_5931,N_5665);
xnor U11309 (N_11309,N_5543,N_6566);
nand U11310 (N_11310,N_9456,N_6849);
or U11311 (N_11311,N_6845,N_8275);
xor U11312 (N_11312,N_7367,N_9808);
and U11313 (N_11313,N_5837,N_8317);
and U11314 (N_11314,N_7073,N_6816);
or U11315 (N_11315,N_8773,N_6422);
or U11316 (N_11316,N_6775,N_8009);
xnor U11317 (N_11317,N_7803,N_5797);
and U11318 (N_11318,N_9195,N_9722);
and U11319 (N_11319,N_7512,N_5857);
nor U11320 (N_11320,N_5723,N_5348);
nand U11321 (N_11321,N_6883,N_7012);
xor U11322 (N_11322,N_7478,N_6207);
nand U11323 (N_11323,N_7101,N_5533);
and U11324 (N_11324,N_7396,N_7946);
and U11325 (N_11325,N_5512,N_5053);
nand U11326 (N_11326,N_9048,N_5638);
nor U11327 (N_11327,N_7776,N_9608);
xnor U11328 (N_11328,N_9043,N_8531);
nor U11329 (N_11329,N_6687,N_5386);
nor U11330 (N_11330,N_5984,N_7230);
or U11331 (N_11331,N_8159,N_7673);
or U11332 (N_11332,N_6942,N_8788);
or U11333 (N_11333,N_8481,N_7102);
xnor U11334 (N_11334,N_7545,N_7439);
and U11335 (N_11335,N_5225,N_9305);
nor U11336 (N_11336,N_7926,N_6251);
or U11337 (N_11337,N_5302,N_9355);
and U11338 (N_11338,N_9498,N_7433);
nor U11339 (N_11339,N_5795,N_6562);
or U11340 (N_11340,N_8763,N_6262);
and U11341 (N_11341,N_5120,N_5501);
xor U11342 (N_11342,N_6781,N_7387);
nor U11343 (N_11343,N_6267,N_9832);
xnor U11344 (N_11344,N_6428,N_6011);
or U11345 (N_11345,N_7932,N_8777);
nand U11346 (N_11346,N_8190,N_7099);
xor U11347 (N_11347,N_7397,N_7910);
nor U11348 (N_11348,N_6318,N_8014);
and U11349 (N_11349,N_9122,N_7018);
or U11350 (N_11350,N_6040,N_7866);
and U11351 (N_11351,N_6595,N_7810);
nand U11352 (N_11352,N_7529,N_8566);
nor U11353 (N_11353,N_5574,N_8077);
xor U11354 (N_11354,N_7856,N_8623);
and U11355 (N_11355,N_5589,N_5983);
and U11356 (N_11356,N_9090,N_5110);
xnor U11357 (N_11357,N_5238,N_6415);
nor U11358 (N_11358,N_6861,N_9214);
or U11359 (N_11359,N_5555,N_8953);
xor U11360 (N_11360,N_5164,N_8607);
nand U11361 (N_11361,N_5911,N_7415);
nand U11362 (N_11362,N_5617,N_6938);
nor U11363 (N_11363,N_9403,N_9942);
nand U11364 (N_11364,N_5193,N_6257);
xor U11365 (N_11365,N_6860,N_7215);
and U11366 (N_11366,N_6676,N_9908);
xor U11367 (N_11367,N_9924,N_9671);
xor U11368 (N_11368,N_6095,N_8305);
and U11369 (N_11369,N_9092,N_9393);
nand U11370 (N_11370,N_8478,N_8115);
nand U11371 (N_11371,N_5275,N_7366);
xor U11372 (N_11372,N_8830,N_7257);
nand U11373 (N_11373,N_8533,N_5749);
nand U11374 (N_11374,N_7552,N_7482);
and U11375 (N_11375,N_8327,N_8377);
nand U11376 (N_11376,N_8754,N_5086);
xnor U11377 (N_11377,N_7418,N_9359);
nor U11378 (N_11378,N_7149,N_5630);
xor U11379 (N_11379,N_7185,N_7998);
nor U11380 (N_11380,N_9193,N_8131);
or U11381 (N_11381,N_7843,N_8177);
xor U11382 (N_11382,N_6166,N_6930);
or U11383 (N_11383,N_8176,N_6272);
xor U11384 (N_11384,N_8999,N_5469);
nand U11385 (N_11385,N_8619,N_7363);
nor U11386 (N_11386,N_5201,N_8289);
or U11387 (N_11387,N_5727,N_7075);
and U11388 (N_11388,N_8625,N_6530);
nand U11389 (N_11389,N_6837,N_6260);
nand U11390 (N_11390,N_7401,N_9630);
or U11391 (N_11391,N_9085,N_8334);
nor U11392 (N_11392,N_9189,N_5962);
xnor U11393 (N_11393,N_6004,N_7912);
or U11394 (N_11394,N_8539,N_5943);
and U11395 (N_11395,N_7891,N_7735);
nor U11396 (N_11396,N_6231,N_5036);
or U11397 (N_11397,N_8698,N_6101);
and U11398 (N_11398,N_8665,N_9267);
xor U11399 (N_11399,N_9198,N_8827);
and U11400 (N_11400,N_5633,N_8300);
or U11401 (N_11401,N_6470,N_5208);
or U11402 (N_11402,N_9318,N_6954);
or U11403 (N_11403,N_7014,N_5686);
or U11404 (N_11404,N_7637,N_6170);
nand U11405 (N_11405,N_9390,N_7491);
xor U11406 (N_11406,N_9952,N_5450);
and U11407 (N_11407,N_7815,N_9000);
and U11408 (N_11408,N_6953,N_8088);
and U11409 (N_11409,N_9761,N_6999);
nor U11410 (N_11410,N_8809,N_7438);
xnor U11411 (N_11411,N_6803,N_6456);
or U11412 (N_11412,N_6018,N_9246);
nor U11413 (N_11413,N_8606,N_5171);
xor U11414 (N_11414,N_9590,N_9182);
xnor U11415 (N_11415,N_5230,N_7237);
or U11416 (N_11416,N_8325,N_5770);
and U11417 (N_11417,N_9564,N_6022);
xnor U11418 (N_11418,N_9086,N_9677);
and U11419 (N_11419,N_8028,N_5884);
and U11420 (N_11420,N_5824,N_7127);
nor U11421 (N_11421,N_9842,N_8903);
nor U11422 (N_11422,N_6420,N_9200);
nand U11423 (N_11423,N_7382,N_8127);
nor U11424 (N_11424,N_6502,N_6419);
nor U11425 (N_11425,N_8216,N_7744);
or U11426 (N_11426,N_9356,N_5987);
nor U11427 (N_11427,N_6249,N_7423);
nand U11428 (N_11428,N_8229,N_9589);
xnor U11429 (N_11429,N_5461,N_9401);
and U11430 (N_11430,N_5667,N_6398);
or U11431 (N_11431,N_5165,N_6939);
nand U11432 (N_11432,N_8271,N_8256);
nor U11433 (N_11433,N_7994,N_6536);
nand U11434 (N_11434,N_7577,N_6283);
nor U11435 (N_11435,N_8331,N_8135);
nand U11436 (N_11436,N_8701,N_8549);
xnor U11437 (N_11437,N_7679,N_7793);
or U11438 (N_11438,N_8767,N_5733);
nand U11439 (N_11439,N_8811,N_5349);
nor U11440 (N_11440,N_9022,N_9873);
nor U11441 (N_11441,N_6607,N_7882);
nand U11442 (N_11442,N_5231,N_6081);
nand U11443 (N_11443,N_6356,N_9223);
and U11444 (N_11444,N_9675,N_8707);
or U11445 (N_11445,N_5838,N_5478);
xor U11446 (N_11446,N_6892,N_9753);
and U11447 (N_11447,N_7904,N_6071);
xor U11448 (N_11448,N_9551,N_6852);
xor U11449 (N_11449,N_8978,N_9817);
xor U11450 (N_11450,N_5028,N_7704);
xor U11451 (N_11451,N_9353,N_7033);
and U11452 (N_11452,N_8730,N_7855);
nor U11453 (N_11453,N_6981,N_9398);
nor U11454 (N_11454,N_8525,N_9437);
xnor U11455 (N_11455,N_6259,N_5941);
or U11456 (N_11456,N_9130,N_7269);
nand U11457 (N_11457,N_6122,N_7613);
nor U11458 (N_11458,N_5055,N_5353);
and U11459 (N_11459,N_7120,N_8806);
nand U11460 (N_11460,N_6238,N_5804);
nor U11461 (N_11461,N_8985,N_9142);
or U11462 (N_11462,N_9641,N_6043);
and U11463 (N_11463,N_9149,N_6657);
nor U11464 (N_11464,N_6518,N_9711);
or U11465 (N_11465,N_6779,N_6269);
or U11466 (N_11466,N_9562,N_7390);
or U11467 (N_11467,N_6823,N_7233);
nand U11468 (N_11468,N_9526,N_6802);
nor U11469 (N_11469,N_9540,N_7908);
nand U11470 (N_11470,N_6784,N_5636);
or U11471 (N_11471,N_7583,N_7178);
nand U11472 (N_11472,N_9723,N_8808);
nand U11473 (N_11473,N_7080,N_9137);
nand U11474 (N_11474,N_5767,N_8394);
or U11475 (N_11475,N_7567,N_5976);
or U11476 (N_11476,N_5285,N_7823);
nor U11477 (N_11477,N_7867,N_7013);
or U11478 (N_11478,N_8712,N_6204);
or U11479 (N_11479,N_6591,N_8675);
nor U11480 (N_11480,N_8050,N_5280);
nor U11481 (N_11481,N_8615,N_5580);
xnor U11482 (N_11482,N_8810,N_5148);
and U11483 (N_11483,N_7517,N_9945);
or U11484 (N_11484,N_9338,N_8915);
nand U11485 (N_11485,N_8870,N_6817);
xnor U11486 (N_11486,N_7527,N_9792);
and U11487 (N_11487,N_7164,N_9482);
nor U11488 (N_11488,N_6144,N_5340);
and U11489 (N_11489,N_7067,N_6214);
nor U11490 (N_11490,N_7667,N_9476);
or U11491 (N_11491,N_5392,N_5559);
xnor U11492 (N_11492,N_8693,N_5692);
xnor U11493 (N_11493,N_7753,N_6155);
xnor U11494 (N_11494,N_7088,N_6787);
or U11495 (N_11495,N_5219,N_9079);
or U11496 (N_11496,N_6328,N_8476);
xnor U11497 (N_11497,N_6534,N_9976);
nor U11498 (N_11498,N_8626,N_9209);
xor U11499 (N_11499,N_6715,N_9940);
nand U11500 (N_11500,N_7718,N_7498);
nor U11501 (N_11501,N_8884,N_8409);
xnor U11502 (N_11502,N_6690,N_7091);
xnor U11503 (N_11503,N_8089,N_5866);
or U11504 (N_11504,N_8507,N_5627);
xor U11505 (N_11505,N_9877,N_5153);
and U11506 (N_11506,N_5888,N_5458);
nor U11507 (N_11507,N_5675,N_7332);
or U11508 (N_11508,N_7093,N_9852);
nor U11509 (N_11509,N_9107,N_9140);
nor U11510 (N_11510,N_7389,N_9417);
xnor U11511 (N_11511,N_7768,N_6825);
nor U11512 (N_11512,N_5807,N_7591);
and U11513 (N_11513,N_5306,N_7110);
and U11514 (N_11514,N_9503,N_6686);
or U11515 (N_11515,N_8580,N_6994);
and U11516 (N_11516,N_8536,N_9611);
nor U11517 (N_11517,N_6359,N_5510);
xor U11518 (N_11518,N_5517,N_5700);
nor U11519 (N_11519,N_8573,N_8694);
nor U11520 (N_11520,N_7736,N_5459);
nand U11521 (N_11521,N_9973,N_7805);
xnor U11522 (N_11522,N_5220,N_8991);
nand U11523 (N_11523,N_7790,N_7264);
xor U11524 (N_11524,N_6640,N_8862);
xor U11525 (N_11525,N_9035,N_5595);
nor U11526 (N_11526,N_6571,N_6315);
nand U11527 (N_11527,N_9116,N_7132);
or U11528 (N_11528,N_6630,N_6865);
xor U11529 (N_11529,N_8656,N_6745);
xnor U11530 (N_11530,N_6483,N_7863);
nand U11531 (N_11531,N_8395,N_7683);
xnor U11532 (N_11532,N_5429,N_6216);
nand U11533 (N_11533,N_5137,N_5188);
nand U11534 (N_11534,N_6031,N_6561);
nor U11535 (N_11535,N_7658,N_5856);
or U11536 (N_11536,N_9411,N_9760);
nor U11537 (N_11537,N_9002,N_5907);
or U11538 (N_11538,N_5726,N_7357);
or U11539 (N_11539,N_8660,N_8230);
xor U11540 (N_11540,N_6684,N_6243);
and U11541 (N_11541,N_9793,N_9688);
nand U11542 (N_11542,N_5396,N_8959);
xor U11543 (N_11543,N_5886,N_6633);
or U11544 (N_11544,N_6459,N_6017);
nand U11545 (N_11545,N_6537,N_8262);
nor U11546 (N_11546,N_8049,N_8680);
xnor U11547 (N_11547,N_8168,N_9016);
xor U11548 (N_11548,N_9402,N_8610);
nand U11549 (N_11549,N_7303,N_7122);
or U11550 (N_11550,N_5986,N_5240);
nor U11551 (N_11551,N_9161,N_6195);
and U11552 (N_11552,N_6695,N_7979);
or U11553 (N_11553,N_9463,N_7905);
nand U11554 (N_11554,N_8528,N_9405);
xor U11555 (N_11555,N_5379,N_6495);
xnor U11556 (N_11556,N_7346,N_7409);
nand U11557 (N_11557,N_5645,N_6046);
and U11558 (N_11558,N_5771,N_7200);
nand U11559 (N_11559,N_9281,N_5103);
nor U11560 (N_11560,N_5793,N_8194);
xnor U11561 (N_11561,N_9991,N_6672);
nand U11562 (N_11562,N_5621,N_7198);
nor U11563 (N_11563,N_5024,N_8706);
or U11564 (N_11564,N_7421,N_8710);
xor U11565 (N_11565,N_8483,N_6351);
nor U11566 (N_11566,N_7824,N_6683);
or U11567 (N_11567,N_5781,N_9291);
nor U11568 (N_11568,N_6127,N_5212);
xnor U11569 (N_11569,N_7974,N_6893);
nand U11570 (N_11570,N_5570,N_7614);
or U11571 (N_11571,N_5710,N_6786);
or U11572 (N_11572,N_6380,N_6458);
xnor U11573 (N_11573,N_9938,N_7696);
nand U11574 (N_11574,N_6444,N_8686);
nand U11575 (N_11575,N_7814,N_5959);
or U11576 (N_11576,N_7819,N_6400);
nor U11577 (N_11577,N_5082,N_9845);
or U11578 (N_11578,N_6625,N_9273);
xor U11579 (N_11579,N_9699,N_8780);
or U11580 (N_11580,N_5742,N_6347);
xor U11581 (N_11581,N_9088,N_5190);
or U11582 (N_11582,N_5114,N_5977);
or U11583 (N_11583,N_7446,N_9133);
and U11584 (N_11584,N_6191,N_9791);
xnor U11585 (N_11585,N_7945,N_9763);
nand U11586 (N_11586,N_9926,N_8333);
xor U11587 (N_11587,N_5761,N_6197);
xor U11588 (N_11588,N_6790,N_7533);
and U11589 (N_11589,N_9061,N_9682);
and U11590 (N_11590,N_9514,N_9073);
or U11591 (N_11591,N_5356,N_9258);
nand U11592 (N_11592,N_9521,N_9897);
nand U11593 (N_11593,N_7777,N_9966);
xnor U11594 (N_11594,N_7076,N_8821);
nand U11595 (N_11595,N_8220,N_5950);
or U11596 (N_11596,N_6667,N_6377);
and U11597 (N_11597,N_8001,N_8163);
or U11598 (N_11598,N_6312,N_8685);
or U11599 (N_11599,N_6750,N_6142);
nor U11600 (N_11600,N_7187,N_9752);
or U11601 (N_11601,N_9794,N_8406);
and U11602 (N_11602,N_5608,N_6866);
or U11603 (N_11603,N_8642,N_6653);
and U11604 (N_11604,N_9754,N_9288);
and U11605 (N_11605,N_6792,N_8738);
xnor U11606 (N_11606,N_9414,N_9748);
nor U11607 (N_11607,N_6244,N_8781);
xnor U11608 (N_11608,N_6107,N_5910);
and U11609 (N_11609,N_5022,N_6304);
and U11610 (N_11610,N_8091,N_6105);
or U11611 (N_11611,N_7100,N_5560);
and U11612 (N_11612,N_6734,N_9905);
xor U11613 (N_11613,N_7000,N_5903);
or U11614 (N_11614,N_7944,N_8678);
and U11615 (N_11615,N_6556,N_9556);
nand U11616 (N_11616,N_7170,N_8032);
nand U11617 (N_11617,N_8017,N_8263);
nor U11618 (N_11618,N_7511,N_8320);
or U11619 (N_11619,N_5753,N_6875);
or U11620 (N_11620,N_8640,N_8303);
nor U11621 (N_11621,N_6689,N_6974);
xor U11622 (N_11622,N_9715,N_7213);
nand U11623 (N_11623,N_8272,N_7459);
and U11624 (N_11624,N_6995,N_6302);
nand U11625 (N_11625,N_5945,N_6568);
nor U11626 (N_11626,N_6677,N_7647);
nor U11627 (N_11627,N_8579,N_7432);
and U11628 (N_11628,N_7663,N_6261);
or U11629 (N_11629,N_5835,N_6737);
and U11630 (N_11630,N_5169,N_8167);
xor U11631 (N_11631,N_5473,N_5843);
nand U11632 (N_11632,N_5023,N_7748);
xnor U11633 (N_11633,N_8421,N_7379);
xor U11634 (N_11634,N_8457,N_9262);
nor U11635 (N_11635,N_9780,N_9272);
nor U11636 (N_11636,N_9077,N_9371);
nand U11637 (N_11637,N_5464,N_6593);
or U11638 (N_11638,N_9146,N_9154);
or U11639 (N_11639,N_6513,N_7995);
nand U11640 (N_11640,N_8350,N_9874);
nand U11641 (N_11641,N_7780,N_7493);
xor U11642 (N_11642,N_5489,N_7589);
and U11643 (N_11643,N_8880,N_8343);
and U11644 (N_11644,N_6949,N_5777);
nor U11645 (N_11645,N_9160,N_7131);
nor U11646 (N_11646,N_5498,N_8994);
nand U11647 (N_11647,N_6997,N_5479);
nor U11648 (N_11648,N_9490,N_8775);
and U11649 (N_11649,N_5662,N_7312);
nor U11650 (N_11650,N_7634,N_8882);
and U11651 (N_11651,N_8723,N_9625);
nand U11652 (N_11652,N_7933,N_5720);
xnor U11653 (N_11653,N_8381,N_7822);
or U11654 (N_11654,N_6535,N_5729);
nand U11655 (N_11655,N_8093,N_8197);
nor U11656 (N_11656,N_9332,N_6162);
xnor U11657 (N_11657,N_8968,N_8174);
or U11658 (N_11658,N_9517,N_8345);
nor U11659 (N_11659,N_8823,N_9961);
nor U11660 (N_11660,N_6111,N_6956);
or U11661 (N_11661,N_9558,N_9171);
nor U11662 (N_11662,N_8702,N_8306);
or U11663 (N_11663,N_5528,N_6174);
nand U11664 (N_11664,N_5897,N_5844);
or U11665 (N_11665,N_8283,N_5211);
nand U11666 (N_11666,N_7893,N_5094);
nor U11667 (N_11667,N_8473,N_7399);
nor U11668 (N_11668,N_6215,N_7687);
and U11669 (N_11669,N_9616,N_5173);
nor U11670 (N_11670,N_8012,N_5368);
xor U11671 (N_11671,N_8679,N_8324);
and U11672 (N_11672,N_5380,N_7169);
and U11673 (N_11673,N_8598,N_7216);
nor U11674 (N_11674,N_5644,N_9487);
nand U11675 (N_11675,N_7738,N_8837);
nor U11676 (N_11676,N_6034,N_6102);
or U11677 (N_11677,N_8506,N_6294);
xnor U11678 (N_11678,N_9472,N_7883);
xor U11679 (N_11679,N_7082,N_6542);
nand U11680 (N_11680,N_8989,N_7105);
nor U11681 (N_11681,N_6943,N_6186);
nor U11682 (N_11682,N_9610,N_7990);
nor U11683 (N_11683,N_8869,N_5673);
and U11684 (N_11684,N_8800,N_8102);
or U11685 (N_11685,N_9265,N_9392);
xor U11686 (N_11686,N_6462,N_5122);
and U11687 (N_11687,N_6868,N_8411);
or U11688 (N_11688,N_5160,N_7789);
nor U11689 (N_11689,N_5425,N_7740);
and U11690 (N_11690,N_9062,N_5100);
nor U11691 (N_11691,N_5815,N_6023);
and U11692 (N_11692,N_8669,N_6001);
nor U11693 (N_11693,N_7566,N_9468);
nor U11694 (N_11694,N_9489,N_5839);
nor U11695 (N_11695,N_5741,N_5278);
nor U11696 (N_11696,N_8687,N_5566);
xor U11697 (N_11697,N_8124,N_6853);
xor U11698 (N_11698,N_5262,N_9533);
xnor U11699 (N_11699,N_8417,N_9731);
xor U11700 (N_11700,N_6025,N_6548);
or U11701 (N_11701,N_6867,N_7061);
or U11702 (N_11702,N_7204,N_5655);
xor U11703 (N_11703,N_8204,N_7413);
and U11704 (N_11704,N_6314,N_8029);
nor U11705 (N_11705,N_6026,N_8055);
or U11706 (N_11706,N_9275,N_9649);
nor U11707 (N_11707,N_9960,N_9609);
nor U11708 (N_11708,N_9795,N_8960);
nand U11709 (N_11709,N_8756,N_6664);
nor U11710 (N_11710,N_8529,N_8970);
nand U11711 (N_11711,N_6659,N_6263);
and U11712 (N_11712,N_8517,N_9827);
nor U11713 (N_11713,N_9993,N_6774);
or U11714 (N_11714,N_5239,N_8866);
or U11715 (N_11715,N_9313,N_9693);
nand U11716 (N_11716,N_7641,N_9755);
and U11717 (N_11717,N_7392,N_7610);
nor U11718 (N_11718,N_9531,N_7378);
xor U11719 (N_11719,N_6732,N_9070);
nor U11720 (N_11720,N_5407,N_5327);
xnor U11721 (N_11721,N_6383,N_8101);
nand U11722 (N_11722,N_9126,N_5413);
nand U11723 (N_11723,N_6921,N_7837);
and U11724 (N_11724,N_6370,N_7770);
and U11725 (N_11725,N_9787,N_5690);
nor U11726 (N_11726,N_8726,N_6116);
nor U11727 (N_11727,N_8489,N_5571);
nand U11728 (N_11728,N_7467,N_6076);
or U11729 (N_11729,N_6323,N_6198);
and U11730 (N_11730,N_6460,N_7486);
xor U11731 (N_11731,N_5688,N_6443);
and U11732 (N_11732,N_7028,N_7612);
nor U11733 (N_11733,N_7887,N_9074);
nor U11734 (N_11734,N_5322,N_6386);
nor U11735 (N_11735,N_9358,N_6120);
nand U11736 (N_11736,N_9882,N_6984);
nand U11737 (N_11737,N_7924,N_6106);
or U11738 (N_11738,N_8222,N_6435);
and U11739 (N_11739,N_5846,N_6099);
nor U11740 (N_11740,N_8365,N_6878);
and U11741 (N_11741,N_9555,N_9900);
nand U11742 (N_11742,N_6585,N_8523);
and U11743 (N_11743,N_6901,N_5354);
nand U11744 (N_11744,N_5993,N_7848);
nor U11745 (N_11745,N_9786,N_6229);
nor U11746 (N_11746,N_8138,N_6225);
or U11747 (N_11747,N_7182,N_7724);
nand U11748 (N_11748,N_5668,N_5256);
nand U11749 (N_11749,N_6538,N_6549);
or U11750 (N_11750,N_6279,N_7694);
nor U11751 (N_11751,N_6355,N_5917);
nor U11752 (N_11752,N_5292,N_6473);
nor U11753 (N_11753,N_9522,N_6900);
or U11754 (N_11754,N_6629,N_7732);
or U11755 (N_11755,N_9271,N_7795);
xnor U11756 (N_11756,N_8716,N_9979);
xor U11757 (N_11757,N_5724,N_8108);
or U11758 (N_11758,N_5812,N_9550);
nand U11759 (N_11759,N_5811,N_8264);
nand U11760 (N_11760,N_8977,N_8826);
xor U11761 (N_11761,N_5980,N_7569);
and U11762 (N_11762,N_7774,N_5541);
xor U11763 (N_11763,N_8973,N_6714);
nand U11764 (N_11764,N_8070,N_5398);
xnor U11765 (N_11765,N_5904,N_5756);
xor U11766 (N_11766,N_8942,N_8184);
nand U11767 (N_11767,N_7983,N_7146);
nand U11768 (N_11768,N_8063,N_7948);
xor U11769 (N_11769,N_6598,N_5549);
nor U11770 (N_11770,N_5719,N_7180);
nand U11771 (N_11771,N_7308,N_9377);
nor U11772 (N_11772,N_9441,N_8550);
nor U11773 (N_11773,N_7685,N_9670);
nor U11774 (N_11774,N_5486,N_6700);
or U11775 (N_11775,N_8570,N_9342);
and U11776 (N_11776,N_7802,N_8941);
xor U11777 (N_11777,N_7341,N_6508);
nand U11778 (N_11778,N_6326,N_6056);
or U11779 (N_11779,N_6129,N_9782);
xnor U11780 (N_11780,N_6036,N_8486);
nor U11781 (N_11781,N_5628,N_8596);
nand U11782 (N_11782,N_7238,N_9906);
or U11783 (N_11783,N_9284,N_5475);
nor U11784 (N_11784,N_8697,N_5677);
nand U11785 (N_11785,N_9668,N_6234);
or U11786 (N_11786,N_6586,N_8412);
or U11787 (N_11787,N_9278,N_5308);
xnor U11788 (N_11788,N_7253,N_6519);
and U11789 (N_11789,N_6181,N_5998);
nor U11790 (N_11790,N_7475,N_8802);
nand U11791 (N_11791,N_9111,N_5191);
and U11792 (N_11792,N_6313,N_7970);
nor U11793 (N_11793,N_8703,N_5883);
nor U11794 (N_11794,N_6253,N_7923);
nand U11795 (N_11795,N_9155,N_7916);
xor U11796 (N_11796,N_7864,N_6471);
nor U11797 (N_11797,N_7601,N_9306);
and U11798 (N_11798,N_8891,N_8842);
and U11799 (N_11799,N_5651,N_5523);
nand U11800 (N_11800,N_8772,N_5374);
nand U11801 (N_11801,N_7313,N_5362);
or U11802 (N_11802,N_7929,N_9060);
and U11803 (N_11803,N_5071,N_5445);
xor U11804 (N_11804,N_6770,N_8605);
or U11805 (N_11805,N_9465,N_6751);
or U11806 (N_11806,N_7880,N_5938);
and U11807 (N_11807,N_9696,N_7407);
nor U11808 (N_11808,N_6452,N_7463);
nand U11809 (N_11809,N_7925,N_7153);
and U11810 (N_11810,N_8067,N_7298);
nand U11811 (N_11811,N_7471,N_9864);
or U11812 (N_11812,N_8430,N_6499);
nor U11813 (N_11813,N_7750,N_8966);
or U11814 (N_11814,N_7602,N_6606);
and U11815 (N_11815,N_5575,N_6648);
and U11816 (N_11816,N_9662,N_8299);
nand U11817 (N_11817,N_6125,N_5518);
xnor U11818 (N_11818,N_7699,N_8948);
and U11819 (N_11819,N_8053,N_9067);
nor U11820 (N_11820,N_9992,N_5062);
nor U11821 (N_11821,N_7003,N_6589);
nand U11822 (N_11822,N_6696,N_7410);
nand U11823 (N_11823,N_7648,N_9775);
and U11824 (N_11824,N_7725,N_7506);
xnor U11825 (N_11825,N_5180,N_5504);
xnor U11826 (N_11826,N_5166,N_8814);
nand U11827 (N_11827,N_8459,N_5369);
or U11828 (N_11828,N_9202,N_8785);
and U11829 (N_11829,N_6931,N_8930);
nor U11830 (N_11830,N_7056,N_8484);
and U11831 (N_11831,N_9602,N_6822);
or U11832 (N_11832,N_6924,N_5119);
and U11833 (N_11833,N_6691,N_6385);
xor U11834 (N_11834,N_9508,N_6705);
nor U11835 (N_11835,N_8895,N_9235);
xnor U11836 (N_11836,N_7159,N_6396);
nor U11837 (N_11837,N_9206,N_8060);
xnor U11838 (N_11838,N_8302,N_8020);
nor U11839 (N_11839,N_9603,N_5294);
and U11840 (N_11840,N_7949,N_5152);
and U11841 (N_11841,N_9621,N_9747);
and U11842 (N_11842,N_6067,N_9865);
xnor U11843 (N_11843,N_8076,N_9844);
nor U11844 (N_11844,N_6871,N_7206);
nand U11845 (N_11845,N_8547,N_9825);
nor U11846 (N_11846,N_7886,N_9876);
and U11847 (N_11847,N_9934,N_7800);
xnor U11848 (N_11848,N_7258,N_8367);
or U11849 (N_11849,N_7826,N_9450);
nand U11850 (N_11850,N_9957,N_7709);
nor U11851 (N_11851,N_9596,N_8024);
and U11852 (N_11852,N_5625,N_9935);
and U11853 (N_11853,N_7240,N_5382);
and U11854 (N_11854,N_8379,N_8995);
or U11855 (N_11855,N_6993,N_9385);
or U11856 (N_11856,N_6303,N_6764);
or U11857 (N_11857,N_5775,N_9879);
xnor U11858 (N_11858,N_6194,N_9959);
and U11859 (N_11859,N_6112,N_6596);
nand U11860 (N_11860,N_8073,N_7052);
and U11861 (N_11861,N_9451,N_9491);
nor U11862 (N_11862,N_7055,N_6540);
nor U11863 (N_11863,N_5388,N_6767);
or U11864 (N_11864,N_8972,N_6821);
and U11865 (N_11865,N_9221,N_8123);
nor U11866 (N_11866,N_5658,N_9261);
xor U11867 (N_11867,N_9075,N_9835);
nor U11868 (N_11868,N_7504,N_6165);
xor U11869 (N_11869,N_8467,N_7060);
nor U11870 (N_11870,N_7064,N_6771);
nand U11871 (N_11871,N_5102,N_5674);
and U11872 (N_11872,N_7359,N_5301);
or U11873 (N_11873,N_6688,N_6008);
xor U11874 (N_11874,N_5660,N_5803);
xnor U11875 (N_11875,N_9412,N_6432);
xor U11876 (N_11876,N_8371,N_9595);
and U11877 (N_11877,N_9290,N_6935);
nand U11878 (N_11878,N_9389,N_5192);
nand U11879 (N_11879,N_5187,N_9050);
and U11880 (N_11880,N_5641,N_9357);
nand U11881 (N_11881,N_7194,N_5635);
nor U11882 (N_11882,N_6602,N_7618);
nor U11883 (N_11883,N_6235,N_8490);
nor U11884 (N_11884,N_8929,N_9889);
and U11885 (N_11885,N_9872,N_9687);
nand U11886 (N_11886,N_8399,N_8085);
or U11887 (N_11887,N_7820,N_9811);
and U11888 (N_11888,N_7871,N_9185);
and U11889 (N_11889,N_6301,N_5303);
nor U11890 (N_11890,N_6208,N_8054);
and U11891 (N_11891,N_9856,N_7645);
or U11892 (N_11892,N_9672,N_5483);
xor U11893 (N_11893,N_7662,N_7857);
xnor U11894 (N_11894,N_8786,N_9816);
nand U11895 (N_11895,N_6352,N_8924);
and U11896 (N_11896,N_5214,N_8812);
nor U11897 (N_11897,N_5377,N_5714);
xor U11898 (N_11898,N_7593,N_6029);
and U11899 (N_11899,N_5258,N_6147);
or U11900 (N_11900,N_5687,N_6275);
nor U11901 (N_11901,N_5244,N_7348);
xor U11902 (N_11902,N_6149,N_8857);
nand U11903 (N_11903,N_6945,N_6365);
and U11904 (N_11904,N_9507,N_7897);
nand U11905 (N_11905,N_6024,N_7626);
or U11906 (N_11906,N_8747,N_5096);
or U11907 (N_11907,N_7023,N_9175);
nor U11908 (N_11908,N_8724,N_8390);
xnor U11909 (N_11909,N_8543,N_5466);
nand U11910 (N_11910,N_6886,N_7917);
xor U11911 (N_11911,N_8719,N_6109);
and U11912 (N_11912,N_8981,N_5503);
and U11913 (N_11913,N_6912,N_5934);
or U11914 (N_11914,N_7225,N_7143);
and U11915 (N_11915,N_9335,N_6307);
nor U11916 (N_11916,N_7015,N_6277);
nor U11917 (N_11917,N_8363,N_6908);
and U11918 (N_11918,N_9858,N_8137);
or U11919 (N_11919,N_6755,N_9520);
and U11920 (N_11920,N_8904,N_6098);
xnor U11921 (N_11921,N_5456,N_6185);
nand U11922 (N_11922,N_8974,N_5282);
nor U11923 (N_11923,N_7711,N_9613);
or U11924 (N_11924,N_6551,N_5990);
or U11925 (N_11925,N_5757,N_8717);
nand U11926 (N_11926,N_7241,N_7557);
nand U11927 (N_11927,N_6582,N_8426);
or U11928 (N_11928,N_8743,N_6335);
xor U11929 (N_11929,N_5031,N_7343);
xnor U11930 (N_11930,N_5040,N_5168);
xor U11931 (N_11931,N_7445,N_9394);
or U11932 (N_11932,N_5895,N_8572);
nor U11933 (N_11933,N_8105,N_7629);
and U11934 (N_11934,N_7001,N_5409);
and U11935 (N_11935,N_7314,N_8361);
nand U11936 (N_11936,N_5794,N_7398);
and U11937 (N_11937,N_8613,N_8433);
and U11938 (N_11938,N_9645,N_8038);
nand U11939 (N_11939,N_6461,N_7989);
nand U11940 (N_11940,N_6791,N_7107);
and U11941 (N_11941,N_9384,N_6557);
nand U11942 (N_11942,N_9869,N_7650);
nor U11943 (N_11943,N_7958,N_6872);
and U11944 (N_11944,N_8804,N_7710);
xor U11945 (N_11945,N_8318,N_6090);
xnor U11946 (N_11946,N_7546,N_6002);
and U11947 (N_11947,N_6936,N_6839);
or U11948 (N_11948,N_9840,N_5885);
nand U11949 (N_11949,N_8455,N_6199);
nor U11950 (N_11950,N_6846,N_9098);
nor U11951 (N_11951,N_9415,N_6060);
nor U11952 (N_11952,N_5058,N_6517);
xor U11953 (N_11953,N_7733,N_6357);
and U11954 (N_11954,N_9216,N_6353);
xor U11955 (N_11955,N_5623,N_8871);
and U11956 (N_11956,N_8357,N_7497);
and U11957 (N_11957,N_6970,N_5434);
and U11958 (N_11958,N_8505,N_7077);
and U11959 (N_11959,N_8913,N_5694);
or U11960 (N_11960,N_5235,N_6926);
nand U11961 (N_11961,N_5954,N_9268);
or U11962 (N_11962,N_6028,N_5791);
or U11963 (N_11963,N_7836,N_9147);
or U11964 (N_11964,N_7548,N_7784);
and U11965 (N_11965,N_6438,N_9544);
nor U11966 (N_11966,N_5133,N_7942);
xnor U11967 (N_11967,N_5485,N_5261);
and U11968 (N_11968,N_8125,N_7535);
nor U11969 (N_11969,N_7305,N_5049);
or U11970 (N_11970,N_7943,N_8021);
or U11971 (N_11971,N_9939,N_7040);
nor U11972 (N_11972,N_6164,N_5985);
or U11973 (N_11973,N_9587,N_5707);
nand U11974 (N_11974,N_7889,N_6773);
nand U11975 (N_11975,N_5217,N_9017);
nand U11976 (N_11976,N_8008,N_9600);
and U11977 (N_11977,N_6590,N_5331);
nand U11978 (N_11978,N_9382,N_9010);
nand U11979 (N_11979,N_8705,N_6989);
xnor U11980 (N_11980,N_8241,N_7117);
and U11981 (N_11981,N_8752,N_8511);
or U11982 (N_11982,N_8000,N_8856);
nand U11983 (N_11983,N_9788,N_6006);
or U11984 (N_11984,N_6287,N_8376);
and U11985 (N_11985,N_7806,N_8725);
nor U11986 (N_11986,N_9326,N_5174);
and U11987 (N_11987,N_6965,N_5763);
and U11988 (N_11988,N_7976,N_8072);
xor U11989 (N_11989,N_9607,N_7344);
and U11990 (N_11990,N_7285,N_7903);
or U11991 (N_11991,N_7041,N_9207);
or U11992 (N_11992,N_6806,N_5653);
nor U11993 (N_11993,N_5789,N_7431);
nand U11994 (N_11994,N_5650,N_9112);
or U11995 (N_11995,N_5460,N_8133);
nand U11996 (N_11996,N_8583,N_6665);
nand U11997 (N_11997,N_7113,N_8817);
or U11998 (N_11998,N_8122,N_5440);
xor U11999 (N_11999,N_8420,N_8997);
and U12000 (N_12000,N_8558,N_6178);
nor U12001 (N_12001,N_7649,N_5289);
and U12002 (N_12002,N_7675,N_5449);
or U12003 (N_12003,N_9511,N_7145);
xnor U12004 (N_12004,N_7168,N_9843);
or U12005 (N_12005,N_7761,N_5098);
xor U12006 (N_12006,N_7072,N_6219);
nor U12007 (N_12007,N_7521,N_7692);
or U12008 (N_12008,N_8016,N_6986);
nand U12009 (N_12009,N_7296,N_8603);
and U12010 (N_12010,N_6626,N_7393);
or U12011 (N_12011,N_9003,N_7834);
or U12012 (N_12012,N_6498,N_8524);
nor U12013 (N_12013,N_6968,N_9381);
nor U12014 (N_12014,N_8797,N_8841);
and U12015 (N_12015,N_5680,N_6547);
nor U12016 (N_12016,N_7172,N_5656);
or U12017 (N_12017,N_7412,N_7081);
nand U12018 (N_12018,N_9654,N_6320);
nand U12019 (N_12019,N_6941,N_5299);
nor U12020 (N_12020,N_9822,N_7509);
or U12021 (N_12021,N_8161,N_6423);
xor U12022 (N_12022,N_8463,N_7500);
or U12023 (N_12023,N_8437,N_6466);
or U12024 (N_12024,N_9014,N_8843);
or U12025 (N_12025,N_6052,N_7460);
and U12026 (N_12026,N_6881,N_8711);
or U12027 (N_12027,N_8316,N_5516);
or U12028 (N_12028,N_9740,N_8901);
nor U12029 (N_12029,N_9099,N_8494);
xor U12030 (N_12030,N_6911,N_8986);
nand U12031 (N_12031,N_9629,N_8011);
xor U12032 (N_12032,N_5312,N_7633);
xnor U12033 (N_12033,N_5234,N_7677);
or U12034 (N_12034,N_8027,N_6555);
nand U12035 (N_12035,N_7452,N_7638);
nand U12036 (N_12036,N_9941,N_8329);
or U12037 (N_12037,N_8407,N_8589);
nor U12038 (N_12038,N_9802,N_5251);
or U12039 (N_12039,N_7868,N_9448);
and U12040 (N_12040,N_5599,N_5003);
nor U12041 (N_12041,N_6885,N_7513);
or U12042 (N_12042,N_5052,N_8209);
and U12043 (N_12043,N_6584,N_7443);
xnor U12044 (N_12044,N_9169,N_8444);
xnor U12045 (N_12045,N_5025,N_6726);
nor U12046 (N_12046,N_7581,N_9201);
or U12047 (N_12047,N_8996,N_5167);
and U12048 (N_12048,N_5257,N_7698);
xor U12049 (N_12049,N_8946,N_5551);
nand U12050 (N_12050,N_6074,N_6877);
nand U12051 (N_12051,N_5996,N_7163);
xor U12052 (N_12052,N_5076,N_9479);
and U12053 (N_12053,N_8192,N_5158);
and U12054 (N_12054,N_7327,N_6869);
or U12055 (N_12055,N_7584,N_9768);
nand U12056 (N_12056,N_9055,N_7544);
and U12057 (N_12057,N_9746,N_6917);
xnor U12058 (N_12058,N_5693,N_6880);
or U12059 (N_12059,N_5708,N_9642);
nand U12060 (N_12060,N_7489,N_9797);
xnor U12061 (N_12061,N_5057,N_5451);
xnor U12062 (N_12062,N_8019,N_5929);
and U12063 (N_12063,N_5887,N_7480);
nand U12064 (N_12064,N_9233,N_9004);
or U12065 (N_12065,N_7906,N_9552);
nor U12066 (N_12066,N_6948,N_6481);
or U12067 (N_12067,N_9547,N_7025);
xnor U12068 (N_12068,N_9040,N_9737);
and U12069 (N_12069,N_8416,N_9708);
or U12070 (N_12070,N_5467,N_9365);
xor U12071 (N_12071,N_5762,N_9834);
or U12072 (N_12072,N_9639,N_6085);
and U12073 (N_12073,N_8639,N_9619);
nor U12074 (N_12074,N_9400,N_7144);
nand U12075 (N_12075,N_6137,N_6321);
xor U12076 (N_12076,N_8425,N_8620);
nand U12077 (N_12077,N_7578,N_5624);
nand U12078 (N_12078,N_8396,N_5669);
nand U12079 (N_12079,N_9851,N_8795);
nand U12080 (N_12080,N_8142,N_8829);
nor U12081 (N_12081,N_7267,N_5131);
and U12082 (N_12082,N_6919,N_6154);
or U12083 (N_12083,N_8150,N_9651);
xor U12084 (N_12084,N_5066,N_5877);
xor U12085 (N_12085,N_6647,N_6505);
xnor U12086 (N_12086,N_5325,N_5424);
nand U12087 (N_12087,N_8188,N_9691);
nor U12088 (N_12088,N_8791,N_7644);
nand U12089 (N_12089,N_6578,N_5587);
and U12090 (N_12090,N_6160,N_7468);
nand U12091 (N_12091,N_9251,N_6228);
nor U12092 (N_12092,N_6493,N_9990);
or U12093 (N_12093,N_8849,N_8248);
nor U12094 (N_12094,N_7239,N_8018);
or U12095 (N_12095,N_9188,N_8195);
or U12096 (N_12096,N_5346,N_6280);
nor U12097 (N_12097,N_6032,N_5751);
or U12098 (N_12098,N_8040,N_7811);
or U12099 (N_12099,N_8709,N_8267);
nor U12100 (N_12100,N_8276,N_7292);
and U12101 (N_12101,N_9601,N_8552);
nand U12102 (N_12102,N_6699,N_7036);
nor U12103 (N_12103,N_7503,N_8532);
and U12104 (N_12104,N_5358,N_9784);
or U12105 (N_12105,N_9427,N_8228);
nor U12106 (N_12106,N_6039,N_8313);
or U12107 (N_12107,N_9127,N_9730);
nor U12108 (N_12108,N_8179,N_8218);
nor U12109 (N_12109,N_7039,N_7362);
nand U12110 (N_12110,N_8649,N_9186);
xor U12111 (N_12111,N_7207,N_6507);
nand U12112 (N_12112,N_8502,N_9316);
or U12113 (N_12113,N_8349,N_5359);
xor U12114 (N_12114,N_8249,N_9094);
nor U12115 (N_12115,N_5778,N_6075);
xor U12116 (N_12116,N_7309,N_9713);
or U12117 (N_12117,N_7426,N_9082);
nor U12118 (N_12118,N_7554,N_8144);
and U12119 (N_12119,N_7106,N_8577);
or U12120 (N_12120,N_8750,N_5394);
or U12121 (N_12121,N_6739,N_5868);
nor U12122 (N_12122,N_8975,N_5557);
and U12123 (N_12123,N_7727,N_5065);
or U12124 (N_12124,N_5610,N_5788);
nor U12125 (N_12125,N_7345,N_6873);
nor U12126 (N_12126,N_6425,N_5128);
xnor U12127 (N_12127,N_7797,N_6899);
xnor U12128 (N_12128,N_6439,N_6998);
or U12129 (N_12129,N_7558,N_5297);
xor U12130 (N_12130,N_7137,N_8368);
nor U12131 (N_12131,N_6565,N_6932);
or U12132 (N_12132,N_8683,N_7226);
nand U12133 (N_12133,N_7862,N_9303);
or U12134 (N_12134,N_5228,N_6828);
and U12135 (N_12135,N_5828,N_8022);
or U12136 (N_12136,N_6410,N_5939);
nor U12137 (N_12137,N_9021,N_6674);
nand U12138 (N_12138,N_9659,N_5129);
and U12139 (N_12139,N_7235,N_7209);
and U12140 (N_12140,N_9170,N_6246);
xor U12141 (N_12141,N_6666,N_7089);
nor U12142 (N_12142,N_9293,N_8662);
or U12143 (N_12143,N_8887,N_6247);
and U12144 (N_12144,N_6717,N_9093);
xnor U12145 (N_12145,N_9716,N_5739);
or U12146 (N_12146,N_5831,N_8129);
xor U12147 (N_12147,N_8734,N_7597);
nor U12148 (N_12148,N_9204,N_7841);
xnor U12149 (N_12149,N_9056,N_6940);
nor U12150 (N_12150,N_7873,N_8048);
nor U12151 (N_12151,N_9315,N_6003);
nor U12152 (N_12152,N_9237,N_8926);
nor U12153 (N_12153,N_7838,N_7937);
nor U12154 (N_12154,N_7266,N_7488);
xor U12155 (N_12155,N_8440,N_5223);
or U12156 (N_12156,N_6641,N_5947);
and U12157 (N_12157,N_9406,N_7441);
and U12158 (N_12158,N_6494,N_5204);
or U12159 (N_12159,N_8282,N_8213);
xnor U12160 (N_12160,N_5826,N_8005);
and U12161 (N_12161,N_8140,N_6736);
and U12162 (N_12162,N_6418,N_5728);
nand U12163 (N_12163,N_5629,N_8715);
or U12164 (N_12164,N_7825,N_6553);
nand U12165 (N_12165,N_7796,N_8820);
xor U12166 (N_12166,N_7176,N_6600);
or U12167 (N_12167,N_7355,N_9553);
nor U12168 (N_12168,N_8385,N_9914);
xor U12169 (N_12169,N_9135,N_7374);
and U12170 (N_12170,N_5097,N_5545);
nand U12171 (N_12171,N_6044,N_7135);
xnor U12172 (N_12172,N_8492,N_9344);
nand U12173 (N_12173,N_7051,N_7333);
xnor U12174 (N_12174,N_5070,N_9407);
nor U12175 (N_12175,N_8378,N_9714);
and U12176 (N_12176,N_6716,N_5898);
and U12177 (N_12177,N_5808,N_9102);
nand U12178 (N_12178,N_7202,N_6614);
and U12179 (N_12179,N_8405,N_7280);
nand U12180 (N_12180,N_7828,N_8265);
nand U12181 (N_12181,N_8186,N_6829);
or U12182 (N_12182,N_5279,N_9943);
xnor U12183 (N_12183,N_7656,N_6054);
and U12184 (N_12184,N_9440,N_8643);
and U12185 (N_12185,N_8645,N_5514);
nor U12186 (N_12186,N_8295,N_9433);
or U12187 (N_12187,N_5284,N_5484);
xor U12188 (N_12188,N_7098,N_5952);
nand U12189 (N_12189,N_9330,N_8033);
xor U12190 (N_12190,N_6844,N_7046);
nand U12191 (N_12191,N_7845,N_6332);
nand U12192 (N_12192,N_5246,N_6697);
or U12193 (N_12193,N_6038,N_8608);
and U12194 (N_12194,N_7141,N_5825);
and U12195 (N_12195,N_7686,N_5875);
or U12196 (N_12196,N_8559,N_7560);
nor U12197 (N_12197,N_5926,N_8311);
xnor U12198 (N_12198,N_5147,N_5252);
nor U12199 (N_12199,N_9378,N_9409);
nand U12200 (N_12200,N_6605,N_6619);
and U12201 (N_12201,N_8840,N_6378);
or U12202 (N_12202,N_9030,N_9009);
xnor U12203 (N_12203,N_5766,N_7993);
nand U12204 (N_12204,N_5332,N_5344);
and U12205 (N_12205,N_9833,N_6179);
nor U12206 (N_12206,N_9469,N_9694);
xor U12207 (N_12207,N_9481,N_6005);
xnor U12208 (N_12208,N_9673,N_8336);
xnor U12209 (N_12209,N_9300,N_6375);
xnor U12210 (N_12210,N_7759,N_5199);
nand U12211 (N_12211,N_5397,N_9105);
xnor U12212 (N_12212,N_9197,N_7922);
nor U12213 (N_12213,N_5691,N_7059);
nor U12214 (N_12214,N_9375,N_9421);
and U12215 (N_12215,N_5210,N_7596);
or U12216 (N_12216,N_6445,N_7715);
nor U12217 (N_12217,N_7037,N_5307);
xor U12218 (N_12218,N_7652,N_8245);
and U12219 (N_12219,N_9397,N_5389);
or U12220 (N_12220,N_9923,N_7935);
and U12221 (N_12221,N_8398,N_5000);
or U12222 (N_12222,N_9532,N_8969);
nor U12223 (N_12223,N_8925,N_6579);
xnor U12224 (N_12224,N_5026,N_9436);
or U12225 (N_12225,N_8927,N_9824);
nor U12226 (N_12226,N_5045,N_9640);
xnor U12227 (N_12227,N_6364,N_6951);
and U12228 (N_12228,N_5290,N_7328);
and U12229 (N_12229,N_7053,N_9120);
and U12230 (N_12230,N_6212,N_7179);
nand U12231 (N_12231,N_9743,N_8253);
xor U12232 (N_12232,N_8104,N_6372);
nor U12233 (N_12233,N_7798,N_6200);
and U12234 (N_12234,N_6136,N_8971);
or U12235 (N_12235,N_5735,N_9453);
xnor U12236 (N_12236,N_9496,N_5482);
or U12237 (N_12237,N_6082,N_9282);
nor U12238 (N_12238,N_6148,N_9299);
xor U12239 (N_12239,N_6019,N_6497);
nand U12240 (N_12240,N_9217,N_6490);
or U12241 (N_12241,N_8261,N_9505);
and U12242 (N_12242,N_6016,N_8359);
nand U12243 (N_12243,N_9656,N_6692);
xnor U12244 (N_12244,N_6632,N_6574);
nor U12245 (N_12245,N_8246,N_8308);
or U12246 (N_12246,N_7121,N_9568);
and U12247 (N_12247,N_9660,N_8092);
or U12248 (N_12248,N_8203,N_6622);
xnor U12249 (N_12249,N_8604,N_6451);
nand U12250 (N_12250,N_6131,N_8047);
or U12251 (N_12251,N_6091,N_5876);
nor U12252 (N_12252,N_8653,N_9657);
nand U12253 (N_12253,N_8851,N_7951);
or U12254 (N_12254,N_6644,N_6065);
or U12255 (N_12255,N_8557,N_5759);
and U12256 (N_12256,N_9266,N_6671);
nor U12257 (N_12257,N_9580,N_5481);
nor U12258 (N_12258,N_5336,N_5276);
or U12259 (N_12259,N_8205,N_6057);
nor U12260 (N_12260,N_7913,N_9174);
nor U12261 (N_12261,N_8402,N_6161);
or U12262 (N_12262,N_5069,N_8631);
and U12263 (N_12263,N_7681,N_7680);
and U12264 (N_12264,N_7657,N_8898);
or U12265 (N_12265,N_7884,N_6211);
nand U12266 (N_12266,N_8191,N_9915);
and U12267 (N_12267,N_5105,N_5654);
nor U12268 (N_12268,N_6658,N_9173);
nand U12269 (N_12269,N_7218,N_9646);
and U12270 (N_12270,N_8238,N_7330);
nor U12271 (N_12271,N_6298,N_9058);
xor U12272 (N_12272,N_8782,N_6887);
nand U12273 (N_12273,N_9653,N_8293);
and U12274 (N_12274,N_9857,N_8657);
nor U12275 (N_12275,N_9969,N_5222);
xor U12276 (N_12276,N_8727,N_5080);
and U12277 (N_12277,N_7250,N_8515);
or U12278 (N_12278,N_5531,N_5701);
or U12279 (N_12279,N_9821,N_9165);
or U12280 (N_12280,N_5254,N_7265);
xnor U12281 (N_12281,N_9829,N_9975);
or U12282 (N_12282,N_9467,N_9636);
xor U12283 (N_12283,N_8950,N_7860);
xor U12284 (N_12284,N_7262,N_7157);
nor U12285 (N_12285,N_8366,N_9612);
nand U12286 (N_12286,N_5496,N_8796);
and U12287 (N_12287,N_7030,N_6248);
and U12288 (N_12288,N_7329,N_9104);
and U12289 (N_12289,N_7256,N_8518);
nor U12290 (N_12290,N_7782,N_8116);
nand U12291 (N_12291,N_6855,N_8553);
or U12292 (N_12292,N_7255,N_6171);
nor U12293 (N_12293,N_9012,N_9634);
xor U12294 (N_12294,N_8629,N_9967);
or U12295 (N_12295,N_5513,N_6979);
nand U12296 (N_12296,N_9813,N_8601);
nor U12297 (N_12297,N_5372,N_5507);
nand U12298 (N_12298,N_9419,N_5116);
nor U12299 (N_12299,N_7676,N_7165);
or U12300 (N_12300,N_6286,N_8824);
or U12301 (N_12301,N_7668,N_6760);
and U12302 (N_12302,N_9510,N_5936);
or U12303 (N_12303,N_5068,N_7050);
xor U12304 (N_12304,N_8908,N_7620);
xnor U12305 (N_12305,N_5499,N_7695);
or U12306 (N_12306,N_6612,N_8844);
and U12307 (N_12307,N_8740,N_7496);
or U12308 (N_12308,N_6293,N_6436);
nand U12309 (N_12309,N_9644,N_5172);
xnor U12310 (N_12310,N_7173,N_9819);
nand U12311 (N_12311,N_6906,N_8878);
nand U12312 (N_12312,N_6114,N_7196);
and U12313 (N_12313,N_7617,N_6271);
nand U12314 (N_12314,N_8403,N_7684);
and U12315 (N_12315,N_6387,N_5802);
nor U12316 (N_12316,N_9545,N_7151);
or U12317 (N_12317,N_5569,N_7454);
nand U12318 (N_12318,N_8291,N_9878);
nor U12319 (N_12319,N_8004,N_9648);
nand U12320 (N_12320,N_7980,N_5704);
nand U12321 (N_12321,N_5360,N_6329);
or U12322 (N_12322,N_9091,N_6929);
nor U12323 (N_12323,N_6381,N_6707);
nor U12324 (N_12324,N_9771,N_8342);
nand U12325 (N_12325,N_7236,N_8301);
xnor U12326 (N_12326,N_8918,N_7388);
nand U12327 (N_12327,N_7785,N_9850);
xnor U12328 (N_12328,N_8187,N_9661);
xnor U12329 (N_12329,N_9242,N_5820);
nand U12330 (N_12330,N_6639,N_6450);
nor U12331 (N_12331,N_8255,N_7600);
xnor U12332 (N_12332,N_6808,N_6511);
or U12333 (N_12333,N_5032,N_7757);
and U12334 (N_12334,N_8594,N_5335);
or U12335 (N_12335,N_9847,N_6824);
or U12336 (N_12336,N_9887,N_6168);
and U12337 (N_12337,N_6843,N_8279);
nand U12338 (N_12338,N_8670,N_8254);
xnor U12339 (N_12339,N_9426,N_6061);
or U12340 (N_12340,N_9783,N_8297);
nor U12341 (N_12341,N_8328,N_6679);
nor U12342 (N_12342,N_9583,N_6408);
xor U12343 (N_12343,N_9989,N_6010);
nor U12344 (N_12344,N_7947,N_8429);
nor U12345 (N_12345,N_7371,N_7440);
or U12346 (N_12346,N_9658,N_7953);
nand U12347 (N_12347,N_7611,N_9995);
or U12348 (N_12348,N_5515,N_7778);
nand U12349 (N_12349,N_5796,N_7248);
xnor U12350 (N_12350,N_8304,N_8207);
nor U12351 (N_12351,N_6920,N_6971);
and U12352 (N_12352,N_5774,N_5259);
nor U12353 (N_12353,N_6643,N_5155);
and U12354 (N_12354,N_9413,N_6757);
or U12355 (N_12355,N_8046,N_8120);
nor U12356 (N_12356,N_9584,N_8894);
nor U12357 (N_12357,N_6662,N_9633);
or U12358 (N_12358,N_6288,N_7027);
nand U12359 (N_12359,N_5689,N_9948);
xor U12360 (N_12360,N_7639,N_7448);
nand U12361 (N_12361,N_6476,N_6270);
nand U12362 (N_12362,N_8154,N_8816);
and U12363 (N_12363,N_8062,N_7984);
nand U12364 (N_12364,N_9684,N_5046);
nand U12365 (N_12365,N_9953,N_6342);
xnor U12366 (N_12366,N_7892,N_9219);
or U12367 (N_12367,N_5579,N_5300);
or U12368 (N_12368,N_6604,N_7045);
xor U12369 (N_12369,N_8362,N_9956);
nand U12370 (N_12370,N_9280,N_8434);
or U12371 (N_12371,N_7047,N_7531);
nor U12372 (N_12372,N_8121,N_8496);
nor U12373 (N_12373,N_5352,N_9627);
nand U12374 (N_12374,N_9921,N_8453);
nand U12375 (N_12375,N_7457,N_8110);
nand U12376 (N_12376,N_8940,N_8514);
or U12377 (N_12377,N_6441,N_5438);
or U12378 (N_12378,N_5444,N_5573);
nand U12379 (N_12379,N_6015,N_9257);
or U12380 (N_12380,N_5964,N_8094);
and U12381 (N_12381,N_5213,N_9841);
xor U12382 (N_12382,N_6723,N_7507);
nand U12383 (N_12383,N_5534,N_7447);
and U12384 (N_12384,N_7227,N_8713);
xor U12385 (N_12385,N_5099,N_5752);
xnor U12386 (N_12386,N_6794,N_7133);
nor U12387 (N_12387,N_5490,N_7807);
and U12388 (N_12388,N_8540,N_8244);
nor U12389 (N_12389,N_7029,N_5615);
xor U12390 (N_12390,N_7070,N_5317);
xor U12391 (N_12391,N_7228,N_5378);
or U12392 (N_12392,N_8485,N_7322);
or U12393 (N_12393,N_8650,N_5836);
nor U12394 (N_12394,N_8298,N_7598);
or U12395 (N_12395,N_6651,N_5181);
nor U12396 (N_12396,N_7582,N_7451);
nand U12397 (N_12397,N_6903,N_7930);
xnor U12398 (N_12398,N_8470,N_7260);
or U12399 (N_12399,N_8667,N_7936);
xor U12400 (N_12400,N_8535,N_8170);
nand U12401 (N_12401,N_9738,N_6749);
nand U12402 (N_12402,N_7536,N_6759);
nand U12403 (N_12403,N_5021,N_8630);
or U12404 (N_12404,N_9836,N_5564);
nor U12405 (N_12405,N_6047,N_7223);
and U12406 (N_12406,N_7874,N_5242);
nand U12407 (N_12407,N_5232,N_6913);
and U12408 (N_12408,N_9031,N_8386);
or U12409 (N_12409,N_9937,N_9084);
xnor U12410 (N_12410,N_5209,N_9789);
or U12411 (N_12411,N_6421,N_5935);
and U12412 (N_12412,N_7619,N_9158);
nor U12413 (N_12413,N_9011,N_8889);
nor U12414 (N_12414,N_6078,N_6522);
or U12415 (N_12415,N_7140,N_7672);
nand U12416 (N_12416,N_9184,N_9674);
xor U12417 (N_12417,N_6501,N_8937);
and U12418 (N_12418,N_6409,N_5737);
nand U12419 (N_12419,N_8744,N_6575);
nor U12420 (N_12420,N_7523,N_8512);
nor U12421 (N_12421,N_9176,N_6613);
xor U12422 (N_12422,N_6904,N_5454);
nand U12423 (N_12423,N_6980,N_5402);
nor U12424 (N_12424,N_7931,N_7981);
nor U12425 (N_12425,N_7326,N_5738);
xor U12426 (N_12426,N_5416,N_5732);
xnor U12427 (N_12427,N_8435,N_8764);
or U12428 (N_12428,N_6187,N_9919);
xor U12429 (N_12429,N_5632,N_7665);
xor U12430 (N_12430,N_5863,N_7918);
and U12431 (N_12431,N_5433,N_7115);
nor U12432 (N_12432,N_6747,N_7717);
xnor U12433 (N_12433,N_5696,N_9528);
or U12434 (N_12434,N_8947,N_9020);
and U12435 (N_12435,N_9543,N_7812);
xor U12436 (N_12436,N_6413,N_5664);
and U12437 (N_12437,N_6305,N_5218);
nor U12438 (N_12438,N_7058,N_6962);
and U12439 (N_12439,N_5419,N_8479);
xor U12440 (N_12440,N_7006,N_9033);
or U12441 (N_12441,N_7044,N_6042);
nor U12442 (N_12442,N_5150,N_7442);
xnor U12443 (N_12443,N_5901,N_6580);
xnor U12444 (N_12444,N_6543,N_6729);
nor U12445 (N_12445,N_9192,N_9626);
xor U12446 (N_12446,N_9080,N_7594);
or U12447 (N_12447,N_6973,N_9777);
nor U12448 (N_12448,N_7707,N_7975);
and U12449 (N_12449,N_6000,N_7801);
xnor U12450 (N_12450,N_5616,N_7992);
nor U12451 (N_12451,N_8146,N_6952);
and U12452 (N_12452,N_9618,N_7682);
nor U12453 (N_12453,N_8976,N_5953);
nand U12454 (N_12454,N_8296,N_9391);
nand U12455 (N_12455,N_6927,N_9025);
nor U12456 (N_12456,N_6349,N_8825);
xor U12457 (N_12457,N_5842,N_8718);
nand U12458 (N_12458,N_5366,N_6937);
nor U12459 (N_12459,N_5862,N_7427);
and U12460 (N_12460,N_7069,N_5054);
and U12461 (N_12461,N_6583,N_6429);
xor U12462 (N_12462,N_8614,N_7960);
or U12463 (N_12463,N_5134,N_9557);
and U12464 (N_12464,N_7400,N_7630);
nand U12465 (N_12465,N_5912,N_9172);
nand U12466 (N_12466,N_5880,N_6062);
nand U12467 (N_12467,N_5814,N_7726);
nor U12468 (N_12468,N_7420,N_8443);
nand U12469 (N_12469,N_5530,N_6175);
or U12470 (N_12470,N_8083,N_5267);
and U12471 (N_12471,N_5553,N_7985);
or U12472 (N_12472,N_8112,N_7817);
and U12473 (N_12473,N_5135,N_6083);
or U12474 (N_12474,N_9733,N_8003);
or U12475 (N_12475,N_7635,N_5149);
or U12476 (N_12476,N_9065,N_7192);
nor U12477 (N_12477,N_8321,N_7853);
xor U12478 (N_12478,N_7580,N_7331);
xnor U12479 (N_12479,N_7914,N_5104);
or U12480 (N_12480,N_6765,N_9895);
xor U12481 (N_12481,N_8269,N_8270);
xnor U12482 (N_12482,N_8833,N_7402);
or U12483 (N_12483,N_7286,N_9226);
nor U12484 (N_12484,N_6446,N_6167);
nor U12485 (N_12485,N_9180,N_7417);
nand U12486 (N_12486,N_5596,N_8219);
and U12487 (N_12487,N_6735,N_8982);
and U12488 (N_12488,N_6701,N_9803);
and U12489 (N_12489,N_8510,N_8961);
xnor U12490 (N_12490,N_7191,N_6072);
nor U12491 (N_12491,N_5957,N_9164);
nand U12492 (N_12492,N_5253,N_9492);
nor U12493 (N_12493,N_8671,N_7428);
xnor U12494 (N_12494,N_8944,N_9709);
xnor U12495 (N_12495,N_5136,N_9917);
and U12496 (N_12496,N_8454,N_8661);
and U12497 (N_12497,N_6454,N_9946);
and U12498 (N_12498,N_9323,N_5801);
or U12499 (N_12499,N_9156,N_6088);
nand U12500 (N_12500,N_7669,N_8347);
nand U12501 (N_12501,N_9900,N_9641);
nor U12502 (N_12502,N_8481,N_5199);
nor U12503 (N_12503,N_7731,N_7792);
nand U12504 (N_12504,N_7925,N_9632);
nand U12505 (N_12505,N_8352,N_6656);
and U12506 (N_12506,N_6124,N_8018);
nand U12507 (N_12507,N_9986,N_7579);
xnor U12508 (N_12508,N_5050,N_6656);
and U12509 (N_12509,N_9430,N_8154);
and U12510 (N_12510,N_6085,N_6131);
nor U12511 (N_12511,N_8387,N_5595);
nand U12512 (N_12512,N_8726,N_9992);
xor U12513 (N_12513,N_6542,N_7845);
nor U12514 (N_12514,N_6219,N_5148);
or U12515 (N_12515,N_8290,N_8023);
xnor U12516 (N_12516,N_8667,N_6394);
and U12517 (N_12517,N_8499,N_9955);
and U12518 (N_12518,N_8033,N_7935);
and U12519 (N_12519,N_8192,N_7947);
xnor U12520 (N_12520,N_9930,N_9712);
nand U12521 (N_12521,N_5342,N_8936);
nor U12522 (N_12522,N_9675,N_5254);
and U12523 (N_12523,N_8423,N_6249);
nor U12524 (N_12524,N_8503,N_9034);
or U12525 (N_12525,N_5674,N_5973);
and U12526 (N_12526,N_6208,N_9066);
nor U12527 (N_12527,N_8645,N_6872);
nand U12528 (N_12528,N_5801,N_5206);
nand U12529 (N_12529,N_5919,N_8324);
and U12530 (N_12530,N_7275,N_8129);
or U12531 (N_12531,N_8855,N_6832);
xnor U12532 (N_12532,N_5480,N_9876);
nand U12533 (N_12533,N_5937,N_9081);
nand U12534 (N_12534,N_7667,N_9839);
nand U12535 (N_12535,N_5867,N_6648);
xnor U12536 (N_12536,N_8181,N_8763);
and U12537 (N_12537,N_5172,N_6703);
xnor U12538 (N_12538,N_6030,N_7720);
nor U12539 (N_12539,N_8737,N_5575);
xor U12540 (N_12540,N_9663,N_5498);
and U12541 (N_12541,N_8409,N_9750);
and U12542 (N_12542,N_5428,N_5214);
nor U12543 (N_12543,N_7834,N_7911);
or U12544 (N_12544,N_8508,N_5545);
xnor U12545 (N_12545,N_8893,N_8276);
and U12546 (N_12546,N_5869,N_8776);
nor U12547 (N_12547,N_9525,N_7411);
and U12548 (N_12548,N_7517,N_5977);
nand U12549 (N_12549,N_5954,N_7297);
nand U12550 (N_12550,N_7926,N_8205);
xnor U12551 (N_12551,N_9506,N_7132);
nor U12552 (N_12552,N_9590,N_7273);
nor U12553 (N_12553,N_8073,N_9269);
nor U12554 (N_12554,N_6270,N_6291);
and U12555 (N_12555,N_7380,N_7653);
and U12556 (N_12556,N_5772,N_7139);
xor U12557 (N_12557,N_9947,N_6157);
nand U12558 (N_12558,N_6860,N_5215);
or U12559 (N_12559,N_5558,N_9917);
xor U12560 (N_12560,N_7303,N_5591);
or U12561 (N_12561,N_9991,N_8397);
xor U12562 (N_12562,N_6802,N_7813);
xor U12563 (N_12563,N_6315,N_5051);
and U12564 (N_12564,N_9441,N_5069);
nand U12565 (N_12565,N_7737,N_6314);
nor U12566 (N_12566,N_8897,N_8616);
and U12567 (N_12567,N_9487,N_8013);
and U12568 (N_12568,N_6345,N_6279);
or U12569 (N_12569,N_5180,N_9609);
and U12570 (N_12570,N_7660,N_9491);
nand U12571 (N_12571,N_8048,N_7484);
or U12572 (N_12572,N_7127,N_6653);
or U12573 (N_12573,N_5193,N_9242);
and U12574 (N_12574,N_7842,N_9657);
xor U12575 (N_12575,N_5988,N_6675);
nand U12576 (N_12576,N_6923,N_8079);
nand U12577 (N_12577,N_6799,N_7000);
and U12578 (N_12578,N_7514,N_7540);
nor U12579 (N_12579,N_9606,N_7449);
and U12580 (N_12580,N_6706,N_9968);
nand U12581 (N_12581,N_7347,N_5431);
nand U12582 (N_12582,N_8603,N_5490);
nand U12583 (N_12583,N_8258,N_7826);
nor U12584 (N_12584,N_8315,N_8016);
nor U12585 (N_12585,N_9307,N_6098);
nor U12586 (N_12586,N_5131,N_8569);
nand U12587 (N_12587,N_8814,N_5566);
or U12588 (N_12588,N_7788,N_5371);
nor U12589 (N_12589,N_6311,N_9256);
and U12590 (N_12590,N_6696,N_9654);
and U12591 (N_12591,N_8935,N_6554);
nor U12592 (N_12592,N_5308,N_5038);
xor U12593 (N_12593,N_5588,N_7765);
nor U12594 (N_12594,N_8976,N_8285);
and U12595 (N_12595,N_6347,N_5981);
nor U12596 (N_12596,N_9120,N_7917);
or U12597 (N_12597,N_7361,N_8668);
nand U12598 (N_12598,N_6679,N_6389);
xnor U12599 (N_12599,N_8171,N_6752);
nor U12600 (N_12600,N_5868,N_6150);
or U12601 (N_12601,N_9334,N_6338);
or U12602 (N_12602,N_8669,N_8261);
or U12603 (N_12603,N_9266,N_7196);
or U12604 (N_12604,N_6963,N_6536);
xor U12605 (N_12605,N_8275,N_8776);
nor U12606 (N_12606,N_6784,N_8189);
nor U12607 (N_12607,N_5226,N_6750);
nor U12608 (N_12608,N_8102,N_5708);
nor U12609 (N_12609,N_6010,N_7088);
nor U12610 (N_12610,N_7292,N_9641);
nand U12611 (N_12611,N_6471,N_9251);
nand U12612 (N_12612,N_5185,N_9000);
and U12613 (N_12613,N_9873,N_6066);
xnor U12614 (N_12614,N_5441,N_6108);
or U12615 (N_12615,N_5655,N_9355);
xnor U12616 (N_12616,N_7032,N_9642);
xnor U12617 (N_12617,N_5073,N_9740);
or U12618 (N_12618,N_5801,N_9252);
or U12619 (N_12619,N_8731,N_8502);
xor U12620 (N_12620,N_6832,N_6738);
and U12621 (N_12621,N_6912,N_7751);
or U12622 (N_12622,N_5427,N_9994);
nand U12623 (N_12623,N_9721,N_5373);
and U12624 (N_12624,N_7654,N_7233);
nand U12625 (N_12625,N_7573,N_6197);
and U12626 (N_12626,N_5743,N_7757);
nor U12627 (N_12627,N_9627,N_6034);
and U12628 (N_12628,N_5017,N_5205);
xor U12629 (N_12629,N_8729,N_5557);
xnor U12630 (N_12630,N_9265,N_5028);
nand U12631 (N_12631,N_8841,N_5832);
and U12632 (N_12632,N_9115,N_8801);
and U12633 (N_12633,N_8267,N_5369);
and U12634 (N_12634,N_9252,N_7565);
and U12635 (N_12635,N_9416,N_5262);
nand U12636 (N_12636,N_5014,N_7605);
nor U12637 (N_12637,N_7038,N_6758);
nor U12638 (N_12638,N_5468,N_9445);
nand U12639 (N_12639,N_5873,N_8719);
and U12640 (N_12640,N_5393,N_6131);
or U12641 (N_12641,N_6950,N_9689);
nor U12642 (N_12642,N_5610,N_5373);
and U12643 (N_12643,N_7577,N_7878);
or U12644 (N_12644,N_9659,N_9835);
xor U12645 (N_12645,N_9086,N_9089);
xnor U12646 (N_12646,N_6723,N_5539);
xor U12647 (N_12647,N_6294,N_7038);
nor U12648 (N_12648,N_9983,N_6250);
xnor U12649 (N_12649,N_9626,N_8107);
and U12650 (N_12650,N_7246,N_9071);
nor U12651 (N_12651,N_7302,N_8738);
nand U12652 (N_12652,N_8066,N_8767);
and U12653 (N_12653,N_7858,N_6256);
nand U12654 (N_12654,N_7025,N_7902);
nand U12655 (N_12655,N_9464,N_8540);
xnor U12656 (N_12656,N_5393,N_8513);
and U12657 (N_12657,N_5721,N_6285);
nor U12658 (N_12658,N_7226,N_7064);
or U12659 (N_12659,N_8102,N_7825);
nor U12660 (N_12660,N_8758,N_5363);
xnor U12661 (N_12661,N_6849,N_8503);
nor U12662 (N_12662,N_8795,N_9976);
xor U12663 (N_12663,N_9995,N_6141);
and U12664 (N_12664,N_7311,N_8417);
or U12665 (N_12665,N_5582,N_5934);
nand U12666 (N_12666,N_8675,N_6018);
nor U12667 (N_12667,N_8086,N_8775);
or U12668 (N_12668,N_8126,N_9873);
or U12669 (N_12669,N_9061,N_6551);
or U12670 (N_12670,N_8219,N_8413);
xnor U12671 (N_12671,N_9171,N_9124);
nand U12672 (N_12672,N_6514,N_5896);
and U12673 (N_12673,N_6139,N_5357);
nor U12674 (N_12674,N_9316,N_5396);
or U12675 (N_12675,N_7025,N_8062);
and U12676 (N_12676,N_5483,N_5419);
nand U12677 (N_12677,N_9064,N_9781);
or U12678 (N_12678,N_9397,N_6017);
or U12679 (N_12679,N_6319,N_6210);
and U12680 (N_12680,N_7103,N_5508);
and U12681 (N_12681,N_8084,N_9771);
and U12682 (N_12682,N_7292,N_7391);
and U12683 (N_12683,N_6772,N_8689);
nand U12684 (N_12684,N_5539,N_5531);
and U12685 (N_12685,N_5443,N_7099);
or U12686 (N_12686,N_7960,N_7173);
nand U12687 (N_12687,N_6209,N_6655);
or U12688 (N_12688,N_9831,N_6643);
nor U12689 (N_12689,N_8975,N_5470);
xor U12690 (N_12690,N_9899,N_7036);
or U12691 (N_12691,N_8891,N_5144);
nand U12692 (N_12692,N_9615,N_7461);
or U12693 (N_12693,N_7994,N_8670);
nand U12694 (N_12694,N_9809,N_9487);
or U12695 (N_12695,N_5671,N_7813);
and U12696 (N_12696,N_9017,N_6045);
nor U12697 (N_12697,N_7580,N_9770);
nand U12698 (N_12698,N_5432,N_9523);
and U12699 (N_12699,N_7144,N_8289);
nand U12700 (N_12700,N_8793,N_6534);
xor U12701 (N_12701,N_8291,N_5836);
xor U12702 (N_12702,N_5859,N_9344);
xnor U12703 (N_12703,N_5746,N_9126);
nor U12704 (N_12704,N_5015,N_9028);
nand U12705 (N_12705,N_8661,N_6460);
and U12706 (N_12706,N_7747,N_9959);
xnor U12707 (N_12707,N_6409,N_6892);
and U12708 (N_12708,N_8481,N_9569);
and U12709 (N_12709,N_5541,N_6821);
or U12710 (N_12710,N_9296,N_9750);
xor U12711 (N_12711,N_9566,N_8514);
or U12712 (N_12712,N_7224,N_8892);
and U12713 (N_12713,N_7154,N_8378);
or U12714 (N_12714,N_7927,N_7807);
and U12715 (N_12715,N_5303,N_5217);
nand U12716 (N_12716,N_9512,N_5641);
nand U12717 (N_12717,N_6202,N_5961);
xnor U12718 (N_12718,N_9112,N_9234);
or U12719 (N_12719,N_9994,N_7589);
nor U12720 (N_12720,N_8994,N_5346);
or U12721 (N_12721,N_7880,N_9283);
nor U12722 (N_12722,N_8034,N_7638);
nand U12723 (N_12723,N_9717,N_8785);
nand U12724 (N_12724,N_5188,N_7560);
or U12725 (N_12725,N_7718,N_6330);
or U12726 (N_12726,N_8082,N_8070);
nor U12727 (N_12727,N_6948,N_9397);
nor U12728 (N_12728,N_7392,N_6500);
or U12729 (N_12729,N_7469,N_8085);
and U12730 (N_12730,N_8065,N_6531);
nand U12731 (N_12731,N_7921,N_5508);
nor U12732 (N_12732,N_6317,N_9366);
nor U12733 (N_12733,N_8673,N_7957);
nor U12734 (N_12734,N_9273,N_6127);
or U12735 (N_12735,N_6596,N_5295);
xnor U12736 (N_12736,N_7391,N_6486);
xor U12737 (N_12737,N_7860,N_5834);
and U12738 (N_12738,N_5982,N_6714);
nand U12739 (N_12739,N_6851,N_5412);
and U12740 (N_12740,N_6384,N_5856);
and U12741 (N_12741,N_7656,N_7375);
xor U12742 (N_12742,N_9223,N_6765);
and U12743 (N_12743,N_8673,N_8254);
or U12744 (N_12744,N_9424,N_8949);
or U12745 (N_12745,N_9787,N_6782);
or U12746 (N_12746,N_6090,N_5311);
nor U12747 (N_12747,N_6983,N_5019);
nor U12748 (N_12748,N_7388,N_6683);
xnor U12749 (N_12749,N_9483,N_7155);
xor U12750 (N_12750,N_8247,N_8273);
xor U12751 (N_12751,N_9341,N_7882);
and U12752 (N_12752,N_9525,N_9168);
or U12753 (N_12753,N_8602,N_8527);
and U12754 (N_12754,N_9140,N_9474);
nor U12755 (N_12755,N_8674,N_5138);
xnor U12756 (N_12756,N_9489,N_9360);
nand U12757 (N_12757,N_6076,N_5101);
and U12758 (N_12758,N_8699,N_7539);
xor U12759 (N_12759,N_5162,N_7787);
or U12760 (N_12760,N_5245,N_5221);
xor U12761 (N_12761,N_7919,N_6728);
xnor U12762 (N_12762,N_7446,N_5548);
nand U12763 (N_12763,N_5301,N_6969);
nand U12764 (N_12764,N_7614,N_7853);
nor U12765 (N_12765,N_7657,N_5167);
nor U12766 (N_12766,N_6999,N_8329);
and U12767 (N_12767,N_9571,N_9526);
xor U12768 (N_12768,N_8622,N_8751);
xnor U12769 (N_12769,N_9550,N_7627);
nand U12770 (N_12770,N_5309,N_6230);
xor U12771 (N_12771,N_6911,N_6113);
and U12772 (N_12772,N_6547,N_5203);
nor U12773 (N_12773,N_5077,N_6003);
nor U12774 (N_12774,N_5189,N_8656);
nand U12775 (N_12775,N_8635,N_9938);
nor U12776 (N_12776,N_7403,N_8508);
and U12777 (N_12777,N_6751,N_8910);
or U12778 (N_12778,N_7905,N_7545);
xor U12779 (N_12779,N_7434,N_6730);
xor U12780 (N_12780,N_7272,N_9720);
or U12781 (N_12781,N_8026,N_8573);
nor U12782 (N_12782,N_8245,N_5756);
nand U12783 (N_12783,N_7788,N_9179);
and U12784 (N_12784,N_6661,N_5405);
and U12785 (N_12785,N_8856,N_9372);
and U12786 (N_12786,N_7465,N_7708);
or U12787 (N_12787,N_9494,N_8394);
nand U12788 (N_12788,N_8398,N_5706);
or U12789 (N_12789,N_7599,N_9390);
nand U12790 (N_12790,N_6717,N_9882);
xor U12791 (N_12791,N_8424,N_9148);
and U12792 (N_12792,N_7624,N_6127);
nor U12793 (N_12793,N_5176,N_5544);
nor U12794 (N_12794,N_9644,N_8350);
xor U12795 (N_12795,N_7020,N_7019);
or U12796 (N_12796,N_6496,N_9888);
and U12797 (N_12797,N_8911,N_6741);
nor U12798 (N_12798,N_6463,N_6929);
and U12799 (N_12799,N_9369,N_7916);
nand U12800 (N_12800,N_7313,N_6060);
xor U12801 (N_12801,N_7960,N_7379);
nand U12802 (N_12802,N_8714,N_5831);
xor U12803 (N_12803,N_8349,N_5026);
xnor U12804 (N_12804,N_9058,N_6787);
nand U12805 (N_12805,N_9344,N_8347);
nand U12806 (N_12806,N_7564,N_5768);
nand U12807 (N_12807,N_5511,N_9128);
xnor U12808 (N_12808,N_9066,N_8939);
and U12809 (N_12809,N_6155,N_6144);
nor U12810 (N_12810,N_9972,N_7480);
nand U12811 (N_12811,N_9316,N_8319);
xnor U12812 (N_12812,N_6481,N_8186);
xnor U12813 (N_12813,N_8062,N_5672);
nand U12814 (N_12814,N_8244,N_7376);
or U12815 (N_12815,N_7944,N_9943);
and U12816 (N_12816,N_8353,N_5689);
nand U12817 (N_12817,N_8429,N_9661);
nand U12818 (N_12818,N_5572,N_7439);
or U12819 (N_12819,N_8331,N_6686);
and U12820 (N_12820,N_5287,N_6353);
nor U12821 (N_12821,N_7466,N_9702);
and U12822 (N_12822,N_8389,N_7376);
and U12823 (N_12823,N_6619,N_9640);
xor U12824 (N_12824,N_7404,N_8236);
or U12825 (N_12825,N_6773,N_7969);
nand U12826 (N_12826,N_7902,N_9005);
and U12827 (N_12827,N_9431,N_5062);
nand U12828 (N_12828,N_5708,N_6847);
and U12829 (N_12829,N_8289,N_8216);
nand U12830 (N_12830,N_6090,N_9484);
nor U12831 (N_12831,N_6664,N_8109);
xor U12832 (N_12832,N_6373,N_7209);
or U12833 (N_12833,N_7847,N_9644);
or U12834 (N_12834,N_5535,N_5797);
xor U12835 (N_12835,N_5090,N_8518);
and U12836 (N_12836,N_6689,N_9608);
nand U12837 (N_12837,N_6372,N_7782);
xor U12838 (N_12838,N_8593,N_6556);
xor U12839 (N_12839,N_9707,N_7261);
nand U12840 (N_12840,N_8671,N_5133);
nor U12841 (N_12841,N_7064,N_5999);
xor U12842 (N_12842,N_7333,N_9333);
and U12843 (N_12843,N_5937,N_9399);
xnor U12844 (N_12844,N_8753,N_6476);
and U12845 (N_12845,N_5721,N_9208);
nand U12846 (N_12846,N_8310,N_6719);
nand U12847 (N_12847,N_8058,N_8245);
nand U12848 (N_12848,N_6057,N_8170);
or U12849 (N_12849,N_6975,N_5721);
and U12850 (N_12850,N_8179,N_7787);
and U12851 (N_12851,N_9727,N_9715);
or U12852 (N_12852,N_8050,N_5013);
nand U12853 (N_12853,N_7358,N_8412);
and U12854 (N_12854,N_7632,N_5163);
and U12855 (N_12855,N_8125,N_7644);
nand U12856 (N_12856,N_5781,N_9724);
nand U12857 (N_12857,N_6169,N_7178);
xnor U12858 (N_12858,N_5848,N_9092);
or U12859 (N_12859,N_8787,N_9392);
nor U12860 (N_12860,N_7894,N_8497);
nand U12861 (N_12861,N_7072,N_9811);
and U12862 (N_12862,N_6041,N_7296);
xor U12863 (N_12863,N_7672,N_5678);
and U12864 (N_12864,N_7568,N_7838);
nand U12865 (N_12865,N_9730,N_7419);
or U12866 (N_12866,N_8524,N_6712);
xor U12867 (N_12867,N_9975,N_5716);
nand U12868 (N_12868,N_8560,N_6728);
xor U12869 (N_12869,N_6493,N_5282);
and U12870 (N_12870,N_8532,N_9333);
and U12871 (N_12871,N_8816,N_5740);
xor U12872 (N_12872,N_9773,N_8979);
or U12873 (N_12873,N_5749,N_7561);
nand U12874 (N_12874,N_9773,N_5804);
and U12875 (N_12875,N_6326,N_6961);
xor U12876 (N_12876,N_9809,N_6729);
and U12877 (N_12877,N_8290,N_8326);
and U12878 (N_12878,N_7189,N_6643);
nor U12879 (N_12879,N_9087,N_7413);
nor U12880 (N_12880,N_9703,N_9882);
and U12881 (N_12881,N_5497,N_9224);
nor U12882 (N_12882,N_9873,N_9518);
nand U12883 (N_12883,N_7377,N_9973);
and U12884 (N_12884,N_7920,N_5600);
and U12885 (N_12885,N_7556,N_7685);
xor U12886 (N_12886,N_8270,N_5555);
nor U12887 (N_12887,N_7469,N_7510);
nand U12888 (N_12888,N_6881,N_5093);
nor U12889 (N_12889,N_5330,N_5792);
nor U12890 (N_12890,N_5484,N_7937);
and U12891 (N_12891,N_9447,N_5625);
and U12892 (N_12892,N_5007,N_6508);
nor U12893 (N_12893,N_9572,N_9012);
xor U12894 (N_12894,N_6767,N_8020);
nand U12895 (N_12895,N_5489,N_7765);
or U12896 (N_12896,N_6409,N_5812);
nand U12897 (N_12897,N_8027,N_9716);
nor U12898 (N_12898,N_8674,N_9672);
nor U12899 (N_12899,N_6758,N_5436);
nand U12900 (N_12900,N_9740,N_7938);
or U12901 (N_12901,N_5228,N_7673);
nand U12902 (N_12902,N_6747,N_7634);
xor U12903 (N_12903,N_5505,N_7637);
or U12904 (N_12904,N_8333,N_8582);
and U12905 (N_12905,N_6251,N_8640);
nand U12906 (N_12906,N_7131,N_6173);
nand U12907 (N_12907,N_7124,N_9252);
and U12908 (N_12908,N_5965,N_5764);
nor U12909 (N_12909,N_7247,N_6180);
xnor U12910 (N_12910,N_9572,N_6228);
or U12911 (N_12911,N_6763,N_7645);
nor U12912 (N_12912,N_9195,N_9027);
nand U12913 (N_12913,N_9932,N_6821);
nand U12914 (N_12914,N_5286,N_7109);
nand U12915 (N_12915,N_9144,N_5968);
nand U12916 (N_12916,N_8246,N_9048);
or U12917 (N_12917,N_6464,N_6297);
nor U12918 (N_12918,N_7775,N_7710);
nand U12919 (N_12919,N_8928,N_6328);
or U12920 (N_12920,N_9156,N_5129);
and U12921 (N_12921,N_8009,N_7535);
nand U12922 (N_12922,N_8661,N_6825);
nor U12923 (N_12923,N_7125,N_8475);
xor U12924 (N_12924,N_6523,N_5551);
nor U12925 (N_12925,N_7354,N_6446);
nand U12926 (N_12926,N_9212,N_9516);
nor U12927 (N_12927,N_6869,N_8860);
or U12928 (N_12928,N_7806,N_5131);
or U12929 (N_12929,N_6363,N_5906);
xnor U12930 (N_12930,N_9742,N_9704);
nor U12931 (N_12931,N_7921,N_8137);
or U12932 (N_12932,N_7318,N_5551);
and U12933 (N_12933,N_7043,N_9334);
or U12934 (N_12934,N_8683,N_8311);
xor U12935 (N_12935,N_7901,N_8654);
nor U12936 (N_12936,N_8372,N_8476);
or U12937 (N_12937,N_6809,N_5720);
nand U12938 (N_12938,N_6369,N_6447);
or U12939 (N_12939,N_9489,N_6325);
nor U12940 (N_12940,N_9619,N_9070);
and U12941 (N_12941,N_9105,N_7185);
or U12942 (N_12942,N_6389,N_6884);
nand U12943 (N_12943,N_8384,N_6517);
nand U12944 (N_12944,N_7707,N_6613);
xnor U12945 (N_12945,N_7385,N_7664);
nor U12946 (N_12946,N_5952,N_9500);
nor U12947 (N_12947,N_7724,N_9840);
and U12948 (N_12948,N_5763,N_5794);
or U12949 (N_12949,N_7995,N_5914);
nor U12950 (N_12950,N_8797,N_9386);
or U12951 (N_12951,N_7936,N_6463);
nor U12952 (N_12952,N_6639,N_9614);
nand U12953 (N_12953,N_5174,N_9004);
and U12954 (N_12954,N_5953,N_7706);
xnor U12955 (N_12955,N_6160,N_8424);
xor U12956 (N_12956,N_9884,N_6774);
nor U12957 (N_12957,N_8764,N_9486);
nand U12958 (N_12958,N_6302,N_8958);
and U12959 (N_12959,N_9794,N_5377);
nand U12960 (N_12960,N_5749,N_6228);
and U12961 (N_12961,N_5413,N_9863);
nand U12962 (N_12962,N_6499,N_9839);
nand U12963 (N_12963,N_8676,N_8133);
nor U12964 (N_12964,N_6962,N_6385);
or U12965 (N_12965,N_8465,N_9246);
xnor U12966 (N_12966,N_8138,N_6837);
and U12967 (N_12967,N_6995,N_9261);
nand U12968 (N_12968,N_5761,N_6905);
nor U12969 (N_12969,N_9149,N_8199);
and U12970 (N_12970,N_7606,N_8719);
nor U12971 (N_12971,N_9817,N_7336);
and U12972 (N_12972,N_9228,N_8672);
xor U12973 (N_12973,N_6542,N_8653);
or U12974 (N_12974,N_6911,N_5369);
or U12975 (N_12975,N_9367,N_8038);
nor U12976 (N_12976,N_9630,N_8330);
or U12977 (N_12977,N_8764,N_5498);
nor U12978 (N_12978,N_5931,N_8647);
and U12979 (N_12979,N_6023,N_9188);
nand U12980 (N_12980,N_7232,N_6743);
nor U12981 (N_12981,N_5310,N_5400);
and U12982 (N_12982,N_6994,N_8328);
or U12983 (N_12983,N_8233,N_8726);
or U12984 (N_12984,N_8038,N_7032);
or U12985 (N_12985,N_7977,N_8600);
nor U12986 (N_12986,N_8466,N_6323);
xor U12987 (N_12987,N_6080,N_7268);
nor U12988 (N_12988,N_9406,N_7206);
nor U12989 (N_12989,N_5956,N_9462);
nand U12990 (N_12990,N_8559,N_8091);
or U12991 (N_12991,N_8706,N_7073);
or U12992 (N_12992,N_6036,N_5573);
nor U12993 (N_12993,N_5810,N_5953);
and U12994 (N_12994,N_6758,N_6241);
nor U12995 (N_12995,N_9359,N_6777);
xnor U12996 (N_12996,N_7934,N_8203);
and U12997 (N_12997,N_9524,N_8207);
and U12998 (N_12998,N_7930,N_5998);
xnor U12999 (N_12999,N_9212,N_9384);
and U13000 (N_13000,N_5044,N_8263);
or U13001 (N_13001,N_8202,N_8047);
xnor U13002 (N_13002,N_5078,N_5700);
nand U13003 (N_13003,N_7197,N_8086);
and U13004 (N_13004,N_8593,N_8186);
nor U13005 (N_13005,N_7240,N_8854);
or U13006 (N_13006,N_6781,N_7070);
nand U13007 (N_13007,N_7565,N_8115);
xnor U13008 (N_13008,N_7145,N_5901);
or U13009 (N_13009,N_9988,N_8775);
and U13010 (N_13010,N_9004,N_5916);
or U13011 (N_13011,N_5124,N_6374);
or U13012 (N_13012,N_9976,N_6965);
and U13013 (N_13013,N_8234,N_8274);
or U13014 (N_13014,N_6936,N_7807);
and U13015 (N_13015,N_7158,N_8455);
xor U13016 (N_13016,N_8364,N_5537);
and U13017 (N_13017,N_6683,N_9674);
or U13018 (N_13018,N_8099,N_6602);
xnor U13019 (N_13019,N_8402,N_8936);
or U13020 (N_13020,N_7106,N_9019);
or U13021 (N_13021,N_7073,N_9425);
nand U13022 (N_13022,N_6381,N_9812);
nand U13023 (N_13023,N_7021,N_5197);
nor U13024 (N_13024,N_9725,N_7107);
xor U13025 (N_13025,N_6687,N_6416);
and U13026 (N_13026,N_6732,N_8922);
and U13027 (N_13027,N_9763,N_5759);
xor U13028 (N_13028,N_5520,N_9923);
or U13029 (N_13029,N_7180,N_8656);
nand U13030 (N_13030,N_7530,N_8600);
xor U13031 (N_13031,N_6212,N_8572);
and U13032 (N_13032,N_7631,N_7704);
xnor U13033 (N_13033,N_9096,N_8000);
nor U13034 (N_13034,N_7504,N_7554);
or U13035 (N_13035,N_5966,N_5487);
or U13036 (N_13036,N_7539,N_9541);
nor U13037 (N_13037,N_9949,N_6112);
nand U13038 (N_13038,N_5402,N_8257);
xnor U13039 (N_13039,N_5436,N_7340);
nor U13040 (N_13040,N_8667,N_5834);
nand U13041 (N_13041,N_7089,N_7407);
xor U13042 (N_13042,N_8430,N_9633);
nand U13043 (N_13043,N_8859,N_8293);
and U13044 (N_13044,N_5358,N_8202);
or U13045 (N_13045,N_6664,N_9585);
xnor U13046 (N_13046,N_5487,N_5085);
nand U13047 (N_13047,N_6752,N_5154);
or U13048 (N_13048,N_7232,N_9840);
and U13049 (N_13049,N_9289,N_7233);
nand U13050 (N_13050,N_8812,N_5953);
and U13051 (N_13051,N_5632,N_9075);
nor U13052 (N_13052,N_8774,N_5750);
nor U13053 (N_13053,N_8270,N_8137);
nand U13054 (N_13054,N_6863,N_8502);
or U13055 (N_13055,N_7875,N_7054);
and U13056 (N_13056,N_9704,N_7348);
and U13057 (N_13057,N_9061,N_8020);
xor U13058 (N_13058,N_5965,N_7919);
xor U13059 (N_13059,N_9400,N_5020);
and U13060 (N_13060,N_9291,N_7309);
nor U13061 (N_13061,N_7849,N_6632);
xnor U13062 (N_13062,N_9253,N_8574);
nor U13063 (N_13063,N_5472,N_8852);
or U13064 (N_13064,N_8789,N_9614);
or U13065 (N_13065,N_8422,N_8737);
and U13066 (N_13066,N_9165,N_6422);
nand U13067 (N_13067,N_8342,N_9415);
xnor U13068 (N_13068,N_9659,N_6781);
and U13069 (N_13069,N_8603,N_6950);
and U13070 (N_13070,N_6771,N_6011);
or U13071 (N_13071,N_8490,N_8107);
nand U13072 (N_13072,N_8438,N_5427);
and U13073 (N_13073,N_9115,N_7329);
nand U13074 (N_13074,N_9746,N_9929);
nor U13075 (N_13075,N_6541,N_5412);
nand U13076 (N_13076,N_8727,N_7003);
or U13077 (N_13077,N_9324,N_6542);
and U13078 (N_13078,N_9829,N_7434);
or U13079 (N_13079,N_9329,N_6997);
or U13080 (N_13080,N_8147,N_9065);
nor U13081 (N_13081,N_9726,N_6216);
nand U13082 (N_13082,N_6142,N_6447);
or U13083 (N_13083,N_5283,N_9848);
nand U13084 (N_13084,N_7311,N_6247);
xnor U13085 (N_13085,N_9582,N_9350);
nand U13086 (N_13086,N_7684,N_5800);
xor U13087 (N_13087,N_7684,N_6990);
and U13088 (N_13088,N_6345,N_5790);
and U13089 (N_13089,N_8688,N_6310);
or U13090 (N_13090,N_6029,N_8493);
and U13091 (N_13091,N_9555,N_9295);
nor U13092 (N_13092,N_9599,N_5281);
or U13093 (N_13093,N_8922,N_9384);
or U13094 (N_13094,N_7940,N_8393);
xor U13095 (N_13095,N_8181,N_9109);
or U13096 (N_13096,N_5133,N_5854);
or U13097 (N_13097,N_9457,N_8815);
nor U13098 (N_13098,N_9028,N_8223);
nand U13099 (N_13099,N_9954,N_8645);
or U13100 (N_13100,N_9081,N_8313);
and U13101 (N_13101,N_6986,N_9345);
nor U13102 (N_13102,N_5516,N_8603);
nand U13103 (N_13103,N_7613,N_7561);
and U13104 (N_13104,N_8642,N_5243);
nor U13105 (N_13105,N_8031,N_8887);
nand U13106 (N_13106,N_5728,N_6430);
and U13107 (N_13107,N_5828,N_5758);
and U13108 (N_13108,N_5677,N_8731);
and U13109 (N_13109,N_5439,N_7767);
and U13110 (N_13110,N_8746,N_7020);
nor U13111 (N_13111,N_9948,N_6585);
xor U13112 (N_13112,N_6993,N_7983);
nor U13113 (N_13113,N_9278,N_5201);
or U13114 (N_13114,N_6075,N_6087);
nor U13115 (N_13115,N_8146,N_8333);
nor U13116 (N_13116,N_7670,N_8167);
xnor U13117 (N_13117,N_7027,N_6283);
or U13118 (N_13118,N_8327,N_8251);
xnor U13119 (N_13119,N_7018,N_8999);
xnor U13120 (N_13120,N_7991,N_9293);
or U13121 (N_13121,N_6520,N_5950);
and U13122 (N_13122,N_7812,N_8880);
or U13123 (N_13123,N_9024,N_7160);
nand U13124 (N_13124,N_8196,N_5035);
and U13125 (N_13125,N_5168,N_5286);
xor U13126 (N_13126,N_6807,N_6149);
or U13127 (N_13127,N_8490,N_7087);
nand U13128 (N_13128,N_9707,N_9055);
or U13129 (N_13129,N_7448,N_8087);
and U13130 (N_13130,N_5598,N_9691);
xor U13131 (N_13131,N_5272,N_7053);
or U13132 (N_13132,N_6611,N_6605);
nand U13133 (N_13133,N_9139,N_7186);
and U13134 (N_13134,N_6009,N_7630);
and U13135 (N_13135,N_7854,N_5775);
nor U13136 (N_13136,N_7133,N_5518);
nor U13137 (N_13137,N_8186,N_6925);
or U13138 (N_13138,N_5438,N_5192);
nor U13139 (N_13139,N_7779,N_9210);
nor U13140 (N_13140,N_7384,N_7338);
nor U13141 (N_13141,N_9701,N_5988);
nand U13142 (N_13142,N_6370,N_6098);
nand U13143 (N_13143,N_7575,N_7552);
nor U13144 (N_13144,N_8052,N_6183);
and U13145 (N_13145,N_7017,N_5118);
or U13146 (N_13146,N_9914,N_5586);
xor U13147 (N_13147,N_9620,N_9333);
xnor U13148 (N_13148,N_9648,N_6503);
or U13149 (N_13149,N_5607,N_6354);
or U13150 (N_13150,N_6956,N_5413);
and U13151 (N_13151,N_8218,N_8870);
xnor U13152 (N_13152,N_9316,N_5344);
xnor U13153 (N_13153,N_5087,N_9444);
nand U13154 (N_13154,N_5550,N_7949);
xor U13155 (N_13155,N_6996,N_5822);
nor U13156 (N_13156,N_9427,N_9451);
nand U13157 (N_13157,N_8118,N_6671);
and U13158 (N_13158,N_7590,N_8467);
nor U13159 (N_13159,N_8577,N_9451);
xnor U13160 (N_13160,N_9503,N_9990);
or U13161 (N_13161,N_9320,N_5053);
nand U13162 (N_13162,N_6737,N_5185);
and U13163 (N_13163,N_6068,N_8570);
nand U13164 (N_13164,N_8710,N_7927);
or U13165 (N_13165,N_8302,N_5032);
and U13166 (N_13166,N_7267,N_6838);
xnor U13167 (N_13167,N_9270,N_6100);
and U13168 (N_13168,N_7706,N_6875);
nor U13169 (N_13169,N_8050,N_8234);
or U13170 (N_13170,N_9716,N_5979);
nor U13171 (N_13171,N_9797,N_6793);
or U13172 (N_13172,N_7639,N_6270);
nand U13173 (N_13173,N_6892,N_8031);
or U13174 (N_13174,N_7355,N_5098);
nand U13175 (N_13175,N_5242,N_9550);
or U13176 (N_13176,N_7910,N_5488);
xnor U13177 (N_13177,N_8324,N_5039);
xnor U13178 (N_13178,N_6532,N_8387);
or U13179 (N_13179,N_6386,N_6982);
xnor U13180 (N_13180,N_7418,N_5812);
or U13181 (N_13181,N_5924,N_7982);
nand U13182 (N_13182,N_8089,N_9810);
xnor U13183 (N_13183,N_8674,N_6734);
or U13184 (N_13184,N_7984,N_8226);
xor U13185 (N_13185,N_5217,N_7704);
nor U13186 (N_13186,N_5891,N_9076);
nor U13187 (N_13187,N_8162,N_7036);
or U13188 (N_13188,N_9246,N_8584);
or U13189 (N_13189,N_9729,N_8298);
or U13190 (N_13190,N_9975,N_6288);
nor U13191 (N_13191,N_6979,N_8209);
or U13192 (N_13192,N_6392,N_7417);
and U13193 (N_13193,N_9831,N_8819);
nor U13194 (N_13194,N_8886,N_8042);
nand U13195 (N_13195,N_9200,N_8906);
xor U13196 (N_13196,N_8696,N_7439);
or U13197 (N_13197,N_8762,N_6260);
nand U13198 (N_13198,N_8249,N_8095);
or U13199 (N_13199,N_8064,N_9864);
and U13200 (N_13200,N_6334,N_8971);
nand U13201 (N_13201,N_5140,N_6442);
xnor U13202 (N_13202,N_6176,N_6683);
nand U13203 (N_13203,N_6258,N_6593);
xnor U13204 (N_13204,N_7013,N_9585);
nand U13205 (N_13205,N_8186,N_9921);
and U13206 (N_13206,N_9553,N_5427);
nand U13207 (N_13207,N_6998,N_8456);
nand U13208 (N_13208,N_8057,N_6484);
xor U13209 (N_13209,N_8529,N_9046);
nor U13210 (N_13210,N_9977,N_7144);
xor U13211 (N_13211,N_7646,N_7084);
and U13212 (N_13212,N_7835,N_9378);
and U13213 (N_13213,N_6428,N_8486);
and U13214 (N_13214,N_7688,N_9823);
nor U13215 (N_13215,N_5916,N_8178);
nand U13216 (N_13216,N_8036,N_7219);
xnor U13217 (N_13217,N_8558,N_8417);
nor U13218 (N_13218,N_7189,N_9718);
or U13219 (N_13219,N_7054,N_9384);
nor U13220 (N_13220,N_7436,N_8219);
and U13221 (N_13221,N_8942,N_8684);
nor U13222 (N_13222,N_8342,N_5475);
nand U13223 (N_13223,N_7603,N_9131);
nand U13224 (N_13224,N_9050,N_5009);
nor U13225 (N_13225,N_5460,N_8703);
and U13226 (N_13226,N_7153,N_5622);
nand U13227 (N_13227,N_9063,N_9094);
and U13228 (N_13228,N_9002,N_9067);
and U13229 (N_13229,N_6234,N_9485);
nor U13230 (N_13230,N_9783,N_8218);
and U13231 (N_13231,N_6688,N_5630);
nand U13232 (N_13232,N_7723,N_5362);
and U13233 (N_13233,N_9196,N_7234);
nand U13234 (N_13234,N_9825,N_9833);
xnor U13235 (N_13235,N_5975,N_5184);
xor U13236 (N_13236,N_5380,N_6771);
or U13237 (N_13237,N_6347,N_6920);
and U13238 (N_13238,N_8306,N_7577);
nand U13239 (N_13239,N_9939,N_9738);
xor U13240 (N_13240,N_8947,N_9110);
nand U13241 (N_13241,N_6445,N_9563);
nor U13242 (N_13242,N_9693,N_7881);
nor U13243 (N_13243,N_8604,N_7339);
xor U13244 (N_13244,N_6933,N_7358);
or U13245 (N_13245,N_5511,N_5207);
and U13246 (N_13246,N_8817,N_9943);
nor U13247 (N_13247,N_8428,N_8458);
xor U13248 (N_13248,N_7451,N_5865);
nand U13249 (N_13249,N_6089,N_7554);
nand U13250 (N_13250,N_7571,N_7513);
and U13251 (N_13251,N_6913,N_5727);
nand U13252 (N_13252,N_9680,N_9300);
nand U13253 (N_13253,N_6079,N_9611);
xor U13254 (N_13254,N_6638,N_6369);
or U13255 (N_13255,N_5658,N_8339);
nor U13256 (N_13256,N_5397,N_9543);
and U13257 (N_13257,N_6846,N_5725);
xnor U13258 (N_13258,N_8526,N_8149);
nand U13259 (N_13259,N_7702,N_5075);
nand U13260 (N_13260,N_7499,N_9324);
and U13261 (N_13261,N_5915,N_6222);
nor U13262 (N_13262,N_5633,N_8302);
and U13263 (N_13263,N_5532,N_5129);
xnor U13264 (N_13264,N_8679,N_7065);
xor U13265 (N_13265,N_6434,N_5630);
nand U13266 (N_13266,N_9449,N_8484);
nand U13267 (N_13267,N_6967,N_5865);
and U13268 (N_13268,N_9839,N_7747);
or U13269 (N_13269,N_5933,N_5715);
or U13270 (N_13270,N_7746,N_9574);
nor U13271 (N_13271,N_6998,N_7808);
or U13272 (N_13272,N_8342,N_5058);
nand U13273 (N_13273,N_6850,N_7766);
or U13274 (N_13274,N_5393,N_5271);
xor U13275 (N_13275,N_9220,N_5648);
nor U13276 (N_13276,N_8946,N_8892);
or U13277 (N_13277,N_7263,N_7158);
xnor U13278 (N_13278,N_7873,N_5397);
nor U13279 (N_13279,N_5698,N_8068);
and U13280 (N_13280,N_9058,N_9536);
nor U13281 (N_13281,N_9031,N_6301);
or U13282 (N_13282,N_7648,N_5242);
or U13283 (N_13283,N_6779,N_5333);
or U13284 (N_13284,N_7148,N_6166);
nand U13285 (N_13285,N_8379,N_8197);
and U13286 (N_13286,N_7495,N_8331);
xor U13287 (N_13287,N_8329,N_6103);
xor U13288 (N_13288,N_9370,N_7914);
nand U13289 (N_13289,N_8602,N_7766);
nand U13290 (N_13290,N_8608,N_7236);
nand U13291 (N_13291,N_8065,N_7696);
xnor U13292 (N_13292,N_9610,N_8899);
nand U13293 (N_13293,N_6776,N_6676);
and U13294 (N_13294,N_5348,N_5645);
nand U13295 (N_13295,N_5096,N_5631);
nand U13296 (N_13296,N_8009,N_5098);
nor U13297 (N_13297,N_8552,N_7813);
and U13298 (N_13298,N_5662,N_6417);
or U13299 (N_13299,N_9937,N_5000);
or U13300 (N_13300,N_7487,N_8472);
and U13301 (N_13301,N_6235,N_7462);
nand U13302 (N_13302,N_7544,N_9605);
xor U13303 (N_13303,N_7213,N_7277);
or U13304 (N_13304,N_8743,N_9008);
nand U13305 (N_13305,N_5405,N_7009);
or U13306 (N_13306,N_9276,N_6847);
xnor U13307 (N_13307,N_6165,N_8451);
xor U13308 (N_13308,N_6382,N_9171);
and U13309 (N_13309,N_6496,N_5920);
nand U13310 (N_13310,N_5962,N_8987);
xor U13311 (N_13311,N_5004,N_6583);
and U13312 (N_13312,N_6647,N_9095);
xor U13313 (N_13313,N_6347,N_5976);
nand U13314 (N_13314,N_7267,N_6134);
nand U13315 (N_13315,N_5299,N_7518);
xor U13316 (N_13316,N_6675,N_6490);
and U13317 (N_13317,N_7676,N_5997);
xnor U13318 (N_13318,N_8803,N_5748);
nor U13319 (N_13319,N_6218,N_6697);
nand U13320 (N_13320,N_9941,N_9804);
or U13321 (N_13321,N_8991,N_5201);
nor U13322 (N_13322,N_9511,N_5203);
xnor U13323 (N_13323,N_8387,N_9208);
nand U13324 (N_13324,N_8188,N_6092);
xnor U13325 (N_13325,N_9910,N_8591);
and U13326 (N_13326,N_8975,N_7717);
nand U13327 (N_13327,N_5706,N_8415);
xor U13328 (N_13328,N_9501,N_5406);
xor U13329 (N_13329,N_5636,N_9832);
nor U13330 (N_13330,N_6032,N_9860);
nor U13331 (N_13331,N_8690,N_8659);
nand U13332 (N_13332,N_5331,N_6516);
or U13333 (N_13333,N_9420,N_9759);
or U13334 (N_13334,N_9214,N_7464);
nand U13335 (N_13335,N_9484,N_5719);
or U13336 (N_13336,N_8962,N_9251);
or U13337 (N_13337,N_9867,N_8560);
nand U13338 (N_13338,N_6783,N_5618);
or U13339 (N_13339,N_8042,N_9170);
nor U13340 (N_13340,N_6498,N_7666);
nand U13341 (N_13341,N_8670,N_6649);
and U13342 (N_13342,N_8156,N_5861);
and U13343 (N_13343,N_9832,N_8163);
or U13344 (N_13344,N_8410,N_7311);
and U13345 (N_13345,N_9727,N_5328);
nor U13346 (N_13346,N_6809,N_5517);
nand U13347 (N_13347,N_5977,N_8627);
nand U13348 (N_13348,N_7674,N_8845);
and U13349 (N_13349,N_6136,N_7652);
nor U13350 (N_13350,N_5453,N_8798);
xor U13351 (N_13351,N_6216,N_6394);
and U13352 (N_13352,N_9815,N_6885);
nor U13353 (N_13353,N_7844,N_9703);
xor U13354 (N_13354,N_5154,N_8126);
or U13355 (N_13355,N_8617,N_5645);
xor U13356 (N_13356,N_6689,N_9720);
nand U13357 (N_13357,N_9656,N_8558);
nor U13358 (N_13358,N_7646,N_8517);
nand U13359 (N_13359,N_6592,N_6349);
nor U13360 (N_13360,N_9861,N_5321);
xnor U13361 (N_13361,N_5066,N_6821);
or U13362 (N_13362,N_6536,N_8278);
nor U13363 (N_13363,N_6109,N_5066);
and U13364 (N_13364,N_7375,N_8973);
nor U13365 (N_13365,N_7994,N_8187);
xnor U13366 (N_13366,N_9182,N_6493);
or U13367 (N_13367,N_9931,N_9866);
or U13368 (N_13368,N_8720,N_9619);
xor U13369 (N_13369,N_7627,N_5187);
or U13370 (N_13370,N_8499,N_8189);
xnor U13371 (N_13371,N_6534,N_9555);
and U13372 (N_13372,N_8634,N_9471);
or U13373 (N_13373,N_8240,N_8845);
and U13374 (N_13374,N_5473,N_5345);
or U13375 (N_13375,N_6801,N_7550);
nor U13376 (N_13376,N_5496,N_5824);
or U13377 (N_13377,N_8862,N_7969);
nand U13378 (N_13378,N_8962,N_7323);
and U13379 (N_13379,N_7053,N_5639);
xor U13380 (N_13380,N_7723,N_8580);
nor U13381 (N_13381,N_5656,N_6941);
xor U13382 (N_13382,N_6382,N_5829);
nor U13383 (N_13383,N_9354,N_5661);
xor U13384 (N_13384,N_7505,N_6373);
and U13385 (N_13385,N_7903,N_8879);
nand U13386 (N_13386,N_9922,N_6503);
or U13387 (N_13387,N_5214,N_8662);
nand U13388 (N_13388,N_8563,N_9748);
nand U13389 (N_13389,N_6831,N_5646);
xor U13390 (N_13390,N_8946,N_8007);
nand U13391 (N_13391,N_8553,N_8449);
nor U13392 (N_13392,N_6406,N_9721);
nand U13393 (N_13393,N_7926,N_8093);
and U13394 (N_13394,N_8293,N_9472);
nor U13395 (N_13395,N_9268,N_5890);
nor U13396 (N_13396,N_8109,N_8733);
and U13397 (N_13397,N_7301,N_9074);
and U13398 (N_13398,N_9508,N_8704);
nor U13399 (N_13399,N_8230,N_8407);
nor U13400 (N_13400,N_8210,N_8408);
nand U13401 (N_13401,N_7373,N_7956);
and U13402 (N_13402,N_5265,N_6405);
or U13403 (N_13403,N_9399,N_9424);
nor U13404 (N_13404,N_9520,N_8384);
or U13405 (N_13405,N_8067,N_7119);
and U13406 (N_13406,N_9494,N_7598);
xor U13407 (N_13407,N_9897,N_6649);
and U13408 (N_13408,N_5114,N_5112);
and U13409 (N_13409,N_5086,N_7258);
or U13410 (N_13410,N_7720,N_8333);
xor U13411 (N_13411,N_5635,N_5769);
xor U13412 (N_13412,N_5947,N_9742);
xnor U13413 (N_13413,N_9751,N_6297);
or U13414 (N_13414,N_6451,N_9785);
and U13415 (N_13415,N_5359,N_6479);
nand U13416 (N_13416,N_8231,N_6311);
nor U13417 (N_13417,N_5201,N_6410);
nand U13418 (N_13418,N_6709,N_9205);
nor U13419 (N_13419,N_8325,N_5081);
xor U13420 (N_13420,N_7921,N_6177);
nor U13421 (N_13421,N_7629,N_8010);
xor U13422 (N_13422,N_5514,N_8318);
or U13423 (N_13423,N_6530,N_6044);
or U13424 (N_13424,N_9309,N_7314);
and U13425 (N_13425,N_6924,N_8233);
nand U13426 (N_13426,N_9256,N_6299);
nand U13427 (N_13427,N_6597,N_5155);
xnor U13428 (N_13428,N_9302,N_9053);
or U13429 (N_13429,N_6465,N_5825);
and U13430 (N_13430,N_5423,N_7234);
xor U13431 (N_13431,N_6620,N_8589);
nand U13432 (N_13432,N_9796,N_7374);
xor U13433 (N_13433,N_8854,N_7223);
nand U13434 (N_13434,N_5765,N_7194);
xor U13435 (N_13435,N_6867,N_7704);
nand U13436 (N_13436,N_5844,N_8579);
or U13437 (N_13437,N_9639,N_5212);
nand U13438 (N_13438,N_6408,N_8130);
nor U13439 (N_13439,N_6371,N_5994);
xnor U13440 (N_13440,N_7089,N_9668);
and U13441 (N_13441,N_6700,N_6496);
or U13442 (N_13442,N_5641,N_7117);
nor U13443 (N_13443,N_6639,N_7947);
and U13444 (N_13444,N_8560,N_9748);
or U13445 (N_13445,N_8110,N_6537);
and U13446 (N_13446,N_9656,N_5302);
nor U13447 (N_13447,N_8580,N_6051);
or U13448 (N_13448,N_5709,N_7195);
or U13449 (N_13449,N_5546,N_9523);
xnor U13450 (N_13450,N_9121,N_6285);
nand U13451 (N_13451,N_9488,N_7278);
and U13452 (N_13452,N_7475,N_5433);
and U13453 (N_13453,N_9791,N_9805);
xor U13454 (N_13454,N_9845,N_7826);
nor U13455 (N_13455,N_5126,N_6738);
xor U13456 (N_13456,N_5630,N_8361);
nand U13457 (N_13457,N_7218,N_5605);
and U13458 (N_13458,N_5251,N_9391);
xor U13459 (N_13459,N_9882,N_7854);
nand U13460 (N_13460,N_8681,N_8917);
xor U13461 (N_13461,N_8128,N_6070);
and U13462 (N_13462,N_7380,N_5167);
and U13463 (N_13463,N_7624,N_8047);
and U13464 (N_13464,N_6312,N_8625);
nor U13465 (N_13465,N_8055,N_5696);
or U13466 (N_13466,N_5317,N_9184);
xnor U13467 (N_13467,N_7290,N_8601);
xnor U13468 (N_13468,N_7010,N_5139);
and U13469 (N_13469,N_7950,N_9745);
nand U13470 (N_13470,N_5337,N_8230);
nand U13471 (N_13471,N_9155,N_6970);
nor U13472 (N_13472,N_5694,N_7220);
nand U13473 (N_13473,N_7924,N_7094);
xnor U13474 (N_13474,N_7269,N_9981);
nand U13475 (N_13475,N_7467,N_6980);
nand U13476 (N_13476,N_7156,N_8232);
or U13477 (N_13477,N_5563,N_5094);
nor U13478 (N_13478,N_7646,N_7567);
nor U13479 (N_13479,N_9567,N_8755);
nand U13480 (N_13480,N_6354,N_6641);
nand U13481 (N_13481,N_7989,N_8469);
nand U13482 (N_13482,N_5125,N_7521);
and U13483 (N_13483,N_7118,N_9825);
nor U13484 (N_13484,N_7647,N_5719);
nor U13485 (N_13485,N_9956,N_9294);
and U13486 (N_13486,N_6682,N_7292);
nor U13487 (N_13487,N_6211,N_5579);
and U13488 (N_13488,N_8413,N_8221);
nand U13489 (N_13489,N_8391,N_9130);
or U13490 (N_13490,N_8059,N_8829);
or U13491 (N_13491,N_6692,N_7407);
nor U13492 (N_13492,N_5614,N_8029);
xor U13493 (N_13493,N_8956,N_6653);
nand U13494 (N_13494,N_7193,N_8944);
xnor U13495 (N_13495,N_9753,N_5514);
and U13496 (N_13496,N_7871,N_6129);
nor U13497 (N_13497,N_9733,N_6074);
nand U13498 (N_13498,N_9483,N_9425);
nor U13499 (N_13499,N_8451,N_7742);
xnor U13500 (N_13500,N_8819,N_9040);
or U13501 (N_13501,N_5068,N_5198);
or U13502 (N_13502,N_7777,N_8254);
nor U13503 (N_13503,N_9483,N_9780);
nand U13504 (N_13504,N_8652,N_5234);
and U13505 (N_13505,N_5593,N_5755);
and U13506 (N_13506,N_8096,N_6836);
nor U13507 (N_13507,N_5235,N_9059);
or U13508 (N_13508,N_7190,N_5261);
nor U13509 (N_13509,N_6171,N_7609);
nor U13510 (N_13510,N_7688,N_6448);
xnor U13511 (N_13511,N_9337,N_7960);
xnor U13512 (N_13512,N_6795,N_8436);
xnor U13513 (N_13513,N_8250,N_9480);
nor U13514 (N_13514,N_5948,N_5532);
and U13515 (N_13515,N_7131,N_6652);
or U13516 (N_13516,N_8869,N_8160);
nor U13517 (N_13517,N_7491,N_7772);
nor U13518 (N_13518,N_8441,N_5651);
nor U13519 (N_13519,N_6018,N_9365);
and U13520 (N_13520,N_8204,N_5650);
or U13521 (N_13521,N_7880,N_7745);
nand U13522 (N_13522,N_7136,N_8151);
and U13523 (N_13523,N_5832,N_8754);
nor U13524 (N_13524,N_7663,N_5977);
nand U13525 (N_13525,N_7756,N_8893);
nand U13526 (N_13526,N_5784,N_6666);
or U13527 (N_13527,N_9980,N_5145);
xor U13528 (N_13528,N_6705,N_8332);
or U13529 (N_13529,N_8205,N_7242);
and U13530 (N_13530,N_8583,N_5591);
or U13531 (N_13531,N_8640,N_8604);
xnor U13532 (N_13532,N_8807,N_8539);
xnor U13533 (N_13533,N_9369,N_5669);
xor U13534 (N_13534,N_5172,N_5058);
nand U13535 (N_13535,N_9333,N_7337);
xnor U13536 (N_13536,N_9998,N_9572);
nand U13537 (N_13537,N_5903,N_9923);
nand U13538 (N_13538,N_6448,N_7135);
xnor U13539 (N_13539,N_5883,N_9956);
xnor U13540 (N_13540,N_8152,N_7973);
or U13541 (N_13541,N_8274,N_7327);
xor U13542 (N_13542,N_7460,N_8015);
xnor U13543 (N_13543,N_9836,N_9111);
nand U13544 (N_13544,N_8858,N_5604);
and U13545 (N_13545,N_5087,N_5330);
and U13546 (N_13546,N_9851,N_7832);
xnor U13547 (N_13547,N_9637,N_7623);
nor U13548 (N_13548,N_7452,N_7486);
and U13549 (N_13549,N_6719,N_9769);
nand U13550 (N_13550,N_9419,N_9061);
or U13551 (N_13551,N_8828,N_8386);
and U13552 (N_13552,N_8174,N_7161);
or U13553 (N_13553,N_9988,N_7342);
nor U13554 (N_13554,N_5658,N_6243);
nand U13555 (N_13555,N_7472,N_7764);
nor U13556 (N_13556,N_9721,N_9716);
or U13557 (N_13557,N_6700,N_5211);
xnor U13558 (N_13558,N_7552,N_9495);
xnor U13559 (N_13559,N_5616,N_7184);
nand U13560 (N_13560,N_7208,N_7192);
or U13561 (N_13561,N_9194,N_9602);
nand U13562 (N_13562,N_6562,N_6736);
or U13563 (N_13563,N_5330,N_9673);
nand U13564 (N_13564,N_7672,N_6439);
nor U13565 (N_13565,N_6078,N_6163);
nand U13566 (N_13566,N_8731,N_9150);
xor U13567 (N_13567,N_9370,N_7181);
or U13568 (N_13568,N_5182,N_5716);
xor U13569 (N_13569,N_6768,N_8926);
or U13570 (N_13570,N_7511,N_9459);
nand U13571 (N_13571,N_8909,N_7813);
and U13572 (N_13572,N_9398,N_5650);
nand U13573 (N_13573,N_6974,N_9755);
and U13574 (N_13574,N_5707,N_9475);
nor U13575 (N_13575,N_6585,N_6576);
nor U13576 (N_13576,N_8868,N_9195);
and U13577 (N_13577,N_6205,N_8021);
and U13578 (N_13578,N_8749,N_6399);
nor U13579 (N_13579,N_9177,N_6495);
xor U13580 (N_13580,N_8827,N_8618);
and U13581 (N_13581,N_5299,N_9664);
and U13582 (N_13582,N_7894,N_5641);
and U13583 (N_13583,N_9135,N_9462);
nor U13584 (N_13584,N_5134,N_8557);
nor U13585 (N_13585,N_8009,N_8303);
or U13586 (N_13586,N_8983,N_6782);
xnor U13587 (N_13587,N_9380,N_5060);
xor U13588 (N_13588,N_7960,N_8957);
and U13589 (N_13589,N_8436,N_7483);
or U13590 (N_13590,N_8190,N_6608);
and U13591 (N_13591,N_9425,N_7662);
nor U13592 (N_13592,N_5367,N_6415);
nand U13593 (N_13593,N_6963,N_6031);
xor U13594 (N_13594,N_6035,N_7752);
nor U13595 (N_13595,N_9274,N_7223);
or U13596 (N_13596,N_9918,N_6755);
xnor U13597 (N_13597,N_6145,N_6088);
and U13598 (N_13598,N_6459,N_8564);
or U13599 (N_13599,N_7584,N_9220);
and U13600 (N_13600,N_7973,N_9702);
xnor U13601 (N_13601,N_6635,N_5265);
nor U13602 (N_13602,N_6842,N_8303);
nand U13603 (N_13603,N_5340,N_7414);
and U13604 (N_13604,N_8952,N_7954);
and U13605 (N_13605,N_6012,N_9813);
and U13606 (N_13606,N_5021,N_5405);
xnor U13607 (N_13607,N_7993,N_6863);
nor U13608 (N_13608,N_7862,N_8645);
xnor U13609 (N_13609,N_9371,N_9876);
nor U13610 (N_13610,N_5952,N_9320);
xor U13611 (N_13611,N_7779,N_9104);
nor U13612 (N_13612,N_9970,N_6997);
nand U13613 (N_13613,N_5880,N_6580);
or U13614 (N_13614,N_7199,N_6760);
nor U13615 (N_13615,N_6501,N_8716);
or U13616 (N_13616,N_9931,N_8211);
xor U13617 (N_13617,N_9080,N_5661);
nor U13618 (N_13618,N_6823,N_6602);
or U13619 (N_13619,N_9057,N_6726);
or U13620 (N_13620,N_7956,N_5619);
xor U13621 (N_13621,N_8807,N_8055);
nand U13622 (N_13622,N_9843,N_9421);
nand U13623 (N_13623,N_6561,N_8912);
nor U13624 (N_13624,N_8311,N_5688);
or U13625 (N_13625,N_7000,N_8378);
or U13626 (N_13626,N_5518,N_7147);
nand U13627 (N_13627,N_5357,N_7292);
or U13628 (N_13628,N_7931,N_8589);
nand U13629 (N_13629,N_6845,N_6811);
or U13630 (N_13630,N_9459,N_6646);
xor U13631 (N_13631,N_6262,N_6842);
nor U13632 (N_13632,N_5602,N_7374);
or U13633 (N_13633,N_8795,N_8312);
nand U13634 (N_13634,N_6737,N_9361);
xnor U13635 (N_13635,N_7588,N_7424);
and U13636 (N_13636,N_9475,N_7133);
nor U13637 (N_13637,N_9245,N_6611);
nand U13638 (N_13638,N_7962,N_5750);
or U13639 (N_13639,N_5887,N_6742);
nand U13640 (N_13640,N_8120,N_6030);
and U13641 (N_13641,N_8639,N_9724);
nand U13642 (N_13642,N_5393,N_6719);
xor U13643 (N_13643,N_9215,N_7592);
nand U13644 (N_13644,N_7483,N_9046);
and U13645 (N_13645,N_6830,N_9424);
and U13646 (N_13646,N_9719,N_9513);
and U13647 (N_13647,N_9406,N_6689);
xor U13648 (N_13648,N_7078,N_6798);
nor U13649 (N_13649,N_7732,N_8573);
nor U13650 (N_13650,N_7475,N_6902);
xnor U13651 (N_13651,N_7423,N_8316);
or U13652 (N_13652,N_8786,N_6930);
xor U13653 (N_13653,N_6623,N_8234);
nor U13654 (N_13654,N_9638,N_9971);
nand U13655 (N_13655,N_5835,N_8640);
xor U13656 (N_13656,N_5754,N_6334);
or U13657 (N_13657,N_6587,N_7997);
or U13658 (N_13658,N_7476,N_9106);
nor U13659 (N_13659,N_8006,N_9592);
nor U13660 (N_13660,N_9538,N_6783);
and U13661 (N_13661,N_8913,N_9110);
nor U13662 (N_13662,N_7719,N_5395);
or U13663 (N_13663,N_5718,N_7763);
or U13664 (N_13664,N_6301,N_5300);
nor U13665 (N_13665,N_8386,N_7445);
nand U13666 (N_13666,N_6295,N_7486);
nand U13667 (N_13667,N_9167,N_7526);
nand U13668 (N_13668,N_9749,N_8116);
and U13669 (N_13669,N_8415,N_9572);
nand U13670 (N_13670,N_9024,N_9640);
or U13671 (N_13671,N_5054,N_7005);
nor U13672 (N_13672,N_8726,N_7981);
and U13673 (N_13673,N_9399,N_7238);
nand U13674 (N_13674,N_5755,N_8412);
xnor U13675 (N_13675,N_8539,N_8406);
nor U13676 (N_13676,N_9946,N_5482);
nor U13677 (N_13677,N_9953,N_8137);
nor U13678 (N_13678,N_9840,N_7179);
nor U13679 (N_13679,N_7732,N_9522);
nor U13680 (N_13680,N_6147,N_9300);
nor U13681 (N_13681,N_9274,N_5289);
nor U13682 (N_13682,N_7479,N_6286);
or U13683 (N_13683,N_5004,N_5005);
nand U13684 (N_13684,N_8998,N_6372);
xnor U13685 (N_13685,N_9497,N_8613);
and U13686 (N_13686,N_5270,N_5547);
or U13687 (N_13687,N_8694,N_5203);
or U13688 (N_13688,N_9696,N_5363);
xor U13689 (N_13689,N_9233,N_7156);
nor U13690 (N_13690,N_8865,N_7586);
or U13691 (N_13691,N_8918,N_6505);
and U13692 (N_13692,N_5673,N_5609);
or U13693 (N_13693,N_6644,N_6216);
nor U13694 (N_13694,N_9817,N_9721);
nor U13695 (N_13695,N_9654,N_5011);
or U13696 (N_13696,N_5493,N_5050);
nor U13697 (N_13697,N_7581,N_6945);
xor U13698 (N_13698,N_5388,N_9032);
nor U13699 (N_13699,N_7388,N_8728);
xor U13700 (N_13700,N_5974,N_6244);
xor U13701 (N_13701,N_7696,N_7188);
xnor U13702 (N_13702,N_9934,N_7662);
and U13703 (N_13703,N_8753,N_8752);
nand U13704 (N_13704,N_6747,N_8778);
nor U13705 (N_13705,N_7829,N_8227);
xnor U13706 (N_13706,N_7383,N_6047);
xor U13707 (N_13707,N_9296,N_7159);
xor U13708 (N_13708,N_5596,N_6846);
or U13709 (N_13709,N_6290,N_6288);
nand U13710 (N_13710,N_9952,N_9984);
or U13711 (N_13711,N_7901,N_6971);
nor U13712 (N_13712,N_9043,N_7889);
or U13713 (N_13713,N_9056,N_7970);
nand U13714 (N_13714,N_9286,N_9993);
xor U13715 (N_13715,N_7221,N_9478);
and U13716 (N_13716,N_6139,N_5601);
nor U13717 (N_13717,N_8752,N_7406);
or U13718 (N_13718,N_6783,N_8695);
nor U13719 (N_13719,N_7605,N_9949);
xnor U13720 (N_13720,N_6036,N_6558);
nor U13721 (N_13721,N_8450,N_7379);
nand U13722 (N_13722,N_9495,N_5886);
xnor U13723 (N_13723,N_7587,N_6438);
xnor U13724 (N_13724,N_5036,N_5882);
and U13725 (N_13725,N_6348,N_6786);
and U13726 (N_13726,N_9233,N_7672);
and U13727 (N_13727,N_7557,N_8576);
or U13728 (N_13728,N_8852,N_9354);
or U13729 (N_13729,N_7661,N_8370);
nor U13730 (N_13730,N_8157,N_8832);
nand U13731 (N_13731,N_8914,N_5508);
nor U13732 (N_13732,N_8379,N_7093);
nor U13733 (N_13733,N_5341,N_6037);
nor U13734 (N_13734,N_6972,N_6327);
xnor U13735 (N_13735,N_5875,N_9920);
or U13736 (N_13736,N_6809,N_9202);
xnor U13737 (N_13737,N_5221,N_6371);
and U13738 (N_13738,N_6919,N_8305);
or U13739 (N_13739,N_6811,N_5336);
nand U13740 (N_13740,N_5189,N_6328);
nor U13741 (N_13741,N_9802,N_9425);
or U13742 (N_13742,N_9909,N_8543);
and U13743 (N_13743,N_6041,N_8312);
nor U13744 (N_13744,N_5712,N_5110);
and U13745 (N_13745,N_7237,N_7702);
nand U13746 (N_13746,N_9843,N_8293);
or U13747 (N_13747,N_5805,N_9869);
nor U13748 (N_13748,N_5168,N_9105);
or U13749 (N_13749,N_8587,N_7042);
nor U13750 (N_13750,N_9338,N_7955);
xnor U13751 (N_13751,N_7657,N_5959);
nor U13752 (N_13752,N_8039,N_8755);
xnor U13753 (N_13753,N_5955,N_7945);
nor U13754 (N_13754,N_9506,N_6924);
nand U13755 (N_13755,N_7629,N_9413);
nand U13756 (N_13756,N_6156,N_7758);
xnor U13757 (N_13757,N_8476,N_7291);
or U13758 (N_13758,N_7920,N_9028);
nor U13759 (N_13759,N_7373,N_9130);
nor U13760 (N_13760,N_6968,N_8592);
xnor U13761 (N_13761,N_6116,N_8626);
nor U13762 (N_13762,N_7532,N_8912);
and U13763 (N_13763,N_8547,N_7890);
nor U13764 (N_13764,N_9623,N_7431);
or U13765 (N_13765,N_6144,N_6172);
nor U13766 (N_13766,N_9711,N_7119);
xor U13767 (N_13767,N_6545,N_8495);
xor U13768 (N_13768,N_5538,N_8178);
and U13769 (N_13769,N_5002,N_7973);
and U13770 (N_13770,N_9834,N_7698);
and U13771 (N_13771,N_7380,N_6493);
or U13772 (N_13772,N_8784,N_9105);
and U13773 (N_13773,N_5553,N_7879);
nor U13774 (N_13774,N_6171,N_8664);
nor U13775 (N_13775,N_8886,N_9821);
nor U13776 (N_13776,N_7666,N_5090);
nor U13777 (N_13777,N_9997,N_8883);
nand U13778 (N_13778,N_5477,N_8509);
or U13779 (N_13779,N_9404,N_7218);
nand U13780 (N_13780,N_5410,N_8991);
xor U13781 (N_13781,N_8395,N_6503);
and U13782 (N_13782,N_5556,N_8485);
nand U13783 (N_13783,N_7044,N_5745);
xor U13784 (N_13784,N_7225,N_7519);
xor U13785 (N_13785,N_7478,N_9753);
and U13786 (N_13786,N_5694,N_5581);
nand U13787 (N_13787,N_5984,N_6325);
and U13788 (N_13788,N_7124,N_6884);
nand U13789 (N_13789,N_5518,N_5281);
xor U13790 (N_13790,N_5108,N_5210);
or U13791 (N_13791,N_6657,N_7263);
and U13792 (N_13792,N_5889,N_8372);
nor U13793 (N_13793,N_5341,N_7868);
nor U13794 (N_13794,N_6271,N_6739);
nor U13795 (N_13795,N_7140,N_5713);
nand U13796 (N_13796,N_5080,N_6248);
nor U13797 (N_13797,N_9967,N_5221);
xor U13798 (N_13798,N_7761,N_6426);
and U13799 (N_13799,N_6417,N_8316);
and U13800 (N_13800,N_7947,N_5550);
and U13801 (N_13801,N_8546,N_7247);
nand U13802 (N_13802,N_9735,N_9537);
xnor U13803 (N_13803,N_8518,N_6772);
xor U13804 (N_13804,N_5544,N_6233);
and U13805 (N_13805,N_8744,N_7487);
or U13806 (N_13806,N_8365,N_6368);
nor U13807 (N_13807,N_7991,N_8290);
and U13808 (N_13808,N_6037,N_8365);
or U13809 (N_13809,N_6304,N_5621);
and U13810 (N_13810,N_7345,N_8626);
nor U13811 (N_13811,N_9241,N_8860);
or U13812 (N_13812,N_6720,N_9210);
and U13813 (N_13813,N_5338,N_7182);
xor U13814 (N_13814,N_5717,N_5974);
xnor U13815 (N_13815,N_6565,N_6055);
xnor U13816 (N_13816,N_9121,N_6328);
xor U13817 (N_13817,N_8336,N_5720);
nor U13818 (N_13818,N_8563,N_5226);
nand U13819 (N_13819,N_7196,N_6287);
nand U13820 (N_13820,N_7108,N_6521);
nor U13821 (N_13821,N_6294,N_7943);
nor U13822 (N_13822,N_9176,N_9161);
nand U13823 (N_13823,N_7722,N_6272);
or U13824 (N_13824,N_7160,N_5242);
nor U13825 (N_13825,N_8717,N_8619);
xnor U13826 (N_13826,N_6247,N_5794);
and U13827 (N_13827,N_6683,N_7234);
xnor U13828 (N_13828,N_9313,N_9974);
xor U13829 (N_13829,N_7794,N_9725);
or U13830 (N_13830,N_7910,N_9387);
nor U13831 (N_13831,N_7462,N_5746);
or U13832 (N_13832,N_8876,N_5787);
or U13833 (N_13833,N_9132,N_8608);
or U13834 (N_13834,N_7315,N_9014);
nor U13835 (N_13835,N_8447,N_9235);
xnor U13836 (N_13836,N_5865,N_9713);
or U13837 (N_13837,N_6373,N_6219);
and U13838 (N_13838,N_5299,N_9057);
or U13839 (N_13839,N_9414,N_8492);
and U13840 (N_13840,N_9752,N_8622);
and U13841 (N_13841,N_9069,N_9131);
or U13842 (N_13842,N_5187,N_7465);
nand U13843 (N_13843,N_9012,N_5821);
xor U13844 (N_13844,N_6374,N_6555);
nand U13845 (N_13845,N_8292,N_5367);
nand U13846 (N_13846,N_9497,N_8950);
nand U13847 (N_13847,N_5551,N_5374);
nor U13848 (N_13848,N_6391,N_9048);
nor U13849 (N_13849,N_9906,N_8832);
nor U13850 (N_13850,N_7185,N_5319);
nor U13851 (N_13851,N_7052,N_7078);
or U13852 (N_13852,N_5304,N_8229);
nor U13853 (N_13853,N_6867,N_5416);
and U13854 (N_13854,N_5360,N_9838);
and U13855 (N_13855,N_7604,N_6879);
nand U13856 (N_13856,N_6343,N_9531);
xor U13857 (N_13857,N_8978,N_5788);
or U13858 (N_13858,N_9143,N_7860);
and U13859 (N_13859,N_8948,N_8831);
nor U13860 (N_13860,N_8142,N_8145);
and U13861 (N_13861,N_7140,N_9965);
and U13862 (N_13862,N_7356,N_6407);
and U13863 (N_13863,N_6719,N_8075);
nor U13864 (N_13864,N_5237,N_5432);
nor U13865 (N_13865,N_5275,N_5042);
or U13866 (N_13866,N_9585,N_7041);
and U13867 (N_13867,N_8735,N_8772);
nor U13868 (N_13868,N_5051,N_7644);
or U13869 (N_13869,N_6938,N_8049);
and U13870 (N_13870,N_6895,N_5401);
nor U13871 (N_13871,N_7685,N_9084);
nor U13872 (N_13872,N_9140,N_7764);
nor U13873 (N_13873,N_7327,N_9247);
or U13874 (N_13874,N_9461,N_6704);
nor U13875 (N_13875,N_8208,N_5162);
and U13876 (N_13876,N_6137,N_7508);
or U13877 (N_13877,N_7363,N_9924);
xor U13878 (N_13878,N_8608,N_9111);
or U13879 (N_13879,N_7307,N_9260);
xor U13880 (N_13880,N_9763,N_9012);
and U13881 (N_13881,N_7986,N_6198);
nand U13882 (N_13882,N_9139,N_7538);
nor U13883 (N_13883,N_7443,N_6374);
nor U13884 (N_13884,N_9406,N_5455);
and U13885 (N_13885,N_7866,N_7155);
and U13886 (N_13886,N_5904,N_8231);
nand U13887 (N_13887,N_7509,N_6232);
xnor U13888 (N_13888,N_8008,N_7770);
xor U13889 (N_13889,N_5793,N_8150);
nor U13890 (N_13890,N_7573,N_7204);
or U13891 (N_13891,N_5043,N_8392);
or U13892 (N_13892,N_7215,N_9912);
nor U13893 (N_13893,N_8095,N_7202);
and U13894 (N_13894,N_6378,N_5794);
nor U13895 (N_13895,N_6284,N_5091);
xor U13896 (N_13896,N_6311,N_5903);
nand U13897 (N_13897,N_5650,N_9797);
and U13898 (N_13898,N_9454,N_9293);
nand U13899 (N_13899,N_6499,N_9540);
nor U13900 (N_13900,N_6841,N_8463);
or U13901 (N_13901,N_9122,N_6345);
or U13902 (N_13902,N_8431,N_8899);
nor U13903 (N_13903,N_7039,N_8707);
nand U13904 (N_13904,N_6674,N_5404);
nand U13905 (N_13905,N_8221,N_6259);
xor U13906 (N_13906,N_9111,N_6021);
and U13907 (N_13907,N_7045,N_5560);
or U13908 (N_13908,N_8839,N_7405);
and U13909 (N_13909,N_7238,N_6539);
nor U13910 (N_13910,N_8915,N_9273);
nor U13911 (N_13911,N_8351,N_8401);
xnor U13912 (N_13912,N_8327,N_9580);
and U13913 (N_13913,N_5324,N_8736);
nor U13914 (N_13914,N_8952,N_9798);
and U13915 (N_13915,N_8961,N_9868);
and U13916 (N_13916,N_8470,N_9791);
nand U13917 (N_13917,N_9914,N_9864);
nor U13918 (N_13918,N_7061,N_9855);
or U13919 (N_13919,N_6299,N_5655);
and U13920 (N_13920,N_7423,N_6429);
or U13921 (N_13921,N_9548,N_8270);
nand U13922 (N_13922,N_9598,N_6131);
nand U13923 (N_13923,N_5199,N_9196);
or U13924 (N_13924,N_8837,N_6818);
nor U13925 (N_13925,N_8555,N_6004);
nor U13926 (N_13926,N_6430,N_6800);
and U13927 (N_13927,N_7432,N_8811);
and U13928 (N_13928,N_9874,N_8610);
xnor U13929 (N_13929,N_5729,N_9791);
or U13930 (N_13930,N_7675,N_7834);
xnor U13931 (N_13931,N_6771,N_6357);
xor U13932 (N_13932,N_8385,N_7666);
nand U13933 (N_13933,N_6847,N_9854);
or U13934 (N_13934,N_9327,N_8053);
xnor U13935 (N_13935,N_7729,N_6055);
nor U13936 (N_13936,N_9123,N_6346);
nand U13937 (N_13937,N_6172,N_5273);
and U13938 (N_13938,N_9334,N_9463);
or U13939 (N_13939,N_6962,N_6438);
nor U13940 (N_13940,N_7920,N_6667);
or U13941 (N_13941,N_9791,N_9149);
xnor U13942 (N_13942,N_8014,N_5460);
xor U13943 (N_13943,N_8657,N_5989);
nor U13944 (N_13944,N_6810,N_6129);
or U13945 (N_13945,N_5323,N_7875);
and U13946 (N_13946,N_6475,N_6081);
nand U13947 (N_13947,N_5111,N_9176);
nand U13948 (N_13948,N_5437,N_5246);
xnor U13949 (N_13949,N_6618,N_5839);
or U13950 (N_13950,N_6999,N_8029);
xor U13951 (N_13951,N_5489,N_8675);
nand U13952 (N_13952,N_9170,N_5606);
nand U13953 (N_13953,N_6476,N_6042);
xnor U13954 (N_13954,N_5870,N_8146);
xnor U13955 (N_13955,N_8627,N_7766);
and U13956 (N_13956,N_8589,N_8561);
and U13957 (N_13957,N_5586,N_9752);
or U13958 (N_13958,N_9337,N_9528);
nor U13959 (N_13959,N_9779,N_7498);
or U13960 (N_13960,N_6466,N_9923);
nor U13961 (N_13961,N_5453,N_9287);
nand U13962 (N_13962,N_5291,N_8490);
and U13963 (N_13963,N_6626,N_5715);
nor U13964 (N_13964,N_8470,N_6768);
xnor U13965 (N_13965,N_9244,N_7442);
nor U13966 (N_13966,N_8563,N_9723);
nand U13967 (N_13967,N_5267,N_8388);
nand U13968 (N_13968,N_8713,N_6718);
or U13969 (N_13969,N_7364,N_9348);
nand U13970 (N_13970,N_7941,N_9989);
and U13971 (N_13971,N_9290,N_9518);
nand U13972 (N_13972,N_8014,N_6329);
nor U13973 (N_13973,N_8571,N_9633);
and U13974 (N_13974,N_8612,N_8197);
or U13975 (N_13975,N_9072,N_7072);
xor U13976 (N_13976,N_9456,N_6342);
xnor U13977 (N_13977,N_8529,N_5096);
nor U13978 (N_13978,N_7196,N_9994);
nand U13979 (N_13979,N_5018,N_7523);
nand U13980 (N_13980,N_5250,N_7013);
nand U13981 (N_13981,N_6921,N_8478);
nor U13982 (N_13982,N_8348,N_9198);
and U13983 (N_13983,N_6739,N_5894);
and U13984 (N_13984,N_5899,N_5204);
nand U13985 (N_13985,N_6582,N_8492);
nor U13986 (N_13986,N_7512,N_5638);
nand U13987 (N_13987,N_5264,N_7320);
xor U13988 (N_13988,N_8954,N_9098);
nor U13989 (N_13989,N_6046,N_7983);
and U13990 (N_13990,N_7622,N_8697);
and U13991 (N_13991,N_8053,N_8809);
nand U13992 (N_13992,N_5374,N_8644);
nand U13993 (N_13993,N_5208,N_8556);
and U13994 (N_13994,N_8207,N_6528);
nand U13995 (N_13995,N_7221,N_6470);
nand U13996 (N_13996,N_5995,N_8696);
xnor U13997 (N_13997,N_8829,N_5851);
nand U13998 (N_13998,N_5569,N_9404);
nor U13999 (N_13999,N_9636,N_6968);
or U14000 (N_14000,N_5074,N_7860);
xnor U14001 (N_14001,N_7604,N_6710);
nor U14002 (N_14002,N_8765,N_9895);
xor U14003 (N_14003,N_8223,N_5982);
or U14004 (N_14004,N_7375,N_6637);
and U14005 (N_14005,N_7576,N_8982);
and U14006 (N_14006,N_5296,N_5451);
nor U14007 (N_14007,N_5888,N_8659);
xor U14008 (N_14008,N_5789,N_7728);
nor U14009 (N_14009,N_8303,N_7307);
nand U14010 (N_14010,N_7871,N_5235);
xor U14011 (N_14011,N_7701,N_5310);
nand U14012 (N_14012,N_6593,N_9787);
and U14013 (N_14013,N_6385,N_7114);
or U14014 (N_14014,N_5758,N_8063);
and U14015 (N_14015,N_5036,N_8762);
nor U14016 (N_14016,N_7368,N_8862);
nor U14017 (N_14017,N_5348,N_7524);
and U14018 (N_14018,N_8780,N_7751);
nand U14019 (N_14019,N_6762,N_9110);
nand U14020 (N_14020,N_6429,N_7101);
xnor U14021 (N_14021,N_9581,N_9173);
or U14022 (N_14022,N_6912,N_8156);
nor U14023 (N_14023,N_9887,N_7116);
xor U14024 (N_14024,N_5322,N_5757);
and U14025 (N_14025,N_5228,N_7980);
or U14026 (N_14026,N_5434,N_8385);
or U14027 (N_14027,N_5380,N_6188);
nand U14028 (N_14028,N_5114,N_6519);
nor U14029 (N_14029,N_7060,N_6015);
nand U14030 (N_14030,N_5093,N_7577);
nor U14031 (N_14031,N_9387,N_9390);
and U14032 (N_14032,N_5940,N_9346);
xor U14033 (N_14033,N_9898,N_7572);
nand U14034 (N_14034,N_6808,N_7657);
or U14035 (N_14035,N_9938,N_5868);
xor U14036 (N_14036,N_5796,N_9704);
and U14037 (N_14037,N_8010,N_5060);
nand U14038 (N_14038,N_8597,N_6793);
xor U14039 (N_14039,N_9034,N_9614);
xor U14040 (N_14040,N_9198,N_8362);
nor U14041 (N_14041,N_9996,N_8237);
nor U14042 (N_14042,N_6299,N_9409);
or U14043 (N_14043,N_6825,N_7927);
or U14044 (N_14044,N_9531,N_6341);
nor U14045 (N_14045,N_5686,N_6075);
xor U14046 (N_14046,N_6015,N_6800);
nor U14047 (N_14047,N_5030,N_8166);
nor U14048 (N_14048,N_5224,N_9006);
nor U14049 (N_14049,N_5504,N_5716);
or U14050 (N_14050,N_7580,N_7366);
and U14051 (N_14051,N_6182,N_5972);
nand U14052 (N_14052,N_6554,N_5979);
nor U14053 (N_14053,N_8137,N_5259);
nand U14054 (N_14054,N_9130,N_9207);
xnor U14055 (N_14055,N_9424,N_8492);
or U14056 (N_14056,N_6785,N_8939);
or U14057 (N_14057,N_8722,N_5676);
or U14058 (N_14058,N_9609,N_6111);
or U14059 (N_14059,N_5989,N_8589);
nand U14060 (N_14060,N_9348,N_8828);
xnor U14061 (N_14061,N_8068,N_7358);
or U14062 (N_14062,N_5888,N_9577);
or U14063 (N_14063,N_8372,N_7531);
nor U14064 (N_14064,N_9814,N_6531);
or U14065 (N_14065,N_6496,N_7257);
nand U14066 (N_14066,N_7256,N_7503);
xor U14067 (N_14067,N_5083,N_7543);
or U14068 (N_14068,N_7896,N_5310);
or U14069 (N_14069,N_9710,N_6154);
and U14070 (N_14070,N_6032,N_5659);
nand U14071 (N_14071,N_9841,N_9660);
nor U14072 (N_14072,N_5861,N_6641);
and U14073 (N_14073,N_8570,N_5222);
or U14074 (N_14074,N_9758,N_6707);
and U14075 (N_14075,N_6851,N_6548);
nand U14076 (N_14076,N_8271,N_6607);
or U14077 (N_14077,N_7912,N_7042);
xnor U14078 (N_14078,N_9819,N_9808);
and U14079 (N_14079,N_6316,N_5006);
xor U14080 (N_14080,N_9380,N_6139);
or U14081 (N_14081,N_8994,N_9233);
nor U14082 (N_14082,N_6206,N_7637);
and U14083 (N_14083,N_7301,N_5150);
xor U14084 (N_14084,N_6922,N_5680);
nand U14085 (N_14085,N_7576,N_9774);
xor U14086 (N_14086,N_6304,N_6198);
or U14087 (N_14087,N_9358,N_7598);
nor U14088 (N_14088,N_6406,N_8698);
and U14089 (N_14089,N_7562,N_9754);
and U14090 (N_14090,N_7141,N_9812);
xnor U14091 (N_14091,N_8292,N_5894);
and U14092 (N_14092,N_8440,N_8095);
or U14093 (N_14093,N_9151,N_9604);
or U14094 (N_14094,N_8670,N_7280);
or U14095 (N_14095,N_9189,N_5743);
and U14096 (N_14096,N_9762,N_7741);
or U14097 (N_14097,N_5005,N_8700);
xnor U14098 (N_14098,N_8840,N_8907);
nand U14099 (N_14099,N_6457,N_8383);
or U14100 (N_14100,N_9322,N_7325);
nor U14101 (N_14101,N_8924,N_5074);
nor U14102 (N_14102,N_5173,N_9179);
nor U14103 (N_14103,N_9116,N_8490);
or U14104 (N_14104,N_7224,N_7094);
or U14105 (N_14105,N_9797,N_8729);
or U14106 (N_14106,N_5989,N_6449);
xor U14107 (N_14107,N_9542,N_5319);
or U14108 (N_14108,N_7137,N_8542);
or U14109 (N_14109,N_5474,N_9016);
and U14110 (N_14110,N_7006,N_8359);
or U14111 (N_14111,N_7941,N_9604);
nor U14112 (N_14112,N_5273,N_6685);
nand U14113 (N_14113,N_7724,N_8338);
and U14114 (N_14114,N_5832,N_5125);
nand U14115 (N_14115,N_6541,N_5531);
nand U14116 (N_14116,N_7851,N_5892);
and U14117 (N_14117,N_7654,N_9864);
or U14118 (N_14118,N_9319,N_6965);
or U14119 (N_14119,N_7341,N_6640);
or U14120 (N_14120,N_8722,N_8993);
xnor U14121 (N_14121,N_6049,N_6223);
or U14122 (N_14122,N_9596,N_6296);
nand U14123 (N_14123,N_5494,N_6593);
nand U14124 (N_14124,N_7093,N_8664);
nor U14125 (N_14125,N_8265,N_5373);
and U14126 (N_14126,N_9063,N_9477);
xor U14127 (N_14127,N_8880,N_5953);
xor U14128 (N_14128,N_6253,N_7540);
and U14129 (N_14129,N_7716,N_9885);
or U14130 (N_14130,N_8106,N_5554);
nand U14131 (N_14131,N_9938,N_9986);
nor U14132 (N_14132,N_7885,N_9032);
and U14133 (N_14133,N_7693,N_8329);
and U14134 (N_14134,N_6095,N_5292);
xor U14135 (N_14135,N_9507,N_5532);
xnor U14136 (N_14136,N_7732,N_8802);
or U14137 (N_14137,N_6600,N_6376);
and U14138 (N_14138,N_8386,N_6721);
and U14139 (N_14139,N_5281,N_9431);
nor U14140 (N_14140,N_8396,N_5833);
or U14141 (N_14141,N_6352,N_9171);
or U14142 (N_14142,N_8326,N_5430);
nand U14143 (N_14143,N_6197,N_8218);
xor U14144 (N_14144,N_8230,N_9906);
nor U14145 (N_14145,N_7884,N_9833);
nand U14146 (N_14146,N_9084,N_7622);
and U14147 (N_14147,N_7578,N_7918);
nor U14148 (N_14148,N_6049,N_5960);
xnor U14149 (N_14149,N_5116,N_7503);
nand U14150 (N_14150,N_5533,N_9919);
or U14151 (N_14151,N_6213,N_9235);
or U14152 (N_14152,N_8461,N_6445);
and U14153 (N_14153,N_6300,N_7909);
or U14154 (N_14154,N_7276,N_9701);
nor U14155 (N_14155,N_9872,N_8567);
nand U14156 (N_14156,N_7361,N_7132);
nor U14157 (N_14157,N_5966,N_5350);
nand U14158 (N_14158,N_6826,N_7821);
xnor U14159 (N_14159,N_9482,N_5793);
and U14160 (N_14160,N_8559,N_6981);
nand U14161 (N_14161,N_9475,N_8657);
xor U14162 (N_14162,N_8321,N_9849);
and U14163 (N_14163,N_9328,N_5522);
and U14164 (N_14164,N_5844,N_7514);
xor U14165 (N_14165,N_5412,N_7592);
and U14166 (N_14166,N_7719,N_5814);
nor U14167 (N_14167,N_8230,N_6384);
or U14168 (N_14168,N_9982,N_7750);
nand U14169 (N_14169,N_8134,N_6106);
or U14170 (N_14170,N_9385,N_7779);
nor U14171 (N_14171,N_9659,N_9581);
nand U14172 (N_14172,N_8154,N_9304);
xor U14173 (N_14173,N_9520,N_7929);
and U14174 (N_14174,N_9061,N_7942);
nand U14175 (N_14175,N_6832,N_9182);
or U14176 (N_14176,N_9202,N_9430);
nor U14177 (N_14177,N_8036,N_9271);
nor U14178 (N_14178,N_9030,N_8034);
xnor U14179 (N_14179,N_7053,N_6938);
nand U14180 (N_14180,N_9660,N_5985);
nor U14181 (N_14181,N_6999,N_8764);
xnor U14182 (N_14182,N_6994,N_7804);
xor U14183 (N_14183,N_5735,N_9614);
and U14184 (N_14184,N_5064,N_5173);
nor U14185 (N_14185,N_8774,N_7916);
nand U14186 (N_14186,N_8061,N_7430);
xnor U14187 (N_14187,N_9769,N_9852);
xor U14188 (N_14188,N_9536,N_9500);
or U14189 (N_14189,N_6030,N_7848);
xor U14190 (N_14190,N_9050,N_6898);
xnor U14191 (N_14191,N_8542,N_6439);
nand U14192 (N_14192,N_8140,N_9989);
and U14193 (N_14193,N_6326,N_6394);
or U14194 (N_14194,N_6324,N_5371);
xnor U14195 (N_14195,N_8261,N_8853);
or U14196 (N_14196,N_6847,N_7501);
xnor U14197 (N_14197,N_9535,N_6772);
nand U14198 (N_14198,N_8216,N_8633);
or U14199 (N_14199,N_9222,N_5403);
xnor U14200 (N_14200,N_5555,N_9894);
xnor U14201 (N_14201,N_5951,N_9102);
nor U14202 (N_14202,N_8789,N_6901);
nor U14203 (N_14203,N_7650,N_9313);
and U14204 (N_14204,N_5483,N_5888);
nand U14205 (N_14205,N_8884,N_5960);
nor U14206 (N_14206,N_8407,N_9156);
nor U14207 (N_14207,N_7766,N_9698);
or U14208 (N_14208,N_6041,N_5153);
or U14209 (N_14209,N_6741,N_6847);
nand U14210 (N_14210,N_9114,N_5885);
or U14211 (N_14211,N_7998,N_8205);
nand U14212 (N_14212,N_7214,N_6165);
nor U14213 (N_14213,N_9939,N_6164);
or U14214 (N_14214,N_9534,N_7883);
nor U14215 (N_14215,N_7816,N_7252);
xnor U14216 (N_14216,N_9685,N_7877);
xor U14217 (N_14217,N_7914,N_6067);
or U14218 (N_14218,N_6748,N_8492);
or U14219 (N_14219,N_9973,N_7428);
and U14220 (N_14220,N_8798,N_5673);
or U14221 (N_14221,N_5455,N_6112);
and U14222 (N_14222,N_6312,N_9675);
xnor U14223 (N_14223,N_5265,N_6808);
and U14224 (N_14224,N_6630,N_8711);
nor U14225 (N_14225,N_5769,N_7520);
nor U14226 (N_14226,N_5293,N_7276);
nand U14227 (N_14227,N_9136,N_9366);
and U14228 (N_14228,N_6790,N_6146);
xor U14229 (N_14229,N_9764,N_6949);
and U14230 (N_14230,N_8535,N_6102);
nor U14231 (N_14231,N_7443,N_5344);
or U14232 (N_14232,N_7342,N_5975);
and U14233 (N_14233,N_6549,N_7130);
xor U14234 (N_14234,N_8418,N_7013);
nand U14235 (N_14235,N_7691,N_8746);
and U14236 (N_14236,N_7887,N_6715);
nor U14237 (N_14237,N_9018,N_7843);
and U14238 (N_14238,N_8200,N_6606);
nor U14239 (N_14239,N_6447,N_9830);
nand U14240 (N_14240,N_6626,N_8048);
and U14241 (N_14241,N_6575,N_9717);
or U14242 (N_14242,N_8495,N_8463);
xor U14243 (N_14243,N_7201,N_7799);
nand U14244 (N_14244,N_8415,N_5030);
nand U14245 (N_14245,N_5638,N_8430);
nand U14246 (N_14246,N_6377,N_8835);
or U14247 (N_14247,N_6710,N_7874);
and U14248 (N_14248,N_6464,N_6305);
nor U14249 (N_14249,N_8391,N_8902);
xnor U14250 (N_14250,N_9890,N_7059);
nand U14251 (N_14251,N_6177,N_9542);
and U14252 (N_14252,N_6448,N_5270);
xnor U14253 (N_14253,N_5025,N_5746);
xnor U14254 (N_14254,N_5164,N_7470);
or U14255 (N_14255,N_9555,N_6339);
or U14256 (N_14256,N_5868,N_7617);
xnor U14257 (N_14257,N_7990,N_5255);
and U14258 (N_14258,N_5348,N_9568);
and U14259 (N_14259,N_8379,N_6715);
nand U14260 (N_14260,N_9955,N_8830);
or U14261 (N_14261,N_9625,N_8281);
nand U14262 (N_14262,N_9790,N_9211);
xor U14263 (N_14263,N_9855,N_6614);
nand U14264 (N_14264,N_6599,N_7229);
or U14265 (N_14265,N_7747,N_9819);
nand U14266 (N_14266,N_8576,N_9524);
and U14267 (N_14267,N_5372,N_6145);
xnor U14268 (N_14268,N_6496,N_9586);
nand U14269 (N_14269,N_7938,N_7056);
xnor U14270 (N_14270,N_6611,N_5531);
nand U14271 (N_14271,N_9420,N_5413);
or U14272 (N_14272,N_9721,N_9078);
xnor U14273 (N_14273,N_6393,N_8928);
and U14274 (N_14274,N_7957,N_8742);
nand U14275 (N_14275,N_8917,N_5226);
xor U14276 (N_14276,N_8997,N_7263);
or U14277 (N_14277,N_9288,N_6644);
nand U14278 (N_14278,N_8454,N_6486);
or U14279 (N_14279,N_7323,N_8895);
nand U14280 (N_14280,N_9894,N_9731);
and U14281 (N_14281,N_6908,N_9273);
and U14282 (N_14282,N_5437,N_5727);
nor U14283 (N_14283,N_5802,N_6717);
xor U14284 (N_14284,N_9670,N_7429);
nand U14285 (N_14285,N_7003,N_5321);
nor U14286 (N_14286,N_5325,N_6771);
and U14287 (N_14287,N_8160,N_7931);
xnor U14288 (N_14288,N_9596,N_6746);
and U14289 (N_14289,N_6895,N_9861);
nor U14290 (N_14290,N_5595,N_9380);
xnor U14291 (N_14291,N_7604,N_5417);
xnor U14292 (N_14292,N_9729,N_6939);
nor U14293 (N_14293,N_8195,N_7378);
xor U14294 (N_14294,N_8812,N_7311);
xor U14295 (N_14295,N_5478,N_7334);
xnor U14296 (N_14296,N_9283,N_6549);
nand U14297 (N_14297,N_5369,N_6202);
or U14298 (N_14298,N_6070,N_8134);
or U14299 (N_14299,N_8823,N_8001);
nand U14300 (N_14300,N_6556,N_6483);
and U14301 (N_14301,N_6145,N_7248);
nand U14302 (N_14302,N_6448,N_9602);
or U14303 (N_14303,N_5213,N_5491);
nor U14304 (N_14304,N_9552,N_8504);
nor U14305 (N_14305,N_9980,N_5518);
nand U14306 (N_14306,N_8307,N_5456);
nor U14307 (N_14307,N_9719,N_5471);
xor U14308 (N_14308,N_8241,N_8059);
xnor U14309 (N_14309,N_8566,N_8595);
nand U14310 (N_14310,N_7428,N_5985);
or U14311 (N_14311,N_7116,N_5151);
nand U14312 (N_14312,N_6167,N_7691);
xor U14313 (N_14313,N_6016,N_8967);
or U14314 (N_14314,N_6263,N_9456);
or U14315 (N_14315,N_7496,N_8037);
or U14316 (N_14316,N_7872,N_5965);
or U14317 (N_14317,N_9707,N_9236);
and U14318 (N_14318,N_5472,N_7206);
nor U14319 (N_14319,N_6988,N_6519);
or U14320 (N_14320,N_6222,N_7044);
and U14321 (N_14321,N_7310,N_8641);
xor U14322 (N_14322,N_9317,N_6947);
or U14323 (N_14323,N_7796,N_8631);
xor U14324 (N_14324,N_6192,N_5365);
or U14325 (N_14325,N_7586,N_5683);
xor U14326 (N_14326,N_6379,N_8691);
and U14327 (N_14327,N_8195,N_9717);
and U14328 (N_14328,N_6496,N_9885);
nand U14329 (N_14329,N_5121,N_8110);
or U14330 (N_14330,N_6317,N_9530);
and U14331 (N_14331,N_8450,N_8386);
nand U14332 (N_14332,N_7911,N_7313);
nand U14333 (N_14333,N_7263,N_5949);
xor U14334 (N_14334,N_7694,N_9295);
nor U14335 (N_14335,N_8376,N_5323);
xnor U14336 (N_14336,N_8182,N_9847);
and U14337 (N_14337,N_7610,N_6758);
and U14338 (N_14338,N_6095,N_7416);
xnor U14339 (N_14339,N_7313,N_6652);
nor U14340 (N_14340,N_6838,N_9191);
nand U14341 (N_14341,N_8472,N_5283);
or U14342 (N_14342,N_8004,N_7064);
nor U14343 (N_14343,N_7716,N_8081);
nor U14344 (N_14344,N_6609,N_6889);
nand U14345 (N_14345,N_5262,N_9879);
or U14346 (N_14346,N_7098,N_5693);
nand U14347 (N_14347,N_9436,N_5165);
xor U14348 (N_14348,N_8220,N_7158);
nor U14349 (N_14349,N_9085,N_6047);
xor U14350 (N_14350,N_5094,N_6198);
and U14351 (N_14351,N_9569,N_8589);
or U14352 (N_14352,N_5986,N_9523);
nor U14353 (N_14353,N_8698,N_6747);
xor U14354 (N_14354,N_6452,N_6515);
or U14355 (N_14355,N_7455,N_8010);
or U14356 (N_14356,N_9529,N_7329);
or U14357 (N_14357,N_5555,N_9589);
xnor U14358 (N_14358,N_6230,N_6522);
nand U14359 (N_14359,N_7248,N_6485);
or U14360 (N_14360,N_8839,N_9221);
or U14361 (N_14361,N_8418,N_9114);
nand U14362 (N_14362,N_5098,N_7403);
nor U14363 (N_14363,N_5745,N_9823);
xor U14364 (N_14364,N_9939,N_6953);
or U14365 (N_14365,N_6083,N_9189);
nor U14366 (N_14366,N_7748,N_5367);
or U14367 (N_14367,N_7552,N_6182);
or U14368 (N_14368,N_5836,N_7788);
nand U14369 (N_14369,N_6874,N_9358);
xor U14370 (N_14370,N_5460,N_8266);
xor U14371 (N_14371,N_6625,N_6435);
nor U14372 (N_14372,N_7132,N_9836);
xor U14373 (N_14373,N_5745,N_6920);
nor U14374 (N_14374,N_8895,N_8525);
and U14375 (N_14375,N_7305,N_7826);
nor U14376 (N_14376,N_5618,N_5398);
nor U14377 (N_14377,N_8291,N_6925);
xnor U14378 (N_14378,N_6805,N_8624);
nor U14379 (N_14379,N_9802,N_8897);
or U14380 (N_14380,N_9170,N_6459);
and U14381 (N_14381,N_6786,N_5786);
xor U14382 (N_14382,N_8243,N_7374);
or U14383 (N_14383,N_8880,N_6729);
nand U14384 (N_14384,N_9335,N_9795);
nor U14385 (N_14385,N_8314,N_9577);
nand U14386 (N_14386,N_5142,N_9953);
or U14387 (N_14387,N_6633,N_9336);
nor U14388 (N_14388,N_6754,N_7714);
or U14389 (N_14389,N_6114,N_5007);
or U14390 (N_14390,N_5486,N_5979);
xnor U14391 (N_14391,N_5987,N_7151);
nor U14392 (N_14392,N_6841,N_5508);
nor U14393 (N_14393,N_7253,N_6271);
xor U14394 (N_14394,N_6920,N_8864);
and U14395 (N_14395,N_9072,N_6424);
or U14396 (N_14396,N_7790,N_5667);
xor U14397 (N_14397,N_7629,N_8441);
or U14398 (N_14398,N_6849,N_8050);
or U14399 (N_14399,N_8357,N_7060);
nand U14400 (N_14400,N_6358,N_6111);
and U14401 (N_14401,N_6639,N_8227);
nor U14402 (N_14402,N_8853,N_5162);
xnor U14403 (N_14403,N_5347,N_6406);
or U14404 (N_14404,N_9628,N_9553);
or U14405 (N_14405,N_9182,N_5240);
xor U14406 (N_14406,N_9590,N_8044);
nor U14407 (N_14407,N_7630,N_5175);
and U14408 (N_14408,N_5719,N_5678);
and U14409 (N_14409,N_5988,N_8198);
xor U14410 (N_14410,N_6976,N_6561);
nor U14411 (N_14411,N_8096,N_5121);
xor U14412 (N_14412,N_7123,N_7415);
xor U14413 (N_14413,N_6985,N_9516);
or U14414 (N_14414,N_6818,N_8286);
nand U14415 (N_14415,N_7608,N_6246);
nor U14416 (N_14416,N_8642,N_6360);
xor U14417 (N_14417,N_9822,N_7581);
and U14418 (N_14418,N_6305,N_7369);
nand U14419 (N_14419,N_7577,N_9113);
xor U14420 (N_14420,N_5600,N_8545);
xnor U14421 (N_14421,N_9988,N_8380);
xnor U14422 (N_14422,N_8382,N_7030);
nor U14423 (N_14423,N_5286,N_6669);
and U14424 (N_14424,N_5195,N_6594);
xor U14425 (N_14425,N_5009,N_5105);
and U14426 (N_14426,N_5118,N_8056);
nor U14427 (N_14427,N_6653,N_6270);
or U14428 (N_14428,N_6092,N_6808);
and U14429 (N_14429,N_8504,N_6495);
nand U14430 (N_14430,N_7019,N_9084);
nor U14431 (N_14431,N_9140,N_8525);
or U14432 (N_14432,N_7628,N_6495);
and U14433 (N_14433,N_8957,N_6492);
nor U14434 (N_14434,N_6711,N_5126);
nand U14435 (N_14435,N_5324,N_8417);
xnor U14436 (N_14436,N_6195,N_6901);
or U14437 (N_14437,N_6558,N_6041);
xnor U14438 (N_14438,N_8707,N_8485);
and U14439 (N_14439,N_7059,N_9632);
xor U14440 (N_14440,N_9416,N_6976);
nor U14441 (N_14441,N_6380,N_8425);
xnor U14442 (N_14442,N_7506,N_7339);
nand U14443 (N_14443,N_9773,N_5099);
nand U14444 (N_14444,N_5872,N_5649);
and U14445 (N_14445,N_7484,N_9609);
nand U14446 (N_14446,N_6870,N_5753);
nor U14447 (N_14447,N_8816,N_6399);
and U14448 (N_14448,N_7685,N_5908);
and U14449 (N_14449,N_7235,N_5558);
or U14450 (N_14450,N_9591,N_7042);
and U14451 (N_14451,N_6279,N_6748);
xnor U14452 (N_14452,N_5104,N_8708);
nand U14453 (N_14453,N_6388,N_6618);
nand U14454 (N_14454,N_9693,N_8658);
and U14455 (N_14455,N_6479,N_8315);
or U14456 (N_14456,N_7557,N_9916);
or U14457 (N_14457,N_6399,N_6454);
or U14458 (N_14458,N_6666,N_5967);
nand U14459 (N_14459,N_8114,N_6653);
and U14460 (N_14460,N_9950,N_8627);
nand U14461 (N_14461,N_6203,N_5433);
or U14462 (N_14462,N_9761,N_9624);
nor U14463 (N_14463,N_6384,N_6042);
nand U14464 (N_14464,N_5012,N_8674);
or U14465 (N_14465,N_5132,N_5532);
nor U14466 (N_14466,N_6602,N_5888);
xnor U14467 (N_14467,N_7645,N_8542);
xor U14468 (N_14468,N_5936,N_7712);
nand U14469 (N_14469,N_8048,N_9611);
or U14470 (N_14470,N_5875,N_9719);
nor U14471 (N_14471,N_8708,N_9577);
and U14472 (N_14472,N_9665,N_8827);
xnor U14473 (N_14473,N_7836,N_9664);
and U14474 (N_14474,N_9545,N_6083);
nor U14475 (N_14475,N_5737,N_6681);
xnor U14476 (N_14476,N_7694,N_5255);
nand U14477 (N_14477,N_6475,N_9875);
and U14478 (N_14478,N_8537,N_6723);
xor U14479 (N_14479,N_5564,N_6989);
xnor U14480 (N_14480,N_8655,N_6947);
or U14481 (N_14481,N_6313,N_7621);
nor U14482 (N_14482,N_6218,N_5881);
nor U14483 (N_14483,N_8634,N_5688);
and U14484 (N_14484,N_9946,N_8261);
nand U14485 (N_14485,N_6269,N_5331);
or U14486 (N_14486,N_7841,N_6725);
nor U14487 (N_14487,N_8469,N_8102);
or U14488 (N_14488,N_9713,N_7335);
xor U14489 (N_14489,N_5983,N_6034);
xor U14490 (N_14490,N_7079,N_5442);
xor U14491 (N_14491,N_7278,N_9190);
xnor U14492 (N_14492,N_8933,N_5217);
and U14493 (N_14493,N_6017,N_8987);
or U14494 (N_14494,N_9637,N_8628);
and U14495 (N_14495,N_9621,N_9506);
nand U14496 (N_14496,N_5921,N_8920);
nand U14497 (N_14497,N_7557,N_8499);
and U14498 (N_14498,N_5120,N_6109);
or U14499 (N_14499,N_7201,N_9682);
and U14500 (N_14500,N_8589,N_7775);
xnor U14501 (N_14501,N_9626,N_9539);
nand U14502 (N_14502,N_5419,N_5593);
xnor U14503 (N_14503,N_5783,N_5592);
nand U14504 (N_14504,N_5036,N_5549);
xor U14505 (N_14505,N_6030,N_8083);
or U14506 (N_14506,N_9432,N_7136);
nor U14507 (N_14507,N_7957,N_6499);
or U14508 (N_14508,N_5218,N_5999);
xnor U14509 (N_14509,N_9791,N_8166);
nand U14510 (N_14510,N_8985,N_6160);
nor U14511 (N_14511,N_8211,N_7477);
nand U14512 (N_14512,N_9126,N_9301);
and U14513 (N_14513,N_7699,N_8269);
or U14514 (N_14514,N_8279,N_6052);
nand U14515 (N_14515,N_8306,N_6321);
nand U14516 (N_14516,N_6225,N_6610);
nand U14517 (N_14517,N_5354,N_6594);
nor U14518 (N_14518,N_5990,N_9757);
nand U14519 (N_14519,N_9030,N_7982);
xnor U14520 (N_14520,N_7015,N_7605);
or U14521 (N_14521,N_7888,N_6233);
xor U14522 (N_14522,N_7219,N_6620);
nand U14523 (N_14523,N_9384,N_8906);
nand U14524 (N_14524,N_9958,N_5209);
and U14525 (N_14525,N_7229,N_8972);
and U14526 (N_14526,N_6510,N_8130);
nand U14527 (N_14527,N_5659,N_6021);
nand U14528 (N_14528,N_9474,N_5424);
and U14529 (N_14529,N_6564,N_6386);
xnor U14530 (N_14530,N_8488,N_8590);
nor U14531 (N_14531,N_5945,N_5736);
xnor U14532 (N_14532,N_7343,N_6114);
nor U14533 (N_14533,N_5107,N_8925);
xnor U14534 (N_14534,N_7979,N_7831);
or U14535 (N_14535,N_5757,N_6509);
and U14536 (N_14536,N_9977,N_6146);
or U14537 (N_14537,N_7310,N_6206);
nor U14538 (N_14538,N_8886,N_5618);
and U14539 (N_14539,N_9116,N_5514);
and U14540 (N_14540,N_7650,N_9617);
xnor U14541 (N_14541,N_6806,N_9778);
nand U14542 (N_14542,N_7774,N_6649);
and U14543 (N_14543,N_9455,N_7156);
or U14544 (N_14544,N_5349,N_6367);
xor U14545 (N_14545,N_6232,N_5938);
nand U14546 (N_14546,N_8905,N_9039);
or U14547 (N_14547,N_5526,N_6599);
and U14548 (N_14548,N_6182,N_7276);
nor U14549 (N_14549,N_9082,N_9302);
nand U14550 (N_14550,N_9195,N_8707);
nor U14551 (N_14551,N_6900,N_6752);
and U14552 (N_14552,N_7248,N_7871);
and U14553 (N_14553,N_7443,N_7285);
nand U14554 (N_14554,N_6825,N_6060);
nand U14555 (N_14555,N_8846,N_8594);
xnor U14556 (N_14556,N_7219,N_5118);
or U14557 (N_14557,N_8768,N_5387);
nor U14558 (N_14558,N_9268,N_6570);
and U14559 (N_14559,N_5993,N_8237);
or U14560 (N_14560,N_8613,N_7238);
xnor U14561 (N_14561,N_9999,N_8389);
nand U14562 (N_14562,N_9197,N_7133);
xor U14563 (N_14563,N_5768,N_5814);
and U14564 (N_14564,N_5194,N_8181);
and U14565 (N_14565,N_6082,N_5090);
nor U14566 (N_14566,N_6995,N_7677);
xor U14567 (N_14567,N_8352,N_6258);
nor U14568 (N_14568,N_8635,N_5177);
nor U14569 (N_14569,N_9969,N_7545);
or U14570 (N_14570,N_7319,N_7128);
or U14571 (N_14571,N_8380,N_9502);
or U14572 (N_14572,N_7905,N_8020);
nor U14573 (N_14573,N_9851,N_8953);
nand U14574 (N_14574,N_9714,N_5374);
nor U14575 (N_14575,N_5524,N_9596);
or U14576 (N_14576,N_7162,N_6410);
nor U14577 (N_14577,N_5489,N_9159);
or U14578 (N_14578,N_7161,N_8440);
nand U14579 (N_14579,N_8319,N_6709);
xor U14580 (N_14580,N_7175,N_5096);
nor U14581 (N_14581,N_7456,N_5458);
and U14582 (N_14582,N_7102,N_8064);
nor U14583 (N_14583,N_8096,N_9073);
nor U14584 (N_14584,N_9148,N_9069);
nand U14585 (N_14585,N_9905,N_6761);
and U14586 (N_14586,N_6156,N_6881);
nor U14587 (N_14587,N_6358,N_5391);
or U14588 (N_14588,N_9340,N_6530);
nor U14589 (N_14589,N_9345,N_5571);
xor U14590 (N_14590,N_6604,N_9163);
or U14591 (N_14591,N_6170,N_5582);
nor U14592 (N_14592,N_5928,N_6351);
nor U14593 (N_14593,N_8624,N_6637);
xor U14594 (N_14594,N_5777,N_9351);
or U14595 (N_14595,N_5746,N_8106);
and U14596 (N_14596,N_6579,N_6436);
or U14597 (N_14597,N_7011,N_9186);
xnor U14598 (N_14598,N_9969,N_5502);
xor U14599 (N_14599,N_8416,N_7849);
nor U14600 (N_14600,N_6213,N_6565);
nand U14601 (N_14601,N_7183,N_7480);
and U14602 (N_14602,N_5220,N_6873);
nor U14603 (N_14603,N_6743,N_6409);
and U14604 (N_14604,N_7609,N_8405);
nor U14605 (N_14605,N_8734,N_5018);
or U14606 (N_14606,N_8484,N_8263);
nand U14607 (N_14607,N_9996,N_5942);
nand U14608 (N_14608,N_7137,N_8402);
or U14609 (N_14609,N_9153,N_7706);
nor U14610 (N_14610,N_5992,N_6251);
xor U14611 (N_14611,N_9569,N_8500);
and U14612 (N_14612,N_7366,N_7552);
nor U14613 (N_14613,N_6238,N_9687);
xor U14614 (N_14614,N_9285,N_5966);
xor U14615 (N_14615,N_6722,N_7104);
or U14616 (N_14616,N_6376,N_9833);
nand U14617 (N_14617,N_8270,N_6299);
or U14618 (N_14618,N_5351,N_9925);
nand U14619 (N_14619,N_6339,N_7767);
xor U14620 (N_14620,N_7991,N_9470);
nand U14621 (N_14621,N_7377,N_9404);
xnor U14622 (N_14622,N_6447,N_7878);
nand U14623 (N_14623,N_8639,N_8392);
nor U14624 (N_14624,N_8616,N_7287);
and U14625 (N_14625,N_5749,N_8199);
nand U14626 (N_14626,N_7828,N_9113);
or U14627 (N_14627,N_8090,N_5937);
nand U14628 (N_14628,N_8195,N_5987);
and U14629 (N_14629,N_5870,N_8145);
or U14630 (N_14630,N_7749,N_9900);
xnor U14631 (N_14631,N_6247,N_9687);
and U14632 (N_14632,N_9898,N_7196);
nand U14633 (N_14633,N_8846,N_7843);
and U14634 (N_14634,N_9415,N_8683);
and U14635 (N_14635,N_7186,N_7808);
nand U14636 (N_14636,N_6111,N_7899);
nor U14637 (N_14637,N_8956,N_5956);
nor U14638 (N_14638,N_9193,N_7977);
or U14639 (N_14639,N_9412,N_7208);
or U14640 (N_14640,N_5058,N_7042);
and U14641 (N_14641,N_5631,N_8662);
nor U14642 (N_14642,N_9059,N_6711);
xnor U14643 (N_14643,N_8595,N_7931);
nor U14644 (N_14644,N_9067,N_7247);
nand U14645 (N_14645,N_6154,N_7996);
nor U14646 (N_14646,N_9157,N_5455);
nor U14647 (N_14647,N_5114,N_8139);
or U14648 (N_14648,N_7050,N_7912);
nand U14649 (N_14649,N_7039,N_9329);
nand U14650 (N_14650,N_8913,N_5976);
xor U14651 (N_14651,N_9415,N_5128);
nand U14652 (N_14652,N_5925,N_5939);
nand U14653 (N_14653,N_5444,N_7811);
and U14654 (N_14654,N_6970,N_6747);
and U14655 (N_14655,N_9168,N_7616);
and U14656 (N_14656,N_9010,N_6483);
and U14657 (N_14657,N_7291,N_9455);
nor U14658 (N_14658,N_5588,N_5345);
and U14659 (N_14659,N_8924,N_9165);
nand U14660 (N_14660,N_7076,N_5037);
nand U14661 (N_14661,N_7164,N_6608);
and U14662 (N_14662,N_5701,N_9438);
and U14663 (N_14663,N_7807,N_8130);
nor U14664 (N_14664,N_6162,N_8611);
nor U14665 (N_14665,N_6440,N_7286);
xor U14666 (N_14666,N_6255,N_9951);
nand U14667 (N_14667,N_6672,N_7023);
xnor U14668 (N_14668,N_8209,N_8204);
nor U14669 (N_14669,N_6485,N_6655);
or U14670 (N_14670,N_6937,N_8207);
nor U14671 (N_14671,N_7188,N_5240);
or U14672 (N_14672,N_8952,N_5524);
xor U14673 (N_14673,N_5225,N_6681);
and U14674 (N_14674,N_5654,N_5499);
nor U14675 (N_14675,N_6178,N_9071);
and U14676 (N_14676,N_8190,N_5250);
nor U14677 (N_14677,N_6766,N_7500);
xnor U14678 (N_14678,N_7300,N_9977);
xor U14679 (N_14679,N_8661,N_5856);
and U14680 (N_14680,N_9023,N_5337);
nand U14681 (N_14681,N_8481,N_5011);
nand U14682 (N_14682,N_6613,N_6090);
and U14683 (N_14683,N_9154,N_6280);
xor U14684 (N_14684,N_7062,N_5620);
or U14685 (N_14685,N_7397,N_9507);
or U14686 (N_14686,N_5703,N_5211);
or U14687 (N_14687,N_8714,N_5603);
and U14688 (N_14688,N_9847,N_9226);
xor U14689 (N_14689,N_6664,N_5701);
and U14690 (N_14690,N_6533,N_8331);
and U14691 (N_14691,N_6884,N_9218);
or U14692 (N_14692,N_8437,N_9666);
xor U14693 (N_14693,N_8921,N_9631);
or U14694 (N_14694,N_5705,N_7696);
nor U14695 (N_14695,N_7645,N_8647);
or U14696 (N_14696,N_6812,N_9685);
nand U14697 (N_14697,N_7873,N_6922);
or U14698 (N_14698,N_9907,N_6545);
nand U14699 (N_14699,N_9285,N_7212);
nand U14700 (N_14700,N_5869,N_8401);
and U14701 (N_14701,N_7847,N_9482);
xor U14702 (N_14702,N_8812,N_5971);
or U14703 (N_14703,N_7522,N_5359);
nand U14704 (N_14704,N_8673,N_6089);
or U14705 (N_14705,N_5212,N_5294);
xor U14706 (N_14706,N_7811,N_9604);
nor U14707 (N_14707,N_8233,N_6304);
nand U14708 (N_14708,N_6259,N_6548);
nand U14709 (N_14709,N_6145,N_8482);
nor U14710 (N_14710,N_5511,N_8461);
or U14711 (N_14711,N_6218,N_9416);
nor U14712 (N_14712,N_7504,N_6182);
xor U14713 (N_14713,N_8289,N_8319);
or U14714 (N_14714,N_8538,N_9846);
xnor U14715 (N_14715,N_7435,N_7853);
nand U14716 (N_14716,N_9837,N_5596);
nor U14717 (N_14717,N_8296,N_7445);
nor U14718 (N_14718,N_7996,N_9841);
xnor U14719 (N_14719,N_8714,N_5781);
xnor U14720 (N_14720,N_9160,N_5401);
xor U14721 (N_14721,N_7783,N_7652);
nand U14722 (N_14722,N_9787,N_6960);
nand U14723 (N_14723,N_5417,N_8649);
nand U14724 (N_14724,N_9729,N_7907);
and U14725 (N_14725,N_9862,N_7989);
xnor U14726 (N_14726,N_9384,N_7027);
xor U14727 (N_14727,N_9142,N_9516);
nand U14728 (N_14728,N_6780,N_6611);
and U14729 (N_14729,N_6479,N_6579);
nor U14730 (N_14730,N_9659,N_5410);
nand U14731 (N_14731,N_8983,N_7991);
xnor U14732 (N_14732,N_7452,N_8877);
nor U14733 (N_14733,N_7444,N_7038);
nor U14734 (N_14734,N_6942,N_6392);
xor U14735 (N_14735,N_5813,N_7527);
xnor U14736 (N_14736,N_5090,N_6249);
nand U14737 (N_14737,N_8403,N_7122);
xor U14738 (N_14738,N_6406,N_5536);
nor U14739 (N_14739,N_9421,N_8496);
xnor U14740 (N_14740,N_5794,N_6969);
or U14741 (N_14741,N_7207,N_8848);
nand U14742 (N_14742,N_8465,N_8226);
nand U14743 (N_14743,N_9954,N_7592);
or U14744 (N_14744,N_9660,N_5166);
xnor U14745 (N_14745,N_8642,N_7172);
and U14746 (N_14746,N_5495,N_5173);
xor U14747 (N_14747,N_6646,N_6311);
or U14748 (N_14748,N_9176,N_5141);
nand U14749 (N_14749,N_7790,N_5494);
xor U14750 (N_14750,N_7219,N_6574);
xnor U14751 (N_14751,N_5056,N_5003);
or U14752 (N_14752,N_8843,N_5750);
xor U14753 (N_14753,N_6536,N_9932);
nor U14754 (N_14754,N_5101,N_7421);
xnor U14755 (N_14755,N_6673,N_7473);
nor U14756 (N_14756,N_9708,N_8059);
nor U14757 (N_14757,N_9259,N_6013);
nor U14758 (N_14758,N_5081,N_8617);
nand U14759 (N_14759,N_6817,N_5574);
and U14760 (N_14760,N_7725,N_9832);
or U14761 (N_14761,N_9538,N_7189);
nand U14762 (N_14762,N_7829,N_7509);
and U14763 (N_14763,N_9685,N_7762);
and U14764 (N_14764,N_8227,N_6971);
or U14765 (N_14765,N_6389,N_6907);
nand U14766 (N_14766,N_7809,N_6899);
xor U14767 (N_14767,N_8112,N_9625);
nor U14768 (N_14768,N_9727,N_5940);
xor U14769 (N_14769,N_6019,N_5732);
xor U14770 (N_14770,N_9269,N_8394);
or U14771 (N_14771,N_5971,N_6971);
and U14772 (N_14772,N_7751,N_7550);
nor U14773 (N_14773,N_8327,N_8813);
and U14774 (N_14774,N_8839,N_7223);
xor U14775 (N_14775,N_6187,N_6299);
xor U14776 (N_14776,N_7718,N_9964);
nor U14777 (N_14777,N_5306,N_7666);
or U14778 (N_14778,N_9446,N_7029);
and U14779 (N_14779,N_6587,N_5631);
nor U14780 (N_14780,N_6916,N_5998);
xnor U14781 (N_14781,N_7457,N_6897);
and U14782 (N_14782,N_7946,N_8230);
xnor U14783 (N_14783,N_5711,N_5994);
and U14784 (N_14784,N_9680,N_8144);
xnor U14785 (N_14785,N_7420,N_6039);
or U14786 (N_14786,N_6863,N_9891);
and U14787 (N_14787,N_6612,N_5279);
nand U14788 (N_14788,N_9172,N_5876);
xnor U14789 (N_14789,N_6134,N_8105);
nand U14790 (N_14790,N_9738,N_9172);
xnor U14791 (N_14791,N_5936,N_9841);
xor U14792 (N_14792,N_9135,N_6302);
nor U14793 (N_14793,N_9191,N_5605);
nor U14794 (N_14794,N_8268,N_7582);
nor U14795 (N_14795,N_5989,N_8087);
and U14796 (N_14796,N_9366,N_6417);
or U14797 (N_14797,N_7481,N_7097);
nand U14798 (N_14798,N_7791,N_8324);
nor U14799 (N_14799,N_9229,N_8650);
xor U14800 (N_14800,N_9748,N_6683);
and U14801 (N_14801,N_9203,N_7463);
and U14802 (N_14802,N_8364,N_8472);
and U14803 (N_14803,N_7472,N_5849);
and U14804 (N_14804,N_5201,N_6791);
nand U14805 (N_14805,N_8003,N_5896);
xor U14806 (N_14806,N_5058,N_8169);
nand U14807 (N_14807,N_8203,N_6760);
nor U14808 (N_14808,N_6966,N_5451);
or U14809 (N_14809,N_5059,N_5743);
xor U14810 (N_14810,N_8320,N_7264);
or U14811 (N_14811,N_9396,N_7777);
nor U14812 (N_14812,N_8113,N_5642);
nand U14813 (N_14813,N_7194,N_9021);
nor U14814 (N_14814,N_7845,N_7684);
xor U14815 (N_14815,N_9564,N_8613);
xor U14816 (N_14816,N_8109,N_5197);
nand U14817 (N_14817,N_8732,N_9489);
nor U14818 (N_14818,N_5206,N_9330);
nand U14819 (N_14819,N_6200,N_6074);
nand U14820 (N_14820,N_5108,N_7711);
nor U14821 (N_14821,N_8043,N_7460);
xor U14822 (N_14822,N_9238,N_8278);
and U14823 (N_14823,N_9922,N_6520);
or U14824 (N_14824,N_9437,N_8169);
and U14825 (N_14825,N_6982,N_5485);
or U14826 (N_14826,N_8828,N_7914);
nor U14827 (N_14827,N_8411,N_5844);
and U14828 (N_14828,N_9297,N_8486);
nor U14829 (N_14829,N_6998,N_8413);
and U14830 (N_14830,N_6813,N_9033);
nand U14831 (N_14831,N_5311,N_6807);
nor U14832 (N_14832,N_9121,N_8185);
or U14833 (N_14833,N_7349,N_9889);
xnor U14834 (N_14834,N_8164,N_8909);
xnor U14835 (N_14835,N_7576,N_8048);
xor U14836 (N_14836,N_7717,N_5834);
nand U14837 (N_14837,N_9848,N_9932);
nand U14838 (N_14838,N_8824,N_8351);
or U14839 (N_14839,N_9956,N_5888);
nor U14840 (N_14840,N_8688,N_5269);
xnor U14841 (N_14841,N_8971,N_8893);
nor U14842 (N_14842,N_9800,N_7594);
nor U14843 (N_14843,N_6676,N_8973);
nand U14844 (N_14844,N_5796,N_5961);
xnor U14845 (N_14845,N_9480,N_5514);
nor U14846 (N_14846,N_7015,N_8269);
nor U14847 (N_14847,N_5594,N_7500);
or U14848 (N_14848,N_8745,N_6681);
and U14849 (N_14849,N_9712,N_5597);
and U14850 (N_14850,N_7194,N_7432);
xnor U14851 (N_14851,N_9253,N_8050);
nor U14852 (N_14852,N_7223,N_6115);
nand U14853 (N_14853,N_5053,N_7402);
and U14854 (N_14854,N_9118,N_8614);
xor U14855 (N_14855,N_9559,N_9869);
nor U14856 (N_14856,N_8085,N_5201);
nor U14857 (N_14857,N_5763,N_8067);
nor U14858 (N_14858,N_6207,N_8547);
nor U14859 (N_14859,N_5243,N_8983);
and U14860 (N_14860,N_5718,N_7112);
and U14861 (N_14861,N_6291,N_9542);
nor U14862 (N_14862,N_9481,N_5784);
and U14863 (N_14863,N_6761,N_7850);
and U14864 (N_14864,N_8343,N_8870);
nor U14865 (N_14865,N_7049,N_6381);
and U14866 (N_14866,N_7014,N_7316);
nor U14867 (N_14867,N_7660,N_6795);
or U14868 (N_14868,N_7422,N_7524);
nand U14869 (N_14869,N_6168,N_8803);
xor U14870 (N_14870,N_5450,N_5778);
nand U14871 (N_14871,N_7758,N_6486);
or U14872 (N_14872,N_5929,N_8298);
nor U14873 (N_14873,N_8446,N_8776);
or U14874 (N_14874,N_6892,N_5072);
nand U14875 (N_14875,N_5411,N_9313);
nor U14876 (N_14876,N_7180,N_7008);
nand U14877 (N_14877,N_6061,N_9664);
xnor U14878 (N_14878,N_6629,N_9527);
nor U14879 (N_14879,N_9791,N_7717);
and U14880 (N_14880,N_9054,N_5687);
or U14881 (N_14881,N_7946,N_9901);
nand U14882 (N_14882,N_5099,N_8431);
nand U14883 (N_14883,N_5081,N_7833);
and U14884 (N_14884,N_5988,N_8347);
nand U14885 (N_14885,N_6974,N_6091);
and U14886 (N_14886,N_8800,N_8725);
or U14887 (N_14887,N_9120,N_7091);
nor U14888 (N_14888,N_7959,N_9091);
nor U14889 (N_14889,N_9947,N_7558);
nand U14890 (N_14890,N_5821,N_6448);
nor U14891 (N_14891,N_7568,N_8215);
nand U14892 (N_14892,N_6501,N_9628);
xor U14893 (N_14893,N_6084,N_6067);
or U14894 (N_14894,N_8685,N_7716);
nor U14895 (N_14895,N_7392,N_5473);
nand U14896 (N_14896,N_7414,N_7940);
or U14897 (N_14897,N_5187,N_6634);
nor U14898 (N_14898,N_9494,N_8284);
or U14899 (N_14899,N_5909,N_8888);
or U14900 (N_14900,N_9141,N_8885);
or U14901 (N_14901,N_7949,N_7240);
nand U14902 (N_14902,N_6427,N_6773);
xor U14903 (N_14903,N_7576,N_5413);
and U14904 (N_14904,N_5206,N_5251);
or U14905 (N_14905,N_7987,N_7081);
nand U14906 (N_14906,N_6042,N_5426);
nor U14907 (N_14907,N_8311,N_6051);
xor U14908 (N_14908,N_8430,N_9647);
xnor U14909 (N_14909,N_5925,N_8752);
nor U14910 (N_14910,N_7716,N_9446);
nand U14911 (N_14911,N_8723,N_6438);
nand U14912 (N_14912,N_6036,N_8236);
xor U14913 (N_14913,N_7837,N_7223);
or U14914 (N_14914,N_8741,N_6635);
xor U14915 (N_14915,N_7427,N_9796);
xor U14916 (N_14916,N_8751,N_5751);
xor U14917 (N_14917,N_5387,N_9062);
nor U14918 (N_14918,N_8183,N_9758);
or U14919 (N_14919,N_6435,N_5107);
nor U14920 (N_14920,N_7181,N_6750);
nand U14921 (N_14921,N_9985,N_8672);
or U14922 (N_14922,N_9006,N_5840);
nand U14923 (N_14923,N_9942,N_8804);
and U14924 (N_14924,N_6969,N_6719);
xnor U14925 (N_14925,N_6633,N_5628);
nand U14926 (N_14926,N_9747,N_5028);
nor U14927 (N_14927,N_6102,N_6682);
and U14928 (N_14928,N_5871,N_7825);
nor U14929 (N_14929,N_5922,N_5846);
nand U14930 (N_14930,N_7286,N_9671);
and U14931 (N_14931,N_8255,N_5888);
nand U14932 (N_14932,N_6135,N_9527);
nor U14933 (N_14933,N_5713,N_9677);
nand U14934 (N_14934,N_6655,N_5997);
nor U14935 (N_14935,N_8608,N_8130);
xor U14936 (N_14936,N_8119,N_7468);
xor U14937 (N_14937,N_7295,N_5894);
nor U14938 (N_14938,N_9360,N_6669);
and U14939 (N_14939,N_7511,N_5436);
nand U14940 (N_14940,N_9967,N_7027);
xnor U14941 (N_14941,N_7746,N_8467);
nor U14942 (N_14942,N_9140,N_8123);
nor U14943 (N_14943,N_6813,N_5056);
nand U14944 (N_14944,N_9458,N_8974);
and U14945 (N_14945,N_7673,N_7133);
nor U14946 (N_14946,N_5615,N_5624);
or U14947 (N_14947,N_6923,N_7261);
xor U14948 (N_14948,N_6692,N_8697);
or U14949 (N_14949,N_5221,N_8387);
nand U14950 (N_14950,N_6540,N_6234);
and U14951 (N_14951,N_9123,N_6882);
xor U14952 (N_14952,N_8527,N_9349);
and U14953 (N_14953,N_9100,N_8803);
nand U14954 (N_14954,N_7893,N_7964);
nor U14955 (N_14955,N_6263,N_5641);
nor U14956 (N_14956,N_9808,N_5700);
xor U14957 (N_14957,N_5427,N_8079);
nand U14958 (N_14958,N_8353,N_7974);
nand U14959 (N_14959,N_6646,N_9735);
nand U14960 (N_14960,N_5750,N_5860);
or U14961 (N_14961,N_8480,N_8233);
and U14962 (N_14962,N_8038,N_7225);
xor U14963 (N_14963,N_6283,N_6386);
or U14964 (N_14964,N_7535,N_7369);
nor U14965 (N_14965,N_6154,N_9678);
and U14966 (N_14966,N_5743,N_5086);
nor U14967 (N_14967,N_8332,N_6127);
nor U14968 (N_14968,N_8621,N_9543);
and U14969 (N_14969,N_8312,N_7782);
or U14970 (N_14970,N_5954,N_6618);
nor U14971 (N_14971,N_8727,N_9336);
and U14972 (N_14972,N_6018,N_9541);
nor U14973 (N_14973,N_5694,N_5868);
nor U14974 (N_14974,N_5333,N_9700);
nand U14975 (N_14975,N_6695,N_5194);
and U14976 (N_14976,N_7014,N_7043);
nand U14977 (N_14977,N_9550,N_6861);
xnor U14978 (N_14978,N_6896,N_6151);
or U14979 (N_14979,N_7695,N_9087);
and U14980 (N_14980,N_8922,N_9823);
xnor U14981 (N_14981,N_9269,N_9340);
nand U14982 (N_14982,N_5138,N_5310);
and U14983 (N_14983,N_9966,N_7890);
nor U14984 (N_14984,N_9939,N_6709);
nand U14985 (N_14985,N_9609,N_6824);
and U14986 (N_14986,N_9179,N_8117);
nor U14987 (N_14987,N_7351,N_5132);
nand U14988 (N_14988,N_5232,N_8323);
xor U14989 (N_14989,N_5021,N_7360);
nor U14990 (N_14990,N_7743,N_8979);
xor U14991 (N_14991,N_8846,N_8593);
nand U14992 (N_14992,N_9088,N_9056);
and U14993 (N_14993,N_6193,N_9635);
nand U14994 (N_14994,N_6622,N_9259);
nor U14995 (N_14995,N_9741,N_6252);
nor U14996 (N_14996,N_9704,N_9873);
nand U14997 (N_14997,N_5689,N_5052);
xor U14998 (N_14998,N_7164,N_9224);
nand U14999 (N_14999,N_5007,N_7139);
nor U15000 (N_15000,N_14002,N_13896);
nand U15001 (N_15001,N_10773,N_13853);
nor U15002 (N_15002,N_11455,N_11832);
xor U15003 (N_15003,N_11061,N_10100);
or U15004 (N_15004,N_13841,N_14411);
nand U15005 (N_15005,N_12730,N_13503);
or U15006 (N_15006,N_11349,N_12590);
or U15007 (N_15007,N_11174,N_11271);
and U15008 (N_15008,N_10785,N_14886);
or U15009 (N_15009,N_11816,N_14908);
or U15010 (N_15010,N_10086,N_10066);
xor U15011 (N_15011,N_10740,N_13565);
nand U15012 (N_15012,N_12923,N_14369);
or U15013 (N_15013,N_10595,N_12431);
and U15014 (N_15014,N_10995,N_13519);
and U15015 (N_15015,N_12703,N_14006);
and U15016 (N_15016,N_14813,N_11328);
nand U15017 (N_15017,N_11430,N_14259);
nor U15018 (N_15018,N_12599,N_12309);
xor U15019 (N_15019,N_11092,N_14168);
xor U15020 (N_15020,N_14590,N_10144);
and U15021 (N_15021,N_11436,N_10273);
nor U15022 (N_15022,N_12582,N_12713);
or U15023 (N_15023,N_12931,N_14156);
xnor U15024 (N_15024,N_12992,N_13569);
xnor U15025 (N_15025,N_14715,N_14619);
and U15026 (N_15026,N_10545,N_11711);
xor U15027 (N_15027,N_10102,N_10991);
or U15028 (N_15028,N_11200,N_14032);
nor U15029 (N_15029,N_13136,N_11093);
nand U15030 (N_15030,N_12917,N_10648);
and U15031 (N_15031,N_12797,N_10658);
nor U15032 (N_15032,N_14422,N_11596);
and U15033 (N_15033,N_11965,N_12249);
nor U15034 (N_15034,N_12860,N_11981);
or U15035 (N_15035,N_13393,N_11834);
nor U15036 (N_15036,N_12436,N_14890);
or U15037 (N_15037,N_10623,N_13485);
xor U15038 (N_15038,N_14687,N_10592);
nor U15039 (N_15039,N_11759,N_12176);
nor U15040 (N_15040,N_13017,N_12990);
nand U15041 (N_15041,N_13492,N_10780);
and U15042 (N_15042,N_12639,N_14141);
and U15043 (N_15043,N_13336,N_12754);
or U15044 (N_15044,N_13927,N_10930);
nor U15045 (N_15045,N_11885,N_11539);
nor U15046 (N_15046,N_13852,N_11382);
and U15047 (N_15047,N_11022,N_11968);
or U15048 (N_15048,N_13030,N_12982);
or U15049 (N_15049,N_14497,N_14031);
or U15050 (N_15050,N_10030,N_10566);
xnor U15051 (N_15051,N_14410,N_14821);
nor U15052 (N_15052,N_12547,N_12246);
xor U15053 (N_15053,N_10862,N_12079);
or U15054 (N_15054,N_14246,N_13862);
or U15055 (N_15055,N_14771,N_11369);
xnor U15056 (N_15056,N_11415,N_12089);
nand U15057 (N_15057,N_11219,N_11859);
nand U15058 (N_15058,N_11334,N_13735);
nor U15059 (N_15059,N_10521,N_14210);
xnor U15060 (N_15060,N_13365,N_10868);
and U15061 (N_15061,N_14625,N_12429);
nor U15062 (N_15062,N_11654,N_13311);
nor U15063 (N_15063,N_10768,N_11672);
and U15064 (N_15064,N_13294,N_13300);
xor U15065 (N_15065,N_12961,N_11168);
and U15066 (N_15066,N_14232,N_11404);
or U15067 (N_15067,N_10399,N_10682);
nor U15068 (N_15068,N_10362,N_12913);
or U15069 (N_15069,N_11838,N_12664);
nor U15070 (N_15070,N_14137,N_12343);
nand U15071 (N_15071,N_14209,N_11141);
or U15072 (N_15072,N_13076,N_13900);
or U15073 (N_15073,N_11634,N_14176);
and U15074 (N_15074,N_14289,N_11083);
xnor U15075 (N_15075,N_10116,N_11163);
nand U15076 (N_15076,N_11228,N_11398);
xor U15077 (N_15077,N_10589,N_12061);
or U15078 (N_15078,N_13967,N_12393);
or U15079 (N_15079,N_13904,N_12051);
nand U15080 (N_15080,N_11622,N_14673);
nor U15081 (N_15081,N_13980,N_11186);
or U15082 (N_15082,N_12954,N_11727);
and U15083 (N_15083,N_13032,N_12877);
xnor U15084 (N_15084,N_13221,N_13186);
xnor U15085 (N_15085,N_11331,N_14728);
xnor U15086 (N_15086,N_12516,N_13845);
and U15087 (N_15087,N_12268,N_12785);
or U15088 (N_15088,N_14303,N_14879);
xor U15089 (N_15089,N_11207,N_14548);
and U15090 (N_15090,N_11172,N_14861);
or U15091 (N_15091,N_14814,N_10817);
nand U15092 (N_15092,N_12311,N_11665);
nor U15093 (N_15093,N_11607,N_13481);
nor U15094 (N_15094,N_11212,N_12213);
nor U15095 (N_15095,N_10774,N_13741);
nand U15096 (N_15096,N_10485,N_12430);
nand U15097 (N_15097,N_10616,N_11114);
or U15098 (N_15098,N_13917,N_10637);
xnor U15099 (N_15099,N_12251,N_12247);
or U15100 (N_15100,N_11515,N_14661);
and U15101 (N_15101,N_11486,N_10530);
and U15102 (N_15102,N_13440,N_12122);
and U15103 (N_15103,N_12910,N_11187);
or U15104 (N_15104,N_11329,N_13228);
and U15105 (N_15105,N_11767,N_10633);
and U15106 (N_15106,N_11267,N_10433);
nor U15107 (N_15107,N_14072,N_14483);
and U15108 (N_15108,N_10560,N_14485);
xnor U15109 (N_15109,N_10668,N_14905);
xnor U15110 (N_15110,N_11009,N_12338);
nor U15111 (N_15111,N_13249,N_12482);
xor U15112 (N_15112,N_13652,N_11919);
or U15113 (N_15113,N_13765,N_13276);
and U15114 (N_15114,N_10925,N_13791);
nor U15115 (N_15115,N_13444,N_10732);
nor U15116 (N_15116,N_13102,N_14866);
xnor U15117 (N_15117,N_11474,N_10992);
xnor U15118 (N_15118,N_12137,N_12867);
nand U15119 (N_15119,N_12541,N_12579);
xor U15120 (N_15120,N_11086,N_11951);
and U15121 (N_15121,N_13745,N_12301);
nand U15122 (N_15122,N_14479,N_10280);
or U15123 (N_15123,N_14591,N_13064);
xor U15124 (N_15124,N_14094,N_13829);
nor U15125 (N_15125,N_10728,N_10120);
and U15126 (N_15126,N_14495,N_10657);
xor U15127 (N_15127,N_10419,N_11161);
xor U15128 (N_15128,N_12386,N_13151);
xor U15129 (N_15129,N_13978,N_14456);
and U15130 (N_15130,N_12654,N_14707);
xnor U15131 (N_15131,N_14835,N_11862);
nand U15132 (N_15132,N_13729,N_13194);
or U15133 (N_15133,N_12971,N_14116);
nor U15134 (N_15134,N_10938,N_10714);
xnor U15135 (N_15135,N_14518,N_11110);
and U15136 (N_15136,N_11211,N_14939);
xnor U15137 (N_15137,N_12648,N_14986);
and U15138 (N_15138,N_13274,N_14837);
xnor U15139 (N_15139,N_12058,N_12084);
nand U15140 (N_15140,N_13783,N_11071);
nand U15141 (N_15141,N_14850,N_11657);
nor U15142 (N_15142,N_10448,N_10157);
and U15143 (N_15143,N_14940,N_14987);
and U15144 (N_15144,N_11117,N_11957);
and U15145 (N_15145,N_11888,N_14616);
nor U15146 (N_15146,N_14952,N_10792);
nand U15147 (N_15147,N_14252,N_14966);
nand U15148 (N_15148,N_11662,N_11264);
nand U15149 (N_15149,N_12820,N_10291);
or U15150 (N_15150,N_14267,N_10161);
nor U15151 (N_15151,N_14104,N_11558);
nor U15152 (N_15152,N_14600,N_13407);
nor U15153 (N_15153,N_13238,N_11350);
nor U15154 (N_15154,N_12161,N_10410);
and U15155 (N_15155,N_14481,N_13286);
xor U15156 (N_15156,N_11223,N_12329);
or U15157 (N_15157,N_14328,N_10617);
nand U15158 (N_15158,N_12824,N_14915);
nor U15159 (N_15159,N_12501,N_11194);
nor U15160 (N_15160,N_14098,N_10618);
nand U15161 (N_15161,N_14585,N_13933);
nand U15162 (N_15162,N_10282,N_13046);
nor U15163 (N_15163,N_10959,N_10756);
and U15164 (N_15164,N_12866,N_11220);
nand U15165 (N_15165,N_11468,N_10487);
and U15166 (N_15166,N_11518,N_13309);
nand U15167 (N_15167,N_14333,N_13807);
nor U15168 (N_15168,N_11709,N_10801);
nand U15169 (N_15169,N_10324,N_14997);
xnor U15170 (N_15170,N_10760,N_14683);
or U15171 (N_15171,N_14877,N_10486);
nand U15172 (N_15172,N_13212,N_11601);
nand U15173 (N_15173,N_14641,N_12916);
nand U15174 (N_15174,N_13441,N_11496);
xor U15175 (N_15175,N_12417,N_10206);
and U15176 (N_15176,N_13074,N_14882);
and U15177 (N_15177,N_11471,N_13546);
nor U15178 (N_15178,N_14774,N_10372);
nor U15179 (N_15179,N_14020,N_11490);
nand U15180 (N_15180,N_13131,N_14659);
nand U15181 (N_15181,N_14164,N_14753);
or U15182 (N_15182,N_13975,N_11538);
and U15183 (N_15183,N_11618,N_10155);
nand U15184 (N_15184,N_12879,N_12463);
and U15185 (N_15185,N_11053,N_13725);
nor U15186 (N_15186,N_13705,N_13338);
and U15187 (N_15187,N_12255,N_14461);
nand U15188 (N_15188,N_14957,N_10705);
and U15189 (N_15189,N_12473,N_11860);
or U15190 (N_15190,N_10869,N_13121);
xor U15191 (N_15191,N_12167,N_13801);
nor U15192 (N_15192,N_12499,N_12160);
or U15193 (N_15193,N_14896,N_10555);
nand U15194 (N_15194,N_13278,N_11313);
nor U15195 (N_15195,N_14484,N_13498);
nor U15196 (N_15196,N_10634,N_12062);
or U15197 (N_15197,N_14414,N_13426);
nor U15198 (N_15198,N_13204,N_14192);
nand U15199 (N_15199,N_11384,N_13491);
xnor U15200 (N_15200,N_14764,N_11611);
nor U15201 (N_15201,N_10824,N_10207);
xnor U15202 (N_15202,N_11362,N_14550);
nand U15203 (N_15203,N_12896,N_11251);
and U15204 (N_15204,N_12583,N_11370);
nand U15205 (N_15205,N_14734,N_12872);
and U15206 (N_15206,N_12569,N_14384);
xnor U15207 (N_15207,N_10584,N_14913);
xnor U15208 (N_15208,N_11333,N_14993);
and U15209 (N_15209,N_10136,N_13699);
xor U15210 (N_15210,N_13193,N_10866);
nor U15211 (N_15211,N_10997,N_13580);
nand U15212 (N_15212,N_14933,N_13944);
or U15213 (N_15213,N_10987,N_10472);
or U15214 (N_15214,N_11300,N_14667);
xnor U15215 (N_15215,N_14489,N_11499);
nor U15216 (N_15216,N_14097,N_10216);
and U15217 (N_15217,N_13717,N_11978);
and U15218 (N_15218,N_10457,N_10802);
or U15219 (N_15219,N_10056,N_14640);
xnor U15220 (N_15220,N_12745,N_12731);
or U15221 (N_15221,N_13614,N_13341);
nand U15222 (N_15222,N_13726,N_12453);
or U15223 (N_15223,N_10495,N_12533);
xnor U15224 (N_15224,N_12447,N_10462);
nor U15225 (N_15225,N_10043,N_14441);
nor U15226 (N_15226,N_12037,N_14371);
xnor U15227 (N_15227,N_11045,N_11853);
nor U15228 (N_15228,N_11507,N_11173);
nor U15229 (N_15229,N_12165,N_11120);
xnor U15230 (N_15230,N_11203,N_13241);
nor U15231 (N_15231,N_12297,N_13357);
and U15232 (N_15232,N_12152,N_12182);
xnor U15233 (N_15233,N_12973,N_14676);
nand U15234 (N_15234,N_13127,N_13130);
or U15235 (N_15235,N_11361,N_13996);
and U15236 (N_15236,N_11376,N_12408);
nor U15237 (N_15237,N_12056,N_14729);
nand U15238 (N_15238,N_10880,N_13335);
nand U15239 (N_15239,N_12668,N_14399);
nor U15240 (N_15240,N_13583,N_10960);
nand U15241 (N_15241,N_11367,N_13720);
nor U15242 (N_15242,N_10272,N_13227);
or U15243 (N_15243,N_14395,N_13409);
nor U15244 (N_15244,N_10420,N_13157);
nor U15245 (N_15245,N_13520,N_11307);
nand U15246 (N_15246,N_10083,N_12966);
or U15247 (N_15247,N_12346,N_13125);
or U15248 (N_15248,N_10827,N_14106);
xor U15249 (N_15249,N_11961,N_11882);
and U15250 (N_15250,N_14705,N_14423);
or U15251 (N_15251,N_14300,N_13708);
and U15252 (N_15252,N_11510,N_14234);
and U15253 (N_15253,N_13758,N_13019);
xnor U15254 (N_15254,N_11438,N_13697);
nand U15255 (N_15255,N_14951,N_14124);
and U15256 (N_15256,N_11210,N_13352);
or U15257 (N_15257,N_13458,N_12018);
xor U15258 (N_15258,N_10830,N_12407);
and U15259 (N_15259,N_14989,N_12324);
xnor U15260 (N_15260,N_13818,N_13464);
xnor U15261 (N_15261,N_10384,N_13921);
or U15262 (N_15262,N_10121,N_12197);
and U15263 (N_15263,N_14457,N_12042);
or U15264 (N_15264,N_11273,N_14128);
or U15265 (N_15265,N_14179,N_13684);
nor U15266 (N_15266,N_10542,N_10076);
and U15267 (N_15267,N_10261,N_10733);
xor U15268 (N_15268,N_11638,N_12738);
and U15269 (N_15269,N_13026,N_14271);
nand U15270 (N_15270,N_11854,N_13898);
nor U15271 (N_15271,N_14108,N_14261);
or U15272 (N_15272,N_11795,N_14779);
and U15273 (N_15273,N_14467,N_13840);
nor U15274 (N_15274,N_13925,N_11498);
nand U15275 (N_15275,N_13468,N_12853);
xor U15276 (N_15276,N_11345,N_14684);
or U15277 (N_15277,N_13993,N_12667);
nand U15278 (N_15278,N_11106,N_14273);
nand U15279 (N_15279,N_11785,N_11419);
xnor U15280 (N_15280,N_13318,N_12315);
nand U15281 (N_15281,N_13218,N_10711);
nor U15282 (N_15282,N_10820,N_14846);
xor U15283 (N_15283,N_13012,N_10323);
or U15284 (N_15284,N_11332,N_14469);
nor U15285 (N_15285,N_11561,N_12674);
and U15286 (N_15286,N_13154,N_12146);
xor U15287 (N_15287,N_14438,N_13501);
xnor U15288 (N_15288,N_11016,N_12722);
xor U15289 (N_15289,N_11732,N_11883);
nand U15290 (N_15290,N_12723,N_14549);
and U15291 (N_15291,N_13532,N_12815);
or U15292 (N_15292,N_14426,N_12168);
nor U15293 (N_15293,N_14722,N_14034);
or U15294 (N_15294,N_14785,N_12227);
nor U15295 (N_15295,N_10832,N_10305);
nor U15296 (N_15296,N_10019,N_11998);
nand U15297 (N_15297,N_13054,N_13346);
nor U15298 (N_15298,N_12865,N_12003);
or U15299 (N_15299,N_13812,N_14322);
nand U15300 (N_15300,N_12323,N_13881);
nand U15301 (N_15301,N_11091,N_12553);
nand U15302 (N_15302,N_12841,N_11397);
nand U15303 (N_15303,N_13786,N_10009);
and U15304 (N_15304,N_11278,N_13764);
xnor U15305 (N_15305,N_13264,N_14150);
nor U15306 (N_15306,N_13727,N_13557);
nand U15307 (N_15307,N_14397,N_13316);
nand U15308 (N_15308,N_14947,N_10748);
nor U15309 (N_15309,N_11060,N_10684);
and U15310 (N_15310,N_10563,N_14567);
nor U15311 (N_15311,N_12871,N_10971);
nand U15312 (N_15312,N_10332,N_10370);
nor U15313 (N_15313,N_14387,N_11427);
and U15314 (N_15314,N_12117,N_12262);
nor U15315 (N_15315,N_10187,N_10726);
or U15316 (N_15316,N_14324,N_13155);
and U15317 (N_15317,N_13522,N_11651);
and U15318 (N_15318,N_11409,N_11437);
or U15319 (N_15319,N_10040,N_12334);
xnor U15320 (N_15320,N_11064,N_13478);
and U15321 (N_15321,N_10177,N_11886);
and U15322 (N_15322,N_10054,N_12012);
and U15323 (N_15323,N_11887,N_13382);
nand U15324 (N_15324,N_13117,N_10226);
xnor U15325 (N_15325,N_11355,N_14162);
or U15326 (N_15326,N_14583,N_13808);
and U15327 (N_15327,N_14242,N_12748);
or U15328 (N_15328,N_13677,N_12376);
nor U15329 (N_15329,N_13998,N_14325);
nor U15330 (N_15330,N_11577,N_14513);
nor U15331 (N_15331,N_14208,N_11390);
xnor U15332 (N_15332,N_13446,N_12783);
or U15333 (N_15333,N_14326,N_10180);
nor U15334 (N_15334,N_13827,N_14768);
nand U15335 (N_15335,N_11279,N_10321);
or U15336 (N_15336,N_13475,N_10425);
nor U15337 (N_15337,N_12318,N_13326);
nor U15338 (N_15338,N_11988,N_12809);
nor U15339 (N_15339,N_13836,N_11542);
and U15340 (N_15340,N_12468,N_10051);
xnor U15341 (N_15341,N_13149,N_14436);
xnor U15342 (N_15342,N_10529,N_10704);
xnor U15343 (N_15343,N_14372,N_14392);
xnor U15344 (N_15344,N_14059,N_10309);
nor U15345 (N_15345,N_10796,N_14664);
nand U15346 (N_15346,N_11516,N_14040);
or U15347 (N_15347,N_11290,N_12229);
nor U15348 (N_15348,N_14043,N_13108);
and U15349 (N_15349,N_11007,N_13083);
and U15350 (N_15350,N_11160,N_12036);
nand U15351 (N_15351,N_11238,N_14375);
or U15352 (N_15352,N_11129,N_10809);
xor U15353 (N_15353,N_13240,N_14201);
or U15354 (N_15354,N_10493,N_12063);
or U15355 (N_15355,N_10843,N_10349);
nor U15356 (N_15356,N_10185,N_12006);
nand U15357 (N_15357,N_12230,N_14736);
and U15358 (N_15358,N_13550,N_12775);
nor U15359 (N_15359,N_11403,N_13771);
or U15360 (N_15360,N_11097,N_14396);
nor U15361 (N_15361,N_12972,N_11572);
nand U15362 (N_15362,N_11915,N_13500);
or U15363 (N_15363,N_14929,N_10856);
xnor U15364 (N_15364,N_12626,N_12921);
nor U15365 (N_15365,N_14749,N_12026);
nand U15366 (N_15366,N_12732,N_11365);
nand U15367 (N_15367,N_11293,N_11426);
nand U15368 (N_15368,N_10652,N_12500);
nor U15369 (N_15369,N_13740,N_13584);
or U15370 (N_15370,N_12127,N_12942);
nand U15371 (N_15371,N_10229,N_12708);
and U15372 (N_15372,N_13502,N_10199);
nor U15373 (N_15373,N_10984,N_11485);
xor U15374 (N_15374,N_13884,N_10779);
nor U15375 (N_15375,N_12620,N_14251);
or U15376 (N_15376,N_13400,N_10787);
or U15377 (N_15377,N_13160,N_14780);
nor U15378 (N_15378,N_14807,N_13627);
xnor U15379 (N_15379,N_10287,N_14649);
nor U15380 (N_15380,N_13695,N_14781);
and U15381 (N_15381,N_14892,N_12939);
and U15382 (N_15382,N_12678,N_11476);
nor U15383 (N_15383,N_12634,N_11694);
nor U15384 (N_15384,N_10769,N_10628);
and U15385 (N_15385,N_11412,N_13516);
and U15386 (N_15386,N_10452,N_14203);
nand U15387 (N_15387,N_14792,N_13182);
nand U15388 (N_15388,N_14697,N_12600);
nand U15389 (N_15389,N_14932,N_10016);
nand U15390 (N_15390,N_11840,N_11484);
and U15391 (N_15391,N_11768,N_13270);
xor U15392 (N_15392,N_12391,N_10639);
and U15393 (N_15393,N_10889,N_10583);
xnor U15394 (N_15394,N_10067,N_12110);
xor U15395 (N_15395,N_13476,N_11813);
or U15396 (N_15396,N_14474,N_11371);
and U15397 (N_15397,N_10114,N_13578);
or U15398 (N_15398,N_11514,N_12039);
or U15399 (N_15399,N_13366,N_12250);
nor U15400 (N_15400,N_10515,N_10148);
and U15401 (N_15401,N_12253,N_10265);
xor U15402 (N_15402,N_12799,N_12098);
xor U15403 (N_15403,N_13126,N_12749);
or U15404 (N_15404,N_14956,N_11015);
nand U15405 (N_15405,N_10597,N_12325);
or U15406 (N_15406,N_10179,N_11924);
nor U15407 (N_15407,N_10979,N_13559);
nor U15408 (N_15408,N_12204,N_11841);
nor U15409 (N_15409,N_10643,N_14775);
and U15410 (N_15410,N_13585,N_12598);
or U15411 (N_15411,N_11557,N_11206);
or U15412 (N_15412,N_11686,N_13200);
or U15413 (N_15413,N_13041,N_11029);
or U15414 (N_15414,N_12631,N_14712);
or U15415 (N_15415,N_13215,N_10808);
nand U15416 (N_15416,N_12969,N_10899);
nor U15417 (N_15417,N_14595,N_12434);
nor U15418 (N_15418,N_13243,N_12739);
or U15419 (N_15419,N_12028,N_12317);
and U15420 (N_15420,N_11353,N_13865);
xor U15421 (N_15421,N_12358,N_10218);
xnor U15422 (N_15422,N_10195,N_11575);
nand U15423 (N_15423,N_11553,N_14727);
and U15424 (N_15424,N_10608,N_12140);
nand U15425 (N_15425,N_13899,N_10708);
xnor U15426 (N_15426,N_13549,N_10197);
or U15427 (N_15427,N_11632,N_10651);
and U15428 (N_15428,N_10154,N_11955);
nor U15429 (N_15429,N_11822,N_11481);
nor U15430 (N_15430,N_14902,N_10262);
nand U15431 (N_15431,N_10205,N_14570);
or U15432 (N_15432,N_11631,N_13308);
nand U15433 (N_15433,N_11900,N_10192);
and U15434 (N_15434,N_10838,N_12478);
nor U15435 (N_15435,N_10319,N_12503);
and U15436 (N_15436,N_10296,N_14965);
xnor U15437 (N_15437,N_11327,N_10847);
or U15438 (N_15438,N_12170,N_11268);
and U15439 (N_15439,N_14158,N_11261);
and U15440 (N_15440,N_12529,N_12145);
nand U15441 (N_15441,N_12616,N_10303);
nand U15442 (N_15442,N_12907,N_13139);
or U15443 (N_15443,N_10193,N_13010);
and U15444 (N_15444,N_12548,N_14972);
xor U15445 (N_15445,N_12491,N_12770);
and U15446 (N_15446,N_14967,N_11150);
and U15447 (N_15447,N_12065,N_14047);
xor U15448 (N_15448,N_11197,N_11044);
and U15449 (N_15449,N_12420,N_12106);
nor U15450 (N_15450,N_13882,N_11950);
or U15451 (N_15451,N_14916,N_12021);
nand U15452 (N_15452,N_10859,N_13329);
or U15453 (N_15453,N_11151,N_12377);
xnor U15454 (N_15454,N_12339,N_10508);
or U15455 (N_15455,N_10675,N_11221);
and U15456 (N_15456,N_12396,N_11942);
xnor U15457 (N_15457,N_12509,N_12153);
or U15458 (N_15458,N_14874,N_11556);
nor U15459 (N_15459,N_14368,N_13534);
or U15460 (N_15460,N_13843,N_13109);
or U15461 (N_15461,N_12245,N_13183);
or U15462 (N_15462,N_14083,N_10867);
xor U15463 (N_15463,N_11454,N_13360);
nor U15464 (N_15464,N_10175,N_13814);
xor U15465 (N_15465,N_14571,N_14769);
or U15466 (N_15466,N_14238,N_10554);
nand U15467 (N_15467,N_14710,N_14257);
nor U15468 (N_15468,N_13872,N_13721);
and U15469 (N_15469,N_14065,N_13613);
and U15470 (N_15470,N_12064,N_12260);
and U15471 (N_15471,N_13061,N_11737);
xor U15472 (N_15472,N_13832,N_11296);
xor U15473 (N_15473,N_13620,N_12873);
nor U15474 (N_15474,N_10887,N_12038);
nor U15475 (N_15475,N_14575,N_14112);
nor U15476 (N_15476,N_12979,N_10517);
and U15477 (N_15477,N_12638,N_13178);
nor U15478 (N_15478,N_11535,N_10833);
xor U15479 (N_15479,N_12228,N_12628);
nor U15480 (N_15480,N_14783,N_10383);
and U15481 (N_15481,N_14134,N_13878);
or U15482 (N_15482,N_14895,N_10596);
nor U15483 (N_15483,N_12926,N_14464);
nor U15484 (N_15484,N_10213,N_12082);
xor U15485 (N_15485,N_13803,N_11435);
xnor U15486 (N_15486,N_12225,N_13903);
xnor U15487 (N_15487,N_14239,N_10547);
xnor U15488 (N_15488,N_14863,N_13486);
nor U15489 (N_15489,N_12151,N_10813);
nor U15490 (N_15490,N_10945,N_10535);
or U15491 (N_15491,N_14638,N_11788);
or U15492 (N_15492,N_12193,N_14307);
nand U15493 (N_15493,N_11823,N_10772);
and U15494 (N_15494,N_11772,N_10638);
and U15495 (N_15495,N_13556,N_10663);
nand U15496 (N_15496,N_10113,N_13566);
nor U15497 (N_15497,N_14284,N_14750);
or U15498 (N_15498,N_11047,N_10721);
nand U15499 (N_15499,N_14602,N_13187);
and U15500 (N_15500,N_14084,N_13573);
nand U15501 (N_15501,N_11241,N_14429);
or U15502 (N_15502,N_13219,N_13391);
nor U15503 (N_15503,N_13624,N_12404);
or U15504 (N_15504,N_12800,N_13135);
nand U15505 (N_15505,N_13298,N_13625);
xor U15506 (N_15506,N_11147,N_10397);
and U15507 (N_15507,N_14144,N_12068);
nor U15508 (N_15508,N_11041,N_14016);
xnor U15509 (N_15509,N_14716,N_12271);
or U15510 (N_15510,N_10137,N_13222);
and U15511 (N_15511,N_10759,N_10334);
xnor U15512 (N_15512,N_13645,N_13088);
nor U15513 (N_15513,N_12461,N_11794);
nand U15514 (N_15514,N_12443,N_12107);
or U15515 (N_15515,N_13632,N_12378);
nand U15516 (N_15516,N_11877,N_11980);
and U15517 (N_15517,N_11928,N_14578);
nor U15518 (N_15518,N_13958,N_13617);
and U15519 (N_15519,N_11380,N_14632);
and U15520 (N_15520,N_14295,N_10480);
nor U15521 (N_15521,N_11844,N_12950);
and U15522 (N_15522,N_11171,N_13604);
and U15523 (N_15523,N_14416,N_10605);
nor U15524 (N_15524,N_12448,N_13422);
xor U15525 (N_15525,N_10128,N_13769);
nor U15526 (N_15526,N_10146,N_14816);
nor U15527 (N_15527,N_13071,N_11655);
xnor U15528 (N_15528,N_10698,N_14378);
xnor U15529 (N_15529,N_13579,N_14671);
nand U15530 (N_15530,N_13715,N_12522);
xor U15531 (N_15531,N_14884,N_12415);
nand U15532 (N_15532,N_14081,N_13377);
nor U15533 (N_15533,N_10249,N_12736);
or U15534 (N_15534,N_10233,N_10574);
nor U15535 (N_15535,N_10174,N_12832);
xnor U15536 (N_15536,N_12205,N_10527);
nand U15537 (N_15537,N_12265,N_11817);
nor U15538 (N_15538,N_14751,N_10473);
nor U15539 (N_15539,N_13761,N_14903);
or U15540 (N_15540,N_13140,N_11994);
nor U15541 (N_15541,N_11982,N_13211);
nand U15542 (N_15542,N_11292,N_13082);
nor U15543 (N_15543,N_10888,N_10791);
and U15544 (N_15544,N_14056,N_13800);
xor U15545 (N_15545,N_12998,N_13355);
xor U15546 (N_15546,N_11080,N_12517);
nand U15547 (N_15547,N_11299,N_11195);
nor U15548 (N_15548,N_12844,N_13959);
xor U15549 (N_15549,N_13641,N_10230);
and U15550 (N_15550,N_11948,N_12008);
nor U15551 (N_15551,N_12915,N_10680);
xor U15552 (N_15552,N_10752,N_12949);
nor U15553 (N_15553,N_12001,N_11581);
nor U15554 (N_15554,N_13749,N_10635);
xor U15555 (N_15555,N_10528,N_11081);
nand U15556 (N_15556,N_12814,N_14596);
xnor U15557 (N_15557,N_12292,N_10520);
and U15558 (N_15558,N_14017,N_11089);
and U15559 (N_15559,N_11265,N_12080);
or U15560 (N_15560,N_11479,N_11399);
or U15561 (N_15561,N_14698,N_10418);
nand U15562 (N_15562,N_13972,N_12774);
or U15563 (N_15563,N_13577,N_11020);
nor U15564 (N_15564,N_14505,N_11494);
xor U15565 (N_15565,N_14470,N_14867);
xor U15566 (N_15566,N_10990,N_14443);
nand U15567 (N_15567,N_11635,N_10660);
and U15568 (N_15568,N_14644,N_11640);
xnor U15569 (N_15569,N_12073,N_13531);
nand U15570 (N_15570,N_14114,N_11964);
xnor U15571 (N_15571,N_10129,N_12696);
and U15572 (N_15572,N_13159,N_11589);
and U15573 (N_15573,N_11578,N_12050);
xnor U15574 (N_15574,N_14213,N_11720);
xor U15575 (N_15575,N_13447,N_12790);
xnor U15576 (N_15576,N_13053,N_14919);
xnor U15577 (N_15577,N_10928,N_13951);
xor U15578 (N_15578,N_10408,N_14421);
xnor U15579 (N_15579,N_11132,N_11179);
and U15580 (N_15580,N_11425,N_12007);
xnor U15581 (N_15581,N_12201,N_13128);
nand U15582 (N_15582,N_10119,N_10696);
nor U15583 (N_15583,N_14336,N_10359);
xor U15584 (N_15584,N_11714,N_13977);
and U15585 (N_15585,N_14878,N_13861);
and U15586 (N_15586,N_14717,N_14844);
and U15587 (N_15587,N_11612,N_13784);
xor U15588 (N_15588,N_13646,N_14431);
and U15589 (N_15589,N_12908,N_12164);
nand U15590 (N_15590,N_10037,N_11528);
or U15591 (N_15591,N_10922,N_12675);
nand U15592 (N_15592,N_13626,N_14459);
and U15593 (N_15593,N_13463,N_14250);
nor U15594 (N_15594,N_12787,N_11930);
nand U15595 (N_15595,N_13428,N_11291);
nor U15596 (N_15596,N_13505,N_14864);
and U15597 (N_15597,N_11028,N_10723);
nand U15598 (N_15598,N_11158,N_13058);
xor U15599 (N_15599,N_10276,N_11843);
nand U15600 (N_15600,N_10565,N_11348);
nand U15601 (N_15601,N_11135,N_11962);
nand U15602 (N_15602,N_11755,N_14747);
xnor U15603 (N_15603,N_12937,N_10736);
and U15604 (N_15604,N_13924,N_11670);
or U15605 (N_15605,N_10818,N_13226);
nand U15606 (N_15606,N_10133,N_14521);
and U15607 (N_15607,N_14102,N_14499);
nand U15608 (N_15608,N_13509,N_14642);
nor U15609 (N_15609,N_10564,N_11146);
xnor U15610 (N_15610,N_11275,N_11431);
and U15611 (N_15611,N_10379,N_11074);
nand U15612 (N_15612,N_14169,N_12746);
nor U15613 (N_15613,N_11923,N_13982);
nand U15614 (N_15614,N_14885,N_12539);
and U15615 (N_15615,N_14822,N_12679);
or U15616 (N_15616,N_13858,N_12554);
nor U15617 (N_15617,N_13886,N_14287);
xnor U15618 (N_15618,N_11855,N_14028);
or U15619 (N_15619,N_13987,N_12763);
nor U15620 (N_15620,N_10151,N_11826);
nor U15621 (N_15621,N_14292,N_12957);
xnor U15622 (N_15622,N_11396,N_13916);
xor U15623 (N_15623,N_14062,N_14331);
xor U15624 (N_15624,N_11692,N_10620);
nor U15625 (N_15625,N_10426,N_13528);
nand U15626 (N_15626,N_13220,N_12768);
nor U15627 (N_15627,N_14757,N_13063);
nand U15628 (N_15628,N_14374,N_13392);
nand U15629 (N_15629,N_14354,N_12901);
or U15630 (N_15630,N_14579,N_11597);
nand U15631 (N_15631,N_13885,N_12072);
xor U15632 (N_15632,N_12411,N_14693);
nand U15633 (N_15633,N_14954,N_13036);
or U15634 (N_15634,N_10488,N_12802);
and U15635 (N_15635,N_14831,N_11311);
xor U15636 (N_15636,N_14334,N_10604);
nand U15637 (N_15637,N_13039,N_14893);
nor U15638 (N_15638,N_14995,N_12066);
nor U15639 (N_15639,N_13539,N_11554);
nand U15640 (N_15640,N_10855,N_12573);
nor U15641 (N_15641,N_13195,N_13177);
nand U15642 (N_15642,N_13794,N_14085);
and U15643 (N_15643,N_12835,N_11598);
nand U15644 (N_15644,N_10568,N_14146);
or U15645 (N_15645,N_14634,N_10252);
nand U15646 (N_15646,N_13045,N_13590);
xnor U15647 (N_15647,N_10719,N_11660);
nand U15648 (N_15648,N_14532,N_12266);
xnor U15649 (N_15649,N_10735,N_12727);
nor U15650 (N_15650,N_13913,N_10613);
nand U15651 (N_15651,N_12485,N_12067);
nor U15652 (N_15652,N_10250,N_11918);
nor U15653 (N_15653,N_11866,N_13804);
and U15654 (N_15654,N_13817,N_14928);
or U15655 (N_15655,N_14612,N_14361);
nor U15656 (N_15656,N_11615,N_10245);
nand U15657 (N_15657,N_10961,N_12948);
nand U15658 (N_15658,N_10156,N_11401);
and U15659 (N_15659,N_10006,N_12629);
or U15660 (N_15660,N_10913,N_14135);
and U15661 (N_15661,N_14796,N_10377);
nor U15662 (N_15662,N_11155,N_14976);
nand U15663 (N_15663,N_11931,N_13162);
nand U15664 (N_15664,N_14451,N_13438);
or U15665 (N_15665,N_10561,N_13024);
nand U15666 (N_15666,N_14581,N_12034);
nor U15667 (N_15667,N_12624,N_13448);
xor U15668 (N_15668,N_13405,N_12904);
and U15669 (N_15669,N_12258,N_14935);
or U15670 (N_15670,N_13621,N_13545);
or U15671 (N_15671,N_12534,N_12511);
and U15672 (N_15672,N_10689,N_10524);
xnor U15673 (N_15673,N_11905,N_13343);
xnor U15674 (N_15674,N_11934,N_14022);
and U15675 (N_15675,N_13815,N_11722);
or U15676 (N_15676,N_14025,N_13388);
and U15677 (N_15677,N_10002,N_11682);
and U15678 (N_15678,N_14131,N_10882);
nor U15679 (N_15679,N_14155,N_11819);
nor U15680 (N_15680,N_11775,N_14068);
and U15681 (N_15681,N_11517,N_13795);
nor U15682 (N_15682,N_12687,N_14811);
or U15683 (N_15683,N_11341,N_14260);
nor U15684 (N_15684,N_11324,N_14560);
nor U15685 (N_15685,N_10118,N_10717);
nor U15686 (N_15686,N_11018,N_14147);
or U15687 (N_15687,N_14924,N_10687);
or U15688 (N_15688,N_10227,N_12162);
nand U15689 (N_15689,N_11216,N_10371);
or U15690 (N_15690,N_12069,N_12196);
and U15691 (N_15691,N_14592,N_10466);
nand U15692 (N_15692,N_14569,N_12221);
nand U15693 (N_15693,N_14115,N_13868);
nor U15694 (N_15694,N_13198,N_11878);
and U15695 (N_15695,N_13709,N_14174);
nand U15696 (N_15696,N_14344,N_12296);
or U15697 (N_15697,N_13537,N_14272);
nand U15698 (N_15698,N_11006,N_10918);
or U15699 (N_15699,N_11815,N_11723);
or U15700 (N_15700,N_13348,N_11017);
xnor U15701 (N_15701,N_13206,N_10800);
nor U15702 (N_15702,N_10621,N_13939);
nor U15703 (N_15703,N_12195,N_10650);
nand U15704 (N_15704,N_13544,N_11449);
and U15705 (N_15705,N_13555,N_10980);
nor U15706 (N_15706,N_12451,N_12640);
nand U15707 (N_15707,N_13176,N_14444);
xor U15708 (N_15708,N_13920,N_10525);
and U15709 (N_15709,N_14278,N_10642);
nand U15710 (N_15710,N_12740,N_12612);
and U15711 (N_15711,N_11154,N_11392);
and U15712 (N_15712,N_13056,N_12041);
xnor U15713 (N_15713,N_12493,N_13390);
and U15714 (N_15714,N_11317,N_10963);
and U15715 (N_15715,N_10729,N_11688);
or U15716 (N_15716,N_10715,N_11895);
nand U15717 (N_15717,N_14502,N_14604);
or U15718 (N_15718,N_13842,N_10944);
nand U15719 (N_15719,N_13575,N_12233);
xnor U15720 (N_15720,N_13770,N_13828);
or U15721 (N_15721,N_13994,N_12498);
xnor U15722 (N_15722,N_10238,N_13028);
and U15723 (N_15723,N_11552,N_11500);
nor U15724 (N_15724,N_13548,N_13322);
nor U15725 (N_15725,N_12103,N_14341);
nand U15726 (N_15726,N_13297,N_14551);
and U15727 (N_15727,N_10412,N_10626);
nor U15728 (N_15728,N_11547,N_12968);
and U15729 (N_15729,N_10586,N_13989);
nor U15730 (N_15730,N_11508,N_12595);
nor U15731 (N_15731,N_12239,N_14576);
and U15732 (N_15732,N_11058,N_13013);
nand U15733 (N_15733,N_11033,N_13313);
xnor U15734 (N_15734,N_12608,N_10876);
nand U15735 (N_15735,N_14911,N_13805);
nand U15736 (N_15736,N_11659,N_11320);
nor U15737 (N_15737,N_12856,N_10263);
nand U15738 (N_15738,N_11712,N_14763);
or U15739 (N_15739,N_12840,N_10405);
or U15740 (N_15740,N_11463,N_13253);
nor U15741 (N_15741,N_10267,N_13239);
xor U15742 (N_15742,N_14172,N_13090);
nand U15743 (N_15743,N_13506,N_10674);
and U15744 (N_15744,N_10911,N_10017);
and U15745 (N_15745,N_13158,N_11927);
and U15746 (N_15746,N_12538,N_13014);
nand U15747 (N_15747,N_12020,N_14733);
xor U15748 (N_15748,N_12752,N_13303);
or U15749 (N_15749,N_14161,N_12693);
and U15750 (N_15750,N_11138,N_14448);
or U15751 (N_15751,N_14759,N_13331);
xor U15752 (N_15752,N_11461,N_10898);
or U15753 (N_15753,N_13619,N_14142);
or U15754 (N_15754,N_13433,N_14803);
nand U15755 (N_15755,N_13831,N_13290);
or U15756 (N_15756,N_12633,N_13395);
or U15757 (N_15757,N_14335,N_13874);
and U15758 (N_15758,N_13928,N_10483);
nor U15759 (N_15759,N_12970,N_10743);
or U15760 (N_15760,N_11691,N_10516);
and U15761 (N_15761,N_14620,N_13582);
and U15762 (N_15762,N_10754,N_14925);
and U15763 (N_15763,N_11909,N_10169);
or U15764 (N_15764,N_10678,N_14855);
xnor U15765 (N_15765,N_12766,N_14478);
or U15766 (N_15766,N_14681,N_11492);
and U15767 (N_15767,N_14180,N_14566);
and U15768 (N_15768,N_14870,N_14332);
xnor U15769 (N_15769,N_12349,N_13615);
or U15770 (N_15770,N_10429,N_11733);
nor U15771 (N_15771,N_10088,N_13603);
nand U15772 (N_15772,N_14523,N_11740);
and U15773 (N_15773,N_11894,N_11989);
and U15774 (N_15774,N_10612,N_10308);
nand U15775 (N_15775,N_11868,N_14206);
or U15776 (N_15776,N_10060,N_14342);
and U15777 (N_15777,N_11266,N_13678);
and U15778 (N_15778,N_11675,N_10346);
nand U15779 (N_15779,N_11102,N_13970);
nor U15780 (N_15780,N_12355,N_11991);
nor U15781 (N_15781,N_14968,N_13034);
nor U15782 (N_15782,N_12584,N_10318);
and U15783 (N_15783,N_14391,N_13260);
xnor U15784 (N_15784,N_12207,N_11683);
xnor U15785 (N_15785,N_14105,N_11012);
or U15786 (N_15786,N_13487,N_13314);
or U15787 (N_15787,N_11448,N_12326);
nand U15788 (N_15788,N_14946,N_11676);
and U15789 (N_15789,N_11019,N_13207);
xor U15790 (N_15790,N_11055,N_12057);
and U15791 (N_15791,N_13022,N_11776);
xnor U15792 (N_15792,N_13702,N_11935);
xnor U15793 (N_15793,N_12997,N_13373);
or U15794 (N_15794,N_13425,N_10921);
and U15795 (N_15795,N_13594,N_11550);
xor U15796 (N_15796,N_14854,N_10531);
nand U15797 (N_15797,N_12779,N_10374);
xor U15798 (N_15798,N_13541,N_12471);
and U15799 (N_15799,N_10697,N_10703);
xor U15800 (N_15800,N_14011,N_14510);
xor U15801 (N_15801,N_14691,N_13662);
and U15802 (N_15802,N_11139,N_12043);
or U15803 (N_15803,N_10012,N_10450);
xnor U15804 (N_15804,N_11407,N_13859);
or U15805 (N_15805,N_10422,N_10923);
nand U15806 (N_15806,N_10077,N_11576);
xor U15807 (N_15807,N_12724,N_11690);
nor U15808 (N_15808,N_13016,N_12278);
and U15809 (N_15809,N_13097,N_14433);
xnor U15810 (N_15810,N_12203,N_10166);
nand U15811 (N_15811,N_14036,N_10367);
and U15812 (N_15812,N_14839,N_10901);
xor U15813 (N_15813,N_11828,N_13340);
nor U15814 (N_15814,N_10393,N_10283);
nand U15815 (N_15815,N_12665,N_13760);
and U15816 (N_15816,N_14291,N_12480);
or U15817 (N_15817,N_13894,N_14794);
nand U15818 (N_15818,N_10631,N_11493);
or U15819 (N_15819,N_13350,N_13184);
or U15820 (N_15820,N_13837,N_10659);
xnor U15821 (N_15821,N_14711,N_10339);
or U15822 (N_15822,N_12010,N_10790);
xnor U15823 (N_15823,N_11594,N_13255);
nand U15824 (N_15824,N_14217,N_13250);
or U15825 (N_15825,N_11356,N_10846);
or U15826 (N_15826,N_11489,N_12422);
nand U15827 (N_15827,N_13597,N_11656);
nor U15828 (N_15828,N_11276,N_14245);
nor U15829 (N_15829,N_13766,N_11588);
nand U15830 (N_15830,N_11534,N_12615);
or U15831 (N_15831,N_13150,N_13423);
and U15832 (N_15832,N_13048,N_14538);
and U15833 (N_15833,N_10603,N_13320);
nand U15834 (N_15834,N_14214,N_12956);
nor U15835 (N_15835,N_14795,N_11075);
nand U15836 (N_15836,N_12914,N_10500);
nor U15837 (N_15837,N_13477,N_14229);
nor U15838 (N_15838,N_12818,N_12549);
or U15839 (N_15839,N_11548,N_11532);
nor U15840 (N_15840,N_12806,N_12644);
nand U15841 (N_15841,N_13706,N_10630);
or U15842 (N_15842,N_11123,N_14541);
nor U15843 (N_15843,N_11562,N_12053);
nand U15844 (N_15844,N_12294,N_12390);
and U15845 (N_15845,N_10976,N_14991);
nor U15846 (N_15846,N_10181,N_10079);
nand U15847 (N_15847,N_11283,N_14139);
or U15848 (N_15848,N_12495,N_14439);
nor U15849 (N_15849,N_12385,N_11717);
or U15850 (N_15850,N_12351,N_12677);
xnor U15851 (N_15851,N_11467,N_10686);
xor U15852 (N_15852,N_11124,N_12235);
xor U15853 (N_15853,N_13301,N_13330);
or U15854 (N_15854,N_14148,N_10214);
and U15855 (N_15855,N_12226,N_10929);
nand U15856 (N_15856,N_10361,N_10475);
nor U15857 (N_15857,N_13907,N_11626);
or U15858 (N_15858,N_14830,N_14730);
or U15859 (N_15859,N_10171,N_13875);
and U15860 (N_15860,N_11600,N_11642);
xor U15861 (N_15861,N_14064,N_11339);
nand U15862 (N_15862,N_10952,N_13156);
and U15863 (N_15863,N_10101,N_12094);
and U15864 (N_15864,N_10806,N_10805);
nor U15865 (N_15865,N_13864,N_13988);
nand U15866 (N_15866,N_10933,N_14367);
xnor U15867 (N_15867,N_10496,N_14808);
nand U15868 (N_15868,N_12150,N_11747);
or U15869 (N_15869,N_14657,N_12384);
nand U15870 (N_15870,N_13553,N_13668);
and U15871 (N_15871,N_11473,N_12218);
nor U15872 (N_15872,N_13623,N_13364);
and U15873 (N_15873,N_14133,N_13798);
xor U15874 (N_15874,N_12627,N_12530);
nand U15875 (N_15875,N_12771,N_13612);
and U15876 (N_15876,N_14437,N_10008);
xor U15877 (N_15877,N_13888,N_14618);
or U15878 (N_15878,N_12943,N_12044);
nor U15879 (N_15879,N_14655,N_14706);
nor U15880 (N_15880,N_12212,N_14556);
or U15881 (N_15881,N_14453,N_10795);
nor U15882 (N_15882,N_14921,N_10610);
or U15883 (N_15883,N_11972,N_13334);
xnor U15884 (N_15884,N_13246,N_10125);
nor U15885 (N_15885,N_11441,N_11130);
nand U15886 (N_15886,N_11766,N_12617);
xnor U15887 (N_15887,N_13421,N_13134);
nand U15888 (N_15888,N_12556,N_11297);
nand U15889 (N_15889,N_10839,N_10018);
or U15890 (N_15890,N_11873,N_12861);
nand U15891 (N_15891,N_12435,N_11804);
nand U15892 (N_15892,N_10579,N_12823);
xor U15893 (N_15893,N_11351,N_11447);
or U15894 (N_15894,N_14506,N_11121);
xor U15895 (N_15895,N_12526,N_10906);
xor U15896 (N_15896,N_10533,N_13530);
nor U15897 (N_15897,N_12348,N_10363);
or U15898 (N_15898,N_12313,N_12935);
nand U15899 (N_15899,N_14183,N_12156);
nand U15900 (N_15900,N_11809,N_13877);
or U15901 (N_15901,N_12630,N_11647);
and U15902 (N_15902,N_12328,N_14293);
xnor U15903 (N_15903,N_14547,N_14406);
and U15904 (N_15904,N_14086,N_10981);
nor U15905 (N_15905,N_14381,N_10821);
nand U15906 (N_15906,N_12208,N_11637);
nor U15907 (N_15907,N_14880,N_13911);
nor U15908 (N_15908,N_13547,N_14454);
xnor U15909 (N_15909,N_13474,N_12097);
and U15910 (N_15910,N_10082,N_11082);
xnor U15911 (N_15911,N_13332,N_13434);
and U15912 (N_15912,N_13739,N_10653);
xor U15913 (N_15913,N_13692,N_14611);
nand U15914 (N_15914,N_12876,N_11530);
nand U15915 (N_15915,N_13767,N_12298);
xor U15916 (N_15916,N_10835,N_12284);
nor U15917 (N_15917,N_13946,N_12424);
nand U15918 (N_15918,N_12414,N_14247);
xor U15919 (N_15919,N_14181,N_13830);
and U15920 (N_15920,N_12647,N_14848);
or U15921 (N_15921,N_13685,N_14403);
nor U15922 (N_15922,N_11803,N_12132);
and U15923 (N_15923,N_14353,N_10170);
and U15924 (N_15924,N_14868,N_14306);
nand U15925 (N_15925,N_14079,N_11242);
or U15926 (N_15926,N_10328,N_13512);
or U15927 (N_15927,N_12192,N_13658);
nand U15928 (N_15928,N_11710,N_13811);
and U15929 (N_15929,N_14961,N_11566);
or U15930 (N_15930,N_11037,N_13504);
nand U15931 (N_15931,N_14277,N_10957);
and U15932 (N_15932,N_10327,N_12959);
and U15933 (N_15933,N_12238,N_13406);
and U15934 (N_15934,N_11643,N_11801);
nor U15935 (N_15935,N_10036,N_10894);
xor U15936 (N_15936,N_11966,N_12852);
or U15937 (N_15937,N_12476,N_13781);
nor U15938 (N_15938,N_13923,N_12593);
nor U15939 (N_15939,N_11864,N_12683);
and U15940 (N_15940,N_12510,N_14832);
or U15941 (N_15941,N_11280,N_13595);
and U15942 (N_15942,N_14988,N_14009);
or U15943 (N_15943,N_10731,N_14624);
or U15944 (N_15944,N_10523,N_11088);
and U15945 (N_15945,N_11798,N_12821);
nand U15946 (N_15946,N_12184,N_13095);
xnor U15947 (N_15947,N_12543,N_14553);
or U15948 (N_15948,N_14498,N_14630);
nor U15949 (N_15949,N_10504,N_14357);
and U15950 (N_15950,N_13835,N_12520);
nand U15951 (N_15951,N_13465,N_11152);
xnor U15952 (N_15952,N_13608,N_12789);
nand U15953 (N_15953,N_13347,N_13363);
and U15954 (N_15954,N_12985,N_12354);
nand U15955 (N_15955,N_12709,N_11940);
nand U15956 (N_15956,N_14745,N_10666);
and U15957 (N_15957,N_14294,N_14847);
nor U15958 (N_15958,N_12905,N_10532);
nand U15959 (N_15959,N_11169,N_12685);
or U15960 (N_15960,N_14024,N_10456);
and U15961 (N_15961,N_10572,N_12402);
nand U15962 (N_15962,N_10546,N_11946);
xnor U15963 (N_15963,N_14752,N_12506);
xnor U15964 (N_15964,N_12356,N_10378);
and U15965 (N_15965,N_14365,N_14101);
and U15966 (N_15966,N_10373,N_13461);
or U15967 (N_15967,N_10004,N_10970);
xor U15968 (N_15968,N_11529,N_12409);
nand U15969 (N_15969,N_13640,N_11190);
xor U15970 (N_15970,N_11364,N_12179);
and U15971 (N_15971,N_13701,N_11459);
or U15972 (N_15972,N_14858,N_14650);
nor U15973 (N_15973,N_11751,N_12382);
xnor U15974 (N_15974,N_11176,N_14171);
nor U15975 (N_15975,N_12040,N_12114);
xor U15976 (N_15976,N_11729,N_10788);
or U15977 (N_15977,N_14674,N_10052);
xnor U15978 (N_15978,N_11830,N_14801);
nand U15979 (N_15979,N_11746,N_12481);
xor U15980 (N_15980,N_14977,N_14580);
nor U15981 (N_15981,N_10254,N_10699);
and U15982 (N_15982,N_10993,N_12883);
and U15983 (N_15983,N_13396,N_12075);
nor U15984 (N_15984,N_11469,N_10982);
nand U15985 (N_15985,N_12563,N_13105);
nand U15986 (N_15986,N_10093,N_12934);
and U15987 (N_15987,N_14643,N_11685);
nand U15988 (N_15988,N_14320,N_12552);
or U15989 (N_15989,N_10896,N_10988);
and U15990 (N_15990,N_14073,N_10489);
and U15991 (N_15991,N_11814,N_12686);
and U15992 (N_15992,N_11143,N_13999);
or U15993 (N_15993,N_14731,N_13107);
and U15994 (N_15994,N_14117,N_11165);
nor U15995 (N_15995,N_10186,N_14770);
or U15996 (N_15996,N_13637,N_14310);
nor U15997 (N_15997,N_11144,N_11116);
nor U15998 (N_15998,N_13321,N_14288);
xnor U15999 (N_15999,N_14672,N_11056);
xnor U16000 (N_16000,N_11752,N_14377);
or U16001 (N_16001,N_14964,N_13315);
and U16002 (N_16002,N_10958,N_13976);
and U16003 (N_16003,N_13572,N_11929);
nand U16004 (N_16004,N_13389,N_13523);
nor U16005 (N_16005,N_12256,N_13232);
or U16006 (N_16006,N_10279,N_12613);
nand U16007 (N_16007,N_10353,N_10571);
nor U16008 (N_16008,N_14748,N_11063);
xor U16009 (N_16009,N_10973,N_14737);
and U16010 (N_16010,N_13797,N_14363);
xnor U16011 (N_16011,N_14626,N_12660);
xnor U16012 (N_16012,N_11936,N_10766);
nor U16013 (N_16013,N_12932,N_14934);
nor U16014 (N_16014,N_10034,N_13483);
nor U16015 (N_16015,N_13981,N_10039);
nor U16016 (N_16016,N_14565,N_14125);
and U16017 (N_16017,N_13436,N_14301);
xnor U16018 (N_16018,N_14512,N_14744);
and U16019 (N_16019,N_11181,N_13605);
nor U16020 (N_16020,N_13170,N_13261);
or U16021 (N_16021,N_14389,N_12588);
xor U16022 (N_16022,N_12711,N_12717);
nor U16023 (N_16023,N_10601,N_14945);
nor U16024 (N_16024,N_13351,N_10068);
nor U16025 (N_16025,N_12138,N_10917);
or U16026 (N_16026,N_12525,N_14688);
or U16027 (N_16027,N_12889,N_10646);
or U16028 (N_16028,N_13554,N_11521);
or U16029 (N_16029,N_14345,N_10135);
or U16030 (N_16030,N_10541,N_12965);
and U16031 (N_16031,N_14601,N_10942);
xnor U16032 (N_16032,N_13292,N_13038);
and U16033 (N_16033,N_13380,N_13728);
and U16034 (N_16034,N_13995,N_11177);
and U16035 (N_16035,N_12248,N_13860);
nand U16036 (N_16036,N_14149,N_11893);
nor U16037 (N_16037,N_14207,N_13990);
nand U16038 (N_16038,N_12839,N_13763);
nor U16039 (N_16039,N_14833,N_12672);
nand U16040 (N_16040,N_12327,N_13536);
xor U16041 (N_16041,N_13023,N_14819);
nand U16042 (N_16042,N_13118,N_12341);
nand U16043 (N_16043,N_11472,N_10277);
or U16044 (N_16044,N_14076,N_12331);
and U16045 (N_16045,N_13636,N_12189);
and U16046 (N_16046,N_11100,N_12131);
nand U16047 (N_16047,N_10046,N_10061);
nand U16048 (N_16048,N_14198,N_14859);
or U16049 (N_16049,N_11702,N_10110);
or U16050 (N_16050,N_13420,N_11406);
nor U16051 (N_16051,N_11906,N_12183);
xnor U16052 (N_16052,N_11026,N_13793);
and U16053 (N_16053,N_10264,N_12211);
xor U16054 (N_16054,N_10602,N_10819);
and U16055 (N_16055,N_11824,N_11395);
nor U16056 (N_16056,N_12898,N_10127);
and U16057 (N_16057,N_13123,N_12088);
and U16058 (N_16058,N_10304,N_10310);
or U16059 (N_16059,N_14520,N_11475);
xor U16060 (N_16060,N_10446,N_14760);
nor U16061 (N_16061,N_12784,N_14472);
or U16062 (N_16062,N_14026,N_13403);
xor U16063 (N_16063,N_12440,N_11366);
nand U16064 (N_16064,N_11708,N_13281);
xnor U16065 (N_16065,N_10270,N_13567);
xor U16066 (N_16066,N_13257,N_10413);
nor U16067 (N_16067,N_12691,N_14978);
nor U16068 (N_16068,N_14442,N_13356);
xor U16069 (N_16069,N_12269,N_11386);
or U16070 (N_16070,N_14542,N_14348);
or U16071 (N_16071,N_14656,N_14936);
nand U16072 (N_16072,N_14742,N_12283);
nand U16073 (N_16073,N_12830,N_14889);
nand U16074 (N_16074,N_11519,N_12244);
or U16075 (N_16075,N_14008,N_13598);
nand U16076 (N_16076,N_10503,N_11555);
and U16077 (N_16077,N_14046,N_12174);
xor U16078 (N_16078,N_10943,N_11305);
nor U16079 (N_16079,N_14953,N_13100);
xnor U16080 (N_16080,N_14515,N_10035);
or U16081 (N_16081,N_10883,N_11715);
and U16082 (N_16082,N_10713,N_12978);
xor U16083 (N_16083,N_12029,N_12335);
xnor U16084 (N_16084,N_13111,N_10700);
or U16085 (N_16085,N_10873,N_14407);
nand U16086 (N_16086,N_12964,N_11704);
xnor U16087 (N_16087,N_14323,N_14998);
nand U16088 (N_16088,N_13214,N_10159);
and U16089 (N_16089,N_13679,N_13971);
nand U16090 (N_16090,N_10306,N_11551);
and U16091 (N_16091,N_11827,N_14963);
or U16092 (N_16092,N_10467,N_11593);
nand U16093 (N_16093,N_13956,N_12136);
xor U16094 (N_16094,N_12989,N_10098);
nand U16095 (N_16095,N_14196,N_10300);
nor U16096 (N_16096,N_10864,N_10407);
or U16097 (N_16097,N_11700,N_10983);
or U16098 (N_16098,N_12287,N_12540);
nor U16099 (N_16099,N_11440,N_12610);
xor U16100 (N_16100,N_13087,N_14069);
nand U16101 (N_16101,N_12129,N_12819);
nand U16102 (N_16102,N_11252,N_14110);
nor U16103 (N_16103,N_10189,N_13435);
nor U16104 (N_16104,N_12653,N_12462);
nand U16105 (N_16105,N_13279,N_11780);
or U16106 (N_16106,N_13248,N_13473);
xnor U16107 (N_16107,N_11763,N_13417);
nand U16108 (N_16108,N_10285,N_12371);
nand U16109 (N_16109,N_10681,N_14299);
nand U16110 (N_16110,N_12981,N_12645);
and U16111 (N_16111,N_14060,N_12795);
and U16112 (N_16112,N_11330,N_10123);
and U16113 (N_16113,N_11408,N_12983);
nor U16114 (N_16114,N_12859,N_10844);
nand U16115 (N_16115,N_10688,N_10085);
nor U16116 (N_16116,N_11095,N_10198);
or U16117 (N_16117,N_10974,N_12187);
and U16118 (N_16118,N_14589,N_13094);
and U16119 (N_16119,N_13750,N_13748);
or U16120 (N_16120,N_12336,N_12304);
or U16121 (N_16121,N_10203,N_14741);
nor U16122 (N_16122,N_14296,N_11170);
nor U16123 (N_16123,N_12101,N_13773);
or U16124 (N_16124,N_14658,N_13362);
and U16125 (N_16125,N_12060,N_10477);
nand U16126 (N_16126,N_10075,N_10588);
xor U16127 (N_16127,N_10096,N_14562);
xnor U16128 (N_16128,N_14123,N_13880);
and U16129 (N_16129,N_14450,N_11137);
or U16130 (N_16130,N_12958,N_13871);
nand U16131 (N_16131,N_14522,N_10712);
nor U16132 (N_16132,N_13431,N_13230);
or U16133 (N_16133,N_12977,N_11543);
or U16134 (N_16134,N_12886,N_12014);
nor U16135 (N_16135,N_10989,N_11050);
nand U16136 (N_16136,N_14660,N_10914);
or U16137 (N_16137,N_11513,N_10954);
and U16138 (N_16138,N_14531,N_10289);
and U16139 (N_16139,N_13683,N_11673);
xor U16140 (N_16140,N_13445,N_10505);
xnor U16141 (N_16141,N_13961,N_12868);
and U16142 (N_16142,N_14975,N_14359);
nor U16143 (N_16143,N_11805,N_10447);
or U16144 (N_16144,N_14668,N_14574);
nand U16145 (N_16145,N_11959,N_12596);
or U16146 (N_16146,N_13168,N_11417);
or U16147 (N_16147,N_13847,N_13707);
xnor U16148 (N_16148,N_13806,N_13167);
nand U16149 (N_16149,N_11793,N_13143);
nand U16150 (N_16150,N_13953,N_10387);
nor U16151 (N_16151,N_11004,N_10023);
nand U16152 (N_16152,N_11584,N_10341);
nor U16153 (N_16153,N_10311,N_10786);
or U16154 (N_16154,N_12929,N_10815);
and U16155 (N_16155,N_10907,N_10509);
nand U16156 (N_16156,N_10271,N_13020);
xnor U16157 (N_16157,N_14045,N_12464);
nor U16158 (N_16158,N_13339,N_11926);
xor U16159 (N_16159,N_11335,N_13876);
or U16160 (N_16160,N_13873,N_13349);
and U16161 (N_16161,N_11487,N_14477);
nor U16162 (N_16162,N_11791,N_14071);
and U16163 (N_16163,N_13217,N_12310);
or U16164 (N_16164,N_10863,N_14388);
and U16165 (N_16165,N_11393,N_14526);
or U16166 (N_16166,N_13651,N_13714);
or U16167 (N_16167,N_11008,N_10365);
nand U16168 (N_16168,N_10402,N_13854);
nand U16169 (N_16169,N_11818,N_10798);
xor U16170 (N_16170,N_13044,N_14087);
xor U16171 (N_16171,N_12303,N_13197);
or U16172 (N_16172,N_13424,N_12483);
and U16173 (N_16173,N_14177,N_11636);
nor U16174 (N_16174,N_13367,N_14637);
xnor U16175 (N_16175,N_13826,N_13152);
nor U16176 (N_16176,N_10053,N_10069);
or U16177 (N_16177,N_13205,N_11617);
nor U16178 (N_16178,N_13952,N_14536);
and U16179 (N_16179,N_13080,N_14004);
or U16180 (N_16180,N_11269,N_13809);
and U16181 (N_16181,N_11232,N_13906);
nand U16182 (N_16182,N_14427,N_13638);
nor U16183 (N_16183,N_14694,N_10622);
and U16184 (N_16184,N_10345,N_12077);
and U16185 (N_16185,N_10459,N_12302);
nand U16186 (N_16186,N_12751,N_13822);
or U16187 (N_16187,N_10567,N_12314);
xor U16188 (N_16188,N_12502,N_13673);
xor U16189 (N_16189,N_13665,N_11898);
nand U16190 (N_16190,N_11402,N_12952);
or U16191 (N_16191,N_10878,N_13201);
and U16192 (N_16192,N_14823,N_14756);
and U16193 (N_16193,N_12720,N_11113);
nand U16194 (N_16194,N_12148,N_10013);
nor U16195 (N_16195,N_11002,N_11567);
xnor U16196 (N_16196,N_11872,N_12512);
or U16197 (N_16197,N_11446,N_14355);
nand U16198 (N_16198,N_13689,N_11738);
xnor U16199 (N_16199,N_14270,N_13789);
or U16200 (N_16200,N_11835,N_14067);
nand U16201 (N_16201,N_10826,N_11956);
or U16202 (N_16202,N_13733,N_12702);
xor U16203 (N_16203,N_10739,N_11072);
nand U16204 (N_16204,N_14445,N_14857);
xor U16205 (N_16205,N_13467,N_10022);
and U16206 (N_16206,N_14049,N_10302);
xor U16207 (N_16207,N_14001,N_13381);
nor U16208 (N_16208,N_11687,N_11503);
nor U16209 (N_16209,N_10382,N_11892);
xnor U16210 (N_16210,N_12048,N_13374);
or U16211 (N_16211,N_13675,N_10232);
nand U16212 (N_16212,N_13589,N_12059);
and U16213 (N_16213,N_13342,N_11209);
xnor U16214 (N_16214,N_14525,N_12273);
nor U16215 (N_16215,N_13242,N_14827);
and U16216 (N_16216,N_11970,N_12974);
and U16217 (N_16217,N_13129,N_12976);
and U16218 (N_16218,N_13676,N_11358);
and U16219 (N_16219,N_12388,N_13732);
or U16220 (N_16220,N_14044,N_11531);
nand U16221 (N_16221,N_13141,N_14603);
or U16222 (N_16222,N_11806,N_10781);
nand U16223 (N_16223,N_10215,N_11323);
xor U16224 (N_16224,N_12515,N_11140);
and U16225 (N_16225,N_12842,N_13460);
nand U16226 (N_16226,N_10011,N_11849);
nand U16227 (N_16227,N_10246,N_11754);
and U16228 (N_16228,N_11347,N_12307);
nand U16229 (N_16229,N_11495,N_13007);
xor U16230 (N_16230,N_13957,N_11452);
xor U16231 (N_16231,N_11314,N_13991);
and U16232 (N_16232,N_10204,N_12782);
or U16233 (N_16233,N_12854,N_13068);
or U16234 (N_16234,N_14543,N_13065);
or U16235 (N_16235,N_12700,N_13323);
xor U16236 (N_16236,N_12902,N_14724);
nand U16237 (N_16237,N_10600,N_14400);
nand U16238 (N_16238,N_13938,N_14552);
xor U16239 (N_16239,N_12803,N_10442);
and U16240 (N_16240,N_11644,N_12488);
nor U16241 (N_16241,N_13225,N_10064);
or U16242 (N_16242,N_11610,N_14418);
nor U16243 (N_16243,N_10167,N_14872);
or U16244 (N_16244,N_11343,N_11731);
xnor U16245 (N_16245,N_10342,N_13496);
xor U16246 (N_16246,N_11587,N_14120);
nand U16247 (N_16247,N_11156,N_10385);
nor U16248 (N_16248,N_10672,N_14480);
and U16249 (N_16249,N_12166,N_13449);
and U16250 (N_16250,N_14941,N_10364);
or U16251 (N_16251,N_13912,N_10150);
nand U16252 (N_16252,N_12350,N_13669);
xnor U16253 (N_16253,N_13778,N_13866);
and U16254 (N_16254,N_11368,N_13780);
nor U16255 (N_16255,N_12903,N_11762);
xnor U16256 (N_16256,N_11857,N_11344);
nand U16257 (N_16257,N_14689,N_12792);
nor U16258 (N_16258,N_14424,N_10152);
nand U16259 (N_16259,N_14849,N_14038);
nor U16260 (N_16260,N_10160,N_10996);
and U16261 (N_16261,N_11641,N_10912);
and U16262 (N_16262,N_10908,N_10939);
nand U16263 (N_16263,N_10080,N_11340);
xnor U16264 (N_16264,N_12000,N_14881);
and U16265 (N_16265,N_14197,N_14651);
xnor U16266 (N_16266,N_11540,N_11914);
nor U16267 (N_16267,N_12076,N_10014);
and U16268 (N_16268,N_12544,N_10506);
nand U16269 (N_16269,N_13459,N_11254);
and U16270 (N_16270,N_10707,N_14487);
and U16271 (N_16271,N_12710,N_14491);
and U16272 (N_16272,N_13593,N_14680);
xor U16273 (N_16273,N_14970,N_12947);
or U16274 (N_16274,N_11730,N_11938);
nor U16275 (N_16275,N_14412,N_14274);
xnor U16276 (N_16276,N_14777,N_12232);
nand U16277 (N_16277,N_14511,N_14041);
or U16278 (N_16278,N_14468,N_14897);
xnor U16279 (N_16279,N_11325,N_11952);
and U16280 (N_16280,N_11753,N_11107);
nor U16281 (N_16281,N_14225,N_11911);
xnor U16282 (N_16282,N_11226,N_14286);
and U16283 (N_16283,N_13688,N_13432);
and U16284 (N_16284,N_11057,N_13648);
xor U16285 (N_16285,N_12862,N_11695);
nand U16286 (N_16286,N_11993,N_10767);
nand U16287 (N_16287,N_11024,N_11568);
xnor U16288 (N_16288,N_10902,N_10969);
or U16289 (N_16289,N_11363,N_11984);
nor U16290 (N_16290,N_11125,N_14027);
nor U16291 (N_16291,N_12769,N_12300);
or U16292 (N_16292,N_12494,N_13490);
or U16293 (N_16293,N_10491,N_11944);
or U16294 (N_16294,N_14826,N_10514);
nand U16295 (N_16295,N_12199,N_10972);
or U16296 (N_16296,N_14366,N_14471);
nand U16297 (N_16297,N_11215,N_14386);
and U16298 (N_16298,N_11633,N_12394);
and U16299 (N_16299,N_13601,N_14996);
xor U16300 (N_16300,N_13273,N_13055);
and U16301 (N_16301,N_13948,N_13493);
nor U16302 (N_16302,N_12719,N_14253);
xor U16303 (N_16303,N_14635,N_10095);
xnor U16304 (N_16304,N_10550,N_13413);
and U16305 (N_16305,N_14107,N_10212);
xnor U16306 (N_16306,N_14191,N_14627);
nor U16307 (N_16307,N_13119,N_10677);
or U16308 (N_16308,N_13289,N_11874);
and U16309 (N_16309,N_12880,N_13963);
xnor U16310 (N_16310,N_11773,N_11052);
nor U16311 (N_16311,N_11003,N_13453);
nor U16312 (N_16312,N_10691,N_11247);
or U16313 (N_16313,N_10811,N_11671);
xor U16314 (N_16314,N_13376,N_14653);
nor U16315 (N_16315,N_14159,N_12874);
and U16316 (N_16316,N_12843,N_13052);
nand U16317 (N_16317,N_11741,N_11941);
nor U16318 (N_16318,N_14440,N_10027);
nand U16319 (N_16319,N_13712,N_10234);
nand U16320 (N_16320,N_10435,N_12545);
or U16321 (N_16321,N_14918,N_11592);
or U16322 (N_16322,N_10162,N_10746);
nor U16323 (N_16323,N_14900,N_12578);
nor U16324 (N_16324,N_11627,N_11501);
nor U16325 (N_16325,N_14237,N_11646);
nor U16326 (N_16326,N_11126,N_14014);
and U16327 (N_16327,N_10117,N_14223);
or U16328 (N_16328,N_14173,N_10257);
nor U16329 (N_16329,N_11580,N_11277);
or U16330 (N_16330,N_13670,N_13192);
xnor U16331 (N_16331,N_10607,N_11298);
nor U16332 (N_16332,N_11105,N_11289);
or U16333 (N_16333,N_13802,N_14720);
xnor U16334 (N_16334,N_12796,N_13535);
and U16335 (N_16335,N_12276,N_13033);
xor U16336 (N_16336,N_14321,N_12133);
nor U16337 (N_16337,N_12878,N_10381);
or U16338 (N_16338,N_12632,N_14494);
or U16339 (N_16339,N_12589,N_14258);
nand U16340 (N_16340,N_14182,N_14462);
xor U16341 (N_16341,N_11761,N_12995);
or U16342 (N_16342,N_14420,N_12134);
xnor U16343 (N_16343,N_13202,N_11639);
xor U16344 (N_16344,N_10070,N_14524);
xnor U16345 (N_16345,N_11115,N_13935);
or U16346 (N_16346,N_12459,N_13050);
and U16347 (N_16347,N_11255,N_10439);
nor U16348 (N_16348,N_12846,N_12410);
nand U16349 (N_16349,N_12364,N_11983);
nor U16350 (N_16350,N_13703,N_13287);
or U16351 (N_16351,N_11719,N_13674);
xnor U16352 (N_16352,N_14241,N_13979);
or U16353 (N_16353,N_12155,N_10755);
or U16354 (N_16354,N_10977,N_10860);
nand U16355 (N_16355,N_14373,N_14063);
nand U16356 (N_16356,N_14200,N_12118);
nor U16357 (N_16357,N_14380,N_11418);
nand U16358 (N_16358,N_13495,N_12100);
or U16359 (N_16359,N_12108,N_13846);
nand U16360 (N_16360,N_14346,N_10975);
nor U16361 (N_16361,N_11689,N_10765);
nor U16362 (N_16362,N_11684,N_14597);
nand U16363 (N_16363,N_11453,N_14690);
nand U16364 (N_16364,N_10909,N_12281);
or U16365 (N_16365,N_12202,N_14235);
and U16366 (N_16366,N_11645,N_14476);
and U16367 (N_16367,N_12572,N_10434);
xnor U16368 (N_16368,N_12762,N_14153);
xnor U16369 (N_16369,N_14615,N_10391);
or U16370 (N_16370,N_12449,N_10440);
xnor U16371 (N_16371,N_13372,N_10891);
nand U16372 (N_16372,N_11405,N_12144);
or U16373 (N_16373,N_14488,N_11073);
or U16374 (N_16374,N_11565,N_14370);
or U16375 (N_16375,N_12527,N_13743);
and U16376 (N_16376,N_13643,N_10956);
or U16377 (N_16377,N_14535,N_12993);
xnor U16378 (N_16378,N_11122,N_13062);
xnor U16379 (N_16379,N_12019,N_14449);
nor U16380 (N_16380,N_13965,N_14309);
nand U16381 (N_16381,N_10316,N_12662);
xor U16382 (N_16382,N_14082,N_14666);
nor U16383 (N_16383,N_14256,N_13251);
or U16384 (N_16384,N_12035,N_10644);
nand U16385 (N_16385,N_11098,N_11545);
nand U16386 (N_16386,N_12810,N_14202);
nand U16387 (N_16387,N_14000,N_12892);
and U16388 (N_16388,N_11526,N_10173);
or U16389 (N_16389,N_14599,N_12047);
xor U16390 (N_16390,N_12365,N_14563);
nand U16391 (N_16391,N_11354,N_11488);
or U16392 (N_16392,N_11850,N_12180);
nand U16393 (N_16393,N_14021,N_13716);
and U16394 (N_16394,N_11204,N_12055);
and U16395 (N_16395,N_13499,N_12280);
and U16396 (N_16396,N_14376,N_11208);
and U16397 (N_16397,N_12927,N_10268);
nor U16398 (N_16398,N_13049,N_13175);
and U16399 (N_16399,N_12725,N_12121);
or U16400 (N_16400,N_11182,N_12778);
or U16401 (N_16401,N_14598,N_12602);
and U16402 (N_16402,N_14804,N_14699);
nor U16403 (N_16403,N_12758,N_13042);
nand U16404 (N_16404,N_13375,N_11274);
nand U16405 (N_16405,N_14984,N_10624);
xor U16406 (N_16406,N_11483,N_14577);
and U16407 (N_16407,N_10380,N_12705);
nand U16408 (N_16408,N_11603,N_12737);
and U16409 (N_16409,N_11250,N_13775);
xnor U16410 (N_16410,N_11693,N_10875);
nor U16411 (N_16411,N_13879,N_10852);
nor U16412 (N_16412,N_12715,N_10431);
nor U16413 (N_16413,N_12267,N_10228);
nor U16414 (N_16414,N_12811,N_11164);
and U16415 (N_16415,N_10443,N_12432);
and U16416 (N_16416,N_14428,N_12930);
and U16417 (N_16417,N_10094,N_12312);
nand U16418 (N_16418,N_10329,N_14948);
or U16419 (N_16419,N_13191,N_12490);
nor U16420 (N_16420,N_10946,N_14290);
nor U16421 (N_16421,N_13887,N_12173);
and U16422 (N_16422,N_14093,N_10343);
xnor U16423 (N_16423,N_13472,N_14088);
xor U16424 (N_16424,N_14834,N_13410);
nor U16425 (N_16425,N_10415,N_14228);
nor U16426 (N_16426,N_13588,N_12922);
xnor U16427 (N_16427,N_12454,N_12813);
xor U16428 (N_16428,N_14871,N_11374);
or U16429 (N_16429,N_14909,N_14514);
or U16430 (N_16430,N_12285,N_10632);
nor U16431 (N_16431,N_12031,N_11385);
and U16432 (N_16432,N_14163,N_11945);
and U16433 (N_16433,N_12105,N_13031);
xnor U16434 (N_16434,N_12154,N_14265);
and U16435 (N_16435,N_10211,N_10145);
or U16436 (N_16436,N_11524,N_14904);
nor U16437 (N_16437,N_14013,N_14958);
nand U16438 (N_16438,N_12528,N_10315);
nor U16439 (N_16439,N_11790,N_12701);
nand U16440 (N_16440,N_10183,N_13429);
xnor U16441 (N_16441,N_14828,N_14621);
nand U16442 (N_16442,N_14136,N_14766);
xor U16443 (N_16443,N_12546,N_12604);
nand U16444 (N_16444,N_13288,N_10416);
nand U16445 (N_16445,N_11191,N_10776);
or U16446 (N_16446,N_12508,N_11870);
nand U16447 (N_16447,N_14057,N_11800);
and U16448 (N_16448,N_14501,N_10122);
nand U16449 (N_16449,N_11696,N_12750);
and U16450 (N_16450,N_14914,N_12216);
and U16451 (N_16451,N_12147,N_11014);
and U16452 (N_16452,N_12816,N_11198);
or U16453 (N_16453,N_10536,N_10576);
xor U16454 (N_16454,N_12744,N_12801);
nor U16455 (N_16455,N_11582,N_11301);
nor U16456 (N_16456,N_14622,N_10131);
nor U16457 (N_16457,N_10401,N_10048);
nand U16458 (N_16458,N_12181,N_13450);
and U16459 (N_16459,N_14906,N_10320);
or U16460 (N_16460,N_12017,N_10549);
or U16461 (N_16461,N_11901,N_12353);
nand U16462 (N_16462,N_14052,N_12444);
and U16463 (N_16463,N_10322,N_13208);
xnor U16464 (N_16464,N_13524,N_14127);
xor U16465 (N_16465,N_11167,N_11922);
nor U16466 (N_16466,N_12286,N_12357);
xnor U16467 (N_16467,N_11705,N_13964);
and U16468 (N_16468,N_13199,N_13344);
nor U16469 (N_16469,N_12373,N_11270);
xor U16470 (N_16470,N_11451,N_11674);
and U16471 (N_16471,N_13592,N_10286);
nor U16472 (N_16472,N_12477,N_13075);
or U16473 (N_16473,N_13568,N_14564);
nor U16474 (N_16474,N_12773,N_11049);
and U16475 (N_16475,N_10823,N_11480);
and U16476 (N_16476,N_11465,N_10103);
and U16477 (N_16477,N_11394,N_11624);
nor U16478 (N_16478,N_13333,N_14054);
or U16479 (N_16479,N_14455,N_10049);
nand U16480 (N_16480,N_13718,N_10962);
or U16481 (N_16481,N_11697,N_13312);
xnor U16482 (N_16482,N_12445,N_13148);
and U16483 (N_16483,N_14788,N_13929);
nand U16484 (N_16484,N_10111,N_14398);
xnor U16485 (N_16485,N_12135,N_11245);
or U16486 (N_16486,N_10240,N_10326);
or U16487 (N_16487,N_12944,N_11411);
xor U16488 (N_16488,N_10444,N_12288);
nor U16489 (N_16489,N_12712,N_13384);
nand U16490 (N_16490,N_13551,N_11030);
nand U16491 (N_16491,N_10184,N_12591);
or U16492 (N_16492,N_10455,N_14452);
nor U16493 (N_16493,N_13690,N_12460);
nand U16494 (N_16494,N_12606,N_14190);
and U16495 (N_16495,N_14723,N_12437);
and U16496 (N_16496,N_11076,N_11921);
and U16497 (N_16497,N_10782,N_12936);
and U16498 (N_16498,N_14220,N_11865);
nand U16499 (N_16499,N_12650,N_10115);
and U16500 (N_16500,N_14540,N_12214);
or U16501 (N_16501,N_13098,N_12535);
nor U16502 (N_16502,N_13091,N_14070);
xor U16503 (N_16503,N_12340,N_14230);
and U16504 (N_16504,N_10492,N_11573);
and U16505 (N_16505,N_11726,N_14647);
or U16506 (N_16506,N_10551,N_11294);
nor U16507 (N_16507,N_10834,N_11101);
nor U16508 (N_16508,N_12689,N_10404);
and U16509 (N_16509,N_11010,N_12045);
nand U16510 (N_16510,N_11821,N_11077);
nand U16511 (N_16511,N_13591,N_13383);
and U16512 (N_16512,N_14738,N_12206);
nand U16513 (N_16513,N_12458,N_14358);
xnor U16514 (N_16514,N_10553,N_10441);
nor U16515 (N_16515,N_14721,N_10920);
or U16516 (N_16516,N_14648,N_13787);
or U16517 (N_16517,N_12405,N_10041);
or U16518 (N_16518,N_12438,N_11414);
nand U16519 (N_16519,N_10020,N_14613);
or U16520 (N_16520,N_12496,N_13096);
nand U16521 (N_16521,N_11416,N_14786);
or U16522 (N_16522,N_11812,N_13756);
nor U16523 (N_16523,N_11149,N_10220);
or U16524 (N_16524,N_12920,N_14675);
or U16525 (N_16525,N_12470,N_12857);
nor U16526 (N_16526,N_12537,N_12395);
or U16527 (N_16527,N_11040,N_11352);
nor U16528 (N_16528,N_11189,N_12807);
and U16529 (N_16529,N_10825,N_10924);
or U16530 (N_16530,N_10097,N_10803);
nand U16531 (N_16531,N_14709,N_12894);
or U16532 (N_16532,N_14430,N_12113);
nor U16533 (N_16533,N_13664,N_11851);
xor U16534 (N_16534,N_13216,N_14645);
nand U16535 (N_16535,N_11457,N_11811);
or U16536 (N_16536,N_12884,N_10274);
or U16537 (N_16537,N_14329,N_14949);
nand U16538 (N_16538,N_12560,N_10298);
nand U16539 (N_16539,N_14089,N_13908);
nor U16540 (N_16540,N_10543,N_10333);
xnor U16541 (N_16541,N_14248,N_11891);
xor U16542 (N_16542,N_11652,N_12659);
and U16543 (N_16543,N_10879,N_11046);
nand U16544 (N_16544,N_12988,N_11614);
nor U16545 (N_16545,N_14227,N_13654);
nor U16546 (N_16546,N_14233,N_11541);
nand U16547 (N_16547,N_11065,N_12109);
xor U16548 (N_16548,N_10694,N_10640);
xnor U16549 (N_16549,N_14840,N_14317);
or U16550 (N_16550,N_14152,N_13629);
or U16551 (N_16551,N_12848,N_11175);
xnor U16552 (N_16552,N_12781,N_11920);
nand U16553 (N_16553,N_13263,N_12071);
xor U16554 (N_16554,N_12504,N_10910);
xor U16555 (N_16555,N_14003,N_13021);
nor U16556 (N_16556,N_12955,N_10482);
nor U16557 (N_16557,N_14670,N_12141);
nand U16558 (N_16558,N_14504,N_12609);
xnor U16559 (N_16559,N_13844,N_10548);
or U16560 (N_16560,N_14974,N_10645);
nand U16561 (N_16561,N_12831,N_13552);
nand U16562 (N_16562,N_11000,N_14339);
or U16563 (N_16563,N_10986,N_10812);
or U16564 (N_16564,N_14798,N_12305);
or U16565 (N_16565,N_14195,N_10112);
and U16566 (N_16566,N_14347,N_12399);
nand U16567 (N_16567,N_10104,N_10669);
nand U16568 (N_16568,N_14937,N_13235);
nor U16569 (N_16569,N_10936,N_14708);
and U16570 (N_16570,N_14633,N_11357);
xor U16571 (N_16571,N_11782,N_13521);
nor U16572 (N_16572,N_10738,N_13719);
nor U16573 (N_16573,N_10580,N_10451);
or U16574 (N_16574,N_11036,N_10582);
nor U16575 (N_16575,N_14187,N_11442);
and U16576 (N_16576,N_14843,N_13497);
nand U16577 (N_16577,N_13115,N_14654);
xnor U16578 (N_16578,N_12158,N_13931);
nor U16579 (N_16579,N_12439,N_12319);
xnor U16580 (N_16580,N_14349,N_11967);
or U16581 (N_16581,N_13008,N_10725);
nor U16582 (N_16582,N_13285,N_14740);
and U16583 (N_16583,N_10905,N_10750);
xnor U16584 (N_16584,N_14305,N_10358);
nor U16585 (N_16585,N_10695,N_12320);
nor U16586 (N_16586,N_10870,N_13073);
or U16587 (N_16587,N_11839,N_12052);
xnor U16588 (N_16588,N_13268,N_13558);
nand U16589 (N_16589,N_14527,N_12308);
nor U16590 (N_16590,N_10396,N_11749);
and U16591 (N_16591,N_10028,N_14019);
nor U16592 (N_16592,N_10337,N_14789);
xnor U16593 (N_16593,N_11912,N_11066);
and U16594 (N_16594,N_10109,N_14739);
nand U16595 (N_16595,N_10350,N_13570);
nand U16596 (N_16596,N_10293,N_11842);
or U16597 (N_16597,N_13518,N_13145);
or U16598 (N_16598,N_12441,N_11445);
nor U16599 (N_16599,N_12352,N_10931);
nor U16600 (N_16600,N_11825,N_12264);
nor U16601 (N_16601,N_12666,N_10941);
and U16602 (N_16602,N_13848,N_12619);
xor U16603 (N_16603,N_12505,N_10627);
and U16604 (N_16604,N_12370,N_10222);
or U16605 (N_16605,N_13188,N_14304);
and U16606 (N_16606,N_10953,N_13576);
xor U16607 (N_16607,N_10886,N_14686);
or U16608 (N_16608,N_10389,N_12906);
xnor U16609 (N_16609,N_12372,N_14762);
or U16610 (N_16610,N_13966,N_12597);
nand U16611 (N_16611,N_14726,N_14092);
nand U16612 (N_16612,N_13694,N_12721);
or U16613 (N_16613,N_14356,N_10757);
nand U16614 (N_16614,N_14519,N_13084);
or U16615 (N_16615,N_10465,N_13319);
nor U16616 (N_16616,N_12086,N_10683);
or U16617 (N_16617,N_14434,N_10837);
and U16618 (N_16618,N_12882,N_14130);
xor U16619 (N_16619,N_11214,N_12951);
xor U16620 (N_16620,N_14231,N_13973);
or U16621 (N_16621,N_13291,N_12900);
nor U16622 (N_16622,N_13269,N_14802);
and U16623 (N_16623,N_10243,N_13244);
or U16624 (N_16624,N_11237,N_14746);
and U16625 (N_16625,N_11013,N_11985);
and U16626 (N_16626,N_14282,N_14824);
xnor U16627 (N_16627,N_14842,N_10999);
and U16628 (N_16628,N_12272,N_14533);
or U16629 (N_16629,N_10578,N_13004);
or U16630 (N_16630,N_13457,N_13856);
nand U16631 (N_16631,N_13002,N_11560);
or U16632 (N_16632,N_11933,N_13015);
or U16633 (N_16633,N_14466,N_11201);
or U16634 (N_16634,N_13722,N_11917);
nor U16635 (N_16635,N_11192,N_12337);
nand U16636 (N_16636,N_11109,N_14319);
and U16637 (N_16637,N_12406,N_13361);
or U16638 (N_16638,N_10763,N_13788);
nor U16639 (N_16639,N_10540,N_14188);
xnor U16640 (N_16640,N_13172,N_11312);
nand U16641 (N_16641,N_11257,N_11910);
xnor U16642 (N_16642,N_11525,N_11316);
xor U16643 (N_16643,N_10258,N_14042);
or U16644 (N_16644,N_10458,N_10662);
xor U16645 (N_16645,N_12083,N_12398);
nand U16646 (N_16646,N_11458,N_12912);
xor U16647 (N_16647,N_12649,N_12646);
and U16648 (N_16648,N_13245,N_12941);
nor U16649 (N_16649,N_10670,N_12027);
or U16650 (N_16650,N_13284,N_12531);
nor U16651 (N_16651,N_11005,N_13796);
and U16652 (N_16652,N_11234,N_13602);
or U16653 (N_16653,N_10409,N_14215);
or U16654 (N_16654,N_12222,N_13762);
and U16655 (N_16655,N_11319,N_13069);
or U16656 (N_16656,N_13471,N_10247);
and U16657 (N_16657,N_13234,N_10926);
nand U16658 (N_16658,N_14930,N_11735);
or U16659 (N_16659,N_11506,N_10730);
or U16660 (N_16660,N_12054,N_13672);
or U16661 (N_16661,N_11025,N_10498);
or U16662 (N_16662,N_12467,N_10994);
nand U16663 (N_16663,N_12209,N_10611);
or U16664 (N_16664,N_10916,N_10655);
or U16665 (N_16665,N_14631,N_13258);
and U16666 (N_16666,N_14109,N_12658);
and U16667 (N_16667,N_12707,N_10484);
nor U16668 (N_16668,N_13736,N_13515);
and U16669 (N_16669,N_12834,N_11239);
xor U16670 (N_16670,N_10275,N_10126);
nor U16671 (N_16671,N_10106,N_14263);
or U16672 (N_16672,N_10978,N_13776);
or U16673 (N_16673,N_12753,N_10021);
and U16674 (N_16674,N_11698,N_13698);
nor U16675 (N_16675,N_13768,N_12684);
nand U16676 (N_16676,N_12111,N_12360);
nand U16677 (N_16677,N_11217,N_12237);
nor U16678 (N_16678,N_14318,N_11707);
xor U16679 (N_16679,N_12092,N_12895);
and U16680 (N_16680,N_13514,N_12759);
nand U16681 (N_16681,N_14922,N_14178);
or U16682 (N_16682,N_10281,N_12946);
and U16683 (N_16683,N_10615,N_14500);
nand U16684 (N_16684,N_13816,N_11848);
nor U16685 (N_16685,N_12963,N_10764);
nand U16686 (N_16686,N_14614,N_14186);
xnor U16687 (N_16687,N_14628,N_14607);
xnor U16688 (N_16688,N_14938,N_11326);
xor U16689 (N_16689,N_14337,N_12728);
nand U16690 (N_16690,N_13751,N_13666);
or U16691 (N_16691,N_10464,N_14119);
or U16692 (N_16692,N_13731,N_11760);
nor U16693 (N_16693,N_10284,N_10411);
xor U16694 (N_16694,N_13057,N_11974);
nand U16695 (N_16695,N_14279,N_14091);
nor U16696 (N_16696,N_13006,N_13525);
xor U16697 (N_16697,N_14817,N_11757);
nor U16698 (N_16698,N_12259,N_10845);
nor U16699 (N_16699,N_11796,N_11903);
xor U16700 (N_16700,N_12524,N_10158);
nor U16701 (N_16701,N_10138,N_12980);
or U16702 (N_16702,N_13252,N_10221);
nor U16703 (N_16703,N_14194,N_10288);
and U16704 (N_16704,N_12387,N_12025);
or U16705 (N_16705,N_13936,N_13482);
and U16706 (N_16706,N_12918,N_10471);
and U16707 (N_16707,N_13634,N_14663);
nor U16708 (N_16708,N_11579,N_14254);
xor U16709 (N_16709,N_11904,N_14702);
and U16710 (N_16710,N_14224,N_12261);
nor U16711 (N_16711,N_14226,N_12523);
nand U16712 (N_16712,N_10848,N_10742);
nand U16713 (N_16713,N_12330,N_10570);
xor U16714 (N_16714,N_14888,N_12456);
and U16715 (N_16715,N_14714,N_11807);
or U16716 (N_16716,N_10935,N_14343);
or U16717 (N_16717,N_14417,N_13943);
and U16718 (N_16718,N_14023,N_10168);
nand U16719 (N_16719,N_13919,N_12836);
nor U16720 (N_16720,N_11544,N_11199);
nor U16721 (N_16721,N_11128,N_12798);
nor U16722 (N_16722,N_12869,N_10015);
nand U16723 (N_16723,N_14075,N_13442);
nand U16724 (N_16724,N_13610,N_10478);
nand U16725 (N_16725,N_14629,N_10884);
xor U16726 (N_16726,N_11990,N_10108);
nor U16727 (N_16727,N_11718,N_10290);
xor U16728 (N_16728,N_10090,N_10499);
nand U16729 (N_16729,N_11744,N_12013);
and U16730 (N_16730,N_12489,N_10139);
nor U16731 (N_16731,N_12940,N_10209);
nor U16732 (N_16732,N_14980,N_14815);
and U16733 (N_16733,N_11664,N_10519);
and U16734 (N_16734,N_11653,N_14166);
nand U16735 (N_16735,N_11721,N_11069);
or U16736 (N_16736,N_13682,N_14700);
xnor U16737 (N_16737,N_13072,N_13047);
and U16738 (N_16738,N_12104,N_14205);
and U16739 (N_16739,N_10360,N_12224);
xnor U16740 (N_16740,N_13401,N_14662);
xnor U16741 (N_16741,N_10223,N_10741);
or U16742 (N_16742,N_14204,N_13813);
xnor U16743 (N_16743,N_13247,N_14145);
nor U16744 (N_16744,N_11756,N_12838);
or U16745 (N_16745,N_14555,N_11054);
xor U16746 (N_16746,N_13962,N_12379);
and U16747 (N_16747,N_10490,N_12690);
and U16748 (N_16748,N_10356,N_11039);
and U16749 (N_16749,N_10087,N_10132);
nor U16750 (N_16750,N_12729,N_10355);
nand U16751 (N_16751,N_13663,N_12706);
nand U16752 (N_16752,N_14390,N_14800);
nor U16753 (N_16753,N_11963,N_14383);
nor U16754 (N_16754,N_10625,N_11605);
nor U16755 (N_16755,N_11119,N_14829);
xor U16756 (N_16756,N_11585,N_11537);
nand U16757 (N_16757,N_11979,N_12863);
or U16758 (N_16758,N_10445,N_11202);
nor U16759 (N_16759,N_12263,N_12381);
xnor U16760 (N_16760,N_12299,N_10718);
or U16761 (N_16761,N_12002,N_11258);
nand U16762 (N_16762,N_12452,N_14415);
nor U16763 (N_16763,N_14776,N_10685);
or U16764 (N_16764,N_13932,N_14103);
nor U16765 (N_16765,N_11213,N_10010);
xor U16766 (N_16766,N_12669,N_10950);
xnor U16767 (N_16767,N_11802,N_13325);
nor U16768 (N_16768,N_11218,N_11087);
xnor U16769 (N_16769,N_10720,N_13079);
xnor U16770 (N_16770,N_10428,N_12178);
nor U16771 (N_16771,N_10934,N_10394);
or U16772 (N_16772,N_11466,N_13611);
or U16773 (N_16773,N_12893,N_11623);
nor U16774 (N_16774,N_12172,N_14677);
and U16775 (N_16775,N_13785,N_12718);
or U16776 (N_16776,N_14588,N_12177);
nand U16777 (N_16777,N_10421,N_11224);
and U16778 (N_16778,N_11282,N_10026);
nand U16779 (N_16779,N_14990,N_11734);
nand U16780 (N_16780,N_13037,N_12682);
xor U16781 (N_16781,N_12881,N_11051);
and U16782 (N_16782,N_12536,N_13089);
xnor U16783 (N_16783,N_10050,N_14608);
and U16784 (N_16784,N_11421,N_12764);
nor U16785 (N_16785,N_10985,N_14308);
and U16786 (N_16786,N_13905,N_12472);
nand U16787 (N_16787,N_11583,N_11432);
nor U16788 (N_16788,N_11183,N_12714);
nor U16789 (N_16789,N_14856,N_11669);
or U16790 (N_16790,N_10130,N_14719);
nand U16791 (N_16791,N_12403,N_10534);
xor U16792 (N_16792,N_12190,N_14061);
xor U16793 (N_16793,N_13947,N_14393);
nor U16794 (N_16794,N_14718,N_10071);
and U16795 (N_16795,N_14351,N_14262);
nor U16796 (N_16796,N_12622,N_12289);
nand U16797 (N_16797,N_12242,N_14528);
and U16798 (N_16798,N_13137,N_14765);
and U16799 (N_16799,N_11285,N_14055);
nor U16800 (N_16800,N_13779,N_10948);
or U16801 (N_16801,N_13855,N_13359);
nor U16802 (N_16802,N_11284,N_12828);
or U16803 (N_16803,N_11322,N_13857);
xnor U16804 (N_16804,N_12558,N_14281);
nor U16805 (N_16805,N_12804,N_12887);
and U16806 (N_16806,N_13262,N_14950);
and U16807 (N_16807,N_10842,N_11410);
nand U16808 (N_16808,N_12215,N_13649);
nand U16809 (N_16809,N_10501,N_11620);
nand U16810 (N_16810,N_11034,N_10892);
xnor U16811 (N_16811,N_12864,N_10344);
nor U16812 (N_16812,N_11428,N_13189);
xor U16813 (N_16813,N_10134,N_11373);
xnor U16814 (N_16814,N_13883,N_11649);
and U16815 (N_16815,N_10398,N_13863);
nand U16816 (N_16816,N_11429,N_12587);
nand U16817 (N_16817,N_12909,N_11608);
and U16818 (N_16818,N_10949,N_11792);
nand U16819 (N_16819,N_13266,N_11564);
xor U16820 (N_16820,N_12562,N_13571);
or U16821 (N_16821,N_11599,N_10336);
nor U16822 (N_16822,N_13277,N_10091);
nand U16823 (N_16823,N_11881,N_12070);
xnor U16824 (N_16824,N_11375,N_13411);
xor U16825 (N_16825,N_10295,N_11434);
nor U16826 (N_16826,N_12519,N_12614);
xnor U16827 (N_16827,N_14838,N_11976);
xor U16828 (N_16828,N_12423,N_13893);
xnor U16829 (N_16829,N_12361,N_11400);
and U16830 (N_16830,N_10751,N_10831);
and U16831 (N_16831,N_12279,N_10575);
xor U16832 (N_16832,N_11381,N_10072);
or U16833 (N_16833,N_14639,N_10771);
nand U16834 (N_16834,N_11724,N_11084);
nand U16835 (N_16835,N_14969,N_14496);
nand U16836 (N_16836,N_10783,N_13630);
or U16837 (N_16837,N_13190,N_14118);
nand U16838 (N_16838,N_10357,N_12015);
nand U16839 (N_16839,N_14901,N_14222);
xor U16840 (N_16840,N_13489,N_14825);
xor U16841 (N_16841,N_14015,N_12788);
or U16842 (N_16842,N_14509,N_14860);
nor U16843 (N_16843,N_13508,N_14539);
and U16844 (N_16844,N_12551,N_12564);
xor U16845 (N_16845,N_12817,N_11378);
xor U16846 (N_16846,N_14360,N_14584);
or U16847 (N_16847,N_13029,N_11318);
and U16848 (N_16848,N_14692,N_13144);
and U16849 (N_16849,N_11505,N_10347);
and U16850 (N_16850,N_14791,N_11262);
nand U16851 (N_16851,N_13909,N_11833);
nand U16852 (N_16852,N_10599,N_10932);
nor U16853 (N_16853,N_14184,N_12657);
nand U16854 (N_16854,N_13233,N_14790);
or U16855 (N_16855,N_11648,N_12605);
nor U16856 (N_16856,N_11153,N_14268);
nand U16857 (N_16857,N_10494,N_12607);
nor U16858 (N_16858,N_14534,N_14266);
xor U16859 (N_16859,N_13328,N_11973);
nand U16860 (N_16860,N_13657,N_12487);
and U16861 (N_16861,N_10710,N_13236);
nand U16862 (N_16862,N_13984,N_13059);
nor U16863 (N_16863,N_12559,N_12217);
nand U16864 (N_16864,N_11259,N_14080);
or U16865 (N_16865,N_14559,N_14077);
nand U16866 (N_16866,N_12474,N_13753);
and U16867 (N_16867,N_13723,N_13369);
and U16868 (N_16868,N_10758,N_13408);
nor U16869 (N_16869,N_13527,N_13533);
nand U16870 (N_16870,N_12652,N_12697);
and U16871 (N_16871,N_13480,N_10593);
xor U16872 (N_16872,N_12450,N_10816);
or U16873 (N_16873,N_11621,N_10609);
nand U16874 (N_16874,N_14425,N_12514);
xnor U16875 (N_16875,N_12282,N_13164);
and U16876 (N_16876,N_10481,N_14537);
nor U16877 (N_16877,N_13267,N_11230);
nand U16878 (N_16878,N_12845,N_12469);
nor U16879 (N_16879,N_10641,N_14586);
nor U16880 (N_16880,N_13644,N_14473);
nor U16881 (N_16881,N_13574,N_13616);
or U16882 (N_16882,N_10224,N_10522);
and U16883 (N_16883,N_11701,N_11388);
xnor U16884 (N_16884,N_12695,N_11462);
nand U16885 (N_16885,N_11286,N_10793);
or U16886 (N_16886,N_10885,N_14189);
xor U16887 (N_16887,N_12676,N_10202);
nor U16888 (N_16888,N_10149,N_11987);
and U16889 (N_16889,N_11157,N_14561);
nand U16890 (N_16890,N_12849,N_10153);
or U16891 (N_16891,N_11287,N_11038);
and U16892 (N_16892,N_10557,N_14276);
nand U16893 (N_16893,N_10716,N_10092);
nand U16894 (N_16894,N_10857,N_12143);
and U16895 (N_16895,N_13542,N_10947);
nor U16896 (N_16896,N_13370,N_13282);
and U16897 (N_16897,N_14898,N_10470);
and U16898 (N_16898,N_10881,N_14154);
or U16899 (N_16899,N_14617,N_13650);
nand U16900 (N_16900,N_11777,N_10807);
or U16901 (N_16901,N_14669,N_12557);
nor U16902 (N_16902,N_12586,N_10737);
and U16903 (N_16903,N_12099,N_13213);
and U16904 (N_16904,N_10078,N_10998);
or U16905 (N_16905,N_13224,N_14249);
nor U16906 (N_16906,N_14943,N_13656);
and U16907 (N_16907,N_14926,N_14129);
nor U16908 (N_16908,N_14095,N_10965);
and U16909 (N_16909,N_13259,N_11613);
nand U16910 (N_16910,N_12928,N_13934);
nor U16911 (N_16911,N_11750,N_10940);
nor U16912 (N_16912,N_13203,N_13451);
nor U16913 (N_16913,N_12890,N_10084);
nor U16914 (N_16914,N_12425,N_11059);
xnor U16915 (N_16915,N_13078,N_14185);
and U16916 (N_16916,N_12277,N_14218);
xor U16917 (N_16917,N_13517,N_10172);
and U16918 (N_16918,N_11808,N_11491);
or U16919 (N_16919,N_12220,N_13106);
or U16920 (N_16920,N_14623,N_13974);
nand U16921 (N_16921,N_13895,N_10479);
or U16922 (N_16922,N_13941,N_10463);
nor U16923 (N_16923,N_10201,N_11658);
nor U16924 (N_16924,N_10647,N_11713);
nand U16925 (N_16925,N_12479,N_12322);
nand U16926 (N_16926,N_10176,N_12875);
and U16927 (N_16927,N_10147,N_14920);
nand U16928 (N_16928,N_12924,N_10392);
nor U16929 (N_16929,N_14529,N_13124);
xnor U16930 (N_16930,N_13181,N_11196);
xor U16931 (N_16931,N_14679,N_12295);
nand U16932 (N_16932,N_11536,N_14609);
nor U16933 (N_16933,N_14917,N_13628);
nor U16934 (N_16934,N_11681,N_12805);
nand U16935 (N_16935,N_12698,N_14030);
xnor U16936 (N_16936,N_11739,N_12567);
nor U16937 (N_16937,N_13513,N_14865);
nand U16938 (N_16938,N_12594,N_11699);
nor U16939 (N_16939,N_10178,N_10236);
and U16940 (N_16940,N_12046,N_13507);
and U16941 (N_16941,N_14314,N_10200);
nand U16942 (N_16942,N_14211,N_14572);
nand U16943 (N_16943,N_10893,N_10208);
nand U16944 (N_16944,N_11001,N_13011);
or U16945 (N_16945,N_14678,N_11764);
nor U16946 (N_16946,N_10636,N_12794);
or U16947 (N_16947,N_14652,N_11591);
or U16948 (N_16948,N_11145,N_12699);
and U16949 (N_16949,N_10526,N_14725);
and U16950 (N_16950,N_10047,N_10903);
xnor U16951 (N_16951,N_13986,N_11770);
and U16952 (N_16952,N_13070,N_12416);
and U16953 (N_16953,N_13671,N_12837);
nor U16954 (N_16954,N_11142,N_10266);
xnor U16955 (N_16955,N_11884,N_11249);
nand U16956 (N_16956,N_10449,N_13307);
nor U16957 (N_16957,N_13223,N_10165);
xnor U16958 (N_16958,N_12891,N_11609);
xnor U16959 (N_16959,N_12306,N_10386);
nand U16960 (N_16960,N_12827,N_11680);
or U16961 (N_16961,N_12484,N_10676);
nand U16962 (N_16962,N_13851,N_13066);
nor U16963 (N_16963,N_13146,N_14401);
xnor U16964 (N_16964,N_10810,N_12566);
or U16965 (N_16965,N_13488,N_13454);
nor U16966 (N_16966,N_11246,N_12911);
nand U16967 (N_16967,N_11288,N_13734);
nand U16968 (N_16968,N_12521,N_11586);
xnor U16969 (N_16969,N_13132,N_11908);
nor U16970 (N_16970,N_13825,N_14869);
and U16971 (N_16971,N_14862,N_12636);
or U16972 (N_16972,N_12033,N_14394);
nand U16973 (N_16973,N_14012,N_11939);
or U16974 (N_16974,N_11090,N_12119);
or U16975 (N_16975,N_12081,N_11377);
xor U16976 (N_16976,N_13051,N_13710);
nor U16977 (N_16977,N_11067,N_13686);
and U16978 (N_16978,N_10460,N_12777);
and U16979 (N_16979,N_13116,N_14404);
xor U16980 (N_16980,N_14413,N_10904);
nand U16981 (N_16981,N_12455,N_12383);
nand U16982 (N_16982,N_13086,N_10432);
nor U16983 (N_16983,N_14460,N_10804);
nand U16984 (N_16984,N_10081,N_12565);
or U16985 (N_16985,N_10777,N_13009);
nand U16986 (N_16986,N_11423,N_13759);
nor U16987 (N_16987,N_12139,N_12009);
or U16988 (N_16988,N_14066,N_13387);
or U16989 (N_16989,N_10513,N_11464);
and U16990 (N_16990,N_13849,N_11112);
and U16991 (N_16991,N_13667,N_11520);
nor U16992 (N_16992,N_13869,N_12655);
nor U16993 (N_16993,N_10044,N_10301);
and U16994 (N_16994,N_11359,N_14350);
or U16995 (N_16995,N_14851,N_10219);
nor U16996 (N_16996,N_12888,N_11159);
or U16997 (N_16997,N_11863,N_12389);
nand U16998 (N_16998,N_13027,N_12747);
or U16999 (N_16999,N_13035,N_14557);
xnor U17000 (N_17000,N_12426,N_14517);
or U17001 (N_17001,N_11243,N_12870);
and U17002 (N_17002,N_12688,N_14960);
or U17003 (N_17003,N_10510,N_13161);
xor U17004 (N_17004,N_10468,N_14696);
xnor U17005 (N_17005,N_12822,N_13930);
xnor U17006 (N_17006,N_13385,N_11233);
nand U17007 (N_17007,N_11969,N_12851);
nand U17008 (N_17008,N_12574,N_13890);
xnor U17009 (N_17009,N_14554,N_13452);
nand U17010 (N_17010,N_12112,N_12611);
nor U17011 (N_17011,N_14907,N_11748);
and U17012 (N_17012,N_12967,N_13415);
xnor U17013 (N_17013,N_10558,N_14313);
nor U17014 (N_17014,N_11450,N_12999);
nand U17015 (N_17015,N_14160,N_10406);
and U17016 (N_17016,N_12397,N_11424);
xor U17017 (N_17017,N_10585,N_10375);
and U17018 (N_17018,N_14587,N_11977);
xor U17019 (N_17019,N_13210,N_10251);
nand U17020 (N_17020,N_14051,N_12986);
or U17021 (N_17021,N_11205,N_11716);
nand U17022 (N_17022,N_10453,N_12757);
xnor U17023 (N_17023,N_13462,N_12428);
or U17024 (N_17024,N_14243,N_10248);
and U17025 (N_17025,N_12234,N_13470);
or U17026 (N_17026,N_13661,N_10656);
or U17027 (N_17027,N_13299,N_11229);
or U17028 (N_17028,N_10105,N_14053);
and U17029 (N_17029,N_13060,N_11522);
nand U17030 (N_17030,N_10784,N_13283);
or U17031 (N_17031,N_14610,N_11996);
xnor U17032 (N_17032,N_13354,N_12925);
nand U17033 (N_17033,N_12243,N_12726);
xor U17034 (N_17034,N_10424,N_14458);
nor U17035 (N_17035,N_13983,N_12960);
or U17036 (N_17036,N_10507,N_10369);
xnor U17037 (N_17037,N_11784,N_12561);
or U17038 (N_17038,N_13757,N_11094);
or U17039 (N_17039,N_14122,N_13398);
xor U17040 (N_17040,N_10877,N_11136);
nor U17041 (N_17041,N_11706,N_14876);
nor U17042 (N_17042,N_13153,N_13092);
nor U17043 (N_17043,N_14732,N_14701);
nor U17044 (N_17044,N_11111,N_12374);
nor U17045 (N_17045,N_10895,N_11337);
and U17046 (N_17046,N_11178,N_13526);
and U17047 (N_17047,N_12542,N_10556);
nand U17048 (N_17048,N_12661,N_12074);
xor U17049 (N_17049,N_11166,N_13737);
and U17050 (N_17050,N_12532,N_13430);
nand U17051 (N_17051,N_13353,N_14806);
nand U17052 (N_17052,N_13003,N_10671);
xnor U17053 (N_17053,N_11048,N_14546);
nand U17054 (N_17054,N_13043,N_13693);
or U17055 (N_17055,N_12623,N_13892);
or U17056 (N_17056,N_10376,N_12850);
and U17057 (N_17057,N_13955,N_14285);
nand U17058 (N_17058,N_11546,N_14735);
and U17059 (N_17059,N_10964,N_12427);
and U17060 (N_17060,N_12005,N_11309);
xor U17061 (N_17061,N_13606,N_12953);
nand U17062 (N_17062,N_13358,N_10325);
nand U17063 (N_17063,N_10822,N_13691);
and U17064 (N_17064,N_11104,N_14910);
xnor U17065 (N_17065,N_10702,N_11315);
and U17066 (N_17066,N_13774,N_12115);
and U17067 (N_17067,N_12492,N_13511);
nand U17068 (N_17068,N_11310,N_12742);
nand U17069 (N_17069,N_10423,N_11820);
or U17070 (N_17070,N_11986,N_11559);
and U17071 (N_17071,N_14121,N_10417);
and U17072 (N_17072,N_13653,N_12175);
xnor U17073 (N_17073,N_11439,N_14782);
or U17074 (N_17074,N_14050,N_13209);
xor U17075 (N_17075,N_13833,N_14773);
nor U17076 (N_17076,N_13700,N_14665);
or U17077 (N_17077,N_12808,N_12829);
nor U17078 (N_17078,N_10338,N_13296);
xnor U17079 (N_17079,N_13622,N_13742);
xnor U17080 (N_17080,N_11281,N_12581);
or U17081 (N_17081,N_13280,N_10897);
and U17082 (N_17082,N_12575,N_13005);
nor U17083 (N_17083,N_11240,N_12091);
nand U17084 (N_17084,N_12333,N_14255);
and U17085 (N_17085,N_14812,N_10966);
nor U17086 (N_17086,N_12991,N_11338);
or U17087 (N_17087,N_14035,N_14379);
and U17088 (N_17088,N_14841,N_13169);
and U17089 (N_17089,N_12316,N_12475);
nor U17090 (N_17090,N_11871,N_14944);
and U17091 (N_17091,N_10706,N_11678);
and U17092 (N_17092,N_11342,N_10661);
or U17093 (N_17093,N_12755,N_13543);
and U17094 (N_17094,N_10598,N_14405);
nor U17095 (N_17095,N_14594,N_11896);
xnor U17096 (N_17096,N_14018,N_13901);
and U17097 (N_17097,N_14219,N_13484);
nand U17098 (N_17098,N_13824,N_13538);
xnor U17099 (N_17099,N_13660,N_10196);
and U17100 (N_17100,N_12412,N_12368);
nand U17101 (N_17101,N_10797,N_11460);
nor U17102 (N_17102,N_10951,N_14315);
nand U17103 (N_17103,N_13914,N_10799);
xnor U17104 (N_17104,N_11630,N_12124);
nand U17105 (N_17105,N_10461,N_12568);
or U17106 (N_17106,N_10395,N_11185);
or U17107 (N_17107,N_11379,N_14805);
xor U17108 (N_17108,N_10538,N_12093);
nand U17109 (N_17109,N_14784,N_11913);
nand U17110 (N_17110,N_11728,N_13581);
nand U17111 (N_17111,N_11078,N_14463);
or U17112 (N_17112,N_12363,N_10190);
nand U17113 (N_17113,N_12332,N_10709);
nor U17114 (N_17114,N_14875,N_11858);
nand U17115 (N_17115,N_11387,N_12032);
or U17116 (N_17116,N_11244,N_11677);
or U17117 (N_17117,N_14312,N_10141);
or U17118 (N_17118,N_10955,N_11511);
nand U17119 (N_17119,N_11512,N_11925);
xor U17120 (N_17120,N_13635,N_12274);
or U17121 (N_17121,N_10762,N_12603);
and U17122 (N_17122,N_11663,N_10191);
and U17123 (N_17123,N_14143,N_13945);
and U17124 (N_17124,N_12366,N_14931);
xor U17125 (N_17125,N_11272,N_13397);
nor U17126 (N_17126,N_10352,N_13304);
or U17127 (N_17127,N_10629,N_11079);
nor U17128 (N_17128,N_11799,N_13772);
nor U17129 (N_17129,N_14327,N_10747);
or U17130 (N_17130,N_12126,N_12240);
xnor U17131 (N_17131,N_12585,N_11916);
xor U17132 (N_17132,N_14033,N_14435);
nand U17133 (N_17133,N_12945,N_14170);
and U17134 (N_17134,N_14126,N_13142);
or U17135 (N_17135,N_12513,N_11958);
or U17136 (N_17136,N_14767,N_14743);
or U17137 (N_17137,N_14778,N_11482);
or U17138 (N_17138,N_11771,N_10307);
nor U17139 (N_17139,N_14408,N_11778);
nand U17140 (N_17140,N_11889,N_14364);
and U17141 (N_17141,N_10872,N_13317);
xor U17142 (N_17142,N_13067,N_11736);
or U17143 (N_17143,N_12625,N_14193);
and U17144 (N_17144,N_12347,N_13179);
xnor U17145 (N_17145,N_10753,N_14682);
xnor U17146 (N_17146,N_13696,N_11876);
nor U17147 (N_17147,N_14982,N_13138);
nand U17148 (N_17148,N_12024,N_11861);
nand U17149 (N_17149,N_14074,N_13293);
nor U17150 (N_17150,N_10029,N_10007);
and U17151 (N_17151,N_12735,N_12780);
xnor U17152 (N_17152,N_11096,N_14157);
nand U17153 (N_17153,N_13324,N_10722);
and U17154 (N_17154,N_10351,N_10253);
xor U17155 (N_17155,N_10861,N_10562);
nor U17156 (N_17156,N_11027,N_10701);
and U17157 (N_17157,N_10829,N_12369);
and U17158 (N_17158,N_14419,N_11523);
nor U17159 (N_17159,N_14151,N_10143);
or U17160 (N_17160,N_10587,N_10967);
nor U17161 (N_17161,N_12022,N_14927);
xor U17162 (N_17162,N_12125,N_13782);
or U17163 (N_17163,N_10537,N_13104);
or U17164 (N_17164,N_10244,N_14503);
or U17165 (N_17165,N_14873,N_12765);
nor U17166 (N_17166,N_11758,N_13950);
nand U17167 (N_17167,N_12897,N_11108);
nor U17168 (N_17168,N_10140,N_10649);
nand U17169 (N_17169,N_11829,N_13112);
xor U17170 (N_17170,N_11527,N_13419);
nand U17171 (N_17171,N_14992,N_10594);
or U17172 (N_17172,N_11661,N_11502);
nor U17173 (N_17173,N_13001,N_13166);
xor U17174 (N_17174,N_14175,N_10591);
nor U17175 (N_17175,N_11856,N_11389);
nor U17176 (N_17176,N_14132,N_14240);
nand U17177 (N_17177,N_10512,N_10414);
xor U17178 (N_17178,N_11563,N_14432);
xnor U17179 (N_17179,N_12772,N_13922);
nor U17180 (N_17180,N_13633,N_13120);
and U17181 (N_17181,N_10606,N_11184);
xnor U17182 (N_17182,N_11070,N_11188);
nor U17183 (N_17183,N_10430,N_14912);
or U17184 (N_17184,N_10217,N_12618);
nand U17185 (N_17185,N_12791,N_14852);
and U17186 (N_17186,N_13738,N_10065);
nor U17187 (N_17187,N_11845,N_14999);
xor U17188 (N_17188,N_12885,N_11321);
nor U17189 (N_17189,N_12497,N_14264);
nand U17190 (N_17190,N_11569,N_13730);
and U17191 (N_17191,N_13850,N_10840);
nand U17192 (N_17192,N_12419,N_11509);
and U17193 (N_17193,N_13371,N_11590);
or U17194 (N_17194,N_14490,N_10059);
nor U17195 (N_17195,N_12651,N_12120);
nor U17196 (N_17196,N_12359,N_13272);
nand U17197 (N_17197,N_12984,N_11902);
xor U17198 (N_17198,N_10673,N_13642);
nand U17199 (N_17199,N_10853,N_12767);
and U17200 (N_17200,N_10073,N_13821);
xnor U17201 (N_17201,N_13379,N_11781);
and U17202 (N_17202,N_10354,N_13174);
and U17203 (N_17203,N_13443,N_14221);
xnor U17204 (N_17204,N_12087,N_14492);
nor U17205 (N_17205,N_14298,N_10025);
xnor U17206 (N_17206,N_12858,N_11478);
and U17207 (N_17207,N_14352,N_12392);
nor U17208 (N_17208,N_14942,N_11604);
nor U17209 (N_17209,N_11456,N_12257);
nor U17210 (N_17210,N_13085,N_11852);
or U17211 (N_17211,N_10552,N_10871);
nor U17212 (N_17212,N_10744,N_11574);
nand U17213 (N_17213,N_14165,N_11306);
xnor U17214 (N_17214,N_11413,N_10474);
and U17215 (N_17215,N_12919,N_11765);
nor U17216 (N_17216,N_13327,N_13618);
xnor U17217 (N_17217,N_14111,N_11133);
or U17218 (N_17218,N_11949,N_12507);
nand U17219 (N_17219,N_14809,N_10778);
xnor U17220 (N_17220,N_11504,N_10299);
or U17221 (N_17221,N_11667,N_14447);
or U17222 (N_17222,N_13077,N_10403);
xor U17223 (N_17223,N_13103,N_11907);
xnor U17224 (N_17224,N_13254,N_14316);
nand U17225 (N_17225,N_11602,N_13081);
nor U17226 (N_17226,N_14606,N_13839);
nor U17227 (N_17227,N_13122,N_14269);
nor U17228 (N_17228,N_10775,N_12576);
and U17229 (N_17229,N_11619,N_13838);
and U17230 (N_17230,N_12344,N_11148);
or U17231 (N_17231,N_10836,N_13469);
or U17232 (N_17232,N_11235,N_14005);
and U17233 (N_17233,N_10544,N_12016);
nand U17234 (N_17234,N_13754,N_10454);
or U17235 (N_17235,N_10038,N_10000);
nand U17236 (N_17236,N_10559,N_14573);
xor U17237 (N_17237,N_10256,N_12743);
and U17238 (N_17238,N_11831,N_12400);
or U17239 (N_17239,N_12442,N_10237);
nand U17240 (N_17240,N_10317,N_14311);
or U17241 (N_17241,N_12704,N_12367);
xnor U17242 (N_17242,N_12142,N_10734);
and U17243 (N_17243,N_10368,N_13681);
nor U17244 (N_17244,N_12734,N_12223);
or U17245 (N_17245,N_13271,N_14605);
xor U17246 (N_17246,N_12123,N_14959);
xnor U17247 (N_17247,N_12733,N_10854);
and U17248 (N_17248,N_14362,N_11975);
and U17249 (N_17249,N_10814,N_14558);
or U17250 (N_17250,N_10851,N_13414);
nor U17251 (N_17251,N_12812,N_13954);
nor U17252 (N_17252,N_10231,N_10476);
nor U17253 (N_17253,N_12149,N_14755);
xnor U17254 (N_17254,N_11595,N_13093);
and U17255 (N_17255,N_11497,N_13777);
xnor U17256 (N_17256,N_13025,N_11628);
or U17257 (N_17257,N_14845,N_10330);
nand U17258 (N_17258,N_10692,N_11869);
and U17259 (N_17259,N_11372,N_13704);
and U17260 (N_17260,N_11236,N_12252);
xnor U17261 (N_17261,N_10927,N_10163);
nand U17262 (N_17262,N_12555,N_11180);
xnor U17263 (N_17263,N_12023,N_11875);
nand U17264 (N_17264,N_13949,N_10005);
xor U17265 (N_17265,N_13891,N_10182);
and U17266 (N_17266,N_13466,N_12102);
xnor U17267 (N_17267,N_14409,N_13960);
nand U17268 (N_17268,N_13114,N_11295);
nor U17269 (N_17269,N_13399,N_11302);
nor U17270 (N_17270,N_10577,N_10259);
and U17271 (N_17271,N_14818,N_13599);
or U17272 (N_17272,N_14962,N_10003);
xnor U17273 (N_17273,N_10427,N_11062);
nand U17274 (N_17274,N_10032,N_11444);
nand U17275 (N_17275,N_12194,N_12291);
nor U17276 (N_17276,N_12760,N_14007);
nand U17277 (N_17277,N_12826,N_11360);
nand U17278 (N_17278,N_13747,N_10573);
nor U17279 (N_17279,N_11947,N_14820);
and U17280 (N_17280,N_11625,N_13529);
nand U17281 (N_17281,N_13790,N_14810);
and U17282 (N_17282,N_10235,N_13237);
xnor U17283 (N_17283,N_13564,N_12741);
or U17284 (N_17284,N_13937,N_12078);
and U17285 (N_17285,N_11960,N_14772);
nor U17286 (N_17286,N_14593,N_11571);
nand U17287 (N_17287,N_12198,N_11789);
and U17288 (N_17288,N_14891,N_12345);
xor U17289 (N_17289,N_11032,N_14465);
xnor U17290 (N_17290,N_13926,N_11679);
nand U17291 (N_17291,N_12825,N_10089);
nand U17292 (N_17292,N_12663,N_13897);
nand U17293 (N_17293,N_10225,N_14582);
or U17294 (N_17294,N_10107,N_14793);
xor U17295 (N_17295,N_12571,N_13744);
nor U17296 (N_17296,N_13110,N_14493);
and U17297 (N_17297,N_13163,N_11897);
nor U17298 (N_17298,N_11336,N_12975);
or U17299 (N_17299,N_12637,N_13305);
and U17300 (N_17300,N_13256,N_12962);
nand U17301 (N_17301,N_13659,N_11774);
nand U17302 (N_17302,N_13479,N_13562);
xnor U17303 (N_17303,N_11629,N_12601);
or U17304 (N_17304,N_12446,N_13596);
xnor U17305 (N_17305,N_14979,N_12833);
and U17306 (N_17306,N_10297,N_12680);
nor U17307 (N_17307,N_13368,N_12855);
nor U17308 (N_17308,N_12159,N_11222);
xor U17309 (N_17309,N_10664,N_10690);
and U17310 (N_17310,N_10581,N_11810);
xnor U17311 (N_17311,N_10124,N_10761);
and U17312 (N_17312,N_14058,N_13639);
and U17313 (N_17313,N_11797,N_13113);
nand U17314 (N_17314,N_12621,N_10770);
xor U17315 (N_17315,N_11999,N_14685);
or U17316 (N_17316,N_10099,N_13306);
xnor U17317 (N_17317,N_10142,N_14486);
nand U17318 (N_17318,N_13275,N_14216);
nand U17319 (N_17319,N_10654,N_10437);
and U17320 (N_17320,N_10255,N_10469);
nand U17321 (N_17321,N_14853,N_10331);
and U17322 (N_17322,N_14516,N_10511);
xnor U17323 (N_17323,N_13231,N_12643);
and U17324 (N_17324,N_12642,N_10693);
or U17325 (N_17325,N_14894,N_11846);
xnor U17326 (N_17326,N_13792,N_13968);
nor U17327 (N_17327,N_11035,N_14482);
nand U17328 (N_17328,N_10045,N_14048);
or U17329 (N_17329,N_14199,N_12375);
or U17330 (N_17330,N_12486,N_10745);
and U17331 (N_17331,N_14508,N_10919);
or U17332 (N_17332,N_13185,N_12004);
or U17333 (N_17333,N_10667,N_13418);
or U17334 (N_17334,N_14754,N_10874);
xor U17335 (N_17335,N_12457,N_13402);
nor U17336 (N_17336,N_14113,N_11769);
nor U17337 (N_17337,N_13940,N_10313);
nand U17338 (N_17338,N_12290,N_10518);
or U17339 (N_17339,N_13810,N_13647);
and U17340 (N_17340,N_14100,N_10968);
xor U17341 (N_17341,N_10438,N_12236);
nand U17342 (N_17342,N_12030,N_13902);
nand U17343 (N_17343,N_10502,N_10278);
nor U17344 (N_17344,N_14981,N_14236);
nor U17345 (N_17345,N_13918,N_12656);
xnor U17346 (N_17346,N_14530,N_12362);
xor U17347 (N_17347,N_13915,N_10436);
xnor U17348 (N_17348,N_11099,N_13229);
nand U17349 (N_17349,N_14140,N_14883);
xnor U17350 (N_17350,N_13819,N_10242);
xnor U17351 (N_17351,N_14713,N_10749);
and U17352 (N_17352,N_10074,N_12570);
nand U17353 (N_17353,N_14302,N_12186);
nand U17354 (N_17354,N_13394,N_11420);
nand U17355 (N_17355,N_12321,N_12756);
xnor U17356 (N_17356,N_11422,N_11443);
nor U17357 (N_17357,N_10055,N_10400);
nand U17358 (N_17358,N_10724,N_13165);
or U17359 (N_17359,N_11433,N_10497);
and U17360 (N_17360,N_13561,N_13755);
or U17361 (N_17361,N_10850,N_11470);
xnor U17362 (N_17362,N_11995,N_11779);
or U17363 (N_17363,N_11880,N_11616);
or U17364 (N_17364,N_11847,N_12577);
nand U17365 (N_17365,N_13302,N_11997);
nand U17366 (N_17366,N_11954,N_12847);
or U17367 (N_17367,N_13799,N_13823);
and U17368 (N_17368,N_14138,N_13456);
or U17369 (N_17369,N_12200,N_12670);
or U17370 (N_17370,N_13969,N_10194);
nor U17371 (N_17371,N_11650,N_13997);
nor U17372 (N_17372,N_10890,N_13310);
xor U17373 (N_17373,N_13655,N_12692);
or U17374 (N_17374,N_11668,N_13412);
xnor U17375 (N_17375,N_13265,N_14037);
xor U17376 (N_17376,N_11193,N_13173);
xor U17377 (N_17377,N_11787,N_13171);
nand U17378 (N_17378,N_12219,N_12580);
and U17379 (N_17379,N_11131,N_13687);
or U17380 (N_17380,N_10031,N_12933);
or U17381 (N_17381,N_14899,N_11021);
nand U17382 (N_17382,N_13540,N_12994);
nand U17383 (N_17383,N_14039,N_13000);
xor U17384 (N_17384,N_10033,N_11227);
or U17385 (N_17385,N_12191,N_12899);
xor U17386 (N_17386,N_11134,N_11391);
nand U17387 (N_17387,N_12275,N_14078);
nand U17388 (N_17388,N_14029,N_11867);
nor U17389 (N_17389,N_11932,N_14695);
nor U17390 (N_17390,N_10849,N_14330);
or U17391 (N_17391,N_14280,N_10241);
xnor U17392 (N_17392,N_10058,N_10590);
nand U17393 (N_17393,N_11303,N_13196);
xor U17394 (N_17394,N_12231,N_13427);
xnor U17395 (N_17395,N_10294,N_11043);
or U17396 (N_17396,N_14985,N_13600);
and U17397 (N_17397,N_12401,N_11225);
nor U17398 (N_17398,N_11042,N_12130);
xnor U17399 (N_17399,N_12157,N_10024);
nand U17400 (N_17400,N_12116,N_11836);
nand U17401 (N_17401,N_12592,N_14275);
nand U17402 (N_17402,N_13889,N_12096);
xor U17403 (N_17403,N_14799,N_10915);
or U17404 (N_17404,N_13560,N_13992);
or U17405 (N_17405,N_14646,N_10348);
and U17406 (N_17406,N_12681,N_10164);
xnor U17407 (N_17407,N_11477,N_10619);
or U17408 (N_17408,N_11879,N_14507);
or U17409 (N_17409,N_10388,N_12938);
xnor U17410 (N_17410,N_12716,N_13378);
nor U17411 (N_17411,N_14836,N_13587);
xor U17412 (N_17412,N_14758,N_14090);
or U17413 (N_17413,N_13910,N_12635);
xor U17414 (N_17414,N_14446,N_12169);
and U17415 (N_17415,N_10665,N_12171);
or U17416 (N_17416,N_10865,N_11943);
or U17417 (N_17417,N_13820,N_13295);
nand U17418 (N_17418,N_14973,N_11127);
or U17419 (N_17419,N_14385,N_14797);
nand U17420 (N_17420,N_14994,N_10858);
and U17421 (N_17421,N_10828,N_10794);
and U17422 (N_17422,N_11786,N_11253);
or U17423 (N_17423,N_13404,N_13985);
and U17424 (N_17424,N_11256,N_13724);
nor U17425 (N_17425,N_10260,N_14568);
or U17426 (N_17426,N_14382,N_12011);
xor U17427 (N_17427,N_10937,N_13040);
nor U17428 (N_17428,N_12085,N_11937);
xnor U17429 (N_17429,N_14704,N_13713);
and U17430 (N_17430,N_10727,N_12210);
nor U17431 (N_17431,N_12996,N_14402);
or U17432 (N_17432,N_12342,N_10062);
and U17433 (N_17433,N_14955,N_13510);
xnor U17434 (N_17434,N_11742,N_10366);
xnor U17435 (N_17435,N_12694,N_14983);
and U17436 (N_17436,N_11231,N_14212);
or U17437 (N_17437,N_12465,N_10841);
xnor U17438 (N_17438,N_12293,N_12270);
and U17439 (N_17439,N_14544,N_13018);
xnor U17440 (N_17440,N_11162,N_10335);
and U17441 (N_17441,N_12049,N_10614);
xnor U17442 (N_17442,N_11890,N_12466);
xor U17443 (N_17443,N_11666,N_14761);
xor U17444 (N_17444,N_10292,N_12433);
and U17445 (N_17445,N_14338,N_12241);
nand U17446 (N_17446,N_14545,N_13345);
xnor U17447 (N_17447,N_12421,N_11606);
nand U17448 (N_17448,N_13180,N_11260);
nand U17449 (N_17449,N_12518,N_10188);
nand U17450 (N_17450,N_13609,N_10679);
or U17451 (N_17451,N_13437,N_11304);
xor U17452 (N_17452,N_13746,N_13834);
nand U17453 (N_17453,N_11031,N_10063);
or U17454 (N_17454,N_13711,N_13607);
xnor U17455 (N_17455,N_14244,N_11783);
and U17456 (N_17456,N_12761,N_13494);
and U17457 (N_17457,N_10057,N_10269);
xnor U17458 (N_17458,N_11011,N_12786);
nor U17459 (N_17459,N_13563,N_14787);
and U17460 (N_17460,N_11118,N_13416);
xnor U17461 (N_17461,N_13337,N_14010);
nor U17462 (N_17462,N_14099,N_12418);
or U17463 (N_17463,N_12671,N_12090);
and U17464 (N_17464,N_13099,N_14340);
nand U17465 (N_17465,N_10042,N_12095);
nor U17466 (N_17466,N_11346,N_11992);
or U17467 (N_17467,N_12987,N_10900);
nand U17468 (N_17468,N_13870,N_11725);
nand U17469 (N_17469,N_11248,N_10314);
nor U17470 (N_17470,N_14096,N_14703);
nand U17471 (N_17471,N_11549,N_13439);
xnor U17472 (N_17472,N_11971,N_13631);
and U17473 (N_17473,N_14636,N_11953);
nor U17474 (N_17474,N_13680,N_11103);
nand U17475 (N_17475,N_10210,N_10001);
and U17476 (N_17476,N_12380,N_12776);
nand U17477 (N_17477,N_13386,N_12188);
nand U17478 (N_17478,N_12185,N_11703);
xor U17479 (N_17479,N_12413,N_10390);
nand U17480 (N_17480,N_13942,N_13867);
and U17481 (N_17481,N_12128,N_12793);
xnor U17482 (N_17482,N_11308,N_12673);
nor U17483 (N_17483,N_14475,N_10340);
xnor U17484 (N_17484,N_12163,N_11570);
nand U17485 (N_17485,N_11899,N_11068);
and U17486 (N_17486,N_14971,N_11745);
nand U17487 (N_17487,N_13752,N_11023);
nand U17488 (N_17488,N_14283,N_12254);
and U17489 (N_17489,N_10569,N_13133);
nor U17490 (N_17490,N_11263,N_11383);
nor U17491 (N_17491,N_10539,N_11533);
nor U17492 (N_17492,N_14297,N_14887);
and U17493 (N_17493,N_13455,N_13586);
or U17494 (N_17494,N_13101,N_11837);
nor U17495 (N_17495,N_13147,N_10789);
nor U17496 (N_17496,N_11743,N_14167);
or U17497 (N_17497,N_14923,N_12641);
or U17498 (N_17498,N_10312,N_12550);
nand U17499 (N_17499,N_11085,N_10239);
nand U17500 (N_17500,N_10215,N_11204);
nand U17501 (N_17501,N_11522,N_12277);
nor U17502 (N_17502,N_12356,N_13263);
and U17503 (N_17503,N_12483,N_11684);
nor U17504 (N_17504,N_11866,N_11138);
nand U17505 (N_17505,N_11988,N_13542);
nor U17506 (N_17506,N_11618,N_13176);
nand U17507 (N_17507,N_11036,N_13119);
nor U17508 (N_17508,N_13764,N_10175);
nor U17509 (N_17509,N_12548,N_13059);
nor U17510 (N_17510,N_10263,N_14992);
nor U17511 (N_17511,N_10926,N_14750);
nor U17512 (N_17512,N_12292,N_10724);
and U17513 (N_17513,N_13610,N_13570);
nor U17514 (N_17514,N_13596,N_11997);
and U17515 (N_17515,N_12442,N_11588);
nor U17516 (N_17516,N_12570,N_13723);
nand U17517 (N_17517,N_13509,N_12367);
nand U17518 (N_17518,N_14927,N_13992);
or U17519 (N_17519,N_13952,N_11582);
or U17520 (N_17520,N_11127,N_12544);
nand U17521 (N_17521,N_13240,N_13447);
nand U17522 (N_17522,N_10898,N_14166);
and U17523 (N_17523,N_12929,N_10262);
xnor U17524 (N_17524,N_10170,N_12302);
nand U17525 (N_17525,N_12401,N_14379);
xor U17526 (N_17526,N_14562,N_12570);
and U17527 (N_17527,N_14161,N_10140);
nand U17528 (N_17528,N_13018,N_14299);
xnor U17529 (N_17529,N_13827,N_11970);
xor U17530 (N_17530,N_13304,N_10883);
and U17531 (N_17531,N_12201,N_13149);
nor U17532 (N_17532,N_12583,N_13984);
xor U17533 (N_17533,N_12695,N_11018);
and U17534 (N_17534,N_10332,N_10187);
nor U17535 (N_17535,N_13179,N_12714);
nor U17536 (N_17536,N_12227,N_11874);
or U17537 (N_17537,N_10809,N_13127);
or U17538 (N_17538,N_10803,N_14336);
and U17539 (N_17539,N_10505,N_13201);
nand U17540 (N_17540,N_11968,N_10738);
or U17541 (N_17541,N_11248,N_13417);
xor U17542 (N_17542,N_14832,N_12530);
xor U17543 (N_17543,N_11275,N_12622);
xnor U17544 (N_17544,N_12342,N_10550);
or U17545 (N_17545,N_14250,N_10592);
and U17546 (N_17546,N_12172,N_10987);
nor U17547 (N_17547,N_12279,N_12848);
or U17548 (N_17548,N_14938,N_14528);
nand U17549 (N_17549,N_10916,N_11571);
nor U17550 (N_17550,N_13695,N_14558);
and U17551 (N_17551,N_13580,N_10319);
and U17552 (N_17552,N_14425,N_11275);
or U17553 (N_17553,N_14608,N_12539);
and U17554 (N_17554,N_13078,N_14326);
or U17555 (N_17555,N_12354,N_12654);
and U17556 (N_17556,N_11810,N_14765);
nand U17557 (N_17557,N_11997,N_11492);
xor U17558 (N_17558,N_11021,N_11503);
and U17559 (N_17559,N_12262,N_12477);
nor U17560 (N_17560,N_10584,N_12828);
nand U17561 (N_17561,N_12828,N_12655);
or U17562 (N_17562,N_10704,N_14599);
nand U17563 (N_17563,N_12282,N_14149);
and U17564 (N_17564,N_12738,N_14354);
and U17565 (N_17565,N_14489,N_13509);
xnor U17566 (N_17566,N_12395,N_14060);
nor U17567 (N_17567,N_13702,N_13443);
or U17568 (N_17568,N_12045,N_10733);
xnor U17569 (N_17569,N_13189,N_13467);
or U17570 (N_17570,N_14696,N_11220);
or U17571 (N_17571,N_13218,N_12302);
and U17572 (N_17572,N_13003,N_10723);
xnor U17573 (N_17573,N_11383,N_14684);
or U17574 (N_17574,N_10984,N_13351);
or U17575 (N_17575,N_12753,N_14155);
nand U17576 (N_17576,N_14783,N_13911);
and U17577 (N_17577,N_11567,N_11969);
and U17578 (N_17578,N_12586,N_11726);
or U17579 (N_17579,N_13414,N_12618);
nor U17580 (N_17580,N_10357,N_13292);
nor U17581 (N_17581,N_10049,N_13195);
nand U17582 (N_17582,N_12816,N_14035);
nand U17583 (N_17583,N_14157,N_13160);
or U17584 (N_17584,N_13782,N_14719);
nand U17585 (N_17585,N_11058,N_11265);
or U17586 (N_17586,N_13651,N_13044);
or U17587 (N_17587,N_13072,N_10557);
or U17588 (N_17588,N_14507,N_14102);
and U17589 (N_17589,N_14630,N_13685);
and U17590 (N_17590,N_13149,N_11334);
and U17591 (N_17591,N_13245,N_11872);
xnor U17592 (N_17592,N_13702,N_13828);
nand U17593 (N_17593,N_12023,N_10075);
nor U17594 (N_17594,N_11635,N_14075);
or U17595 (N_17595,N_14351,N_13616);
nand U17596 (N_17596,N_14608,N_12910);
xnor U17597 (N_17597,N_14490,N_14133);
or U17598 (N_17598,N_10673,N_11342);
nor U17599 (N_17599,N_11239,N_11534);
or U17600 (N_17600,N_10945,N_11863);
nor U17601 (N_17601,N_14411,N_12380);
nand U17602 (N_17602,N_10995,N_11369);
nor U17603 (N_17603,N_10911,N_10862);
xor U17604 (N_17604,N_12096,N_14748);
nand U17605 (N_17605,N_12831,N_13321);
nor U17606 (N_17606,N_11712,N_11835);
or U17607 (N_17607,N_13008,N_10964);
or U17608 (N_17608,N_14255,N_13121);
xor U17609 (N_17609,N_14282,N_12795);
xnor U17610 (N_17610,N_11558,N_11651);
xor U17611 (N_17611,N_11819,N_14240);
nand U17612 (N_17612,N_12029,N_11560);
nor U17613 (N_17613,N_14313,N_12091);
or U17614 (N_17614,N_12099,N_13985);
nand U17615 (N_17615,N_14144,N_14295);
nor U17616 (N_17616,N_11871,N_12788);
or U17617 (N_17617,N_12255,N_14691);
nor U17618 (N_17618,N_14308,N_14405);
and U17619 (N_17619,N_11816,N_12908);
nor U17620 (N_17620,N_11017,N_12583);
xnor U17621 (N_17621,N_11688,N_12788);
or U17622 (N_17622,N_14891,N_11399);
or U17623 (N_17623,N_11734,N_11954);
nor U17624 (N_17624,N_10132,N_14628);
nor U17625 (N_17625,N_14422,N_10720);
or U17626 (N_17626,N_14987,N_13502);
or U17627 (N_17627,N_11092,N_14792);
nand U17628 (N_17628,N_13392,N_10056);
or U17629 (N_17629,N_12126,N_11822);
xnor U17630 (N_17630,N_13724,N_11517);
and U17631 (N_17631,N_14017,N_12200);
nand U17632 (N_17632,N_12061,N_11157);
or U17633 (N_17633,N_14515,N_14348);
or U17634 (N_17634,N_14289,N_14137);
and U17635 (N_17635,N_12325,N_14457);
xor U17636 (N_17636,N_10886,N_13263);
xnor U17637 (N_17637,N_11053,N_11638);
or U17638 (N_17638,N_14602,N_11783);
nand U17639 (N_17639,N_13306,N_11445);
xnor U17640 (N_17640,N_13365,N_12318);
nor U17641 (N_17641,N_12794,N_13039);
and U17642 (N_17642,N_14508,N_10125);
xnor U17643 (N_17643,N_14542,N_10527);
nor U17644 (N_17644,N_12863,N_10710);
nor U17645 (N_17645,N_11122,N_12872);
nor U17646 (N_17646,N_12710,N_13956);
or U17647 (N_17647,N_14928,N_14664);
xnor U17648 (N_17648,N_14514,N_11924);
and U17649 (N_17649,N_14116,N_10913);
nor U17650 (N_17650,N_14682,N_12298);
xnor U17651 (N_17651,N_11670,N_10015);
nor U17652 (N_17652,N_12549,N_10396);
or U17653 (N_17653,N_10906,N_14045);
nand U17654 (N_17654,N_14277,N_13853);
nor U17655 (N_17655,N_14619,N_12827);
and U17656 (N_17656,N_14637,N_13398);
nor U17657 (N_17657,N_11103,N_13372);
xor U17658 (N_17658,N_13953,N_13489);
xor U17659 (N_17659,N_10352,N_14846);
or U17660 (N_17660,N_11150,N_14069);
nand U17661 (N_17661,N_14542,N_14641);
and U17662 (N_17662,N_13939,N_14875);
nor U17663 (N_17663,N_12200,N_11648);
or U17664 (N_17664,N_12293,N_12022);
and U17665 (N_17665,N_11612,N_10899);
nand U17666 (N_17666,N_12261,N_14074);
xnor U17667 (N_17667,N_12610,N_14254);
xor U17668 (N_17668,N_10063,N_13331);
or U17669 (N_17669,N_13137,N_10938);
xor U17670 (N_17670,N_14995,N_11754);
or U17671 (N_17671,N_10663,N_13193);
or U17672 (N_17672,N_11683,N_12326);
nor U17673 (N_17673,N_12380,N_13370);
or U17674 (N_17674,N_13296,N_11616);
nor U17675 (N_17675,N_11855,N_10818);
nand U17676 (N_17676,N_13328,N_14217);
xor U17677 (N_17677,N_11145,N_11081);
or U17678 (N_17678,N_12710,N_12197);
and U17679 (N_17679,N_11091,N_12890);
nor U17680 (N_17680,N_12308,N_12542);
nor U17681 (N_17681,N_10011,N_14085);
nor U17682 (N_17682,N_12411,N_11957);
or U17683 (N_17683,N_13463,N_11972);
and U17684 (N_17684,N_12686,N_13865);
nor U17685 (N_17685,N_14019,N_12171);
or U17686 (N_17686,N_11030,N_11614);
xor U17687 (N_17687,N_11734,N_13777);
or U17688 (N_17688,N_12118,N_10646);
and U17689 (N_17689,N_11630,N_11145);
nand U17690 (N_17690,N_11243,N_14700);
and U17691 (N_17691,N_11792,N_13018);
or U17692 (N_17692,N_11031,N_14623);
and U17693 (N_17693,N_10219,N_14506);
xor U17694 (N_17694,N_14701,N_12867);
nor U17695 (N_17695,N_12968,N_13775);
xnor U17696 (N_17696,N_11277,N_11364);
or U17697 (N_17697,N_10682,N_13397);
nand U17698 (N_17698,N_10856,N_12309);
nor U17699 (N_17699,N_10562,N_10490);
xnor U17700 (N_17700,N_13995,N_11727);
and U17701 (N_17701,N_10322,N_12108);
nor U17702 (N_17702,N_10567,N_12752);
or U17703 (N_17703,N_12336,N_10447);
nand U17704 (N_17704,N_14077,N_12602);
or U17705 (N_17705,N_14247,N_13758);
or U17706 (N_17706,N_10519,N_14827);
and U17707 (N_17707,N_14195,N_14213);
xnor U17708 (N_17708,N_10985,N_12688);
or U17709 (N_17709,N_12633,N_11726);
and U17710 (N_17710,N_10971,N_13680);
and U17711 (N_17711,N_11571,N_12613);
nor U17712 (N_17712,N_13929,N_11510);
nand U17713 (N_17713,N_14580,N_14195);
or U17714 (N_17714,N_10304,N_14928);
and U17715 (N_17715,N_14807,N_10610);
xnor U17716 (N_17716,N_12590,N_14763);
xor U17717 (N_17717,N_12935,N_10193);
nor U17718 (N_17718,N_12947,N_10320);
nor U17719 (N_17719,N_12302,N_10853);
xnor U17720 (N_17720,N_13558,N_14775);
or U17721 (N_17721,N_14658,N_12515);
nand U17722 (N_17722,N_14208,N_12539);
nor U17723 (N_17723,N_12351,N_14837);
or U17724 (N_17724,N_10769,N_12834);
or U17725 (N_17725,N_10770,N_13763);
and U17726 (N_17726,N_11016,N_13155);
xor U17727 (N_17727,N_14240,N_12931);
or U17728 (N_17728,N_10458,N_11369);
nand U17729 (N_17729,N_12630,N_11842);
nor U17730 (N_17730,N_12259,N_12323);
and U17731 (N_17731,N_11697,N_12041);
and U17732 (N_17732,N_12709,N_14719);
and U17733 (N_17733,N_14542,N_12210);
and U17734 (N_17734,N_10822,N_13223);
or U17735 (N_17735,N_10156,N_14900);
nor U17736 (N_17736,N_13307,N_13263);
and U17737 (N_17737,N_10160,N_12353);
nor U17738 (N_17738,N_12802,N_11176);
and U17739 (N_17739,N_12195,N_12995);
and U17740 (N_17740,N_10296,N_10381);
and U17741 (N_17741,N_13513,N_10488);
and U17742 (N_17742,N_10340,N_12031);
or U17743 (N_17743,N_14738,N_10920);
or U17744 (N_17744,N_11046,N_11124);
and U17745 (N_17745,N_12456,N_10759);
or U17746 (N_17746,N_10269,N_14592);
xor U17747 (N_17747,N_13537,N_10839);
nor U17748 (N_17748,N_14809,N_14573);
nor U17749 (N_17749,N_11939,N_10399);
and U17750 (N_17750,N_11721,N_14295);
and U17751 (N_17751,N_11022,N_10800);
xor U17752 (N_17752,N_12427,N_12717);
or U17753 (N_17753,N_11115,N_14436);
xnor U17754 (N_17754,N_13629,N_13837);
nor U17755 (N_17755,N_10164,N_13212);
nor U17756 (N_17756,N_11180,N_14719);
and U17757 (N_17757,N_14847,N_12776);
and U17758 (N_17758,N_14700,N_11967);
xor U17759 (N_17759,N_14560,N_10707);
nor U17760 (N_17760,N_10714,N_13535);
and U17761 (N_17761,N_14268,N_10260);
nor U17762 (N_17762,N_12149,N_10976);
or U17763 (N_17763,N_12880,N_11597);
or U17764 (N_17764,N_14496,N_13292);
nor U17765 (N_17765,N_13777,N_12331);
nand U17766 (N_17766,N_14982,N_12700);
nand U17767 (N_17767,N_12284,N_11576);
nand U17768 (N_17768,N_10183,N_14479);
xor U17769 (N_17769,N_10416,N_11391);
nor U17770 (N_17770,N_14416,N_10223);
or U17771 (N_17771,N_13238,N_12208);
nand U17772 (N_17772,N_11768,N_14413);
and U17773 (N_17773,N_13875,N_14894);
nor U17774 (N_17774,N_13744,N_12194);
or U17775 (N_17775,N_13390,N_12484);
xnor U17776 (N_17776,N_13967,N_11695);
nor U17777 (N_17777,N_12679,N_13876);
nand U17778 (N_17778,N_14657,N_14792);
or U17779 (N_17779,N_12852,N_12385);
nor U17780 (N_17780,N_10585,N_10343);
or U17781 (N_17781,N_10283,N_12636);
nor U17782 (N_17782,N_10721,N_13023);
nor U17783 (N_17783,N_11263,N_14219);
and U17784 (N_17784,N_13402,N_12869);
xnor U17785 (N_17785,N_14246,N_11397);
nor U17786 (N_17786,N_14232,N_10042);
xnor U17787 (N_17787,N_12410,N_12996);
or U17788 (N_17788,N_14429,N_11935);
nor U17789 (N_17789,N_13782,N_12790);
nor U17790 (N_17790,N_14191,N_13389);
nor U17791 (N_17791,N_12532,N_12392);
or U17792 (N_17792,N_13203,N_13124);
or U17793 (N_17793,N_10715,N_11312);
or U17794 (N_17794,N_11685,N_12288);
nor U17795 (N_17795,N_14746,N_11813);
nor U17796 (N_17796,N_10625,N_11830);
and U17797 (N_17797,N_11428,N_13112);
nand U17798 (N_17798,N_14477,N_11298);
and U17799 (N_17799,N_10563,N_13826);
nor U17800 (N_17800,N_13891,N_10645);
and U17801 (N_17801,N_11495,N_12469);
nor U17802 (N_17802,N_13886,N_14134);
xor U17803 (N_17803,N_10785,N_14422);
nand U17804 (N_17804,N_14342,N_10312);
or U17805 (N_17805,N_11116,N_14811);
xnor U17806 (N_17806,N_14869,N_10571);
nor U17807 (N_17807,N_13706,N_13553);
nand U17808 (N_17808,N_14155,N_11096);
or U17809 (N_17809,N_11196,N_13799);
nand U17810 (N_17810,N_12323,N_10940);
nor U17811 (N_17811,N_11270,N_10779);
or U17812 (N_17812,N_13281,N_13839);
nand U17813 (N_17813,N_11163,N_13045);
xnor U17814 (N_17814,N_14885,N_11981);
nor U17815 (N_17815,N_13985,N_13640);
and U17816 (N_17816,N_11751,N_14191);
nand U17817 (N_17817,N_11591,N_13034);
or U17818 (N_17818,N_14328,N_13869);
or U17819 (N_17819,N_11486,N_14357);
and U17820 (N_17820,N_12729,N_12245);
and U17821 (N_17821,N_14772,N_11921);
nand U17822 (N_17822,N_13523,N_10194);
and U17823 (N_17823,N_14807,N_14259);
nor U17824 (N_17824,N_12440,N_11067);
xor U17825 (N_17825,N_10203,N_11472);
and U17826 (N_17826,N_13962,N_13964);
xor U17827 (N_17827,N_11318,N_12837);
xnor U17828 (N_17828,N_12119,N_10146);
xor U17829 (N_17829,N_10254,N_12680);
xor U17830 (N_17830,N_10452,N_10617);
and U17831 (N_17831,N_13972,N_10601);
or U17832 (N_17832,N_14528,N_10228);
or U17833 (N_17833,N_14012,N_11900);
nand U17834 (N_17834,N_14951,N_14253);
nand U17835 (N_17835,N_10868,N_14876);
nand U17836 (N_17836,N_13427,N_12631);
nor U17837 (N_17837,N_13436,N_10173);
and U17838 (N_17838,N_12012,N_10835);
and U17839 (N_17839,N_14324,N_13843);
nor U17840 (N_17840,N_11345,N_12315);
and U17841 (N_17841,N_10357,N_12074);
xor U17842 (N_17842,N_13872,N_10937);
nand U17843 (N_17843,N_11635,N_10547);
nor U17844 (N_17844,N_11310,N_12613);
or U17845 (N_17845,N_12712,N_10637);
and U17846 (N_17846,N_12918,N_13522);
xnor U17847 (N_17847,N_10578,N_14029);
xor U17848 (N_17848,N_13858,N_13535);
or U17849 (N_17849,N_11035,N_11708);
or U17850 (N_17850,N_14866,N_11507);
xor U17851 (N_17851,N_12282,N_11171);
nand U17852 (N_17852,N_14442,N_10503);
and U17853 (N_17853,N_11128,N_14065);
and U17854 (N_17854,N_11867,N_11783);
nand U17855 (N_17855,N_12462,N_12276);
and U17856 (N_17856,N_10687,N_14576);
nand U17857 (N_17857,N_11602,N_13060);
nor U17858 (N_17858,N_12963,N_13918);
nor U17859 (N_17859,N_14839,N_10772);
nand U17860 (N_17860,N_11572,N_14272);
nand U17861 (N_17861,N_11304,N_11764);
nor U17862 (N_17862,N_13329,N_13148);
and U17863 (N_17863,N_12899,N_11767);
nor U17864 (N_17864,N_12634,N_11108);
nand U17865 (N_17865,N_12152,N_12338);
and U17866 (N_17866,N_10097,N_13311);
nand U17867 (N_17867,N_12549,N_12813);
nand U17868 (N_17868,N_11255,N_14441);
nor U17869 (N_17869,N_11856,N_13014);
or U17870 (N_17870,N_14490,N_11441);
nor U17871 (N_17871,N_14367,N_14182);
xor U17872 (N_17872,N_12479,N_10027);
or U17873 (N_17873,N_14516,N_13041);
nor U17874 (N_17874,N_10540,N_13196);
xor U17875 (N_17875,N_12691,N_14021);
and U17876 (N_17876,N_10713,N_13223);
nand U17877 (N_17877,N_10159,N_14367);
nor U17878 (N_17878,N_10531,N_11398);
nor U17879 (N_17879,N_13285,N_13268);
or U17880 (N_17880,N_14896,N_14327);
nand U17881 (N_17881,N_12238,N_14948);
nor U17882 (N_17882,N_13976,N_13350);
and U17883 (N_17883,N_11143,N_14524);
xor U17884 (N_17884,N_14099,N_14773);
nor U17885 (N_17885,N_13738,N_14516);
or U17886 (N_17886,N_12162,N_14597);
xnor U17887 (N_17887,N_13095,N_12223);
and U17888 (N_17888,N_10499,N_13959);
xor U17889 (N_17889,N_14446,N_12619);
or U17890 (N_17890,N_13994,N_13132);
nor U17891 (N_17891,N_11162,N_10880);
or U17892 (N_17892,N_10538,N_14153);
nand U17893 (N_17893,N_14225,N_14881);
xor U17894 (N_17894,N_14730,N_14173);
and U17895 (N_17895,N_13817,N_13641);
or U17896 (N_17896,N_12414,N_10040);
nand U17897 (N_17897,N_11794,N_12653);
or U17898 (N_17898,N_12183,N_13709);
nor U17899 (N_17899,N_12254,N_13933);
nor U17900 (N_17900,N_11681,N_11234);
or U17901 (N_17901,N_12088,N_11130);
nor U17902 (N_17902,N_14617,N_10574);
xor U17903 (N_17903,N_13875,N_14675);
and U17904 (N_17904,N_12538,N_12211);
nand U17905 (N_17905,N_11240,N_12085);
nor U17906 (N_17906,N_12512,N_12635);
nor U17907 (N_17907,N_12696,N_14884);
and U17908 (N_17908,N_12975,N_14767);
and U17909 (N_17909,N_10966,N_13062);
or U17910 (N_17910,N_11643,N_12792);
nor U17911 (N_17911,N_10946,N_10594);
and U17912 (N_17912,N_12553,N_12766);
or U17913 (N_17913,N_10002,N_11910);
and U17914 (N_17914,N_14460,N_13660);
or U17915 (N_17915,N_12586,N_12086);
or U17916 (N_17916,N_11412,N_14097);
xnor U17917 (N_17917,N_14748,N_12601);
and U17918 (N_17918,N_13679,N_13891);
nor U17919 (N_17919,N_10821,N_13850);
and U17920 (N_17920,N_10441,N_12880);
or U17921 (N_17921,N_12744,N_12949);
nor U17922 (N_17922,N_14019,N_12474);
nand U17923 (N_17923,N_14180,N_11936);
xnor U17924 (N_17924,N_11447,N_10368);
xor U17925 (N_17925,N_11322,N_14836);
nand U17926 (N_17926,N_13706,N_10006);
nand U17927 (N_17927,N_12199,N_13030);
xor U17928 (N_17928,N_14576,N_12299);
xor U17929 (N_17929,N_11114,N_14980);
nor U17930 (N_17930,N_13334,N_13640);
and U17931 (N_17931,N_11922,N_10554);
nor U17932 (N_17932,N_10603,N_10231);
and U17933 (N_17933,N_10182,N_14774);
nand U17934 (N_17934,N_13931,N_11455);
xnor U17935 (N_17935,N_12074,N_14278);
nor U17936 (N_17936,N_13513,N_11891);
or U17937 (N_17937,N_10510,N_13110);
nand U17938 (N_17938,N_12354,N_11943);
or U17939 (N_17939,N_13894,N_10455);
nand U17940 (N_17940,N_11461,N_12684);
or U17941 (N_17941,N_10549,N_11850);
nor U17942 (N_17942,N_13720,N_10893);
xor U17943 (N_17943,N_11408,N_11497);
nand U17944 (N_17944,N_12796,N_11284);
nor U17945 (N_17945,N_11573,N_11490);
xor U17946 (N_17946,N_13983,N_13830);
xor U17947 (N_17947,N_14975,N_11743);
nand U17948 (N_17948,N_10687,N_12855);
nor U17949 (N_17949,N_10181,N_12989);
xnor U17950 (N_17950,N_13313,N_13179);
or U17951 (N_17951,N_10445,N_11440);
or U17952 (N_17952,N_14613,N_10148);
nor U17953 (N_17953,N_14931,N_13059);
and U17954 (N_17954,N_10008,N_12361);
xnor U17955 (N_17955,N_11081,N_10425);
nor U17956 (N_17956,N_14326,N_13513);
xor U17957 (N_17957,N_14926,N_11066);
or U17958 (N_17958,N_12728,N_14782);
or U17959 (N_17959,N_11531,N_12955);
or U17960 (N_17960,N_13356,N_14324);
nor U17961 (N_17961,N_12820,N_13987);
nand U17962 (N_17962,N_14573,N_13282);
and U17963 (N_17963,N_14531,N_14134);
nor U17964 (N_17964,N_11425,N_11605);
nor U17965 (N_17965,N_11181,N_14701);
nor U17966 (N_17966,N_10586,N_11740);
nand U17967 (N_17967,N_12462,N_10114);
nand U17968 (N_17968,N_12491,N_14826);
nor U17969 (N_17969,N_12140,N_11068);
xor U17970 (N_17970,N_14562,N_14295);
nand U17971 (N_17971,N_10763,N_11189);
nor U17972 (N_17972,N_13070,N_11293);
nand U17973 (N_17973,N_12034,N_10128);
nor U17974 (N_17974,N_11760,N_13352);
nor U17975 (N_17975,N_14937,N_10729);
nand U17976 (N_17976,N_14202,N_11286);
nand U17977 (N_17977,N_13675,N_13255);
xnor U17978 (N_17978,N_10696,N_11904);
and U17979 (N_17979,N_12555,N_10691);
nor U17980 (N_17980,N_12116,N_12691);
and U17981 (N_17981,N_14602,N_14794);
nand U17982 (N_17982,N_11425,N_14274);
and U17983 (N_17983,N_10646,N_14805);
or U17984 (N_17984,N_13347,N_11923);
xor U17985 (N_17985,N_11540,N_11668);
and U17986 (N_17986,N_10774,N_10689);
xor U17987 (N_17987,N_14838,N_11941);
nand U17988 (N_17988,N_11897,N_14647);
xor U17989 (N_17989,N_12365,N_10406);
or U17990 (N_17990,N_14196,N_12724);
nand U17991 (N_17991,N_10799,N_10469);
nor U17992 (N_17992,N_13871,N_10962);
nand U17993 (N_17993,N_13232,N_12828);
xnor U17994 (N_17994,N_13151,N_12308);
and U17995 (N_17995,N_10217,N_10861);
nor U17996 (N_17996,N_10442,N_12760);
or U17997 (N_17997,N_13564,N_14932);
or U17998 (N_17998,N_13242,N_11713);
and U17999 (N_17999,N_11154,N_13497);
nor U18000 (N_18000,N_11915,N_10912);
nor U18001 (N_18001,N_10044,N_12092);
or U18002 (N_18002,N_14184,N_13784);
xor U18003 (N_18003,N_13153,N_14185);
or U18004 (N_18004,N_14314,N_11354);
xor U18005 (N_18005,N_10118,N_12515);
and U18006 (N_18006,N_13331,N_11122);
nor U18007 (N_18007,N_13508,N_11485);
or U18008 (N_18008,N_13979,N_12577);
nor U18009 (N_18009,N_13599,N_13041);
nand U18010 (N_18010,N_11676,N_14023);
xor U18011 (N_18011,N_10525,N_14396);
nand U18012 (N_18012,N_14902,N_12099);
or U18013 (N_18013,N_12123,N_13056);
and U18014 (N_18014,N_10184,N_11736);
nor U18015 (N_18015,N_10126,N_14959);
nor U18016 (N_18016,N_11083,N_10457);
nand U18017 (N_18017,N_13694,N_11826);
nand U18018 (N_18018,N_12852,N_12119);
nand U18019 (N_18019,N_11671,N_13408);
and U18020 (N_18020,N_11554,N_14199);
xnor U18021 (N_18021,N_13058,N_13893);
nand U18022 (N_18022,N_10630,N_14065);
nand U18023 (N_18023,N_13194,N_11102);
nor U18024 (N_18024,N_12440,N_11730);
nor U18025 (N_18025,N_11472,N_10397);
xor U18026 (N_18026,N_11003,N_10223);
nand U18027 (N_18027,N_10534,N_11549);
nand U18028 (N_18028,N_10698,N_12597);
xnor U18029 (N_18029,N_12900,N_11036);
nand U18030 (N_18030,N_14611,N_13027);
xnor U18031 (N_18031,N_13308,N_12492);
xnor U18032 (N_18032,N_10942,N_11143);
nand U18033 (N_18033,N_12520,N_11644);
nand U18034 (N_18034,N_14985,N_14979);
nor U18035 (N_18035,N_13530,N_12416);
xnor U18036 (N_18036,N_10120,N_10670);
nor U18037 (N_18037,N_14466,N_12282);
and U18038 (N_18038,N_11592,N_10355);
xor U18039 (N_18039,N_11678,N_13261);
and U18040 (N_18040,N_14302,N_11564);
or U18041 (N_18041,N_10385,N_14561);
nand U18042 (N_18042,N_12121,N_11833);
and U18043 (N_18043,N_10320,N_10153);
nand U18044 (N_18044,N_12961,N_10682);
xor U18045 (N_18045,N_13989,N_13343);
xor U18046 (N_18046,N_12579,N_13870);
and U18047 (N_18047,N_12959,N_14872);
or U18048 (N_18048,N_14256,N_11956);
nor U18049 (N_18049,N_10728,N_10453);
nor U18050 (N_18050,N_10425,N_14472);
nor U18051 (N_18051,N_14877,N_11221);
xnor U18052 (N_18052,N_10076,N_13292);
nand U18053 (N_18053,N_11493,N_11810);
or U18054 (N_18054,N_11988,N_11807);
xnor U18055 (N_18055,N_11588,N_13515);
nor U18056 (N_18056,N_14337,N_14003);
or U18057 (N_18057,N_11050,N_12788);
and U18058 (N_18058,N_14794,N_12522);
xnor U18059 (N_18059,N_13473,N_12399);
nand U18060 (N_18060,N_11768,N_10873);
xnor U18061 (N_18061,N_14742,N_10301);
nor U18062 (N_18062,N_11915,N_13368);
nor U18063 (N_18063,N_14319,N_14414);
nand U18064 (N_18064,N_10957,N_11981);
xnor U18065 (N_18065,N_11657,N_11121);
nor U18066 (N_18066,N_10853,N_10834);
nand U18067 (N_18067,N_13862,N_13977);
nor U18068 (N_18068,N_12148,N_11571);
nand U18069 (N_18069,N_10510,N_14202);
and U18070 (N_18070,N_14535,N_14030);
or U18071 (N_18071,N_13215,N_13268);
nor U18072 (N_18072,N_13528,N_13414);
nor U18073 (N_18073,N_13355,N_12497);
nor U18074 (N_18074,N_14330,N_12989);
and U18075 (N_18075,N_14966,N_14545);
xor U18076 (N_18076,N_11841,N_13938);
nor U18077 (N_18077,N_13398,N_10702);
nand U18078 (N_18078,N_13627,N_13992);
nand U18079 (N_18079,N_12819,N_12452);
nor U18080 (N_18080,N_10645,N_11636);
and U18081 (N_18081,N_11942,N_10625);
or U18082 (N_18082,N_10385,N_14835);
or U18083 (N_18083,N_14547,N_12539);
nor U18084 (N_18084,N_13507,N_13492);
nand U18085 (N_18085,N_13256,N_14496);
xnor U18086 (N_18086,N_11331,N_14766);
nor U18087 (N_18087,N_14867,N_14559);
nor U18088 (N_18088,N_10326,N_11650);
nor U18089 (N_18089,N_11324,N_11276);
nand U18090 (N_18090,N_11214,N_12826);
and U18091 (N_18091,N_10208,N_11705);
and U18092 (N_18092,N_11717,N_13874);
nor U18093 (N_18093,N_12372,N_12929);
and U18094 (N_18094,N_14399,N_12473);
and U18095 (N_18095,N_14745,N_12255);
nand U18096 (N_18096,N_11171,N_10106);
or U18097 (N_18097,N_13634,N_12946);
xor U18098 (N_18098,N_13128,N_14445);
xnor U18099 (N_18099,N_13194,N_14469);
and U18100 (N_18100,N_10378,N_13857);
and U18101 (N_18101,N_11139,N_14845);
nand U18102 (N_18102,N_14507,N_14739);
nand U18103 (N_18103,N_13641,N_11714);
nand U18104 (N_18104,N_14901,N_11477);
nand U18105 (N_18105,N_11757,N_12166);
nand U18106 (N_18106,N_14383,N_12052);
or U18107 (N_18107,N_11591,N_12864);
and U18108 (N_18108,N_14580,N_10045);
nor U18109 (N_18109,N_11340,N_12205);
xnor U18110 (N_18110,N_10927,N_13568);
nand U18111 (N_18111,N_12168,N_11338);
nor U18112 (N_18112,N_13712,N_10317);
nand U18113 (N_18113,N_10352,N_11995);
nor U18114 (N_18114,N_14063,N_13611);
and U18115 (N_18115,N_11227,N_11259);
nand U18116 (N_18116,N_13181,N_11055);
or U18117 (N_18117,N_12518,N_10674);
or U18118 (N_18118,N_11414,N_12709);
xor U18119 (N_18119,N_13326,N_13744);
or U18120 (N_18120,N_11800,N_13551);
or U18121 (N_18121,N_13793,N_11117);
or U18122 (N_18122,N_11855,N_13291);
nor U18123 (N_18123,N_13263,N_11873);
or U18124 (N_18124,N_10483,N_10797);
and U18125 (N_18125,N_11368,N_13157);
and U18126 (N_18126,N_10261,N_10154);
or U18127 (N_18127,N_12402,N_14167);
or U18128 (N_18128,N_14026,N_10092);
nand U18129 (N_18129,N_13625,N_13583);
or U18130 (N_18130,N_14908,N_10188);
and U18131 (N_18131,N_11199,N_14387);
xor U18132 (N_18132,N_11294,N_14298);
xor U18133 (N_18133,N_11479,N_14248);
nand U18134 (N_18134,N_14099,N_10732);
xor U18135 (N_18135,N_10129,N_14760);
nor U18136 (N_18136,N_13832,N_10928);
nand U18137 (N_18137,N_13031,N_13748);
xnor U18138 (N_18138,N_14274,N_10455);
nor U18139 (N_18139,N_12880,N_13240);
xor U18140 (N_18140,N_10252,N_10000);
and U18141 (N_18141,N_13176,N_13608);
nor U18142 (N_18142,N_13945,N_10912);
nor U18143 (N_18143,N_10045,N_12061);
nand U18144 (N_18144,N_14431,N_12941);
nor U18145 (N_18145,N_14524,N_12824);
xnor U18146 (N_18146,N_14590,N_14324);
nand U18147 (N_18147,N_13952,N_10593);
nand U18148 (N_18148,N_12212,N_10497);
and U18149 (N_18149,N_14296,N_11317);
xnor U18150 (N_18150,N_11432,N_10280);
nor U18151 (N_18151,N_11389,N_13087);
nor U18152 (N_18152,N_14684,N_11285);
or U18153 (N_18153,N_12147,N_13305);
xnor U18154 (N_18154,N_13434,N_11500);
nand U18155 (N_18155,N_14107,N_10412);
and U18156 (N_18156,N_14736,N_10162);
and U18157 (N_18157,N_11494,N_12796);
nor U18158 (N_18158,N_14390,N_12157);
xnor U18159 (N_18159,N_14726,N_10153);
and U18160 (N_18160,N_12725,N_11561);
xor U18161 (N_18161,N_14948,N_10368);
and U18162 (N_18162,N_14957,N_13858);
or U18163 (N_18163,N_10779,N_10166);
nand U18164 (N_18164,N_13018,N_10956);
xor U18165 (N_18165,N_14900,N_12701);
nand U18166 (N_18166,N_10736,N_13115);
nand U18167 (N_18167,N_13583,N_13808);
or U18168 (N_18168,N_14490,N_10549);
xnor U18169 (N_18169,N_13703,N_12065);
xnor U18170 (N_18170,N_11759,N_13258);
or U18171 (N_18171,N_14737,N_12700);
nor U18172 (N_18172,N_13240,N_12904);
and U18173 (N_18173,N_11298,N_13976);
and U18174 (N_18174,N_11691,N_14902);
nor U18175 (N_18175,N_10909,N_10545);
xnor U18176 (N_18176,N_10493,N_12663);
or U18177 (N_18177,N_14261,N_14635);
xnor U18178 (N_18178,N_11659,N_14274);
nand U18179 (N_18179,N_11707,N_10739);
or U18180 (N_18180,N_12475,N_12653);
and U18181 (N_18181,N_14210,N_10305);
nand U18182 (N_18182,N_14501,N_14727);
and U18183 (N_18183,N_10022,N_10884);
xor U18184 (N_18184,N_12730,N_12390);
xnor U18185 (N_18185,N_14818,N_13329);
and U18186 (N_18186,N_12076,N_12843);
xor U18187 (N_18187,N_12126,N_11194);
or U18188 (N_18188,N_10520,N_10892);
or U18189 (N_18189,N_10829,N_11482);
and U18190 (N_18190,N_10350,N_10080);
xor U18191 (N_18191,N_11982,N_12375);
nor U18192 (N_18192,N_11453,N_11041);
or U18193 (N_18193,N_12308,N_13568);
or U18194 (N_18194,N_12363,N_11419);
and U18195 (N_18195,N_11841,N_10985);
and U18196 (N_18196,N_12930,N_11630);
and U18197 (N_18197,N_10569,N_11451);
xnor U18198 (N_18198,N_11098,N_13665);
or U18199 (N_18199,N_11993,N_10892);
nor U18200 (N_18200,N_12908,N_14361);
xnor U18201 (N_18201,N_10818,N_14116);
xnor U18202 (N_18202,N_10741,N_13562);
nand U18203 (N_18203,N_11103,N_12165);
nand U18204 (N_18204,N_12601,N_13055);
xnor U18205 (N_18205,N_14634,N_14023);
or U18206 (N_18206,N_13338,N_12977);
xor U18207 (N_18207,N_13172,N_14538);
xnor U18208 (N_18208,N_12425,N_14770);
xnor U18209 (N_18209,N_10045,N_14634);
or U18210 (N_18210,N_13111,N_14173);
nor U18211 (N_18211,N_10596,N_10321);
nor U18212 (N_18212,N_12193,N_14675);
nor U18213 (N_18213,N_10630,N_12752);
or U18214 (N_18214,N_13116,N_14588);
nand U18215 (N_18215,N_13374,N_14294);
xnor U18216 (N_18216,N_12238,N_14509);
or U18217 (N_18217,N_13766,N_14269);
nor U18218 (N_18218,N_11856,N_12299);
or U18219 (N_18219,N_12844,N_11354);
and U18220 (N_18220,N_10773,N_11941);
or U18221 (N_18221,N_10505,N_12671);
or U18222 (N_18222,N_10594,N_11952);
xor U18223 (N_18223,N_13394,N_10417);
and U18224 (N_18224,N_11971,N_11114);
and U18225 (N_18225,N_11507,N_13207);
nand U18226 (N_18226,N_11621,N_13088);
xor U18227 (N_18227,N_11381,N_11854);
nor U18228 (N_18228,N_11717,N_14174);
or U18229 (N_18229,N_12586,N_13808);
or U18230 (N_18230,N_13274,N_12222);
or U18231 (N_18231,N_10359,N_11889);
and U18232 (N_18232,N_11434,N_12708);
or U18233 (N_18233,N_11451,N_11683);
or U18234 (N_18234,N_13353,N_12458);
nor U18235 (N_18235,N_11465,N_13656);
or U18236 (N_18236,N_11133,N_13633);
nand U18237 (N_18237,N_14764,N_14588);
nand U18238 (N_18238,N_10693,N_14967);
nand U18239 (N_18239,N_12563,N_10949);
xor U18240 (N_18240,N_13924,N_10673);
and U18241 (N_18241,N_12170,N_13471);
and U18242 (N_18242,N_13455,N_10098);
nand U18243 (N_18243,N_10729,N_11871);
nor U18244 (N_18244,N_14593,N_14339);
and U18245 (N_18245,N_10426,N_14419);
or U18246 (N_18246,N_14112,N_12282);
and U18247 (N_18247,N_10913,N_14605);
xnor U18248 (N_18248,N_10720,N_13963);
and U18249 (N_18249,N_14521,N_13531);
xor U18250 (N_18250,N_11188,N_12450);
nor U18251 (N_18251,N_13710,N_11399);
xnor U18252 (N_18252,N_11642,N_13263);
xnor U18253 (N_18253,N_10862,N_12297);
and U18254 (N_18254,N_11650,N_12233);
nor U18255 (N_18255,N_13429,N_10282);
or U18256 (N_18256,N_11065,N_12625);
and U18257 (N_18257,N_11822,N_12573);
xnor U18258 (N_18258,N_11152,N_12737);
and U18259 (N_18259,N_11291,N_13328);
or U18260 (N_18260,N_14078,N_13073);
nand U18261 (N_18261,N_10078,N_13326);
nand U18262 (N_18262,N_13495,N_11661);
xnor U18263 (N_18263,N_12326,N_12344);
nand U18264 (N_18264,N_14087,N_11774);
and U18265 (N_18265,N_11370,N_10623);
xor U18266 (N_18266,N_11526,N_12870);
and U18267 (N_18267,N_14693,N_11629);
or U18268 (N_18268,N_11527,N_12643);
nand U18269 (N_18269,N_14288,N_10957);
xnor U18270 (N_18270,N_14147,N_12127);
nand U18271 (N_18271,N_11773,N_11749);
nand U18272 (N_18272,N_13469,N_13523);
and U18273 (N_18273,N_13699,N_12020);
nand U18274 (N_18274,N_11992,N_13303);
or U18275 (N_18275,N_14069,N_14750);
xor U18276 (N_18276,N_10551,N_11438);
nor U18277 (N_18277,N_14754,N_13804);
nand U18278 (N_18278,N_14570,N_14032);
or U18279 (N_18279,N_13691,N_10943);
or U18280 (N_18280,N_14712,N_13582);
nor U18281 (N_18281,N_13412,N_14479);
xnor U18282 (N_18282,N_11421,N_12264);
nand U18283 (N_18283,N_11187,N_12911);
nand U18284 (N_18284,N_14395,N_10583);
and U18285 (N_18285,N_14301,N_14466);
xor U18286 (N_18286,N_12115,N_14163);
xor U18287 (N_18287,N_14455,N_14217);
nand U18288 (N_18288,N_10701,N_10055);
nand U18289 (N_18289,N_13552,N_14645);
or U18290 (N_18290,N_14871,N_11797);
nand U18291 (N_18291,N_10930,N_10270);
and U18292 (N_18292,N_12184,N_11960);
nand U18293 (N_18293,N_11776,N_12700);
and U18294 (N_18294,N_14967,N_14665);
nand U18295 (N_18295,N_10380,N_14748);
and U18296 (N_18296,N_13295,N_11801);
xnor U18297 (N_18297,N_12115,N_12414);
nor U18298 (N_18298,N_12384,N_12019);
xor U18299 (N_18299,N_12407,N_11030);
nand U18300 (N_18300,N_12530,N_12496);
nor U18301 (N_18301,N_14854,N_14948);
or U18302 (N_18302,N_14050,N_13217);
and U18303 (N_18303,N_14278,N_12735);
nor U18304 (N_18304,N_10892,N_10051);
and U18305 (N_18305,N_13616,N_13337);
or U18306 (N_18306,N_12343,N_14807);
nand U18307 (N_18307,N_11464,N_14383);
and U18308 (N_18308,N_12040,N_10810);
and U18309 (N_18309,N_14954,N_13635);
and U18310 (N_18310,N_11440,N_12305);
nor U18311 (N_18311,N_11976,N_14971);
or U18312 (N_18312,N_12075,N_10548);
xor U18313 (N_18313,N_11657,N_13409);
nand U18314 (N_18314,N_11168,N_10214);
xor U18315 (N_18315,N_14764,N_13844);
and U18316 (N_18316,N_14200,N_13438);
or U18317 (N_18317,N_11019,N_11759);
xnor U18318 (N_18318,N_11515,N_10526);
or U18319 (N_18319,N_14292,N_12320);
and U18320 (N_18320,N_11345,N_14345);
and U18321 (N_18321,N_11840,N_13044);
xor U18322 (N_18322,N_12558,N_13081);
xor U18323 (N_18323,N_14726,N_11741);
nand U18324 (N_18324,N_14025,N_10098);
or U18325 (N_18325,N_14277,N_14575);
nand U18326 (N_18326,N_11659,N_11471);
nand U18327 (N_18327,N_10386,N_12261);
nand U18328 (N_18328,N_11759,N_13688);
nor U18329 (N_18329,N_14968,N_11158);
and U18330 (N_18330,N_12907,N_12521);
xnor U18331 (N_18331,N_12158,N_10191);
or U18332 (N_18332,N_11765,N_14325);
and U18333 (N_18333,N_11287,N_12801);
xor U18334 (N_18334,N_10824,N_10208);
or U18335 (N_18335,N_10800,N_13826);
and U18336 (N_18336,N_13583,N_13187);
nand U18337 (N_18337,N_11589,N_11490);
xor U18338 (N_18338,N_10651,N_13568);
or U18339 (N_18339,N_11986,N_11364);
nand U18340 (N_18340,N_12347,N_14741);
or U18341 (N_18341,N_12384,N_10555);
and U18342 (N_18342,N_14588,N_11232);
nor U18343 (N_18343,N_13576,N_11406);
nand U18344 (N_18344,N_10742,N_12615);
or U18345 (N_18345,N_12885,N_11109);
or U18346 (N_18346,N_11944,N_12330);
and U18347 (N_18347,N_12402,N_13419);
and U18348 (N_18348,N_10020,N_12954);
or U18349 (N_18349,N_11998,N_14848);
and U18350 (N_18350,N_12308,N_13994);
xnor U18351 (N_18351,N_10648,N_10573);
nand U18352 (N_18352,N_13215,N_11752);
nand U18353 (N_18353,N_10893,N_11328);
and U18354 (N_18354,N_10578,N_10946);
and U18355 (N_18355,N_13779,N_11277);
and U18356 (N_18356,N_12068,N_10305);
and U18357 (N_18357,N_13571,N_14246);
xnor U18358 (N_18358,N_11984,N_13331);
and U18359 (N_18359,N_11765,N_11800);
xor U18360 (N_18360,N_13017,N_13160);
or U18361 (N_18361,N_12597,N_14967);
or U18362 (N_18362,N_14022,N_10450);
nand U18363 (N_18363,N_11385,N_10662);
nand U18364 (N_18364,N_12439,N_10200);
or U18365 (N_18365,N_10655,N_13493);
nand U18366 (N_18366,N_13901,N_13246);
and U18367 (N_18367,N_13457,N_13530);
and U18368 (N_18368,N_13452,N_12604);
or U18369 (N_18369,N_13309,N_10402);
or U18370 (N_18370,N_14098,N_13598);
and U18371 (N_18371,N_13060,N_12938);
and U18372 (N_18372,N_12094,N_14293);
xor U18373 (N_18373,N_12332,N_12595);
and U18374 (N_18374,N_14024,N_13492);
or U18375 (N_18375,N_13373,N_14778);
nand U18376 (N_18376,N_12338,N_11499);
nand U18377 (N_18377,N_13529,N_10254);
xor U18378 (N_18378,N_12525,N_12610);
xnor U18379 (N_18379,N_14374,N_12195);
or U18380 (N_18380,N_10845,N_10057);
xor U18381 (N_18381,N_12312,N_10758);
nor U18382 (N_18382,N_11996,N_13053);
xnor U18383 (N_18383,N_12506,N_12098);
xnor U18384 (N_18384,N_12556,N_11019);
or U18385 (N_18385,N_14303,N_12372);
or U18386 (N_18386,N_13029,N_12007);
nand U18387 (N_18387,N_13059,N_12625);
nand U18388 (N_18388,N_13449,N_14010);
nand U18389 (N_18389,N_12543,N_11744);
xnor U18390 (N_18390,N_10009,N_12460);
nor U18391 (N_18391,N_12875,N_12221);
nor U18392 (N_18392,N_14005,N_10693);
xor U18393 (N_18393,N_14939,N_11205);
or U18394 (N_18394,N_12109,N_10855);
nand U18395 (N_18395,N_10166,N_13531);
or U18396 (N_18396,N_13748,N_12701);
nand U18397 (N_18397,N_10588,N_12193);
nor U18398 (N_18398,N_12086,N_12542);
nor U18399 (N_18399,N_13231,N_12204);
nand U18400 (N_18400,N_10915,N_14353);
nor U18401 (N_18401,N_10999,N_12475);
nand U18402 (N_18402,N_11172,N_13057);
nor U18403 (N_18403,N_10456,N_11283);
and U18404 (N_18404,N_13891,N_12595);
or U18405 (N_18405,N_11058,N_10144);
nand U18406 (N_18406,N_13536,N_11269);
or U18407 (N_18407,N_14850,N_13517);
xor U18408 (N_18408,N_11176,N_11780);
xnor U18409 (N_18409,N_11505,N_12140);
or U18410 (N_18410,N_10077,N_10440);
and U18411 (N_18411,N_11346,N_14114);
nor U18412 (N_18412,N_13125,N_11014);
xor U18413 (N_18413,N_11747,N_10786);
or U18414 (N_18414,N_10869,N_12239);
and U18415 (N_18415,N_11846,N_13572);
nand U18416 (N_18416,N_11664,N_11790);
nand U18417 (N_18417,N_11532,N_10613);
or U18418 (N_18418,N_11687,N_11814);
and U18419 (N_18419,N_12021,N_11757);
xor U18420 (N_18420,N_11539,N_14070);
nand U18421 (N_18421,N_10416,N_12752);
xor U18422 (N_18422,N_14668,N_11288);
or U18423 (N_18423,N_14740,N_11107);
xnor U18424 (N_18424,N_11004,N_13278);
nand U18425 (N_18425,N_12575,N_12562);
and U18426 (N_18426,N_12771,N_11447);
nand U18427 (N_18427,N_13385,N_14609);
or U18428 (N_18428,N_14752,N_11034);
or U18429 (N_18429,N_11474,N_10451);
nand U18430 (N_18430,N_12874,N_14546);
xor U18431 (N_18431,N_10356,N_10408);
xnor U18432 (N_18432,N_11829,N_14043);
and U18433 (N_18433,N_12339,N_12660);
or U18434 (N_18434,N_14564,N_14236);
or U18435 (N_18435,N_13003,N_10383);
nor U18436 (N_18436,N_10103,N_14516);
nand U18437 (N_18437,N_12278,N_12779);
and U18438 (N_18438,N_10868,N_11769);
xnor U18439 (N_18439,N_14086,N_14944);
nand U18440 (N_18440,N_12704,N_13022);
nand U18441 (N_18441,N_14551,N_10921);
or U18442 (N_18442,N_12849,N_10324);
or U18443 (N_18443,N_14131,N_13636);
or U18444 (N_18444,N_14520,N_11994);
or U18445 (N_18445,N_12523,N_14265);
and U18446 (N_18446,N_12361,N_11799);
xnor U18447 (N_18447,N_13315,N_13208);
nor U18448 (N_18448,N_12055,N_14470);
nand U18449 (N_18449,N_11588,N_12198);
nor U18450 (N_18450,N_12707,N_14662);
xnor U18451 (N_18451,N_14786,N_11733);
nor U18452 (N_18452,N_12254,N_11279);
or U18453 (N_18453,N_10219,N_10599);
nand U18454 (N_18454,N_13475,N_14963);
nand U18455 (N_18455,N_14953,N_11716);
and U18456 (N_18456,N_14497,N_14196);
or U18457 (N_18457,N_13849,N_10226);
nand U18458 (N_18458,N_11728,N_10867);
or U18459 (N_18459,N_14814,N_13283);
nor U18460 (N_18460,N_11295,N_10118);
xnor U18461 (N_18461,N_10279,N_13066);
xnor U18462 (N_18462,N_10604,N_10828);
and U18463 (N_18463,N_11836,N_10528);
and U18464 (N_18464,N_13542,N_14854);
nor U18465 (N_18465,N_13606,N_11484);
nor U18466 (N_18466,N_12844,N_10685);
or U18467 (N_18467,N_14141,N_12477);
and U18468 (N_18468,N_14386,N_13841);
nand U18469 (N_18469,N_14945,N_10614);
xor U18470 (N_18470,N_12050,N_13678);
xor U18471 (N_18471,N_11060,N_11436);
and U18472 (N_18472,N_14842,N_14380);
xor U18473 (N_18473,N_13804,N_14689);
nand U18474 (N_18474,N_11965,N_13145);
and U18475 (N_18475,N_11035,N_10991);
nand U18476 (N_18476,N_12158,N_12794);
nor U18477 (N_18477,N_12801,N_10522);
nand U18478 (N_18478,N_12352,N_13773);
and U18479 (N_18479,N_11149,N_14771);
and U18480 (N_18480,N_10960,N_10894);
xnor U18481 (N_18481,N_12166,N_11323);
or U18482 (N_18482,N_14061,N_12429);
nor U18483 (N_18483,N_14797,N_11192);
nor U18484 (N_18484,N_14225,N_14760);
or U18485 (N_18485,N_10450,N_11166);
nand U18486 (N_18486,N_13044,N_11649);
and U18487 (N_18487,N_14832,N_14105);
nor U18488 (N_18488,N_12697,N_12382);
nor U18489 (N_18489,N_14300,N_12314);
xor U18490 (N_18490,N_13185,N_14997);
or U18491 (N_18491,N_11311,N_12593);
nand U18492 (N_18492,N_11329,N_10059);
nor U18493 (N_18493,N_10870,N_14495);
and U18494 (N_18494,N_14896,N_13380);
and U18495 (N_18495,N_10708,N_11691);
or U18496 (N_18496,N_14551,N_13479);
or U18497 (N_18497,N_12873,N_13653);
xor U18498 (N_18498,N_12495,N_11905);
or U18499 (N_18499,N_12878,N_12598);
and U18500 (N_18500,N_14888,N_14111);
and U18501 (N_18501,N_13130,N_11723);
and U18502 (N_18502,N_10076,N_12675);
nand U18503 (N_18503,N_11771,N_11264);
nor U18504 (N_18504,N_11022,N_11658);
and U18505 (N_18505,N_12998,N_11025);
xor U18506 (N_18506,N_10114,N_13123);
xor U18507 (N_18507,N_14823,N_13547);
xnor U18508 (N_18508,N_12329,N_13042);
or U18509 (N_18509,N_10794,N_10107);
and U18510 (N_18510,N_13405,N_14940);
and U18511 (N_18511,N_11246,N_12381);
nor U18512 (N_18512,N_14748,N_14761);
nand U18513 (N_18513,N_13763,N_13391);
nor U18514 (N_18514,N_13802,N_14770);
xor U18515 (N_18515,N_13474,N_12572);
nand U18516 (N_18516,N_12447,N_12341);
xnor U18517 (N_18517,N_10528,N_14124);
xor U18518 (N_18518,N_13585,N_12407);
nand U18519 (N_18519,N_14037,N_11546);
and U18520 (N_18520,N_12104,N_11072);
xor U18521 (N_18521,N_12701,N_10311);
xor U18522 (N_18522,N_13206,N_10650);
xnor U18523 (N_18523,N_10467,N_12060);
nand U18524 (N_18524,N_13757,N_11041);
nand U18525 (N_18525,N_12790,N_13269);
nand U18526 (N_18526,N_13168,N_11237);
nand U18527 (N_18527,N_14719,N_12539);
nor U18528 (N_18528,N_10145,N_10323);
or U18529 (N_18529,N_14517,N_12146);
nor U18530 (N_18530,N_10962,N_11549);
and U18531 (N_18531,N_10148,N_13391);
and U18532 (N_18532,N_10395,N_11818);
and U18533 (N_18533,N_12537,N_10013);
or U18534 (N_18534,N_12301,N_11451);
nor U18535 (N_18535,N_10293,N_11983);
nand U18536 (N_18536,N_12541,N_14052);
or U18537 (N_18537,N_12424,N_14446);
and U18538 (N_18538,N_10547,N_13998);
xor U18539 (N_18539,N_10267,N_14321);
and U18540 (N_18540,N_10425,N_12092);
nor U18541 (N_18541,N_12437,N_13053);
xnor U18542 (N_18542,N_14199,N_13467);
nor U18543 (N_18543,N_14840,N_10482);
and U18544 (N_18544,N_10714,N_13172);
xnor U18545 (N_18545,N_13518,N_12915);
nor U18546 (N_18546,N_12622,N_12042);
and U18547 (N_18547,N_13209,N_10133);
or U18548 (N_18548,N_13843,N_13899);
or U18549 (N_18549,N_14604,N_12434);
or U18550 (N_18550,N_10421,N_11102);
nor U18551 (N_18551,N_11034,N_10125);
or U18552 (N_18552,N_11428,N_10612);
and U18553 (N_18553,N_10253,N_11219);
xnor U18554 (N_18554,N_13751,N_14526);
nor U18555 (N_18555,N_13610,N_12729);
or U18556 (N_18556,N_12902,N_12455);
nand U18557 (N_18557,N_13481,N_14988);
xor U18558 (N_18558,N_14599,N_10105);
or U18559 (N_18559,N_10988,N_14637);
or U18560 (N_18560,N_13471,N_10103);
nor U18561 (N_18561,N_10738,N_12887);
xnor U18562 (N_18562,N_12370,N_12653);
xnor U18563 (N_18563,N_11373,N_12218);
or U18564 (N_18564,N_13453,N_14952);
or U18565 (N_18565,N_13998,N_10112);
and U18566 (N_18566,N_14677,N_14993);
nor U18567 (N_18567,N_11351,N_11649);
nor U18568 (N_18568,N_13502,N_13370);
xor U18569 (N_18569,N_10154,N_13982);
nor U18570 (N_18570,N_13137,N_12478);
nor U18571 (N_18571,N_12580,N_12603);
or U18572 (N_18572,N_13553,N_13599);
xor U18573 (N_18573,N_11753,N_10902);
xnor U18574 (N_18574,N_10827,N_10108);
and U18575 (N_18575,N_11560,N_14143);
nand U18576 (N_18576,N_10985,N_12058);
nor U18577 (N_18577,N_12357,N_12850);
and U18578 (N_18578,N_13289,N_13904);
and U18579 (N_18579,N_11926,N_10517);
xor U18580 (N_18580,N_10692,N_13967);
and U18581 (N_18581,N_10179,N_13945);
nand U18582 (N_18582,N_12439,N_13240);
xor U18583 (N_18583,N_13460,N_13504);
xnor U18584 (N_18584,N_10303,N_13833);
and U18585 (N_18585,N_14073,N_11023);
or U18586 (N_18586,N_13170,N_14155);
and U18587 (N_18587,N_14114,N_11709);
xor U18588 (N_18588,N_12389,N_11124);
xnor U18589 (N_18589,N_13087,N_11728);
nand U18590 (N_18590,N_13499,N_11657);
xor U18591 (N_18591,N_12383,N_12066);
nor U18592 (N_18592,N_14746,N_11497);
and U18593 (N_18593,N_14056,N_10310);
or U18594 (N_18594,N_13123,N_12737);
or U18595 (N_18595,N_13988,N_11782);
or U18596 (N_18596,N_12621,N_10904);
and U18597 (N_18597,N_13807,N_13261);
nand U18598 (N_18598,N_11293,N_13373);
xnor U18599 (N_18599,N_14727,N_11326);
nand U18600 (N_18600,N_14896,N_10319);
nor U18601 (N_18601,N_10253,N_14858);
nand U18602 (N_18602,N_11031,N_13933);
or U18603 (N_18603,N_13340,N_10437);
and U18604 (N_18604,N_13360,N_12162);
or U18605 (N_18605,N_14039,N_12800);
and U18606 (N_18606,N_13298,N_10984);
or U18607 (N_18607,N_11094,N_11762);
nor U18608 (N_18608,N_10805,N_10656);
and U18609 (N_18609,N_12184,N_13746);
nand U18610 (N_18610,N_13568,N_11849);
and U18611 (N_18611,N_11489,N_11719);
and U18612 (N_18612,N_10922,N_12194);
and U18613 (N_18613,N_14221,N_12435);
or U18614 (N_18614,N_12376,N_12040);
xor U18615 (N_18615,N_10987,N_10537);
nand U18616 (N_18616,N_13920,N_11872);
or U18617 (N_18617,N_13894,N_14350);
xnor U18618 (N_18618,N_10596,N_13389);
nor U18619 (N_18619,N_11796,N_11953);
xnor U18620 (N_18620,N_14359,N_14747);
nand U18621 (N_18621,N_10528,N_12296);
xnor U18622 (N_18622,N_11830,N_10795);
xor U18623 (N_18623,N_12836,N_10444);
xnor U18624 (N_18624,N_11495,N_10752);
nor U18625 (N_18625,N_14676,N_13982);
and U18626 (N_18626,N_12532,N_10308);
or U18627 (N_18627,N_11581,N_10841);
nor U18628 (N_18628,N_12245,N_12337);
nand U18629 (N_18629,N_12764,N_11980);
nand U18630 (N_18630,N_10904,N_10542);
and U18631 (N_18631,N_11177,N_10095);
or U18632 (N_18632,N_12945,N_14439);
and U18633 (N_18633,N_13044,N_10967);
nor U18634 (N_18634,N_10674,N_10751);
and U18635 (N_18635,N_14749,N_10566);
xnor U18636 (N_18636,N_10424,N_11098);
and U18637 (N_18637,N_13940,N_11341);
nand U18638 (N_18638,N_11497,N_10472);
nor U18639 (N_18639,N_10190,N_11163);
xnor U18640 (N_18640,N_12893,N_13469);
xnor U18641 (N_18641,N_14331,N_11135);
nor U18642 (N_18642,N_10722,N_14179);
xor U18643 (N_18643,N_11002,N_11948);
nor U18644 (N_18644,N_13554,N_11569);
xor U18645 (N_18645,N_11140,N_14383);
xor U18646 (N_18646,N_13132,N_10904);
xor U18647 (N_18647,N_11745,N_12367);
and U18648 (N_18648,N_13021,N_10964);
nand U18649 (N_18649,N_14079,N_13547);
nand U18650 (N_18650,N_13499,N_12475);
nand U18651 (N_18651,N_10413,N_11021);
nor U18652 (N_18652,N_11765,N_14589);
nor U18653 (N_18653,N_11928,N_13126);
and U18654 (N_18654,N_10409,N_11531);
nor U18655 (N_18655,N_10305,N_12085);
nand U18656 (N_18656,N_11070,N_12001);
or U18657 (N_18657,N_10235,N_12188);
and U18658 (N_18658,N_10049,N_10375);
xnor U18659 (N_18659,N_12599,N_13112);
nand U18660 (N_18660,N_12735,N_11627);
nor U18661 (N_18661,N_13213,N_12423);
nand U18662 (N_18662,N_12588,N_13784);
xnor U18663 (N_18663,N_12163,N_11117);
nand U18664 (N_18664,N_10457,N_12268);
nand U18665 (N_18665,N_13339,N_10756);
and U18666 (N_18666,N_14580,N_13494);
xnor U18667 (N_18667,N_13404,N_11966);
nand U18668 (N_18668,N_10354,N_12207);
or U18669 (N_18669,N_10761,N_12802);
or U18670 (N_18670,N_13783,N_13518);
xor U18671 (N_18671,N_11618,N_10091);
nand U18672 (N_18672,N_13010,N_12148);
nand U18673 (N_18673,N_13038,N_13384);
nor U18674 (N_18674,N_14427,N_10483);
nor U18675 (N_18675,N_14044,N_14768);
nand U18676 (N_18676,N_12866,N_12403);
xnor U18677 (N_18677,N_10079,N_10606);
or U18678 (N_18678,N_12330,N_10567);
and U18679 (N_18679,N_14424,N_11560);
and U18680 (N_18680,N_13084,N_10174);
nand U18681 (N_18681,N_10163,N_10843);
xor U18682 (N_18682,N_13090,N_11855);
nand U18683 (N_18683,N_13786,N_12460);
nor U18684 (N_18684,N_11285,N_12324);
nor U18685 (N_18685,N_13654,N_13896);
or U18686 (N_18686,N_13820,N_14697);
nor U18687 (N_18687,N_13689,N_13277);
and U18688 (N_18688,N_11911,N_14896);
nor U18689 (N_18689,N_11481,N_12572);
and U18690 (N_18690,N_14420,N_11469);
nor U18691 (N_18691,N_11660,N_10709);
or U18692 (N_18692,N_14719,N_11875);
nand U18693 (N_18693,N_12018,N_12510);
or U18694 (N_18694,N_11008,N_13134);
nor U18695 (N_18695,N_13022,N_12173);
xnor U18696 (N_18696,N_13057,N_11727);
nand U18697 (N_18697,N_12292,N_14873);
nand U18698 (N_18698,N_12880,N_11033);
or U18699 (N_18699,N_11295,N_10297);
and U18700 (N_18700,N_10762,N_13882);
nor U18701 (N_18701,N_11882,N_13559);
nor U18702 (N_18702,N_10767,N_14342);
nor U18703 (N_18703,N_14597,N_10064);
nor U18704 (N_18704,N_10785,N_12775);
and U18705 (N_18705,N_11218,N_12502);
xnor U18706 (N_18706,N_14283,N_11584);
xor U18707 (N_18707,N_14797,N_14309);
and U18708 (N_18708,N_14892,N_14532);
nor U18709 (N_18709,N_11449,N_12256);
xor U18710 (N_18710,N_12058,N_13272);
xor U18711 (N_18711,N_14144,N_10093);
or U18712 (N_18712,N_12603,N_11541);
xnor U18713 (N_18713,N_11230,N_14485);
or U18714 (N_18714,N_13008,N_10320);
and U18715 (N_18715,N_12686,N_10085);
and U18716 (N_18716,N_10078,N_12714);
nor U18717 (N_18717,N_14106,N_10531);
and U18718 (N_18718,N_13564,N_12185);
xnor U18719 (N_18719,N_14054,N_10728);
nand U18720 (N_18720,N_14742,N_14537);
nand U18721 (N_18721,N_14345,N_12544);
nor U18722 (N_18722,N_13969,N_13489);
or U18723 (N_18723,N_11336,N_12651);
and U18724 (N_18724,N_14983,N_11122);
xor U18725 (N_18725,N_13479,N_12114);
nand U18726 (N_18726,N_12206,N_10948);
or U18727 (N_18727,N_14327,N_11418);
and U18728 (N_18728,N_10607,N_10316);
and U18729 (N_18729,N_14125,N_11008);
nand U18730 (N_18730,N_11676,N_14273);
or U18731 (N_18731,N_13985,N_12696);
nor U18732 (N_18732,N_10857,N_12891);
xor U18733 (N_18733,N_13821,N_12540);
or U18734 (N_18734,N_13297,N_14411);
or U18735 (N_18735,N_12416,N_14294);
and U18736 (N_18736,N_14377,N_14549);
xor U18737 (N_18737,N_12264,N_12121);
nand U18738 (N_18738,N_11789,N_12119);
nand U18739 (N_18739,N_12522,N_11843);
xor U18740 (N_18740,N_10890,N_11661);
nand U18741 (N_18741,N_14517,N_12780);
or U18742 (N_18742,N_13937,N_11460);
xnor U18743 (N_18743,N_12850,N_13098);
or U18744 (N_18744,N_14226,N_13324);
nand U18745 (N_18745,N_10464,N_11232);
or U18746 (N_18746,N_12359,N_12157);
nor U18747 (N_18747,N_13223,N_10802);
nand U18748 (N_18748,N_14240,N_13566);
nor U18749 (N_18749,N_12798,N_14477);
or U18750 (N_18750,N_12469,N_11010);
nor U18751 (N_18751,N_14542,N_12208);
and U18752 (N_18752,N_14650,N_13474);
or U18753 (N_18753,N_12082,N_12893);
and U18754 (N_18754,N_11439,N_11729);
xnor U18755 (N_18755,N_13835,N_10332);
xor U18756 (N_18756,N_11799,N_10426);
nor U18757 (N_18757,N_10272,N_14248);
nor U18758 (N_18758,N_13384,N_11117);
nor U18759 (N_18759,N_13784,N_11335);
xnor U18760 (N_18760,N_12137,N_10135);
xnor U18761 (N_18761,N_10352,N_13365);
nand U18762 (N_18762,N_11568,N_14716);
and U18763 (N_18763,N_11921,N_14358);
nand U18764 (N_18764,N_12437,N_11335);
nor U18765 (N_18765,N_12837,N_13388);
nand U18766 (N_18766,N_12572,N_11272);
xnor U18767 (N_18767,N_10981,N_10548);
xor U18768 (N_18768,N_10031,N_12004);
and U18769 (N_18769,N_11046,N_10701);
or U18770 (N_18770,N_11279,N_14894);
xnor U18771 (N_18771,N_14346,N_10812);
nand U18772 (N_18772,N_10896,N_11269);
and U18773 (N_18773,N_14207,N_12608);
or U18774 (N_18774,N_13970,N_10858);
or U18775 (N_18775,N_14856,N_13921);
nand U18776 (N_18776,N_10844,N_10211);
xnor U18777 (N_18777,N_14078,N_13769);
nand U18778 (N_18778,N_13820,N_13470);
or U18779 (N_18779,N_14433,N_12406);
nor U18780 (N_18780,N_14916,N_12357);
or U18781 (N_18781,N_10420,N_13025);
xnor U18782 (N_18782,N_11679,N_12430);
xnor U18783 (N_18783,N_12635,N_12276);
and U18784 (N_18784,N_10365,N_12695);
nand U18785 (N_18785,N_11649,N_12222);
and U18786 (N_18786,N_10266,N_14350);
or U18787 (N_18787,N_11850,N_14546);
xor U18788 (N_18788,N_12480,N_11446);
xnor U18789 (N_18789,N_11513,N_12790);
nor U18790 (N_18790,N_10280,N_11455);
xor U18791 (N_18791,N_14974,N_12915);
nand U18792 (N_18792,N_12957,N_11760);
xor U18793 (N_18793,N_14899,N_14631);
nor U18794 (N_18794,N_13732,N_12224);
nand U18795 (N_18795,N_10767,N_13449);
or U18796 (N_18796,N_12713,N_10128);
nor U18797 (N_18797,N_12447,N_11513);
and U18798 (N_18798,N_11861,N_14314);
nor U18799 (N_18799,N_10729,N_12278);
nand U18800 (N_18800,N_12783,N_10331);
and U18801 (N_18801,N_13255,N_12704);
or U18802 (N_18802,N_13597,N_12893);
and U18803 (N_18803,N_10763,N_14987);
xnor U18804 (N_18804,N_12118,N_10186);
or U18805 (N_18805,N_11333,N_12011);
nand U18806 (N_18806,N_10489,N_12874);
and U18807 (N_18807,N_12763,N_10251);
nand U18808 (N_18808,N_12174,N_11788);
xnor U18809 (N_18809,N_13907,N_12554);
nor U18810 (N_18810,N_10052,N_10160);
and U18811 (N_18811,N_14212,N_14129);
xnor U18812 (N_18812,N_14062,N_12725);
nor U18813 (N_18813,N_11614,N_14446);
nand U18814 (N_18814,N_13968,N_13803);
and U18815 (N_18815,N_14271,N_14338);
nand U18816 (N_18816,N_10674,N_14484);
xor U18817 (N_18817,N_11976,N_10369);
and U18818 (N_18818,N_11902,N_12001);
xnor U18819 (N_18819,N_12205,N_10581);
or U18820 (N_18820,N_11106,N_11213);
xor U18821 (N_18821,N_11899,N_11897);
nor U18822 (N_18822,N_12863,N_10951);
nand U18823 (N_18823,N_10227,N_13167);
and U18824 (N_18824,N_10395,N_11755);
and U18825 (N_18825,N_14356,N_11650);
nand U18826 (N_18826,N_12462,N_11501);
nand U18827 (N_18827,N_12857,N_11080);
nand U18828 (N_18828,N_13536,N_13687);
and U18829 (N_18829,N_13004,N_11657);
nor U18830 (N_18830,N_13738,N_11114);
nor U18831 (N_18831,N_14715,N_13726);
nor U18832 (N_18832,N_11788,N_12050);
xor U18833 (N_18833,N_10579,N_12308);
and U18834 (N_18834,N_13489,N_13388);
nand U18835 (N_18835,N_11334,N_13463);
or U18836 (N_18836,N_11254,N_13142);
and U18837 (N_18837,N_14663,N_14180);
nand U18838 (N_18838,N_13047,N_10570);
or U18839 (N_18839,N_13227,N_14447);
or U18840 (N_18840,N_12427,N_10911);
xnor U18841 (N_18841,N_10718,N_13938);
nand U18842 (N_18842,N_11814,N_10168);
xor U18843 (N_18843,N_11824,N_13258);
xnor U18844 (N_18844,N_14883,N_10459);
nand U18845 (N_18845,N_13611,N_12797);
or U18846 (N_18846,N_12089,N_12835);
nor U18847 (N_18847,N_10167,N_11877);
xor U18848 (N_18848,N_11671,N_11318);
or U18849 (N_18849,N_11568,N_13174);
xor U18850 (N_18850,N_10168,N_10405);
and U18851 (N_18851,N_10841,N_13348);
or U18852 (N_18852,N_12587,N_10156);
and U18853 (N_18853,N_12742,N_14921);
nand U18854 (N_18854,N_13722,N_12981);
nand U18855 (N_18855,N_12311,N_14361);
xor U18856 (N_18856,N_11994,N_10685);
nor U18857 (N_18857,N_11099,N_13428);
or U18858 (N_18858,N_11398,N_11772);
nand U18859 (N_18859,N_13476,N_12248);
or U18860 (N_18860,N_14126,N_10874);
nand U18861 (N_18861,N_10298,N_11816);
xnor U18862 (N_18862,N_12796,N_14726);
and U18863 (N_18863,N_10065,N_14655);
xnor U18864 (N_18864,N_10593,N_13302);
and U18865 (N_18865,N_13602,N_12192);
nand U18866 (N_18866,N_10682,N_10971);
and U18867 (N_18867,N_13249,N_11084);
nor U18868 (N_18868,N_10492,N_13464);
and U18869 (N_18869,N_10799,N_12732);
and U18870 (N_18870,N_10037,N_10768);
or U18871 (N_18871,N_11234,N_14882);
nand U18872 (N_18872,N_10711,N_10091);
nand U18873 (N_18873,N_10683,N_10109);
nand U18874 (N_18874,N_10674,N_11896);
or U18875 (N_18875,N_11438,N_14142);
xnor U18876 (N_18876,N_10689,N_14718);
or U18877 (N_18877,N_11731,N_10736);
xnor U18878 (N_18878,N_11494,N_14424);
nand U18879 (N_18879,N_11943,N_13290);
and U18880 (N_18880,N_10358,N_11342);
or U18881 (N_18881,N_10632,N_14695);
or U18882 (N_18882,N_12098,N_14013);
or U18883 (N_18883,N_10802,N_13943);
nor U18884 (N_18884,N_12712,N_11712);
nor U18885 (N_18885,N_13128,N_10393);
and U18886 (N_18886,N_10355,N_11857);
nand U18887 (N_18887,N_12035,N_14257);
nand U18888 (N_18888,N_11148,N_14126);
nand U18889 (N_18889,N_12267,N_11538);
xnor U18890 (N_18890,N_10647,N_10670);
nor U18891 (N_18891,N_14269,N_11902);
nor U18892 (N_18892,N_12214,N_13427);
nor U18893 (N_18893,N_13305,N_11865);
and U18894 (N_18894,N_13416,N_10486);
or U18895 (N_18895,N_11779,N_13938);
xor U18896 (N_18896,N_11670,N_12476);
and U18897 (N_18897,N_10869,N_14803);
xnor U18898 (N_18898,N_11413,N_10965);
and U18899 (N_18899,N_12985,N_11158);
nand U18900 (N_18900,N_12495,N_13193);
nand U18901 (N_18901,N_13711,N_12145);
or U18902 (N_18902,N_13299,N_10623);
or U18903 (N_18903,N_13736,N_12696);
nor U18904 (N_18904,N_13167,N_13383);
xnor U18905 (N_18905,N_13441,N_11981);
nor U18906 (N_18906,N_14252,N_10563);
or U18907 (N_18907,N_11135,N_12707);
nor U18908 (N_18908,N_13086,N_10672);
or U18909 (N_18909,N_13377,N_14689);
or U18910 (N_18910,N_12694,N_12907);
and U18911 (N_18911,N_10146,N_11876);
or U18912 (N_18912,N_14823,N_10517);
and U18913 (N_18913,N_14708,N_14877);
and U18914 (N_18914,N_14718,N_11981);
xnor U18915 (N_18915,N_10764,N_12529);
xnor U18916 (N_18916,N_10339,N_12821);
nor U18917 (N_18917,N_12041,N_10629);
nor U18918 (N_18918,N_13760,N_10911);
or U18919 (N_18919,N_10283,N_14771);
nor U18920 (N_18920,N_13396,N_10646);
nand U18921 (N_18921,N_13799,N_12326);
or U18922 (N_18922,N_12154,N_12631);
xnor U18923 (N_18923,N_10263,N_14298);
xor U18924 (N_18924,N_13217,N_14990);
and U18925 (N_18925,N_14597,N_14750);
nor U18926 (N_18926,N_11049,N_14673);
nor U18927 (N_18927,N_11825,N_10934);
nor U18928 (N_18928,N_12145,N_11208);
xnor U18929 (N_18929,N_12995,N_13372);
and U18930 (N_18930,N_14559,N_13408);
nor U18931 (N_18931,N_11877,N_14803);
xor U18932 (N_18932,N_11264,N_10078);
nor U18933 (N_18933,N_13889,N_13888);
and U18934 (N_18934,N_12465,N_14414);
xor U18935 (N_18935,N_13702,N_10918);
xnor U18936 (N_18936,N_14105,N_12970);
xor U18937 (N_18937,N_11577,N_14060);
and U18938 (N_18938,N_14989,N_14499);
and U18939 (N_18939,N_11370,N_11518);
xnor U18940 (N_18940,N_10050,N_10317);
nor U18941 (N_18941,N_12868,N_12060);
xnor U18942 (N_18942,N_14498,N_14459);
nor U18943 (N_18943,N_12875,N_13076);
nor U18944 (N_18944,N_14373,N_10211);
or U18945 (N_18945,N_11941,N_14108);
xor U18946 (N_18946,N_14157,N_11029);
or U18947 (N_18947,N_10569,N_10612);
and U18948 (N_18948,N_11807,N_11451);
nor U18949 (N_18949,N_13613,N_13340);
or U18950 (N_18950,N_14736,N_12917);
xor U18951 (N_18951,N_12203,N_14728);
xnor U18952 (N_18952,N_14862,N_10215);
nor U18953 (N_18953,N_10617,N_11323);
nor U18954 (N_18954,N_12447,N_14699);
and U18955 (N_18955,N_11275,N_14709);
and U18956 (N_18956,N_12417,N_14886);
nor U18957 (N_18957,N_14596,N_11420);
and U18958 (N_18958,N_10670,N_10811);
nand U18959 (N_18959,N_13030,N_13375);
xnor U18960 (N_18960,N_10205,N_13863);
nor U18961 (N_18961,N_13898,N_13206);
nand U18962 (N_18962,N_13765,N_14344);
xnor U18963 (N_18963,N_11753,N_11451);
xnor U18964 (N_18964,N_10530,N_10323);
xnor U18965 (N_18965,N_10201,N_13251);
xor U18966 (N_18966,N_10227,N_12090);
and U18967 (N_18967,N_11886,N_13369);
nor U18968 (N_18968,N_12618,N_11722);
xor U18969 (N_18969,N_12518,N_14362);
nand U18970 (N_18970,N_12954,N_13043);
nor U18971 (N_18971,N_11406,N_14685);
or U18972 (N_18972,N_12883,N_11383);
nor U18973 (N_18973,N_13352,N_13390);
and U18974 (N_18974,N_10254,N_11274);
or U18975 (N_18975,N_12196,N_11783);
nand U18976 (N_18976,N_14865,N_14189);
or U18977 (N_18977,N_11507,N_13900);
nor U18978 (N_18978,N_12523,N_14654);
or U18979 (N_18979,N_11490,N_10513);
or U18980 (N_18980,N_11173,N_11748);
nor U18981 (N_18981,N_12639,N_10161);
nand U18982 (N_18982,N_14196,N_14758);
or U18983 (N_18983,N_12343,N_11509);
nor U18984 (N_18984,N_12682,N_12770);
and U18985 (N_18985,N_14641,N_14910);
and U18986 (N_18986,N_11031,N_14045);
and U18987 (N_18987,N_10822,N_10652);
nand U18988 (N_18988,N_14078,N_13136);
nand U18989 (N_18989,N_14069,N_10446);
nor U18990 (N_18990,N_11925,N_11115);
nand U18991 (N_18991,N_11595,N_11189);
xnor U18992 (N_18992,N_12197,N_14099);
nor U18993 (N_18993,N_14290,N_14774);
and U18994 (N_18994,N_11607,N_11140);
and U18995 (N_18995,N_10825,N_14780);
nand U18996 (N_18996,N_12639,N_12848);
xor U18997 (N_18997,N_14685,N_14939);
nor U18998 (N_18998,N_11124,N_11932);
nor U18999 (N_18999,N_11412,N_14015);
nand U19000 (N_19000,N_14158,N_10132);
or U19001 (N_19001,N_12433,N_12835);
xor U19002 (N_19002,N_12539,N_11644);
and U19003 (N_19003,N_13332,N_14576);
nor U19004 (N_19004,N_14464,N_13136);
nand U19005 (N_19005,N_12505,N_12594);
or U19006 (N_19006,N_13423,N_12603);
or U19007 (N_19007,N_11707,N_12151);
and U19008 (N_19008,N_13177,N_11920);
nor U19009 (N_19009,N_10497,N_10502);
nand U19010 (N_19010,N_14241,N_10176);
xor U19011 (N_19011,N_13907,N_14632);
nand U19012 (N_19012,N_11158,N_14905);
nand U19013 (N_19013,N_14699,N_12679);
nor U19014 (N_19014,N_14424,N_10192);
xnor U19015 (N_19015,N_13991,N_14925);
or U19016 (N_19016,N_14355,N_11010);
nand U19017 (N_19017,N_13284,N_11555);
and U19018 (N_19018,N_14054,N_12693);
and U19019 (N_19019,N_11469,N_11005);
nor U19020 (N_19020,N_12955,N_11390);
and U19021 (N_19021,N_12909,N_10447);
nor U19022 (N_19022,N_14267,N_14339);
and U19023 (N_19023,N_10286,N_11694);
and U19024 (N_19024,N_14528,N_11953);
and U19025 (N_19025,N_11874,N_12737);
nor U19026 (N_19026,N_10184,N_11728);
nand U19027 (N_19027,N_10117,N_10428);
and U19028 (N_19028,N_13568,N_12049);
or U19029 (N_19029,N_14593,N_12162);
nand U19030 (N_19030,N_12657,N_12531);
nand U19031 (N_19031,N_13028,N_14723);
xnor U19032 (N_19032,N_10434,N_14653);
nand U19033 (N_19033,N_11847,N_10389);
nand U19034 (N_19034,N_12310,N_11823);
nand U19035 (N_19035,N_12141,N_13018);
xnor U19036 (N_19036,N_11403,N_13571);
xnor U19037 (N_19037,N_14801,N_12554);
and U19038 (N_19038,N_13397,N_14934);
xnor U19039 (N_19039,N_14351,N_12210);
nor U19040 (N_19040,N_11177,N_11503);
or U19041 (N_19041,N_11543,N_12236);
or U19042 (N_19042,N_12961,N_11973);
and U19043 (N_19043,N_12787,N_10021);
and U19044 (N_19044,N_14106,N_13731);
nor U19045 (N_19045,N_12332,N_14039);
nor U19046 (N_19046,N_11943,N_10263);
nor U19047 (N_19047,N_13446,N_10854);
or U19048 (N_19048,N_12174,N_10280);
or U19049 (N_19049,N_13097,N_13342);
nor U19050 (N_19050,N_13010,N_12189);
nor U19051 (N_19051,N_12791,N_13260);
or U19052 (N_19052,N_13784,N_12353);
or U19053 (N_19053,N_10087,N_13952);
xnor U19054 (N_19054,N_13165,N_14895);
or U19055 (N_19055,N_14335,N_10069);
nand U19056 (N_19056,N_10736,N_10247);
or U19057 (N_19057,N_12753,N_10875);
xor U19058 (N_19058,N_11569,N_11760);
and U19059 (N_19059,N_12955,N_11101);
and U19060 (N_19060,N_13358,N_12719);
nor U19061 (N_19061,N_10155,N_14669);
or U19062 (N_19062,N_14992,N_11003);
or U19063 (N_19063,N_13915,N_11760);
nor U19064 (N_19064,N_10311,N_13223);
xor U19065 (N_19065,N_12131,N_14400);
xor U19066 (N_19066,N_11868,N_12064);
nand U19067 (N_19067,N_14502,N_11872);
nor U19068 (N_19068,N_14346,N_14768);
nand U19069 (N_19069,N_13116,N_10642);
nand U19070 (N_19070,N_14736,N_12811);
or U19071 (N_19071,N_14146,N_14627);
nor U19072 (N_19072,N_14804,N_14159);
or U19073 (N_19073,N_14341,N_10671);
nor U19074 (N_19074,N_12730,N_11483);
nand U19075 (N_19075,N_14407,N_14031);
xnor U19076 (N_19076,N_14569,N_13052);
xor U19077 (N_19077,N_11141,N_12535);
and U19078 (N_19078,N_12885,N_14505);
nand U19079 (N_19079,N_13743,N_14870);
nor U19080 (N_19080,N_12752,N_14985);
nor U19081 (N_19081,N_11446,N_12827);
and U19082 (N_19082,N_14938,N_13739);
nand U19083 (N_19083,N_13682,N_12864);
xnor U19084 (N_19084,N_10749,N_11661);
or U19085 (N_19085,N_13718,N_14074);
nor U19086 (N_19086,N_14894,N_11823);
nand U19087 (N_19087,N_12828,N_14385);
nor U19088 (N_19088,N_11314,N_10479);
xnor U19089 (N_19089,N_12556,N_14382);
or U19090 (N_19090,N_12788,N_12098);
or U19091 (N_19091,N_14021,N_14550);
nand U19092 (N_19092,N_12496,N_11378);
nand U19093 (N_19093,N_14103,N_11265);
xnor U19094 (N_19094,N_14709,N_12399);
or U19095 (N_19095,N_13978,N_13191);
and U19096 (N_19096,N_11128,N_11650);
xor U19097 (N_19097,N_13845,N_12746);
and U19098 (N_19098,N_12987,N_11145);
nand U19099 (N_19099,N_14892,N_13270);
xor U19100 (N_19100,N_14893,N_12480);
and U19101 (N_19101,N_11902,N_11885);
xnor U19102 (N_19102,N_14317,N_12312);
and U19103 (N_19103,N_13256,N_11935);
or U19104 (N_19104,N_10804,N_11766);
nor U19105 (N_19105,N_14540,N_14100);
nor U19106 (N_19106,N_11841,N_14345);
xor U19107 (N_19107,N_13654,N_13938);
or U19108 (N_19108,N_14712,N_13787);
nor U19109 (N_19109,N_12158,N_13371);
or U19110 (N_19110,N_12259,N_12738);
nor U19111 (N_19111,N_13072,N_10851);
nor U19112 (N_19112,N_11286,N_11101);
and U19113 (N_19113,N_10526,N_14850);
nand U19114 (N_19114,N_14877,N_13568);
nand U19115 (N_19115,N_12811,N_13783);
nand U19116 (N_19116,N_10933,N_10203);
or U19117 (N_19117,N_10505,N_14704);
nor U19118 (N_19118,N_10710,N_12748);
xnor U19119 (N_19119,N_10670,N_11956);
and U19120 (N_19120,N_11817,N_13543);
nand U19121 (N_19121,N_12645,N_13468);
and U19122 (N_19122,N_12114,N_13913);
xor U19123 (N_19123,N_10430,N_11988);
nor U19124 (N_19124,N_10646,N_11554);
and U19125 (N_19125,N_11996,N_11186);
or U19126 (N_19126,N_12095,N_11982);
nor U19127 (N_19127,N_11812,N_12059);
nand U19128 (N_19128,N_13940,N_10158);
or U19129 (N_19129,N_13200,N_13079);
or U19130 (N_19130,N_11442,N_14362);
xor U19131 (N_19131,N_10803,N_14093);
nor U19132 (N_19132,N_13737,N_12486);
nor U19133 (N_19133,N_14644,N_14929);
and U19134 (N_19134,N_12375,N_10726);
nor U19135 (N_19135,N_12092,N_13738);
and U19136 (N_19136,N_11588,N_14231);
nor U19137 (N_19137,N_12787,N_14556);
nor U19138 (N_19138,N_14347,N_11783);
or U19139 (N_19139,N_12057,N_11717);
and U19140 (N_19140,N_13607,N_13966);
and U19141 (N_19141,N_10316,N_12145);
nor U19142 (N_19142,N_13083,N_14239);
or U19143 (N_19143,N_11000,N_12697);
nor U19144 (N_19144,N_14407,N_13823);
or U19145 (N_19145,N_12569,N_12097);
or U19146 (N_19146,N_12669,N_12443);
nor U19147 (N_19147,N_12651,N_12221);
xnor U19148 (N_19148,N_14391,N_14825);
or U19149 (N_19149,N_11851,N_12020);
nand U19150 (N_19150,N_13396,N_14699);
or U19151 (N_19151,N_13409,N_11285);
xnor U19152 (N_19152,N_13004,N_11528);
nor U19153 (N_19153,N_13700,N_11056);
xnor U19154 (N_19154,N_10938,N_12340);
or U19155 (N_19155,N_13160,N_11514);
or U19156 (N_19156,N_11477,N_13743);
nand U19157 (N_19157,N_12843,N_11103);
or U19158 (N_19158,N_13313,N_14814);
and U19159 (N_19159,N_14943,N_11477);
and U19160 (N_19160,N_14883,N_11007);
nor U19161 (N_19161,N_13125,N_10735);
nand U19162 (N_19162,N_12346,N_13306);
or U19163 (N_19163,N_13101,N_10336);
or U19164 (N_19164,N_10637,N_13730);
nor U19165 (N_19165,N_13389,N_14599);
nor U19166 (N_19166,N_13850,N_14313);
nand U19167 (N_19167,N_14900,N_12779);
and U19168 (N_19168,N_14564,N_10054);
and U19169 (N_19169,N_11596,N_12338);
and U19170 (N_19170,N_14863,N_13576);
xor U19171 (N_19171,N_13620,N_11380);
or U19172 (N_19172,N_10605,N_10769);
and U19173 (N_19173,N_11837,N_12776);
or U19174 (N_19174,N_13153,N_12820);
xor U19175 (N_19175,N_12931,N_13261);
nand U19176 (N_19176,N_13962,N_11977);
nor U19177 (N_19177,N_12424,N_10749);
or U19178 (N_19178,N_10810,N_14327);
nor U19179 (N_19179,N_11468,N_13431);
xnor U19180 (N_19180,N_14326,N_14943);
xnor U19181 (N_19181,N_13994,N_11976);
xnor U19182 (N_19182,N_10121,N_12476);
nand U19183 (N_19183,N_10718,N_13621);
and U19184 (N_19184,N_11825,N_10142);
xnor U19185 (N_19185,N_10218,N_14021);
and U19186 (N_19186,N_11487,N_14377);
nor U19187 (N_19187,N_10041,N_11154);
or U19188 (N_19188,N_11081,N_14257);
nor U19189 (N_19189,N_13840,N_14883);
or U19190 (N_19190,N_13317,N_14379);
nor U19191 (N_19191,N_11582,N_14448);
and U19192 (N_19192,N_13434,N_11783);
nand U19193 (N_19193,N_10858,N_12981);
and U19194 (N_19194,N_14678,N_14926);
xnor U19195 (N_19195,N_14886,N_12401);
xor U19196 (N_19196,N_13002,N_12742);
or U19197 (N_19197,N_11216,N_14367);
xnor U19198 (N_19198,N_12476,N_14847);
nor U19199 (N_19199,N_10790,N_11608);
nand U19200 (N_19200,N_10912,N_10500);
and U19201 (N_19201,N_10452,N_14414);
or U19202 (N_19202,N_14316,N_13840);
xor U19203 (N_19203,N_14813,N_14538);
or U19204 (N_19204,N_12597,N_11472);
nor U19205 (N_19205,N_10793,N_14307);
and U19206 (N_19206,N_11006,N_10745);
and U19207 (N_19207,N_14959,N_13373);
or U19208 (N_19208,N_14113,N_11368);
or U19209 (N_19209,N_10514,N_11932);
and U19210 (N_19210,N_13142,N_11193);
xnor U19211 (N_19211,N_12598,N_10677);
xnor U19212 (N_19212,N_14528,N_14170);
or U19213 (N_19213,N_14354,N_14949);
xor U19214 (N_19214,N_14524,N_10388);
and U19215 (N_19215,N_13178,N_12251);
nor U19216 (N_19216,N_11277,N_13984);
or U19217 (N_19217,N_12738,N_12921);
and U19218 (N_19218,N_10491,N_14577);
nor U19219 (N_19219,N_14006,N_11093);
xor U19220 (N_19220,N_14454,N_10664);
xor U19221 (N_19221,N_11220,N_11075);
nor U19222 (N_19222,N_11501,N_14865);
or U19223 (N_19223,N_14313,N_12703);
and U19224 (N_19224,N_11797,N_10143);
nand U19225 (N_19225,N_13111,N_13502);
or U19226 (N_19226,N_11779,N_10836);
nand U19227 (N_19227,N_14637,N_11933);
nand U19228 (N_19228,N_10332,N_10615);
xor U19229 (N_19229,N_14565,N_14344);
xor U19230 (N_19230,N_13849,N_12984);
or U19231 (N_19231,N_13522,N_10631);
nand U19232 (N_19232,N_11172,N_14581);
and U19233 (N_19233,N_14579,N_12786);
and U19234 (N_19234,N_14946,N_10112);
nand U19235 (N_19235,N_14694,N_13871);
and U19236 (N_19236,N_12583,N_14947);
or U19237 (N_19237,N_14573,N_14288);
or U19238 (N_19238,N_10175,N_14151);
nand U19239 (N_19239,N_11784,N_11624);
or U19240 (N_19240,N_12334,N_12716);
or U19241 (N_19241,N_10420,N_13789);
and U19242 (N_19242,N_12090,N_11103);
or U19243 (N_19243,N_11805,N_14825);
nand U19244 (N_19244,N_14801,N_11906);
nor U19245 (N_19245,N_10311,N_14510);
nor U19246 (N_19246,N_13261,N_11095);
and U19247 (N_19247,N_10992,N_14590);
and U19248 (N_19248,N_10397,N_10223);
xor U19249 (N_19249,N_11289,N_10691);
or U19250 (N_19250,N_13753,N_11508);
nand U19251 (N_19251,N_11988,N_10578);
xnor U19252 (N_19252,N_10603,N_12471);
and U19253 (N_19253,N_14253,N_12240);
xnor U19254 (N_19254,N_11191,N_14794);
nand U19255 (N_19255,N_11019,N_13528);
nor U19256 (N_19256,N_13354,N_12770);
nor U19257 (N_19257,N_12250,N_13193);
nor U19258 (N_19258,N_14014,N_14310);
nand U19259 (N_19259,N_12411,N_14450);
or U19260 (N_19260,N_14602,N_10031);
xnor U19261 (N_19261,N_11222,N_14260);
nand U19262 (N_19262,N_13045,N_10225);
xnor U19263 (N_19263,N_10526,N_12604);
nand U19264 (N_19264,N_11566,N_12144);
or U19265 (N_19265,N_13280,N_10049);
nor U19266 (N_19266,N_10088,N_10731);
and U19267 (N_19267,N_14049,N_12811);
or U19268 (N_19268,N_12441,N_12026);
xnor U19269 (N_19269,N_12769,N_13145);
xor U19270 (N_19270,N_11014,N_14457);
xnor U19271 (N_19271,N_10509,N_13671);
nand U19272 (N_19272,N_14080,N_12449);
and U19273 (N_19273,N_12228,N_13572);
nand U19274 (N_19274,N_13472,N_14561);
nor U19275 (N_19275,N_12981,N_10092);
and U19276 (N_19276,N_10810,N_10327);
and U19277 (N_19277,N_13511,N_11744);
and U19278 (N_19278,N_11925,N_13882);
nand U19279 (N_19279,N_12305,N_13297);
or U19280 (N_19280,N_14736,N_10929);
and U19281 (N_19281,N_14008,N_14711);
or U19282 (N_19282,N_12092,N_11977);
or U19283 (N_19283,N_11063,N_14778);
xor U19284 (N_19284,N_11355,N_12487);
nand U19285 (N_19285,N_10043,N_10125);
nor U19286 (N_19286,N_14684,N_12946);
nor U19287 (N_19287,N_10963,N_10126);
nand U19288 (N_19288,N_11156,N_14747);
xor U19289 (N_19289,N_12797,N_13438);
nand U19290 (N_19290,N_11639,N_10447);
nand U19291 (N_19291,N_13085,N_11807);
nor U19292 (N_19292,N_13342,N_10029);
nand U19293 (N_19293,N_14916,N_13166);
nand U19294 (N_19294,N_10513,N_14232);
nor U19295 (N_19295,N_14501,N_10766);
nor U19296 (N_19296,N_11489,N_14428);
or U19297 (N_19297,N_10308,N_11423);
nor U19298 (N_19298,N_10062,N_12839);
nand U19299 (N_19299,N_14538,N_12612);
and U19300 (N_19300,N_13198,N_10922);
nand U19301 (N_19301,N_13165,N_10698);
nor U19302 (N_19302,N_12264,N_10918);
nor U19303 (N_19303,N_11881,N_13286);
nand U19304 (N_19304,N_10290,N_10570);
nand U19305 (N_19305,N_10080,N_14656);
xor U19306 (N_19306,N_11117,N_13874);
xnor U19307 (N_19307,N_12621,N_13933);
xnor U19308 (N_19308,N_10923,N_11713);
nor U19309 (N_19309,N_12284,N_12454);
and U19310 (N_19310,N_10853,N_13657);
or U19311 (N_19311,N_12898,N_13683);
nor U19312 (N_19312,N_14610,N_10080);
nand U19313 (N_19313,N_10840,N_12352);
or U19314 (N_19314,N_13182,N_14084);
nand U19315 (N_19315,N_13008,N_13498);
nor U19316 (N_19316,N_14465,N_14516);
xor U19317 (N_19317,N_14977,N_13063);
nand U19318 (N_19318,N_12903,N_11164);
xor U19319 (N_19319,N_11026,N_13843);
nor U19320 (N_19320,N_14940,N_14770);
nor U19321 (N_19321,N_11301,N_13786);
nor U19322 (N_19322,N_11767,N_12483);
nand U19323 (N_19323,N_13914,N_10145);
and U19324 (N_19324,N_10486,N_10212);
nor U19325 (N_19325,N_14311,N_13784);
xnor U19326 (N_19326,N_11375,N_12435);
and U19327 (N_19327,N_10843,N_14437);
xor U19328 (N_19328,N_11786,N_13066);
xnor U19329 (N_19329,N_12841,N_13950);
nand U19330 (N_19330,N_11866,N_11909);
nand U19331 (N_19331,N_13517,N_14641);
xor U19332 (N_19332,N_11214,N_13201);
xnor U19333 (N_19333,N_13005,N_11011);
and U19334 (N_19334,N_10084,N_13773);
and U19335 (N_19335,N_13375,N_13731);
nor U19336 (N_19336,N_13194,N_10289);
nand U19337 (N_19337,N_12211,N_10893);
xor U19338 (N_19338,N_13313,N_12062);
xor U19339 (N_19339,N_13954,N_13948);
nor U19340 (N_19340,N_13768,N_14083);
or U19341 (N_19341,N_11951,N_13288);
nor U19342 (N_19342,N_14237,N_11782);
and U19343 (N_19343,N_11937,N_10911);
nor U19344 (N_19344,N_12535,N_12084);
xor U19345 (N_19345,N_10525,N_13796);
or U19346 (N_19346,N_10026,N_12179);
nor U19347 (N_19347,N_12842,N_10998);
xor U19348 (N_19348,N_14022,N_10507);
nor U19349 (N_19349,N_11774,N_14067);
and U19350 (N_19350,N_10123,N_12187);
and U19351 (N_19351,N_14660,N_12942);
xnor U19352 (N_19352,N_10307,N_11249);
xnor U19353 (N_19353,N_13469,N_11057);
nor U19354 (N_19354,N_14555,N_14958);
or U19355 (N_19355,N_12283,N_14121);
nor U19356 (N_19356,N_14039,N_14772);
xnor U19357 (N_19357,N_12645,N_13059);
nor U19358 (N_19358,N_10245,N_10307);
nand U19359 (N_19359,N_10855,N_12935);
nand U19360 (N_19360,N_11947,N_11315);
and U19361 (N_19361,N_12510,N_12939);
nor U19362 (N_19362,N_11054,N_14320);
nor U19363 (N_19363,N_14166,N_13175);
and U19364 (N_19364,N_11452,N_13113);
xor U19365 (N_19365,N_13601,N_12722);
xor U19366 (N_19366,N_10186,N_14694);
and U19367 (N_19367,N_13620,N_12484);
nand U19368 (N_19368,N_13117,N_12232);
and U19369 (N_19369,N_10265,N_12411);
and U19370 (N_19370,N_11824,N_12277);
nand U19371 (N_19371,N_11357,N_13318);
nor U19372 (N_19372,N_13576,N_11483);
xnor U19373 (N_19373,N_14066,N_12761);
nor U19374 (N_19374,N_14579,N_13718);
and U19375 (N_19375,N_10198,N_13294);
or U19376 (N_19376,N_13396,N_10611);
nor U19377 (N_19377,N_14187,N_12227);
nor U19378 (N_19378,N_13500,N_13256);
nor U19379 (N_19379,N_13401,N_10890);
xnor U19380 (N_19380,N_14899,N_14866);
or U19381 (N_19381,N_12805,N_12161);
or U19382 (N_19382,N_10164,N_10333);
and U19383 (N_19383,N_10455,N_13357);
or U19384 (N_19384,N_10671,N_13625);
nor U19385 (N_19385,N_13457,N_13969);
or U19386 (N_19386,N_13684,N_14182);
xnor U19387 (N_19387,N_12038,N_14297);
nor U19388 (N_19388,N_12204,N_11627);
nand U19389 (N_19389,N_14318,N_10594);
nor U19390 (N_19390,N_12619,N_13944);
and U19391 (N_19391,N_10263,N_14280);
and U19392 (N_19392,N_14465,N_11541);
nor U19393 (N_19393,N_14611,N_13356);
or U19394 (N_19394,N_14889,N_14219);
nor U19395 (N_19395,N_10989,N_12375);
or U19396 (N_19396,N_14002,N_14790);
and U19397 (N_19397,N_11700,N_11423);
nor U19398 (N_19398,N_10624,N_11783);
nand U19399 (N_19399,N_13513,N_12185);
nor U19400 (N_19400,N_10637,N_10144);
and U19401 (N_19401,N_14697,N_11812);
or U19402 (N_19402,N_14095,N_10072);
nor U19403 (N_19403,N_14595,N_11315);
nor U19404 (N_19404,N_13474,N_11426);
nand U19405 (N_19405,N_11914,N_14683);
xnor U19406 (N_19406,N_10787,N_11940);
or U19407 (N_19407,N_11745,N_10866);
and U19408 (N_19408,N_13640,N_10415);
nor U19409 (N_19409,N_11722,N_10437);
or U19410 (N_19410,N_13894,N_14439);
nor U19411 (N_19411,N_12907,N_13777);
xnor U19412 (N_19412,N_14299,N_12034);
nor U19413 (N_19413,N_13197,N_12608);
nand U19414 (N_19414,N_13762,N_14244);
xnor U19415 (N_19415,N_13970,N_10646);
and U19416 (N_19416,N_13484,N_11455);
xnor U19417 (N_19417,N_13363,N_10335);
nor U19418 (N_19418,N_10530,N_14450);
or U19419 (N_19419,N_10920,N_13256);
xnor U19420 (N_19420,N_10697,N_14779);
nand U19421 (N_19421,N_11389,N_11007);
nor U19422 (N_19422,N_12232,N_13246);
xor U19423 (N_19423,N_13797,N_13263);
and U19424 (N_19424,N_13064,N_13291);
or U19425 (N_19425,N_13061,N_13586);
nor U19426 (N_19426,N_11163,N_13196);
nand U19427 (N_19427,N_14952,N_13899);
xnor U19428 (N_19428,N_13690,N_10272);
nand U19429 (N_19429,N_11008,N_12681);
nand U19430 (N_19430,N_13306,N_13336);
or U19431 (N_19431,N_13975,N_11991);
and U19432 (N_19432,N_11053,N_14052);
and U19433 (N_19433,N_10039,N_11851);
or U19434 (N_19434,N_14743,N_10070);
nand U19435 (N_19435,N_12622,N_10626);
or U19436 (N_19436,N_12281,N_14954);
xnor U19437 (N_19437,N_13555,N_13344);
nand U19438 (N_19438,N_11819,N_11384);
or U19439 (N_19439,N_11218,N_12866);
xnor U19440 (N_19440,N_14637,N_14038);
or U19441 (N_19441,N_11170,N_12468);
nand U19442 (N_19442,N_13597,N_11791);
nor U19443 (N_19443,N_10867,N_12889);
nor U19444 (N_19444,N_12851,N_14771);
xor U19445 (N_19445,N_10805,N_12149);
xnor U19446 (N_19446,N_10654,N_11370);
nor U19447 (N_19447,N_14775,N_14879);
xor U19448 (N_19448,N_12764,N_13553);
or U19449 (N_19449,N_14301,N_12096);
xnor U19450 (N_19450,N_13054,N_12405);
xnor U19451 (N_19451,N_12570,N_10195);
and U19452 (N_19452,N_14139,N_14981);
nor U19453 (N_19453,N_11320,N_10365);
nor U19454 (N_19454,N_11561,N_12047);
nand U19455 (N_19455,N_13659,N_14280);
and U19456 (N_19456,N_14296,N_10177);
or U19457 (N_19457,N_11216,N_14822);
nand U19458 (N_19458,N_12193,N_11041);
xor U19459 (N_19459,N_13788,N_12006);
and U19460 (N_19460,N_14383,N_11930);
xnor U19461 (N_19461,N_11857,N_11006);
or U19462 (N_19462,N_11306,N_14810);
and U19463 (N_19463,N_13110,N_12374);
and U19464 (N_19464,N_12134,N_13515);
xnor U19465 (N_19465,N_10435,N_12274);
and U19466 (N_19466,N_10009,N_12374);
and U19467 (N_19467,N_10612,N_14059);
or U19468 (N_19468,N_11642,N_13800);
nor U19469 (N_19469,N_10787,N_12098);
xnor U19470 (N_19470,N_14449,N_14759);
nor U19471 (N_19471,N_14054,N_11886);
and U19472 (N_19472,N_13043,N_11976);
nor U19473 (N_19473,N_12741,N_10566);
nand U19474 (N_19474,N_14237,N_12849);
and U19475 (N_19475,N_11685,N_13963);
and U19476 (N_19476,N_11320,N_14327);
xor U19477 (N_19477,N_14639,N_12772);
nor U19478 (N_19478,N_11815,N_11714);
and U19479 (N_19479,N_14175,N_13273);
nand U19480 (N_19480,N_13423,N_12855);
nand U19481 (N_19481,N_14969,N_14324);
nand U19482 (N_19482,N_14537,N_14079);
and U19483 (N_19483,N_10119,N_12044);
nor U19484 (N_19484,N_11972,N_13881);
and U19485 (N_19485,N_13067,N_12895);
or U19486 (N_19486,N_12040,N_11505);
nor U19487 (N_19487,N_10488,N_11434);
and U19488 (N_19488,N_13162,N_14514);
nand U19489 (N_19489,N_11554,N_13873);
xor U19490 (N_19490,N_12963,N_12894);
nor U19491 (N_19491,N_13152,N_13657);
nand U19492 (N_19492,N_12400,N_13449);
and U19493 (N_19493,N_10451,N_12213);
xnor U19494 (N_19494,N_11253,N_11964);
nor U19495 (N_19495,N_11521,N_14481);
and U19496 (N_19496,N_13236,N_10393);
nand U19497 (N_19497,N_14112,N_12286);
xnor U19498 (N_19498,N_14151,N_13450);
and U19499 (N_19499,N_11855,N_13355);
or U19500 (N_19500,N_12624,N_11298);
or U19501 (N_19501,N_11549,N_14239);
xnor U19502 (N_19502,N_12578,N_12076);
xnor U19503 (N_19503,N_10318,N_14571);
xor U19504 (N_19504,N_10761,N_13266);
and U19505 (N_19505,N_14504,N_12596);
and U19506 (N_19506,N_10710,N_10152);
nand U19507 (N_19507,N_13206,N_10975);
nand U19508 (N_19508,N_13102,N_10725);
nand U19509 (N_19509,N_10489,N_14612);
xor U19510 (N_19510,N_11130,N_12025);
xor U19511 (N_19511,N_12580,N_13324);
and U19512 (N_19512,N_13996,N_10398);
nor U19513 (N_19513,N_14210,N_10126);
and U19514 (N_19514,N_14796,N_10209);
and U19515 (N_19515,N_14806,N_13464);
xnor U19516 (N_19516,N_10112,N_13433);
or U19517 (N_19517,N_14282,N_14483);
xnor U19518 (N_19518,N_12639,N_10383);
xnor U19519 (N_19519,N_14482,N_10073);
xor U19520 (N_19520,N_11646,N_10407);
or U19521 (N_19521,N_12332,N_12981);
xnor U19522 (N_19522,N_10923,N_13740);
and U19523 (N_19523,N_12448,N_14261);
xnor U19524 (N_19524,N_13714,N_10184);
and U19525 (N_19525,N_12670,N_13733);
nor U19526 (N_19526,N_13639,N_10310);
or U19527 (N_19527,N_14507,N_13402);
and U19528 (N_19528,N_13826,N_11780);
nor U19529 (N_19529,N_11498,N_10206);
xnor U19530 (N_19530,N_14618,N_13115);
or U19531 (N_19531,N_11993,N_13239);
xor U19532 (N_19532,N_13415,N_12353);
nand U19533 (N_19533,N_10035,N_14595);
nand U19534 (N_19534,N_10771,N_14894);
or U19535 (N_19535,N_14140,N_10217);
nor U19536 (N_19536,N_11183,N_11875);
nor U19537 (N_19537,N_13890,N_13211);
nor U19538 (N_19538,N_11198,N_13329);
nand U19539 (N_19539,N_12086,N_14940);
nand U19540 (N_19540,N_11306,N_10027);
or U19541 (N_19541,N_11117,N_12814);
nor U19542 (N_19542,N_11522,N_10693);
xor U19543 (N_19543,N_13367,N_14606);
nor U19544 (N_19544,N_12549,N_10275);
and U19545 (N_19545,N_14600,N_10128);
or U19546 (N_19546,N_14318,N_12709);
nand U19547 (N_19547,N_10624,N_10819);
nor U19548 (N_19548,N_12506,N_14751);
nor U19549 (N_19549,N_12955,N_12462);
xor U19550 (N_19550,N_10329,N_11407);
xor U19551 (N_19551,N_10734,N_10084);
and U19552 (N_19552,N_13309,N_10460);
nand U19553 (N_19553,N_10140,N_12124);
nand U19554 (N_19554,N_14114,N_12910);
or U19555 (N_19555,N_11190,N_13159);
nand U19556 (N_19556,N_11511,N_13591);
nand U19557 (N_19557,N_14307,N_11438);
nand U19558 (N_19558,N_12646,N_12276);
xor U19559 (N_19559,N_11553,N_12332);
nor U19560 (N_19560,N_12296,N_13363);
xnor U19561 (N_19561,N_13267,N_14930);
and U19562 (N_19562,N_11800,N_12637);
nor U19563 (N_19563,N_14058,N_10995);
or U19564 (N_19564,N_11328,N_13496);
and U19565 (N_19565,N_13740,N_12542);
or U19566 (N_19566,N_10858,N_13117);
xor U19567 (N_19567,N_14467,N_11686);
xor U19568 (N_19568,N_14976,N_14291);
xnor U19569 (N_19569,N_13264,N_14760);
or U19570 (N_19570,N_14750,N_12394);
xor U19571 (N_19571,N_11985,N_14807);
xor U19572 (N_19572,N_13912,N_13313);
nand U19573 (N_19573,N_11563,N_13742);
or U19574 (N_19574,N_14997,N_12785);
nor U19575 (N_19575,N_14053,N_12174);
and U19576 (N_19576,N_14732,N_11933);
xor U19577 (N_19577,N_10336,N_14556);
nand U19578 (N_19578,N_11367,N_11447);
nand U19579 (N_19579,N_13408,N_12538);
nand U19580 (N_19580,N_11731,N_10415);
and U19581 (N_19581,N_14881,N_10336);
xor U19582 (N_19582,N_11644,N_12058);
or U19583 (N_19583,N_11680,N_11636);
or U19584 (N_19584,N_12987,N_10623);
nor U19585 (N_19585,N_14451,N_12872);
and U19586 (N_19586,N_11065,N_11244);
nand U19587 (N_19587,N_11342,N_14721);
or U19588 (N_19588,N_11309,N_11680);
or U19589 (N_19589,N_11574,N_12203);
xor U19590 (N_19590,N_10413,N_13545);
and U19591 (N_19591,N_12108,N_10782);
xor U19592 (N_19592,N_12607,N_13366);
nor U19593 (N_19593,N_11599,N_11902);
nor U19594 (N_19594,N_11338,N_11033);
and U19595 (N_19595,N_12385,N_14337);
and U19596 (N_19596,N_11688,N_11452);
and U19597 (N_19597,N_13351,N_14293);
xor U19598 (N_19598,N_10584,N_11129);
or U19599 (N_19599,N_14905,N_12595);
xnor U19600 (N_19600,N_13665,N_12514);
xor U19601 (N_19601,N_13041,N_12392);
xnor U19602 (N_19602,N_13024,N_14201);
xor U19603 (N_19603,N_12331,N_12221);
and U19604 (N_19604,N_13627,N_13307);
xnor U19605 (N_19605,N_10590,N_10718);
nand U19606 (N_19606,N_13841,N_13465);
or U19607 (N_19607,N_13344,N_11512);
or U19608 (N_19608,N_14757,N_14735);
nand U19609 (N_19609,N_10178,N_11107);
nand U19610 (N_19610,N_10812,N_11513);
nor U19611 (N_19611,N_10488,N_14965);
nand U19612 (N_19612,N_14410,N_12441);
nor U19613 (N_19613,N_10141,N_12147);
nand U19614 (N_19614,N_13035,N_11890);
and U19615 (N_19615,N_11387,N_12578);
nor U19616 (N_19616,N_12381,N_10903);
or U19617 (N_19617,N_10296,N_12511);
or U19618 (N_19618,N_14939,N_10379);
nand U19619 (N_19619,N_14345,N_12802);
nor U19620 (N_19620,N_13408,N_10055);
xor U19621 (N_19621,N_10609,N_11500);
nor U19622 (N_19622,N_14031,N_11335);
and U19623 (N_19623,N_12493,N_12589);
nor U19624 (N_19624,N_14789,N_14069);
nor U19625 (N_19625,N_13525,N_12061);
nand U19626 (N_19626,N_10753,N_10191);
or U19627 (N_19627,N_14959,N_14726);
nor U19628 (N_19628,N_12906,N_10870);
and U19629 (N_19629,N_11178,N_12524);
and U19630 (N_19630,N_11676,N_13561);
xor U19631 (N_19631,N_14819,N_12933);
and U19632 (N_19632,N_13592,N_11460);
xor U19633 (N_19633,N_10655,N_10152);
and U19634 (N_19634,N_12251,N_12878);
nor U19635 (N_19635,N_13607,N_10556);
nand U19636 (N_19636,N_14632,N_12249);
xor U19637 (N_19637,N_14949,N_12493);
nor U19638 (N_19638,N_10818,N_14148);
xnor U19639 (N_19639,N_12856,N_13753);
and U19640 (N_19640,N_11475,N_11820);
nor U19641 (N_19641,N_14680,N_13348);
nand U19642 (N_19642,N_12360,N_10174);
nor U19643 (N_19643,N_14811,N_12077);
and U19644 (N_19644,N_14073,N_10256);
nor U19645 (N_19645,N_10713,N_14631);
xor U19646 (N_19646,N_12142,N_14411);
and U19647 (N_19647,N_10114,N_12751);
and U19648 (N_19648,N_14639,N_12539);
xnor U19649 (N_19649,N_14179,N_10433);
or U19650 (N_19650,N_10369,N_10174);
nand U19651 (N_19651,N_14204,N_10064);
and U19652 (N_19652,N_11733,N_12037);
xnor U19653 (N_19653,N_10953,N_10474);
nand U19654 (N_19654,N_10927,N_13857);
xor U19655 (N_19655,N_12982,N_12652);
xnor U19656 (N_19656,N_10350,N_10490);
and U19657 (N_19657,N_10506,N_12835);
nand U19658 (N_19658,N_12255,N_11402);
xnor U19659 (N_19659,N_10680,N_12345);
nand U19660 (N_19660,N_14587,N_10163);
or U19661 (N_19661,N_14290,N_14593);
xor U19662 (N_19662,N_10531,N_11180);
or U19663 (N_19663,N_12748,N_11236);
or U19664 (N_19664,N_10347,N_10480);
xnor U19665 (N_19665,N_11685,N_13673);
nor U19666 (N_19666,N_11833,N_12667);
nand U19667 (N_19667,N_11616,N_12670);
xnor U19668 (N_19668,N_11534,N_10020);
xnor U19669 (N_19669,N_12521,N_14831);
and U19670 (N_19670,N_12812,N_13736);
or U19671 (N_19671,N_12998,N_11731);
nand U19672 (N_19672,N_13320,N_14349);
or U19673 (N_19673,N_14749,N_10244);
nand U19674 (N_19674,N_14181,N_12084);
nor U19675 (N_19675,N_13095,N_11929);
xnor U19676 (N_19676,N_10349,N_13663);
and U19677 (N_19677,N_14952,N_11451);
nand U19678 (N_19678,N_13249,N_10141);
nor U19679 (N_19679,N_14208,N_14954);
and U19680 (N_19680,N_10933,N_14155);
or U19681 (N_19681,N_12957,N_13660);
and U19682 (N_19682,N_10906,N_14422);
nor U19683 (N_19683,N_11996,N_12435);
xnor U19684 (N_19684,N_13874,N_11701);
and U19685 (N_19685,N_14833,N_13908);
or U19686 (N_19686,N_11052,N_14109);
and U19687 (N_19687,N_11577,N_12614);
nor U19688 (N_19688,N_14641,N_10633);
and U19689 (N_19689,N_11115,N_12710);
or U19690 (N_19690,N_12982,N_13678);
nor U19691 (N_19691,N_11178,N_14891);
and U19692 (N_19692,N_10950,N_12076);
xnor U19693 (N_19693,N_12129,N_13403);
xnor U19694 (N_19694,N_13570,N_12559);
and U19695 (N_19695,N_14344,N_11341);
nor U19696 (N_19696,N_11063,N_10715);
nor U19697 (N_19697,N_12354,N_12013);
nand U19698 (N_19698,N_14216,N_13510);
nand U19699 (N_19699,N_11784,N_12466);
nand U19700 (N_19700,N_14104,N_10180);
or U19701 (N_19701,N_14090,N_14384);
and U19702 (N_19702,N_10313,N_14817);
nand U19703 (N_19703,N_14876,N_13626);
nor U19704 (N_19704,N_12508,N_14324);
nand U19705 (N_19705,N_12914,N_12215);
and U19706 (N_19706,N_12455,N_13464);
and U19707 (N_19707,N_11848,N_11266);
xor U19708 (N_19708,N_12847,N_10435);
xnor U19709 (N_19709,N_13234,N_14824);
nor U19710 (N_19710,N_14020,N_11851);
nor U19711 (N_19711,N_14084,N_11218);
nand U19712 (N_19712,N_12197,N_11178);
xor U19713 (N_19713,N_11530,N_13601);
or U19714 (N_19714,N_14433,N_10461);
or U19715 (N_19715,N_14933,N_12340);
nor U19716 (N_19716,N_14835,N_10879);
and U19717 (N_19717,N_10358,N_14322);
nor U19718 (N_19718,N_11768,N_10203);
xnor U19719 (N_19719,N_13973,N_12668);
nor U19720 (N_19720,N_14958,N_14575);
and U19721 (N_19721,N_12534,N_12496);
nor U19722 (N_19722,N_14180,N_12336);
xnor U19723 (N_19723,N_11427,N_10812);
and U19724 (N_19724,N_11145,N_14005);
nor U19725 (N_19725,N_14132,N_12182);
xnor U19726 (N_19726,N_12579,N_10744);
or U19727 (N_19727,N_14687,N_12906);
nor U19728 (N_19728,N_11998,N_14055);
or U19729 (N_19729,N_14371,N_13731);
and U19730 (N_19730,N_11308,N_11399);
xor U19731 (N_19731,N_14977,N_14087);
nand U19732 (N_19732,N_11341,N_11470);
and U19733 (N_19733,N_10281,N_14643);
xnor U19734 (N_19734,N_13927,N_13292);
and U19735 (N_19735,N_11169,N_11096);
nand U19736 (N_19736,N_13895,N_11855);
or U19737 (N_19737,N_13392,N_12367);
or U19738 (N_19738,N_12315,N_14732);
nand U19739 (N_19739,N_12813,N_11691);
nor U19740 (N_19740,N_11478,N_12746);
nand U19741 (N_19741,N_12530,N_14213);
nor U19742 (N_19742,N_12482,N_11844);
or U19743 (N_19743,N_10692,N_13908);
and U19744 (N_19744,N_14505,N_11798);
xor U19745 (N_19745,N_10683,N_11819);
xor U19746 (N_19746,N_10608,N_12402);
nand U19747 (N_19747,N_10794,N_11143);
xnor U19748 (N_19748,N_12936,N_10403);
or U19749 (N_19749,N_14456,N_13736);
nand U19750 (N_19750,N_13749,N_11038);
nand U19751 (N_19751,N_13203,N_10509);
or U19752 (N_19752,N_11911,N_13422);
xor U19753 (N_19753,N_14430,N_11857);
nor U19754 (N_19754,N_11098,N_11412);
nand U19755 (N_19755,N_10360,N_10110);
and U19756 (N_19756,N_10981,N_14587);
xor U19757 (N_19757,N_10567,N_12818);
or U19758 (N_19758,N_14919,N_10610);
nor U19759 (N_19759,N_14271,N_14676);
and U19760 (N_19760,N_13527,N_14406);
or U19761 (N_19761,N_10419,N_11839);
xnor U19762 (N_19762,N_12904,N_11262);
nor U19763 (N_19763,N_14261,N_13457);
nor U19764 (N_19764,N_13199,N_13494);
or U19765 (N_19765,N_14811,N_11416);
and U19766 (N_19766,N_13091,N_11780);
nand U19767 (N_19767,N_12609,N_12887);
and U19768 (N_19768,N_14734,N_12657);
and U19769 (N_19769,N_14619,N_14416);
xor U19770 (N_19770,N_12773,N_12669);
nor U19771 (N_19771,N_12616,N_12627);
and U19772 (N_19772,N_14335,N_11893);
or U19773 (N_19773,N_14079,N_13070);
xnor U19774 (N_19774,N_11237,N_13837);
or U19775 (N_19775,N_11816,N_14869);
nor U19776 (N_19776,N_10431,N_11740);
and U19777 (N_19777,N_13367,N_12925);
nor U19778 (N_19778,N_12196,N_12581);
nand U19779 (N_19779,N_14035,N_11841);
nor U19780 (N_19780,N_14076,N_11977);
and U19781 (N_19781,N_12808,N_11959);
xnor U19782 (N_19782,N_14920,N_11337);
xnor U19783 (N_19783,N_13492,N_12741);
xor U19784 (N_19784,N_12783,N_12279);
xor U19785 (N_19785,N_14605,N_10630);
nand U19786 (N_19786,N_13595,N_11419);
nor U19787 (N_19787,N_14983,N_10576);
nand U19788 (N_19788,N_12770,N_14593);
nand U19789 (N_19789,N_13668,N_12421);
or U19790 (N_19790,N_12498,N_10620);
xnor U19791 (N_19791,N_12484,N_12652);
or U19792 (N_19792,N_11545,N_11514);
or U19793 (N_19793,N_13648,N_11032);
xnor U19794 (N_19794,N_14024,N_11015);
or U19795 (N_19795,N_14852,N_13176);
nand U19796 (N_19796,N_12384,N_11514);
or U19797 (N_19797,N_11831,N_13560);
or U19798 (N_19798,N_13665,N_11566);
nor U19799 (N_19799,N_11780,N_13338);
and U19800 (N_19800,N_13629,N_13314);
nor U19801 (N_19801,N_12221,N_10982);
xor U19802 (N_19802,N_10630,N_12025);
xor U19803 (N_19803,N_12782,N_12403);
xor U19804 (N_19804,N_12056,N_13056);
or U19805 (N_19805,N_12616,N_14965);
nand U19806 (N_19806,N_10732,N_10161);
nor U19807 (N_19807,N_14775,N_13995);
and U19808 (N_19808,N_14737,N_12389);
xnor U19809 (N_19809,N_14328,N_12282);
and U19810 (N_19810,N_11641,N_12133);
nand U19811 (N_19811,N_13959,N_12495);
or U19812 (N_19812,N_12659,N_12519);
xnor U19813 (N_19813,N_14697,N_11463);
or U19814 (N_19814,N_13450,N_14459);
nand U19815 (N_19815,N_12255,N_14019);
or U19816 (N_19816,N_10336,N_13876);
and U19817 (N_19817,N_10317,N_11922);
or U19818 (N_19818,N_11690,N_14230);
and U19819 (N_19819,N_14935,N_14141);
and U19820 (N_19820,N_13975,N_14527);
nand U19821 (N_19821,N_14340,N_12019);
or U19822 (N_19822,N_13810,N_12541);
or U19823 (N_19823,N_11515,N_10877);
or U19824 (N_19824,N_14095,N_10736);
nor U19825 (N_19825,N_14878,N_13010);
and U19826 (N_19826,N_13125,N_11482);
nor U19827 (N_19827,N_13591,N_10495);
or U19828 (N_19828,N_11593,N_14913);
nor U19829 (N_19829,N_12438,N_14661);
nor U19830 (N_19830,N_12390,N_13019);
nor U19831 (N_19831,N_11710,N_11966);
or U19832 (N_19832,N_14779,N_12144);
or U19833 (N_19833,N_11557,N_14413);
nand U19834 (N_19834,N_12296,N_12495);
and U19835 (N_19835,N_10283,N_11881);
nor U19836 (N_19836,N_13534,N_14175);
or U19837 (N_19837,N_11662,N_12035);
nor U19838 (N_19838,N_12035,N_11095);
nor U19839 (N_19839,N_12276,N_10663);
or U19840 (N_19840,N_13355,N_10671);
nor U19841 (N_19841,N_14138,N_11506);
or U19842 (N_19842,N_11258,N_12235);
or U19843 (N_19843,N_10922,N_12013);
nor U19844 (N_19844,N_10663,N_10728);
and U19845 (N_19845,N_10205,N_12417);
nor U19846 (N_19846,N_14082,N_10288);
nor U19847 (N_19847,N_12467,N_13037);
and U19848 (N_19848,N_12314,N_11637);
nor U19849 (N_19849,N_11725,N_10766);
nand U19850 (N_19850,N_11631,N_13928);
nor U19851 (N_19851,N_11049,N_12525);
nand U19852 (N_19852,N_10232,N_10466);
nand U19853 (N_19853,N_12617,N_10980);
and U19854 (N_19854,N_13850,N_10588);
or U19855 (N_19855,N_10194,N_14889);
and U19856 (N_19856,N_12448,N_10966);
nor U19857 (N_19857,N_13267,N_11162);
nand U19858 (N_19858,N_13828,N_10720);
nand U19859 (N_19859,N_11932,N_12298);
nand U19860 (N_19860,N_12414,N_12728);
or U19861 (N_19861,N_12492,N_13138);
nor U19862 (N_19862,N_14894,N_12883);
nor U19863 (N_19863,N_10714,N_11012);
xor U19864 (N_19864,N_10957,N_14522);
and U19865 (N_19865,N_10426,N_13405);
nor U19866 (N_19866,N_11410,N_14969);
nand U19867 (N_19867,N_12761,N_14163);
nor U19868 (N_19868,N_10491,N_12196);
or U19869 (N_19869,N_12586,N_12179);
xnor U19870 (N_19870,N_12666,N_10596);
or U19871 (N_19871,N_11262,N_14371);
nor U19872 (N_19872,N_13586,N_11753);
xor U19873 (N_19873,N_12570,N_14704);
nor U19874 (N_19874,N_13810,N_12986);
nand U19875 (N_19875,N_13277,N_10796);
xnor U19876 (N_19876,N_14466,N_14701);
nand U19877 (N_19877,N_13572,N_14819);
nand U19878 (N_19878,N_12157,N_13043);
and U19879 (N_19879,N_12447,N_12881);
and U19880 (N_19880,N_10668,N_13673);
nor U19881 (N_19881,N_10583,N_13326);
nand U19882 (N_19882,N_14638,N_11317);
or U19883 (N_19883,N_12403,N_10248);
xor U19884 (N_19884,N_14671,N_13903);
and U19885 (N_19885,N_13433,N_11979);
xnor U19886 (N_19886,N_11620,N_13873);
or U19887 (N_19887,N_10910,N_12125);
or U19888 (N_19888,N_14369,N_11760);
nor U19889 (N_19889,N_12098,N_12097);
xor U19890 (N_19890,N_11043,N_14197);
nor U19891 (N_19891,N_10103,N_12343);
nor U19892 (N_19892,N_11333,N_14247);
nor U19893 (N_19893,N_12492,N_13272);
and U19894 (N_19894,N_12118,N_11221);
nand U19895 (N_19895,N_11046,N_12580);
xor U19896 (N_19896,N_10481,N_10863);
xor U19897 (N_19897,N_12271,N_10334);
and U19898 (N_19898,N_11200,N_10850);
or U19899 (N_19899,N_12451,N_10136);
xnor U19900 (N_19900,N_14028,N_14515);
or U19901 (N_19901,N_10637,N_11060);
nand U19902 (N_19902,N_12556,N_10975);
nor U19903 (N_19903,N_14295,N_14193);
nor U19904 (N_19904,N_14503,N_11424);
or U19905 (N_19905,N_13692,N_12296);
xnor U19906 (N_19906,N_14585,N_12237);
xnor U19907 (N_19907,N_12172,N_12200);
or U19908 (N_19908,N_14202,N_12890);
nor U19909 (N_19909,N_13303,N_13429);
and U19910 (N_19910,N_10774,N_11384);
xnor U19911 (N_19911,N_13171,N_10787);
or U19912 (N_19912,N_12388,N_10002);
or U19913 (N_19913,N_10765,N_13473);
nand U19914 (N_19914,N_13079,N_11677);
or U19915 (N_19915,N_10024,N_10206);
nor U19916 (N_19916,N_14837,N_10706);
and U19917 (N_19917,N_11356,N_12835);
or U19918 (N_19918,N_13116,N_10268);
or U19919 (N_19919,N_13993,N_13259);
and U19920 (N_19920,N_12187,N_12169);
or U19921 (N_19921,N_11979,N_10869);
or U19922 (N_19922,N_12342,N_11717);
or U19923 (N_19923,N_10718,N_10191);
or U19924 (N_19924,N_12398,N_14569);
nor U19925 (N_19925,N_12755,N_10455);
nor U19926 (N_19926,N_12159,N_12391);
or U19927 (N_19927,N_14719,N_14806);
xor U19928 (N_19928,N_12937,N_14930);
and U19929 (N_19929,N_11113,N_11358);
or U19930 (N_19930,N_13042,N_14791);
nand U19931 (N_19931,N_11037,N_14216);
nor U19932 (N_19932,N_10013,N_10988);
and U19933 (N_19933,N_13774,N_13175);
xor U19934 (N_19934,N_14338,N_11760);
xnor U19935 (N_19935,N_11578,N_14649);
nand U19936 (N_19936,N_13033,N_11546);
xnor U19937 (N_19937,N_10653,N_11830);
and U19938 (N_19938,N_14553,N_13259);
xor U19939 (N_19939,N_13270,N_12137);
nand U19940 (N_19940,N_12747,N_12587);
nor U19941 (N_19941,N_10225,N_11892);
nor U19942 (N_19942,N_10426,N_14250);
and U19943 (N_19943,N_12744,N_14524);
xnor U19944 (N_19944,N_11847,N_12396);
xnor U19945 (N_19945,N_11101,N_14894);
nand U19946 (N_19946,N_14802,N_11661);
or U19947 (N_19947,N_11964,N_10703);
and U19948 (N_19948,N_12091,N_11097);
and U19949 (N_19949,N_12164,N_11067);
and U19950 (N_19950,N_11295,N_11431);
xor U19951 (N_19951,N_11091,N_10134);
nand U19952 (N_19952,N_12283,N_12153);
nor U19953 (N_19953,N_12229,N_10000);
xnor U19954 (N_19954,N_14667,N_13081);
nor U19955 (N_19955,N_12126,N_10272);
nand U19956 (N_19956,N_11804,N_11140);
nor U19957 (N_19957,N_10606,N_12730);
nor U19958 (N_19958,N_11581,N_10968);
and U19959 (N_19959,N_10567,N_10343);
nor U19960 (N_19960,N_12264,N_10432);
nor U19961 (N_19961,N_11560,N_10677);
nand U19962 (N_19962,N_10780,N_14519);
nand U19963 (N_19963,N_11444,N_12598);
nand U19964 (N_19964,N_10557,N_14126);
or U19965 (N_19965,N_12019,N_13830);
nand U19966 (N_19966,N_11074,N_11114);
nor U19967 (N_19967,N_13208,N_13114);
nor U19968 (N_19968,N_13973,N_14223);
nand U19969 (N_19969,N_10484,N_11066);
or U19970 (N_19970,N_11481,N_14572);
nand U19971 (N_19971,N_12832,N_12981);
xor U19972 (N_19972,N_13343,N_13722);
and U19973 (N_19973,N_12879,N_10674);
or U19974 (N_19974,N_13536,N_10216);
or U19975 (N_19975,N_10555,N_14803);
nor U19976 (N_19976,N_10658,N_13849);
nor U19977 (N_19977,N_10922,N_13996);
nand U19978 (N_19978,N_10332,N_13896);
or U19979 (N_19979,N_12852,N_14649);
or U19980 (N_19980,N_13998,N_13416);
nand U19981 (N_19981,N_13266,N_14140);
and U19982 (N_19982,N_11495,N_12084);
xor U19983 (N_19983,N_13502,N_11132);
nand U19984 (N_19984,N_14447,N_13773);
xor U19985 (N_19985,N_11759,N_13719);
xor U19986 (N_19986,N_14761,N_12068);
nor U19987 (N_19987,N_13462,N_10156);
nand U19988 (N_19988,N_14756,N_12511);
or U19989 (N_19989,N_13379,N_13964);
or U19990 (N_19990,N_13265,N_10177);
xnor U19991 (N_19991,N_10584,N_13905);
nor U19992 (N_19992,N_13085,N_12487);
nor U19993 (N_19993,N_11131,N_10317);
xnor U19994 (N_19994,N_12458,N_10773);
xor U19995 (N_19995,N_10371,N_11692);
xor U19996 (N_19996,N_12812,N_12521);
xor U19997 (N_19997,N_13840,N_12587);
xnor U19998 (N_19998,N_11979,N_13332);
and U19999 (N_19999,N_10935,N_13811);
nand UO_0 (O_0,N_16965,N_19073);
xnor UO_1 (O_1,N_17335,N_17755);
xor UO_2 (O_2,N_16209,N_16700);
xor UO_3 (O_3,N_16605,N_17164);
nand UO_4 (O_4,N_15535,N_19571);
and UO_5 (O_5,N_17757,N_17891);
and UO_6 (O_6,N_16816,N_15603);
nand UO_7 (O_7,N_19859,N_17798);
and UO_8 (O_8,N_18514,N_19965);
and UO_9 (O_9,N_19489,N_17660);
nand UO_10 (O_10,N_15375,N_17868);
and UO_11 (O_11,N_19088,N_16592);
nor UO_12 (O_12,N_17106,N_18490);
or UO_13 (O_13,N_17621,N_17321);
nor UO_14 (O_14,N_18629,N_16405);
nand UO_15 (O_15,N_18900,N_18021);
nand UO_16 (O_16,N_15287,N_15421);
and UO_17 (O_17,N_19492,N_17005);
and UO_18 (O_18,N_16773,N_16305);
nand UO_19 (O_19,N_16634,N_17664);
nor UO_20 (O_20,N_15538,N_19519);
xnor UO_21 (O_21,N_18234,N_15916);
nor UO_22 (O_22,N_19289,N_19649);
and UO_23 (O_23,N_18006,N_17021);
and UO_24 (O_24,N_16022,N_19243);
nor UO_25 (O_25,N_18979,N_16653);
xor UO_26 (O_26,N_17327,N_15076);
xor UO_27 (O_27,N_18618,N_17825);
or UO_28 (O_28,N_16990,N_17315);
nor UO_29 (O_29,N_17107,N_19895);
and UO_30 (O_30,N_18496,N_15181);
xnor UO_31 (O_31,N_18232,N_15308);
or UO_32 (O_32,N_17690,N_16230);
nor UO_33 (O_33,N_17665,N_18414);
xnor UO_34 (O_34,N_19525,N_15092);
nand UO_35 (O_35,N_16658,N_17003);
xnor UO_36 (O_36,N_19761,N_18740);
nand UO_37 (O_37,N_17175,N_19939);
and UO_38 (O_38,N_16543,N_19904);
or UO_39 (O_39,N_18755,N_19844);
nand UO_40 (O_40,N_17914,N_15631);
or UO_41 (O_41,N_18507,N_16900);
or UO_42 (O_42,N_19559,N_16250);
or UO_43 (O_43,N_18696,N_16876);
nand UO_44 (O_44,N_18619,N_15472);
nor UO_45 (O_45,N_15911,N_15992);
nor UO_46 (O_46,N_15401,N_18277);
or UO_47 (O_47,N_16312,N_16124);
nand UO_48 (O_48,N_19150,N_19179);
and UO_49 (O_49,N_16763,N_19295);
nor UO_50 (O_50,N_19343,N_15902);
or UO_51 (O_51,N_18446,N_19254);
and UO_52 (O_52,N_19326,N_17976);
and UO_53 (O_53,N_18298,N_19934);
or UO_54 (O_54,N_16884,N_17401);
or UO_55 (O_55,N_16721,N_15410);
nor UO_56 (O_56,N_15235,N_19167);
and UO_57 (O_57,N_15494,N_17795);
and UO_58 (O_58,N_18066,N_19183);
xnor UO_59 (O_59,N_19849,N_16636);
nand UO_60 (O_60,N_16943,N_18138);
nand UO_61 (O_61,N_19759,N_17622);
or UO_62 (O_62,N_19261,N_16954);
nand UO_63 (O_63,N_16602,N_17812);
xor UO_64 (O_64,N_15719,N_18864);
nand UO_65 (O_65,N_15079,N_18879);
and UO_66 (O_66,N_16383,N_17927);
and UO_67 (O_67,N_15377,N_19540);
or UO_68 (O_68,N_15748,N_15716);
nor UO_69 (O_69,N_18031,N_15269);
or UO_70 (O_70,N_16366,N_19958);
nand UO_71 (O_71,N_19432,N_15143);
xor UO_72 (O_72,N_19257,N_18665);
xnor UO_73 (O_73,N_19810,N_17864);
or UO_74 (O_74,N_15641,N_15470);
nand UO_75 (O_75,N_19842,N_19941);
nor UO_76 (O_76,N_19349,N_15214);
or UO_77 (O_77,N_19359,N_17410);
nand UO_78 (O_78,N_17793,N_19703);
xnor UO_79 (O_79,N_17531,N_15386);
xor UO_80 (O_80,N_16915,N_17648);
nor UO_81 (O_81,N_18017,N_15717);
or UO_82 (O_82,N_18447,N_18626);
nor UO_83 (O_83,N_17781,N_15735);
or UO_84 (O_84,N_17115,N_19505);
nand UO_85 (O_85,N_15511,N_17211);
and UO_86 (O_86,N_19338,N_15651);
or UO_87 (O_87,N_17370,N_16745);
or UO_88 (O_88,N_15014,N_16604);
and UO_89 (O_89,N_15579,N_19832);
and UO_90 (O_90,N_19056,N_16493);
or UO_91 (O_91,N_15407,N_16030);
xnor UO_92 (O_92,N_17871,N_16709);
and UO_93 (O_93,N_16938,N_15282);
xnor UO_94 (O_94,N_15489,N_17380);
xor UO_95 (O_95,N_16216,N_19841);
or UO_96 (O_96,N_19210,N_17212);
nor UO_97 (O_97,N_18393,N_19995);
xor UO_98 (O_98,N_15322,N_16425);
or UO_99 (O_99,N_16574,N_19371);
xor UO_100 (O_100,N_16142,N_19395);
nand UO_101 (O_101,N_16883,N_15905);
xor UO_102 (O_102,N_19990,N_18673);
nor UO_103 (O_103,N_19457,N_17904);
and UO_104 (O_104,N_16765,N_16572);
nor UO_105 (O_105,N_16245,N_17202);
nand UO_106 (O_106,N_18702,N_16200);
and UO_107 (O_107,N_19421,N_16109);
nand UO_108 (O_108,N_16754,N_19134);
and UO_109 (O_109,N_18759,N_16524);
nand UO_110 (O_110,N_19181,N_17899);
xor UO_111 (O_111,N_16307,N_18628);
nand UO_112 (O_112,N_17997,N_15926);
nor UO_113 (O_113,N_15586,N_17076);
xnor UO_114 (O_114,N_18047,N_19109);
and UO_115 (O_115,N_19807,N_17847);
and UO_116 (O_116,N_18376,N_16337);
nand UO_117 (O_117,N_19866,N_18027);
nor UO_118 (O_118,N_17672,N_18334);
or UO_119 (O_119,N_18279,N_18976);
or UO_120 (O_120,N_18373,N_18191);
and UO_121 (O_121,N_17097,N_16346);
nor UO_122 (O_122,N_19704,N_17708);
xnor UO_123 (O_123,N_18459,N_18061);
and UO_124 (O_124,N_15257,N_16238);
xor UO_125 (O_125,N_19597,N_18916);
xor UO_126 (O_126,N_16770,N_16823);
or UO_127 (O_127,N_15276,N_16614);
nor UO_128 (O_128,N_15029,N_16912);
nor UO_129 (O_129,N_17906,N_16006);
xor UO_130 (O_130,N_17921,N_15499);
nor UO_131 (O_131,N_19118,N_15175);
and UO_132 (O_132,N_18065,N_18125);
nand UO_133 (O_133,N_17023,N_17201);
or UO_134 (O_134,N_17736,N_16423);
nand UO_135 (O_135,N_18775,N_15464);
or UO_136 (O_136,N_19798,N_18337);
or UO_137 (O_137,N_15187,N_16304);
and UO_138 (O_138,N_15453,N_17247);
and UO_139 (O_139,N_19237,N_18478);
nand UO_140 (O_140,N_17326,N_17210);
xnor UO_141 (O_141,N_18560,N_19607);
and UO_142 (O_142,N_17192,N_19213);
nor UO_143 (O_143,N_19872,N_19443);
nand UO_144 (O_144,N_17070,N_18651);
xor UO_145 (O_145,N_17198,N_17287);
or UO_146 (O_146,N_17993,N_15388);
nor UO_147 (O_147,N_19923,N_19174);
and UO_148 (O_148,N_17886,N_17544);
xnor UO_149 (O_149,N_19960,N_16083);
or UO_150 (O_150,N_18904,N_18307);
xor UO_151 (O_151,N_16847,N_15712);
and UO_152 (O_152,N_17249,N_17581);
nor UO_153 (O_153,N_19630,N_18932);
and UO_154 (O_154,N_16065,N_17160);
or UO_155 (O_155,N_18647,N_16739);
or UO_156 (O_156,N_16373,N_17880);
or UO_157 (O_157,N_15742,N_17064);
or UO_158 (O_158,N_18533,N_17592);
xnor UO_159 (O_159,N_16828,N_19191);
nor UO_160 (O_160,N_18971,N_15506);
or UO_161 (O_161,N_16635,N_16835);
or UO_162 (O_162,N_18293,N_15786);
or UO_163 (O_163,N_18103,N_19802);
nand UO_164 (O_164,N_16212,N_15979);
nand UO_165 (O_165,N_17417,N_17985);
or UO_166 (O_166,N_16435,N_18348);
or UO_167 (O_167,N_18018,N_19555);
nand UO_168 (O_168,N_18427,N_19216);
xnor UO_169 (O_169,N_15823,N_19306);
nor UO_170 (O_170,N_15856,N_16067);
nor UO_171 (O_171,N_15596,N_16386);
or UO_172 (O_172,N_18720,N_18660);
xor UO_173 (O_173,N_15928,N_15057);
nor UO_174 (O_174,N_19907,N_15790);
nand UO_175 (O_175,N_15339,N_15554);
and UO_176 (O_176,N_17749,N_16338);
or UO_177 (O_177,N_15915,N_18952);
nand UO_178 (O_178,N_17088,N_19817);
xnor UO_179 (O_179,N_18413,N_16039);
nand UO_180 (O_180,N_19650,N_19901);
xnor UO_181 (O_181,N_18195,N_18513);
nor UO_182 (O_182,N_18625,N_19335);
nand UO_183 (O_183,N_19409,N_19446);
and UO_184 (O_184,N_19985,N_18617);
or UO_185 (O_185,N_15784,N_15879);
or UO_186 (O_186,N_16452,N_19594);
or UO_187 (O_187,N_16177,N_18402);
or UO_188 (O_188,N_17322,N_16603);
and UO_189 (O_189,N_17197,N_17360);
xnor UO_190 (O_190,N_18523,N_18784);
or UO_191 (O_191,N_19975,N_18477);
nor UO_192 (O_192,N_19885,N_18273);
nand UO_193 (O_193,N_18164,N_16045);
or UO_194 (O_194,N_18052,N_15259);
nor UO_195 (O_195,N_17228,N_19544);
and UO_196 (O_196,N_18147,N_19850);
nand UO_197 (O_197,N_19998,N_16797);
or UO_198 (O_198,N_16401,N_19935);
xnor UO_199 (O_199,N_15274,N_15542);
and UO_200 (O_200,N_16005,N_18936);
or UO_201 (O_201,N_16742,N_15700);
xor UO_202 (O_202,N_16479,N_17908);
and UO_203 (O_203,N_18291,N_15302);
and UO_204 (O_204,N_19081,N_17207);
xor UO_205 (O_205,N_16132,N_17451);
nor UO_206 (O_206,N_15771,N_19804);
nand UO_207 (O_207,N_19994,N_15679);
nand UO_208 (O_208,N_16474,N_18221);
xnor UO_209 (O_209,N_18358,N_19422);
nor UO_210 (O_210,N_15875,N_15424);
nand UO_211 (O_211,N_19404,N_17912);
nand UO_212 (O_212,N_16372,N_18753);
xor UO_213 (O_213,N_19330,N_17389);
or UO_214 (O_214,N_16936,N_15415);
xnor UO_215 (O_215,N_16907,N_18497);
and UO_216 (O_216,N_17834,N_16253);
nand UO_217 (O_217,N_19380,N_18611);
nor UO_218 (O_218,N_15537,N_17139);
or UO_219 (O_219,N_16855,N_16568);
nor UO_220 (O_220,N_15291,N_19442);
and UO_221 (O_221,N_19373,N_15625);
or UO_222 (O_222,N_16406,N_17391);
or UO_223 (O_223,N_18268,N_19689);
nand UO_224 (O_224,N_15277,N_19632);
and UO_225 (O_225,N_17116,N_17213);
and UO_226 (O_226,N_19893,N_17521);
nor UO_227 (O_227,N_16573,N_19546);
xor UO_228 (O_228,N_18118,N_18733);
and UO_229 (O_229,N_19613,N_17551);
nand UO_230 (O_230,N_17461,N_19493);
and UO_231 (O_231,N_19346,N_16813);
and UO_232 (O_232,N_17636,N_16606);
or UO_233 (O_233,N_16613,N_15253);
and UO_234 (O_234,N_15144,N_17136);
nand UO_235 (O_235,N_16066,N_15458);
or UO_236 (O_236,N_15686,N_16637);
or UO_237 (O_237,N_15907,N_16193);
or UO_238 (O_238,N_18394,N_17585);
and UO_239 (O_239,N_17733,N_17859);
nand UO_240 (O_240,N_16601,N_18008);
nand UO_241 (O_241,N_18874,N_18917);
xnor UO_242 (O_242,N_16159,N_19482);
xnor UO_243 (O_243,N_16453,N_16444);
and UO_244 (O_244,N_17361,N_19193);
or UO_245 (O_245,N_15056,N_17355);
xnor UO_246 (O_246,N_17274,N_18656);
nor UO_247 (O_247,N_17220,N_15395);
xnor UO_248 (O_248,N_19793,N_17447);
nor UO_249 (O_249,N_16928,N_16724);
and UO_250 (O_250,N_17369,N_18214);
and UO_251 (O_251,N_15229,N_18173);
nand UO_252 (O_252,N_15261,N_15313);
or UO_253 (O_253,N_19256,N_18303);
or UO_254 (O_254,N_17513,N_18860);
xor UO_255 (O_255,N_15370,N_16345);
or UO_256 (O_256,N_16623,N_17289);
xor UO_257 (O_257,N_17049,N_17727);
nor UO_258 (O_258,N_16420,N_19940);
and UO_259 (O_259,N_16344,N_18817);
xnor UO_260 (O_260,N_19105,N_19120);
and UO_261 (O_261,N_15987,N_16962);
or UO_262 (O_262,N_17712,N_17381);
and UO_263 (O_263,N_18395,N_15732);
or UO_264 (O_264,N_16911,N_15062);
or UO_265 (O_265,N_19561,N_18081);
or UO_266 (O_266,N_16695,N_19333);
xnor UO_267 (O_267,N_18687,N_17922);
xor UO_268 (O_268,N_15025,N_16903);
and UO_269 (O_269,N_15919,N_19470);
or UO_270 (O_270,N_17769,N_18750);
nor UO_271 (O_271,N_19287,N_18470);
nand UO_272 (O_272,N_19248,N_16061);
nand UO_273 (O_273,N_16378,N_18312);
and UO_274 (O_274,N_16660,N_18100);
nand UO_275 (O_275,N_16904,N_18010);
nand UO_276 (O_276,N_19004,N_15619);
nand UO_277 (O_277,N_18282,N_16424);
xnor UO_278 (O_278,N_17485,N_19751);
or UO_279 (O_279,N_17400,N_18857);
or UO_280 (O_280,N_17692,N_19671);
nand UO_281 (O_281,N_16485,N_15846);
and UO_282 (O_282,N_19430,N_19161);
or UO_283 (O_283,N_15240,N_15951);
nor UO_284 (O_284,N_19244,N_15148);
and UO_285 (O_285,N_18441,N_17445);
and UO_286 (O_286,N_19000,N_16003);
xor UO_287 (O_287,N_17264,N_16008);
nor UO_288 (O_288,N_16678,N_19483);
nand UO_289 (O_289,N_16272,N_15923);
nand UO_290 (O_290,N_16716,N_15460);
or UO_291 (O_291,N_17307,N_19427);
nor UO_292 (O_292,N_18505,N_15425);
or UO_293 (O_293,N_16978,N_18317);
and UO_294 (O_294,N_15435,N_15167);
and UO_295 (O_295,N_15706,N_19236);
nor UO_296 (O_296,N_19032,N_17570);
and UO_297 (O_297,N_17406,N_15011);
nor UO_298 (O_298,N_16254,N_18235);
and UO_299 (O_299,N_17556,N_19739);
nor UO_300 (O_300,N_18676,N_17158);
nand UO_301 (O_301,N_16897,N_18315);
xnor UO_302 (O_302,N_15135,N_15184);
nand UO_303 (O_303,N_19580,N_18175);
xnor UO_304 (O_304,N_17561,N_15970);
and UO_305 (O_305,N_19005,N_16382);
nand UO_306 (O_306,N_18335,N_16343);
nor UO_307 (O_307,N_15575,N_17881);
nor UO_308 (O_308,N_16171,N_15747);
nor UO_309 (O_309,N_19410,N_15985);
or UO_310 (O_310,N_18452,N_15637);
nor UO_311 (O_311,N_15505,N_16248);
nand UO_312 (O_312,N_15147,N_19063);
nor UO_313 (O_313,N_19777,N_18368);
nor UO_314 (O_314,N_16644,N_18422);
or UO_315 (O_315,N_18791,N_17087);
or UO_316 (O_316,N_15848,N_16808);
and UO_317 (O_317,N_15994,N_17935);
or UO_318 (O_318,N_15461,N_18415);
or UO_319 (O_319,N_19862,N_18893);
nor UO_320 (O_320,N_15945,N_16199);
nor UO_321 (O_321,N_17980,N_17071);
xor UO_322 (O_322,N_18126,N_16752);
xnor UO_323 (O_323,N_19121,N_15493);
xor UO_324 (O_324,N_15677,N_16916);
xor UO_325 (O_325,N_16888,N_16487);
nor UO_326 (O_326,N_18901,N_17500);
and UO_327 (O_327,N_15636,N_17366);
xor UO_328 (O_328,N_16454,N_18638);
xnor UO_329 (O_329,N_18834,N_15295);
or UO_330 (O_330,N_15614,N_18553);
xor UO_331 (O_331,N_19677,N_18922);
and UO_332 (O_332,N_16821,N_15367);
or UO_333 (O_333,N_16779,N_15394);
nor UO_334 (O_334,N_19401,N_18949);
nand UO_335 (O_335,N_17449,N_18658);
and UO_336 (O_336,N_19714,N_15806);
and UO_337 (O_337,N_16099,N_15122);
nand UO_338 (O_338,N_17078,N_18225);
and UO_339 (O_339,N_18377,N_18453);
and UO_340 (O_340,N_19917,N_19082);
nand UO_341 (O_341,N_15795,N_19246);
nor UO_342 (O_342,N_15446,N_15210);
nand UO_343 (O_343,N_16328,N_19783);
xor UO_344 (O_344,N_15929,N_17655);
and UO_345 (O_345,N_17635,N_17024);
nand UO_346 (O_346,N_18152,N_16351);
nand UO_347 (O_347,N_16924,N_15382);
and UO_348 (O_348,N_16131,N_16786);
and UO_349 (O_349,N_15528,N_17553);
and UO_350 (O_350,N_17583,N_17718);
nor UO_351 (O_351,N_16627,N_18948);
nor UO_352 (O_352,N_17863,N_18005);
and UO_353 (O_353,N_16078,N_16046);
xor UO_354 (O_354,N_16802,N_18501);
nand UO_355 (O_355,N_19983,N_16037);
nand UO_356 (O_356,N_17128,N_17044);
or UO_357 (O_357,N_18559,N_15720);
xnor UO_358 (O_358,N_19076,N_18633);
or UO_359 (O_359,N_19241,N_19723);
nand UO_360 (O_360,N_17893,N_19787);
nand UO_361 (O_361,N_16718,N_18862);
nand UO_362 (O_362,N_18104,N_18251);
nand UO_363 (O_363,N_16581,N_15899);
xnor UO_364 (O_364,N_18378,N_15616);
nor UO_365 (O_365,N_19265,N_16295);
nor UO_366 (O_366,N_16190,N_15449);
or UO_367 (O_367,N_15519,N_16398);
nor UO_368 (O_368,N_17497,N_17143);
xnor UO_369 (O_369,N_17227,N_18653);
or UO_370 (O_370,N_17262,N_16955);
and UO_371 (O_371,N_16858,N_17861);
nand UO_372 (O_372,N_16436,N_18153);
nand UO_373 (O_373,N_19881,N_17134);
xor UO_374 (O_374,N_19294,N_18991);
and UO_375 (O_375,N_18727,N_17481);
and UO_376 (O_376,N_19262,N_19222);
nand UO_377 (O_377,N_15590,N_18576);
nand UO_378 (O_378,N_18794,N_19423);
and UO_379 (O_379,N_16923,N_18231);
and UO_380 (O_380,N_18830,N_18326);
xnor UO_381 (O_381,N_16240,N_17177);
and UO_382 (O_382,N_15065,N_19038);
and UO_383 (O_383,N_18370,N_15389);
or UO_384 (O_384,N_19581,N_15558);
nand UO_385 (O_385,N_17495,N_16280);
nand UO_386 (O_386,N_19218,N_17946);
nand UO_387 (O_387,N_18230,N_19416);
or UO_388 (O_388,N_19406,N_16150);
nor UO_389 (O_389,N_17180,N_15185);
nand UO_390 (O_390,N_18072,N_19537);
nand UO_391 (O_391,N_15782,N_19054);
or UO_392 (O_392,N_18499,N_16587);
nand UO_393 (O_393,N_18581,N_16844);
nor UO_394 (O_394,N_18743,N_16442);
xnor UO_395 (O_395,N_19447,N_19745);
nand UO_396 (O_396,N_19285,N_18908);
nand UO_397 (O_397,N_18258,N_19033);
and UO_398 (O_398,N_17552,N_18709);
xor UO_399 (O_399,N_17316,N_16628);
xor UO_400 (O_400,N_16090,N_18799);
or UO_401 (O_401,N_16194,N_16784);
nand UO_402 (O_402,N_16300,N_19645);
and UO_403 (O_403,N_17932,N_19507);
nand UO_404 (O_404,N_19575,N_18518);
or UO_405 (O_405,N_17193,N_17883);
xor UO_406 (O_406,N_18200,N_16134);
xnor UO_407 (O_407,N_18101,N_15220);
or UO_408 (O_408,N_15871,N_15520);
nand UO_409 (O_409,N_17027,N_17028);
nand UO_410 (O_410,N_18713,N_16977);
or UO_411 (O_411,N_17701,N_16314);
nand UO_412 (O_412,N_15164,N_18295);
nand UO_413 (O_413,N_16749,N_17702);
nand UO_414 (O_414,N_15508,N_15171);
xnor UO_415 (O_415,N_17444,N_18624);
or UO_416 (O_416,N_18804,N_16685);
xor UO_417 (O_417,N_19838,N_19992);
xor UO_418 (O_418,N_15281,N_18412);
or UO_419 (O_419,N_18590,N_17966);
nand UO_420 (O_420,N_15172,N_15933);
xnor UO_421 (O_421,N_16275,N_16147);
or UO_422 (O_422,N_16694,N_16692);
nor UO_423 (O_423,N_17971,N_15134);
xnor UO_424 (O_424,N_19822,N_16859);
and UO_425 (O_425,N_16014,N_16617);
nor UO_426 (O_426,N_15352,N_19159);
nor UO_427 (O_427,N_19317,N_18838);
and UO_428 (O_428,N_16467,N_16713);
nand UO_429 (O_429,N_15202,N_19593);
or UO_430 (O_430,N_17297,N_19846);
xnor UO_431 (O_431,N_18340,N_17074);
xnor UO_432 (O_432,N_18328,N_18179);
or UO_433 (O_433,N_18265,N_15141);
and UO_434 (O_434,N_16680,N_19288);
nand UO_435 (O_435,N_16533,N_15102);
or UO_436 (O_436,N_16963,N_15208);
and UO_437 (O_437,N_18706,N_18439);
or UO_438 (O_438,N_18354,N_18958);
nor UO_439 (O_439,N_15480,N_18756);
and UO_440 (O_440,N_15814,N_19982);
or UO_441 (O_441,N_15682,N_15288);
nor UO_442 (O_442,N_16495,N_16416);
and UO_443 (O_443,N_17382,N_15789);
nand UO_444 (O_444,N_16669,N_17931);
nor UO_445 (O_445,N_16504,N_16176);
nand UO_446 (O_446,N_17813,N_15910);
or UO_447 (O_447,N_18278,N_19131);
or UO_448 (O_448,N_18375,N_17318);
nor UO_449 (O_449,N_19878,N_17545);
xor UO_450 (O_450,N_16670,N_16381);
nand UO_451 (O_451,N_16273,N_19439);
nor UO_452 (O_452,N_15294,N_15653);
xnor UO_453 (O_453,N_19557,N_16882);
or UO_454 (O_454,N_18451,N_17214);
or UO_455 (O_455,N_18181,N_17338);
and UO_456 (O_456,N_16320,N_19768);
nand UO_457 (O_457,N_18284,N_17826);
and UO_458 (O_458,N_15560,N_19280);
or UO_459 (O_459,N_18313,N_17794);
and UO_460 (O_460,N_15778,N_17385);
xnor UO_461 (O_461,N_18102,N_19496);
nand UO_462 (O_462,N_16158,N_16024);
xor UO_463 (O_463,N_17279,N_15661);
nor UO_464 (O_464,N_18531,N_18973);
xnor UO_465 (O_465,N_19153,N_17367);
or UO_466 (O_466,N_16326,N_18489);
nor UO_467 (O_467,N_15695,N_18053);
xor UO_468 (O_468,N_18690,N_16554);
and UO_469 (O_469,N_18261,N_17696);
nand UO_470 (O_470,N_19454,N_18616);
and UO_471 (O_471,N_16011,N_17694);
nand UO_472 (O_472,N_15454,N_17245);
nand UO_473 (O_473,N_16334,N_16917);
or UO_474 (O_474,N_17190,N_19903);
nand UO_475 (O_475,N_16015,N_17359);
xor UO_476 (O_476,N_16983,N_18526);
or UO_477 (O_477,N_19785,N_16531);
or UO_478 (O_478,N_15110,N_19047);
nor UO_479 (O_479,N_18024,N_16927);
or UO_480 (O_480,N_18736,N_15640);
xor UO_481 (O_481,N_19046,N_16322);
nand UO_482 (O_482,N_17740,N_15117);
and UO_483 (O_483,N_16033,N_17715);
nand UO_484 (O_484,N_15047,N_17129);
xnor UO_485 (O_485,N_16957,N_15342);
nor UO_486 (O_486,N_19364,N_18554);
or UO_487 (O_487,N_17066,N_16782);
nand UO_488 (O_488,N_19360,N_18982);
and UO_489 (O_489,N_15635,N_17114);
or UO_490 (O_490,N_15965,N_18620);
nor UO_491 (O_491,N_15290,N_18579);
nor UO_492 (O_492,N_17095,N_16086);
nor UO_493 (O_493,N_16129,N_16775);
and UO_494 (O_494,N_15063,N_15217);
nor UO_495 (O_495,N_15317,N_17007);
and UO_496 (O_496,N_17761,N_17343);
nor UO_497 (O_497,N_19176,N_15310);
and UO_498 (O_498,N_17748,N_18931);
or UO_499 (O_499,N_16117,N_17586);
or UO_500 (O_500,N_16010,N_16455);
nor UO_501 (O_501,N_18831,N_16926);
nand UO_502 (O_502,N_19465,N_15649);
xor UO_503 (O_503,N_18462,N_19201);
and UO_504 (O_504,N_19968,N_15545);
xor UO_505 (O_505,N_15468,N_16068);
nand UO_506 (O_506,N_18613,N_18567);
nor UO_507 (O_507,N_17598,N_19926);
xor UO_508 (O_508,N_18498,N_17772);
and UO_509 (O_509,N_15192,N_19532);
nand UO_510 (O_510,N_18994,N_17077);
and UO_511 (O_511,N_19303,N_19884);
or UO_512 (O_512,N_15158,N_19586);
nand UO_513 (O_513,N_15130,N_16542);
nand UO_514 (O_514,N_15084,N_16564);
nor UO_515 (O_515,N_17855,N_16885);
xor UO_516 (O_516,N_18212,N_16899);
and UO_517 (O_517,N_18873,N_17771);
nand UO_518 (O_518,N_15691,N_19328);
xnor UO_519 (O_519,N_18694,N_17758);
xnor UO_520 (O_520,N_19068,N_19057);
and UO_521 (O_521,N_18585,N_17093);
nor UO_522 (O_522,N_19808,N_16397);
and UO_523 (O_523,N_19882,N_19945);
nand UO_524 (O_524,N_15772,N_16428);
and UO_525 (O_525,N_16297,N_17530);
and UO_526 (O_526,N_15054,N_19378);
and UO_527 (O_527,N_19831,N_16691);
nor UO_528 (O_528,N_18172,N_15088);
and UO_529 (O_529,N_17800,N_19639);
xor UO_530 (O_530,N_19400,N_16615);
xnor UO_531 (O_531,N_18963,N_18409);
xnor UO_532 (O_532,N_17527,N_18782);
nand UO_533 (O_533,N_16266,N_17808);
nand UO_534 (O_534,N_16481,N_17423);
nand UO_535 (O_535,N_15569,N_15236);
nor UO_536 (O_536,N_17675,N_18699);
xnor UO_537 (O_537,N_18670,N_19315);
and UO_538 (O_538,N_16879,N_15566);
nand UO_539 (O_539,N_18964,N_19839);
xor UO_540 (O_540,N_18621,N_17843);
and UO_541 (O_541,N_19436,N_18168);
nand UO_542 (O_542,N_15002,N_15658);
xnor UO_543 (O_543,N_18255,N_19756);
xor UO_544 (O_544,N_17988,N_18711);
and UO_545 (O_545,N_19437,N_19170);
or UO_546 (O_546,N_18188,N_16550);
nand UO_547 (O_547,N_16832,N_17719);
and UO_548 (O_548,N_18674,N_19864);
and UO_549 (O_549,N_19906,N_15660);
nor UO_550 (O_550,N_17890,N_18851);
xor UO_551 (O_551,N_16873,N_18539);
xnor UO_552 (O_552,N_18210,N_17962);
xor UO_553 (O_553,N_19096,N_19976);
or UO_554 (O_554,N_15309,N_15019);
xnor UO_555 (O_555,N_15422,N_18990);
nor UO_556 (O_556,N_18848,N_16997);
or UO_557 (O_557,N_17091,N_15477);
and UO_558 (O_558,N_16089,N_15120);
nand UO_559 (O_559,N_16350,N_19471);
or UO_560 (O_560,N_17833,N_19075);
nand UO_561 (O_561,N_19717,N_19771);
nor UO_562 (O_562,N_17725,N_19002);
nand UO_563 (O_563,N_18920,N_17409);
nand UO_564 (O_564,N_19847,N_17742);
and UO_565 (O_565,N_18416,N_18096);
nor UO_566 (O_566,N_17995,N_17973);
or UO_567 (O_567,N_18826,N_17832);
nand UO_568 (O_568,N_16756,N_19684);
or UO_569 (O_569,N_15114,N_18944);
nand UO_570 (O_570,N_15633,N_15250);
nor UO_571 (O_571,N_18464,N_18071);
and UO_572 (O_572,N_15222,N_17186);
and UO_573 (O_573,N_18504,N_18520);
and UO_574 (O_574,N_15623,N_19009);
or UO_575 (O_575,N_17419,N_16120);
xnor UO_576 (O_576,N_15021,N_15251);
or UO_577 (O_577,N_16909,N_18663);
or UO_578 (O_578,N_19177,N_15896);
or UO_579 (O_579,N_17089,N_15195);
or UO_580 (O_580,N_15412,N_19616);
or UO_581 (O_581,N_17756,N_18816);
nand UO_582 (O_582,N_17432,N_17068);
and UO_583 (O_583,N_18300,N_17779);
or UO_584 (O_584,N_15152,N_16865);
nor UO_585 (O_585,N_15751,N_15306);
or UO_586 (O_586,N_18582,N_18306);
xor UO_587 (O_587,N_18798,N_15197);
or UO_588 (O_588,N_17339,N_15602);
xnor UO_589 (O_589,N_17103,N_18465);
xnor UO_590 (O_590,N_15589,N_16895);
nand UO_591 (O_591,N_17356,N_19172);
or UO_592 (O_592,N_15263,N_16994);
nand UO_593 (O_593,N_15906,N_16594);
and UO_594 (O_594,N_19577,N_18137);
and UO_595 (O_595,N_15364,N_19195);
nor UO_596 (O_596,N_15360,N_19931);
nand UO_597 (O_597,N_16421,N_17149);
nor UO_598 (O_598,N_19981,N_18591);
nor UO_599 (O_599,N_15805,N_16875);
nor UO_600 (O_600,N_17975,N_17244);
and UO_601 (O_601,N_18623,N_19387);
and UO_602 (O_602,N_17348,N_16591);
or UO_603 (O_603,N_17872,N_15901);
and UO_604 (O_604,N_15385,N_15865);
xnor UO_605 (O_605,N_15275,N_16210);
xnor UO_606 (O_606,N_19008,N_15909);
xnor UO_607 (O_607,N_18744,N_17809);
nor UO_608 (O_608,N_17480,N_15842);
or UO_609 (O_609,N_16755,N_16993);
xor UO_610 (O_610,N_18970,N_19463);
xnor UO_611 (O_611,N_19080,N_15857);
and UO_612 (O_612,N_17000,N_15647);
nor UO_613 (O_613,N_19135,N_19833);
nor UO_614 (O_614,N_16016,N_19059);
nand UO_615 (O_615,N_18686,N_15954);
and UO_616 (O_616,N_18583,N_18009);
xnor UO_617 (O_617,N_17413,N_19520);
nand UO_618 (O_618,N_16112,N_17025);
and UO_619 (O_619,N_16357,N_18111);
nor UO_620 (O_620,N_17970,N_17476);
xnor UO_621 (O_621,N_15803,N_17486);
and UO_622 (O_622,N_18601,N_17836);
or UO_623 (O_623,N_18903,N_17310);
nor UO_624 (O_624,N_16448,N_15634);
and UO_625 (O_625,N_16640,N_17818);
xor UO_626 (O_626,N_19765,N_19536);
nand UO_627 (O_627,N_18547,N_16837);
nand UO_628 (O_628,N_19018,N_15927);
nor UO_629 (O_629,N_15289,N_18309);
or UO_630 (O_630,N_17189,N_15196);
nor UO_631 (O_631,N_15340,N_16179);
or UO_632 (O_632,N_19823,N_17231);
nor UO_633 (O_633,N_17567,N_16968);
and UO_634 (O_634,N_19066,N_18492);
xnor UO_635 (O_635,N_19103,N_19706);
or UO_636 (O_636,N_15746,N_15479);
xnor UO_637 (O_637,N_17607,N_19466);
nor UO_638 (O_638,N_18032,N_18097);
nand UO_639 (O_639,N_15301,N_17487);
or UO_640 (O_640,N_18042,N_15498);
nor UO_641 (O_641,N_18158,N_16409);
xor UO_642 (O_642,N_15280,N_15834);
and UO_643 (O_643,N_18002,N_18192);
or UO_644 (O_644,N_19845,N_15138);
nor UO_645 (O_645,N_19012,N_19786);
nand UO_646 (O_646,N_19171,N_17127);
nand UO_647 (O_647,N_16135,N_16539);
or UO_648 (O_648,N_18603,N_18332);
xnor UO_649 (O_649,N_17435,N_19414);
nand UO_650 (O_650,N_18972,N_18712);
or UO_651 (O_651,N_16947,N_16433);
nor UO_652 (O_652,N_17119,N_16103);
or UO_653 (O_653,N_16647,N_18321);
nor UO_654 (O_654,N_16047,N_17765);
xor UO_655 (O_655,N_19726,N_18177);
nor UO_656 (O_656,N_18789,N_16681);
xnor UO_657 (O_657,N_16703,N_16469);
nor UO_658 (O_658,N_15572,N_15471);
nand UO_659 (O_659,N_15972,N_16494);
and UO_660 (O_660,N_15484,N_17875);
nor UO_661 (O_661,N_19665,N_18128);
and UO_662 (O_662,N_18742,N_15708);
nor UO_663 (O_663,N_19920,N_18406);
or UO_664 (O_664,N_16157,N_17388);
xnor UO_665 (O_665,N_15199,N_16940);
and UO_666 (O_666,N_18450,N_19342);
or UO_667 (O_667,N_16298,N_19168);
or UO_668 (O_668,N_16403,N_17543);
nand UO_669 (O_669,N_19925,N_16437);
xor UO_670 (O_670,N_17250,N_17033);
or UO_671 (O_671,N_18156,N_18909);
nor UO_672 (O_672,N_19155,N_16289);
or UO_673 (O_673,N_18614,N_19648);
nand UO_674 (O_674,N_17457,N_19498);
xor UO_675 (O_675,N_18218,N_15017);
or UO_676 (O_676,N_18530,N_19554);
xnor UO_677 (O_677,N_19776,N_19578);
or UO_678 (O_678,N_16466,N_15930);
xnor UO_679 (O_679,N_17365,N_18985);
or UO_680 (O_680,N_17503,N_19816);
nor UO_681 (O_681,N_16862,N_19238);
nand UO_682 (O_682,N_19944,N_18692);
xnor UO_683 (O_683,N_15701,N_16064);
nand UO_684 (O_684,N_19137,N_19770);
nor UO_685 (O_685,N_16804,N_19725);
nor UO_686 (O_686,N_18463,N_16417);
xor UO_687 (O_687,N_18992,N_15159);
and UO_688 (O_688,N_17564,N_18974);
and UO_689 (O_689,N_16522,N_18345);
nand UO_690 (O_690,N_19952,N_19962);
xnor UO_691 (O_691,N_15399,N_19874);
and UO_692 (O_692,N_15817,N_19426);
and UO_693 (O_693,N_19988,N_15737);
nand UO_694 (O_694,N_18580,N_18271);
and UO_695 (O_695,N_18850,N_16563);
and UO_696 (O_696,N_15252,N_16569);
and UO_697 (O_697,N_18068,N_17887);
xnor UO_698 (O_698,N_18171,N_18786);
nand UO_699 (O_699,N_18781,N_18678);
or UO_700 (O_700,N_17936,N_17810);
or UO_701 (O_701,N_16380,N_19865);
xor UO_702 (O_702,N_18436,N_19980);
nor UO_703 (O_703,N_16062,N_19245);
nor UO_704 (O_704,N_18304,N_15881);
nor UO_705 (O_705,N_15878,N_15839);
and UO_706 (O_706,N_19870,N_17153);
xnor UO_707 (O_707,N_19718,N_17443);
nand UO_708 (O_708,N_15146,N_17700);
nand UO_709 (O_709,N_19367,N_18962);
and UO_710 (O_710,N_17547,N_16013);
and UO_711 (O_711,N_17477,N_16683);
nand UO_712 (O_712,N_17048,N_17408);
xnor UO_713 (O_713,N_19044,N_17200);
nor UO_714 (O_714,N_16607,N_19381);
nand UO_715 (O_715,N_15201,N_15870);
nor UO_716 (O_716,N_18718,N_18995);
and UO_717 (O_717,N_19397,N_18146);
nand UO_718 (O_718,N_18534,N_18389);
nand UO_719 (O_719,N_16490,N_18013);
xor UO_720 (O_720,N_16002,N_15264);
xor UO_721 (O_721,N_15696,N_15440);
and UO_722 (O_722,N_17398,N_15361);
and UO_723 (O_723,N_15327,N_15664);
nand UO_724 (O_724,N_16044,N_15628);
nor UO_725 (O_725,N_19619,N_15721);
xor UO_726 (O_726,N_18937,N_15205);
and UO_727 (O_727,N_16622,N_18911);
and UO_728 (O_728,N_18596,N_19654);
or UO_729 (O_729,N_18881,N_15487);
or UO_730 (O_730,N_17479,N_15955);
nor UO_731 (O_731,N_15826,N_17098);
nand UO_732 (O_732,N_16556,N_19861);
nand UO_733 (O_733,N_19408,N_18193);
and UO_734 (O_734,N_15042,N_18359);
nor UO_735 (O_735,N_16166,N_17471);
and UO_736 (O_736,N_16975,N_16740);
xnor UO_737 (O_737,N_17296,N_17351);
xnor UO_738 (O_738,N_17332,N_16822);
xor UO_739 (O_739,N_16666,N_17014);
nor UO_740 (O_740,N_19921,N_19220);
xor UO_741 (O_741,N_15140,N_19247);
and UO_742 (O_742,N_15648,N_17004);
nand UO_743 (O_743,N_15934,N_17953);
nand UO_744 (O_744,N_19058,N_18430);
nor UO_745 (O_745,N_15966,N_19748);
and UO_746 (O_746,N_18959,N_18311);
nor UO_747 (O_747,N_19078,N_19743);
nor UO_748 (O_748,N_16359,N_19698);
nand UO_749 (O_749,N_18083,N_16352);
or UO_750 (O_750,N_17610,N_18067);
nor UO_751 (O_751,N_15568,N_16141);
and UO_752 (O_752,N_18122,N_15882);
nand UO_753 (O_753,N_18889,N_15587);
and UO_754 (O_754,N_18770,N_15093);
and UO_755 (O_755,N_19321,N_17155);
xor UO_756 (O_756,N_17142,N_17523);
or UO_757 (O_757,N_16404,N_17083);
nor UO_758 (O_758,N_17254,N_19633);
or UO_759 (O_759,N_15813,N_15536);
and UO_760 (O_760,N_16243,N_18793);
xnor UO_761 (O_761,N_18527,N_17942);
nor UO_762 (O_762,N_17301,N_18528);
or UO_763 (O_763,N_17763,N_16475);
nor UO_764 (O_764,N_15591,N_15445);
and UO_765 (O_765,N_15527,N_18790);
nand UO_766 (O_766,N_17240,N_15086);
nand UO_767 (O_767,N_15335,N_16562);
nor UO_768 (O_768,N_17357,N_16901);
nand UO_769 (O_769,N_17109,N_18350);
nand UO_770 (O_770,N_18110,N_17869);
xor UO_771 (O_771,N_19235,N_19252);
nor UO_772 (O_772,N_16654,N_17992);
or UO_773 (O_773,N_15761,N_18532);
xnor UO_774 (O_774,N_16799,N_17161);
and UO_775 (O_775,N_16445,N_16515);
nor UO_776 (O_776,N_17169,N_16723);
xor UO_777 (O_777,N_15133,N_16609);
xor UO_778 (O_778,N_17061,N_15015);
xor UO_779 (O_779,N_17731,N_18561);
xnor UO_780 (O_780,N_19311,N_16282);
or UO_781 (O_781,N_17528,N_19673);
nand UO_782 (O_782,N_17823,N_16087);
and UO_783 (O_783,N_15559,N_19548);
nand UO_784 (O_784,N_19614,N_17628);
nor UO_785 (O_785,N_18646,N_16471);
nand UO_786 (O_786,N_17498,N_16390);
nand UO_787 (O_787,N_19258,N_17344);
and UO_788 (O_788,N_18762,N_15510);
nor UO_789 (O_789,N_15791,N_16501);
nor UO_790 (O_790,N_16113,N_19271);
or UO_791 (O_791,N_15504,N_17276);
nand UO_792 (O_792,N_16559,N_19738);
or UO_793 (O_793,N_19890,N_19564);
nand UO_794 (O_794,N_19264,N_19455);
or UO_795 (O_795,N_17767,N_18408);
nand UO_796 (O_796,N_17502,N_15877);
nor UO_797 (O_797,N_19001,N_19209);
or UO_798 (O_798,N_19565,N_15315);
nor UO_799 (O_799,N_17358,N_15976);
xor UO_800 (O_800,N_18033,N_17637);
nand UO_801 (O_801,N_19450,N_15977);
xnor UO_802 (O_802,N_17156,N_19867);
and UO_803 (O_803,N_19425,N_16929);
and UO_804 (O_804,N_17804,N_19886);
xnor UO_805 (O_805,N_17587,N_15323);
and UO_806 (O_806,N_19977,N_18248);
nand UO_807 (O_807,N_18652,N_16139);
nor UO_808 (O_808,N_16729,N_17724);
and UO_809 (O_809,N_16427,N_19268);
nor UO_810 (O_810,N_16529,N_17840);
nand UO_811 (O_811,N_17407,N_15434);
and UO_812 (O_812,N_19101,N_19782);
nand UO_813 (O_813,N_17595,N_18640);
and UO_814 (O_814,N_18189,N_17792);
nand UO_815 (O_815,N_16831,N_18419);
or UO_816 (O_816,N_19693,N_17789);
nand UO_817 (O_817,N_17263,N_19194);
xnor UO_818 (O_818,N_18803,N_18812);
and UO_819 (O_819,N_16412,N_17303);
nand UO_820 (O_820,N_19871,N_17514);
nor UO_821 (O_821,N_15853,N_15420);
or UO_822 (O_822,N_19646,N_15441);
or UO_823 (O_823,N_15032,N_17372);
and UO_824 (O_824,N_17669,N_17069);
and UO_825 (O_825,N_17753,N_19668);
xnor UO_826 (O_826,N_18247,N_19514);
nand UO_827 (O_827,N_19927,N_17099);
or UO_828 (O_828,N_19755,N_18751);
and UO_829 (O_829,N_17349,N_15874);
xnor UO_830 (O_830,N_19628,N_18872);
and UO_831 (O_831,N_17375,N_16872);
nor UO_832 (O_832,N_17693,N_16095);
and UO_833 (O_833,N_17280,N_16668);
or UO_834 (O_834,N_15451,N_17805);
xor UO_835 (O_835,N_17363,N_18346);
xnor UO_836 (O_836,N_19284,N_16701);
and UO_837 (O_837,N_19211,N_17260);
and UO_838 (O_838,N_18259,N_17125);
xnor UO_839 (O_839,N_18723,N_15920);
xor UO_840 (O_840,N_18546,N_17283);
nand UO_841 (O_841,N_15863,N_15639);
and UO_842 (O_842,N_16889,N_18557);
nand UO_843 (O_843,N_16984,N_17463);
or UO_844 (O_844,N_19302,N_17600);
and UO_845 (O_845,N_17999,N_19909);
and UO_846 (O_846,N_18595,N_17052);
or UO_847 (O_847,N_18543,N_15962);
or UO_848 (O_848,N_19928,N_16023);
nor UO_849 (O_849,N_18767,N_15113);
and UO_850 (O_850,N_17824,N_16126);
xnor UO_851 (O_851,N_15003,N_15242);
nor UO_852 (O_852,N_15904,N_16905);
nand UO_853 (O_853,N_15749,N_16316);
xor UO_854 (O_854,N_16394,N_18469);
and UO_855 (O_855,N_16271,N_18134);
nand UO_856 (O_856,N_17802,N_17434);
nand UO_857 (O_857,N_17294,N_17852);
or UO_858 (O_858,N_18069,N_18832);
nand UO_859 (O_859,N_19835,N_19731);
nand UO_860 (O_860,N_19621,N_15239);
or UO_861 (O_861,N_18242,N_15858);
nor UO_862 (O_862,N_18584,N_19249);
nand UO_863 (O_863,N_16484,N_19757);
nand UO_864 (O_864,N_16093,N_15840);
nor UO_865 (O_865,N_17184,N_19605);
xor UO_866 (O_866,N_16235,N_17803);
nor UO_867 (O_867,N_16355,N_17785);
nor UO_868 (O_868,N_15330,N_15889);
nand UO_869 (O_869,N_18440,N_18837);
nand UO_870 (O_870,N_19686,N_15040);
or UO_871 (O_871,N_18203,N_16952);
or UO_872 (O_872,N_19352,N_16107);
nor UO_873 (O_873,N_18688,N_18897);
and UO_874 (O_874,N_17703,N_15338);
xor UO_875 (O_875,N_18105,N_19805);
and UO_876 (O_876,N_15298,N_18392);
xor UO_877 (O_877,N_16110,N_16265);
or UO_878 (O_878,N_15822,N_19722);
or UO_879 (O_879,N_15785,N_18682);
nor UO_880 (O_880,N_17229,N_17846);
xor UO_881 (O_881,N_19583,N_19966);
or UO_882 (O_882,N_16203,N_18763);
or UO_883 (O_883,N_19898,N_17989);
or UO_884 (O_884,N_19379,N_19438);
nand UO_885 (O_885,N_19658,N_16431);
xor UO_886 (O_886,N_18276,N_17392);
xor UO_887 (O_887,N_16215,N_19143);
nor UO_888 (O_888,N_15781,N_16525);
and UO_889 (O_889,N_15615,N_16146);
and UO_890 (O_890,N_18382,N_17347);
or UO_891 (O_891,N_16811,N_16375);
and UO_892 (O_892,N_18383,N_16100);
xor UO_893 (O_893,N_19970,N_16801);
nor UO_894 (O_894,N_18927,N_19711);
xnor UO_895 (O_895,N_19572,N_16017);
or UO_896 (O_896,N_16426,N_18724);
and UO_897 (O_897,N_15485,N_15750);
xnor UO_898 (O_898,N_16869,N_18266);
xor UO_899 (O_899,N_16287,N_15864);
xnor UO_900 (O_900,N_15442,N_16526);
nand UO_901 (O_901,N_19398,N_18019);
or UO_902 (O_902,N_18697,N_16812);
nand UO_903 (O_903,N_15474,N_18761);
nor UO_904 (O_904,N_15550,N_17266);
nor UO_905 (O_905,N_19741,N_16430);
nand UO_906 (O_906,N_19453,N_19314);
nor UO_907 (O_907,N_16656,N_16687);
or UO_908 (O_908,N_16679,N_17752);
nor UO_909 (O_909,N_19946,N_16296);
nand UO_910 (O_910,N_16202,N_18049);
nand UO_911 (O_911,N_18746,N_16119);
or UO_912 (O_912,N_19913,N_16846);
or UO_913 (O_913,N_15270,N_18672);
xnor UO_914 (O_914,N_15430,N_17159);
or UO_915 (O_915,N_15755,N_18915);
or UO_916 (O_916,N_17697,N_15983);
or UO_917 (O_917,N_18129,N_15157);
nor UO_918 (O_918,N_19896,N_16973);
xor UO_919 (O_919,N_19007,N_17402);
or UO_920 (O_920,N_15331,N_17617);
xor UO_921 (O_921,N_16422,N_19089);
or UO_922 (O_922,N_16162,N_16720);
and UO_923 (O_923,N_18854,N_15867);
nor UO_924 (O_924,N_19899,N_18121);
and UO_925 (O_925,N_17377,N_16118);
nand UO_926 (O_926,N_19813,N_16585);
nor UO_927 (O_927,N_16787,N_18715);
or UO_928 (O_928,N_19233,N_17569);
nand UO_929 (O_929,N_17286,N_18883);
xnor UO_930 (O_930,N_17633,N_17896);
and UO_931 (O_931,N_15312,N_16356);
nor UO_932 (O_932,N_17465,N_19523);
or UO_933 (O_933,N_17517,N_15812);
nor UO_934 (O_934,N_18327,N_19461);
xor UO_935 (O_935,N_16056,N_15265);
nand UO_936 (O_936,N_15443,N_19186);
and UO_937 (O_937,N_16339,N_16362);
xor UO_938 (O_938,N_15481,N_17707);
xor UO_939 (O_939,N_15160,N_15503);
nor UO_940 (O_940,N_17654,N_18131);
xor UO_941 (O_941,N_15573,N_15428);
nand UO_942 (O_942,N_19857,N_15168);
nor UO_943 (O_943,N_16578,N_17221);
xor UO_944 (O_944,N_17121,N_17858);
and UO_945 (O_945,N_17462,N_16456);
nor UO_946 (O_946,N_19133,N_17258);
and UO_947 (O_947,N_17483,N_18041);
xor UO_948 (O_948,N_15754,N_15467);
and UO_949 (O_949,N_17611,N_15922);
nand UO_950 (O_950,N_16949,N_18938);
nor UO_951 (O_951,N_17459,N_19510);
nor UO_952 (O_952,N_15512,N_15358);
or UO_953 (O_953,N_16229,N_19071);
or UO_954 (O_954,N_18442,N_18026);
nor UO_955 (O_955,N_19972,N_17848);
xor UO_956 (O_956,N_18515,N_17426);
nand UO_957 (O_957,N_17860,N_18197);
or UO_958 (O_958,N_15403,N_15738);
nor UO_959 (O_959,N_15283,N_19747);
xor UO_960 (O_960,N_15577,N_19488);
nor UO_961 (O_961,N_18997,N_19700);
or UO_962 (O_962,N_16341,N_16268);
or UO_963 (O_963,N_18929,N_18865);
nand UO_964 (O_964,N_19100,N_19799);
xnor UO_965 (O_965,N_15576,N_17362);
or UO_966 (O_966,N_19221,N_16985);
and UO_967 (O_967,N_15556,N_19277);
nand UO_968 (O_968,N_18352,N_19279);
or UO_969 (O_969,N_15775,N_19644);
nand UO_970 (O_970,N_15238,N_16817);
nor UO_971 (O_971,N_16727,N_17524);
xnor UO_972 (O_972,N_17952,N_15548);
nor UO_973 (O_973,N_18649,N_18410);
xnor UO_974 (O_974,N_16315,N_17778);
nor UO_975 (O_975,N_17278,N_18432);
and UO_976 (O_976,N_19339,N_18046);
nand UO_977 (O_977,N_18000,N_15213);
nor UO_978 (O_978,N_19929,N_15013);
or UO_979 (O_979,N_16057,N_17797);
xnor UO_980 (O_980,N_19830,N_18821);
nor UO_981 (O_981,N_18599,N_17905);
or UO_982 (O_982,N_15072,N_17716);
or UO_983 (O_983,N_15773,N_19467);
and UO_984 (O_984,N_19764,N_16565);
and UO_985 (O_985,N_18257,N_15108);
nand UO_986 (O_986,N_19062,N_18677);
xor UO_987 (O_987,N_15917,N_16561);
and UO_988 (O_988,N_19337,N_16234);
nor UO_989 (O_989,N_19464,N_18833);
and UO_990 (O_990,N_15849,N_18542);
and UO_991 (O_991,N_15836,N_18977);
and UO_992 (O_992,N_16309,N_19132);
and UO_993 (O_993,N_17194,N_17591);
and UO_994 (O_994,N_19019,N_16319);
nor UO_995 (O_995,N_15496,N_15227);
xor UO_996 (O_996,N_19158,N_19790);
or UO_997 (O_997,N_15876,N_17352);
xor UO_998 (O_998,N_16255,N_15123);
and UO_999 (O_999,N_19242,N_19060);
nor UO_1000 (O_1000,N_18486,N_18039);
and UO_1001 (O_1001,N_17594,N_19039);
and UO_1002 (O_1002,N_15262,N_17154);
xnor UO_1003 (O_1003,N_16794,N_15398);
and UO_1004 (O_1004,N_18167,N_17609);
and UO_1005 (O_1005,N_16182,N_19412);
xor UO_1006 (O_1006,N_18867,N_18792);
xnor UO_1007 (O_1007,N_18943,N_17302);
xnor UO_1008 (O_1008,N_16767,N_19129);
or UO_1009 (O_1009,N_19301,N_17754);
xor UO_1010 (O_1010,N_17967,N_17060);
xnor UO_1011 (O_1011,N_17384,N_16964);
nand UO_1012 (O_1012,N_19547,N_16028);
and UO_1013 (O_1013,N_16508,N_17882);
nor UO_1014 (O_1014,N_17208,N_18241);
or UO_1015 (O_1015,N_16937,N_19327);
or UO_1016 (O_1016,N_19163,N_15426);
nor UO_1017 (O_1017,N_19735,N_16620);
or UO_1018 (O_1018,N_16535,N_19185);
nor UO_1019 (O_1019,N_15931,N_17043);
and UO_1020 (O_1020,N_18941,N_19950);
xor UO_1021 (O_1021,N_16094,N_16021);
xor UO_1022 (O_1022,N_16769,N_17658);
nor UO_1023 (O_1023,N_17991,N_19366);
xnor UO_1024 (O_1024,N_18574,N_15897);
or UO_1025 (O_1025,N_18166,N_18745);
and UO_1026 (O_1026,N_16633,N_15727);
and UO_1027 (O_1027,N_16566,N_19662);
or UO_1028 (O_1028,N_16321,N_17118);
nor UO_1029 (O_1029,N_15074,N_17933);
or UO_1030 (O_1030,N_15678,N_17026);
xor UO_1031 (O_1031,N_17820,N_17849);
and UO_1032 (O_1032,N_15765,N_17507);
nand UO_1033 (O_1033,N_18999,N_19720);
nor UO_1034 (O_1034,N_16091,N_19037);
or UO_1035 (O_1035,N_17036,N_16646);
nor UO_1036 (O_1036,N_19641,N_18159);
nand UO_1037 (O_1037,N_18059,N_15482);
nand UO_1038 (O_1038,N_17295,N_18411);
or UO_1039 (O_1039,N_19993,N_16389);
nor UO_1040 (O_1040,N_15843,N_17557);
or UO_1041 (O_1041,N_18776,N_19647);
or UO_1042 (O_1042,N_19991,N_15580);
nor UO_1043 (O_1043,N_15642,N_19856);
nor UO_1044 (O_1044,N_19511,N_15085);
or UO_1045 (O_1045,N_15689,N_16026);
or UO_1046 (O_1046,N_18684,N_17122);
and UO_1047 (O_1047,N_15232,N_17403);
nor UO_1048 (O_1048,N_18233,N_16116);
or UO_1049 (O_1049,N_19708,N_17750);
nand UO_1050 (O_1050,N_18878,N_16153);
xnor UO_1051 (O_1051,N_15783,N_16922);
nand UO_1052 (O_1052,N_17590,N_18239);
or UO_1053 (O_1053,N_18921,N_15961);
xnor UO_1054 (O_1054,N_17102,N_18267);
xor UO_1055 (O_1055,N_16597,N_18907);
xor UO_1056 (O_1056,N_19678,N_19479);
nor UO_1057 (O_1057,N_16621,N_19858);
nor UO_1058 (O_1058,N_16612,N_19542);
and UO_1059 (O_1059,N_16746,N_16473);
and UO_1060 (O_1060,N_17442,N_17168);
xnor UO_1061 (O_1061,N_19502,N_15203);
nand UO_1062 (O_1062,N_16673,N_16227);
or UO_1063 (O_1063,N_15759,N_16301);
nor UO_1064 (O_1064,N_19915,N_18764);
or UO_1065 (O_1065,N_18374,N_19815);
nand UO_1066 (O_1066,N_18732,N_18578);
or UO_1067 (O_1067,N_15165,N_16115);
xnor UO_1068 (O_1068,N_16902,N_15609);
and UO_1069 (O_1069,N_15245,N_16370);
nand UO_1070 (O_1070,N_16659,N_16735);
xor UO_1071 (O_1071,N_19336,N_18956);
nand UO_1072 (O_1072,N_19006,N_19957);
nor UO_1073 (O_1073,N_17039,N_19556);
nand UO_1074 (O_1074,N_15004,N_16864);
xor UO_1075 (O_1075,N_17944,N_17268);
xnor UO_1076 (O_1076,N_16035,N_17783);
xnor UO_1077 (O_1077,N_15091,N_19638);
nand UO_1078 (O_1078,N_18512,N_16736);
or UO_1079 (O_1079,N_19854,N_17131);
nor UO_1080 (O_1080,N_19967,N_17559);
or UO_1081 (O_1081,N_17242,N_17885);
xnor UO_1082 (O_1082,N_16213,N_17799);
nand UO_1083 (O_1083,N_17271,N_18935);
nor UO_1084 (O_1084,N_18163,N_18853);
or UO_1085 (O_1085,N_16665,N_18187);
xor UO_1086 (O_1086,N_17350,N_19687);
nor UO_1087 (O_1087,N_15433,N_19978);
xnor UO_1088 (O_1088,N_19484,N_18036);
and UO_1089 (O_1089,N_16001,N_17150);
and UO_1090 (O_1090,N_17050,N_18779);
or UO_1091 (O_1091,N_15762,N_16499);
xor UO_1092 (O_1092,N_17634,N_17346);
nand UO_1093 (O_1093,N_19724,N_18818);
xnor UO_1094 (O_1094,N_17917,N_18635);
xnor UO_1095 (O_1095,N_18116,N_17830);
nand UO_1096 (O_1096,N_18087,N_18034);
and UO_1097 (O_1097,N_16891,N_15219);
xor UO_1098 (O_1098,N_16070,N_18890);
nor UO_1099 (O_1099,N_19809,N_18186);
and UO_1100 (O_1100,N_19157,N_15343);
or UO_1101 (O_1101,N_16324,N_17233);
and UO_1102 (O_1102,N_15106,N_17456);
and UO_1103 (O_1103,N_18675,N_16178);
xor UO_1104 (O_1104,N_19772,N_17990);
nand UO_1105 (O_1105,N_19513,N_17290);
xnor UO_1106 (O_1106,N_17618,N_16530);
and UO_1107 (O_1107,N_18407,N_17839);
nand UO_1108 (O_1108,N_15788,N_15326);
xnor UO_1109 (O_1109,N_16639,N_15337);
xor UO_1110 (O_1110,N_17482,N_15183);
nor UO_1111 (O_1111,N_16547,N_16519);
or UO_1112 (O_1112,N_17790,N_17441);
or UO_1113 (O_1113,N_18815,N_19240);
and UO_1114 (O_1114,N_17383,N_18139);
xor UO_1115 (O_1115,N_18381,N_18305);
xor UO_1116 (O_1116,N_19022,N_18001);
or UO_1117 (O_1117,N_15687,N_18856);
or UO_1118 (O_1118,N_16232,N_18443);
nor UO_1119 (O_1119,N_17685,N_15873);
or UO_1120 (O_1120,N_18198,N_17938);
xnor UO_1121 (O_1121,N_15612,N_17342);
or UO_1122 (O_1122,N_18178,N_15188);
or UO_1123 (O_1123,N_17491,N_18535);
and UO_1124 (O_1124,N_17791,N_16365);
nand UO_1125 (O_1125,N_17673,N_16826);
or UO_1126 (O_1126,N_15346,N_19231);
nor UO_1127 (O_1127,N_16123,N_18048);
nor UO_1128 (O_1128,N_15404,N_17851);
nor UO_1129 (O_1129,N_17151,N_15957);
or UO_1130 (O_1130,N_16629,N_17536);
nor UO_1131 (O_1131,N_15390,N_18895);
or UO_1132 (O_1132,N_19269,N_16588);
xor UO_1133 (O_1133,N_18014,N_19627);
nand UO_1134 (O_1134,N_16077,N_18570);
xnor UO_1135 (O_1135,N_17934,N_15278);
nor UO_1136 (O_1136,N_16852,N_18939);
and UO_1137 (O_1137,N_15866,N_18981);
nor UO_1138 (O_1138,N_18882,N_18088);
nand UO_1139 (O_1139,N_17219,N_16986);
and UO_1140 (O_1140,N_17907,N_16233);
or UO_1141 (O_1141,N_17364,N_15341);
nor UO_1142 (O_1142,N_19811,N_19819);
xor UO_1143 (O_1143,N_18314,N_18367);
xor UO_1144 (O_1144,N_19803,N_16958);
nor UO_1145 (O_1145,N_18206,N_18758);
and UO_1146 (O_1146,N_16418,N_15365);
nand UO_1147 (O_1147,N_15378,N_19224);
nor UO_1148 (O_1148,N_17167,N_18863);
xnor UO_1149 (O_1149,N_17575,N_15830);
nand UO_1150 (O_1150,N_17775,N_18285);
nor UO_1151 (O_1151,N_17499,N_16935);
or UO_1152 (O_1152,N_15000,N_17281);
or UO_1153 (O_1153,N_15176,N_19477);
nor UO_1154 (O_1154,N_17404,N_18517);
xor UO_1155 (O_1155,N_18357,N_17945);
xnor UO_1156 (O_1156,N_16071,N_16661);
xnor UO_1157 (O_1157,N_15553,N_17589);
xnor UO_1158 (O_1158,N_17065,N_16969);
nor UO_1159 (O_1159,N_19313,N_18906);
xor UO_1160 (O_1160,N_19591,N_19043);
or UO_1161 (O_1161,N_19732,N_17196);
xor UO_1162 (O_1162,N_18602,N_17336);
nand UO_1163 (O_1163,N_16032,N_18728);
nor UO_1164 (O_1164,N_17172,N_17954);
xnor UO_1165 (O_1165,N_18364,N_16377);
nand UO_1166 (O_1166,N_19227,N_15861);
nand UO_1167 (O_1167,N_18437,N_15583);
xnor UO_1168 (O_1168,N_19377,N_15571);
or UO_1169 (O_1169,N_18466,N_15173);
or UO_1170 (O_1170,N_19035,N_15109);
xnor UO_1171 (O_1171,N_15073,N_17040);
nor UO_1172 (O_1172,N_15036,N_18077);
or UO_1173 (O_1173,N_19651,N_16815);
nand UO_1174 (O_1174,N_15100,N_16102);
nor UO_1175 (O_1175,N_15466,N_19694);
and UO_1176 (O_1176,N_15507,N_19309);
and UO_1177 (O_1177,N_19543,N_15734);
or UO_1178 (O_1178,N_15570,N_18556);
or UO_1179 (O_1179,N_15942,N_15186);
and UO_1180 (O_1180,N_19435,N_18783);
nand UO_1181 (O_1181,N_16231,N_19682);
and UO_1182 (O_1182,N_18797,N_15562);
and UO_1183 (O_1183,N_19922,N_16851);
nand UO_1184 (O_1184,N_16441,N_19602);
nor UO_1185 (O_1185,N_17203,N_15177);
xor UO_1186 (O_1186,N_15131,N_16443);
and UO_1187 (O_1187,N_16195,N_17512);
or UO_1188 (O_1188,N_18124,N_15296);
and UO_1189 (O_1189,N_19282,N_17965);
or UO_1190 (O_1190,N_19117,N_16995);
nor UO_1191 (O_1191,N_16619,N_15847);
or UO_1192 (O_1192,N_15126,N_16570);
xor UO_1193 (O_1193,N_19589,N_15359);
xnor UO_1194 (O_1194,N_19272,N_17205);
and UO_1195 (O_1195,N_18598,N_16144);
nand UO_1196 (O_1196,N_15497,N_15726);
xnor UO_1197 (O_1197,N_19017,N_18562);
xnor UO_1198 (O_1198,N_18928,N_18645);
or UO_1199 (O_1199,N_15601,N_16459);
and UO_1200 (O_1200,N_18301,N_19259);
xor UO_1201 (O_1201,N_18708,N_17619);
nand UO_1202 (O_1202,N_17079,N_19792);
nand UO_1203 (O_1203,N_17722,N_19260);
xor UO_1204 (O_1204,N_15200,N_15694);
and UO_1205 (O_1205,N_18571,N_17178);
xnor UO_1206 (O_1206,N_17680,N_16058);
and UO_1207 (O_1207,N_17341,N_18905);
nor UO_1208 (O_1208,N_18577,N_15659);
and UO_1209 (O_1209,N_19754,N_17615);
nand UO_1210 (O_1210,N_19049,N_15774);
and UO_1211 (O_1211,N_18721,N_19382);
and UO_1212 (O_1212,N_18519,N_16311);
and UO_1213 (O_1213,N_19198,N_15704);
nor UO_1214 (O_1214,N_17215,N_15835);
nand UO_1215 (O_1215,N_17225,N_18714);
nand UO_1216 (O_1216,N_19855,N_18605);
or UO_1217 (O_1217,N_18092,N_16385);
or UO_1218 (O_1218,N_17539,N_17165);
xor UO_1219 (O_1219,N_18737,N_19522);
nand UO_1220 (O_1220,N_19052,N_18246);
or UO_1221 (O_1221,N_19579,N_15212);
xor UO_1222 (O_1222,N_16914,N_16192);
nor UO_1223 (O_1223,N_19894,N_19386);
xor UO_1224 (O_1224,N_15692,N_17100);
nor UO_1225 (O_1225,N_18270,N_15392);
xnor UO_1226 (O_1226,N_15303,N_16136);
nand UO_1227 (O_1227,N_17185,N_16778);
or UO_1228 (O_1228,N_15533,N_16850);
nor UO_1229 (O_1229,N_19331,N_15319);
and UO_1230 (O_1230,N_17029,N_16645);
nor UO_1231 (O_1231,N_16523,N_17811);
and UO_1232 (O_1232,N_19362,N_15516);
nand UO_1233 (O_1233,N_19215,N_17522);
nor UO_1234 (O_1234,N_18642,N_19506);
xnor UO_1235 (O_1235,N_19250,N_19024);
xnor UO_1236 (O_1236,N_19911,N_19462);
xnor UO_1237 (O_1237,N_15038,N_16264);
nor UO_1238 (O_1238,N_15832,N_19919);
nor UO_1239 (O_1239,N_15432,N_18228);
or UO_1240 (O_1240,N_15027,N_16890);
and UO_1241 (O_1241,N_16830,N_17222);
and UO_1242 (O_1242,N_19208,N_15055);
or UO_1243 (O_1243,N_15787,N_17056);
nand UO_1244 (O_1244,N_19156,N_19740);
and UO_1245 (O_1245,N_17766,N_19368);
or UO_1246 (O_1246,N_18217,N_19266);
and UO_1247 (O_1247,N_15190,N_15475);
or UO_1248 (O_1248,N_19986,N_17170);
or UO_1249 (O_1249,N_19608,N_17019);
xor UO_1250 (O_1250,N_15939,N_19392);
and UO_1251 (O_1251,N_18154,N_15452);
xnor UO_1252 (O_1252,N_17920,N_17827);
and UO_1253 (O_1253,N_16063,N_19356);
nor UO_1254 (O_1254,N_15518,N_18264);
and UO_1255 (O_1255,N_15083,N_17578);
nand UO_1256 (O_1256,N_18521,N_19875);
nand UO_1257 (O_1257,N_19791,N_15728);
xor UO_1258 (O_1258,N_17597,N_19228);
nand UO_1259 (O_1259,N_18685,N_17866);
nand UO_1260 (O_1260,N_17996,N_19214);
and UO_1261 (O_1261,N_18045,N_16191);
or UO_1262 (O_1262,N_16470,N_15667);
xnor UO_1263 (O_1263,N_16308,N_16055);
nor UO_1264 (O_1264,N_18028,N_17630);
nor UO_1265 (O_1265,N_19323,N_15592);
nor UO_1266 (O_1266,N_18185,N_18236);
nor UO_1267 (O_1267,N_18423,N_18487);
nor UO_1268 (O_1268,N_16511,N_16419);
xnor UO_1269 (O_1269,N_19051,N_18075);
nor UO_1270 (O_1270,N_15960,N_17374);
and UO_1271 (O_1271,N_18063,N_17224);
xnor UO_1272 (O_1272,N_18500,N_15082);
nand UO_1273 (O_1273,N_16824,N_19729);
and UO_1274 (O_1274,N_19758,N_18109);
nor UO_1275 (O_1275,N_15714,N_15947);
xnor UO_1276 (O_1276,N_17474,N_17187);
nor UO_1277 (O_1277,N_15118,N_19595);
or UO_1278 (O_1278,N_16860,N_18454);
nor UO_1279 (O_1279,N_18918,N_15119);
nor UO_1280 (O_1280,N_19042,N_15632);
nand UO_1281 (O_1281,N_15796,N_16776);
nand UO_1282 (O_1282,N_19239,N_15539);
nand UO_1283 (O_1283,N_19558,N_16181);
xor UO_1284 (O_1284,N_18495,N_15457);
and UO_1285 (O_1285,N_17856,N_16211);
xnor UO_1286 (O_1286,N_17010,N_17626);
xnor UO_1287 (O_1287,N_19106,N_18885);
nor UO_1288 (O_1288,N_15486,N_17016);
xor UO_1289 (O_1289,N_17051,N_19276);
and UO_1290 (O_1290,N_15174,N_19473);
xnor UO_1291 (O_1291,N_15872,N_16306);
xnor UO_1292 (O_1292,N_18811,N_16439);
nor UO_1293 (O_1293,N_17546,N_15672);
xor UO_1294 (O_1294,N_15952,N_15900);
and UO_1295 (O_1295,N_17427,N_18161);
xnor UO_1296 (O_1296,N_19517,N_17698);
xnor UO_1297 (O_1297,N_17889,N_18208);
nor UO_1298 (O_1298,N_19097,N_18951);
nor UO_1299 (O_1299,N_17505,N_15949);
or UO_1300 (O_1300,N_16781,N_17862);
nor UO_1301 (O_1301,N_17042,N_15669);
nor UO_1302 (O_1302,N_17470,N_19521);
nor UO_1303 (O_1303,N_19403,N_15618);
or UO_1304 (O_1304,N_19031,N_18333);
or UO_1305 (O_1305,N_17238,N_15982);
or UO_1306 (O_1306,N_19582,N_17488);
nor UO_1307 (O_1307,N_19300,N_16154);
nand UO_1308 (O_1308,N_17191,N_17418);
or UO_1309 (O_1309,N_18076,N_15741);
xor UO_1310 (O_1310,N_19077,N_16360);
or UO_1311 (O_1311,N_15009,N_15355);
xnor UO_1312 (O_1312,N_17854,N_18112);
xor UO_1313 (O_1313,N_15582,N_19020);
nor UO_1314 (O_1314,N_17845,N_15739);
nor UO_1315 (O_1315,N_17340,N_18898);
xnor UO_1316 (O_1316,N_19286,N_19734);
and UO_1317 (O_1317,N_18237,N_16509);
nor UO_1318 (O_1318,N_19625,N_17608);
and UO_1319 (O_1319,N_15546,N_18871);
and UO_1320 (O_1320,N_17639,N_18604);
nor UO_1321 (O_1321,N_17084,N_16138);
nand UO_1322 (O_1322,N_17959,N_16976);
or UO_1323 (O_1323,N_16029,N_18176);
nor UO_1324 (O_1324,N_18957,N_19460);
nor UO_1325 (O_1325,N_15794,N_18302);
and UO_1326 (O_1326,N_15948,N_18953);
or UO_1327 (O_1327,N_18224,N_18204);
nand UO_1328 (O_1328,N_18288,N_19273);
nor UO_1329 (O_1329,N_17478,N_15097);
or UO_1330 (O_1330,N_19737,N_15137);
or UO_1331 (O_1331,N_19933,N_16842);
or UO_1332 (O_1332,N_18632,N_19657);
and UO_1333 (O_1333,N_16478,N_18945);
xnor UO_1334 (O_1334,N_16348,N_16318);
or UO_1335 (O_1335,N_17720,N_15995);
nor UO_1336 (O_1336,N_19860,N_18253);
nor UO_1337 (O_1337,N_17678,N_16999);
and UO_1338 (O_1338,N_19316,N_15444);
and UO_1339 (O_1339,N_17492,N_19021);
nand UO_1340 (O_1340,N_19036,N_16910);
and UO_1341 (O_1341,N_16682,N_18435);
xnor UO_1342 (O_1342,N_17518,N_15941);
xnor UO_1343 (O_1343,N_17735,N_16121);
xor UO_1344 (O_1344,N_19162,N_16145);
xor UO_1345 (O_1345,N_19192,N_17002);
nand UO_1346 (O_1346,N_18385,N_18144);
and UO_1347 (O_1347,N_17311,N_15980);
xor UO_1348 (O_1348,N_15483,N_18456);
xnor UO_1349 (O_1349,N_17555,N_15455);
and UO_1350 (O_1350,N_15650,N_16052);
nand UO_1351 (O_1351,N_16766,N_19469);
nor UO_1352 (O_1352,N_18510,N_15827);
nor UO_1353 (O_1353,N_16079,N_19495);
and UO_1354 (O_1354,N_16518,N_15492);
and UO_1355 (O_1355,N_16128,N_18593);
xnor UO_1356 (O_1356,N_16599,N_15151);
nand UO_1357 (O_1357,N_17509,N_15101);
xor UO_1358 (O_1358,N_17504,N_15324);
nand UO_1359 (O_1359,N_16279,N_17455);
and UO_1360 (O_1360,N_17429,N_15766);
xor UO_1361 (O_1361,N_16688,N_18765);
nor UO_1362 (O_1362,N_19061,N_15400);
and UO_1363 (O_1363,N_18361,N_16946);
xor UO_1364 (O_1364,N_17166,N_17613);
nor UO_1365 (O_1365,N_15702,N_18780);
and UO_1366 (O_1366,N_18142,N_19365);
nor UO_1367 (O_1367,N_15023,N_16942);
nor UO_1368 (O_1368,N_17624,N_19016);
nor UO_1369 (O_1369,N_19319,N_16457);
or UO_1370 (O_1370,N_15638,N_16881);
xor UO_1371 (O_1371,N_19278,N_18425);
nand UO_1372 (O_1372,N_18540,N_15709);
nand UO_1373 (O_1373,N_15080,N_18592);
or UO_1374 (O_1374,N_17415,N_16358);
nor UO_1375 (O_1375,N_16532,N_15431);
nand UO_1376 (O_1376,N_19345,N_19428);
and UO_1377 (O_1377,N_17270,N_15332);
and UO_1378 (O_1378,N_19824,N_19545);
xor UO_1379 (O_1379,N_18717,N_17096);
nand UO_1380 (O_1380,N_17568,N_17140);
nand UO_1381 (O_1381,N_15690,N_15041);
xnor UO_1382 (O_1382,N_19490,N_17562);
xnor UO_1383 (O_1383,N_17644,N_18705);
xnor UO_1384 (O_1384,N_16734,N_15351);
xnor UO_1385 (O_1385,N_17554,N_15007);
and UO_1386 (O_1386,N_18729,N_16391);
xor UO_1387 (O_1387,N_16677,N_17516);
xnor UO_1388 (O_1388,N_19569,N_16738);
and UO_1389 (O_1389,N_15804,N_16122);
nor UO_1390 (O_1390,N_17057,N_19449);
and UO_1391 (O_1391,N_15924,N_18448);
nor UO_1392 (O_1392,N_17239,N_17062);
nor UO_1393 (O_1393,N_16722,N_19552);
and UO_1394 (O_1394,N_18822,N_16353);
and UO_1395 (O_1395,N_16327,N_19670);
and UO_1396 (O_1396,N_18844,N_19573);
nand UO_1397 (O_1397,N_19390,N_17865);
nand UO_1398 (O_1398,N_17746,N_19620);
or UO_1399 (O_1399,N_15473,N_15798);
nor UO_1400 (O_1400,N_19937,N_18399);
or UO_1401 (O_1401,N_15162,N_19590);
xnor UO_1402 (O_1402,N_16836,N_17558);
xor UO_1403 (O_1403,N_16038,N_16887);
and UO_1404 (O_1404,N_15293,N_16270);
nor UO_1405 (O_1405,N_17412,N_17054);
nand UO_1406 (O_1406,N_19090,N_17870);
and UO_1407 (O_1407,N_16502,N_15450);
nor UO_1408 (O_1408,N_15673,N_18145);
or UO_1409 (O_1409,N_17430,N_15663);
and UO_1410 (O_1410,N_17844,N_16034);
or UO_1411 (O_1411,N_17838,N_15427);
or UO_1412 (O_1412,N_19126,N_15286);
xor UO_1413 (O_1413,N_16256,N_19481);
nand UO_1414 (O_1414,N_18558,N_18502);
or UO_1415 (O_1415,N_16125,N_17436);
or UO_1416 (O_1416,N_19415,N_18365);
or UO_1417 (O_1417,N_18254,N_18091);
xnor UO_1418 (O_1418,N_18297,N_15608);
nand UO_1419 (O_1419,N_18657,N_16854);
xnor UO_1420 (O_1420,N_16206,N_18240);
or UO_1421 (O_1421,N_16638,N_15621);
xor UO_1422 (O_1422,N_18829,N_18787);
nand UO_1423 (O_1423,N_16291,N_18037);
xnor UO_1424 (O_1424,N_19312,N_16580);
or UO_1425 (O_1425,N_17674,N_15316);
nor UO_1426 (O_1426,N_15833,N_16294);
nand UO_1427 (O_1427,N_18114,N_17873);
xnor UO_1428 (O_1428,N_15888,N_15053);
xor UO_1429 (O_1429,N_16163,N_17330);
xor UO_1430 (O_1430,N_15383,N_15035);
nand UO_1431 (O_1431,N_19969,N_18079);
nand UO_1432 (O_1432,N_15731,N_19879);
and UO_1433 (O_1433,N_16208,N_18886);
xnor UO_1434 (O_1434,N_15713,N_15743);
nor UO_1435 (O_1435,N_18064,N_15600);
nor UO_1436 (O_1436,N_17574,N_19797);
nand UO_1437 (O_1437,N_17857,N_15049);
and UO_1438 (O_1438,N_18555,N_18630);
nor UO_1439 (O_1439,N_19504,N_17072);
nor UO_1440 (O_1440,N_15150,N_15525);
nand UO_1441 (O_1441,N_19014,N_18330);
nor UO_1442 (O_1442,N_17041,N_15089);
xor UO_1443 (O_1443,N_18749,N_16582);
xnor UO_1444 (O_1444,N_19094,N_19932);
nor UO_1445 (O_1445,N_15675,N_16283);
nor UO_1446 (O_1446,N_19393,N_16169);
and UO_1447 (O_1447,N_18207,N_17895);
and UO_1448 (O_1448,N_16671,N_15078);
nand UO_1449 (O_1449,N_18281,N_15305);
nor UO_1450 (O_1450,N_17493,N_18960);
and UO_1451 (O_1451,N_18324,N_17897);
or UO_1452 (O_1452,N_18607,N_18220);
nor UO_1453 (O_1453,N_17642,N_19876);
nand UO_1454 (O_1454,N_16558,N_17919);
and UO_1455 (O_1455,N_18356,N_19667);
nor UO_1456 (O_1456,N_17623,N_15285);
nand UO_1457 (O_1457,N_16737,N_16396);
nand UO_1458 (O_1458,N_19391,N_19763);
or UO_1459 (O_1459,N_17560,N_15311);
nor UO_1460 (O_1460,N_15655,N_17267);
xnor UO_1461 (O_1461,N_16299,N_16080);
and UO_1462 (O_1462,N_16189,N_18925);
xor UO_1463 (O_1463,N_16263,N_18481);
xor UO_1464 (O_1464,N_17162,N_19541);
or UO_1465 (O_1465,N_15045,N_19606);
xnor UO_1466 (O_1466,N_19232,N_16950);
nand UO_1467 (O_1467,N_17282,N_19104);
nor UO_1468 (O_1468,N_18926,N_19818);
xnor UO_1469 (O_1469,N_17334,N_16160);
xor UO_1470 (O_1470,N_15249,N_17683);
nor UO_1471 (O_1471,N_15121,N_16708);
and UO_1472 (O_1472,N_15320,N_16505);
nand UO_1473 (O_1473,N_15374,N_17928);
nor UO_1474 (O_1474,N_15328,N_17437);
and UO_1475 (O_1475,N_19190,N_17661);
nor UO_1476 (O_1476,N_16898,N_16728);
or UO_1477 (O_1477,N_16686,N_18353);
nor UO_1478 (O_1478,N_19322,N_19027);
or UO_1479 (O_1479,N_15476,N_16590);
and UO_1480 (O_1480,N_17460,N_17706);
nand UO_1481 (O_1481,N_17073,N_15304);
nand UO_1482 (O_1482,N_16262,N_17182);
or UO_1483 (O_1483,N_15997,N_17034);
and UO_1484 (O_1484,N_19750,N_15500);
nor UO_1485 (O_1485,N_16959,N_18741);
xor UO_1486 (O_1486,N_18524,N_15883);
nand UO_1487 (O_1487,N_17067,N_16042);
or UO_1488 (O_1488,N_17393,N_15348);
nor UO_1489 (O_1489,N_19663,N_18030);
nor UO_1490 (O_1490,N_17729,N_16185);
nand UO_1491 (O_1491,N_15740,N_16643);
nor UO_1492 (O_1492,N_17183,N_19034);
nor UO_1493 (O_1493,N_16241,N_15620);
xor UO_1494 (O_1494,N_17230,N_15845);
or UO_1495 (O_1495,N_16966,N_19848);
xnor UO_1496 (O_1496,N_16376,N_19778);
xor UO_1497 (O_1497,N_16610,N_18796);
and UO_1498 (O_1498,N_17484,N_15607);
nand UO_1499 (O_1499,N_18150,N_16247);
nor UO_1500 (O_1500,N_16750,N_16527);
or UO_1501 (O_1501,N_16161,N_18089);
and UO_1502 (O_1502,N_15662,N_17031);
or UO_1503 (O_1503,N_18434,N_17663);
xnor UO_1504 (O_1504,N_17038,N_19585);
nor UO_1505 (O_1505,N_16552,N_16082);
or UO_1506 (O_1506,N_16867,N_17776);
and UO_1507 (O_1507,N_19497,N_17013);
xor UO_1508 (O_1508,N_17741,N_18165);
or UO_1509 (O_1509,N_15495,N_16249);
xnor UO_1510 (O_1510,N_18184,N_16967);
and UO_1511 (O_1511,N_19701,N_17940);
xnor UO_1512 (O_1512,N_17252,N_16939);
or UO_1513 (O_1513,N_16197,N_16451);
nand UO_1514 (O_1514,N_17320,N_18004);
nand UO_1515 (O_1515,N_16274,N_18476);
and UO_1516 (O_1516,N_19683,N_19064);
or UO_1517 (O_1517,N_18606,N_15008);
or UO_1518 (O_1518,N_19883,N_18308);
xnor UO_1519 (O_1519,N_17132,N_15764);
nor UO_1520 (O_1520,N_18627,N_17691);
and UO_1521 (O_1521,N_18249,N_18130);
nand UO_1522 (O_1522,N_15393,N_16838);
xor UO_1523 (O_1523,N_19140,N_16944);
and UO_1524 (O_1524,N_18998,N_19095);
or UO_1525 (O_1525,N_17796,N_19130);
xor UO_1526 (O_1526,N_16463,N_18148);
nor UO_1527 (O_1527,N_15116,N_19475);
xnor UO_1528 (O_1528,N_18483,N_15975);
xor UO_1529 (O_1529,N_18379,N_19152);
nor UO_1530 (O_1530,N_19653,N_17390);
nand UO_1531 (O_1531,N_17548,N_16440);
nor UO_1532 (O_1532,N_17532,N_15155);
xor UO_1533 (O_1533,N_16111,N_15191);
and UO_1534 (O_1534,N_18731,N_15629);
xor UO_1535 (O_1535,N_17237,N_15020);
and UO_1536 (O_1536,N_16167,N_19528);
nand UO_1537 (O_1537,N_15408,N_17345);
and UO_1538 (O_1538,N_17689,N_19779);
and UO_1539 (O_1539,N_17137,N_15908);
or UO_1540 (O_1540,N_15292,N_18855);
xor UO_1541 (O_1541,N_15567,N_15831);
or UO_1542 (O_1542,N_19509,N_18923);
or UO_1543 (O_1543,N_19452,N_18445);
and UO_1544 (O_1544,N_16097,N_17710);
nor UO_1545 (O_1545,N_18771,N_18631);
nand UO_1546 (O_1546,N_18719,N_16388);
nor UO_1547 (O_1547,N_19399,N_19938);
xor UO_1548 (O_1548,N_19789,N_16541);
xor UO_1549 (O_1549,N_17304,N_16548);
xor UO_1550 (O_1550,N_17520,N_15409);
nand UO_1551 (O_1551,N_16488,N_19165);
xnor UO_1552 (O_1552,N_18484,N_19480);
xor UO_1553 (O_1553,N_15018,N_15974);
xnor UO_1554 (O_1554,N_18993,N_18029);
nor UO_1555 (O_1555,N_19598,N_18420);
or UO_1556 (O_1556,N_16829,N_18106);
and UO_1557 (O_1557,N_16760,N_18734);
xor UO_1558 (O_1558,N_17163,N_15898);
and UO_1559 (O_1559,N_15299,N_16790);
and UO_1560 (O_1560,N_17773,N_17533);
and UO_1561 (O_1561,N_15723,N_15417);
or UO_1562 (O_1562,N_19026,N_17877);
or UO_1563 (O_1563,N_15622,N_16586);
and UO_1564 (O_1564,N_16663,N_15223);
or UO_1565 (O_1565,N_16258,N_19661);
nor UO_1566 (O_1566,N_18090,N_16217);
and UO_1567 (O_1567,N_18482,N_15935);
nor UO_1568 (O_1568,N_18272,N_19394);
and UO_1569 (O_1569,N_17653,N_16500);
nor UO_1570 (O_1570,N_18572,N_17659);
xor UO_1571 (O_1571,N_15626,N_15391);
xnor UO_1572 (O_1572,N_19753,N_18460);
nor UO_1573 (O_1573,N_18987,N_16236);
xor UO_1574 (O_1574,N_18424,N_15768);
or UO_1575 (O_1575,N_17006,N_19713);
xnor UO_1576 (O_1576,N_19767,N_19702);
xor UO_1577 (O_1577,N_17657,N_18747);
nand UO_1578 (O_1578,N_19204,N_16513);
nor UO_1579 (O_1579,N_15161,N_17424);
and UO_1580 (O_1580,N_16432,N_17620);
nand UO_1581 (O_1581,N_15153,N_15599);
or UO_1582 (O_1582,N_17055,N_17807);
xor UO_1583 (O_1583,N_16918,N_16697);
xor UO_1584 (O_1584,N_18545,N_15071);
nor UO_1585 (O_1585,N_17821,N_19512);
nand UO_1586 (O_1586,N_19888,N_15752);
nand UO_1587 (O_1587,N_17501,N_19124);
xnor UO_1588 (O_1588,N_17082,N_17910);
nand UO_1589 (O_1589,N_18661,N_19128);
nor UO_1590 (O_1590,N_19973,N_18852);
or UO_1591 (O_1591,N_16290,N_15103);
nand UO_1592 (O_1592,N_18722,N_19746);
nor UO_1593 (O_1593,N_15254,N_15224);
or UO_1594 (O_1594,N_18095,N_15284);
nand UO_1595 (O_1595,N_18174,N_17094);
xor UO_1596 (O_1596,N_16948,N_19984);
nor UO_1597 (O_1597,N_18564,N_17236);
nand UO_1598 (O_1598,N_17469,N_19099);
xnor UO_1599 (O_1599,N_17982,N_16371);
nor UO_1600 (O_1600,N_18155,N_15617);
nand UO_1601 (O_1601,N_19253,N_16810);
nand UO_1602 (O_1602,N_19806,N_18438);
xor UO_1603 (O_1603,N_16689,N_15624);
or UO_1604 (O_1604,N_16180,N_19098);
or UO_1605 (O_1605,N_15606,N_18896);
xor UO_1606 (O_1606,N_16460,N_16598);
and UO_1607 (O_1607,N_18824,N_16819);
and UO_1608 (O_1608,N_18202,N_19916);
xor UO_1609 (O_1609,N_19182,N_18491);
and UO_1610 (O_1610,N_16183,N_15001);
or UO_1611 (O_1611,N_17251,N_15396);
and UO_1612 (O_1612,N_16096,N_15336);
nor UO_1613 (O_1613,N_16317,N_15986);
or UO_1614 (O_1614,N_19025,N_15478);
nand UO_1615 (O_1615,N_16225,N_19154);
nand UO_1616 (O_1616,N_19196,N_16168);
or UO_1617 (O_1617,N_15885,N_16710);
and UO_1618 (O_1618,N_17328,N_19604);
nand UO_1619 (O_1619,N_15850,N_17682);
and UO_1620 (O_1620,N_15462,N_15598);
nor UO_1621 (O_1621,N_18398,N_16744);
nor UO_1622 (O_1622,N_16712,N_18600);
xnor UO_1623 (O_1623,N_17045,N_15260);
xor UO_1624 (O_1624,N_16600,N_16845);
xor UO_1625 (O_1625,N_19069,N_19407);
or UO_1626 (O_1626,N_19924,N_17987);
or UO_1627 (O_1627,N_15387,N_17631);
nand UO_1628 (O_1628,N_16277,N_15170);
nand UO_1629 (O_1629,N_17325,N_16589);
nand UO_1630 (O_1630,N_18211,N_18418);
nor UO_1631 (O_1631,N_18707,N_17898);
nand UO_1632 (O_1632,N_18182,N_17593);
xnor UO_1633 (O_1633,N_18169,N_16075);
or UO_1634 (O_1634,N_19015,N_15869);
nor UO_1635 (O_1635,N_19320,N_17969);
and UO_1636 (O_1636,N_17625,N_18380);
nand UO_1637 (O_1637,N_17822,N_15903);
nand UO_1638 (O_1638,N_17148,N_15345);
and UO_1639 (O_1639,N_17086,N_19655);
nand UO_1640 (O_1640,N_19675,N_16834);
and UO_1641 (O_1641,N_18698,N_15584);
and UO_1642 (O_1642,N_18084,N_18038);
or UO_1643 (O_1643,N_16222,N_16156);
and UO_1644 (O_1644,N_18828,N_17974);
or UO_1645 (O_1645,N_16207,N_16908);
or UO_1646 (O_1646,N_17641,N_15234);
or UO_1647 (O_1647,N_19529,N_18485);
or UO_1648 (O_1648,N_19147,N_15156);
nand UO_1649 (O_1649,N_18516,N_15350);
nor UO_1650 (O_1650,N_18269,N_19942);
nand UO_1651 (O_1651,N_18769,N_17179);
xor UO_1652 (O_1652,N_17941,N_15095);
xor UO_1653 (O_1653,N_18342,N_19951);
or UO_1654 (O_1654,N_17145,N_16951);
nand UO_1655 (O_1655,N_16108,N_18054);
or UO_1656 (O_1656,N_19298,N_16863);
xor UO_1657 (O_1657,N_19187,N_16447);
nand UO_1658 (O_1658,N_18119,N_15522);
nor UO_1659 (O_1659,N_16632,N_15333);
and UO_1660 (O_1660,N_18785,N_15801);
or UO_1661 (O_1661,N_19801,N_19897);
nor UO_1662 (O_1662,N_16151,N_17379);
nor UO_1663 (O_1663,N_19766,N_19419);
and UO_1664 (O_1664,N_19344,N_18566);
nor UO_1665 (O_1665,N_19889,N_16027);
or UO_1666 (O_1666,N_15893,N_17984);
nand UO_1667 (O_1667,N_19048,N_17645);
xor UO_1668 (O_1668,N_17453,N_18810);
and UO_1669 (O_1669,N_16048,N_17784);
nor UO_1670 (O_1670,N_16868,N_17111);
nand UO_1671 (O_1671,N_17216,N_17466);
nand UO_1672 (O_1672,N_19293,N_17964);
nand UO_1673 (O_1673,N_16521,N_17770);
or UO_1674 (O_1674,N_19877,N_18473);
and UO_1675 (O_1675,N_19592,N_17018);
nor UO_1676 (O_1676,N_15414,N_17529);
and UO_1677 (O_1677,N_19013,N_18641);
and UO_1678 (O_1678,N_16618,N_16878);
and UO_1679 (O_1679,N_15194,N_17947);
xnor UO_1680 (O_1680,N_15757,N_15981);
nand UO_1681 (O_1681,N_17454,N_17035);
xor UO_1682 (O_1682,N_16293,N_16332);
or UO_1683 (O_1683,N_17709,N_19795);
and UO_1684 (O_1684,N_15932,N_19576);
nand UO_1685 (O_1685,N_18565,N_16931);
and UO_1686 (O_1686,N_16719,N_16285);
xnor UO_1687 (O_1687,N_18250,N_18287);
nand UO_1688 (O_1688,N_18151,N_16818);
nor UO_1689 (O_1689,N_17255,N_19955);
and UO_1690 (O_1690,N_15758,N_19169);
xnor UO_1691 (O_1691,N_15469,N_17955);
or UO_1692 (O_1692,N_15034,N_19263);
or UO_1693 (O_1693,N_18339,N_16803);
xor UO_1694 (O_1694,N_16877,N_18222);
nand UO_1695 (O_1695,N_17126,N_19527);
nor UO_1696 (O_1696,N_16148,N_18060);
nor UO_1697 (O_1697,N_16707,N_15613);
xor UO_1698 (O_1698,N_15776,N_16450);
or UO_1699 (O_1699,N_15209,N_16989);
nor UO_1700 (O_1700,N_16853,N_18814);
nor UO_1701 (O_1701,N_19596,N_17842);
or UO_1702 (O_1702,N_15544,N_19553);
xnor UO_1703 (O_1703,N_19762,N_17929);
and UO_1704 (O_1704,N_18768,N_16310);
xor UO_1705 (O_1705,N_16953,N_16399);
xnor UO_1706 (O_1706,N_15329,N_18813);
nor UO_1707 (O_1707,N_16674,N_18868);
and UO_1708 (O_1708,N_18351,N_17420);
nand UO_1709 (O_1709,N_16173,N_16667);
or UO_1710 (O_1710,N_16886,N_15792);
and UO_1711 (O_1711,N_17667,N_18704);
and UO_1712 (O_1712,N_16050,N_16833);
and UO_1713 (O_1713,N_18919,N_16932);
or UO_1714 (O_1714,N_19551,N_15060);
nor UO_1715 (O_1715,N_19491,N_15357);
or UO_1716 (O_1716,N_17396,N_18802);
nand UO_1717 (O_1717,N_16127,N_18471);
nor UO_1718 (O_1718,N_16468,N_19011);
or UO_1719 (O_1719,N_18849,N_19110);
nor UO_1720 (O_1720,N_18597,N_16237);
and UO_1721 (O_1721,N_18643,N_16595);
and UO_1722 (O_1722,N_18975,N_19318);
or UO_1723 (O_1723,N_19305,N_16414);
or UO_1724 (O_1724,N_17108,N_16060);
nor UO_1725 (O_1725,N_19900,N_18325);
and UO_1726 (O_1726,N_18322,N_18347);
nand UO_1727 (O_1727,N_16514,N_15543);
or UO_1728 (O_1728,N_17760,N_17032);
nand UO_1729 (O_1729,N_18055,N_15646);
or UO_1730 (O_1730,N_15521,N_19567);
nand UO_1731 (O_1731,N_16651,N_19852);
nor UO_1732 (O_1732,N_18143,N_17337);
nor UO_1733 (O_1733,N_16069,N_19308);
xnor UO_1734 (O_1734,N_16624,N_15066);
nand UO_1735 (O_1735,N_18426,N_17446);
nor UO_1736 (O_1736,N_16880,N_15465);
nand UO_1737 (O_1737,N_19223,N_18760);
and UO_1738 (O_1738,N_19560,N_17537);
nand UO_1739 (O_1739,N_17884,N_17981);
nand UO_1740 (O_1740,N_16303,N_19652);
nand UO_1741 (O_1741,N_19963,N_18362);
nor UO_1742 (O_1742,N_19468,N_15215);
and UO_1743 (O_1743,N_16364,N_16392);
nor UO_1744 (O_1744,N_16593,N_19752);
and UO_1745 (O_1745,N_18986,N_18480);
xnor UO_1746 (O_1746,N_18417,N_17371);
xor UO_1747 (O_1747,N_15654,N_19643);
nor UO_1748 (O_1748,N_18205,N_16960);
and UO_1749 (O_1749,N_16941,N_16921);
nand UO_1750 (O_1750,N_17472,N_18876);
nand UO_1751 (O_1751,N_17135,N_16101);
nor UO_1752 (O_1752,N_17695,N_18180);
and UO_1753 (O_1753,N_17573,N_17892);
and UO_1754 (O_1754,N_16625,N_17902);
or UO_1755 (O_1755,N_15189,N_19623);
xor UO_1756 (O_1756,N_16188,N_15693);
and UO_1757 (O_1757,N_16839,N_19429);
and UO_1758 (O_1758,N_19672,N_19500);
xor UO_1759 (O_1759,N_16347,N_19539);
nand UO_1760 (O_1760,N_15255,N_18319);
or UO_1761 (O_1761,N_15563,N_16464);
nor UO_1762 (O_1762,N_15006,N_16991);
and UO_1763 (O_1763,N_19562,N_19478);
and UO_1764 (O_1764,N_17248,N_15707);
nor UO_1765 (O_1765,N_19203,N_19930);
or UO_1766 (O_1766,N_19050,N_16748);
nor UO_1767 (O_1767,N_15547,N_17814);
nand UO_1768 (O_1768,N_19699,N_18120);
nor UO_1769 (O_1769,N_16806,N_17565);
or UO_1770 (O_1770,N_19736,N_16702);
and UO_1771 (O_1771,N_18752,N_16544);
and UO_1772 (O_1772,N_15456,N_15943);
xor UO_1773 (O_1773,N_17253,N_16329);
or UO_1774 (O_1774,N_15852,N_16220);
nand UO_1775 (O_1775,N_15820,N_17728);
nand UO_1776 (O_1776,N_18875,N_18094);
or UO_1777 (O_1777,N_19296,N_17308);
xor UO_1778 (O_1778,N_16971,N_18294);
nand UO_1779 (O_1779,N_18003,N_16384);
nor UO_1780 (O_1780,N_19115,N_18843);
and UO_1781 (O_1781,N_19383,N_17133);
nand UO_1782 (O_1782,N_16785,N_19712);
or UO_1783 (O_1783,N_19676,N_15022);
or UO_1784 (O_1784,N_19563,N_15154);
or UO_1785 (O_1785,N_19640,N_18669);
nor UO_1786 (O_1786,N_18404,N_16516);
nor UO_1787 (O_1787,N_18274,N_18671);
nor UO_1788 (O_1788,N_16896,N_17277);
nand UO_1789 (O_1789,N_15318,N_17171);
nand UO_1790 (O_1790,N_15207,N_16438);
xor UO_1791 (O_1791,N_19324,N_18140);
and UO_1792 (O_1792,N_18290,N_18025);
nand UO_1793 (O_1793,N_19570,N_18020);
and UO_1794 (O_1794,N_16476,N_15541);
and UO_1795 (O_1795,N_19456,N_19499);
or UO_1796 (O_1796,N_16540,N_18608);
xor UO_1797 (O_1797,N_15354,N_16172);
or UO_1798 (O_1798,N_17879,N_16893);
or UO_1799 (O_1799,N_16996,N_19029);
xor UO_1800 (O_1800,N_18080,N_18086);
xnor UO_1801 (O_1801,N_19354,N_15973);
or UO_1802 (O_1802,N_17909,N_17714);
or UO_1803 (O_1803,N_17640,N_18479);
and UO_1804 (O_1804,N_17744,N_15179);
or UO_1805 (O_1805,N_16342,N_19680);
xor UO_1806 (O_1806,N_16492,N_17815);
xnor UO_1807 (O_1807,N_15880,N_16009);
xnor UO_1808 (O_1808,N_17092,N_17265);
and UO_1809 (O_1809,N_16313,N_16704);
nor UO_1810 (O_1810,N_16496,N_19173);
nor UO_1811 (O_1811,N_17939,N_17475);
nor UO_1812 (O_1812,N_18615,N_18503);
nor UO_1813 (O_1813,N_15314,N_16489);
nor UO_1814 (O_1814,N_19474,N_15334);
nand UO_1815 (O_1815,N_16517,N_15268);
nand UO_1816 (O_1816,N_19624,N_17292);
nand UO_1817 (O_1817,N_19715,N_19448);
xor UO_1818 (O_1818,N_19144,N_18133);
nor UO_1819 (O_1819,N_19361,N_18157);
and UO_1820 (O_1820,N_16498,N_15090);
and UO_1821 (O_1821,N_19634,N_18880);
and UO_1822 (O_1822,N_15703,N_18283);
and UO_1823 (O_1823,N_18421,N_15715);
xor UO_1824 (O_1824,N_19180,N_16393);
xnor UO_1825 (O_1825,N_15859,N_18983);
xnor UO_1826 (O_1826,N_17983,N_19325);
or UO_1827 (O_1827,N_18766,N_17723);
xnor UO_1828 (O_1828,N_17012,N_17666);
nor UO_1829 (O_1829,N_19405,N_16930);
nand UO_1830 (O_1830,N_18934,N_18840);
nor UO_1831 (O_1831,N_19669,N_17105);
and UO_1832 (O_1832,N_16792,N_17616);
and UO_1833 (O_1833,N_16085,N_17913);
nor UO_1834 (O_1834,N_19353,N_16462);
xnor UO_1835 (O_1835,N_16992,N_19451);
and UO_1836 (O_1836,N_15241,N_19341);
or UO_1837 (O_1837,N_19175,N_19290);
xnor UO_1838 (O_1838,N_18899,N_18933);
nand UO_1839 (O_1839,N_16198,N_17878);
xnor UO_1840 (O_1840,N_16461,N_19402);
nand UO_1841 (O_1841,N_18040,N_18892);
xnor UO_1842 (O_1842,N_19749,N_16979);
or UO_1843 (O_1843,N_18836,N_17571);
nand UO_1844 (O_1844,N_19827,N_19445);
nor UO_1845 (O_1845,N_19996,N_17144);
xnor UO_1846 (O_1846,N_15818,N_16269);
nand UO_1847 (O_1847,N_18634,N_19145);
nand UO_1848 (O_1848,N_19775,N_17828);
and UO_1849 (O_1849,N_19943,N_18194);
nand UO_1850 (O_1850,N_15991,N_18511);
nand UO_1851 (O_1851,N_17900,N_17047);
nor UO_1852 (O_1852,N_16187,N_15129);
nor UO_1853 (O_1853,N_15971,N_15266);
or UO_1854 (O_1854,N_17961,N_17686);
nor UO_1855 (O_1855,N_17448,N_15081);
nor UO_1856 (O_1856,N_17063,N_17958);
or UO_1857 (O_1857,N_17717,N_15413);
or UO_1858 (O_1858,N_18795,N_19297);
nand UO_1859 (O_1859,N_19612,N_19524);
nor UO_1860 (O_1860,N_16025,N_19164);
nor UO_1861 (O_1861,N_19742,N_15046);
xnor UO_1862 (O_1862,N_17110,N_15744);
and UO_1863 (O_1863,N_18924,N_18431);
and UO_1864 (O_1864,N_17017,N_18544);
and UO_1865 (O_1865,N_16219,N_19113);
and UO_1866 (O_1866,N_15211,N_17743);
or UO_1867 (O_1867,N_16201,N_15956);
nand UO_1868 (O_1868,N_15136,N_18573);
nand UO_1869 (O_1869,N_17780,N_17831);
xnor UO_1870 (O_1870,N_18586,N_15605);
and UO_1871 (O_1871,N_19166,N_19887);
and UO_1872 (O_1872,N_15862,N_19611);
nand UO_1873 (O_1873,N_19526,N_18390);
nand UO_1874 (O_1874,N_17075,N_19826);
xnor UO_1875 (O_1875,N_16486,N_18847);
and UO_1876 (O_1876,N_17726,N_17331);
and UO_1877 (O_1877,N_19892,N_18428);
xnor UO_1878 (O_1878,N_15145,N_15953);
and UO_1879 (O_1879,N_15656,N_18093);
and UO_1880 (O_1880,N_17450,N_19083);
xor UO_1881 (O_1881,N_16657,N_18757);
nand UO_1882 (O_1882,N_17354,N_16655);
nand UO_1883 (O_1883,N_19045,N_16165);
xnor UO_1884 (O_1884,N_19587,N_18012);
or UO_1885 (O_1885,N_16870,N_19369);
and UO_1886 (O_1886,N_19207,N_17768);
or UO_1887 (O_1887,N_17174,N_17515);
xor UO_1888 (O_1888,N_19053,N_15297);
nand UO_1889 (O_1889,N_19728,N_15988);
or UO_1890 (O_1890,N_15216,N_16843);
nand UO_1891 (O_1891,N_19600,N_17232);
nor UO_1892 (O_1892,N_19055,N_17113);
xnor UO_1893 (O_1893,N_16267,N_16567);
nand UO_1894 (O_1894,N_16140,N_18117);
and UO_1895 (O_1895,N_19355,N_15884);
or UO_1896 (O_1896,N_16186,N_15059);
and UO_1897 (O_1897,N_18588,N_16363);
xnor UO_1898 (O_1898,N_19125,N_15010);
xor UO_1899 (O_1899,N_19821,N_17738);
nor UO_1900 (O_1900,N_19987,N_17572);
and UO_1901 (O_1901,N_19114,N_17926);
nor UO_1902 (O_1902,N_15067,N_19727);
nand UO_1903 (O_1903,N_15681,N_18772);
nand UO_1904 (O_1904,N_17141,N_17234);
nand UO_1905 (O_1905,N_16711,N_15524);
nor UO_1906 (O_1906,N_16925,N_15218);
or UO_1907 (O_1907,N_15890,N_19065);
or UO_1908 (O_1908,N_17901,N_17699);
nor UO_1909 (O_1909,N_17606,N_17643);
nand UO_1910 (O_1910,N_15225,N_17386);
or UO_1911 (O_1911,N_15710,N_16367);
nor UO_1912 (O_1912,N_18548,N_17612);
and UO_1913 (O_1913,N_15166,N_18575);
nand UO_1914 (O_1914,N_17972,N_18056);
nor UO_1915 (O_1915,N_17739,N_18123);
or UO_1916 (O_1916,N_15459,N_15593);
xnor UO_1917 (O_1917,N_15724,N_17123);
nor UO_1918 (O_1918,N_17930,N_17269);
nand UO_1919 (O_1919,N_17376,N_15780);
nor UO_1920 (O_1920,N_18226,N_19151);
nor UO_1921 (O_1921,N_16302,N_18467);
xor UO_1922 (O_1922,N_16330,N_18058);
nor UO_1923 (O_1923,N_15142,N_19119);
and UO_1924 (O_1924,N_17662,N_15125);
and UO_1925 (O_1925,N_19971,N_18022);
or UO_1926 (O_1926,N_17257,N_19148);
xor UO_1927 (O_1927,N_15555,N_15860);
nor UO_1928 (O_1928,N_19696,N_16012);
nand UO_1929 (O_1929,N_17960,N_17011);
nand UO_1930 (O_1930,N_16175,N_17978);
nand UO_1931 (O_1931,N_19441,N_18372);
nand UO_1932 (O_1932,N_15237,N_18219);
nor UO_1933 (O_1933,N_18778,N_19074);
nand UO_1934 (O_1934,N_19622,N_18612);
and UO_1935 (O_1935,N_18057,N_17676);
xnor UO_1936 (O_1936,N_15644,N_15799);
xnor UO_1937 (O_1937,N_19709,N_17468);
or UO_1938 (O_1938,N_18329,N_15940);
or UO_1939 (O_1939,N_18968,N_15944);
nand UO_1940 (O_1940,N_18213,N_19629);
xnor UO_1941 (O_1941,N_17534,N_19666);
and UO_1942 (O_1942,N_15610,N_16982);
or UO_1943 (O_1943,N_16429,N_18827);
or UO_1944 (O_1944,N_15574,N_19707);
nand UO_1945 (O_1945,N_17576,N_19486);
and UO_1946 (O_1946,N_18070,N_17994);
nand UO_1947 (O_1947,N_15810,N_17605);
and UO_1948 (O_1948,N_15098,N_17649);
xor UO_1949 (O_1949,N_16743,N_17704);
and UO_1950 (O_1950,N_18695,N_18858);
nand UO_1951 (O_1951,N_18914,N_17206);
nor UO_1952 (O_1952,N_19800,N_15652);
or UO_1953 (O_1953,N_15730,N_19417);
or UO_1954 (O_1954,N_15815,N_18622);
xor UO_1955 (O_1955,N_19184,N_17627);
nand UO_1956 (O_1956,N_19769,N_19964);
xor UO_1957 (O_1957,N_18455,N_18666);
and UO_1958 (O_1958,N_15061,N_18299);
or UO_1959 (O_1959,N_16260,N_16998);
xnor UO_1960 (O_1960,N_17876,N_15124);
nand UO_1961 (O_1961,N_17298,N_19092);
xnor UO_1962 (O_1962,N_15030,N_15683);
nor UO_1963 (O_1963,N_19234,N_15604);
xnor UO_1964 (O_1964,N_16483,N_15829);
nor UO_1965 (O_1965,N_15697,N_17272);
nor UO_1966 (O_1966,N_16714,N_19626);
or UO_1967 (O_1967,N_15397,N_17651);
xnor UO_1968 (O_1968,N_16733,N_19947);
and UO_1969 (O_1969,N_15069,N_16807);
or UO_1970 (O_1970,N_17494,N_15244);
nand UO_1971 (O_1971,N_18363,N_18807);
nand UO_1972 (O_1972,N_17705,N_18894);
nor UO_1973 (O_1973,N_17806,N_16020);
nand UO_1974 (O_1974,N_19396,N_17519);
nor UO_1975 (O_1975,N_18683,N_16934);
and UO_1976 (O_1976,N_19853,N_19010);
and UO_1977 (O_1977,N_15680,N_18902);
or UO_1978 (O_1978,N_15104,N_16041);
or UO_1979 (O_1979,N_17541,N_16649);
xor UO_1980 (O_1980,N_19116,N_16286);
xnor UO_1981 (O_1981,N_17579,N_17138);
xor UO_1982 (O_1982,N_16732,N_15668);
xor UO_1983 (O_1983,N_18397,N_18659);
or UO_1984 (O_1984,N_18725,N_18401);
xnor UO_1985 (O_1985,N_18458,N_19642);
xor UO_1986 (O_1986,N_16945,N_18667);
xnor UO_1987 (O_1987,N_19918,N_16098);
nor UO_1988 (O_1988,N_18739,N_17195);
or UO_1989 (O_1989,N_17957,N_16410);
nand UO_1990 (O_1990,N_16323,N_16751);
nor UO_1991 (O_1991,N_18529,N_15868);
xor UO_1992 (O_1992,N_15925,N_18107);
or UO_1993 (O_1993,N_16726,N_17157);
nand UO_1994 (O_1994,N_16395,N_18700);
nand UO_1995 (O_1995,N_19370,N_19997);
nor UO_1996 (O_1996,N_18449,N_17496);
or UO_1997 (O_1997,N_16933,N_18947);
and UO_1998 (O_1998,N_17525,N_18011);
or UO_1999 (O_1999,N_19084,N_18457);
or UO_2000 (O_2000,N_18280,N_16340);
and UO_2001 (O_2001,N_16239,N_19108);
nor UO_2002 (O_2002,N_18331,N_16648);
xor UO_2003 (O_2003,N_19566,N_17299);
xor UO_2004 (O_2004,N_16809,N_15530);
or UO_2005 (O_2005,N_18823,N_16825);
and UO_2006 (O_2006,N_17786,N_17577);
or UO_2007 (O_2007,N_18569,N_18648);
and UO_2008 (O_2008,N_17425,N_19160);
nor UO_2009 (O_2009,N_16278,N_15031);
xnor UO_2010 (O_2010,N_19615,N_16892);
xnor UO_2011 (O_2011,N_16411,N_19067);
nand UO_2012 (O_2012,N_17949,N_19961);
or UO_2013 (O_2013,N_15779,N_17416);
nand UO_2014 (O_2014,N_15705,N_19936);
nor UO_2015 (O_2015,N_18216,N_19836);
nand UO_2016 (O_2016,N_15447,N_17968);
nand UO_2017 (O_2017,N_15423,N_18808);
or UO_2018 (O_2018,N_17387,N_19780);
or UO_2019 (O_2019,N_19389,N_17473);
and UO_2020 (O_2020,N_18183,N_15745);
nor UO_2021 (O_2021,N_19656,N_15077);
nor UO_2022 (O_2022,N_17314,N_19660);
nand UO_2023 (O_2023,N_16800,N_17428);
nor UO_2024 (O_2024,N_15128,N_15448);
and UO_2025 (O_2025,N_16434,N_15733);
nor UO_2026 (O_2026,N_17681,N_17788);
xor UO_2027 (O_2027,N_18366,N_18343);
and UO_2028 (O_2028,N_18777,N_15416);
xnor UO_2029 (O_2029,N_17241,N_15699);
xor UO_2030 (O_2030,N_16174,N_16374);
nand UO_2031 (O_2031,N_17837,N_16906);
nor UO_2032 (O_2032,N_17688,N_17584);
nor UO_2033 (O_2033,N_16871,N_16631);
nand UO_2034 (O_2034,N_19603,N_16805);
nand UO_2035 (O_2035,N_16081,N_17549);
xnor UO_2036 (O_2036,N_15050,N_19744);
and UO_2037 (O_2037,N_15371,N_16848);
and UO_2038 (O_2038,N_19206,N_15984);
nand UO_2039 (O_2039,N_16919,N_15564);
xor UO_2040 (O_2040,N_18961,N_18429);
xnor UO_2041 (O_2041,N_17440,N_16076);
nor UO_2042 (O_2042,N_18774,N_16407);
nor UO_2043 (O_2043,N_15132,N_15855);
xor UO_2044 (O_2044,N_15139,N_18199);
or UO_2045 (O_2045,N_19781,N_15684);
or UO_2046 (O_2046,N_18788,N_17923);
xor UO_2047 (O_2047,N_17874,N_16972);
nand UO_2048 (O_2048,N_16706,N_16717);
nor UO_2049 (O_2049,N_18245,N_18387);
or UO_2050 (O_2050,N_17022,N_17540);
and UO_2051 (O_2051,N_15226,N_19230);
and UO_2052 (O_2052,N_15044,N_17223);
or UO_2053 (O_2053,N_18955,N_17526);
nand UO_2054 (O_2054,N_19003,N_15488);
nor UO_2055 (O_2055,N_17259,N_19784);
nand UO_2056 (O_2056,N_17414,N_18716);
xor UO_2057 (O_2057,N_17596,N_18433);
xnor UO_2058 (O_2058,N_16780,N_18654);
or UO_2059 (O_2059,N_16149,N_18887);
or UO_2060 (O_2060,N_16777,N_17209);
or UO_2061 (O_2061,N_16387,N_15248);
nand UO_2062 (O_2062,N_18461,N_19431);
nand UO_2063 (O_2063,N_16018,N_16798);
or UO_2064 (O_2064,N_16536,N_16762);
and UO_2065 (O_2065,N_17580,N_19659);
nor UO_2066 (O_2066,N_16053,N_16184);
xor UO_2067 (O_2067,N_19531,N_17563);
and UO_2068 (O_2068,N_17053,N_15272);
xor UO_2069 (O_2069,N_17319,N_18035);
nand UO_2070 (O_2070,N_15892,N_17246);
xor UO_2071 (O_2071,N_16981,N_19599);
or UO_2072 (O_2072,N_19347,N_16284);
nand UO_2073 (O_2073,N_16672,N_15325);
xnor UO_2074 (O_2074,N_19304,N_16759);
nor UO_2075 (O_2075,N_18336,N_16789);
and UO_2076 (O_2076,N_19440,N_16051);
nor UO_2077 (O_2077,N_17261,N_16788);
and UO_2078 (O_2078,N_15999,N_16214);
nor UO_2079 (O_2079,N_15912,N_17306);
xor UO_2080 (O_2080,N_17668,N_16768);
or UO_2081 (O_2081,N_16676,N_16259);
and UO_2082 (O_2082,N_18127,N_17656);
or UO_2083 (O_2083,N_17588,N_15671);
nor UO_2084 (O_2084,N_19721,N_18726);
xnor UO_2085 (O_2085,N_19912,N_16491);
xor UO_2086 (O_2086,N_17305,N_16772);
nand UO_2087 (O_2087,N_16827,N_19601);
nor UO_2088 (O_2088,N_16849,N_19695);
nor UO_2089 (O_2089,N_16031,N_17782);
or UO_2090 (O_2090,N_16796,N_16874);
nand UO_2091 (O_2091,N_15978,N_16795);
nor UO_2092 (O_2092,N_15094,N_16857);
xnor UO_2093 (O_2093,N_16257,N_17894);
or UO_2094 (O_2094,N_15964,N_18215);
nand UO_2095 (O_2095,N_15206,N_15376);
xnor UO_2096 (O_2096,N_16073,N_17762);
nor UO_2097 (O_2097,N_17059,N_16408);
and UO_2098 (O_2098,N_15770,N_18710);
or UO_2099 (O_2099,N_18946,N_18859);
nor UO_2100 (O_2100,N_15051,N_15107);
nor UO_2101 (O_2101,N_17081,N_16137);
nor UO_2102 (O_2102,N_17421,N_16608);
and UO_2103 (O_2103,N_18655,N_19028);
or UO_2104 (O_2104,N_18805,N_18371);
nor UO_2105 (O_2105,N_15588,N_19086);
xnor UO_2106 (O_2106,N_17293,N_18738);
nor UO_2107 (O_2107,N_17256,N_17817);
xor UO_2108 (O_2108,N_16244,N_15837);
nor UO_2109 (O_2109,N_15501,N_19202);
or UO_2110 (O_2110,N_17291,N_15666);
and UO_2111 (O_2111,N_19332,N_16472);
or UO_2112 (O_2112,N_19674,N_15012);
nand UO_2113 (O_2113,N_18289,N_16731);
nor UO_2114 (O_2114,N_19840,N_19087);
and UO_2115 (O_2115,N_17582,N_18988);
nand UO_2116 (O_2116,N_16980,N_19348);
or UO_2117 (O_2117,N_16696,N_15419);
or UO_2118 (O_2118,N_17439,N_19200);
nand UO_2119 (O_2119,N_15918,N_19030);
nor UO_2120 (O_2120,N_19255,N_18488);
xor UO_2121 (O_2121,N_16866,N_18292);
xor UO_2122 (O_2122,N_19834,N_19433);
nand UO_2123 (O_2123,N_15767,N_18691);
xnor UO_2124 (O_2124,N_17602,N_19358);
nand UO_2125 (O_2125,N_17009,N_18506);
xor UO_2126 (O_2126,N_19376,N_17130);
and UO_2127 (O_2127,N_15549,N_17285);
nand UO_2128 (O_2128,N_18260,N_17734);
and UO_2129 (O_2129,N_16764,N_19664);
nor UO_2130 (O_2130,N_18238,N_18355);
nand UO_2131 (O_2131,N_16251,N_19340);
or UO_2132 (O_2132,N_15463,N_17841);
and UO_2133 (O_2133,N_15645,N_18263);
and UO_2134 (O_2134,N_16043,N_19979);
xor UO_2135 (O_2135,N_18996,N_15028);
xnor UO_2136 (O_2136,N_15585,N_15033);
xnor UO_2137 (O_2137,N_17986,N_19375);
nor UO_2138 (O_2138,N_16368,N_19574);
nand UO_2139 (O_2139,N_15523,N_16553);
nor UO_2140 (O_2140,N_18384,N_15729);
xor UO_2141 (O_2141,N_17275,N_18493);
xor UO_2142 (O_2142,N_15221,N_18841);
nor UO_2143 (O_2143,N_18689,N_17173);
nor UO_2144 (O_2144,N_17120,N_18773);
or UO_2145 (O_2145,N_18969,N_19617);
xnor UO_2146 (O_2146,N_15233,N_16576);
nand UO_2147 (O_2147,N_16894,N_18196);
and UO_2148 (O_2148,N_15800,N_15115);
nand UO_2149 (O_2149,N_16049,N_16331);
or UO_2150 (O_2150,N_18835,N_17638);
nor UO_2151 (O_2151,N_15366,N_18388);
nand UO_2152 (O_2152,N_16596,N_18693);
and UO_2153 (O_2153,N_15802,N_15271);
and UO_2154 (O_2154,N_15243,N_19363);
or UO_2155 (O_2155,N_17309,N_15676);
nor UO_2156 (O_2156,N_16664,N_17284);
nor UO_2157 (O_2157,N_16059,N_18884);
nand UO_2158 (O_2158,N_15362,N_15578);
or UO_2159 (O_2159,N_15436,N_18494);
nand UO_2160 (O_2160,N_16335,N_18730);
or UO_2161 (O_2161,N_15279,N_15180);
and UO_2162 (O_2162,N_19618,N_16354);
nor UO_2163 (O_2163,N_19487,N_18170);
or UO_2164 (O_2164,N_16261,N_15698);
nand UO_2165 (O_2165,N_19102,N_19189);
nor UO_2166 (O_2166,N_19299,N_15969);
xnor UO_2167 (O_2167,N_19637,N_15552);
or UO_2168 (O_2168,N_16793,N_17601);
nor UO_2169 (O_2169,N_15198,N_15711);
xor UO_2170 (O_2170,N_15363,N_18050);
and UO_2171 (O_2171,N_19796,N_16557);
nor UO_2172 (O_2172,N_16616,N_17903);
nand UO_2173 (O_2173,N_15163,N_16242);
and UO_2174 (O_2174,N_15075,N_15968);
or UO_2175 (O_2175,N_17506,N_15439);
and UO_2176 (O_2176,N_18051,N_17199);
and UO_2177 (O_2177,N_19820,N_16675);
nor UO_2178 (O_2178,N_17001,N_18341);
and UO_2179 (O_2179,N_17950,N_18256);
xor UO_2180 (O_2180,N_17433,N_16506);
or UO_2181 (O_2181,N_16510,N_15627);
and UO_2182 (O_2182,N_19679,N_17925);
nand UO_2183 (O_2183,N_17535,N_16480);
nor UO_2184 (O_2184,N_19217,N_16446);
nand UO_2185 (O_2185,N_15886,N_19226);
nor UO_2186 (O_2186,N_15258,N_15127);
xor UO_2187 (O_2187,N_15491,N_19413);
nand UO_2188 (O_2188,N_18115,N_16662);
nand UO_2189 (O_2189,N_19111,N_15998);
nand UO_2190 (O_2190,N_19685,N_17550);
nand UO_2191 (O_2191,N_16626,N_19334);
xnor UO_2192 (O_2192,N_18360,N_15438);
nand UO_2193 (O_2193,N_15753,N_18160);
nand UO_2194 (O_2194,N_17948,N_15561);
or UO_2195 (O_2195,N_17732,N_16753);
xnor UO_2196 (O_2196,N_16577,N_16288);
and UO_2197 (O_2197,N_18316,N_16549);
nand UO_2198 (O_2198,N_17300,N_16856);
and UO_2199 (O_2199,N_19851,N_19503);
and UO_2200 (O_2200,N_15825,N_16503);
nand UO_2201 (O_2201,N_19070,N_15267);
xnor UO_2202 (O_2202,N_16252,N_19692);
nor UO_2203 (O_2203,N_18015,N_19794);
nand UO_2204 (O_2204,N_18965,N_15368);
and UO_2205 (O_2205,N_15630,N_18113);
nor UO_2206 (O_2206,N_15816,N_17538);
nand UO_2207 (O_2207,N_17288,N_18825);
and UO_2208 (O_2208,N_18839,N_16106);
nor UO_2209 (O_2209,N_18108,N_17235);
nand UO_2210 (O_2210,N_18468,N_18475);
xnor UO_2211 (O_2211,N_19212,N_16040);
xnor UO_2212 (O_2212,N_19476,N_15418);
xor UO_2213 (O_2213,N_19902,N_18323);
nor UO_2214 (O_2214,N_19122,N_17979);
nand UO_2215 (O_2215,N_15946,N_18444);
and UO_2216 (O_2216,N_16228,N_19825);
and UO_2217 (O_2217,N_19205,N_19275);
nand UO_2218 (O_2218,N_15016,N_18637);
xor UO_2219 (O_2219,N_18016,N_16730);
or UO_2220 (O_2220,N_17911,N_18190);
xor UO_2221 (O_2221,N_17721,N_17333);
nor UO_2222 (O_2222,N_17037,N_18589);
nor UO_2223 (O_2223,N_17850,N_15597);
nand UO_2224 (O_2224,N_15557,N_16520);
nand UO_2225 (O_2225,N_18989,N_17937);
nor UO_2226 (O_2226,N_16369,N_17652);
xnor UO_2227 (O_2227,N_19910,N_16114);
xnor UO_2228 (O_2228,N_18664,N_15405);
xor UO_2229 (O_2229,N_16379,N_16699);
nand UO_2230 (O_2230,N_15096,N_17819);
xnor UO_2231 (O_2231,N_18861,N_15026);
or UO_2232 (O_2232,N_15058,N_16196);
xor UO_2233 (O_2233,N_16072,N_17317);
nand UO_2234 (O_2234,N_19530,N_19444);
nor UO_2235 (O_2235,N_17124,N_15838);
or UO_2236 (O_2236,N_15807,N_18680);
or UO_2237 (O_2237,N_18801,N_15321);
nor UO_2238 (O_2238,N_17777,N_16970);
xor UO_2239 (O_2239,N_15760,N_16084);
or UO_2240 (O_2240,N_18537,N_19251);
or UO_2241 (O_2241,N_16584,N_15369);
nor UO_2242 (O_2242,N_19274,N_18662);
or UO_2243 (O_2243,N_15819,N_19188);
nand UO_2244 (O_2244,N_16000,N_15099);
xnor UO_2245 (O_2245,N_16088,N_15402);
nand UO_2246 (O_2246,N_16004,N_18244);
nor UO_2247 (O_2247,N_18472,N_19829);
nor UO_2248 (O_2248,N_19374,N_16725);
nand UO_2249 (O_2249,N_15064,N_17015);
nor UO_2250 (O_2250,N_19773,N_16074);
nand UO_2251 (O_2251,N_17378,N_17112);
nor UO_2252 (O_2252,N_16761,N_17373);
or UO_2253 (O_2253,N_16861,N_17243);
nor UO_2254 (O_2254,N_17395,N_15990);
or UO_2255 (O_2255,N_15854,N_17943);
and UO_2256 (O_2256,N_18078,N_18074);
or UO_2257 (O_2257,N_17008,N_16690);
or UO_2258 (O_2258,N_16092,N_18984);
nand UO_2259 (O_2259,N_15989,N_15048);
nor UO_2260 (O_2260,N_15851,N_19411);
xor UO_2261 (O_2261,N_19229,N_16555);
and UO_2262 (O_2262,N_18369,N_18820);
nor UO_2263 (O_2263,N_16105,N_15052);
nand UO_2264 (O_2264,N_15039,N_17181);
nand UO_2265 (O_2265,N_17324,N_19384);
nand UO_2266 (O_2266,N_16155,N_19812);
or UO_2267 (O_2267,N_19636,N_19549);
xnor UO_2268 (O_2268,N_16221,N_19485);
xor UO_2269 (O_2269,N_19999,N_17147);
and UO_2270 (O_2270,N_18668,N_18735);
nor UO_2271 (O_2271,N_18082,N_17711);
xnor UO_2272 (O_2272,N_17397,N_18043);
or UO_2273 (O_2273,N_15688,N_19880);
or UO_2274 (O_2274,N_18275,N_15894);
or UO_2275 (O_2275,N_17464,N_16840);
or UO_2276 (O_2276,N_18930,N_15514);
and UO_2277 (O_2277,N_17438,N_18044);
nor UO_2278 (O_2278,N_16054,N_16920);
nor UO_2279 (O_2279,N_19609,N_19774);
xor UO_2280 (O_2280,N_16820,N_18980);
nand UO_2281 (O_2281,N_15246,N_19515);
nand UO_2282 (O_2282,N_16226,N_15429);
and UO_2283 (O_2283,N_16458,N_19719);
or UO_2284 (O_2284,N_18748,N_19873);
nand UO_2285 (O_2285,N_15763,N_19814);
nand UO_2286 (O_2286,N_18243,N_16224);
nor UO_2287 (O_2287,N_19535,N_17566);
or UO_2288 (O_2288,N_19199,N_18136);
xor UO_2289 (O_2289,N_18162,N_15111);
or UO_2290 (O_2290,N_16698,N_17915);
or UO_2291 (O_2291,N_18978,N_16741);
xor UO_2292 (O_2292,N_19372,N_18201);
nand UO_2293 (O_2293,N_19146,N_17918);
and UO_2294 (O_2294,N_19568,N_17829);
or UO_2295 (O_2295,N_18349,N_16336);
nand UO_2296 (O_2296,N_15182,N_16036);
and UO_2297 (O_2297,N_16497,N_16956);
xnor UO_2298 (O_2298,N_17188,N_17090);
nand UO_2299 (O_2299,N_18229,N_16652);
nor UO_2300 (O_2300,N_15532,N_17273);
nor UO_2301 (O_2301,N_19584,N_15821);
and UO_2302 (O_2302,N_18950,N_17020);
and UO_2303 (O_2303,N_15070,N_17713);
or UO_2304 (O_2304,N_17684,N_16512);
nor UO_2305 (O_2305,N_15043,N_17687);
or UO_2306 (O_2306,N_18942,N_19949);
nand UO_2307 (O_2307,N_17104,N_15844);
or UO_2308 (O_2308,N_19631,N_15565);
or UO_2309 (O_2309,N_19041,N_17951);
nor UO_2310 (O_2310,N_19828,N_18209);
xnor UO_2311 (O_2311,N_18062,N_16579);
xnor UO_2312 (O_2312,N_16218,N_15665);
xor UO_2313 (O_2313,N_19178,N_18296);
or UO_2314 (O_2314,N_18701,N_19357);
xor UO_2315 (O_2315,N_19136,N_17313);
nand UO_2316 (O_2316,N_15913,N_15777);
and UO_2317 (O_2317,N_15513,N_18536);
or UO_2318 (O_2318,N_19281,N_19959);
nor UO_2319 (O_2319,N_16415,N_15204);
xor UO_2320 (O_2320,N_17998,N_15657);
or UO_2321 (O_2321,N_16507,N_17916);
or UO_2322 (O_2322,N_15736,N_18912);
nand UO_2323 (O_2323,N_18252,N_18552);
nand UO_2324 (O_2324,N_15531,N_17085);
nor UO_2325 (O_2325,N_17816,N_15891);
xor UO_2326 (O_2326,N_18320,N_19079);
or UO_2327 (O_2327,N_19139,N_16246);
nand UO_2328 (O_2328,N_19908,N_17226);
nand UO_2329 (O_2329,N_17030,N_18391);
and UO_2330 (O_2330,N_15406,N_16402);
nand UO_2331 (O_2331,N_15437,N_15824);
and UO_2332 (O_2332,N_19072,N_17603);
and UO_2333 (O_2333,N_15005,N_15381);
xnor UO_2334 (O_2334,N_17411,N_17431);
and UO_2335 (O_2335,N_19197,N_16482);
nor UO_2336 (O_2336,N_16757,N_17963);
and UO_2337 (O_2337,N_18132,N_16988);
nand UO_2338 (O_2338,N_15384,N_15540);
and UO_2339 (O_2339,N_19518,N_19091);
nor UO_2340 (O_2340,N_15372,N_19350);
nor UO_2341 (O_2341,N_18400,N_19516);
and UO_2342 (O_2342,N_19023,N_15411);
and UO_2343 (O_2343,N_18549,N_16630);
and UO_2344 (O_2344,N_18568,N_16974);
nor UO_2345 (O_2345,N_16538,N_18866);
and UO_2346 (O_2346,N_15551,N_18007);
or UO_2347 (O_2347,N_15356,N_16413);
or UO_2348 (O_2348,N_18891,N_18538);
xnor UO_2349 (O_2349,N_19085,N_18845);
and UO_2350 (O_2350,N_15895,N_15950);
xnor UO_2351 (O_2351,N_17511,N_15914);
and UO_2352 (O_2352,N_18800,N_19472);
or UO_2353 (O_2353,N_16130,N_15515);
nor UO_2354 (O_2354,N_17489,N_18085);
nor UO_2355 (O_2355,N_15963,N_19040);
or UO_2356 (O_2356,N_19974,N_16571);
and UO_2357 (O_2357,N_15967,N_19635);
and UO_2358 (O_2358,N_19730,N_19138);
xnor UO_2359 (O_2359,N_17368,N_19837);
nand UO_2360 (O_2360,N_17646,N_19710);
or UO_2361 (O_2361,N_19420,N_18099);
nor UO_2362 (O_2362,N_17405,N_16560);
or UO_2363 (O_2363,N_16611,N_17614);
nor UO_2364 (O_2364,N_15228,N_17510);
xnor UO_2365 (O_2365,N_18396,N_15828);
or UO_2366 (O_2366,N_15112,N_15379);
xnor UO_2367 (O_2367,N_19093,N_15509);
or UO_2368 (O_2368,N_18610,N_18098);
xnor UO_2369 (O_2369,N_18819,N_19868);
xnor UO_2370 (O_2370,N_17888,N_18223);
xor UO_2371 (O_2371,N_15068,N_15643);
nand UO_2372 (O_2372,N_15193,N_19501);
nor UO_2373 (O_2373,N_17924,N_18940);
or UO_2374 (O_2374,N_16841,N_16545);
nand UO_2375 (O_2375,N_17542,N_18023);
and UO_2376 (O_2376,N_17323,N_15808);
and UO_2377 (O_2377,N_18910,N_15517);
nor UO_2378 (O_2378,N_15756,N_15996);
nand UO_2379 (O_2379,N_16693,N_19948);
nand UO_2380 (O_2380,N_15105,N_18403);
xnor UO_2381 (O_2381,N_17650,N_17956);
xor UO_2382 (O_2382,N_19610,N_16164);
and UO_2383 (O_2383,N_18541,N_17853);
xnor UO_2384 (O_2384,N_15594,N_18286);
and UO_2385 (O_2385,N_15347,N_17080);
xnor UO_2386 (O_2386,N_16747,N_15300);
nor UO_2387 (O_2387,N_16642,N_15809);
and UO_2388 (O_2388,N_19550,N_18135);
nand UO_2389 (O_2389,N_15344,N_18405);
xor UO_2390 (O_2390,N_16684,N_19688);
nor UO_2391 (O_2391,N_17117,N_15670);
nand UO_2392 (O_2392,N_19283,N_19292);
nor UO_2393 (O_2393,N_17604,N_18149);
and UO_2394 (O_2394,N_16641,N_15169);
nor UO_2395 (O_2395,N_17176,N_19788);
and UO_2396 (O_2396,N_17399,N_19989);
or UO_2397 (O_2397,N_19914,N_19219);
and UO_2398 (O_2398,N_19127,N_17747);
nor UO_2399 (O_2399,N_17677,N_15718);
xnor UO_2400 (O_2400,N_18639,N_19760);
and UO_2401 (O_2401,N_16705,N_15938);
xor UO_2402 (O_2402,N_15231,N_18754);
nand UO_2403 (O_2403,N_18508,N_19459);
nor UO_2404 (O_2404,N_18310,N_19123);
and UO_2405 (O_2405,N_16575,N_17329);
or UO_2406 (O_2406,N_19869,N_17730);
or UO_2407 (O_2407,N_15256,N_19716);
nand UO_2408 (O_2408,N_16546,N_18806);
xor UO_2409 (O_2409,N_15529,N_15993);
and UO_2410 (O_2410,N_19388,N_17312);
nor UO_2411 (O_2411,N_18594,N_18386);
and UO_2412 (O_2412,N_16987,N_19458);
xnor UO_2413 (O_2413,N_16400,N_19534);
and UO_2414 (O_2414,N_15811,N_16152);
nor UO_2415 (O_2415,N_15674,N_18842);
xor UO_2416 (O_2416,N_15349,N_16477);
nor UO_2417 (O_2417,N_17058,N_16715);
or UO_2418 (O_2418,N_19891,N_19588);
and UO_2419 (O_2419,N_17835,N_19267);
nand UO_2420 (O_2420,N_17101,N_16961);
xnor UO_2421 (O_2421,N_15273,N_19270);
and UO_2422 (O_2422,N_18262,N_17353);
xnor UO_2423 (O_2423,N_18344,N_17801);
nand UO_2424 (O_2424,N_15024,N_19291);
nor UO_2425 (O_2425,N_18587,N_16007);
and UO_2426 (O_2426,N_15581,N_16913);
or UO_2427 (O_2427,N_16758,N_15380);
xor UO_2428 (O_2428,N_18141,N_17759);
nand UO_2429 (O_2429,N_16528,N_15685);
xnor UO_2430 (O_2430,N_18636,N_18703);
xor UO_2431 (O_2431,N_19307,N_15725);
nor UO_2432 (O_2432,N_17629,N_18913);
xor UO_2433 (O_2433,N_19954,N_19225);
xor UO_2434 (O_2434,N_16814,N_17751);
and UO_2435 (O_2435,N_15534,N_18846);
nand UO_2436 (O_2436,N_16465,N_18073);
or UO_2437 (O_2437,N_17774,N_16333);
and UO_2438 (O_2438,N_17218,N_16783);
and UO_2439 (O_2439,N_16325,N_17679);
or UO_2440 (O_2440,N_15793,N_18888);
or UO_2441 (O_2441,N_16349,N_18954);
or UO_2442 (O_2442,N_15611,N_19508);
nand UO_2443 (O_2443,N_16019,N_18509);
xnor UO_2444 (O_2444,N_16771,N_19424);
nor UO_2445 (O_2445,N_18609,N_15936);
or UO_2446 (O_2446,N_19494,N_19434);
xnor UO_2447 (O_2447,N_16774,N_19681);
xor UO_2448 (O_2448,N_17647,N_16205);
xnor UO_2449 (O_2449,N_16276,N_15841);
nand UO_2450 (O_2450,N_17632,N_15373);
nor UO_2451 (O_2451,N_15502,N_19112);
xor UO_2452 (O_2452,N_19533,N_19385);
nor UO_2453 (O_2453,N_19956,N_19863);
or UO_2454 (O_2454,N_15490,N_17394);
or UO_2455 (O_2455,N_15959,N_17745);
nor UO_2456 (O_2456,N_17467,N_16143);
and UO_2457 (O_2457,N_15353,N_18525);
and UO_2458 (O_2458,N_15230,N_16537);
xor UO_2459 (O_2459,N_19843,N_16534);
nor UO_2460 (O_2460,N_18474,N_17204);
and UO_2461 (O_2461,N_19538,N_15307);
nand UO_2462 (O_2462,N_18338,N_17490);
nand UO_2463 (O_2463,N_16281,N_16292);
and UO_2464 (O_2464,N_16551,N_17599);
nor UO_2465 (O_2465,N_17508,N_15087);
nor UO_2466 (O_2466,N_17787,N_15769);
nand UO_2467 (O_2467,N_19690,N_17146);
or UO_2468 (O_2468,N_16650,N_17737);
and UO_2469 (O_2469,N_17046,N_15178);
and UO_2470 (O_2470,N_17152,N_16583);
nor UO_2471 (O_2471,N_16223,N_18869);
nor UO_2472 (O_2472,N_19310,N_17670);
and UO_2473 (O_2473,N_16361,N_18550);
xnor UO_2474 (O_2474,N_19691,N_19351);
nor UO_2475 (O_2475,N_19697,N_19329);
or UO_2476 (O_2476,N_15595,N_16133);
xor UO_2477 (O_2477,N_17867,N_19141);
nand UO_2478 (O_2478,N_17422,N_17671);
and UO_2479 (O_2479,N_19418,N_18967);
nand UO_2480 (O_2480,N_18318,N_18966);
xnor UO_2481 (O_2481,N_18563,N_15958);
and UO_2482 (O_2482,N_18877,N_15149);
nand UO_2483 (O_2483,N_18644,N_18679);
and UO_2484 (O_2484,N_15797,N_15921);
and UO_2485 (O_2485,N_17452,N_19107);
or UO_2486 (O_2486,N_18809,N_19733);
xor UO_2487 (O_2487,N_19705,N_16204);
nor UO_2488 (O_2488,N_15037,N_16104);
and UO_2489 (O_2489,N_16449,N_17217);
or UO_2490 (O_2490,N_17977,N_19142);
and UO_2491 (O_2491,N_18551,N_17764);
and UO_2492 (O_2492,N_15247,N_18227);
or UO_2493 (O_2493,N_16170,N_19149);
nor UO_2494 (O_2494,N_18522,N_19905);
nand UO_2495 (O_2495,N_15887,N_18650);
nor UO_2496 (O_2496,N_15937,N_19953);
and UO_2497 (O_2497,N_16791,N_17458);
xor UO_2498 (O_2498,N_18681,N_15722);
nand UO_2499 (O_2499,N_15526,N_18870);
endmodule