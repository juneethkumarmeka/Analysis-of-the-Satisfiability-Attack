module basic_1000_10000_1500_10_levels_2xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_724,In_766);
nor U1 (N_1,In_24,In_32);
nor U2 (N_2,In_147,In_9);
nand U3 (N_3,In_607,In_291);
and U4 (N_4,In_519,In_102);
nand U5 (N_5,In_581,In_702);
or U6 (N_6,In_606,In_103);
nand U7 (N_7,In_719,In_962);
nand U8 (N_8,In_514,In_474);
nand U9 (N_9,In_359,In_559);
or U10 (N_10,In_735,In_859);
nor U11 (N_11,In_941,In_57);
and U12 (N_12,In_897,In_840);
nand U13 (N_13,In_882,In_881);
and U14 (N_14,In_139,In_178);
and U15 (N_15,In_876,In_444);
or U16 (N_16,In_931,In_682);
nor U17 (N_17,In_903,In_647);
nand U18 (N_18,In_642,In_200);
nand U19 (N_19,In_553,In_81);
and U20 (N_20,In_68,In_341);
or U21 (N_21,In_908,In_93);
or U22 (N_22,In_796,In_53);
and U23 (N_23,In_853,In_75);
and U24 (N_24,In_65,In_163);
and U25 (N_25,In_532,In_873);
or U26 (N_26,In_942,In_856);
nand U27 (N_27,In_621,In_170);
or U28 (N_28,In_401,In_36);
nor U29 (N_29,In_728,In_248);
nand U30 (N_30,In_723,In_874);
or U31 (N_31,In_323,In_535);
nand U32 (N_32,In_598,In_822);
or U33 (N_33,In_925,In_218);
nor U34 (N_34,In_370,In_386);
or U35 (N_35,In_83,In_107);
or U36 (N_36,In_928,In_453);
nand U37 (N_37,In_989,In_515);
and U38 (N_38,In_570,In_288);
nand U39 (N_39,In_590,In_596);
nor U40 (N_40,In_828,In_551);
xor U41 (N_41,In_141,In_660);
and U42 (N_42,In_466,In_354);
nand U43 (N_43,In_130,In_584);
nand U44 (N_44,In_297,In_933);
or U45 (N_45,In_233,In_87);
and U46 (N_46,In_605,In_373);
nor U47 (N_47,In_977,In_738);
and U48 (N_48,In_499,In_135);
nand U49 (N_49,In_754,In_312);
nand U50 (N_50,In_43,In_831);
nor U51 (N_51,In_184,In_531);
and U52 (N_52,In_516,In_74);
nand U53 (N_53,In_802,In_174);
nor U54 (N_54,In_430,In_571);
or U55 (N_55,In_648,In_990);
nand U56 (N_56,In_587,In_543);
and U57 (N_57,In_943,In_619);
nand U58 (N_58,In_827,In_661);
and U59 (N_59,In_191,In_149);
nor U60 (N_60,In_637,In_157);
and U61 (N_61,In_592,In_109);
or U62 (N_62,In_310,In_525);
nor U63 (N_63,In_402,In_106);
xnor U64 (N_64,In_975,In_123);
nand U65 (N_65,In_818,In_47);
nand U66 (N_66,In_755,In_971);
or U67 (N_67,In_387,In_437);
nor U68 (N_68,In_739,In_599);
or U69 (N_69,In_722,In_825);
nand U70 (N_70,In_131,In_995);
and U71 (N_71,In_238,In_90);
or U72 (N_72,In_650,In_557);
nand U73 (N_73,In_253,In_765);
nand U74 (N_74,In_226,In_936);
or U75 (N_75,In_336,In_481);
and U76 (N_76,In_55,In_451);
nand U77 (N_77,In_817,In_980);
nor U78 (N_78,In_440,In_717);
nor U79 (N_79,In_677,In_947);
or U80 (N_80,In_665,In_568);
or U81 (N_81,In_194,In_114);
nand U82 (N_82,In_573,In_711);
or U83 (N_83,In_527,In_270);
and U84 (N_84,In_835,In_364);
and U85 (N_85,In_449,In_643);
nor U86 (N_86,In_976,In_877);
and U87 (N_87,In_8,In_829);
nand U88 (N_88,In_888,In_916);
nand U89 (N_89,In_128,In_795);
nand U90 (N_90,In_731,In_871);
or U91 (N_91,In_476,In_506);
nor U92 (N_92,In_306,In_472);
nor U93 (N_93,In_763,In_22);
or U94 (N_94,In_917,In_545);
nand U95 (N_95,In_448,In_815);
and U96 (N_96,In_246,In_945);
nor U97 (N_97,In_264,In_800);
and U98 (N_98,In_646,In_582);
nand U99 (N_99,In_845,In_477);
nand U100 (N_100,In_999,In_424);
and U101 (N_101,In_222,In_14);
and U102 (N_102,In_392,In_372);
or U103 (N_103,In_169,In_992);
nand U104 (N_104,In_961,In_979);
or U105 (N_105,In_922,In_281);
and U106 (N_106,In_59,In_811);
nand U107 (N_107,In_578,In_816);
nand U108 (N_108,In_788,In_681);
nor U109 (N_109,In_358,In_921);
or U110 (N_110,In_688,In_764);
nor U111 (N_111,In_241,In_985);
nor U112 (N_112,In_741,In_207);
or U113 (N_113,In_549,In_991);
or U114 (N_114,In_342,In_113);
nor U115 (N_115,In_693,In_574);
nor U116 (N_116,In_61,In_389);
or U117 (N_117,In_772,In_957);
or U118 (N_118,In_664,In_313);
and U119 (N_119,In_21,In_691);
nand U120 (N_120,In_436,In_186);
and U121 (N_121,In_552,In_641);
nor U122 (N_122,In_199,In_683);
nand U123 (N_123,In_29,In_547);
or U124 (N_124,In_217,In_585);
and U125 (N_125,In_132,In_508);
and U126 (N_126,In_280,In_537);
or U127 (N_127,In_858,In_517);
or U128 (N_128,In_697,In_413);
nand U129 (N_129,In_467,In_620);
and U130 (N_130,In_875,In_397);
xor U131 (N_131,In_40,In_912);
or U132 (N_132,In_834,In_100);
and U133 (N_133,In_416,In_227);
and U134 (N_134,In_396,In_631);
or U135 (N_135,In_564,In_899);
or U136 (N_136,In_165,In_98);
nor U137 (N_137,In_27,In_981);
or U138 (N_138,In_744,In_484);
nor U139 (N_139,In_320,In_303);
and U140 (N_140,In_459,In_580);
nor U141 (N_141,In_890,In_761);
or U142 (N_142,In_409,In_880);
nand U143 (N_143,In_234,In_544);
nor U144 (N_144,In_949,In_346);
nand U145 (N_145,In_565,In_263);
and U146 (N_146,In_91,In_694);
nor U147 (N_147,In_208,In_318);
or U148 (N_148,In_232,In_460);
and U149 (N_149,In_632,In_381);
nor U150 (N_150,In_566,In_279);
or U151 (N_151,In_80,In_548);
nand U152 (N_152,In_707,In_569);
and U153 (N_153,In_775,In_630);
nor U154 (N_154,In_277,In_932);
nand U155 (N_155,In_363,In_299);
or U156 (N_156,In_973,In_910);
nand U157 (N_157,In_0,In_972);
nor U158 (N_158,In_144,In_645);
and U159 (N_159,In_356,In_804);
and U160 (N_160,In_628,In_797);
nor U161 (N_161,In_750,In_202);
or U162 (N_162,In_901,In_58);
and U163 (N_163,In_92,In_421);
nand U164 (N_164,In_623,In_798);
and U165 (N_165,In_117,In_555);
nor U166 (N_166,In_177,In_528);
or U167 (N_167,In_478,In_920);
and U168 (N_168,In_562,In_13);
nand U169 (N_169,In_950,In_287);
or U170 (N_170,In_210,In_806);
nor U171 (N_171,In_30,In_377);
or U172 (N_172,In_770,In_304);
and U173 (N_173,In_777,In_616);
and U174 (N_174,In_46,In_867);
and U175 (N_175,In_913,In_333);
or U176 (N_176,In_240,In_205);
and U177 (N_177,In_322,In_355);
and U178 (N_178,In_196,In_382);
and U179 (N_179,In_894,In_679);
nand U180 (N_180,In_725,In_586);
nor U181 (N_181,In_340,In_457);
or U182 (N_182,In_809,In_134);
or U183 (N_183,In_629,In_690);
or U184 (N_184,In_610,In_930);
nor U185 (N_185,In_733,In_583);
and U186 (N_186,In_640,In_31);
xor U187 (N_187,In_133,In_790);
nor U188 (N_188,In_345,In_667);
or U189 (N_189,In_635,In_309);
and U190 (N_190,In_511,In_969);
or U191 (N_191,In_706,In_471);
nor U192 (N_192,In_497,In_420);
and U193 (N_193,In_452,In_496);
or U194 (N_194,In_450,In_110);
nor U195 (N_195,In_563,In_332);
or U196 (N_196,In_161,In_151);
and U197 (N_197,In_203,In_572);
nand U198 (N_198,In_812,In_305);
xnor U199 (N_199,In_316,In_101);
and U200 (N_200,In_197,In_791);
and U201 (N_201,In_625,In_35);
nor U202 (N_202,In_42,In_813);
nor U203 (N_203,In_403,In_51);
nand U204 (N_204,In_771,In_849);
nor U205 (N_205,In_275,In_521);
and U206 (N_206,In_824,In_940);
or U207 (N_207,In_339,In_172);
nand U208 (N_208,In_366,In_231);
nand U209 (N_209,In_984,In_844);
nand U210 (N_210,In_236,In_575);
nand U211 (N_211,In_352,In_863);
nand U212 (N_212,In_896,In_162);
nand U213 (N_213,In_948,In_39);
nand U214 (N_214,In_404,In_745);
and U215 (N_215,In_311,In_864);
and U216 (N_216,In_252,In_823);
nand U217 (N_217,In_997,In_768);
xnor U218 (N_218,In_594,In_70);
nor U219 (N_219,In_793,In_893);
nor U220 (N_220,In_77,In_736);
nand U221 (N_221,In_814,In_257);
or U222 (N_222,In_78,In_400);
xor U223 (N_223,In_353,In_529);
nor U224 (N_224,In_307,In_490);
nand U225 (N_225,In_410,In_656);
and U226 (N_226,In_613,In_368);
nand U227 (N_227,In_126,In_747);
and U228 (N_228,In_657,In_730);
nand U229 (N_229,In_603,In_485);
or U230 (N_230,In_308,In_180);
nand U231 (N_231,In_50,In_699);
or U232 (N_232,In_314,In_369);
and U233 (N_233,In_965,In_455);
nor U234 (N_234,In_335,In_810);
nor U235 (N_235,In_668,In_622);
and U236 (N_236,In_250,In_636);
xnor U237 (N_237,In_425,In_964);
and U238 (N_238,In_887,In_638);
nand U239 (N_239,In_493,In_468);
nor U240 (N_240,In_282,In_495);
nor U241 (N_241,In_266,In_841);
and U242 (N_242,In_429,In_998);
and U243 (N_243,In_680,In_480);
xor U244 (N_244,In_380,In_504);
nand U245 (N_245,In_385,In_442);
and U246 (N_246,In_28,In_136);
nor U247 (N_247,In_255,In_685);
and U248 (N_248,In_97,In_225);
and U249 (N_249,In_249,In_301);
nor U250 (N_250,In_522,In_6);
nand U251 (N_251,In_538,In_546);
nor U252 (N_252,In_627,In_153);
and U253 (N_253,In_294,In_82);
nand U254 (N_254,In_715,In_787);
or U255 (N_255,In_179,In_300);
or U256 (N_256,In_60,In_261);
nor U257 (N_257,In_315,In_684);
or U258 (N_258,In_762,In_904);
or U259 (N_259,In_862,In_938);
and U260 (N_260,In_391,In_639);
nor U261 (N_261,In_915,In_351);
or U262 (N_262,In_918,In_461);
and U263 (N_263,In_748,In_749);
and U264 (N_264,In_978,In_321);
nand U265 (N_265,In_937,In_89);
nor U266 (N_266,In_362,In_379);
nor U267 (N_267,In_520,In_669);
and U268 (N_268,In_394,In_689);
nor U269 (N_269,In_434,In_869);
nand U270 (N_270,In_432,In_854);
nor U271 (N_271,In_489,In_406);
nor U272 (N_272,In_152,In_884);
and U273 (N_273,In_601,In_150);
or U274 (N_274,In_944,In_125);
nor U275 (N_275,In_967,In_924);
nand U276 (N_276,In_376,In_794);
nor U277 (N_277,In_122,In_2);
and U278 (N_278,In_456,In_883);
nor U279 (N_279,In_542,In_142);
nand U280 (N_280,In_419,In_491);
nor U281 (N_281,In_716,In_168);
or U282 (N_282,In_143,In_63);
nand U283 (N_283,In_338,In_435);
nor U284 (N_284,In_792,In_41);
nor U285 (N_285,In_758,In_588);
nand U286 (N_286,In_192,In_17);
xor U287 (N_287,In_709,In_742);
or U288 (N_288,In_591,In_367);
and U289 (N_289,In_734,In_659);
nor U290 (N_290,In_617,In_95);
or U291 (N_291,In_433,In_900);
nand U292 (N_292,In_502,In_720);
or U293 (N_293,In_868,In_25);
nor U294 (N_294,In_26,In_780);
and U295 (N_295,In_350,In_462);
and U296 (N_296,In_618,In_268);
and U297 (N_297,In_820,In_789);
nand U298 (N_298,In_33,In_889);
and U299 (N_299,In_272,In_64);
and U300 (N_300,In_954,In_360);
nand U301 (N_301,In_963,In_176);
nand U302 (N_302,In_258,In_411);
nor U303 (N_303,In_348,In_295);
and U304 (N_304,In_260,In_526);
or U305 (N_305,In_686,In_16);
or U306 (N_306,In_673,In_159);
nor U307 (N_307,In_454,In_79);
or U308 (N_308,In_45,In_510);
nand U309 (N_309,In_73,In_513);
nand U310 (N_310,In_838,In_129);
nor U311 (N_311,In_422,In_533);
and U312 (N_312,In_447,In_395);
nand U313 (N_313,In_327,In_146);
and U314 (N_314,In_776,In_700);
and U315 (N_315,In_34,In_914);
or U316 (N_316,In_124,In_76);
nand U317 (N_317,In_173,In_672);
xor U318 (N_318,In_383,In_498);
nand U319 (N_319,In_955,In_751);
nor U320 (N_320,In_185,In_952);
nand U321 (N_321,In_567,In_96);
and U322 (N_322,In_254,In_469);
nand U323 (N_323,In_198,In_783);
or U324 (N_324,In_221,In_614);
or U325 (N_325,In_778,In_774);
nor U326 (N_326,In_705,In_654);
nand U327 (N_327,In_104,In_228);
and U328 (N_328,In_66,In_166);
or U329 (N_329,In_674,In_273);
and U330 (N_330,In_675,In_120);
or U331 (N_331,In_302,In_757);
nand U332 (N_332,In_843,In_269);
nor U333 (N_333,In_852,In_953);
nor U334 (N_334,In_259,In_906);
or U335 (N_335,In_140,In_213);
or U336 (N_336,In_986,In_785);
and U337 (N_337,In_326,In_215);
and U338 (N_338,In_836,In_958);
nor U339 (N_339,In_767,In_577);
xor U340 (N_340,In_600,In_801);
nor U341 (N_341,In_204,In_127);
nor U342 (N_342,In_371,In_56);
or U343 (N_343,In_99,In_927);
or U344 (N_344,In_704,In_740);
nand U345 (N_345,In_116,In_446);
nor U346 (N_346,In_826,In_760);
nand U347 (N_347,In_651,In_84);
nand U348 (N_348,In_407,In_865);
nor U349 (N_349,In_408,In_317);
and U350 (N_350,In_885,In_540);
nand U351 (N_351,In_833,In_220);
or U352 (N_352,In_968,In_54);
nand U353 (N_353,In_443,In_224);
nor U354 (N_354,In_781,In_753);
nand U355 (N_355,In_155,In_1);
nand U356 (N_356,In_283,In_439);
nor U357 (N_357,In_219,In_799);
nor U358 (N_358,In_743,In_426);
xnor U359 (N_359,In_509,In_518);
nand U360 (N_360,In_939,In_848);
and U361 (N_361,In_145,In_415);
nor U362 (N_362,In_188,In_94);
and U363 (N_363,In_653,In_898);
nand U364 (N_364,In_597,In_866);
and U365 (N_365,In_708,In_417);
nor U366 (N_366,In_251,In_769);
or U367 (N_367,In_727,In_934);
or U368 (N_368,In_615,In_759);
nor U369 (N_369,In_530,In_698);
or U370 (N_370,In_678,In_445);
and U371 (N_371,In_69,In_154);
and U372 (N_372,In_703,In_119);
nand U373 (N_373,In_365,In_523);
nand U374 (N_374,In_554,In_167);
nor U375 (N_375,In_996,In_160);
xnor U376 (N_376,In_105,In_331);
nand U377 (N_377,In_602,In_644);
and U378 (N_378,In_983,In_713);
or U379 (N_379,In_649,In_441);
or U380 (N_380,In_658,In_819);
nor U381 (N_381,In_247,In_712);
or U382 (N_382,In_48,In_687);
nand U383 (N_383,In_483,In_206);
nor U384 (N_384,In_399,In_121);
nor U385 (N_385,In_88,In_286);
nor U386 (N_386,In_909,In_714);
or U387 (N_387,In_701,In_935);
and U388 (N_388,In_482,In_663);
nand U389 (N_389,In_216,In_847);
and U390 (N_390,In_427,In_595);
or U391 (N_391,In_746,In_37);
xor U392 (N_392,In_12,In_604);
nor U393 (N_393,In_463,In_465);
nand U394 (N_394,In_62,In_556);
nand U395 (N_395,In_431,In_337);
or U396 (N_396,In_851,In_821);
or U397 (N_397,In_756,In_494);
xor U398 (N_398,In_3,In_211);
and U399 (N_399,In_138,In_611);
or U400 (N_400,In_256,In_267);
nand U401 (N_401,In_112,In_52);
or U402 (N_402,In_589,In_324);
nor U403 (N_403,In_512,In_223);
xnor U404 (N_404,In_44,In_946);
or U405 (N_405,In_891,In_633);
or U406 (N_406,In_902,In_438);
and U407 (N_407,In_919,In_729);
or U408 (N_408,In_993,In_807);
or U409 (N_409,In_966,In_970);
and U410 (N_410,In_190,In_229);
and U411 (N_411,In_670,In_929);
and U412 (N_412,In_558,In_737);
or U413 (N_413,In_710,In_374);
or U414 (N_414,In_837,In_608);
xor U415 (N_415,In_108,In_18);
and U416 (N_416,In_846,In_860);
or U417 (N_417,In_343,In_458);
nand U418 (N_418,In_329,In_325);
or U419 (N_419,In_696,In_830);
and U420 (N_420,In_662,In_156);
or U421 (N_421,In_892,In_384);
nor U422 (N_422,In_561,In_982);
nor U423 (N_423,In_473,In_959);
or U424 (N_424,In_414,In_671);
and U425 (N_425,In_289,In_189);
or U426 (N_426,In_726,In_390);
or U427 (N_427,In_560,In_666);
nand U428 (N_428,In_655,In_803);
xnor U429 (N_429,In_137,In_576);
or U430 (N_430,In_7,In_19);
nand U431 (N_431,In_243,In_11);
nand U432 (N_432,In_361,In_895);
nor U433 (N_433,In_405,In_951);
xnor U434 (N_434,In_181,In_388);
or U435 (N_435,In_148,In_245);
or U436 (N_436,In_271,In_230);
nor U437 (N_437,In_956,In_634);
nor U438 (N_438,In_212,In_773);
nand U439 (N_439,In_244,In_870);
or U440 (N_440,In_330,In_49);
and U441 (N_441,In_464,In_923);
and U442 (N_442,In_872,In_183);
or U443 (N_443,In_534,In_265);
nand U444 (N_444,In_470,In_861);
or U445 (N_445,In_718,In_237);
and U446 (N_446,In_926,In_71);
nand U447 (N_447,In_20,In_784);
or U448 (N_448,In_974,In_732);
and U449 (N_449,In_721,In_182);
nand U450 (N_450,In_626,In_652);
nor U451 (N_451,In_839,In_23);
nor U452 (N_452,In_503,In_290);
and U453 (N_453,In_214,In_118);
xnor U454 (N_454,In_344,In_193);
and U455 (N_455,In_72,In_187);
or U456 (N_456,In_85,In_857);
or U457 (N_457,In_805,In_86);
and U458 (N_458,In_550,In_695);
nor U459 (N_459,In_479,In_832);
or U460 (N_460,In_692,In_487);
nor U461 (N_461,In_334,In_475);
nor U462 (N_462,In_988,In_782);
and U463 (N_463,In_239,In_209);
and U464 (N_464,In_878,In_398);
nor U465 (N_465,In_115,In_507);
and U466 (N_466,In_201,In_505);
or U467 (N_467,In_905,In_850);
and U468 (N_468,In_67,In_158);
or U469 (N_469,In_676,In_298);
nor U470 (N_470,In_195,In_319);
and U471 (N_471,In_486,In_274);
or U472 (N_472,In_15,In_808);
nor U473 (N_473,In_752,In_579);
and U474 (N_474,In_262,In_879);
nand U475 (N_475,In_612,In_349);
nor U476 (N_476,In_357,In_378);
xnor U477 (N_477,In_296,In_284);
and U478 (N_478,In_855,In_987);
and U479 (N_479,In_492,In_500);
nand U480 (N_480,In_292,In_541);
and U481 (N_481,In_4,In_293);
or U482 (N_482,In_412,In_960);
or U483 (N_483,In_886,In_418);
or U484 (N_484,In_10,In_393);
and U485 (N_485,In_428,In_842);
nor U486 (N_486,In_536,In_423);
nor U487 (N_487,In_276,In_609);
xor U488 (N_488,In_164,In_375);
nand U489 (N_489,In_994,In_242);
nand U490 (N_490,In_278,In_779);
xor U491 (N_491,In_501,In_911);
nand U492 (N_492,In_539,In_285);
and U493 (N_493,In_235,In_38);
or U494 (N_494,In_328,In_171);
xnor U495 (N_495,In_5,In_111);
nand U496 (N_496,In_488,In_175);
and U497 (N_497,In_347,In_624);
nor U498 (N_498,In_524,In_907);
and U499 (N_499,In_593,In_786);
xnor U500 (N_500,In_926,In_218);
nand U501 (N_501,In_337,In_382);
or U502 (N_502,In_163,In_819);
nand U503 (N_503,In_141,In_958);
nor U504 (N_504,In_294,In_609);
nand U505 (N_505,In_984,In_57);
nor U506 (N_506,In_738,In_191);
nand U507 (N_507,In_701,In_257);
nor U508 (N_508,In_728,In_24);
and U509 (N_509,In_119,In_679);
nand U510 (N_510,In_158,In_256);
nand U511 (N_511,In_593,In_379);
and U512 (N_512,In_769,In_46);
and U513 (N_513,In_150,In_596);
nor U514 (N_514,In_137,In_715);
nand U515 (N_515,In_869,In_580);
and U516 (N_516,In_214,In_59);
nand U517 (N_517,In_624,In_43);
and U518 (N_518,In_91,In_388);
and U519 (N_519,In_585,In_690);
nand U520 (N_520,In_569,In_71);
or U521 (N_521,In_35,In_615);
nand U522 (N_522,In_581,In_513);
nand U523 (N_523,In_788,In_219);
nor U524 (N_524,In_227,In_6);
nand U525 (N_525,In_785,In_564);
nand U526 (N_526,In_381,In_819);
or U527 (N_527,In_284,In_495);
nand U528 (N_528,In_829,In_337);
nand U529 (N_529,In_291,In_341);
nor U530 (N_530,In_348,In_853);
nor U531 (N_531,In_227,In_464);
nor U532 (N_532,In_26,In_339);
or U533 (N_533,In_473,In_845);
nand U534 (N_534,In_234,In_872);
nand U535 (N_535,In_703,In_694);
or U536 (N_536,In_2,In_98);
nand U537 (N_537,In_99,In_889);
and U538 (N_538,In_415,In_668);
nor U539 (N_539,In_952,In_145);
and U540 (N_540,In_896,In_769);
nand U541 (N_541,In_938,In_703);
nand U542 (N_542,In_915,In_173);
or U543 (N_543,In_125,In_804);
nand U544 (N_544,In_989,In_206);
xor U545 (N_545,In_496,In_917);
and U546 (N_546,In_550,In_982);
nand U547 (N_547,In_364,In_578);
or U548 (N_548,In_743,In_691);
and U549 (N_549,In_13,In_325);
and U550 (N_550,In_785,In_379);
and U551 (N_551,In_149,In_247);
xor U552 (N_552,In_916,In_573);
nor U553 (N_553,In_575,In_295);
nor U554 (N_554,In_511,In_623);
nand U555 (N_555,In_68,In_51);
xnor U556 (N_556,In_47,In_243);
nand U557 (N_557,In_393,In_975);
or U558 (N_558,In_377,In_346);
or U559 (N_559,In_707,In_127);
nor U560 (N_560,In_127,In_854);
and U561 (N_561,In_583,In_92);
nor U562 (N_562,In_481,In_665);
xor U563 (N_563,In_883,In_514);
or U564 (N_564,In_586,In_109);
nor U565 (N_565,In_884,In_259);
nand U566 (N_566,In_518,In_432);
and U567 (N_567,In_51,In_83);
nor U568 (N_568,In_368,In_754);
nand U569 (N_569,In_740,In_181);
nor U570 (N_570,In_375,In_48);
nor U571 (N_571,In_774,In_347);
xor U572 (N_572,In_466,In_230);
or U573 (N_573,In_232,In_696);
or U574 (N_574,In_319,In_484);
nand U575 (N_575,In_95,In_247);
nand U576 (N_576,In_507,In_391);
nor U577 (N_577,In_469,In_703);
nand U578 (N_578,In_255,In_41);
nor U579 (N_579,In_973,In_721);
or U580 (N_580,In_546,In_572);
and U581 (N_581,In_780,In_114);
or U582 (N_582,In_752,In_394);
and U583 (N_583,In_43,In_81);
nand U584 (N_584,In_483,In_767);
and U585 (N_585,In_925,In_261);
nand U586 (N_586,In_181,In_96);
or U587 (N_587,In_656,In_244);
and U588 (N_588,In_292,In_190);
or U589 (N_589,In_703,In_125);
nor U590 (N_590,In_769,In_172);
nor U591 (N_591,In_667,In_477);
or U592 (N_592,In_212,In_460);
xor U593 (N_593,In_800,In_229);
nor U594 (N_594,In_322,In_255);
and U595 (N_595,In_583,In_359);
nand U596 (N_596,In_957,In_856);
and U597 (N_597,In_150,In_764);
nor U598 (N_598,In_384,In_542);
or U599 (N_599,In_169,In_320);
nor U600 (N_600,In_232,In_298);
or U601 (N_601,In_318,In_749);
or U602 (N_602,In_741,In_595);
nor U603 (N_603,In_174,In_250);
nand U604 (N_604,In_877,In_676);
nor U605 (N_605,In_951,In_103);
nor U606 (N_606,In_1,In_397);
nand U607 (N_607,In_615,In_527);
or U608 (N_608,In_111,In_303);
or U609 (N_609,In_177,In_805);
nand U610 (N_610,In_983,In_726);
nand U611 (N_611,In_643,In_175);
or U612 (N_612,In_634,In_123);
and U613 (N_613,In_288,In_576);
nand U614 (N_614,In_636,In_940);
nor U615 (N_615,In_684,In_740);
and U616 (N_616,In_53,In_3);
nor U617 (N_617,In_313,In_615);
nor U618 (N_618,In_447,In_985);
or U619 (N_619,In_741,In_483);
or U620 (N_620,In_643,In_239);
nor U621 (N_621,In_714,In_141);
and U622 (N_622,In_892,In_24);
xor U623 (N_623,In_944,In_386);
nor U624 (N_624,In_583,In_308);
nor U625 (N_625,In_184,In_37);
nand U626 (N_626,In_333,In_685);
nand U627 (N_627,In_893,In_100);
nand U628 (N_628,In_295,In_320);
and U629 (N_629,In_581,In_754);
nand U630 (N_630,In_978,In_128);
or U631 (N_631,In_598,In_199);
or U632 (N_632,In_320,In_754);
and U633 (N_633,In_245,In_817);
and U634 (N_634,In_955,In_464);
nor U635 (N_635,In_628,In_696);
nor U636 (N_636,In_692,In_299);
or U637 (N_637,In_343,In_418);
or U638 (N_638,In_545,In_13);
and U639 (N_639,In_256,In_203);
or U640 (N_640,In_69,In_314);
nand U641 (N_641,In_167,In_148);
nor U642 (N_642,In_372,In_203);
nor U643 (N_643,In_643,In_637);
nand U644 (N_644,In_218,In_378);
and U645 (N_645,In_334,In_467);
and U646 (N_646,In_803,In_664);
nor U647 (N_647,In_930,In_116);
or U648 (N_648,In_692,In_130);
and U649 (N_649,In_388,In_39);
nand U650 (N_650,In_169,In_296);
or U651 (N_651,In_286,In_989);
and U652 (N_652,In_104,In_840);
or U653 (N_653,In_324,In_160);
nor U654 (N_654,In_194,In_197);
nor U655 (N_655,In_507,In_506);
xnor U656 (N_656,In_676,In_776);
or U657 (N_657,In_510,In_266);
and U658 (N_658,In_627,In_115);
nand U659 (N_659,In_528,In_98);
and U660 (N_660,In_739,In_888);
nand U661 (N_661,In_108,In_811);
nand U662 (N_662,In_460,In_686);
xor U663 (N_663,In_719,In_302);
and U664 (N_664,In_331,In_663);
and U665 (N_665,In_418,In_92);
nor U666 (N_666,In_47,In_950);
nand U667 (N_667,In_816,In_976);
and U668 (N_668,In_220,In_776);
or U669 (N_669,In_115,In_14);
or U670 (N_670,In_233,In_890);
nand U671 (N_671,In_943,In_158);
nor U672 (N_672,In_285,In_284);
or U673 (N_673,In_3,In_134);
nor U674 (N_674,In_723,In_638);
nand U675 (N_675,In_786,In_611);
nand U676 (N_676,In_962,In_738);
or U677 (N_677,In_151,In_595);
or U678 (N_678,In_236,In_290);
or U679 (N_679,In_326,In_300);
or U680 (N_680,In_930,In_682);
nand U681 (N_681,In_131,In_215);
and U682 (N_682,In_371,In_880);
and U683 (N_683,In_597,In_981);
and U684 (N_684,In_11,In_503);
or U685 (N_685,In_336,In_496);
nand U686 (N_686,In_57,In_196);
nand U687 (N_687,In_541,In_295);
nor U688 (N_688,In_609,In_519);
and U689 (N_689,In_749,In_726);
and U690 (N_690,In_509,In_697);
nor U691 (N_691,In_136,In_722);
nor U692 (N_692,In_3,In_381);
nor U693 (N_693,In_650,In_896);
xnor U694 (N_694,In_438,In_155);
nor U695 (N_695,In_361,In_258);
or U696 (N_696,In_722,In_443);
nand U697 (N_697,In_871,In_759);
and U698 (N_698,In_406,In_279);
nand U699 (N_699,In_316,In_949);
or U700 (N_700,In_565,In_12);
nor U701 (N_701,In_18,In_144);
nand U702 (N_702,In_653,In_940);
or U703 (N_703,In_821,In_34);
xor U704 (N_704,In_187,In_516);
and U705 (N_705,In_126,In_16);
or U706 (N_706,In_771,In_53);
nor U707 (N_707,In_123,In_457);
nor U708 (N_708,In_958,In_672);
nor U709 (N_709,In_785,In_52);
and U710 (N_710,In_513,In_848);
or U711 (N_711,In_446,In_903);
nor U712 (N_712,In_58,In_549);
or U713 (N_713,In_914,In_338);
nand U714 (N_714,In_515,In_413);
nand U715 (N_715,In_609,In_963);
nand U716 (N_716,In_979,In_521);
xnor U717 (N_717,In_301,In_834);
nor U718 (N_718,In_110,In_87);
nor U719 (N_719,In_889,In_288);
or U720 (N_720,In_634,In_959);
nand U721 (N_721,In_494,In_931);
nand U722 (N_722,In_25,In_156);
and U723 (N_723,In_939,In_37);
nand U724 (N_724,In_407,In_680);
and U725 (N_725,In_102,In_945);
or U726 (N_726,In_878,In_942);
nor U727 (N_727,In_209,In_448);
or U728 (N_728,In_374,In_798);
and U729 (N_729,In_182,In_369);
and U730 (N_730,In_344,In_543);
and U731 (N_731,In_133,In_610);
nand U732 (N_732,In_127,In_400);
nand U733 (N_733,In_665,In_23);
nor U734 (N_734,In_564,In_415);
nand U735 (N_735,In_833,In_232);
xnor U736 (N_736,In_820,In_555);
or U737 (N_737,In_699,In_192);
nor U738 (N_738,In_439,In_424);
nor U739 (N_739,In_992,In_329);
nor U740 (N_740,In_757,In_826);
nor U741 (N_741,In_443,In_277);
or U742 (N_742,In_665,In_748);
and U743 (N_743,In_20,In_341);
and U744 (N_744,In_752,In_348);
nor U745 (N_745,In_73,In_739);
and U746 (N_746,In_767,In_447);
or U747 (N_747,In_746,In_241);
nand U748 (N_748,In_887,In_218);
xor U749 (N_749,In_754,In_456);
nor U750 (N_750,In_799,In_355);
nor U751 (N_751,In_571,In_833);
or U752 (N_752,In_589,In_557);
nor U753 (N_753,In_473,In_789);
or U754 (N_754,In_992,In_716);
xor U755 (N_755,In_203,In_873);
and U756 (N_756,In_57,In_556);
nand U757 (N_757,In_530,In_608);
nor U758 (N_758,In_541,In_213);
xor U759 (N_759,In_942,In_610);
nor U760 (N_760,In_534,In_752);
nor U761 (N_761,In_468,In_276);
nor U762 (N_762,In_542,In_646);
and U763 (N_763,In_472,In_585);
and U764 (N_764,In_761,In_914);
and U765 (N_765,In_437,In_311);
nor U766 (N_766,In_441,In_558);
nor U767 (N_767,In_999,In_634);
nand U768 (N_768,In_498,In_116);
and U769 (N_769,In_478,In_35);
nand U770 (N_770,In_545,In_346);
or U771 (N_771,In_53,In_435);
xnor U772 (N_772,In_409,In_652);
nand U773 (N_773,In_214,In_447);
nand U774 (N_774,In_9,In_907);
and U775 (N_775,In_18,In_691);
or U776 (N_776,In_353,In_850);
or U777 (N_777,In_118,In_986);
and U778 (N_778,In_194,In_176);
or U779 (N_779,In_700,In_540);
nor U780 (N_780,In_638,In_922);
and U781 (N_781,In_635,In_746);
and U782 (N_782,In_67,In_122);
nor U783 (N_783,In_725,In_201);
or U784 (N_784,In_117,In_201);
xor U785 (N_785,In_464,In_853);
xor U786 (N_786,In_644,In_333);
or U787 (N_787,In_249,In_78);
and U788 (N_788,In_21,In_372);
nor U789 (N_789,In_810,In_779);
and U790 (N_790,In_485,In_834);
and U791 (N_791,In_377,In_974);
nor U792 (N_792,In_789,In_905);
nor U793 (N_793,In_238,In_228);
nand U794 (N_794,In_92,In_325);
nor U795 (N_795,In_608,In_20);
or U796 (N_796,In_706,In_379);
or U797 (N_797,In_125,In_988);
nand U798 (N_798,In_439,In_890);
nand U799 (N_799,In_141,In_464);
and U800 (N_800,In_32,In_289);
nor U801 (N_801,In_856,In_869);
nor U802 (N_802,In_518,In_441);
nor U803 (N_803,In_631,In_66);
and U804 (N_804,In_511,In_95);
and U805 (N_805,In_865,In_836);
or U806 (N_806,In_328,In_872);
or U807 (N_807,In_699,In_695);
nand U808 (N_808,In_714,In_990);
nor U809 (N_809,In_736,In_730);
nand U810 (N_810,In_518,In_256);
or U811 (N_811,In_459,In_871);
nor U812 (N_812,In_293,In_783);
nand U813 (N_813,In_939,In_879);
or U814 (N_814,In_694,In_934);
nand U815 (N_815,In_141,In_337);
nor U816 (N_816,In_568,In_564);
nand U817 (N_817,In_578,In_236);
and U818 (N_818,In_479,In_127);
nor U819 (N_819,In_825,In_339);
nor U820 (N_820,In_385,In_576);
or U821 (N_821,In_261,In_200);
and U822 (N_822,In_396,In_443);
or U823 (N_823,In_203,In_709);
nand U824 (N_824,In_574,In_59);
and U825 (N_825,In_273,In_372);
or U826 (N_826,In_320,In_956);
nand U827 (N_827,In_189,In_716);
or U828 (N_828,In_547,In_445);
or U829 (N_829,In_360,In_685);
and U830 (N_830,In_315,In_311);
nor U831 (N_831,In_678,In_467);
nand U832 (N_832,In_428,In_876);
nand U833 (N_833,In_914,In_619);
nor U834 (N_834,In_256,In_989);
nor U835 (N_835,In_825,In_980);
or U836 (N_836,In_890,In_108);
nor U837 (N_837,In_986,In_301);
or U838 (N_838,In_920,In_116);
or U839 (N_839,In_147,In_349);
or U840 (N_840,In_862,In_581);
and U841 (N_841,In_300,In_451);
nor U842 (N_842,In_697,In_695);
or U843 (N_843,In_333,In_199);
and U844 (N_844,In_726,In_936);
or U845 (N_845,In_675,In_547);
or U846 (N_846,In_674,In_461);
nor U847 (N_847,In_325,In_913);
and U848 (N_848,In_316,In_93);
nor U849 (N_849,In_467,In_995);
nand U850 (N_850,In_247,In_832);
and U851 (N_851,In_791,In_720);
nand U852 (N_852,In_721,In_986);
nand U853 (N_853,In_783,In_268);
or U854 (N_854,In_734,In_911);
or U855 (N_855,In_450,In_311);
nand U856 (N_856,In_191,In_812);
nand U857 (N_857,In_75,In_674);
nand U858 (N_858,In_188,In_825);
nor U859 (N_859,In_799,In_447);
nand U860 (N_860,In_923,In_21);
nand U861 (N_861,In_866,In_932);
xor U862 (N_862,In_459,In_61);
nor U863 (N_863,In_80,In_118);
nor U864 (N_864,In_437,In_801);
nand U865 (N_865,In_3,In_182);
nand U866 (N_866,In_451,In_345);
or U867 (N_867,In_330,In_758);
or U868 (N_868,In_787,In_632);
or U869 (N_869,In_49,In_631);
nor U870 (N_870,In_95,In_123);
nand U871 (N_871,In_581,In_204);
or U872 (N_872,In_322,In_68);
or U873 (N_873,In_596,In_251);
nand U874 (N_874,In_337,In_822);
nand U875 (N_875,In_723,In_331);
nor U876 (N_876,In_246,In_705);
nor U877 (N_877,In_99,In_455);
nand U878 (N_878,In_279,In_983);
or U879 (N_879,In_810,In_872);
or U880 (N_880,In_384,In_226);
and U881 (N_881,In_115,In_488);
or U882 (N_882,In_524,In_49);
or U883 (N_883,In_477,In_305);
nor U884 (N_884,In_400,In_174);
nor U885 (N_885,In_71,In_793);
nor U886 (N_886,In_469,In_24);
or U887 (N_887,In_905,In_976);
nand U888 (N_888,In_9,In_75);
and U889 (N_889,In_284,In_789);
or U890 (N_890,In_875,In_7);
nor U891 (N_891,In_728,In_584);
or U892 (N_892,In_77,In_637);
or U893 (N_893,In_301,In_661);
nor U894 (N_894,In_271,In_163);
nand U895 (N_895,In_238,In_192);
and U896 (N_896,In_846,In_340);
nor U897 (N_897,In_304,In_209);
or U898 (N_898,In_981,In_543);
xnor U899 (N_899,In_928,In_253);
nand U900 (N_900,In_31,In_902);
or U901 (N_901,In_640,In_432);
xnor U902 (N_902,In_177,In_452);
or U903 (N_903,In_205,In_632);
or U904 (N_904,In_643,In_972);
nor U905 (N_905,In_324,In_577);
xor U906 (N_906,In_972,In_935);
and U907 (N_907,In_467,In_60);
xnor U908 (N_908,In_972,In_546);
and U909 (N_909,In_170,In_570);
nor U910 (N_910,In_662,In_500);
nand U911 (N_911,In_621,In_220);
or U912 (N_912,In_493,In_145);
or U913 (N_913,In_914,In_48);
and U914 (N_914,In_45,In_934);
or U915 (N_915,In_194,In_91);
and U916 (N_916,In_459,In_218);
and U917 (N_917,In_834,In_183);
or U918 (N_918,In_792,In_719);
and U919 (N_919,In_692,In_325);
and U920 (N_920,In_577,In_977);
nor U921 (N_921,In_501,In_60);
and U922 (N_922,In_769,In_41);
nor U923 (N_923,In_420,In_802);
and U924 (N_924,In_182,In_664);
and U925 (N_925,In_101,In_338);
or U926 (N_926,In_892,In_755);
and U927 (N_927,In_430,In_541);
and U928 (N_928,In_999,In_682);
nand U929 (N_929,In_910,In_16);
nand U930 (N_930,In_510,In_770);
nor U931 (N_931,In_924,In_33);
or U932 (N_932,In_925,In_377);
nand U933 (N_933,In_76,In_472);
and U934 (N_934,In_68,In_237);
nand U935 (N_935,In_109,In_916);
or U936 (N_936,In_790,In_631);
and U937 (N_937,In_847,In_358);
nand U938 (N_938,In_437,In_303);
nand U939 (N_939,In_275,In_297);
or U940 (N_940,In_916,In_683);
or U941 (N_941,In_597,In_200);
or U942 (N_942,In_393,In_994);
nor U943 (N_943,In_449,In_256);
nand U944 (N_944,In_793,In_54);
and U945 (N_945,In_250,In_208);
nor U946 (N_946,In_109,In_23);
nand U947 (N_947,In_762,In_464);
and U948 (N_948,In_343,In_260);
or U949 (N_949,In_953,In_970);
and U950 (N_950,In_64,In_834);
and U951 (N_951,In_218,In_157);
or U952 (N_952,In_163,In_155);
or U953 (N_953,In_287,In_316);
nor U954 (N_954,In_988,In_969);
nor U955 (N_955,In_749,In_918);
and U956 (N_956,In_406,In_725);
or U957 (N_957,In_702,In_759);
and U958 (N_958,In_42,In_52);
or U959 (N_959,In_979,In_806);
nand U960 (N_960,In_857,In_388);
nand U961 (N_961,In_595,In_39);
and U962 (N_962,In_424,In_468);
and U963 (N_963,In_912,In_586);
or U964 (N_964,In_577,In_973);
or U965 (N_965,In_195,In_346);
and U966 (N_966,In_144,In_275);
and U967 (N_967,In_786,In_671);
nor U968 (N_968,In_997,In_430);
or U969 (N_969,In_13,In_90);
or U970 (N_970,In_736,In_121);
nor U971 (N_971,In_451,In_369);
nand U972 (N_972,In_588,In_829);
and U973 (N_973,In_810,In_276);
nand U974 (N_974,In_802,In_226);
or U975 (N_975,In_634,In_183);
nand U976 (N_976,In_398,In_544);
nor U977 (N_977,In_513,In_266);
or U978 (N_978,In_101,In_858);
or U979 (N_979,In_204,In_234);
nand U980 (N_980,In_424,In_125);
nand U981 (N_981,In_710,In_741);
and U982 (N_982,In_441,In_43);
nand U983 (N_983,In_532,In_417);
and U984 (N_984,In_95,In_500);
nor U985 (N_985,In_314,In_119);
nor U986 (N_986,In_950,In_876);
and U987 (N_987,In_55,In_6);
and U988 (N_988,In_165,In_791);
nor U989 (N_989,In_307,In_605);
and U990 (N_990,In_943,In_183);
nand U991 (N_991,In_249,In_769);
nand U992 (N_992,In_694,In_763);
nor U993 (N_993,In_648,In_55);
nand U994 (N_994,In_45,In_355);
nand U995 (N_995,In_806,In_202);
nor U996 (N_996,In_6,In_713);
nand U997 (N_997,In_768,In_268);
nand U998 (N_998,In_709,In_137);
or U999 (N_999,In_866,In_236);
nor U1000 (N_1000,N_848,N_513);
nor U1001 (N_1001,N_244,N_90);
nand U1002 (N_1002,N_84,N_169);
nor U1003 (N_1003,N_544,N_316);
and U1004 (N_1004,N_844,N_407);
nor U1005 (N_1005,N_473,N_594);
nand U1006 (N_1006,N_215,N_734);
nand U1007 (N_1007,N_797,N_649);
and U1008 (N_1008,N_871,N_166);
and U1009 (N_1009,N_918,N_961);
nor U1010 (N_1010,N_261,N_647);
and U1011 (N_1011,N_6,N_706);
and U1012 (N_1012,N_672,N_278);
or U1013 (N_1013,N_348,N_122);
nand U1014 (N_1014,N_980,N_144);
or U1015 (N_1015,N_895,N_605);
nand U1016 (N_1016,N_521,N_638);
and U1017 (N_1017,N_220,N_661);
or U1018 (N_1018,N_861,N_164);
nor U1019 (N_1019,N_623,N_905);
and U1020 (N_1020,N_387,N_602);
nand U1021 (N_1021,N_221,N_385);
or U1022 (N_1022,N_753,N_63);
and U1023 (N_1023,N_763,N_588);
and U1024 (N_1024,N_398,N_366);
nand U1025 (N_1025,N_947,N_194);
nand U1026 (N_1026,N_449,N_486);
nor U1027 (N_1027,N_81,N_991);
nor U1028 (N_1028,N_318,N_276);
or U1029 (N_1029,N_162,N_746);
and U1030 (N_1030,N_802,N_670);
nand U1031 (N_1031,N_765,N_560);
or U1032 (N_1032,N_152,N_48);
nor U1033 (N_1033,N_279,N_774);
or U1034 (N_1034,N_798,N_756);
or U1035 (N_1035,N_264,N_552);
and U1036 (N_1036,N_703,N_754);
or U1037 (N_1037,N_858,N_102);
nor U1038 (N_1038,N_241,N_381);
nand U1039 (N_1039,N_572,N_755);
nor U1040 (N_1040,N_474,N_21);
or U1041 (N_1041,N_416,N_826);
or U1042 (N_1042,N_729,N_543);
xnor U1043 (N_1043,N_738,N_614);
or U1044 (N_1044,N_863,N_38);
nand U1045 (N_1045,N_663,N_659);
xor U1046 (N_1046,N_996,N_35);
nor U1047 (N_1047,N_460,N_549);
nor U1048 (N_1048,N_740,N_862);
or U1049 (N_1049,N_520,N_396);
or U1050 (N_1050,N_444,N_469);
or U1051 (N_1051,N_491,N_0);
nor U1052 (N_1052,N_187,N_333);
nand U1053 (N_1053,N_28,N_232);
nor U1054 (N_1054,N_646,N_626);
and U1055 (N_1055,N_301,N_104);
nor U1056 (N_1056,N_482,N_843);
and U1057 (N_1057,N_7,N_977);
nand U1058 (N_1058,N_712,N_294);
nand U1059 (N_1059,N_155,N_682);
and U1060 (N_1060,N_983,N_849);
or U1061 (N_1061,N_950,N_457);
nand U1062 (N_1062,N_37,N_54);
or U1063 (N_1063,N_511,N_405);
and U1064 (N_1064,N_693,N_424);
and U1065 (N_1065,N_314,N_694);
nor U1066 (N_1066,N_466,N_379);
nand U1067 (N_1067,N_696,N_33);
and U1068 (N_1068,N_368,N_46);
and U1069 (N_1069,N_837,N_408);
nor U1070 (N_1070,N_321,N_404);
nor U1071 (N_1071,N_807,N_923);
and U1072 (N_1072,N_135,N_395);
xor U1073 (N_1073,N_822,N_870);
nor U1074 (N_1074,N_804,N_69);
nand U1075 (N_1075,N_496,N_391);
or U1076 (N_1076,N_954,N_539);
or U1077 (N_1077,N_850,N_4);
nand U1078 (N_1078,N_43,N_953);
nor U1079 (N_1079,N_574,N_845);
nand U1080 (N_1080,N_838,N_213);
nand U1081 (N_1081,N_372,N_906);
or U1082 (N_1082,N_943,N_867);
and U1083 (N_1083,N_642,N_675);
and U1084 (N_1084,N_12,N_847);
nand U1085 (N_1085,N_132,N_230);
and U1086 (N_1086,N_128,N_402);
nand U1087 (N_1087,N_591,N_624);
nor U1088 (N_1088,N_172,N_175);
or U1089 (N_1089,N_309,N_226);
nor U1090 (N_1090,N_79,N_188);
nand U1091 (N_1091,N_205,N_914);
and U1092 (N_1092,N_358,N_32);
or U1093 (N_1093,N_665,N_470);
and U1094 (N_1094,N_208,N_65);
nand U1095 (N_1095,N_251,N_744);
or U1096 (N_1096,N_242,N_620);
nor U1097 (N_1097,N_999,N_655);
nand U1098 (N_1098,N_699,N_958);
nand U1099 (N_1099,N_422,N_742);
nand U1100 (N_1100,N_23,N_970);
and U1101 (N_1101,N_978,N_758);
and U1102 (N_1102,N_553,N_471);
nand U1103 (N_1103,N_489,N_165);
and U1104 (N_1104,N_692,N_218);
nand U1105 (N_1105,N_566,N_13);
nor U1106 (N_1106,N_210,N_153);
nor U1107 (N_1107,N_394,N_736);
and U1108 (N_1108,N_965,N_779);
and U1109 (N_1109,N_903,N_115);
nand U1110 (N_1110,N_722,N_201);
nor U1111 (N_1111,N_877,N_963);
or U1112 (N_1112,N_537,N_141);
or U1113 (N_1113,N_564,N_435);
or U1114 (N_1114,N_308,N_635);
nand U1115 (N_1115,N_417,N_322);
or U1116 (N_1116,N_487,N_897);
nand U1117 (N_1117,N_446,N_691);
and U1118 (N_1118,N_993,N_180);
nand U1119 (N_1119,N_973,N_500);
and U1120 (N_1120,N_982,N_16);
and U1121 (N_1121,N_558,N_428);
and U1122 (N_1122,N_270,N_91);
nand U1123 (N_1123,N_501,N_618);
nor U1124 (N_1124,N_669,N_995);
nor U1125 (N_1125,N_932,N_812);
nor U1126 (N_1126,N_476,N_881);
nor U1127 (N_1127,N_448,N_687);
nand U1128 (N_1128,N_595,N_203);
nor U1129 (N_1129,N_854,N_179);
or U1130 (N_1130,N_632,N_362);
nand U1131 (N_1131,N_83,N_787);
and U1132 (N_1132,N_835,N_832);
and U1133 (N_1133,N_727,N_250);
and U1134 (N_1134,N_206,N_431);
nand U1135 (N_1135,N_393,N_894);
or U1136 (N_1136,N_582,N_26);
and U1137 (N_1137,N_904,N_505);
or U1138 (N_1138,N_168,N_525);
or U1139 (N_1139,N_613,N_374);
nor U1140 (N_1140,N_370,N_445);
nand U1141 (N_1141,N_283,N_77);
nor U1142 (N_1142,N_129,N_150);
nand U1143 (N_1143,N_523,N_545);
or U1144 (N_1144,N_781,N_600);
and U1145 (N_1145,N_8,N_258);
and U1146 (N_1146,N_96,N_89);
nor U1147 (N_1147,N_979,N_879);
nand U1148 (N_1148,N_484,N_355);
or U1149 (N_1149,N_608,N_71);
or U1150 (N_1150,N_938,N_820);
nor U1151 (N_1151,N_430,N_698);
nand U1152 (N_1152,N_184,N_956);
nor U1153 (N_1153,N_823,N_942);
or U1154 (N_1154,N_793,N_481);
or U1155 (N_1155,N_610,N_328);
xor U1156 (N_1156,N_809,N_332);
and U1157 (N_1157,N_516,N_522);
nand U1158 (N_1158,N_195,N_778);
or U1159 (N_1159,N_936,N_593);
nor U1160 (N_1160,N_711,N_262);
and U1161 (N_1161,N_714,N_299);
nand U1162 (N_1162,N_719,N_792);
xor U1163 (N_1163,N_578,N_361);
nor U1164 (N_1164,N_266,N_263);
nor U1165 (N_1165,N_327,N_454);
nor U1166 (N_1166,N_625,N_890);
nor U1167 (N_1167,N_493,N_645);
or U1168 (N_1168,N_151,N_36);
or U1169 (N_1169,N_688,N_127);
or U1170 (N_1170,N_873,N_64);
nor U1171 (N_1171,N_944,N_531);
nand U1172 (N_1172,N_783,N_312);
nand U1173 (N_1173,N_427,N_580);
nand U1174 (N_1174,N_173,N_341);
nor U1175 (N_1175,N_211,N_57);
nand U1176 (N_1176,N_926,N_479);
nor U1177 (N_1177,N_750,N_842);
and U1178 (N_1178,N_653,N_869);
nor U1179 (N_1179,N_410,N_419);
xor U1180 (N_1180,N_74,N_627);
nor U1181 (N_1181,N_751,N_42);
or U1182 (N_1182,N_273,N_737);
and U1183 (N_1183,N_159,N_528);
and U1184 (N_1184,N_229,N_384);
or U1185 (N_1185,N_799,N_900);
nor U1186 (N_1186,N_930,N_868);
and U1187 (N_1187,N_291,N_828);
nor U1188 (N_1188,N_243,N_452);
nand U1189 (N_1189,N_24,N_371);
nand U1190 (N_1190,N_640,N_246);
or U1191 (N_1191,N_612,N_677);
nor U1192 (N_1192,N_733,N_643);
or U1193 (N_1193,N_514,N_93);
and U1194 (N_1194,N_725,N_51);
nor U1195 (N_1195,N_388,N_498);
nor U1196 (N_1196,N_401,N_878);
and U1197 (N_1197,N_617,N_284);
nand U1198 (N_1198,N_885,N_443);
and U1199 (N_1199,N_217,N_922);
nand U1200 (N_1200,N_536,N_542);
and U1201 (N_1201,N_386,N_782);
xor U1202 (N_1202,N_403,N_800);
and U1203 (N_1203,N_785,N_925);
nand U1204 (N_1204,N_198,N_437);
or U1205 (N_1205,N_376,N_145);
or U1206 (N_1206,N_569,N_61);
or U1207 (N_1207,N_30,N_62);
or U1208 (N_1208,N_757,N_976);
nor U1209 (N_1209,N_860,N_356);
nor U1210 (N_1210,N_654,N_87);
nand U1211 (N_1211,N_865,N_161);
nor U1212 (N_1212,N_360,N_931);
nor U1213 (N_1213,N_636,N_777);
nand U1214 (N_1214,N_607,N_507);
nand U1215 (N_1215,N_550,N_546);
nand U1216 (N_1216,N_88,N_534);
nor U1217 (N_1217,N_584,N_256);
nand U1218 (N_1218,N_95,N_154);
nor U1219 (N_1219,N_197,N_724);
and U1220 (N_1220,N_859,N_939);
nor U1221 (N_1221,N_921,N_690);
nand U1222 (N_1222,N_700,N_794);
and U1223 (N_1223,N_510,N_648);
and U1224 (N_1224,N_429,N_888);
or U1225 (N_1225,N_351,N_49);
nand U1226 (N_1226,N_805,N_14);
and U1227 (N_1227,N_269,N_120);
and U1228 (N_1228,N_801,N_293);
nor U1229 (N_1229,N_941,N_415);
and U1230 (N_1230,N_816,N_236);
and U1231 (N_1231,N_27,N_167);
nor U1232 (N_1232,N_465,N_667);
nand U1233 (N_1233,N_767,N_85);
nand U1234 (N_1234,N_323,N_960);
and U1235 (N_1235,N_156,N_108);
nor U1236 (N_1236,N_840,N_726);
nand U1237 (N_1237,N_772,N_331);
nor U1238 (N_1238,N_106,N_515);
nand U1239 (N_1239,N_573,N_228);
and U1240 (N_1240,N_409,N_780);
or U1241 (N_1241,N_946,N_66);
nand U1242 (N_1242,N_260,N_606);
nor U1243 (N_1243,N_193,N_604);
nand U1244 (N_1244,N_615,N_234);
nor U1245 (N_1245,N_125,N_502);
and U1246 (N_1246,N_53,N_439);
and U1247 (N_1247,N_296,N_363);
nor U1248 (N_1248,N_257,N_597);
nor U1249 (N_1249,N_909,N_559);
nor U1250 (N_1250,N_303,N_238);
or U1251 (N_1251,N_784,N_40);
or U1252 (N_1252,N_347,N_771);
nor U1253 (N_1253,N_821,N_22);
xor U1254 (N_1254,N_247,N_806);
nand U1255 (N_1255,N_86,N_883);
nor U1256 (N_1256,N_92,N_796);
nand U1257 (N_1257,N_789,N_275);
or U1258 (N_1258,N_680,N_111);
or U1259 (N_1259,N_907,N_997);
nand U1260 (N_1260,N_852,N_240);
nor U1261 (N_1261,N_715,N_373);
nand U1262 (N_1262,N_810,N_773);
nor U1263 (N_1263,N_412,N_519);
and U1264 (N_1264,N_335,N_998);
nand U1265 (N_1265,N_60,N_107);
nor U1266 (N_1266,N_18,N_329);
nor U1267 (N_1267,N_532,N_836);
and U1268 (N_1268,N_629,N_683);
or U1269 (N_1269,N_59,N_399);
nand U1270 (N_1270,N_813,N_9);
and U1271 (N_1271,N_307,N_192);
and U1272 (N_1272,N_720,N_55);
nand U1273 (N_1273,N_311,N_400);
xor U1274 (N_1274,N_652,N_815);
or U1275 (N_1275,N_686,N_529);
and U1276 (N_1276,N_5,N_786);
or U1277 (N_1277,N_577,N_178);
nand U1278 (N_1278,N_186,N_948);
or U1279 (N_1279,N_472,N_524);
xor U1280 (N_1280,N_143,N_492);
or U1281 (N_1281,N_124,N_298);
nand U1282 (N_1282,N_350,N_344);
nand U1283 (N_1283,N_34,N_31);
and U1284 (N_1284,N_752,N_834);
and U1285 (N_1285,N_237,N_819);
nor U1286 (N_1286,N_585,N_245);
and U1287 (N_1287,N_920,N_547);
or U1288 (N_1288,N_349,N_506);
and U1289 (N_1289,N_281,N_641);
or U1290 (N_1290,N_764,N_679);
and U1291 (N_1291,N_44,N_908);
or U1292 (N_1292,N_451,N_222);
or U1293 (N_1293,N_252,N_512);
xnor U1294 (N_1294,N_662,N_933);
or U1295 (N_1295,N_568,N_11);
nand U1296 (N_1296,N_684,N_319);
nor U1297 (N_1297,N_105,N_418);
nor U1298 (N_1298,N_39,N_880);
or U1299 (N_1299,N_535,N_775);
nand U1300 (N_1300,N_110,N_112);
nand U1301 (N_1301,N_45,N_78);
nor U1302 (N_1302,N_717,N_919);
nand U1303 (N_1303,N_587,N_274);
and U1304 (N_1304,N_488,N_109);
nor U1305 (N_1305,N_200,N_884);
and U1306 (N_1306,N_576,N_825);
or U1307 (N_1307,N_503,N_338);
nand U1308 (N_1308,N_872,N_456);
or U1309 (N_1309,N_113,N_138);
and U1310 (N_1310,N_716,N_509);
nand U1311 (N_1311,N_962,N_177);
and U1312 (N_1312,N_940,N_817);
nor U1313 (N_1313,N_436,N_841);
nand U1314 (N_1314,N_876,N_901);
xor U1315 (N_1315,N_839,N_121);
or U1316 (N_1316,N_285,N_434);
nor U1317 (N_1317,N_317,N_440);
or U1318 (N_1318,N_389,N_286);
and U1319 (N_1319,N_829,N_123);
or U1320 (N_1320,N_557,N_392);
nand U1321 (N_1321,N_985,N_814);
nand U1322 (N_1322,N_769,N_297);
and U1323 (N_1323,N_477,N_204);
nor U1324 (N_1324,N_267,N_526);
and U1325 (N_1325,N_499,N_898);
nand U1326 (N_1326,N_310,N_721);
or U1327 (N_1327,N_171,N_146);
and U1328 (N_1328,N_882,N_548);
or U1329 (N_1329,N_887,N_413);
or U1330 (N_1330,N_735,N_934);
nand U1331 (N_1331,N_334,N_455);
nor U1332 (N_1332,N_75,N_330);
nor U1333 (N_1333,N_795,N_136);
nor U1334 (N_1334,N_739,N_831);
and U1335 (N_1335,N_411,N_369);
nor U1336 (N_1336,N_598,N_98);
or U1337 (N_1337,N_745,N_853);
nand U1338 (N_1338,N_567,N_540);
nor U1339 (N_1339,N_433,N_357);
and U1340 (N_1340,N_216,N_660);
nand U1341 (N_1341,N_56,N_117);
nor U1342 (N_1342,N_20,N_857);
and U1343 (N_1343,N_17,N_749);
or U1344 (N_1344,N_271,N_280);
nand U1345 (N_1345,N_131,N_565);
and U1346 (N_1346,N_517,N_987);
nor U1347 (N_1347,N_342,N_732);
nand U1348 (N_1348,N_685,N_214);
xor U1349 (N_1349,N_495,N_592);
nand U1350 (N_1350,N_191,N_268);
and U1351 (N_1351,N_899,N_972);
nand U1352 (N_1352,N_3,N_975);
nor U1353 (N_1353,N_718,N_289);
or U1354 (N_1354,N_974,N_438);
nand U1355 (N_1355,N_461,N_855);
nand U1356 (N_1356,N_300,N_29);
nor U1357 (N_1357,N_80,N_609);
or U1358 (N_1358,N_657,N_354);
nor U1359 (N_1359,N_352,N_917);
and U1360 (N_1360,N_119,N_530);
nor U1361 (N_1361,N_380,N_555);
nand U1362 (N_1362,N_730,N_741);
and U1363 (N_1363,N_114,N_916);
and U1364 (N_1364,N_72,N_695);
nor U1365 (N_1365,N_575,N_15);
or U1366 (N_1366,N_326,N_52);
nand U1367 (N_1367,N_760,N_989);
or U1368 (N_1368,N_377,N_340);
nor U1369 (N_1369,N_345,N_689);
nand U1370 (N_1370,N_704,N_485);
or U1371 (N_1371,N_833,N_101);
and U1372 (N_1372,N_551,N_76);
and U1373 (N_1373,N_896,N_248);
and U1374 (N_1374,N_874,N_619);
or U1375 (N_1375,N_731,N_571);
and U1376 (N_1376,N_255,N_981);
nand U1377 (N_1377,N_325,N_994);
nand U1378 (N_1378,N_912,N_227);
nand U1379 (N_1379,N_1,N_728);
or U1380 (N_1380,N_966,N_346);
or U1381 (N_1381,N_935,N_464);
or U1382 (N_1382,N_490,N_463);
nand U1383 (N_1383,N_631,N_803);
or U1384 (N_1384,N_601,N_992);
xor U1385 (N_1385,N_518,N_126);
nor U1386 (N_1386,N_678,N_148);
nor U1387 (N_1387,N_259,N_827);
nand U1388 (N_1388,N_527,N_459);
or U1389 (N_1389,N_302,N_673);
nand U1390 (N_1390,N_924,N_915);
nand U1391 (N_1391,N_776,N_189);
and U1392 (N_1392,N_599,N_292);
or U1393 (N_1393,N_570,N_157);
or U1394 (N_1394,N_927,N_462);
nor U1395 (N_1395,N_364,N_209);
and U1396 (N_1396,N_713,N_701);
nor U1397 (N_1397,N_304,N_945);
or U1398 (N_1398,N_10,N_766);
and U1399 (N_1399,N_359,N_748);
nand U1400 (N_1400,N_556,N_249);
nor U1401 (N_1401,N_637,N_911);
xor U1402 (N_1402,N_160,N_681);
nand U1403 (N_1403,N_589,N_99);
and U1404 (N_1404,N_891,N_324);
nor U1405 (N_1405,N_759,N_761);
or U1406 (N_1406,N_447,N_199);
nor U1407 (N_1407,N_19,N_697);
or U1408 (N_1408,N_140,N_658);
and U1409 (N_1409,N_181,N_282);
or U1410 (N_1410,N_339,N_82);
nand U1411 (N_1411,N_158,N_533);
nor U1412 (N_1412,N_497,N_202);
nor U1413 (N_1413,N_277,N_94);
nand U1414 (N_1414,N_442,N_420);
nor U1415 (N_1415,N_951,N_949);
nor U1416 (N_1416,N_818,N_233);
and U1417 (N_1417,N_223,N_287);
xnor U1418 (N_1418,N_70,N_174);
nor U1419 (N_1419,N_478,N_467);
or U1420 (N_1420,N_219,N_622);
nand U1421 (N_1421,N_710,N_142);
nand U1422 (N_1422,N_163,N_382);
xor U1423 (N_1423,N_207,N_475);
and U1424 (N_1424,N_235,N_541);
nor U1425 (N_1425,N_353,N_494);
nor U1426 (N_1426,N_886,N_383);
and U1427 (N_1427,N_130,N_768);
nand U1428 (N_1428,N_133,N_139);
or U1429 (N_1429,N_708,N_137);
or U1430 (N_1430,N_709,N_928);
nor U1431 (N_1431,N_603,N_889);
and U1432 (N_1432,N_378,N_633);
nand U1433 (N_1433,N_290,N_483);
nand U1434 (N_1434,N_504,N_929);
nand U1435 (N_1435,N_73,N_423);
or U1436 (N_1436,N_134,N_103);
and U1437 (N_1437,N_705,N_770);
nor U1438 (N_1438,N_336,N_902);
nand U1439 (N_1439,N_183,N_170);
or U1440 (N_1440,N_762,N_554);
and U1441 (N_1441,N_25,N_586);
nor U1442 (N_1442,N_147,N_952);
and U1443 (N_1443,N_986,N_650);
nor U1444 (N_1444,N_190,N_561);
nand U1445 (N_1445,N_651,N_116);
nor U1446 (N_1446,N_583,N_68);
and U1447 (N_1447,N_808,N_790);
nor U1448 (N_1448,N_2,N_581);
nand U1449 (N_1449,N_666,N_984);
nand U1450 (N_1450,N_628,N_97);
or U1451 (N_1451,N_414,N_967);
and U1452 (N_1452,N_674,N_937);
or U1453 (N_1453,N_315,N_231);
or U1454 (N_1454,N_955,N_367);
or U1455 (N_1455,N_791,N_47);
or U1456 (N_1456,N_458,N_432);
or U1457 (N_1457,N_305,N_851);
or U1458 (N_1458,N_656,N_959);
and U1459 (N_1459,N_390,N_182);
nor U1460 (N_1460,N_616,N_176);
or U1461 (N_1461,N_957,N_453);
or U1462 (N_1462,N_811,N_747);
and U1463 (N_1463,N_254,N_830);
or U1464 (N_1464,N_337,N_988);
nor U1465 (N_1465,N_320,N_630);
nand U1466 (N_1466,N_893,N_425);
or U1467 (N_1467,N_702,N_306);
nand U1468 (N_1468,N_295,N_313);
nand U1469 (N_1469,N_224,N_611);
nor U1470 (N_1470,N_50,N_596);
xnor U1471 (N_1471,N_196,N_468);
or U1472 (N_1472,N_824,N_990);
nand U1473 (N_1473,N_621,N_910);
or U1474 (N_1474,N_634,N_707);
nand U1475 (N_1475,N_100,N_639);
nor U1476 (N_1476,N_149,N_671);
nand U1477 (N_1477,N_67,N_664);
nand U1478 (N_1478,N_375,N_964);
nor U1479 (N_1479,N_441,N_856);
nand U1480 (N_1480,N_892,N_579);
nand U1481 (N_1481,N_343,N_397);
nand U1482 (N_1482,N_118,N_875);
nand U1483 (N_1483,N_866,N_968);
or U1484 (N_1484,N_239,N_288);
nor U1485 (N_1485,N_272,N_508);
nand U1486 (N_1486,N_480,N_421);
and U1487 (N_1487,N_58,N_676);
nand U1488 (N_1488,N_253,N_743);
and U1489 (N_1489,N_788,N_41);
nor U1490 (N_1490,N_644,N_450);
or U1491 (N_1491,N_426,N_723);
nor U1492 (N_1492,N_225,N_212);
nand U1493 (N_1493,N_406,N_265);
nand U1494 (N_1494,N_563,N_971);
nor U1495 (N_1495,N_969,N_864);
or U1496 (N_1496,N_846,N_668);
nand U1497 (N_1497,N_590,N_913);
and U1498 (N_1498,N_365,N_562);
or U1499 (N_1499,N_538,N_185);
nand U1500 (N_1500,N_496,N_634);
nor U1501 (N_1501,N_169,N_63);
and U1502 (N_1502,N_294,N_26);
nand U1503 (N_1503,N_509,N_969);
nor U1504 (N_1504,N_196,N_360);
or U1505 (N_1505,N_446,N_225);
nand U1506 (N_1506,N_533,N_432);
nand U1507 (N_1507,N_347,N_769);
and U1508 (N_1508,N_281,N_844);
nand U1509 (N_1509,N_123,N_106);
nor U1510 (N_1510,N_227,N_192);
nor U1511 (N_1511,N_399,N_385);
and U1512 (N_1512,N_315,N_886);
nand U1513 (N_1513,N_959,N_750);
nor U1514 (N_1514,N_945,N_759);
and U1515 (N_1515,N_674,N_432);
or U1516 (N_1516,N_291,N_411);
and U1517 (N_1517,N_422,N_432);
or U1518 (N_1518,N_248,N_366);
and U1519 (N_1519,N_753,N_180);
nor U1520 (N_1520,N_29,N_928);
and U1521 (N_1521,N_63,N_698);
and U1522 (N_1522,N_860,N_276);
nor U1523 (N_1523,N_851,N_591);
and U1524 (N_1524,N_905,N_438);
nand U1525 (N_1525,N_211,N_165);
nor U1526 (N_1526,N_203,N_748);
nor U1527 (N_1527,N_471,N_315);
and U1528 (N_1528,N_687,N_867);
or U1529 (N_1529,N_588,N_259);
or U1530 (N_1530,N_229,N_494);
or U1531 (N_1531,N_121,N_530);
and U1532 (N_1532,N_130,N_211);
nor U1533 (N_1533,N_124,N_290);
and U1534 (N_1534,N_996,N_731);
nor U1535 (N_1535,N_260,N_923);
nor U1536 (N_1536,N_354,N_726);
nor U1537 (N_1537,N_967,N_261);
or U1538 (N_1538,N_836,N_717);
or U1539 (N_1539,N_864,N_872);
or U1540 (N_1540,N_500,N_423);
and U1541 (N_1541,N_152,N_535);
and U1542 (N_1542,N_793,N_893);
nand U1543 (N_1543,N_288,N_911);
nand U1544 (N_1544,N_41,N_188);
xnor U1545 (N_1545,N_91,N_53);
nor U1546 (N_1546,N_910,N_104);
or U1547 (N_1547,N_834,N_942);
nand U1548 (N_1548,N_358,N_840);
and U1549 (N_1549,N_305,N_898);
nand U1550 (N_1550,N_544,N_686);
nand U1551 (N_1551,N_823,N_871);
nand U1552 (N_1552,N_655,N_475);
nor U1553 (N_1553,N_168,N_492);
or U1554 (N_1554,N_508,N_664);
nor U1555 (N_1555,N_777,N_16);
nand U1556 (N_1556,N_787,N_688);
nand U1557 (N_1557,N_910,N_451);
nand U1558 (N_1558,N_613,N_156);
nor U1559 (N_1559,N_981,N_169);
or U1560 (N_1560,N_417,N_885);
nor U1561 (N_1561,N_248,N_493);
nor U1562 (N_1562,N_429,N_428);
nand U1563 (N_1563,N_73,N_801);
nand U1564 (N_1564,N_801,N_679);
and U1565 (N_1565,N_44,N_430);
nor U1566 (N_1566,N_75,N_155);
and U1567 (N_1567,N_749,N_903);
nand U1568 (N_1568,N_539,N_255);
nand U1569 (N_1569,N_666,N_469);
and U1570 (N_1570,N_651,N_909);
nand U1571 (N_1571,N_173,N_17);
and U1572 (N_1572,N_690,N_463);
or U1573 (N_1573,N_939,N_812);
xor U1574 (N_1574,N_562,N_72);
nand U1575 (N_1575,N_581,N_408);
or U1576 (N_1576,N_459,N_6);
and U1577 (N_1577,N_371,N_377);
nor U1578 (N_1578,N_82,N_826);
nor U1579 (N_1579,N_429,N_339);
nor U1580 (N_1580,N_963,N_500);
nor U1581 (N_1581,N_913,N_206);
nand U1582 (N_1582,N_983,N_161);
nor U1583 (N_1583,N_133,N_932);
and U1584 (N_1584,N_686,N_97);
and U1585 (N_1585,N_707,N_376);
nor U1586 (N_1586,N_949,N_214);
nor U1587 (N_1587,N_667,N_361);
nand U1588 (N_1588,N_516,N_795);
and U1589 (N_1589,N_969,N_71);
or U1590 (N_1590,N_964,N_603);
and U1591 (N_1591,N_680,N_958);
nand U1592 (N_1592,N_303,N_20);
or U1593 (N_1593,N_261,N_856);
or U1594 (N_1594,N_101,N_595);
nor U1595 (N_1595,N_233,N_35);
nor U1596 (N_1596,N_851,N_21);
and U1597 (N_1597,N_722,N_927);
and U1598 (N_1598,N_740,N_551);
nand U1599 (N_1599,N_520,N_366);
nand U1600 (N_1600,N_284,N_408);
or U1601 (N_1601,N_462,N_472);
or U1602 (N_1602,N_294,N_449);
and U1603 (N_1603,N_598,N_26);
nand U1604 (N_1604,N_964,N_411);
nor U1605 (N_1605,N_338,N_387);
or U1606 (N_1606,N_427,N_964);
nand U1607 (N_1607,N_503,N_463);
nor U1608 (N_1608,N_179,N_641);
nand U1609 (N_1609,N_511,N_73);
and U1610 (N_1610,N_388,N_560);
or U1611 (N_1611,N_450,N_697);
or U1612 (N_1612,N_816,N_878);
or U1613 (N_1613,N_801,N_432);
nor U1614 (N_1614,N_709,N_489);
and U1615 (N_1615,N_898,N_926);
nand U1616 (N_1616,N_725,N_949);
nor U1617 (N_1617,N_135,N_578);
nand U1618 (N_1618,N_408,N_253);
nand U1619 (N_1619,N_827,N_183);
nand U1620 (N_1620,N_426,N_429);
nor U1621 (N_1621,N_186,N_206);
nand U1622 (N_1622,N_215,N_363);
xnor U1623 (N_1623,N_738,N_459);
and U1624 (N_1624,N_274,N_196);
xnor U1625 (N_1625,N_67,N_239);
or U1626 (N_1626,N_928,N_861);
and U1627 (N_1627,N_811,N_993);
nor U1628 (N_1628,N_398,N_599);
nand U1629 (N_1629,N_411,N_132);
and U1630 (N_1630,N_292,N_114);
nand U1631 (N_1631,N_854,N_177);
nor U1632 (N_1632,N_997,N_150);
and U1633 (N_1633,N_945,N_830);
nor U1634 (N_1634,N_982,N_232);
nand U1635 (N_1635,N_400,N_78);
or U1636 (N_1636,N_70,N_350);
nand U1637 (N_1637,N_138,N_429);
or U1638 (N_1638,N_260,N_83);
nand U1639 (N_1639,N_234,N_897);
nand U1640 (N_1640,N_387,N_594);
or U1641 (N_1641,N_533,N_430);
and U1642 (N_1642,N_838,N_945);
and U1643 (N_1643,N_27,N_664);
nor U1644 (N_1644,N_763,N_416);
and U1645 (N_1645,N_106,N_230);
nand U1646 (N_1646,N_463,N_369);
and U1647 (N_1647,N_52,N_328);
or U1648 (N_1648,N_337,N_390);
nand U1649 (N_1649,N_697,N_448);
nor U1650 (N_1650,N_796,N_730);
nor U1651 (N_1651,N_915,N_886);
nor U1652 (N_1652,N_290,N_181);
or U1653 (N_1653,N_310,N_416);
nand U1654 (N_1654,N_626,N_822);
or U1655 (N_1655,N_263,N_254);
nand U1656 (N_1656,N_421,N_453);
nor U1657 (N_1657,N_833,N_664);
or U1658 (N_1658,N_815,N_608);
nand U1659 (N_1659,N_454,N_47);
or U1660 (N_1660,N_355,N_216);
nand U1661 (N_1661,N_872,N_269);
nand U1662 (N_1662,N_59,N_157);
or U1663 (N_1663,N_0,N_6);
nor U1664 (N_1664,N_779,N_94);
nor U1665 (N_1665,N_378,N_553);
or U1666 (N_1666,N_825,N_137);
or U1667 (N_1667,N_47,N_829);
nand U1668 (N_1668,N_605,N_748);
nor U1669 (N_1669,N_140,N_971);
and U1670 (N_1670,N_597,N_916);
and U1671 (N_1671,N_589,N_531);
or U1672 (N_1672,N_407,N_232);
or U1673 (N_1673,N_76,N_65);
and U1674 (N_1674,N_262,N_452);
nor U1675 (N_1675,N_450,N_99);
nor U1676 (N_1676,N_307,N_976);
and U1677 (N_1677,N_955,N_385);
or U1678 (N_1678,N_299,N_334);
and U1679 (N_1679,N_892,N_527);
or U1680 (N_1680,N_584,N_291);
and U1681 (N_1681,N_864,N_398);
and U1682 (N_1682,N_879,N_399);
nor U1683 (N_1683,N_87,N_949);
nand U1684 (N_1684,N_676,N_664);
or U1685 (N_1685,N_812,N_930);
nor U1686 (N_1686,N_689,N_870);
nand U1687 (N_1687,N_775,N_979);
and U1688 (N_1688,N_202,N_883);
or U1689 (N_1689,N_925,N_765);
nand U1690 (N_1690,N_155,N_532);
nand U1691 (N_1691,N_41,N_725);
nor U1692 (N_1692,N_333,N_202);
and U1693 (N_1693,N_63,N_580);
nor U1694 (N_1694,N_664,N_263);
or U1695 (N_1695,N_612,N_515);
and U1696 (N_1696,N_525,N_830);
nor U1697 (N_1697,N_66,N_911);
and U1698 (N_1698,N_821,N_484);
or U1699 (N_1699,N_266,N_288);
nor U1700 (N_1700,N_808,N_861);
xnor U1701 (N_1701,N_204,N_633);
nand U1702 (N_1702,N_37,N_345);
nand U1703 (N_1703,N_800,N_317);
and U1704 (N_1704,N_887,N_785);
nand U1705 (N_1705,N_550,N_282);
nand U1706 (N_1706,N_148,N_325);
nand U1707 (N_1707,N_159,N_199);
nor U1708 (N_1708,N_912,N_81);
nand U1709 (N_1709,N_43,N_164);
or U1710 (N_1710,N_131,N_442);
or U1711 (N_1711,N_671,N_282);
and U1712 (N_1712,N_634,N_862);
and U1713 (N_1713,N_110,N_979);
or U1714 (N_1714,N_704,N_406);
or U1715 (N_1715,N_719,N_371);
and U1716 (N_1716,N_810,N_561);
or U1717 (N_1717,N_361,N_671);
nand U1718 (N_1718,N_553,N_426);
or U1719 (N_1719,N_971,N_189);
xnor U1720 (N_1720,N_658,N_94);
and U1721 (N_1721,N_133,N_580);
nor U1722 (N_1722,N_752,N_700);
or U1723 (N_1723,N_858,N_207);
or U1724 (N_1724,N_735,N_725);
nand U1725 (N_1725,N_3,N_461);
and U1726 (N_1726,N_885,N_665);
nand U1727 (N_1727,N_625,N_322);
nand U1728 (N_1728,N_827,N_848);
nand U1729 (N_1729,N_9,N_686);
and U1730 (N_1730,N_460,N_796);
nor U1731 (N_1731,N_85,N_668);
or U1732 (N_1732,N_500,N_759);
xor U1733 (N_1733,N_679,N_454);
nor U1734 (N_1734,N_973,N_131);
and U1735 (N_1735,N_653,N_191);
and U1736 (N_1736,N_543,N_181);
and U1737 (N_1737,N_915,N_688);
nor U1738 (N_1738,N_779,N_78);
or U1739 (N_1739,N_881,N_988);
or U1740 (N_1740,N_978,N_209);
or U1741 (N_1741,N_687,N_284);
nor U1742 (N_1742,N_662,N_292);
or U1743 (N_1743,N_610,N_384);
or U1744 (N_1744,N_970,N_100);
nand U1745 (N_1745,N_772,N_390);
and U1746 (N_1746,N_311,N_692);
and U1747 (N_1747,N_291,N_212);
and U1748 (N_1748,N_985,N_603);
nor U1749 (N_1749,N_913,N_204);
or U1750 (N_1750,N_199,N_136);
nand U1751 (N_1751,N_550,N_242);
nor U1752 (N_1752,N_239,N_504);
nand U1753 (N_1753,N_899,N_908);
nor U1754 (N_1754,N_179,N_998);
nor U1755 (N_1755,N_616,N_881);
or U1756 (N_1756,N_43,N_325);
or U1757 (N_1757,N_942,N_332);
and U1758 (N_1758,N_94,N_480);
nor U1759 (N_1759,N_428,N_397);
nor U1760 (N_1760,N_679,N_740);
nor U1761 (N_1761,N_495,N_960);
nor U1762 (N_1762,N_450,N_97);
nor U1763 (N_1763,N_33,N_551);
or U1764 (N_1764,N_213,N_112);
and U1765 (N_1765,N_746,N_330);
nand U1766 (N_1766,N_761,N_835);
or U1767 (N_1767,N_218,N_528);
nor U1768 (N_1768,N_660,N_954);
nand U1769 (N_1769,N_231,N_472);
nor U1770 (N_1770,N_961,N_179);
and U1771 (N_1771,N_644,N_172);
nand U1772 (N_1772,N_425,N_859);
nand U1773 (N_1773,N_871,N_916);
nand U1774 (N_1774,N_995,N_358);
nor U1775 (N_1775,N_99,N_36);
nor U1776 (N_1776,N_80,N_849);
or U1777 (N_1777,N_757,N_844);
nand U1778 (N_1778,N_565,N_503);
or U1779 (N_1779,N_327,N_672);
and U1780 (N_1780,N_912,N_246);
nand U1781 (N_1781,N_527,N_736);
xor U1782 (N_1782,N_124,N_338);
or U1783 (N_1783,N_352,N_635);
nand U1784 (N_1784,N_738,N_632);
or U1785 (N_1785,N_957,N_384);
nor U1786 (N_1786,N_998,N_952);
and U1787 (N_1787,N_213,N_961);
and U1788 (N_1788,N_488,N_220);
or U1789 (N_1789,N_45,N_115);
and U1790 (N_1790,N_170,N_139);
or U1791 (N_1791,N_723,N_983);
and U1792 (N_1792,N_164,N_992);
and U1793 (N_1793,N_650,N_284);
and U1794 (N_1794,N_985,N_397);
nand U1795 (N_1795,N_939,N_774);
nor U1796 (N_1796,N_852,N_796);
nor U1797 (N_1797,N_129,N_98);
and U1798 (N_1798,N_51,N_669);
nor U1799 (N_1799,N_790,N_968);
nand U1800 (N_1800,N_599,N_207);
nand U1801 (N_1801,N_191,N_982);
and U1802 (N_1802,N_940,N_412);
nor U1803 (N_1803,N_548,N_55);
xnor U1804 (N_1804,N_493,N_126);
nor U1805 (N_1805,N_658,N_365);
and U1806 (N_1806,N_198,N_712);
or U1807 (N_1807,N_146,N_603);
nand U1808 (N_1808,N_383,N_797);
nor U1809 (N_1809,N_294,N_93);
nand U1810 (N_1810,N_809,N_64);
and U1811 (N_1811,N_813,N_545);
and U1812 (N_1812,N_709,N_947);
and U1813 (N_1813,N_807,N_204);
nor U1814 (N_1814,N_340,N_109);
and U1815 (N_1815,N_184,N_303);
or U1816 (N_1816,N_116,N_826);
and U1817 (N_1817,N_154,N_315);
and U1818 (N_1818,N_899,N_737);
and U1819 (N_1819,N_520,N_203);
nor U1820 (N_1820,N_430,N_997);
nor U1821 (N_1821,N_673,N_811);
nand U1822 (N_1822,N_848,N_289);
and U1823 (N_1823,N_665,N_446);
nand U1824 (N_1824,N_600,N_509);
nand U1825 (N_1825,N_667,N_187);
nand U1826 (N_1826,N_809,N_240);
and U1827 (N_1827,N_616,N_576);
nor U1828 (N_1828,N_533,N_200);
or U1829 (N_1829,N_696,N_533);
and U1830 (N_1830,N_157,N_514);
and U1831 (N_1831,N_891,N_131);
and U1832 (N_1832,N_262,N_505);
or U1833 (N_1833,N_671,N_445);
or U1834 (N_1834,N_748,N_165);
nand U1835 (N_1835,N_619,N_228);
xor U1836 (N_1836,N_935,N_923);
and U1837 (N_1837,N_322,N_552);
and U1838 (N_1838,N_531,N_401);
and U1839 (N_1839,N_345,N_143);
or U1840 (N_1840,N_412,N_348);
or U1841 (N_1841,N_623,N_402);
and U1842 (N_1842,N_994,N_649);
and U1843 (N_1843,N_19,N_742);
or U1844 (N_1844,N_952,N_269);
nor U1845 (N_1845,N_952,N_442);
nand U1846 (N_1846,N_619,N_904);
and U1847 (N_1847,N_435,N_434);
or U1848 (N_1848,N_468,N_58);
nor U1849 (N_1849,N_514,N_189);
nor U1850 (N_1850,N_196,N_853);
and U1851 (N_1851,N_784,N_877);
or U1852 (N_1852,N_116,N_664);
or U1853 (N_1853,N_82,N_139);
or U1854 (N_1854,N_478,N_180);
nor U1855 (N_1855,N_610,N_289);
or U1856 (N_1856,N_736,N_511);
nor U1857 (N_1857,N_166,N_5);
or U1858 (N_1858,N_292,N_679);
or U1859 (N_1859,N_641,N_67);
nor U1860 (N_1860,N_646,N_593);
and U1861 (N_1861,N_328,N_414);
or U1862 (N_1862,N_974,N_944);
xor U1863 (N_1863,N_263,N_94);
and U1864 (N_1864,N_758,N_219);
or U1865 (N_1865,N_347,N_38);
or U1866 (N_1866,N_765,N_195);
or U1867 (N_1867,N_561,N_761);
nor U1868 (N_1868,N_337,N_449);
or U1869 (N_1869,N_645,N_884);
or U1870 (N_1870,N_699,N_531);
or U1871 (N_1871,N_380,N_720);
nand U1872 (N_1872,N_443,N_704);
xor U1873 (N_1873,N_119,N_336);
and U1874 (N_1874,N_567,N_641);
or U1875 (N_1875,N_455,N_861);
and U1876 (N_1876,N_464,N_754);
or U1877 (N_1877,N_340,N_561);
or U1878 (N_1878,N_997,N_512);
and U1879 (N_1879,N_824,N_330);
nand U1880 (N_1880,N_600,N_547);
or U1881 (N_1881,N_931,N_699);
nor U1882 (N_1882,N_991,N_118);
nor U1883 (N_1883,N_953,N_264);
and U1884 (N_1884,N_330,N_395);
and U1885 (N_1885,N_403,N_594);
or U1886 (N_1886,N_5,N_555);
or U1887 (N_1887,N_275,N_783);
nor U1888 (N_1888,N_436,N_365);
or U1889 (N_1889,N_894,N_206);
nand U1890 (N_1890,N_473,N_973);
or U1891 (N_1891,N_220,N_352);
nand U1892 (N_1892,N_321,N_569);
nor U1893 (N_1893,N_391,N_369);
or U1894 (N_1894,N_885,N_20);
or U1895 (N_1895,N_275,N_786);
or U1896 (N_1896,N_262,N_967);
nand U1897 (N_1897,N_489,N_967);
and U1898 (N_1898,N_269,N_408);
nand U1899 (N_1899,N_285,N_321);
nor U1900 (N_1900,N_24,N_10);
nand U1901 (N_1901,N_726,N_240);
and U1902 (N_1902,N_39,N_231);
or U1903 (N_1903,N_604,N_798);
or U1904 (N_1904,N_680,N_808);
nor U1905 (N_1905,N_817,N_665);
nor U1906 (N_1906,N_291,N_659);
nor U1907 (N_1907,N_973,N_525);
xnor U1908 (N_1908,N_292,N_340);
or U1909 (N_1909,N_754,N_773);
or U1910 (N_1910,N_884,N_364);
nand U1911 (N_1911,N_392,N_955);
or U1912 (N_1912,N_962,N_572);
nand U1913 (N_1913,N_270,N_831);
nand U1914 (N_1914,N_710,N_486);
nor U1915 (N_1915,N_574,N_962);
and U1916 (N_1916,N_450,N_378);
nand U1917 (N_1917,N_783,N_704);
nor U1918 (N_1918,N_548,N_509);
or U1919 (N_1919,N_469,N_798);
nor U1920 (N_1920,N_285,N_344);
and U1921 (N_1921,N_322,N_474);
nor U1922 (N_1922,N_436,N_590);
or U1923 (N_1923,N_257,N_580);
nand U1924 (N_1924,N_470,N_14);
nand U1925 (N_1925,N_286,N_206);
nor U1926 (N_1926,N_974,N_209);
and U1927 (N_1927,N_310,N_955);
nor U1928 (N_1928,N_593,N_971);
or U1929 (N_1929,N_384,N_82);
or U1930 (N_1930,N_410,N_382);
or U1931 (N_1931,N_707,N_851);
or U1932 (N_1932,N_384,N_588);
or U1933 (N_1933,N_120,N_602);
or U1934 (N_1934,N_719,N_528);
nand U1935 (N_1935,N_661,N_588);
and U1936 (N_1936,N_742,N_466);
nand U1937 (N_1937,N_646,N_864);
or U1938 (N_1938,N_591,N_674);
and U1939 (N_1939,N_771,N_220);
and U1940 (N_1940,N_600,N_797);
or U1941 (N_1941,N_24,N_516);
and U1942 (N_1942,N_514,N_530);
nand U1943 (N_1943,N_321,N_66);
and U1944 (N_1944,N_748,N_803);
or U1945 (N_1945,N_755,N_802);
nor U1946 (N_1946,N_262,N_214);
nor U1947 (N_1947,N_665,N_814);
and U1948 (N_1948,N_320,N_201);
and U1949 (N_1949,N_343,N_26);
or U1950 (N_1950,N_819,N_654);
or U1951 (N_1951,N_411,N_147);
and U1952 (N_1952,N_769,N_610);
nor U1953 (N_1953,N_135,N_170);
or U1954 (N_1954,N_937,N_99);
nand U1955 (N_1955,N_645,N_216);
and U1956 (N_1956,N_462,N_747);
and U1957 (N_1957,N_87,N_878);
and U1958 (N_1958,N_588,N_198);
and U1959 (N_1959,N_109,N_618);
and U1960 (N_1960,N_967,N_520);
nor U1961 (N_1961,N_391,N_339);
and U1962 (N_1962,N_835,N_868);
nor U1963 (N_1963,N_233,N_921);
and U1964 (N_1964,N_721,N_183);
or U1965 (N_1965,N_661,N_854);
and U1966 (N_1966,N_943,N_787);
nor U1967 (N_1967,N_159,N_278);
and U1968 (N_1968,N_192,N_104);
nor U1969 (N_1969,N_49,N_25);
or U1970 (N_1970,N_492,N_396);
and U1971 (N_1971,N_216,N_846);
nand U1972 (N_1972,N_224,N_146);
nand U1973 (N_1973,N_541,N_195);
xnor U1974 (N_1974,N_538,N_381);
and U1975 (N_1975,N_708,N_179);
and U1976 (N_1976,N_661,N_272);
nor U1977 (N_1977,N_41,N_235);
or U1978 (N_1978,N_265,N_6);
nor U1979 (N_1979,N_590,N_266);
or U1980 (N_1980,N_570,N_870);
or U1981 (N_1981,N_589,N_544);
nor U1982 (N_1982,N_720,N_316);
or U1983 (N_1983,N_243,N_605);
nand U1984 (N_1984,N_486,N_737);
xnor U1985 (N_1985,N_281,N_683);
and U1986 (N_1986,N_280,N_781);
nand U1987 (N_1987,N_554,N_791);
and U1988 (N_1988,N_484,N_956);
and U1989 (N_1989,N_248,N_232);
or U1990 (N_1990,N_508,N_167);
or U1991 (N_1991,N_9,N_297);
and U1992 (N_1992,N_751,N_743);
or U1993 (N_1993,N_962,N_300);
nand U1994 (N_1994,N_434,N_249);
and U1995 (N_1995,N_382,N_391);
nor U1996 (N_1996,N_731,N_694);
nand U1997 (N_1997,N_194,N_433);
or U1998 (N_1998,N_873,N_510);
nand U1999 (N_1999,N_192,N_270);
or U2000 (N_2000,N_1099,N_1056);
nand U2001 (N_2001,N_1304,N_1272);
and U2002 (N_2002,N_1326,N_1197);
or U2003 (N_2003,N_1030,N_1042);
nor U2004 (N_2004,N_1496,N_1307);
nand U2005 (N_2005,N_1605,N_1606);
or U2006 (N_2006,N_1413,N_1624);
nor U2007 (N_2007,N_1767,N_1227);
or U2008 (N_2008,N_1128,N_1271);
nand U2009 (N_2009,N_1064,N_1560);
nand U2010 (N_2010,N_1852,N_1512);
xor U2011 (N_2011,N_1415,N_1266);
nand U2012 (N_2012,N_1650,N_1361);
or U2013 (N_2013,N_1894,N_1747);
or U2014 (N_2014,N_1303,N_1455);
or U2015 (N_2015,N_1832,N_1929);
nor U2016 (N_2016,N_1074,N_1363);
nor U2017 (N_2017,N_1092,N_1398);
nor U2018 (N_2018,N_1598,N_1634);
nor U2019 (N_2019,N_1258,N_1163);
or U2020 (N_2020,N_1773,N_1007);
nand U2021 (N_2021,N_1887,N_1502);
nor U2022 (N_2022,N_1636,N_1527);
or U2023 (N_2023,N_1790,N_1223);
nand U2024 (N_2024,N_1618,N_1426);
and U2025 (N_2025,N_1824,N_1222);
xnor U2026 (N_2026,N_1802,N_1559);
nor U2027 (N_2027,N_1759,N_1620);
and U2028 (N_2028,N_1692,N_1509);
nand U2029 (N_2029,N_1148,N_1242);
and U2030 (N_2030,N_1275,N_1281);
nand U2031 (N_2031,N_1172,N_1943);
nand U2032 (N_2032,N_1269,N_1633);
nor U2033 (N_2033,N_1193,N_1318);
and U2034 (N_2034,N_1651,N_1595);
nor U2035 (N_2035,N_1245,N_1554);
nand U2036 (N_2036,N_1609,N_1553);
xor U2037 (N_2037,N_1126,N_1395);
or U2038 (N_2038,N_1424,N_1623);
and U2039 (N_2039,N_1966,N_1780);
nor U2040 (N_2040,N_1050,N_1334);
or U2041 (N_2041,N_1120,N_1340);
or U2042 (N_2042,N_1836,N_1255);
or U2043 (N_2043,N_1377,N_1231);
nand U2044 (N_2044,N_1571,N_1751);
or U2045 (N_2045,N_1775,N_1820);
nand U2046 (N_2046,N_1762,N_1501);
nor U2047 (N_2047,N_1167,N_1044);
nand U2048 (N_2048,N_1814,N_1290);
nand U2049 (N_2049,N_1719,N_1433);
nor U2050 (N_2050,N_1243,N_1503);
nor U2051 (N_2051,N_1933,N_1582);
or U2052 (N_2052,N_1277,N_1165);
nor U2053 (N_2053,N_1194,N_1524);
nand U2054 (N_2054,N_1815,N_1043);
or U2055 (N_2055,N_1338,N_1722);
nor U2056 (N_2056,N_1001,N_1123);
nand U2057 (N_2057,N_1434,N_1577);
or U2058 (N_2058,N_1990,N_1487);
and U2059 (N_2059,N_1541,N_1694);
nand U2060 (N_2060,N_1071,N_1573);
and U2061 (N_2061,N_1965,N_1195);
nand U2062 (N_2062,N_1584,N_1282);
or U2063 (N_2063,N_1017,N_1339);
and U2064 (N_2064,N_1312,N_1793);
or U2065 (N_2065,N_1689,N_1729);
xnor U2066 (N_2066,N_1508,N_1484);
or U2067 (N_2067,N_1717,N_1350);
and U2068 (N_2068,N_1569,N_1770);
and U2069 (N_2069,N_1886,N_1495);
nor U2070 (N_2070,N_1918,N_1107);
xor U2071 (N_2071,N_1497,N_1839);
or U2072 (N_2072,N_1146,N_1898);
nand U2073 (N_2073,N_1038,N_1109);
nor U2074 (N_2074,N_1853,N_1649);
nor U2075 (N_2075,N_1332,N_1586);
nand U2076 (N_2076,N_1319,N_1536);
nand U2077 (N_2077,N_1488,N_1701);
nand U2078 (N_2078,N_1486,N_1766);
and U2079 (N_2079,N_1593,N_1628);
nor U2080 (N_2080,N_1783,N_1530);
and U2081 (N_2081,N_1670,N_1666);
and U2082 (N_2082,N_1130,N_1441);
nand U2083 (N_2083,N_1024,N_1088);
nor U2084 (N_2084,N_1500,N_1947);
and U2085 (N_2085,N_1678,N_1254);
nand U2086 (N_2086,N_1122,N_1868);
xnor U2087 (N_2087,N_1962,N_1283);
and U2088 (N_2088,N_1768,N_1860);
nor U2089 (N_2089,N_1669,N_1671);
and U2090 (N_2090,N_1925,N_1972);
or U2091 (N_2091,N_1854,N_1199);
or U2092 (N_2092,N_1084,N_1108);
or U2093 (N_2093,N_1520,N_1481);
and U2094 (N_2094,N_1556,N_1543);
or U2095 (N_2095,N_1233,N_1951);
or U2096 (N_2096,N_1238,N_1405);
and U2097 (N_2097,N_1708,N_1732);
nor U2098 (N_2098,N_1629,N_1461);
or U2099 (N_2099,N_1993,N_1330);
nand U2100 (N_2100,N_1058,N_1881);
or U2101 (N_2101,N_1117,N_1012);
nand U2102 (N_2102,N_1858,N_1013);
or U2103 (N_2103,N_1466,N_1869);
nand U2104 (N_2104,N_1119,N_1826);
nand U2105 (N_2105,N_1029,N_1305);
nand U2106 (N_2106,N_1156,N_1346);
and U2107 (N_2107,N_1856,N_1944);
and U2108 (N_2108,N_1257,N_1080);
and U2109 (N_2109,N_1190,N_1412);
or U2110 (N_2110,N_1677,N_1637);
nor U2111 (N_2111,N_1592,N_1958);
and U2112 (N_2112,N_1704,N_1366);
nor U2113 (N_2113,N_1519,N_1955);
nor U2114 (N_2114,N_1796,N_1798);
nor U2115 (N_2115,N_1381,N_1622);
nand U2116 (N_2116,N_1507,N_1781);
and U2117 (N_2117,N_1752,N_1237);
nand U2118 (N_2118,N_1895,N_1081);
and U2119 (N_2119,N_1679,N_1260);
or U2120 (N_2120,N_1136,N_1331);
and U2121 (N_2121,N_1574,N_1535);
and U2122 (N_2122,N_1162,N_1157);
and U2123 (N_2123,N_1110,N_1794);
and U2124 (N_2124,N_1871,N_1511);
nand U2125 (N_2125,N_1475,N_1444);
nand U2126 (N_2126,N_1922,N_1842);
nor U2127 (N_2127,N_1224,N_1268);
or U2128 (N_2128,N_1370,N_1915);
or U2129 (N_2129,N_1063,N_1896);
and U2130 (N_2130,N_1387,N_1207);
nand U2131 (N_2131,N_1600,N_1758);
or U2132 (N_2132,N_1323,N_1037);
and U2133 (N_2133,N_1548,N_1378);
and U2134 (N_2134,N_1129,N_1928);
nor U2135 (N_2135,N_1386,N_1036);
and U2136 (N_2136,N_1923,N_1604);
and U2137 (N_2137,N_1292,N_1220);
xnor U2138 (N_2138,N_1082,N_1362);
nor U2139 (N_2139,N_1427,N_1716);
or U2140 (N_2140,N_1893,N_1125);
or U2141 (N_2141,N_1875,N_1186);
nor U2142 (N_2142,N_1464,N_1799);
nand U2143 (N_2143,N_1632,N_1429);
nor U2144 (N_2144,N_1391,N_1472);
or U2145 (N_2145,N_1919,N_1921);
nor U2146 (N_2146,N_1838,N_1959);
nor U2147 (N_2147,N_1355,N_1336);
or U2148 (N_2148,N_1217,N_1187);
xnor U2149 (N_2149,N_1714,N_1971);
nor U2150 (N_2150,N_1792,N_1211);
nand U2151 (N_2151,N_1137,N_1937);
or U2152 (N_2152,N_1544,N_1698);
and U2153 (N_2153,N_1450,N_1189);
nor U2154 (N_2154,N_1096,N_1251);
xor U2155 (N_2155,N_1969,N_1494);
or U2156 (N_2156,N_1440,N_1451);
or U2157 (N_2157,N_1695,N_1383);
nor U2158 (N_2158,N_1141,N_1968);
or U2159 (N_2159,N_1053,N_1308);
and U2160 (N_2160,N_1754,N_1685);
and U2161 (N_2161,N_1952,N_1542);
nor U2162 (N_2162,N_1483,N_1499);
nand U2163 (N_2163,N_1159,N_1841);
nand U2164 (N_2164,N_1314,N_1745);
and U2165 (N_2165,N_1720,N_1562);
or U2166 (N_2166,N_1003,N_1675);
or U2167 (N_2167,N_1421,N_1811);
nor U2168 (N_2168,N_1528,N_1351);
and U2169 (N_2169,N_1612,N_1996);
and U2170 (N_2170,N_1219,N_1713);
nand U2171 (N_2171,N_1152,N_1899);
and U2172 (N_2172,N_1801,N_1178);
and U2173 (N_2173,N_1347,N_1205);
nor U2174 (N_2174,N_1927,N_1910);
nand U2175 (N_2175,N_1756,N_1552);
and U2176 (N_2176,N_1806,N_1010);
xor U2177 (N_2177,N_1158,N_1791);
or U2178 (N_2178,N_1023,N_1452);
nor U2179 (N_2179,N_1912,N_1170);
nor U2180 (N_2180,N_1179,N_1828);
and U2181 (N_2181,N_1564,N_1845);
and U2182 (N_2182,N_1216,N_1953);
nor U2183 (N_2183,N_1712,N_1660);
nor U2184 (N_2184,N_1069,N_1594);
nor U2185 (N_2185,N_1862,N_1135);
and U2186 (N_2186,N_1437,N_1373);
nand U2187 (N_2187,N_1999,N_1655);
nor U2188 (N_2188,N_1934,N_1550);
nand U2189 (N_2189,N_1786,N_1748);
nand U2190 (N_2190,N_1626,N_1104);
or U2191 (N_2191,N_1196,N_1143);
and U2192 (N_2192,N_1491,N_1880);
nor U2193 (N_2193,N_1705,N_1516);
nand U2194 (N_2194,N_1396,N_1213);
and U2195 (N_2195,N_1394,N_1737);
or U2196 (N_2196,N_1407,N_1435);
nand U2197 (N_2197,N_1776,N_1480);
nor U2198 (N_2198,N_1686,N_1575);
nor U2199 (N_2199,N_1133,N_1454);
nor U2200 (N_2200,N_1973,N_1872);
and U2201 (N_2201,N_1093,N_1324);
nor U2202 (N_2202,N_1161,N_1425);
and U2203 (N_2203,N_1328,N_1981);
nor U2204 (N_2204,N_1335,N_1124);
nor U2205 (N_2205,N_1567,N_1420);
nand U2206 (N_2206,N_1411,N_1585);
or U2207 (N_2207,N_1684,N_1960);
nor U2208 (N_2208,N_1568,N_1975);
or U2209 (N_2209,N_1149,N_1368);
and U2210 (N_2210,N_1371,N_1343);
nand U2211 (N_2211,N_1089,N_1627);
or U2212 (N_2212,N_1359,N_1252);
nor U2213 (N_2213,N_1325,N_1111);
nand U2214 (N_2214,N_1907,N_1565);
and U2215 (N_2215,N_1631,N_1865);
and U2216 (N_2216,N_1457,N_1474);
or U2217 (N_2217,N_1306,N_1376);
nor U2218 (N_2218,N_1635,N_1239);
nand U2219 (N_2219,N_1859,N_1070);
nor U2220 (N_2220,N_1772,N_1293);
nand U2221 (N_2221,N_1734,N_1337);
xor U2222 (N_2222,N_1221,N_1462);
and U2223 (N_2223,N_1068,N_1674);
nand U2224 (N_2224,N_1611,N_1823);
and U2225 (N_2225,N_1344,N_1028);
nor U2226 (N_2226,N_1436,N_1809);
and U2227 (N_2227,N_1103,N_1563);
or U2228 (N_2228,N_1721,N_1816);
and U2229 (N_2229,N_1738,N_1715);
nand U2230 (N_2230,N_1062,N_1288);
nor U2231 (N_2231,N_1296,N_1442);
nand U2232 (N_2232,N_1735,N_1613);
and U2233 (N_2233,N_1225,N_1203);
and U2234 (N_2234,N_1778,N_1743);
or U2235 (N_2235,N_1446,N_1757);
or U2236 (N_2236,N_1286,N_1358);
nor U2237 (N_2237,N_1803,N_1939);
or U2238 (N_2238,N_1579,N_1982);
nand U2239 (N_2239,N_1279,N_1739);
nor U2240 (N_2240,N_1206,N_1289);
nand U2241 (N_2241,N_1904,N_1805);
or U2242 (N_2242,N_1078,N_1460);
nor U2243 (N_2243,N_1406,N_1764);
nand U2244 (N_2244,N_1182,N_1851);
and U2245 (N_2245,N_1936,N_1278);
and U2246 (N_2246,N_1097,N_1986);
or U2247 (N_2247,N_1645,N_1587);
nor U2248 (N_2248,N_1341,N_1322);
and U2249 (N_2249,N_1646,N_1850);
and U2250 (N_2250,N_1664,N_1883);
and U2251 (N_2251,N_1547,N_1034);
nand U2252 (N_2252,N_1945,N_1882);
nor U2253 (N_2253,N_1769,N_1040);
nand U2254 (N_2254,N_1234,N_1009);
and U2255 (N_2255,N_1049,N_1202);
nor U2256 (N_2256,N_1513,N_1169);
nor U2257 (N_2257,N_1212,N_1490);
nand U2258 (N_2258,N_1113,N_1379);
nand U2259 (N_2259,N_1987,N_1320);
nand U2260 (N_2260,N_1285,N_1215);
nand U2261 (N_2261,N_1984,N_1310);
or U2262 (N_2262,N_1035,N_1132);
and U2263 (N_2263,N_1526,N_1948);
and U2264 (N_2264,N_1913,N_1834);
and U2265 (N_2265,N_1537,N_1821);
nor U2266 (N_2266,N_1602,N_1911);
nand U2267 (N_2267,N_1517,N_1329);
and U2268 (N_2268,N_1116,N_1192);
nor U2269 (N_2269,N_1866,N_1848);
nor U2270 (N_2270,N_1558,N_1901);
or U2271 (N_2271,N_1808,N_1638);
and U2272 (N_2272,N_1997,N_1438);
or U2273 (N_2273,N_1284,N_1549);
and U2274 (N_2274,N_1625,N_1864);
nor U2275 (N_2275,N_1015,N_1797);
nand U2276 (N_2276,N_1188,N_1873);
and U2277 (N_2277,N_1085,N_1051);
and U2278 (N_2278,N_1014,N_1094);
nor U2279 (N_2279,N_1505,N_1138);
nor U2280 (N_2280,N_1447,N_1348);
xnor U2281 (N_2281,N_1967,N_1707);
nor U2282 (N_2282,N_1905,N_1617);
nand U2283 (N_2283,N_1448,N_1291);
nor U2284 (N_2284,N_1788,N_1090);
or U2285 (N_2285,N_1531,N_1970);
or U2286 (N_2286,N_1261,N_1800);
nor U2287 (N_2287,N_1065,N_1771);
nand U2288 (N_2288,N_1367,N_1393);
and U2289 (N_2289,N_1557,N_1259);
and U2290 (N_2290,N_1777,N_1054);
nor U2291 (N_2291,N_1833,N_1048);
and U2292 (N_2292,N_1957,N_1214);
or U2293 (N_2293,N_1870,N_1353);
or U2294 (N_2294,N_1736,N_1687);
and U2295 (N_2295,N_1027,N_1249);
or U2296 (N_2296,N_1682,N_1693);
nor U2297 (N_2297,N_1401,N_1198);
xor U2298 (N_2298,N_1144,N_1356);
or U2299 (N_2299,N_1004,N_1404);
nand U2300 (N_2300,N_1256,N_1931);
or U2301 (N_2301,N_1112,N_1031);
and U2302 (N_2302,N_1264,N_1384);
nor U2303 (N_2303,N_1818,N_1647);
and U2304 (N_2304,N_1658,N_1016);
nand U2305 (N_2305,N_1963,N_1827);
and U2306 (N_2306,N_1232,N_1661);
and U2307 (N_2307,N_1599,N_1208);
or U2308 (N_2308,N_1057,N_1978);
or U2309 (N_2309,N_1855,N_1020);
nand U2310 (N_2310,N_1974,N_1956);
or U2311 (N_2311,N_1603,N_1164);
or U2312 (N_2312,N_1300,N_1134);
nor U2313 (N_2313,N_1498,N_1066);
nand U2314 (N_2314,N_1008,N_1696);
nor U2315 (N_2315,N_1608,N_1876);
nor U2316 (N_2316,N_1374,N_1482);
or U2317 (N_2317,N_1861,N_1656);
nor U2318 (N_2318,N_1744,N_1313);
nand U2319 (N_2319,N_1155,N_1139);
or U2320 (N_2320,N_1465,N_1153);
xor U2321 (N_2321,N_1410,N_1891);
xor U2322 (N_2322,N_1473,N_1654);
or U2323 (N_2323,N_1201,N_1725);
nand U2324 (N_2324,N_1443,N_1240);
and U2325 (N_2325,N_1640,N_1000);
xnor U2326 (N_2326,N_1075,N_1022);
nand U2327 (N_2327,N_1857,N_1403);
and U2328 (N_2328,N_1697,N_1485);
or U2329 (N_2329,N_1884,N_1619);
nor U2330 (N_2330,N_1659,N_1414);
nand U2331 (N_2331,N_1690,N_1382);
or U2332 (N_2332,N_1785,N_1700);
and U2333 (N_2333,N_1807,N_1241);
nor U2334 (N_2334,N_1601,N_1392);
or U2335 (N_2335,N_1365,N_1369);
nor U2336 (N_2336,N_1301,N_1115);
or U2337 (N_2337,N_1273,N_1514);
and U2338 (N_2338,N_1428,N_1668);
or U2339 (N_2339,N_1317,N_1349);
nand U2340 (N_2340,N_1311,N_1964);
nor U2341 (N_2341,N_1262,N_1749);
nand U2342 (N_2342,N_1810,N_1295);
nor U2343 (N_2343,N_1127,N_1784);
nor U2344 (N_2344,N_1087,N_1765);
and U2345 (N_2345,N_1309,N_1354);
and U2346 (N_2346,N_1315,N_1449);
and U2347 (N_2347,N_1072,N_1782);
nand U2348 (N_2348,N_1648,N_1538);
and U2349 (N_2349,N_1372,N_1529);
nor U2350 (N_2350,N_1218,N_1045);
nand U2351 (N_2351,N_1662,N_1253);
nand U2352 (N_2352,N_1812,N_1879);
and U2353 (N_2353,N_1900,N_1246);
nand U2354 (N_2354,N_1375,N_1002);
or U2355 (N_2355,N_1493,N_1706);
nand U2356 (N_2356,N_1703,N_1710);
nor U2357 (N_2357,N_1525,N_1546);
or U2358 (N_2358,N_1950,N_1431);
nor U2359 (N_2359,N_1731,N_1941);
nand U2360 (N_2360,N_1863,N_1006);
or U2361 (N_2361,N_1025,N_1930);
or U2362 (N_2362,N_1813,N_1106);
or U2363 (N_2363,N_1247,N_1641);
or U2364 (N_2364,N_1357,N_1327);
and U2365 (N_2365,N_1229,N_1991);
or U2366 (N_2366,N_1479,N_1418);
and U2367 (N_2367,N_1924,N_1095);
or U2368 (N_2368,N_1630,N_1976);
nor U2369 (N_2369,N_1607,N_1977);
nand U2370 (N_2370,N_1100,N_1299);
and U2371 (N_2371,N_1297,N_1011);
or U2372 (N_2372,N_1615,N_1302);
or U2373 (N_2373,N_1091,N_1908);
nand U2374 (N_2374,N_1998,N_1992);
nand U2375 (N_2375,N_1470,N_1345);
nor U2376 (N_2376,N_1079,N_1683);
nand U2377 (N_2377,N_1985,N_1021);
nand U2378 (N_2378,N_1760,N_1055);
and U2379 (N_2379,N_1702,N_1168);
nand U2380 (N_2380,N_1026,N_1102);
nand U2381 (N_2381,N_1018,N_1105);
or U2382 (N_2382,N_1995,N_1580);
or U2383 (N_2383,N_1166,N_1204);
and U2384 (N_2384,N_1920,N_1724);
or U2385 (N_2385,N_1667,N_1763);
nand U2386 (N_2386,N_1572,N_1545);
nand U2387 (N_2387,N_1316,N_1831);
nand U2388 (N_2388,N_1360,N_1774);
nand U2389 (N_2389,N_1954,N_1114);
xor U2390 (N_2390,N_1730,N_1847);
or U2391 (N_2391,N_1175,N_1267);
or U2392 (N_2392,N_1742,N_1039);
and U2393 (N_2393,N_1076,N_1566);
or U2394 (N_2394,N_1523,N_1352);
or U2395 (N_2395,N_1422,N_1610);
nand U2396 (N_2396,N_1576,N_1263);
nor U2397 (N_2397,N_1949,N_1423);
and U2398 (N_2398,N_1902,N_1333);
and U2399 (N_2399,N_1644,N_1621);
and U2400 (N_2400,N_1210,N_1476);
nand U2401 (N_2401,N_1532,N_1101);
and U2402 (N_2402,N_1614,N_1728);
nor U2403 (N_2403,N_1581,N_1469);
nor U2404 (N_2404,N_1226,N_1878);
and U2405 (N_2405,N_1150,N_1019);
nand U2406 (N_2406,N_1699,N_1463);
and U2407 (N_2407,N_1843,N_1276);
nand U2408 (N_2408,N_1830,N_1551);
nand U2409 (N_2409,N_1154,N_1657);
xor U2410 (N_2410,N_1840,N_1534);
nor U2411 (N_2411,N_1709,N_1032);
and U2412 (N_2412,N_1399,N_1181);
nand U2413 (N_2413,N_1061,N_1672);
or U2414 (N_2414,N_1746,N_1183);
or U2415 (N_2415,N_1979,N_1244);
nand U2416 (N_2416,N_1121,N_1439);
nor U2417 (N_2417,N_1942,N_1118);
or U2418 (N_2418,N_1589,N_1098);
nor U2419 (N_2419,N_1673,N_1835);
or U2420 (N_2420,N_1209,N_1515);
and U2421 (N_2421,N_1280,N_1230);
or U2422 (N_2422,N_1639,N_1946);
and U2423 (N_2423,N_1726,N_1147);
or U2424 (N_2424,N_1380,N_1753);
nand U2425 (N_2425,N_1321,N_1789);
and U2426 (N_2426,N_1665,N_1177);
and U2427 (N_2427,N_1073,N_1596);
nand U2428 (N_2428,N_1077,N_1236);
and U2429 (N_2429,N_1409,N_1795);
or U2430 (N_2430,N_1888,N_1539);
or U2431 (N_2431,N_1926,N_1779);
nand U2432 (N_2432,N_1265,N_1510);
nand U2433 (N_2433,N_1397,N_1897);
or U2434 (N_2434,N_1733,N_1588);
nor U2435 (N_2435,N_1390,N_1142);
or U2436 (N_2436,N_1846,N_1471);
nand U2437 (N_2437,N_1468,N_1235);
or U2438 (N_2438,N_1890,N_1173);
nand U2439 (N_2439,N_1822,N_1046);
and U2440 (N_2440,N_1445,N_1385);
nor U2441 (N_2441,N_1578,N_1829);
nand U2442 (N_2442,N_1453,N_1432);
nand U2443 (N_2443,N_1583,N_1458);
or U2444 (N_2444,N_1430,N_1653);
nor U2445 (N_2445,N_1663,N_1691);
nand U2446 (N_2446,N_1989,N_1533);
nor U2447 (N_2447,N_1518,N_1591);
or U2448 (N_2448,N_1506,N_1867);
nand U2449 (N_2449,N_1988,N_1849);
nor U2450 (N_2450,N_1711,N_1688);
nand U2451 (N_2451,N_1740,N_1961);
and U2452 (N_2452,N_1342,N_1804);
nor U2453 (N_2453,N_1643,N_1909);
or U2454 (N_2454,N_1086,N_1844);
or U2455 (N_2455,N_1914,N_1892);
and U2456 (N_2456,N_1298,N_1994);
and U2457 (N_2457,N_1492,N_1417);
nand U2458 (N_2458,N_1478,N_1185);
or U2459 (N_2459,N_1932,N_1228);
nor U2460 (N_2460,N_1459,N_1787);
nor U2461 (N_2461,N_1642,N_1145);
nand U2462 (N_2462,N_1889,N_1151);
nor U2463 (N_2463,N_1248,N_1817);
and U2464 (N_2464,N_1176,N_1489);
or U2465 (N_2465,N_1060,N_1819);
nor U2466 (N_2466,N_1597,N_1067);
or U2467 (N_2467,N_1083,N_1676);
nor U2468 (N_2468,N_1184,N_1400);
and U2469 (N_2469,N_1041,N_1416);
or U2470 (N_2470,N_1561,N_1274);
or U2471 (N_2471,N_1364,N_1590);
nand U2472 (N_2472,N_1456,N_1504);
nor U2473 (N_2473,N_1033,N_1467);
nand U2474 (N_2474,N_1916,N_1200);
nor U2475 (N_2475,N_1877,N_1761);
nor U2476 (N_2476,N_1825,N_1741);
or U2477 (N_2477,N_1906,N_1723);
or U2478 (N_2478,N_1837,N_1059);
nand U2479 (N_2479,N_1652,N_1755);
nand U2480 (N_2480,N_1160,N_1938);
xor U2481 (N_2481,N_1191,N_1408);
or U2482 (N_2482,N_1570,N_1521);
nand U2483 (N_2483,N_1171,N_1287);
nor U2484 (N_2484,N_1917,N_1616);
and U2485 (N_2485,N_1980,N_1983);
nor U2486 (N_2486,N_1388,N_1935);
and U2487 (N_2487,N_1180,N_1522);
and U2488 (N_2488,N_1140,N_1540);
or U2489 (N_2489,N_1389,N_1005);
and U2490 (N_2490,N_1750,N_1681);
or U2491 (N_2491,N_1270,N_1131);
or U2492 (N_2492,N_1727,N_1874);
nand U2493 (N_2493,N_1402,N_1885);
nor U2494 (N_2494,N_1052,N_1555);
nand U2495 (N_2495,N_1419,N_1718);
or U2496 (N_2496,N_1903,N_1477);
nor U2497 (N_2497,N_1940,N_1047);
nor U2498 (N_2498,N_1174,N_1294);
nand U2499 (N_2499,N_1250,N_1680);
or U2500 (N_2500,N_1586,N_1090);
nor U2501 (N_2501,N_1580,N_1292);
and U2502 (N_2502,N_1082,N_1269);
and U2503 (N_2503,N_1751,N_1145);
or U2504 (N_2504,N_1546,N_1570);
nand U2505 (N_2505,N_1439,N_1244);
or U2506 (N_2506,N_1019,N_1239);
xnor U2507 (N_2507,N_1179,N_1076);
and U2508 (N_2508,N_1457,N_1098);
and U2509 (N_2509,N_1867,N_1591);
xor U2510 (N_2510,N_1247,N_1882);
and U2511 (N_2511,N_1641,N_1659);
nand U2512 (N_2512,N_1270,N_1592);
nand U2513 (N_2513,N_1198,N_1846);
nor U2514 (N_2514,N_1947,N_1087);
nor U2515 (N_2515,N_1656,N_1766);
nor U2516 (N_2516,N_1522,N_1307);
or U2517 (N_2517,N_1678,N_1284);
nand U2518 (N_2518,N_1089,N_1872);
nand U2519 (N_2519,N_1929,N_1659);
and U2520 (N_2520,N_1453,N_1065);
xor U2521 (N_2521,N_1282,N_1927);
nor U2522 (N_2522,N_1446,N_1050);
or U2523 (N_2523,N_1632,N_1543);
nor U2524 (N_2524,N_1485,N_1959);
or U2525 (N_2525,N_1722,N_1478);
or U2526 (N_2526,N_1960,N_1396);
and U2527 (N_2527,N_1924,N_1431);
nor U2528 (N_2528,N_1566,N_1714);
or U2529 (N_2529,N_1796,N_1327);
nand U2530 (N_2530,N_1726,N_1795);
nand U2531 (N_2531,N_1644,N_1652);
nand U2532 (N_2532,N_1036,N_1666);
nand U2533 (N_2533,N_1339,N_1735);
or U2534 (N_2534,N_1676,N_1274);
and U2535 (N_2535,N_1386,N_1057);
nand U2536 (N_2536,N_1632,N_1071);
and U2537 (N_2537,N_1877,N_1116);
nand U2538 (N_2538,N_1076,N_1845);
nor U2539 (N_2539,N_1270,N_1048);
and U2540 (N_2540,N_1810,N_1093);
nand U2541 (N_2541,N_1458,N_1004);
and U2542 (N_2542,N_1834,N_1381);
nand U2543 (N_2543,N_1948,N_1625);
nor U2544 (N_2544,N_1829,N_1106);
or U2545 (N_2545,N_1004,N_1429);
nand U2546 (N_2546,N_1927,N_1977);
and U2547 (N_2547,N_1768,N_1433);
nor U2548 (N_2548,N_1986,N_1323);
or U2549 (N_2549,N_1492,N_1077);
nor U2550 (N_2550,N_1191,N_1337);
and U2551 (N_2551,N_1329,N_1701);
nand U2552 (N_2552,N_1904,N_1479);
nor U2553 (N_2553,N_1727,N_1447);
nand U2554 (N_2554,N_1973,N_1763);
nand U2555 (N_2555,N_1786,N_1069);
and U2556 (N_2556,N_1870,N_1942);
nand U2557 (N_2557,N_1687,N_1894);
and U2558 (N_2558,N_1533,N_1130);
and U2559 (N_2559,N_1789,N_1531);
nand U2560 (N_2560,N_1059,N_1371);
nor U2561 (N_2561,N_1961,N_1959);
or U2562 (N_2562,N_1605,N_1705);
nand U2563 (N_2563,N_1819,N_1269);
nand U2564 (N_2564,N_1339,N_1578);
nor U2565 (N_2565,N_1203,N_1290);
and U2566 (N_2566,N_1481,N_1792);
and U2567 (N_2567,N_1514,N_1175);
or U2568 (N_2568,N_1171,N_1533);
and U2569 (N_2569,N_1962,N_1138);
nor U2570 (N_2570,N_1872,N_1155);
nor U2571 (N_2571,N_1057,N_1418);
or U2572 (N_2572,N_1110,N_1901);
nand U2573 (N_2573,N_1924,N_1846);
nor U2574 (N_2574,N_1252,N_1221);
or U2575 (N_2575,N_1192,N_1813);
xor U2576 (N_2576,N_1805,N_1750);
or U2577 (N_2577,N_1528,N_1525);
nand U2578 (N_2578,N_1048,N_1512);
and U2579 (N_2579,N_1610,N_1012);
or U2580 (N_2580,N_1027,N_1368);
or U2581 (N_2581,N_1079,N_1988);
nand U2582 (N_2582,N_1487,N_1539);
and U2583 (N_2583,N_1898,N_1607);
nor U2584 (N_2584,N_1386,N_1884);
nand U2585 (N_2585,N_1909,N_1608);
nand U2586 (N_2586,N_1913,N_1212);
and U2587 (N_2587,N_1310,N_1750);
or U2588 (N_2588,N_1793,N_1380);
or U2589 (N_2589,N_1247,N_1710);
xnor U2590 (N_2590,N_1687,N_1997);
nor U2591 (N_2591,N_1347,N_1187);
nand U2592 (N_2592,N_1514,N_1305);
or U2593 (N_2593,N_1597,N_1283);
nand U2594 (N_2594,N_1168,N_1018);
and U2595 (N_2595,N_1006,N_1477);
and U2596 (N_2596,N_1291,N_1014);
nor U2597 (N_2597,N_1387,N_1086);
nand U2598 (N_2598,N_1109,N_1759);
or U2599 (N_2599,N_1942,N_1147);
or U2600 (N_2600,N_1103,N_1048);
nand U2601 (N_2601,N_1619,N_1400);
nand U2602 (N_2602,N_1438,N_1690);
nor U2603 (N_2603,N_1054,N_1240);
nor U2604 (N_2604,N_1878,N_1484);
or U2605 (N_2605,N_1537,N_1884);
and U2606 (N_2606,N_1258,N_1814);
nor U2607 (N_2607,N_1208,N_1771);
nor U2608 (N_2608,N_1924,N_1655);
or U2609 (N_2609,N_1059,N_1439);
or U2610 (N_2610,N_1689,N_1117);
and U2611 (N_2611,N_1284,N_1992);
nor U2612 (N_2612,N_1229,N_1576);
and U2613 (N_2613,N_1677,N_1789);
nand U2614 (N_2614,N_1599,N_1568);
nand U2615 (N_2615,N_1372,N_1205);
and U2616 (N_2616,N_1686,N_1129);
or U2617 (N_2617,N_1366,N_1637);
nand U2618 (N_2618,N_1539,N_1520);
nand U2619 (N_2619,N_1590,N_1645);
and U2620 (N_2620,N_1937,N_1243);
or U2621 (N_2621,N_1471,N_1056);
nor U2622 (N_2622,N_1623,N_1317);
nor U2623 (N_2623,N_1448,N_1407);
nor U2624 (N_2624,N_1284,N_1115);
nand U2625 (N_2625,N_1421,N_1290);
and U2626 (N_2626,N_1270,N_1993);
or U2627 (N_2627,N_1914,N_1690);
xor U2628 (N_2628,N_1782,N_1022);
nor U2629 (N_2629,N_1158,N_1969);
nor U2630 (N_2630,N_1951,N_1005);
and U2631 (N_2631,N_1474,N_1399);
nand U2632 (N_2632,N_1241,N_1527);
nand U2633 (N_2633,N_1157,N_1441);
or U2634 (N_2634,N_1049,N_1488);
nor U2635 (N_2635,N_1019,N_1931);
and U2636 (N_2636,N_1518,N_1471);
and U2637 (N_2637,N_1880,N_1150);
xor U2638 (N_2638,N_1148,N_1136);
nor U2639 (N_2639,N_1719,N_1503);
nand U2640 (N_2640,N_1632,N_1337);
nand U2641 (N_2641,N_1774,N_1104);
and U2642 (N_2642,N_1588,N_1963);
and U2643 (N_2643,N_1033,N_1040);
and U2644 (N_2644,N_1427,N_1027);
nand U2645 (N_2645,N_1573,N_1615);
xnor U2646 (N_2646,N_1118,N_1896);
and U2647 (N_2647,N_1233,N_1848);
nand U2648 (N_2648,N_1811,N_1173);
nor U2649 (N_2649,N_1797,N_1396);
and U2650 (N_2650,N_1484,N_1456);
or U2651 (N_2651,N_1822,N_1079);
xor U2652 (N_2652,N_1137,N_1666);
nand U2653 (N_2653,N_1853,N_1029);
nor U2654 (N_2654,N_1248,N_1390);
nand U2655 (N_2655,N_1788,N_1449);
nor U2656 (N_2656,N_1002,N_1119);
and U2657 (N_2657,N_1211,N_1788);
or U2658 (N_2658,N_1594,N_1370);
nor U2659 (N_2659,N_1902,N_1206);
nor U2660 (N_2660,N_1412,N_1448);
nand U2661 (N_2661,N_1475,N_1726);
nor U2662 (N_2662,N_1874,N_1597);
or U2663 (N_2663,N_1816,N_1800);
or U2664 (N_2664,N_1906,N_1542);
or U2665 (N_2665,N_1161,N_1318);
and U2666 (N_2666,N_1642,N_1771);
xor U2667 (N_2667,N_1788,N_1060);
nor U2668 (N_2668,N_1313,N_1412);
nor U2669 (N_2669,N_1158,N_1819);
and U2670 (N_2670,N_1964,N_1479);
or U2671 (N_2671,N_1120,N_1776);
nand U2672 (N_2672,N_1576,N_1677);
and U2673 (N_2673,N_1700,N_1006);
nand U2674 (N_2674,N_1754,N_1484);
nand U2675 (N_2675,N_1710,N_1585);
nand U2676 (N_2676,N_1225,N_1924);
nor U2677 (N_2677,N_1619,N_1447);
nor U2678 (N_2678,N_1785,N_1169);
or U2679 (N_2679,N_1254,N_1714);
or U2680 (N_2680,N_1645,N_1263);
nor U2681 (N_2681,N_1543,N_1343);
or U2682 (N_2682,N_1844,N_1361);
or U2683 (N_2683,N_1602,N_1819);
or U2684 (N_2684,N_1862,N_1767);
nand U2685 (N_2685,N_1234,N_1502);
nor U2686 (N_2686,N_1116,N_1939);
or U2687 (N_2687,N_1432,N_1776);
nor U2688 (N_2688,N_1481,N_1848);
nand U2689 (N_2689,N_1239,N_1066);
nand U2690 (N_2690,N_1076,N_1190);
nor U2691 (N_2691,N_1052,N_1774);
nor U2692 (N_2692,N_1086,N_1629);
xnor U2693 (N_2693,N_1869,N_1341);
nor U2694 (N_2694,N_1540,N_1119);
and U2695 (N_2695,N_1904,N_1218);
or U2696 (N_2696,N_1391,N_1695);
nor U2697 (N_2697,N_1642,N_1019);
nand U2698 (N_2698,N_1746,N_1269);
nor U2699 (N_2699,N_1887,N_1823);
or U2700 (N_2700,N_1725,N_1052);
and U2701 (N_2701,N_1253,N_1503);
and U2702 (N_2702,N_1211,N_1899);
nor U2703 (N_2703,N_1007,N_1610);
nor U2704 (N_2704,N_1784,N_1034);
nor U2705 (N_2705,N_1279,N_1779);
or U2706 (N_2706,N_1368,N_1253);
nand U2707 (N_2707,N_1100,N_1721);
and U2708 (N_2708,N_1660,N_1064);
or U2709 (N_2709,N_1077,N_1508);
nor U2710 (N_2710,N_1505,N_1681);
nand U2711 (N_2711,N_1935,N_1129);
nand U2712 (N_2712,N_1483,N_1758);
nor U2713 (N_2713,N_1285,N_1661);
nand U2714 (N_2714,N_1891,N_1659);
nand U2715 (N_2715,N_1375,N_1766);
and U2716 (N_2716,N_1742,N_1170);
or U2717 (N_2717,N_1079,N_1339);
nor U2718 (N_2718,N_1356,N_1540);
nor U2719 (N_2719,N_1338,N_1033);
or U2720 (N_2720,N_1704,N_1682);
nand U2721 (N_2721,N_1023,N_1746);
and U2722 (N_2722,N_1503,N_1394);
nand U2723 (N_2723,N_1133,N_1028);
or U2724 (N_2724,N_1400,N_1254);
and U2725 (N_2725,N_1643,N_1980);
or U2726 (N_2726,N_1573,N_1389);
nand U2727 (N_2727,N_1354,N_1628);
xor U2728 (N_2728,N_1858,N_1632);
nor U2729 (N_2729,N_1382,N_1412);
nor U2730 (N_2730,N_1471,N_1465);
and U2731 (N_2731,N_1710,N_1674);
and U2732 (N_2732,N_1900,N_1082);
nor U2733 (N_2733,N_1284,N_1065);
nand U2734 (N_2734,N_1656,N_1852);
nor U2735 (N_2735,N_1840,N_1495);
nand U2736 (N_2736,N_1494,N_1424);
nand U2737 (N_2737,N_1883,N_1054);
or U2738 (N_2738,N_1076,N_1871);
nand U2739 (N_2739,N_1204,N_1716);
and U2740 (N_2740,N_1185,N_1798);
or U2741 (N_2741,N_1937,N_1107);
or U2742 (N_2742,N_1373,N_1625);
nand U2743 (N_2743,N_1799,N_1621);
or U2744 (N_2744,N_1268,N_1000);
or U2745 (N_2745,N_1873,N_1248);
nor U2746 (N_2746,N_1930,N_1262);
nor U2747 (N_2747,N_1698,N_1183);
nand U2748 (N_2748,N_1142,N_1955);
and U2749 (N_2749,N_1480,N_1933);
or U2750 (N_2750,N_1310,N_1634);
and U2751 (N_2751,N_1951,N_1839);
nor U2752 (N_2752,N_1908,N_1098);
nand U2753 (N_2753,N_1706,N_1060);
or U2754 (N_2754,N_1092,N_1762);
nand U2755 (N_2755,N_1078,N_1770);
nand U2756 (N_2756,N_1945,N_1013);
or U2757 (N_2757,N_1136,N_1930);
nand U2758 (N_2758,N_1098,N_1066);
nand U2759 (N_2759,N_1497,N_1029);
nand U2760 (N_2760,N_1409,N_1353);
or U2761 (N_2761,N_1680,N_1451);
nor U2762 (N_2762,N_1600,N_1128);
and U2763 (N_2763,N_1966,N_1984);
and U2764 (N_2764,N_1997,N_1196);
nor U2765 (N_2765,N_1935,N_1957);
nor U2766 (N_2766,N_1887,N_1531);
nand U2767 (N_2767,N_1109,N_1410);
and U2768 (N_2768,N_1276,N_1825);
nor U2769 (N_2769,N_1837,N_1760);
nor U2770 (N_2770,N_1976,N_1049);
nand U2771 (N_2771,N_1016,N_1099);
and U2772 (N_2772,N_1689,N_1781);
or U2773 (N_2773,N_1481,N_1661);
and U2774 (N_2774,N_1912,N_1459);
and U2775 (N_2775,N_1832,N_1797);
or U2776 (N_2776,N_1673,N_1146);
and U2777 (N_2777,N_1792,N_1724);
and U2778 (N_2778,N_1364,N_1013);
nor U2779 (N_2779,N_1840,N_1439);
and U2780 (N_2780,N_1309,N_1740);
or U2781 (N_2781,N_1282,N_1013);
or U2782 (N_2782,N_1987,N_1344);
nor U2783 (N_2783,N_1025,N_1978);
nor U2784 (N_2784,N_1975,N_1062);
nand U2785 (N_2785,N_1041,N_1252);
and U2786 (N_2786,N_1208,N_1443);
xor U2787 (N_2787,N_1377,N_1303);
and U2788 (N_2788,N_1679,N_1401);
nand U2789 (N_2789,N_1706,N_1786);
nor U2790 (N_2790,N_1164,N_1340);
and U2791 (N_2791,N_1469,N_1018);
and U2792 (N_2792,N_1694,N_1127);
and U2793 (N_2793,N_1310,N_1269);
nand U2794 (N_2794,N_1979,N_1709);
nor U2795 (N_2795,N_1490,N_1600);
nand U2796 (N_2796,N_1538,N_1564);
nand U2797 (N_2797,N_1907,N_1258);
and U2798 (N_2798,N_1747,N_1791);
and U2799 (N_2799,N_1188,N_1112);
nand U2800 (N_2800,N_1916,N_1400);
xor U2801 (N_2801,N_1810,N_1559);
nor U2802 (N_2802,N_1896,N_1512);
or U2803 (N_2803,N_1883,N_1200);
nor U2804 (N_2804,N_1851,N_1823);
nand U2805 (N_2805,N_1814,N_1891);
nor U2806 (N_2806,N_1881,N_1414);
or U2807 (N_2807,N_1395,N_1994);
or U2808 (N_2808,N_1953,N_1210);
nor U2809 (N_2809,N_1207,N_1962);
or U2810 (N_2810,N_1385,N_1500);
or U2811 (N_2811,N_1362,N_1284);
nand U2812 (N_2812,N_1118,N_1156);
nand U2813 (N_2813,N_1705,N_1894);
or U2814 (N_2814,N_1854,N_1455);
nand U2815 (N_2815,N_1093,N_1194);
nor U2816 (N_2816,N_1805,N_1199);
nand U2817 (N_2817,N_1629,N_1647);
or U2818 (N_2818,N_1652,N_1370);
nor U2819 (N_2819,N_1417,N_1536);
nor U2820 (N_2820,N_1519,N_1822);
or U2821 (N_2821,N_1169,N_1611);
and U2822 (N_2822,N_1075,N_1057);
and U2823 (N_2823,N_1878,N_1651);
and U2824 (N_2824,N_1550,N_1389);
or U2825 (N_2825,N_1137,N_1978);
xnor U2826 (N_2826,N_1966,N_1792);
nand U2827 (N_2827,N_1555,N_1190);
nor U2828 (N_2828,N_1532,N_1034);
nor U2829 (N_2829,N_1822,N_1983);
nor U2830 (N_2830,N_1886,N_1210);
or U2831 (N_2831,N_1515,N_1706);
nor U2832 (N_2832,N_1052,N_1116);
or U2833 (N_2833,N_1345,N_1660);
and U2834 (N_2834,N_1145,N_1161);
nor U2835 (N_2835,N_1094,N_1917);
and U2836 (N_2836,N_1431,N_1929);
or U2837 (N_2837,N_1845,N_1656);
nand U2838 (N_2838,N_1127,N_1178);
nor U2839 (N_2839,N_1516,N_1444);
xnor U2840 (N_2840,N_1276,N_1034);
or U2841 (N_2841,N_1765,N_1815);
nand U2842 (N_2842,N_1826,N_1800);
nand U2843 (N_2843,N_1036,N_1024);
or U2844 (N_2844,N_1930,N_1420);
and U2845 (N_2845,N_1837,N_1621);
and U2846 (N_2846,N_1067,N_1519);
nand U2847 (N_2847,N_1951,N_1076);
and U2848 (N_2848,N_1663,N_1799);
and U2849 (N_2849,N_1316,N_1043);
and U2850 (N_2850,N_1395,N_1225);
xor U2851 (N_2851,N_1855,N_1958);
nor U2852 (N_2852,N_1845,N_1954);
and U2853 (N_2853,N_1818,N_1671);
nor U2854 (N_2854,N_1106,N_1606);
or U2855 (N_2855,N_1776,N_1858);
and U2856 (N_2856,N_1969,N_1544);
or U2857 (N_2857,N_1718,N_1301);
and U2858 (N_2858,N_1653,N_1672);
nor U2859 (N_2859,N_1883,N_1634);
or U2860 (N_2860,N_1082,N_1958);
or U2861 (N_2861,N_1369,N_1727);
nor U2862 (N_2862,N_1775,N_1519);
and U2863 (N_2863,N_1367,N_1303);
and U2864 (N_2864,N_1383,N_1209);
and U2865 (N_2865,N_1247,N_1307);
and U2866 (N_2866,N_1061,N_1607);
nor U2867 (N_2867,N_1925,N_1747);
nor U2868 (N_2868,N_1150,N_1836);
and U2869 (N_2869,N_1301,N_1314);
or U2870 (N_2870,N_1669,N_1705);
xor U2871 (N_2871,N_1168,N_1745);
nor U2872 (N_2872,N_1731,N_1342);
nand U2873 (N_2873,N_1721,N_1195);
and U2874 (N_2874,N_1859,N_1700);
or U2875 (N_2875,N_1156,N_1418);
nand U2876 (N_2876,N_1561,N_1739);
nor U2877 (N_2877,N_1923,N_1046);
and U2878 (N_2878,N_1020,N_1806);
and U2879 (N_2879,N_1814,N_1103);
and U2880 (N_2880,N_1829,N_1534);
or U2881 (N_2881,N_1767,N_1068);
and U2882 (N_2882,N_1782,N_1999);
nor U2883 (N_2883,N_1743,N_1663);
nand U2884 (N_2884,N_1488,N_1089);
and U2885 (N_2885,N_1587,N_1029);
and U2886 (N_2886,N_1958,N_1807);
nor U2887 (N_2887,N_1056,N_1549);
nand U2888 (N_2888,N_1713,N_1752);
and U2889 (N_2889,N_1011,N_1024);
or U2890 (N_2890,N_1317,N_1499);
nand U2891 (N_2891,N_1967,N_1889);
and U2892 (N_2892,N_1724,N_1819);
nand U2893 (N_2893,N_1856,N_1357);
and U2894 (N_2894,N_1882,N_1215);
or U2895 (N_2895,N_1252,N_1681);
and U2896 (N_2896,N_1694,N_1848);
nand U2897 (N_2897,N_1672,N_1639);
and U2898 (N_2898,N_1748,N_1869);
nor U2899 (N_2899,N_1232,N_1211);
and U2900 (N_2900,N_1035,N_1009);
nand U2901 (N_2901,N_1246,N_1262);
or U2902 (N_2902,N_1484,N_1924);
nor U2903 (N_2903,N_1477,N_1221);
and U2904 (N_2904,N_1109,N_1533);
and U2905 (N_2905,N_1385,N_1788);
nand U2906 (N_2906,N_1174,N_1090);
or U2907 (N_2907,N_1204,N_1042);
nand U2908 (N_2908,N_1117,N_1873);
nand U2909 (N_2909,N_1972,N_1545);
xnor U2910 (N_2910,N_1192,N_1005);
or U2911 (N_2911,N_1492,N_1463);
nand U2912 (N_2912,N_1364,N_1454);
nand U2913 (N_2913,N_1358,N_1245);
or U2914 (N_2914,N_1444,N_1024);
nor U2915 (N_2915,N_1136,N_1423);
and U2916 (N_2916,N_1118,N_1802);
nand U2917 (N_2917,N_1553,N_1563);
or U2918 (N_2918,N_1931,N_1787);
or U2919 (N_2919,N_1838,N_1480);
or U2920 (N_2920,N_1385,N_1183);
and U2921 (N_2921,N_1381,N_1667);
and U2922 (N_2922,N_1276,N_1824);
nor U2923 (N_2923,N_1591,N_1315);
nand U2924 (N_2924,N_1126,N_1575);
nor U2925 (N_2925,N_1010,N_1527);
nor U2926 (N_2926,N_1926,N_1047);
nand U2927 (N_2927,N_1432,N_1092);
nor U2928 (N_2928,N_1645,N_1912);
nor U2929 (N_2929,N_1067,N_1108);
nor U2930 (N_2930,N_1702,N_1144);
nor U2931 (N_2931,N_1241,N_1758);
nand U2932 (N_2932,N_1579,N_1616);
and U2933 (N_2933,N_1665,N_1714);
nor U2934 (N_2934,N_1734,N_1522);
nand U2935 (N_2935,N_1614,N_1295);
and U2936 (N_2936,N_1035,N_1582);
and U2937 (N_2937,N_1510,N_1883);
nor U2938 (N_2938,N_1117,N_1085);
and U2939 (N_2939,N_1720,N_1920);
or U2940 (N_2940,N_1648,N_1881);
nor U2941 (N_2941,N_1485,N_1413);
or U2942 (N_2942,N_1139,N_1290);
and U2943 (N_2943,N_1864,N_1796);
nand U2944 (N_2944,N_1208,N_1372);
nor U2945 (N_2945,N_1977,N_1596);
and U2946 (N_2946,N_1127,N_1039);
or U2947 (N_2947,N_1953,N_1260);
or U2948 (N_2948,N_1656,N_1833);
nand U2949 (N_2949,N_1350,N_1193);
or U2950 (N_2950,N_1800,N_1033);
nor U2951 (N_2951,N_1376,N_1716);
nand U2952 (N_2952,N_1708,N_1040);
and U2953 (N_2953,N_1980,N_1306);
and U2954 (N_2954,N_1810,N_1610);
or U2955 (N_2955,N_1397,N_1930);
or U2956 (N_2956,N_1580,N_1642);
or U2957 (N_2957,N_1878,N_1607);
nand U2958 (N_2958,N_1066,N_1178);
and U2959 (N_2959,N_1059,N_1064);
nor U2960 (N_2960,N_1320,N_1776);
nand U2961 (N_2961,N_1685,N_1777);
nand U2962 (N_2962,N_1416,N_1025);
or U2963 (N_2963,N_1881,N_1017);
and U2964 (N_2964,N_1722,N_1368);
and U2965 (N_2965,N_1446,N_1833);
and U2966 (N_2966,N_1080,N_1063);
and U2967 (N_2967,N_1906,N_1218);
and U2968 (N_2968,N_1154,N_1991);
nor U2969 (N_2969,N_1199,N_1177);
xor U2970 (N_2970,N_1255,N_1901);
nor U2971 (N_2971,N_1996,N_1225);
xor U2972 (N_2972,N_1162,N_1923);
nor U2973 (N_2973,N_1858,N_1603);
nand U2974 (N_2974,N_1895,N_1693);
xnor U2975 (N_2975,N_1420,N_1438);
or U2976 (N_2976,N_1193,N_1280);
and U2977 (N_2977,N_1492,N_1495);
or U2978 (N_2978,N_1664,N_1746);
nor U2979 (N_2979,N_1588,N_1581);
nor U2980 (N_2980,N_1976,N_1741);
or U2981 (N_2981,N_1461,N_1893);
nand U2982 (N_2982,N_1543,N_1530);
nand U2983 (N_2983,N_1392,N_1018);
nor U2984 (N_2984,N_1447,N_1724);
nand U2985 (N_2985,N_1468,N_1438);
and U2986 (N_2986,N_1316,N_1123);
xor U2987 (N_2987,N_1548,N_1726);
nor U2988 (N_2988,N_1334,N_1191);
nor U2989 (N_2989,N_1721,N_1037);
nand U2990 (N_2990,N_1109,N_1977);
xor U2991 (N_2991,N_1853,N_1598);
or U2992 (N_2992,N_1819,N_1616);
and U2993 (N_2993,N_1223,N_1010);
or U2994 (N_2994,N_1713,N_1584);
nor U2995 (N_2995,N_1960,N_1737);
nand U2996 (N_2996,N_1790,N_1287);
nor U2997 (N_2997,N_1734,N_1058);
nand U2998 (N_2998,N_1943,N_1244);
or U2999 (N_2999,N_1277,N_1603);
nand U3000 (N_3000,N_2721,N_2559);
nor U3001 (N_3001,N_2623,N_2614);
nand U3002 (N_3002,N_2628,N_2199);
and U3003 (N_3003,N_2536,N_2544);
nor U3004 (N_3004,N_2481,N_2941);
and U3005 (N_3005,N_2736,N_2165);
nand U3006 (N_3006,N_2786,N_2032);
xnor U3007 (N_3007,N_2316,N_2490);
or U3008 (N_3008,N_2065,N_2627);
nor U3009 (N_3009,N_2500,N_2903);
or U3010 (N_3010,N_2475,N_2154);
and U3011 (N_3011,N_2135,N_2867);
and U3012 (N_3012,N_2970,N_2625);
nor U3013 (N_3013,N_2979,N_2428);
or U3014 (N_3014,N_2422,N_2804);
and U3015 (N_3015,N_2247,N_2450);
nand U3016 (N_3016,N_2752,N_2373);
and U3017 (N_3017,N_2133,N_2036);
nor U3018 (N_3018,N_2261,N_2895);
nand U3019 (N_3019,N_2781,N_2576);
or U3020 (N_3020,N_2965,N_2825);
or U3021 (N_3021,N_2547,N_2122);
nand U3022 (N_3022,N_2933,N_2866);
and U3023 (N_3023,N_2580,N_2792);
nor U3024 (N_3024,N_2185,N_2279);
nor U3025 (N_3025,N_2458,N_2912);
or U3026 (N_3026,N_2655,N_2177);
and U3027 (N_3027,N_2106,N_2692);
nand U3028 (N_3028,N_2553,N_2515);
and U3029 (N_3029,N_2451,N_2534);
nor U3030 (N_3030,N_2243,N_2820);
nand U3031 (N_3031,N_2972,N_2691);
xor U3032 (N_3032,N_2893,N_2677);
nor U3033 (N_3033,N_2558,N_2026);
and U3034 (N_3034,N_2349,N_2619);
and U3035 (N_3035,N_2277,N_2267);
and U3036 (N_3036,N_2822,N_2003);
or U3037 (N_3037,N_2667,N_2717);
nor U3038 (N_3038,N_2735,N_2410);
or U3039 (N_3039,N_2022,N_2439);
and U3040 (N_3040,N_2270,N_2732);
nand U3041 (N_3041,N_2125,N_2132);
nand U3042 (N_3042,N_2287,N_2303);
nor U3043 (N_3043,N_2603,N_2230);
or U3044 (N_3044,N_2711,N_2621);
nor U3045 (N_3045,N_2528,N_2636);
and U3046 (N_3046,N_2518,N_2063);
nand U3047 (N_3047,N_2974,N_2309);
nor U3048 (N_3048,N_2016,N_2266);
nor U3049 (N_3049,N_2187,N_2632);
or U3050 (N_3050,N_2761,N_2138);
nor U3051 (N_3051,N_2326,N_2115);
nor U3052 (N_3052,N_2673,N_2955);
nor U3053 (N_3053,N_2647,N_2396);
xor U3054 (N_3054,N_2504,N_2447);
nor U3055 (N_3055,N_2976,N_2890);
nand U3056 (N_3056,N_2159,N_2850);
or U3057 (N_3057,N_2999,N_2669);
nand U3058 (N_3058,N_2409,N_2479);
and U3059 (N_3059,N_2947,N_2201);
nand U3060 (N_3060,N_2521,N_2973);
or U3061 (N_3061,N_2174,N_2189);
nand U3062 (N_3062,N_2148,N_2662);
or U3063 (N_3063,N_2010,N_2212);
or U3064 (N_3064,N_2314,N_2545);
or U3065 (N_3065,N_2367,N_2995);
and U3066 (N_3066,N_2363,N_2998);
and U3067 (N_3067,N_2771,N_2078);
xnor U3068 (N_3068,N_2502,N_2682);
xor U3069 (N_3069,N_2723,N_2334);
nand U3070 (N_3070,N_2983,N_2910);
nand U3071 (N_3071,N_2718,N_2206);
nand U3072 (N_3072,N_2555,N_2835);
nand U3073 (N_3073,N_2378,N_2264);
nand U3074 (N_3074,N_2787,N_2809);
or U3075 (N_3075,N_2250,N_2220);
and U3076 (N_3076,N_2629,N_2986);
and U3077 (N_3077,N_2901,N_2511);
nor U3078 (N_3078,N_2612,N_2760);
and U3079 (N_3079,N_2529,N_2088);
nand U3080 (N_3080,N_2488,N_2640);
or U3081 (N_3081,N_2676,N_2634);
nor U3082 (N_3082,N_2501,N_2366);
and U3083 (N_3083,N_2519,N_2195);
nand U3084 (N_3084,N_2100,N_2802);
or U3085 (N_3085,N_2228,N_2620);
nor U3086 (N_3086,N_2925,N_2008);
nor U3087 (N_3087,N_2583,N_2005);
or U3088 (N_3088,N_2126,N_2858);
or U3089 (N_3089,N_2778,N_2171);
nor U3090 (N_3090,N_2437,N_2921);
nand U3091 (N_3091,N_2840,N_2432);
nand U3092 (N_3092,N_2427,N_2375);
nand U3093 (N_3093,N_2800,N_2729);
or U3094 (N_3094,N_2307,N_2202);
nand U3095 (N_3095,N_2790,N_2320);
nand U3096 (N_3096,N_2384,N_2224);
and U3097 (N_3097,N_2184,N_2687);
and U3098 (N_3098,N_2932,N_2724);
and U3099 (N_3099,N_2522,N_2770);
and U3100 (N_3100,N_2657,N_2433);
or U3101 (N_3101,N_2728,N_2313);
nand U3102 (N_3102,N_2332,N_2953);
and U3103 (N_3103,N_2104,N_2915);
and U3104 (N_3104,N_2937,N_2856);
nor U3105 (N_3105,N_2278,N_2922);
and U3106 (N_3106,N_2872,N_2743);
or U3107 (N_3107,N_2219,N_2606);
nand U3108 (N_3108,N_2837,N_2507);
and U3109 (N_3109,N_2703,N_2613);
nor U3110 (N_3110,N_2441,N_2110);
nor U3111 (N_3111,N_2158,N_2830);
nor U3112 (N_3112,N_2844,N_2557);
nor U3113 (N_3113,N_2819,N_2763);
nor U3114 (N_3114,N_2582,N_2783);
or U3115 (N_3115,N_2714,N_2672);
nand U3116 (N_3116,N_2664,N_2896);
and U3117 (N_3117,N_2406,N_2708);
nand U3118 (N_3118,N_2531,N_2203);
nand U3119 (N_3119,N_2340,N_2197);
or U3120 (N_3120,N_2116,N_2080);
and U3121 (N_3121,N_2989,N_2460);
nand U3122 (N_3122,N_2288,N_2058);
nand U3123 (N_3123,N_2549,N_2855);
nor U3124 (N_3124,N_2646,N_2702);
nor U3125 (N_3125,N_2149,N_2643);
nand U3126 (N_3126,N_2767,N_2930);
nand U3127 (N_3127,N_2157,N_2801);
and U3128 (N_3128,N_2175,N_2130);
xnor U3129 (N_3129,N_2982,N_2961);
nand U3130 (N_3130,N_2674,N_2275);
and U3131 (N_3131,N_2524,N_2306);
nor U3132 (N_3132,N_2794,N_2793);
nand U3133 (N_3133,N_2814,N_2353);
nor U3134 (N_3134,N_2959,N_2269);
nand U3135 (N_3135,N_2235,N_2217);
nand U3136 (N_3136,N_2618,N_2879);
and U3137 (N_3137,N_2807,N_2570);
and U3138 (N_3138,N_2284,N_2079);
nor U3139 (N_3139,N_2376,N_2889);
nand U3140 (N_3140,N_2734,N_2514);
nand U3141 (N_3141,N_2888,N_2486);
and U3142 (N_3142,N_2589,N_2556);
or U3143 (N_3143,N_2412,N_2315);
and U3144 (N_3144,N_2321,N_2745);
nor U3145 (N_3145,N_2540,N_2000);
and U3146 (N_3146,N_2865,N_2299);
or U3147 (N_3147,N_2887,N_2136);
or U3148 (N_3148,N_2040,N_2607);
nor U3149 (N_3149,N_2706,N_2004);
and U3150 (N_3150,N_2142,N_2824);
nand U3151 (N_3151,N_2435,N_2851);
or U3152 (N_3152,N_2928,N_2029);
or U3153 (N_3153,N_2909,N_2103);
xor U3154 (N_3154,N_2030,N_2360);
or U3155 (N_3155,N_2311,N_2601);
or U3156 (N_3156,N_2140,N_2497);
nor U3157 (N_3157,N_2537,N_2805);
or U3158 (N_3158,N_2352,N_2407);
nand U3159 (N_3159,N_2411,N_2469);
nor U3160 (N_3160,N_2838,N_2225);
nand U3161 (N_3161,N_2649,N_2906);
and U3162 (N_3162,N_2654,N_2949);
and U3163 (N_3163,N_2641,N_2190);
or U3164 (N_3164,N_2948,N_2810);
and U3165 (N_3165,N_2483,N_2747);
or U3166 (N_3166,N_2290,N_2473);
or U3167 (N_3167,N_2054,N_2459);
nand U3168 (N_3168,N_2255,N_2689);
nor U3169 (N_3169,N_2684,N_2017);
nor U3170 (N_3170,N_2400,N_2957);
and U3171 (N_3171,N_2463,N_2806);
or U3172 (N_3172,N_2121,N_2695);
nand U3173 (N_3173,N_2902,N_2907);
nor U3174 (N_3174,N_2464,N_2686);
and U3175 (N_3175,N_2462,N_2826);
xor U3176 (N_3176,N_2834,N_2927);
nor U3177 (N_3177,N_2214,N_2129);
nand U3178 (N_3178,N_2229,N_2091);
or U3179 (N_3179,N_2211,N_2087);
nand U3180 (N_3180,N_2616,N_2213);
or U3181 (N_3181,N_2420,N_2938);
nand U3182 (N_3182,N_2337,N_2923);
nand U3183 (N_3183,N_2204,N_2652);
nand U3184 (N_3184,N_2798,N_2071);
nor U3185 (N_3185,N_2797,N_2942);
or U3186 (N_3186,N_2162,N_2449);
and U3187 (N_3187,N_2848,N_2232);
or U3188 (N_3188,N_2722,N_2064);
nand U3189 (N_3189,N_2997,N_2538);
nor U3190 (N_3190,N_2574,N_2585);
nor U3191 (N_3191,N_2594,N_2358);
nor U3192 (N_3192,N_2845,N_2429);
nor U3193 (N_3193,N_2759,N_2535);
or U3194 (N_3194,N_2526,N_2119);
and U3195 (N_3195,N_2050,N_2495);
and U3196 (N_3196,N_2466,N_2622);
and U3197 (N_3197,N_2045,N_2829);
or U3198 (N_3198,N_2552,N_2383);
nor U3199 (N_3199,N_2296,N_2341);
and U3200 (N_3200,N_2147,N_2234);
nor U3201 (N_3201,N_2823,N_2221);
nand U3202 (N_3202,N_2413,N_2393);
nor U3203 (N_3203,N_2985,N_2139);
nand U3204 (N_3204,N_2991,N_2283);
nand U3205 (N_3205,N_2155,N_2394);
and U3206 (N_3206,N_2775,N_2156);
nand U3207 (N_3207,N_2741,N_2263);
and U3208 (N_3208,N_2342,N_2572);
nor U3209 (N_3209,N_2812,N_2757);
nand U3210 (N_3210,N_2756,N_2963);
nand U3211 (N_3211,N_2060,N_2052);
nand U3212 (N_3212,N_2633,N_2878);
nor U3213 (N_3213,N_2239,N_2994);
and U3214 (N_3214,N_2870,N_2492);
nor U3215 (N_3215,N_2282,N_2359);
nor U3216 (N_3216,N_2874,N_2444);
nand U3217 (N_3217,N_2832,N_2681);
nand U3218 (N_3218,N_2569,N_2563);
and U3219 (N_3219,N_2385,N_2818);
nand U3220 (N_3220,N_2871,N_2018);
nor U3221 (N_3221,N_2170,N_2587);
nand U3222 (N_3222,N_2044,N_2405);
nand U3223 (N_3223,N_2377,N_2262);
nor U3224 (N_3224,N_2038,N_2461);
and U3225 (N_3225,N_2271,N_2929);
or U3226 (N_3226,N_2386,N_2470);
nor U3227 (N_3227,N_2295,N_2300);
nand U3228 (N_3228,N_2072,N_2317);
nor U3229 (N_3229,N_2608,N_2670);
or U3230 (N_3230,N_2491,N_2506);
nand U3231 (N_3231,N_2143,N_2318);
and U3232 (N_3232,N_2056,N_2426);
or U3233 (N_3233,N_2615,N_2624);
or U3234 (N_3234,N_2127,N_2176);
nor U3235 (N_3235,N_2249,N_2020);
nand U3236 (N_3236,N_2298,N_2112);
nand U3237 (N_3237,N_2180,N_2758);
nand U3238 (N_3238,N_2852,N_2988);
nor U3239 (N_3239,N_2754,N_2591);
nor U3240 (N_3240,N_2236,N_2019);
nor U3241 (N_3241,N_2712,N_2904);
and U3242 (N_3242,N_2392,N_2920);
or U3243 (N_3243,N_2274,N_2465);
and U3244 (N_3244,N_2579,N_2821);
or U3245 (N_3245,N_2877,N_2635);
nor U3246 (N_3246,N_2581,N_2251);
and U3247 (N_3247,N_2354,N_2371);
and U3248 (N_3248,N_2048,N_2067);
nand U3249 (N_3249,N_2530,N_2182);
and U3250 (N_3250,N_2053,N_2968);
and U3251 (N_3251,N_2609,N_2408);
or U3252 (N_3252,N_2561,N_2550);
nand U3253 (N_3253,N_2630,N_2006);
or U3254 (N_3254,N_2726,N_2445);
nor U3255 (N_3255,N_2338,N_2551);
nand U3256 (N_3256,N_2339,N_2859);
nor U3257 (N_3257,N_2943,N_2685);
and U3258 (N_3258,N_2323,N_2179);
nand U3259 (N_3259,N_2846,N_2192);
nand U3260 (N_3260,N_2510,N_2782);
or U3261 (N_3261,N_2764,N_2012);
and U3262 (N_3262,N_2679,N_2241);
or U3263 (N_3263,N_2543,N_2484);
and U3264 (N_3264,N_2525,N_2967);
or U3265 (N_3265,N_2931,N_2128);
and U3266 (N_3266,N_2853,N_2242);
nor U3267 (N_3267,N_2913,N_2969);
and U3268 (N_3268,N_2899,N_2467);
nor U3269 (N_3269,N_2028,N_2578);
and U3270 (N_3270,N_2161,N_2813);
nand U3271 (N_3271,N_2694,N_2472);
and U3272 (N_3272,N_2924,N_2457);
xnor U3273 (N_3273,N_2595,N_2114);
nand U3274 (N_3274,N_2671,N_2193);
nand U3275 (N_3275,N_2841,N_2645);
xnor U3276 (N_3276,N_2285,N_2831);
nor U3277 (N_3277,N_2586,N_2828);
or U3278 (N_3278,N_2259,N_2061);
nand U3279 (N_3279,N_2222,N_2885);
nor U3280 (N_3280,N_2876,N_2194);
and U3281 (N_3281,N_2597,N_2739);
nor U3282 (N_3282,N_2984,N_2066);
nand U3283 (N_3283,N_2791,N_2699);
or U3284 (N_3284,N_2697,N_2099);
nand U3285 (N_3285,N_2939,N_2293);
nand U3286 (N_3286,N_2291,N_2742);
or U3287 (N_3287,N_2057,N_2577);
or U3288 (N_3288,N_2150,N_2839);
or U3289 (N_3289,N_2328,N_2744);
nor U3290 (N_3290,N_2077,N_2868);
and U3291 (N_3291,N_2434,N_2748);
nand U3292 (N_3292,N_2978,N_2862);
or U3293 (N_3293,N_2346,N_2704);
nand U3294 (N_3294,N_2567,N_2322);
and U3295 (N_3295,N_2389,N_2568);
nor U3296 (N_3296,N_2169,N_2539);
nand U3297 (N_3297,N_2118,N_2513);
or U3298 (N_3298,N_2560,N_2663);
and U3299 (N_3299,N_2493,N_2768);
nand U3300 (N_3300,N_2404,N_2911);
and U3301 (N_3301,N_2992,N_2145);
nand U3302 (N_3302,N_2489,N_2245);
nor U3303 (N_3303,N_2163,N_2533);
and U3304 (N_3304,N_2253,N_2886);
nand U3305 (N_3305,N_2720,N_2356);
or U3306 (N_3306,N_2849,N_2546);
nand U3307 (N_3307,N_2996,N_2380);
or U3308 (N_3308,N_2598,N_2592);
nor U3309 (N_3309,N_2733,N_2120);
nand U3310 (N_3310,N_2073,N_2709);
nand U3311 (N_3311,N_2329,N_2713);
nand U3312 (N_3312,N_2951,N_2105);
and U3313 (N_3313,N_2041,N_2520);
and U3314 (N_3314,N_2842,N_2683);
nand U3315 (N_3315,N_2883,N_2347);
nand U3316 (N_3316,N_2926,N_2398);
and U3317 (N_3317,N_2207,N_2863);
nand U3318 (N_3318,N_2021,N_2059);
nor U3319 (N_3319,N_2361,N_2402);
nand U3320 (N_3320,N_2914,N_2861);
or U3321 (N_3321,N_2209,N_2715);
nor U3322 (N_3322,N_2631,N_2166);
and U3323 (N_3323,N_2095,N_2160);
and U3324 (N_3324,N_2777,N_2765);
or U3325 (N_3325,N_2651,N_2789);
nand U3326 (N_3326,N_2035,N_2456);
or U3327 (N_3327,N_2505,N_2123);
nor U3328 (N_3328,N_2496,N_2395);
or U3329 (N_3329,N_2302,N_2368);
or U3330 (N_3330,N_2605,N_2956);
nand U3331 (N_3331,N_2333,N_2331);
nor U3332 (N_3332,N_2419,N_2265);
nor U3333 (N_3333,N_2094,N_2391);
and U3334 (N_3334,N_2980,N_2693);
nor U3335 (N_3335,N_2455,N_2882);
nand U3336 (N_3336,N_2638,N_2934);
and U3337 (N_3337,N_2705,N_2575);
nand U3338 (N_3338,N_2370,N_2324);
nand U3339 (N_3339,N_2074,N_2258);
nand U3340 (N_3340,N_2892,N_2517);
nand U3341 (N_3341,N_2365,N_2590);
nand U3342 (N_3342,N_2257,N_2565);
nand U3343 (N_3343,N_2769,N_2244);
and U3344 (N_3344,N_2661,N_2372);
nor U3345 (N_3345,N_2975,N_2610);
nand U3346 (N_3346,N_2600,N_2477);
and U3347 (N_3347,N_2788,N_2289);
and U3348 (N_3348,N_2815,N_2873);
or U3349 (N_3349,N_2716,N_2131);
nor U3350 (N_3350,N_2847,N_2260);
nor U3351 (N_3351,N_2898,N_2725);
nand U3352 (N_3352,N_2098,N_2357);
nor U3353 (N_3353,N_2111,N_2113);
nand U3354 (N_3354,N_2541,N_2381);
and U3355 (N_3355,N_2678,N_2401);
nor U3356 (N_3356,N_2216,N_2109);
or U3357 (N_3357,N_2799,N_2962);
and U3358 (N_3358,N_2987,N_2141);
or U3359 (N_3359,N_2031,N_2092);
nand U3360 (N_3360,N_2055,N_2916);
and U3361 (N_3361,N_2604,N_2208);
and U3362 (N_3362,N_2237,N_2200);
and U3363 (N_3363,N_2438,N_2512);
nand U3364 (N_3364,N_2102,N_2564);
nor U3365 (N_3365,N_2548,N_2101);
nand U3366 (N_3366,N_2369,N_2144);
nor U3367 (N_3367,N_2090,N_2738);
and U3368 (N_3368,N_2780,N_2795);
and U3369 (N_3369,N_2573,N_2675);
nor U3370 (N_3370,N_2746,N_2891);
nand U3371 (N_3371,N_2453,N_2542);
or U3372 (N_3372,N_2964,N_2069);
and U3373 (N_3373,N_2343,N_2108);
nor U3374 (N_3374,N_2039,N_2919);
and U3375 (N_3375,N_2081,N_2593);
or U3376 (N_3376,N_2416,N_2656);
nor U3377 (N_3377,N_2509,N_2944);
or U3378 (N_3378,N_2917,N_2990);
nor U3379 (N_3379,N_2344,N_2700);
or U3380 (N_3380,N_2482,N_2068);
or U3381 (N_3381,N_2776,N_2042);
nor U3382 (N_3382,N_2562,N_2227);
and U3383 (N_3383,N_2796,N_2710);
nor U3384 (N_3384,N_2246,N_2226);
or U3385 (N_3385,N_2471,N_2894);
nor U3386 (N_3386,N_2854,N_2082);
or U3387 (N_3387,N_2033,N_2146);
nand U3388 (N_3388,N_2362,N_2454);
nor U3389 (N_3389,N_2336,N_2273);
and U3390 (N_3390,N_2981,N_2751);
nand U3391 (N_3391,N_2626,N_2107);
nor U3392 (N_3392,N_2173,N_2762);
or U3393 (N_3393,N_2037,N_2355);
or U3394 (N_3394,N_2025,N_2644);
and U3395 (N_3395,N_2452,N_2124);
nand U3396 (N_3396,N_2516,N_2966);
nor U3397 (N_3397,N_2294,N_2223);
nand U3398 (N_3398,N_2869,N_2688);
nor U3399 (N_3399,N_2740,N_2013);
nor U3400 (N_3400,N_2117,N_2240);
nand U3401 (N_3401,N_2875,N_2414);
or U3402 (N_3402,N_2364,N_2617);
and U3403 (N_3403,N_2905,N_2946);
xnor U3404 (N_3404,N_2046,N_2297);
and U3405 (N_3405,N_2276,N_2881);
and U3406 (N_3406,N_2774,N_2864);
or U3407 (N_3407,N_2468,N_2698);
and U3408 (N_3408,N_2730,N_2785);
or U3409 (N_3409,N_2503,N_2588);
or U3410 (N_3410,N_2476,N_2808);
and U3411 (N_3411,N_2690,N_2554);
nor U3412 (N_3412,N_2183,N_2137);
and U3413 (N_3413,N_2602,N_2084);
nand U3414 (N_3414,N_2350,N_2658);
nor U3415 (N_3415,N_2043,N_2024);
nor U3416 (N_3416,N_2047,N_2833);
nand U3417 (N_3417,N_2399,N_2430);
or U3418 (N_3418,N_2330,N_2281);
nor U3419 (N_3419,N_2034,N_2134);
nand U3420 (N_3420,N_2319,N_2415);
nor U3421 (N_3421,N_2936,N_2181);
and U3422 (N_3422,N_2374,N_2952);
nand U3423 (N_3423,N_2950,N_2523);
and U3424 (N_3424,N_2425,N_2977);
and U3425 (N_3425,N_2719,N_2773);
nor U3426 (N_3426,N_2766,N_2478);
or U3427 (N_3427,N_2960,N_2487);
nor U3428 (N_3428,N_2015,N_2571);
and U3429 (N_3429,N_2252,N_2935);
and U3430 (N_3430,N_2880,N_2784);
nor U3431 (N_3431,N_2248,N_2164);
nand U3432 (N_3432,N_2167,N_2049);
or U3433 (N_3433,N_2418,N_2945);
or U3434 (N_3434,N_2827,N_2191);
nor U3435 (N_3435,N_2308,N_2417);
and U3436 (N_3436,N_2660,N_2186);
nand U3437 (N_3437,N_2817,N_2566);
nand U3438 (N_3438,N_2954,N_2286);
or U3439 (N_3439,N_2659,N_2480);
and U3440 (N_3440,N_2231,N_2325);
and U3441 (N_3441,N_2062,N_2254);
nor U3442 (N_3442,N_2803,N_2908);
nand U3443 (N_3443,N_2648,N_2280);
or U3444 (N_3444,N_2153,N_2508);
and U3445 (N_3445,N_2218,N_2027);
nand U3446 (N_3446,N_2611,N_2215);
and U3447 (N_3447,N_2351,N_2083);
nand U3448 (N_3448,N_2993,N_2075);
and U3449 (N_3449,N_2639,N_2304);
or U3450 (N_3450,N_2527,N_2680);
xnor U3451 (N_3451,N_2755,N_2093);
nor U3452 (N_3452,N_2474,N_2707);
nand U3453 (N_3453,N_2335,N_2188);
nand U3454 (N_3454,N_2379,N_2431);
nand U3455 (N_3455,N_2390,N_2305);
nand U3456 (N_3456,N_2014,N_2498);
and U3457 (N_3457,N_2009,N_2196);
nand U3458 (N_3458,N_2151,N_2387);
or U3459 (N_3459,N_2811,N_2940);
or U3460 (N_3460,N_2696,N_2327);
nor U3461 (N_3461,N_2172,N_2011);
nor U3462 (N_3462,N_2001,N_2446);
nand U3463 (N_3463,N_2485,N_2198);
nor U3464 (N_3464,N_2421,N_2918);
or U3465 (N_3465,N_2665,N_2494);
nand U3466 (N_3466,N_2836,N_2749);
nor U3467 (N_3467,N_2268,N_2884);
nand U3468 (N_3468,N_2152,N_2584);
nand U3469 (N_3469,N_2210,N_2168);
nand U3470 (N_3470,N_2007,N_2701);
or U3471 (N_3471,N_2205,N_2971);
or U3472 (N_3472,N_2737,N_2397);
nor U3473 (N_3473,N_2436,N_2637);
nor U3474 (N_3474,N_2382,N_2097);
or U3475 (N_3475,N_2002,N_2653);
or U3476 (N_3476,N_2233,N_2023);
and U3477 (N_3477,N_2816,N_2440);
nand U3478 (N_3478,N_2085,N_2301);
and U3479 (N_3479,N_2086,N_2668);
nand U3480 (N_3480,N_2843,N_2348);
xor U3481 (N_3481,N_2345,N_2448);
or U3482 (N_3482,N_2897,N_2051);
nand U3483 (N_3483,N_2857,N_2089);
xor U3484 (N_3484,N_2238,N_2958);
or U3485 (N_3485,N_2860,N_2599);
nor U3486 (N_3486,N_2424,N_2753);
nor U3487 (N_3487,N_2070,N_2403);
nand U3488 (N_3488,N_2442,N_2076);
nor U3489 (N_3489,N_2731,N_2727);
nor U3490 (N_3490,N_2532,N_2750);
or U3491 (N_3491,N_2596,N_2312);
or U3492 (N_3492,N_2096,N_2650);
nor U3493 (N_3493,N_2779,N_2178);
nand U3494 (N_3494,N_2272,N_2499);
nand U3495 (N_3495,N_2900,N_2443);
or U3496 (N_3496,N_2310,N_2772);
nor U3497 (N_3497,N_2256,N_2388);
and U3498 (N_3498,N_2642,N_2666);
nor U3499 (N_3499,N_2292,N_2423);
nand U3500 (N_3500,N_2539,N_2025);
nand U3501 (N_3501,N_2339,N_2018);
and U3502 (N_3502,N_2945,N_2443);
or U3503 (N_3503,N_2784,N_2037);
nor U3504 (N_3504,N_2806,N_2284);
or U3505 (N_3505,N_2293,N_2643);
or U3506 (N_3506,N_2189,N_2442);
and U3507 (N_3507,N_2985,N_2765);
xor U3508 (N_3508,N_2204,N_2873);
and U3509 (N_3509,N_2456,N_2313);
nor U3510 (N_3510,N_2872,N_2676);
or U3511 (N_3511,N_2526,N_2721);
nand U3512 (N_3512,N_2821,N_2989);
or U3513 (N_3513,N_2990,N_2030);
or U3514 (N_3514,N_2828,N_2923);
nor U3515 (N_3515,N_2514,N_2164);
and U3516 (N_3516,N_2704,N_2008);
nand U3517 (N_3517,N_2133,N_2800);
and U3518 (N_3518,N_2107,N_2337);
nor U3519 (N_3519,N_2352,N_2099);
or U3520 (N_3520,N_2904,N_2586);
or U3521 (N_3521,N_2262,N_2118);
nor U3522 (N_3522,N_2510,N_2629);
and U3523 (N_3523,N_2771,N_2868);
or U3524 (N_3524,N_2071,N_2534);
nand U3525 (N_3525,N_2579,N_2685);
or U3526 (N_3526,N_2884,N_2049);
nand U3527 (N_3527,N_2127,N_2910);
nor U3528 (N_3528,N_2482,N_2546);
and U3529 (N_3529,N_2182,N_2195);
nor U3530 (N_3530,N_2787,N_2451);
or U3531 (N_3531,N_2040,N_2691);
and U3532 (N_3532,N_2228,N_2422);
and U3533 (N_3533,N_2005,N_2448);
nand U3534 (N_3534,N_2754,N_2265);
and U3535 (N_3535,N_2886,N_2101);
or U3536 (N_3536,N_2095,N_2924);
nor U3537 (N_3537,N_2543,N_2152);
or U3538 (N_3538,N_2196,N_2806);
or U3539 (N_3539,N_2923,N_2378);
nor U3540 (N_3540,N_2811,N_2112);
nor U3541 (N_3541,N_2171,N_2517);
nand U3542 (N_3542,N_2428,N_2010);
or U3543 (N_3543,N_2333,N_2581);
and U3544 (N_3544,N_2718,N_2264);
nor U3545 (N_3545,N_2316,N_2056);
and U3546 (N_3546,N_2848,N_2527);
nand U3547 (N_3547,N_2101,N_2283);
and U3548 (N_3548,N_2653,N_2384);
nor U3549 (N_3549,N_2289,N_2705);
nand U3550 (N_3550,N_2490,N_2905);
nand U3551 (N_3551,N_2519,N_2313);
nor U3552 (N_3552,N_2574,N_2641);
nand U3553 (N_3553,N_2705,N_2089);
or U3554 (N_3554,N_2142,N_2846);
nand U3555 (N_3555,N_2871,N_2048);
nand U3556 (N_3556,N_2305,N_2366);
or U3557 (N_3557,N_2467,N_2451);
or U3558 (N_3558,N_2404,N_2965);
xnor U3559 (N_3559,N_2425,N_2056);
nor U3560 (N_3560,N_2033,N_2230);
nor U3561 (N_3561,N_2158,N_2638);
and U3562 (N_3562,N_2149,N_2142);
and U3563 (N_3563,N_2731,N_2284);
nand U3564 (N_3564,N_2416,N_2851);
or U3565 (N_3565,N_2990,N_2036);
or U3566 (N_3566,N_2401,N_2740);
nand U3567 (N_3567,N_2445,N_2357);
or U3568 (N_3568,N_2155,N_2082);
or U3569 (N_3569,N_2437,N_2067);
nor U3570 (N_3570,N_2660,N_2604);
or U3571 (N_3571,N_2904,N_2591);
and U3572 (N_3572,N_2367,N_2445);
nor U3573 (N_3573,N_2292,N_2243);
nand U3574 (N_3574,N_2777,N_2169);
nor U3575 (N_3575,N_2097,N_2203);
or U3576 (N_3576,N_2138,N_2269);
or U3577 (N_3577,N_2958,N_2548);
nor U3578 (N_3578,N_2826,N_2728);
xnor U3579 (N_3579,N_2734,N_2083);
nand U3580 (N_3580,N_2233,N_2881);
and U3581 (N_3581,N_2085,N_2379);
nand U3582 (N_3582,N_2269,N_2580);
and U3583 (N_3583,N_2038,N_2257);
and U3584 (N_3584,N_2977,N_2845);
or U3585 (N_3585,N_2142,N_2701);
or U3586 (N_3586,N_2124,N_2617);
and U3587 (N_3587,N_2719,N_2177);
nand U3588 (N_3588,N_2258,N_2920);
or U3589 (N_3589,N_2642,N_2476);
or U3590 (N_3590,N_2586,N_2702);
nor U3591 (N_3591,N_2628,N_2313);
and U3592 (N_3592,N_2697,N_2405);
or U3593 (N_3593,N_2737,N_2571);
or U3594 (N_3594,N_2658,N_2114);
and U3595 (N_3595,N_2103,N_2046);
or U3596 (N_3596,N_2759,N_2638);
xnor U3597 (N_3597,N_2711,N_2238);
and U3598 (N_3598,N_2265,N_2576);
or U3599 (N_3599,N_2194,N_2619);
or U3600 (N_3600,N_2390,N_2383);
or U3601 (N_3601,N_2661,N_2431);
nand U3602 (N_3602,N_2284,N_2583);
and U3603 (N_3603,N_2368,N_2047);
nor U3604 (N_3604,N_2080,N_2231);
nand U3605 (N_3605,N_2261,N_2541);
or U3606 (N_3606,N_2310,N_2659);
and U3607 (N_3607,N_2736,N_2336);
nor U3608 (N_3608,N_2782,N_2349);
and U3609 (N_3609,N_2500,N_2461);
nand U3610 (N_3610,N_2582,N_2760);
or U3611 (N_3611,N_2848,N_2437);
or U3612 (N_3612,N_2180,N_2992);
or U3613 (N_3613,N_2364,N_2383);
nor U3614 (N_3614,N_2259,N_2774);
and U3615 (N_3615,N_2064,N_2051);
or U3616 (N_3616,N_2086,N_2467);
or U3617 (N_3617,N_2331,N_2667);
nand U3618 (N_3618,N_2863,N_2584);
nand U3619 (N_3619,N_2052,N_2613);
or U3620 (N_3620,N_2544,N_2168);
or U3621 (N_3621,N_2946,N_2630);
nand U3622 (N_3622,N_2842,N_2449);
nand U3623 (N_3623,N_2494,N_2543);
or U3624 (N_3624,N_2239,N_2591);
and U3625 (N_3625,N_2441,N_2759);
or U3626 (N_3626,N_2048,N_2769);
nand U3627 (N_3627,N_2483,N_2374);
nand U3628 (N_3628,N_2417,N_2563);
nand U3629 (N_3629,N_2251,N_2335);
xnor U3630 (N_3630,N_2870,N_2922);
nor U3631 (N_3631,N_2032,N_2746);
nor U3632 (N_3632,N_2487,N_2287);
and U3633 (N_3633,N_2241,N_2803);
or U3634 (N_3634,N_2912,N_2197);
or U3635 (N_3635,N_2919,N_2668);
or U3636 (N_3636,N_2351,N_2909);
nor U3637 (N_3637,N_2253,N_2528);
and U3638 (N_3638,N_2740,N_2368);
and U3639 (N_3639,N_2347,N_2517);
and U3640 (N_3640,N_2089,N_2812);
nor U3641 (N_3641,N_2868,N_2016);
or U3642 (N_3642,N_2600,N_2271);
nand U3643 (N_3643,N_2786,N_2792);
and U3644 (N_3644,N_2482,N_2806);
nand U3645 (N_3645,N_2278,N_2300);
or U3646 (N_3646,N_2339,N_2973);
or U3647 (N_3647,N_2620,N_2782);
nor U3648 (N_3648,N_2893,N_2005);
or U3649 (N_3649,N_2232,N_2182);
and U3650 (N_3650,N_2543,N_2448);
and U3651 (N_3651,N_2089,N_2825);
or U3652 (N_3652,N_2530,N_2930);
nand U3653 (N_3653,N_2812,N_2283);
nor U3654 (N_3654,N_2144,N_2613);
and U3655 (N_3655,N_2696,N_2186);
and U3656 (N_3656,N_2623,N_2680);
nand U3657 (N_3657,N_2981,N_2735);
nor U3658 (N_3658,N_2563,N_2286);
nor U3659 (N_3659,N_2798,N_2452);
nor U3660 (N_3660,N_2357,N_2105);
nand U3661 (N_3661,N_2238,N_2485);
nand U3662 (N_3662,N_2520,N_2619);
or U3663 (N_3663,N_2597,N_2645);
or U3664 (N_3664,N_2372,N_2335);
xnor U3665 (N_3665,N_2346,N_2229);
and U3666 (N_3666,N_2144,N_2226);
and U3667 (N_3667,N_2202,N_2182);
or U3668 (N_3668,N_2979,N_2030);
or U3669 (N_3669,N_2243,N_2118);
nor U3670 (N_3670,N_2165,N_2162);
or U3671 (N_3671,N_2859,N_2914);
nand U3672 (N_3672,N_2567,N_2054);
nor U3673 (N_3673,N_2886,N_2527);
nor U3674 (N_3674,N_2826,N_2721);
or U3675 (N_3675,N_2318,N_2464);
and U3676 (N_3676,N_2555,N_2187);
nor U3677 (N_3677,N_2934,N_2736);
nor U3678 (N_3678,N_2393,N_2590);
nand U3679 (N_3679,N_2012,N_2918);
and U3680 (N_3680,N_2016,N_2028);
xor U3681 (N_3681,N_2250,N_2390);
and U3682 (N_3682,N_2385,N_2354);
or U3683 (N_3683,N_2679,N_2406);
and U3684 (N_3684,N_2796,N_2519);
and U3685 (N_3685,N_2153,N_2074);
and U3686 (N_3686,N_2998,N_2602);
and U3687 (N_3687,N_2926,N_2158);
nand U3688 (N_3688,N_2575,N_2300);
or U3689 (N_3689,N_2380,N_2113);
nor U3690 (N_3690,N_2648,N_2875);
and U3691 (N_3691,N_2847,N_2878);
or U3692 (N_3692,N_2778,N_2800);
nand U3693 (N_3693,N_2841,N_2812);
and U3694 (N_3694,N_2558,N_2796);
nand U3695 (N_3695,N_2367,N_2294);
and U3696 (N_3696,N_2442,N_2629);
nor U3697 (N_3697,N_2239,N_2217);
nand U3698 (N_3698,N_2962,N_2678);
or U3699 (N_3699,N_2238,N_2414);
or U3700 (N_3700,N_2990,N_2641);
nand U3701 (N_3701,N_2001,N_2461);
and U3702 (N_3702,N_2045,N_2853);
and U3703 (N_3703,N_2002,N_2977);
nor U3704 (N_3704,N_2012,N_2787);
nor U3705 (N_3705,N_2259,N_2669);
and U3706 (N_3706,N_2656,N_2074);
or U3707 (N_3707,N_2468,N_2965);
nand U3708 (N_3708,N_2262,N_2369);
or U3709 (N_3709,N_2801,N_2578);
nor U3710 (N_3710,N_2756,N_2657);
nor U3711 (N_3711,N_2487,N_2228);
and U3712 (N_3712,N_2117,N_2332);
or U3713 (N_3713,N_2418,N_2826);
and U3714 (N_3714,N_2995,N_2298);
nor U3715 (N_3715,N_2050,N_2011);
and U3716 (N_3716,N_2270,N_2831);
and U3717 (N_3717,N_2849,N_2972);
and U3718 (N_3718,N_2194,N_2590);
and U3719 (N_3719,N_2379,N_2539);
nor U3720 (N_3720,N_2575,N_2307);
or U3721 (N_3721,N_2284,N_2396);
or U3722 (N_3722,N_2755,N_2466);
and U3723 (N_3723,N_2155,N_2962);
and U3724 (N_3724,N_2502,N_2960);
nand U3725 (N_3725,N_2033,N_2038);
or U3726 (N_3726,N_2235,N_2900);
nor U3727 (N_3727,N_2824,N_2627);
nor U3728 (N_3728,N_2620,N_2253);
or U3729 (N_3729,N_2128,N_2812);
nand U3730 (N_3730,N_2499,N_2540);
nand U3731 (N_3731,N_2345,N_2010);
and U3732 (N_3732,N_2974,N_2473);
or U3733 (N_3733,N_2016,N_2054);
and U3734 (N_3734,N_2140,N_2278);
and U3735 (N_3735,N_2653,N_2319);
xor U3736 (N_3736,N_2042,N_2394);
nand U3737 (N_3737,N_2383,N_2951);
or U3738 (N_3738,N_2712,N_2733);
and U3739 (N_3739,N_2907,N_2640);
or U3740 (N_3740,N_2009,N_2433);
nand U3741 (N_3741,N_2522,N_2340);
or U3742 (N_3742,N_2476,N_2877);
nand U3743 (N_3743,N_2473,N_2730);
or U3744 (N_3744,N_2660,N_2651);
xnor U3745 (N_3745,N_2015,N_2248);
and U3746 (N_3746,N_2955,N_2194);
xnor U3747 (N_3747,N_2466,N_2750);
and U3748 (N_3748,N_2477,N_2233);
and U3749 (N_3749,N_2923,N_2434);
nor U3750 (N_3750,N_2126,N_2001);
and U3751 (N_3751,N_2255,N_2304);
nand U3752 (N_3752,N_2499,N_2841);
and U3753 (N_3753,N_2685,N_2598);
and U3754 (N_3754,N_2933,N_2525);
or U3755 (N_3755,N_2268,N_2127);
nand U3756 (N_3756,N_2922,N_2365);
nor U3757 (N_3757,N_2269,N_2603);
nand U3758 (N_3758,N_2028,N_2374);
nand U3759 (N_3759,N_2588,N_2997);
or U3760 (N_3760,N_2993,N_2445);
xor U3761 (N_3761,N_2062,N_2029);
and U3762 (N_3762,N_2091,N_2910);
and U3763 (N_3763,N_2310,N_2019);
nor U3764 (N_3764,N_2407,N_2867);
nor U3765 (N_3765,N_2904,N_2387);
and U3766 (N_3766,N_2151,N_2078);
nor U3767 (N_3767,N_2163,N_2991);
and U3768 (N_3768,N_2135,N_2786);
and U3769 (N_3769,N_2551,N_2505);
and U3770 (N_3770,N_2822,N_2560);
nor U3771 (N_3771,N_2008,N_2443);
nand U3772 (N_3772,N_2961,N_2425);
xnor U3773 (N_3773,N_2767,N_2695);
and U3774 (N_3774,N_2020,N_2857);
nor U3775 (N_3775,N_2648,N_2445);
nor U3776 (N_3776,N_2505,N_2707);
or U3777 (N_3777,N_2313,N_2619);
and U3778 (N_3778,N_2834,N_2622);
nand U3779 (N_3779,N_2332,N_2871);
or U3780 (N_3780,N_2472,N_2048);
and U3781 (N_3781,N_2200,N_2586);
nand U3782 (N_3782,N_2051,N_2644);
or U3783 (N_3783,N_2940,N_2715);
nand U3784 (N_3784,N_2881,N_2567);
or U3785 (N_3785,N_2078,N_2818);
xnor U3786 (N_3786,N_2767,N_2647);
nand U3787 (N_3787,N_2805,N_2853);
or U3788 (N_3788,N_2312,N_2689);
or U3789 (N_3789,N_2663,N_2059);
and U3790 (N_3790,N_2558,N_2865);
xnor U3791 (N_3791,N_2591,N_2725);
or U3792 (N_3792,N_2988,N_2938);
nand U3793 (N_3793,N_2649,N_2480);
xor U3794 (N_3794,N_2783,N_2847);
or U3795 (N_3795,N_2349,N_2461);
and U3796 (N_3796,N_2064,N_2544);
or U3797 (N_3797,N_2916,N_2193);
xor U3798 (N_3798,N_2634,N_2463);
nand U3799 (N_3799,N_2887,N_2396);
or U3800 (N_3800,N_2052,N_2687);
nor U3801 (N_3801,N_2296,N_2551);
or U3802 (N_3802,N_2701,N_2864);
nand U3803 (N_3803,N_2221,N_2361);
xor U3804 (N_3804,N_2526,N_2866);
or U3805 (N_3805,N_2418,N_2248);
or U3806 (N_3806,N_2587,N_2441);
and U3807 (N_3807,N_2723,N_2744);
and U3808 (N_3808,N_2116,N_2446);
and U3809 (N_3809,N_2454,N_2960);
or U3810 (N_3810,N_2157,N_2386);
nand U3811 (N_3811,N_2431,N_2939);
nand U3812 (N_3812,N_2985,N_2831);
nor U3813 (N_3813,N_2134,N_2986);
and U3814 (N_3814,N_2028,N_2612);
or U3815 (N_3815,N_2958,N_2200);
or U3816 (N_3816,N_2504,N_2822);
nand U3817 (N_3817,N_2382,N_2680);
or U3818 (N_3818,N_2157,N_2804);
nand U3819 (N_3819,N_2098,N_2479);
and U3820 (N_3820,N_2099,N_2515);
xor U3821 (N_3821,N_2336,N_2089);
and U3822 (N_3822,N_2423,N_2718);
or U3823 (N_3823,N_2984,N_2424);
nand U3824 (N_3824,N_2356,N_2701);
nor U3825 (N_3825,N_2827,N_2777);
and U3826 (N_3826,N_2465,N_2816);
nand U3827 (N_3827,N_2540,N_2996);
xnor U3828 (N_3828,N_2583,N_2664);
or U3829 (N_3829,N_2695,N_2754);
nand U3830 (N_3830,N_2238,N_2159);
and U3831 (N_3831,N_2644,N_2156);
or U3832 (N_3832,N_2625,N_2527);
xnor U3833 (N_3833,N_2270,N_2182);
or U3834 (N_3834,N_2112,N_2343);
and U3835 (N_3835,N_2377,N_2871);
or U3836 (N_3836,N_2362,N_2623);
or U3837 (N_3837,N_2707,N_2800);
and U3838 (N_3838,N_2435,N_2663);
and U3839 (N_3839,N_2949,N_2133);
or U3840 (N_3840,N_2282,N_2751);
and U3841 (N_3841,N_2005,N_2867);
nand U3842 (N_3842,N_2685,N_2416);
nand U3843 (N_3843,N_2668,N_2417);
nand U3844 (N_3844,N_2904,N_2318);
or U3845 (N_3845,N_2598,N_2535);
nor U3846 (N_3846,N_2373,N_2582);
or U3847 (N_3847,N_2718,N_2064);
nand U3848 (N_3848,N_2813,N_2288);
nor U3849 (N_3849,N_2900,N_2296);
and U3850 (N_3850,N_2612,N_2508);
nor U3851 (N_3851,N_2913,N_2764);
nand U3852 (N_3852,N_2725,N_2689);
nor U3853 (N_3853,N_2115,N_2334);
nor U3854 (N_3854,N_2472,N_2454);
nor U3855 (N_3855,N_2410,N_2229);
nand U3856 (N_3856,N_2495,N_2855);
and U3857 (N_3857,N_2150,N_2092);
and U3858 (N_3858,N_2705,N_2852);
or U3859 (N_3859,N_2807,N_2524);
or U3860 (N_3860,N_2568,N_2357);
or U3861 (N_3861,N_2019,N_2199);
nand U3862 (N_3862,N_2896,N_2253);
and U3863 (N_3863,N_2972,N_2992);
nand U3864 (N_3864,N_2774,N_2245);
and U3865 (N_3865,N_2915,N_2087);
nor U3866 (N_3866,N_2468,N_2163);
and U3867 (N_3867,N_2610,N_2344);
nand U3868 (N_3868,N_2695,N_2126);
or U3869 (N_3869,N_2929,N_2840);
or U3870 (N_3870,N_2209,N_2430);
or U3871 (N_3871,N_2344,N_2293);
nand U3872 (N_3872,N_2963,N_2349);
nand U3873 (N_3873,N_2726,N_2296);
and U3874 (N_3874,N_2097,N_2058);
nor U3875 (N_3875,N_2193,N_2549);
nand U3876 (N_3876,N_2609,N_2592);
or U3877 (N_3877,N_2969,N_2236);
nor U3878 (N_3878,N_2961,N_2217);
and U3879 (N_3879,N_2780,N_2309);
and U3880 (N_3880,N_2783,N_2107);
nand U3881 (N_3881,N_2619,N_2813);
or U3882 (N_3882,N_2158,N_2342);
nand U3883 (N_3883,N_2381,N_2503);
or U3884 (N_3884,N_2997,N_2736);
or U3885 (N_3885,N_2883,N_2693);
and U3886 (N_3886,N_2521,N_2347);
nand U3887 (N_3887,N_2459,N_2404);
nand U3888 (N_3888,N_2691,N_2468);
or U3889 (N_3889,N_2792,N_2859);
and U3890 (N_3890,N_2370,N_2383);
and U3891 (N_3891,N_2308,N_2450);
nand U3892 (N_3892,N_2276,N_2709);
nand U3893 (N_3893,N_2951,N_2175);
or U3894 (N_3894,N_2795,N_2679);
nand U3895 (N_3895,N_2722,N_2098);
nor U3896 (N_3896,N_2343,N_2885);
and U3897 (N_3897,N_2284,N_2642);
and U3898 (N_3898,N_2401,N_2965);
nor U3899 (N_3899,N_2877,N_2147);
nor U3900 (N_3900,N_2797,N_2878);
nor U3901 (N_3901,N_2462,N_2011);
nand U3902 (N_3902,N_2160,N_2441);
or U3903 (N_3903,N_2279,N_2073);
and U3904 (N_3904,N_2698,N_2736);
and U3905 (N_3905,N_2086,N_2929);
and U3906 (N_3906,N_2794,N_2630);
nand U3907 (N_3907,N_2147,N_2996);
nand U3908 (N_3908,N_2726,N_2806);
nand U3909 (N_3909,N_2943,N_2052);
or U3910 (N_3910,N_2485,N_2340);
nor U3911 (N_3911,N_2422,N_2448);
or U3912 (N_3912,N_2396,N_2518);
or U3913 (N_3913,N_2238,N_2890);
nor U3914 (N_3914,N_2521,N_2334);
nor U3915 (N_3915,N_2975,N_2675);
or U3916 (N_3916,N_2082,N_2823);
or U3917 (N_3917,N_2018,N_2311);
nor U3918 (N_3918,N_2493,N_2607);
or U3919 (N_3919,N_2816,N_2426);
and U3920 (N_3920,N_2232,N_2356);
and U3921 (N_3921,N_2860,N_2996);
nor U3922 (N_3922,N_2917,N_2092);
and U3923 (N_3923,N_2087,N_2989);
or U3924 (N_3924,N_2541,N_2669);
nor U3925 (N_3925,N_2925,N_2014);
nor U3926 (N_3926,N_2263,N_2641);
nand U3927 (N_3927,N_2233,N_2162);
or U3928 (N_3928,N_2151,N_2521);
and U3929 (N_3929,N_2051,N_2689);
and U3930 (N_3930,N_2356,N_2519);
nand U3931 (N_3931,N_2891,N_2734);
or U3932 (N_3932,N_2460,N_2632);
or U3933 (N_3933,N_2357,N_2856);
nand U3934 (N_3934,N_2767,N_2314);
nor U3935 (N_3935,N_2620,N_2165);
or U3936 (N_3936,N_2352,N_2313);
or U3937 (N_3937,N_2475,N_2949);
nor U3938 (N_3938,N_2582,N_2806);
nor U3939 (N_3939,N_2472,N_2143);
and U3940 (N_3940,N_2860,N_2568);
nor U3941 (N_3941,N_2610,N_2948);
and U3942 (N_3942,N_2989,N_2740);
and U3943 (N_3943,N_2356,N_2192);
and U3944 (N_3944,N_2541,N_2568);
or U3945 (N_3945,N_2990,N_2718);
nand U3946 (N_3946,N_2836,N_2570);
nor U3947 (N_3947,N_2462,N_2969);
nor U3948 (N_3948,N_2175,N_2337);
nand U3949 (N_3949,N_2798,N_2714);
nor U3950 (N_3950,N_2566,N_2231);
nor U3951 (N_3951,N_2877,N_2875);
nor U3952 (N_3952,N_2325,N_2206);
and U3953 (N_3953,N_2052,N_2164);
nand U3954 (N_3954,N_2525,N_2845);
nor U3955 (N_3955,N_2514,N_2857);
nor U3956 (N_3956,N_2304,N_2244);
or U3957 (N_3957,N_2098,N_2383);
nand U3958 (N_3958,N_2839,N_2770);
nand U3959 (N_3959,N_2551,N_2929);
nor U3960 (N_3960,N_2660,N_2500);
nor U3961 (N_3961,N_2701,N_2128);
or U3962 (N_3962,N_2046,N_2776);
or U3963 (N_3963,N_2157,N_2860);
or U3964 (N_3964,N_2040,N_2131);
nand U3965 (N_3965,N_2762,N_2777);
nand U3966 (N_3966,N_2338,N_2298);
or U3967 (N_3967,N_2996,N_2605);
xnor U3968 (N_3968,N_2279,N_2628);
and U3969 (N_3969,N_2645,N_2470);
and U3970 (N_3970,N_2294,N_2659);
or U3971 (N_3971,N_2370,N_2218);
nand U3972 (N_3972,N_2622,N_2451);
and U3973 (N_3973,N_2181,N_2645);
nand U3974 (N_3974,N_2076,N_2941);
or U3975 (N_3975,N_2768,N_2215);
nor U3976 (N_3976,N_2909,N_2756);
or U3977 (N_3977,N_2221,N_2375);
nand U3978 (N_3978,N_2361,N_2040);
and U3979 (N_3979,N_2963,N_2771);
nor U3980 (N_3980,N_2379,N_2898);
nand U3981 (N_3981,N_2038,N_2755);
or U3982 (N_3982,N_2666,N_2129);
and U3983 (N_3983,N_2144,N_2850);
nand U3984 (N_3984,N_2713,N_2505);
or U3985 (N_3985,N_2756,N_2302);
and U3986 (N_3986,N_2632,N_2493);
nor U3987 (N_3987,N_2939,N_2618);
nand U3988 (N_3988,N_2467,N_2125);
nor U3989 (N_3989,N_2497,N_2217);
nand U3990 (N_3990,N_2165,N_2591);
nor U3991 (N_3991,N_2010,N_2818);
nor U3992 (N_3992,N_2218,N_2212);
nand U3993 (N_3993,N_2982,N_2627);
nor U3994 (N_3994,N_2265,N_2899);
xor U3995 (N_3995,N_2281,N_2229);
or U3996 (N_3996,N_2716,N_2738);
or U3997 (N_3997,N_2473,N_2751);
or U3998 (N_3998,N_2019,N_2345);
nand U3999 (N_3999,N_2627,N_2039);
nand U4000 (N_4000,N_3453,N_3238);
or U4001 (N_4001,N_3035,N_3278);
and U4002 (N_4002,N_3855,N_3875);
and U4003 (N_4003,N_3448,N_3868);
nor U4004 (N_4004,N_3378,N_3679);
nor U4005 (N_4005,N_3016,N_3173);
nand U4006 (N_4006,N_3252,N_3121);
or U4007 (N_4007,N_3330,N_3223);
nand U4008 (N_4008,N_3407,N_3484);
nand U4009 (N_4009,N_3648,N_3400);
nor U4010 (N_4010,N_3753,N_3233);
or U4011 (N_4011,N_3549,N_3327);
and U4012 (N_4012,N_3915,N_3879);
and U4013 (N_4013,N_3161,N_3669);
nand U4014 (N_4014,N_3235,N_3073);
and U4015 (N_4015,N_3214,N_3272);
or U4016 (N_4016,N_3187,N_3156);
xnor U4017 (N_4017,N_3832,N_3478);
nand U4018 (N_4018,N_3998,N_3396);
nand U4019 (N_4019,N_3019,N_3319);
and U4020 (N_4020,N_3629,N_3651);
nor U4021 (N_4021,N_3772,N_3706);
xnor U4022 (N_4022,N_3236,N_3819);
and U4023 (N_4023,N_3461,N_3215);
or U4024 (N_4024,N_3137,N_3477);
nand U4025 (N_4025,N_3863,N_3334);
nor U4026 (N_4026,N_3425,N_3075);
and U4027 (N_4027,N_3259,N_3899);
nor U4028 (N_4028,N_3661,N_3471);
and U4029 (N_4029,N_3514,N_3351);
nand U4030 (N_4030,N_3206,N_3147);
nand U4031 (N_4031,N_3049,N_3690);
nand U4032 (N_4032,N_3548,N_3050);
or U4033 (N_4033,N_3650,N_3955);
or U4034 (N_4034,N_3796,N_3129);
or U4035 (N_4035,N_3495,N_3540);
or U4036 (N_4036,N_3560,N_3285);
or U4037 (N_4037,N_3139,N_3784);
nor U4038 (N_4038,N_3756,N_3555);
nand U4039 (N_4039,N_3444,N_3992);
nor U4040 (N_4040,N_3126,N_3810);
or U4041 (N_4041,N_3601,N_3339);
and U4042 (N_4042,N_3504,N_3685);
nand U4043 (N_4043,N_3397,N_3506);
nand U4044 (N_4044,N_3467,N_3956);
xor U4045 (N_4045,N_3482,N_3203);
and U4046 (N_4046,N_3036,N_3337);
nand U4047 (N_4047,N_3011,N_3503);
xor U4048 (N_4048,N_3727,N_3287);
and U4049 (N_4049,N_3441,N_3342);
nor U4050 (N_4050,N_3698,N_3054);
xor U4051 (N_4051,N_3553,N_3394);
nor U4052 (N_4052,N_3304,N_3057);
and U4053 (N_4053,N_3204,N_3313);
nand U4054 (N_4054,N_3346,N_3357);
nand U4055 (N_4055,N_3616,N_3686);
nor U4056 (N_4056,N_3886,N_3427);
and U4057 (N_4057,N_3020,N_3547);
and U4058 (N_4058,N_3712,N_3390);
nand U4059 (N_4059,N_3635,N_3680);
nor U4060 (N_4060,N_3314,N_3537);
and U4061 (N_4061,N_3360,N_3530);
nand U4062 (N_4062,N_3100,N_3527);
and U4063 (N_4063,N_3630,N_3830);
and U4064 (N_4064,N_3306,N_3595);
or U4065 (N_4065,N_3406,N_3789);
nor U4066 (N_4066,N_3300,N_3438);
and U4067 (N_4067,N_3095,N_3571);
and U4068 (N_4068,N_3762,N_3133);
or U4069 (N_4069,N_3399,N_3625);
nand U4070 (N_4070,N_3589,N_3802);
and U4071 (N_4071,N_3740,N_3115);
or U4072 (N_4072,N_3212,N_3485);
or U4073 (N_4073,N_3720,N_3920);
and U4074 (N_4074,N_3454,N_3801);
nor U4075 (N_4075,N_3096,N_3561);
and U4076 (N_4076,N_3528,N_3646);
or U4077 (N_4077,N_3568,N_3183);
nor U4078 (N_4078,N_3492,N_3715);
nor U4079 (N_4079,N_3499,N_3718);
nor U4080 (N_4080,N_3055,N_3457);
and U4081 (N_4081,N_3961,N_3687);
and U4082 (N_4082,N_3490,N_3671);
nand U4083 (N_4083,N_3769,N_3930);
nor U4084 (N_4084,N_3613,N_3475);
nor U4085 (N_4085,N_3840,N_3729);
nand U4086 (N_4086,N_3984,N_3921);
and U4087 (N_4087,N_3246,N_3231);
nor U4088 (N_4088,N_3140,N_3089);
nand U4089 (N_4089,N_3315,N_3615);
nor U4090 (N_4090,N_3431,N_3426);
and U4091 (N_4091,N_3531,N_3277);
nor U4092 (N_4092,N_3888,N_3707);
or U4093 (N_4093,N_3710,N_3048);
and U4094 (N_4094,N_3436,N_3655);
nand U4095 (N_4095,N_3579,N_3437);
nor U4096 (N_4096,N_3744,N_3349);
nor U4097 (N_4097,N_3205,N_3385);
and U4098 (N_4098,N_3823,N_3312);
nand U4099 (N_4099,N_3544,N_3507);
and U4100 (N_4100,N_3626,N_3760);
and U4101 (N_4101,N_3132,N_3862);
nor U4102 (N_4102,N_3329,N_3127);
nand U4103 (N_4103,N_3853,N_3841);
nand U4104 (N_4104,N_3083,N_3825);
nand U4105 (N_4105,N_3415,N_3939);
nand U4106 (N_4106,N_3505,N_3751);
nand U4107 (N_4107,N_3014,N_3642);
nand U4108 (N_4108,N_3747,N_3692);
and U4109 (N_4109,N_3344,N_3367);
or U4110 (N_4110,N_3979,N_3456);
nor U4111 (N_4111,N_3632,N_3382);
nor U4112 (N_4112,N_3901,N_3827);
and U4113 (N_4113,N_3677,N_3617);
nor U4114 (N_4114,N_3150,N_3067);
nor U4115 (N_4115,N_3084,N_3764);
nor U4116 (N_4116,N_3276,N_3237);
and U4117 (N_4117,N_3922,N_3975);
and U4118 (N_4118,N_3874,N_3416);
nor U4119 (N_4119,N_3672,N_3366);
nor U4120 (N_4120,N_3573,N_3852);
or U4121 (N_4121,N_3638,N_3871);
and U4122 (N_4122,N_3608,N_3804);
or U4123 (N_4123,N_3216,N_3972);
or U4124 (N_4124,N_3009,N_3820);
nand U4125 (N_4125,N_3146,N_3105);
or U4126 (N_4126,N_3594,N_3887);
nor U4127 (N_4127,N_3917,N_3192);
nor U4128 (N_4128,N_3567,N_3848);
nor U4129 (N_4129,N_3502,N_3576);
nor U4130 (N_4130,N_3501,N_3128);
nor U4131 (N_4131,N_3213,N_3986);
or U4132 (N_4132,N_3976,N_3735);
xor U4133 (N_4133,N_3851,N_3022);
nor U4134 (N_4134,N_3045,N_3843);
or U4135 (N_4135,N_3417,N_3782);
nor U4136 (N_4136,N_3834,N_3535);
and U4137 (N_4137,N_3299,N_3383);
nand U4138 (N_4138,N_3470,N_3831);
nand U4139 (N_4139,N_3713,N_3645);
and U4140 (N_4140,N_3934,N_3787);
and U4141 (N_4141,N_3565,N_3509);
or U4142 (N_4142,N_3323,N_3420);
and U4143 (N_4143,N_3186,N_3633);
and U4144 (N_4144,N_3451,N_3062);
nor U4145 (N_4145,N_3781,N_3480);
nor U4146 (N_4146,N_3167,N_3592);
nand U4147 (N_4147,N_3119,N_3861);
or U4148 (N_4148,N_3041,N_3900);
or U4149 (N_4149,N_3987,N_3380);
and U4150 (N_4150,N_3963,N_3971);
nand U4151 (N_4151,N_3335,N_3890);
and U4152 (N_4152,N_3941,N_3950);
or U4153 (N_4153,N_3010,N_3993);
or U4154 (N_4154,N_3389,N_3379);
or U4155 (N_4155,N_3556,N_3908);
or U4156 (N_4156,N_3469,N_3533);
xnor U4157 (N_4157,N_3865,N_3893);
nand U4158 (N_4158,N_3543,N_3051);
or U4159 (N_4159,N_3234,N_3190);
or U4160 (N_4160,N_3464,N_3809);
nand U4161 (N_4161,N_3878,N_3797);
and U4162 (N_4162,N_3138,N_3085);
nand U4163 (N_4163,N_3824,N_3008);
and U4164 (N_4164,N_3116,N_3157);
and U4165 (N_4165,N_3726,N_3557);
nor U4166 (N_4166,N_3130,N_3208);
or U4167 (N_4167,N_3402,N_3948);
and U4168 (N_4168,N_3585,N_3295);
xor U4169 (N_4169,N_3230,N_3359);
nand U4170 (N_4170,N_3826,N_3224);
nand U4171 (N_4171,N_3962,N_3714);
or U4172 (N_4172,N_3700,N_3298);
and U4173 (N_4173,N_3405,N_3012);
nand U4174 (N_4174,N_3967,N_3310);
nor U4175 (N_4175,N_3813,N_3375);
and U4176 (N_4176,N_3099,N_3833);
nand U4177 (N_4177,N_3933,N_3628);
or U4178 (N_4178,N_3763,N_3184);
or U4179 (N_4179,N_3404,N_3732);
nand U4180 (N_4180,N_3191,N_3725);
nand U4181 (N_4181,N_3551,N_3286);
or U4182 (N_4182,N_3609,N_3989);
and U4183 (N_4183,N_3403,N_3430);
or U4184 (N_4184,N_3957,N_3822);
nand U4185 (N_4185,N_3786,N_3031);
nor U4186 (N_4186,N_3268,N_3296);
and U4187 (N_4187,N_3262,N_3421);
nand U4188 (N_4188,N_3949,N_3766);
and U4189 (N_4189,N_3973,N_3647);
nand U4190 (N_4190,N_3952,N_3331);
nand U4191 (N_4191,N_3711,N_3866);
nor U4192 (N_4192,N_3068,N_3450);
nand U4193 (N_4193,N_3355,N_3123);
nor U4194 (N_4194,N_3033,N_3520);
or U4195 (N_4195,N_3256,N_3736);
or U4196 (N_4196,N_3369,N_3472);
xor U4197 (N_4197,N_3688,N_3927);
and U4198 (N_4198,N_3023,N_3552);
and U4199 (N_4199,N_3596,N_3985);
and U4200 (N_4200,N_3284,N_3515);
and U4201 (N_4201,N_3704,N_3320);
nand U4202 (N_4202,N_3293,N_3849);
and U4203 (N_4203,N_3336,N_3294);
or U4204 (N_4204,N_3829,N_3353);
nand U4205 (N_4205,N_3523,N_3244);
nor U4206 (N_4206,N_3429,N_3869);
xor U4207 (N_4207,N_3065,N_3803);
and U4208 (N_4208,N_3498,N_3850);
and U4209 (N_4209,N_3303,N_3525);
or U4210 (N_4210,N_3649,N_3876);
nand U4211 (N_4211,N_3697,N_3247);
or U4212 (N_4212,N_3860,N_3978);
and U4213 (N_4213,N_3667,N_3932);
and U4214 (N_4214,N_3542,N_3025);
and U4215 (N_4215,N_3053,N_3343);
nor U4216 (N_4216,N_3828,N_3643);
nor U4217 (N_4217,N_3266,N_3746);
nand U4218 (N_4218,N_3015,N_3027);
or U4219 (N_4219,N_3665,N_3196);
nand U4220 (N_4220,N_3659,N_3269);
or U4221 (N_4221,N_3386,N_3856);
or U4222 (N_4222,N_3546,N_3193);
or U4223 (N_4223,N_3977,N_3462);
or U4224 (N_4224,N_3563,N_3097);
nor U4225 (N_4225,N_3951,N_3775);
or U4226 (N_4226,N_3522,N_3757);
and U4227 (N_4227,N_3370,N_3728);
or U4228 (N_4228,N_3107,N_3974);
and U4229 (N_4229,N_3674,N_3148);
and U4230 (N_4230,N_3142,N_3924);
or U4231 (N_4231,N_3220,N_3481);
xor U4232 (N_4232,N_3063,N_3905);
nand U4233 (N_4233,N_3812,N_3603);
or U4234 (N_4234,N_3254,N_3854);
or U4235 (N_4235,N_3722,N_3814);
and U4236 (N_4236,N_3387,N_3612);
and U4237 (N_4237,N_3703,N_3047);
or U4238 (N_4238,N_3108,N_3424);
nand U4239 (N_4239,N_3326,N_3037);
or U4240 (N_4240,N_3516,N_3241);
nand U4241 (N_4241,N_3903,N_3322);
xor U4242 (N_4242,N_3889,N_3759);
and U4243 (N_4243,N_3496,N_3258);
and U4244 (N_4244,N_3474,N_3719);
nor U4245 (N_4245,N_3926,N_3584);
or U4246 (N_4246,N_3837,N_3434);
and U4247 (N_4247,N_3572,N_3311);
nor U4248 (N_4248,N_3906,N_3101);
nand U4249 (N_4249,N_3885,N_3811);
and U4250 (N_4250,N_3966,N_3188);
nand U4251 (N_4251,N_3517,N_3001);
or U4252 (N_4252,N_3449,N_3122);
or U4253 (N_4253,N_3656,N_3884);
and U4254 (N_4254,N_3578,N_3857);
nor U4255 (N_4255,N_3169,N_3182);
nand U4256 (N_4256,N_3080,N_3172);
or U4257 (N_4257,N_3468,N_3755);
nor U4258 (N_4258,N_3701,N_3566);
nor U4259 (N_4259,N_3634,N_3816);
and U4260 (N_4260,N_3891,N_3730);
nand U4261 (N_4261,N_3705,N_3631);
nand U4262 (N_4262,N_3070,N_3093);
nor U4263 (N_4263,N_3131,N_3597);
nand U4264 (N_4264,N_3271,N_3770);
nor U4265 (N_4265,N_3219,N_3491);
or U4266 (N_4266,N_3393,N_3395);
nand U4267 (N_4267,N_3078,N_3873);
and U4268 (N_4268,N_3221,N_3748);
and U4269 (N_4269,N_3145,N_3297);
or U4270 (N_4270,N_3724,N_3897);
nand U4271 (N_4271,N_3177,N_3652);
and U4272 (N_4272,N_3739,N_3338);
and U4273 (N_4273,N_3800,N_3526);
or U4274 (N_4274,N_3524,N_3895);
or U4275 (N_4275,N_3004,N_3202);
or U4276 (N_4276,N_3198,N_3185);
and U4277 (N_4277,N_3006,N_3087);
or U4278 (N_4278,N_3788,N_3153);
and U4279 (N_4279,N_3919,N_3489);
nor U4280 (N_4280,N_3239,N_3529);
nand U4281 (N_4281,N_3281,N_3500);
and U4282 (N_4282,N_3721,N_3301);
or U4283 (N_4283,N_3799,N_3898);
and U4284 (N_4284,N_3743,N_3681);
nor U4285 (N_4285,N_3569,N_3280);
or U4286 (N_4286,N_3918,N_3110);
nor U4287 (N_4287,N_3002,N_3066);
or U4288 (N_4288,N_3162,N_3991);
and U4289 (N_4289,N_3733,N_3088);
nand U4290 (N_4290,N_3793,N_3668);
or U4291 (N_4291,N_3790,N_3061);
or U4292 (N_4292,N_3845,N_3442);
or U4293 (N_4293,N_3988,N_3154);
nand U4294 (N_4294,N_3414,N_3767);
xnor U4295 (N_4295,N_3494,N_3654);
or U4296 (N_4296,N_3175,N_3745);
nor U4297 (N_4297,N_3624,N_3664);
and U4298 (N_4298,N_3550,N_3410);
or U4299 (N_4299,N_3907,N_3598);
nor U4300 (N_4300,N_3689,N_3465);
nor U4301 (N_4301,N_3493,N_3124);
nor U4302 (N_4302,N_3316,N_3373);
nor U4303 (N_4303,N_3279,N_3639);
xor U4304 (N_4304,N_3534,N_3640);
nor U4305 (N_4305,N_3980,N_3290);
nand U4306 (N_4306,N_3602,N_3452);
and U4307 (N_4307,N_3518,N_3805);
nand U4308 (N_4308,N_3846,N_3362);
nor U4309 (N_4309,N_3257,N_3159);
nand U4310 (N_4310,N_3925,N_3968);
nor U4311 (N_4311,N_3513,N_3808);
nor U4312 (N_4312,N_3384,N_3605);
or U4313 (N_4313,N_3479,N_3345);
nor U4314 (N_4314,N_3752,N_3263);
and U4315 (N_4315,N_3350,N_3283);
nand U4316 (N_4316,N_3731,N_3248);
or U4317 (N_4317,N_3443,N_3488);
or U4318 (N_4318,N_3435,N_3013);
or U4319 (N_4319,N_3821,N_3069);
or U4320 (N_4320,N_3892,N_3195);
or U4321 (N_4321,N_3094,N_3372);
or U4322 (N_4322,N_3942,N_3199);
and U4323 (N_4323,N_3699,N_3780);
nor U4324 (N_4324,N_3928,N_3694);
nor U4325 (N_4325,N_3910,N_3909);
or U4326 (N_4326,N_3684,N_3670);
nor U4327 (N_4327,N_3682,N_3997);
nor U4328 (N_4328,N_3381,N_3305);
nor U4329 (N_4329,N_3459,N_3914);
and U4330 (N_4330,N_3189,N_3916);
and U4331 (N_4331,N_3676,N_3622);
nand U4332 (N_4332,N_3896,N_3620);
and U4333 (N_4333,N_3582,N_3842);
or U4334 (N_4334,N_3398,N_3113);
or U4335 (N_4335,N_3970,N_3619);
or U4336 (N_4336,N_3749,N_3599);
nor U4337 (N_4337,N_3377,N_3365);
and U4338 (N_4338,N_3447,N_3940);
or U4339 (N_4339,N_3463,N_3858);
nand U4340 (N_4340,N_3614,N_3432);
or U4341 (N_4341,N_3894,N_3695);
nor U4342 (N_4342,N_3064,N_3611);
and U4343 (N_4343,N_3792,N_3693);
nor U4344 (N_4344,N_3758,N_3902);
nand U4345 (N_4345,N_3176,N_3912);
xor U4346 (N_4346,N_3455,N_3794);
or U4347 (N_4347,N_3795,N_3742);
and U4348 (N_4348,N_3791,N_3696);
and U4349 (N_4349,N_3046,N_3593);
or U4350 (N_4350,N_3709,N_3024);
or U4351 (N_4351,N_3155,N_3662);
nand U4352 (N_4352,N_3151,N_3883);
and U4353 (N_4353,N_3125,N_3445);
nor U4354 (N_4354,N_3815,N_3923);
nor U4355 (N_4355,N_3818,N_3486);
nand U4356 (N_4356,N_3356,N_3723);
or U4357 (N_4357,N_3460,N_3240);
nand U4358 (N_4358,N_3060,N_3000);
or U4359 (N_4359,N_3765,N_3412);
nor U4360 (N_4360,N_3959,N_3392);
or U4361 (N_4361,N_3943,N_3242);
and U4362 (N_4362,N_3082,N_3043);
nand U4363 (N_4363,N_3164,N_3983);
nand U4364 (N_4364,N_3904,N_3409);
and U4365 (N_4365,N_3267,N_3870);
and U4366 (N_4366,N_3347,N_3783);
or U4367 (N_4367,N_3166,N_3207);
or U4368 (N_4368,N_3251,N_3586);
and U4369 (N_4369,N_3321,N_3229);
nor U4370 (N_4370,N_3243,N_3368);
and U4371 (N_4371,N_3274,N_3141);
or U4372 (N_4372,N_3171,N_3641);
nor U4373 (N_4373,N_3143,N_3358);
nand U4374 (N_4374,N_3636,N_3777);
nand U4375 (N_4375,N_3044,N_3228);
nor U4376 (N_4376,N_3798,N_3030);
and U4377 (N_4377,N_3034,N_3994);
nand U4378 (N_4378,N_3017,N_3965);
nand U4379 (N_4379,N_3090,N_3076);
and U4380 (N_4380,N_3134,N_3564);
nor U4381 (N_4381,N_3741,N_3497);
or U4382 (N_4382,N_3785,N_3413);
nor U4383 (N_4383,N_3931,N_3750);
nand U4384 (N_4384,N_3282,N_3117);
and U4385 (N_4385,N_3265,N_3483);
nor U4386 (N_4386,N_3104,N_3181);
nand U4387 (N_4387,N_3005,N_3981);
nand U4388 (N_4388,N_3768,N_3374);
or U4389 (N_4389,N_3149,N_3318);
nor U4390 (N_4390,N_3440,N_3021);
nand U4391 (N_4391,N_3180,N_3581);
xor U4392 (N_4392,N_3194,N_3702);
and U4393 (N_4393,N_3964,N_3817);
or U4394 (N_4394,N_3859,N_3371);
nand U4395 (N_4395,N_3077,N_3644);
or U4396 (N_4396,N_3738,N_3040);
nand U4397 (N_4397,N_3209,N_3559);
nor U4398 (N_4398,N_3273,N_3953);
nor U4399 (N_4399,N_3519,N_3056);
and U4400 (N_4400,N_3847,N_3999);
or U4401 (N_4401,N_3419,N_3913);
or U4402 (N_4402,N_3039,N_3408);
nand U4403 (N_4403,N_3324,N_3807);
nor U4404 (N_4404,N_3653,N_3937);
and U4405 (N_4405,N_3118,N_3604);
nand U4406 (N_4406,N_3958,N_3771);
and U4407 (N_4407,N_3938,N_3275);
or U4408 (N_4408,N_3838,N_3178);
and U4409 (N_4409,N_3264,N_3144);
and U4410 (N_4410,N_3052,N_3683);
and U4411 (N_4411,N_3081,N_3328);
or U4412 (N_4412,N_3778,N_3836);
or U4413 (N_4413,N_3532,N_3545);
nor U4414 (N_4414,N_3754,N_3106);
nor U4415 (N_4415,N_3446,N_3245);
nor U4416 (N_4416,N_3071,N_3291);
nor U4417 (N_4417,N_3135,N_3288);
nand U4418 (N_4418,N_3880,N_3418);
nand U4419 (N_4419,N_3007,N_3102);
nor U4420 (N_4420,N_3708,N_3388);
nor U4421 (N_4421,N_3072,N_3307);
or U4422 (N_4422,N_3225,N_3536);
or U4423 (N_4423,N_3098,N_3361);
or U4424 (N_4424,N_3982,N_3332);
or U4425 (N_4425,N_3174,N_3411);
nand U4426 (N_4426,N_3211,N_3660);
nor U4427 (N_4427,N_3111,N_3621);
nor U4428 (N_4428,N_3773,N_3222);
nor U4429 (N_4429,N_3774,N_3734);
nand U4430 (N_4430,N_3844,N_3317);
and U4431 (N_4431,N_3588,N_3340);
nor U4432 (N_4432,N_3610,N_3201);
nand U4433 (N_4433,N_3929,N_3839);
nand U4434 (N_4434,N_3210,N_3354);
or U4435 (N_4435,N_3541,N_3877);
and U4436 (N_4436,N_3574,N_3364);
nor U4437 (N_4437,N_3945,N_3112);
and U4438 (N_4438,N_3627,N_3558);
nand U4439 (N_4439,N_3990,N_3250);
nor U4440 (N_4440,N_3348,N_3675);
nand U4441 (N_4441,N_3570,N_3308);
and U4442 (N_4442,N_3423,N_3580);
and U4443 (N_4443,N_3867,N_3562);
or U4444 (N_4444,N_3539,N_3761);
nand U4445 (N_4445,N_3032,N_3200);
nand U4446 (N_4446,N_3946,N_3954);
nor U4447 (N_4447,N_3577,N_3341);
nand U4448 (N_4448,N_3120,N_3168);
or U4449 (N_4449,N_3260,N_3969);
nor U4450 (N_4450,N_3476,N_3936);
or U4451 (N_4451,N_3618,N_3114);
and U4452 (N_4452,N_3292,N_3091);
nand U4453 (N_4453,N_3217,N_3512);
and U4454 (N_4454,N_3607,N_3458);
xnor U4455 (N_4455,N_3227,N_3554);
and U4456 (N_4456,N_3197,N_3466);
and U4457 (N_4457,N_3508,N_3439);
nor U4458 (N_4458,N_3935,N_3658);
nor U4459 (N_4459,N_3170,N_3666);
nor U4460 (N_4460,N_3253,N_3673);
nand U4461 (N_4461,N_3779,N_3881);
or U4462 (N_4462,N_3678,N_3591);
nand U4463 (N_4463,N_3663,N_3109);
or U4464 (N_4464,N_3042,N_3302);
and U4465 (N_4465,N_3059,N_3103);
xnor U4466 (N_4466,N_3261,N_3510);
nor U4467 (N_4467,N_3864,N_3590);
and U4468 (N_4468,N_3029,N_3160);
nor U4469 (N_4469,N_3152,N_3163);
nor U4470 (N_4470,N_3911,N_3600);
and U4471 (N_4471,N_3309,N_3623);
or U4472 (N_4472,N_3575,N_3944);
or U4473 (N_4473,N_3218,N_3333);
nor U4474 (N_4474,N_3058,N_3538);
and U4475 (N_4475,N_3018,N_3074);
and U4476 (N_4476,N_3717,N_3158);
nand U4477 (N_4477,N_3511,N_3835);
and U4478 (N_4478,N_3996,N_3363);
nand U4479 (N_4479,N_3882,N_3376);
nand U4480 (N_4480,N_3226,N_3289);
nor U4481 (N_4481,N_3473,N_3776);
nand U4482 (N_4482,N_3352,N_3038);
nor U4483 (N_4483,N_3995,N_3806);
nand U4484 (N_4484,N_3391,N_3637);
nor U4485 (N_4485,N_3433,N_3487);
nor U4486 (N_4486,N_3428,N_3947);
or U4487 (N_4487,N_3079,N_3092);
and U4488 (N_4488,N_3136,N_3401);
nand U4489 (N_4489,N_3583,N_3325);
nor U4490 (N_4490,N_3716,N_3657);
and U4491 (N_4491,N_3691,N_3872);
and U4492 (N_4492,N_3003,N_3960);
and U4493 (N_4493,N_3587,N_3232);
nor U4494 (N_4494,N_3606,N_3165);
or U4495 (N_4495,N_3521,N_3086);
nor U4496 (N_4496,N_3255,N_3249);
or U4497 (N_4497,N_3028,N_3737);
and U4498 (N_4498,N_3422,N_3026);
and U4499 (N_4499,N_3179,N_3270);
nor U4500 (N_4500,N_3745,N_3035);
and U4501 (N_4501,N_3916,N_3739);
and U4502 (N_4502,N_3202,N_3296);
and U4503 (N_4503,N_3166,N_3084);
nand U4504 (N_4504,N_3572,N_3886);
nor U4505 (N_4505,N_3376,N_3080);
nand U4506 (N_4506,N_3053,N_3155);
nor U4507 (N_4507,N_3208,N_3110);
or U4508 (N_4508,N_3748,N_3115);
or U4509 (N_4509,N_3802,N_3138);
nor U4510 (N_4510,N_3010,N_3595);
or U4511 (N_4511,N_3497,N_3219);
or U4512 (N_4512,N_3756,N_3559);
nand U4513 (N_4513,N_3651,N_3889);
nand U4514 (N_4514,N_3781,N_3989);
nor U4515 (N_4515,N_3921,N_3766);
nand U4516 (N_4516,N_3757,N_3217);
nand U4517 (N_4517,N_3101,N_3573);
nor U4518 (N_4518,N_3614,N_3983);
nand U4519 (N_4519,N_3945,N_3923);
nand U4520 (N_4520,N_3978,N_3989);
or U4521 (N_4521,N_3899,N_3212);
nand U4522 (N_4522,N_3112,N_3594);
and U4523 (N_4523,N_3018,N_3620);
nand U4524 (N_4524,N_3428,N_3547);
nand U4525 (N_4525,N_3578,N_3096);
nor U4526 (N_4526,N_3731,N_3203);
nor U4527 (N_4527,N_3037,N_3359);
or U4528 (N_4528,N_3360,N_3974);
xnor U4529 (N_4529,N_3659,N_3301);
nor U4530 (N_4530,N_3179,N_3768);
xnor U4531 (N_4531,N_3673,N_3339);
or U4532 (N_4532,N_3489,N_3539);
nor U4533 (N_4533,N_3965,N_3736);
nand U4534 (N_4534,N_3902,N_3019);
xnor U4535 (N_4535,N_3614,N_3018);
nor U4536 (N_4536,N_3949,N_3751);
nor U4537 (N_4537,N_3451,N_3399);
and U4538 (N_4538,N_3522,N_3270);
nor U4539 (N_4539,N_3109,N_3202);
nand U4540 (N_4540,N_3173,N_3703);
nand U4541 (N_4541,N_3407,N_3566);
xor U4542 (N_4542,N_3038,N_3551);
nor U4543 (N_4543,N_3288,N_3463);
and U4544 (N_4544,N_3028,N_3720);
nor U4545 (N_4545,N_3220,N_3604);
or U4546 (N_4546,N_3439,N_3516);
or U4547 (N_4547,N_3220,N_3473);
nor U4548 (N_4548,N_3776,N_3564);
nor U4549 (N_4549,N_3915,N_3756);
or U4550 (N_4550,N_3110,N_3178);
nor U4551 (N_4551,N_3402,N_3342);
or U4552 (N_4552,N_3832,N_3055);
nor U4553 (N_4553,N_3268,N_3945);
nor U4554 (N_4554,N_3269,N_3196);
or U4555 (N_4555,N_3344,N_3129);
nor U4556 (N_4556,N_3105,N_3716);
nand U4557 (N_4557,N_3128,N_3952);
or U4558 (N_4558,N_3460,N_3554);
nor U4559 (N_4559,N_3258,N_3280);
nand U4560 (N_4560,N_3799,N_3844);
and U4561 (N_4561,N_3088,N_3370);
nand U4562 (N_4562,N_3737,N_3142);
nand U4563 (N_4563,N_3020,N_3523);
nor U4564 (N_4564,N_3655,N_3289);
or U4565 (N_4565,N_3744,N_3831);
or U4566 (N_4566,N_3771,N_3225);
and U4567 (N_4567,N_3195,N_3230);
nor U4568 (N_4568,N_3519,N_3748);
or U4569 (N_4569,N_3456,N_3864);
or U4570 (N_4570,N_3259,N_3579);
nand U4571 (N_4571,N_3027,N_3651);
and U4572 (N_4572,N_3055,N_3388);
nor U4573 (N_4573,N_3768,N_3134);
xnor U4574 (N_4574,N_3205,N_3948);
or U4575 (N_4575,N_3127,N_3341);
nand U4576 (N_4576,N_3122,N_3233);
nor U4577 (N_4577,N_3076,N_3629);
nor U4578 (N_4578,N_3870,N_3284);
and U4579 (N_4579,N_3877,N_3580);
nor U4580 (N_4580,N_3759,N_3764);
nor U4581 (N_4581,N_3735,N_3015);
and U4582 (N_4582,N_3469,N_3854);
nor U4583 (N_4583,N_3497,N_3402);
nand U4584 (N_4584,N_3099,N_3676);
or U4585 (N_4585,N_3913,N_3531);
nand U4586 (N_4586,N_3026,N_3603);
and U4587 (N_4587,N_3097,N_3668);
or U4588 (N_4588,N_3727,N_3014);
or U4589 (N_4589,N_3134,N_3602);
or U4590 (N_4590,N_3703,N_3377);
nand U4591 (N_4591,N_3762,N_3755);
nor U4592 (N_4592,N_3138,N_3953);
nand U4593 (N_4593,N_3306,N_3058);
or U4594 (N_4594,N_3833,N_3215);
nand U4595 (N_4595,N_3211,N_3396);
nand U4596 (N_4596,N_3664,N_3800);
nor U4597 (N_4597,N_3066,N_3740);
nand U4598 (N_4598,N_3143,N_3061);
or U4599 (N_4599,N_3702,N_3679);
or U4600 (N_4600,N_3134,N_3765);
nor U4601 (N_4601,N_3952,N_3581);
or U4602 (N_4602,N_3159,N_3752);
and U4603 (N_4603,N_3761,N_3686);
nand U4604 (N_4604,N_3018,N_3436);
and U4605 (N_4605,N_3091,N_3342);
nand U4606 (N_4606,N_3515,N_3359);
nor U4607 (N_4607,N_3724,N_3340);
or U4608 (N_4608,N_3850,N_3463);
or U4609 (N_4609,N_3016,N_3264);
and U4610 (N_4610,N_3867,N_3519);
nand U4611 (N_4611,N_3682,N_3593);
nand U4612 (N_4612,N_3824,N_3207);
nand U4613 (N_4613,N_3656,N_3017);
nand U4614 (N_4614,N_3084,N_3829);
nand U4615 (N_4615,N_3417,N_3262);
or U4616 (N_4616,N_3207,N_3015);
nand U4617 (N_4617,N_3861,N_3351);
nor U4618 (N_4618,N_3196,N_3120);
nand U4619 (N_4619,N_3653,N_3491);
or U4620 (N_4620,N_3481,N_3976);
nor U4621 (N_4621,N_3480,N_3565);
nand U4622 (N_4622,N_3229,N_3070);
nand U4623 (N_4623,N_3191,N_3682);
and U4624 (N_4624,N_3289,N_3860);
nor U4625 (N_4625,N_3499,N_3823);
or U4626 (N_4626,N_3704,N_3981);
nand U4627 (N_4627,N_3107,N_3166);
xor U4628 (N_4628,N_3595,N_3113);
or U4629 (N_4629,N_3994,N_3882);
and U4630 (N_4630,N_3399,N_3001);
and U4631 (N_4631,N_3028,N_3525);
nand U4632 (N_4632,N_3379,N_3565);
and U4633 (N_4633,N_3269,N_3164);
nor U4634 (N_4634,N_3159,N_3170);
and U4635 (N_4635,N_3511,N_3937);
or U4636 (N_4636,N_3178,N_3192);
nand U4637 (N_4637,N_3558,N_3211);
or U4638 (N_4638,N_3850,N_3718);
nor U4639 (N_4639,N_3183,N_3625);
nor U4640 (N_4640,N_3412,N_3267);
nand U4641 (N_4641,N_3418,N_3053);
and U4642 (N_4642,N_3549,N_3336);
or U4643 (N_4643,N_3749,N_3852);
and U4644 (N_4644,N_3556,N_3519);
and U4645 (N_4645,N_3617,N_3767);
nor U4646 (N_4646,N_3583,N_3592);
nand U4647 (N_4647,N_3720,N_3715);
or U4648 (N_4648,N_3326,N_3579);
nor U4649 (N_4649,N_3155,N_3485);
nand U4650 (N_4650,N_3225,N_3149);
or U4651 (N_4651,N_3733,N_3447);
or U4652 (N_4652,N_3003,N_3025);
and U4653 (N_4653,N_3272,N_3738);
nor U4654 (N_4654,N_3679,N_3897);
nor U4655 (N_4655,N_3559,N_3166);
or U4656 (N_4656,N_3927,N_3972);
or U4657 (N_4657,N_3843,N_3201);
nor U4658 (N_4658,N_3876,N_3478);
nand U4659 (N_4659,N_3740,N_3189);
nand U4660 (N_4660,N_3444,N_3201);
and U4661 (N_4661,N_3632,N_3241);
nor U4662 (N_4662,N_3573,N_3436);
and U4663 (N_4663,N_3402,N_3270);
or U4664 (N_4664,N_3765,N_3962);
and U4665 (N_4665,N_3351,N_3504);
nand U4666 (N_4666,N_3155,N_3266);
and U4667 (N_4667,N_3371,N_3477);
nor U4668 (N_4668,N_3002,N_3603);
or U4669 (N_4669,N_3410,N_3479);
xnor U4670 (N_4670,N_3788,N_3443);
or U4671 (N_4671,N_3879,N_3443);
nand U4672 (N_4672,N_3449,N_3208);
or U4673 (N_4673,N_3110,N_3545);
and U4674 (N_4674,N_3557,N_3393);
and U4675 (N_4675,N_3739,N_3271);
nand U4676 (N_4676,N_3503,N_3275);
nor U4677 (N_4677,N_3122,N_3368);
xnor U4678 (N_4678,N_3040,N_3127);
and U4679 (N_4679,N_3783,N_3877);
nand U4680 (N_4680,N_3987,N_3344);
nand U4681 (N_4681,N_3378,N_3685);
nand U4682 (N_4682,N_3247,N_3639);
and U4683 (N_4683,N_3297,N_3528);
and U4684 (N_4684,N_3228,N_3653);
or U4685 (N_4685,N_3983,N_3055);
or U4686 (N_4686,N_3205,N_3669);
xnor U4687 (N_4687,N_3236,N_3499);
and U4688 (N_4688,N_3613,N_3979);
or U4689 (N_4689,N_3311,N_3237);
and U4690 (N_4690,N_3567,N_3827);
nand U4691 (N_4691,N_3237,N_3275);
nand U4692 (N_4692,N_3510,N_3041);
and U4693 (N_4693,N_3268,N_3875);
nand U4694 (N_4694,N_3878,N_3059);
nor U4695 (N_4695,N_3348,N_3848);
nand U4696 (N_4696,N_3693,N_3969);
nor U4697 (N_4697,N_3709,N_3981);
nor U4698 (N_4698,N_3420,N_3392);
nor U4699 (N_4699,N_3694,N_3454);
nor U4700 (N_4700,N_3251,N_3397);
xor U4701 (N_4701,N_3482,N_3091);
or U4702 (N_4702,N_3133,N_3043);
and U4703 (N_4703,N_3431,N_3935);
nor U4704 (N_4704,N_3592,N_3939);
nand U4705 (N_4705,N_3999,N_3597);
nand U4706 (N_4706,N_3667,N_3143);
nor U4707 (N_4707,N_3171,N_3832);
or U4708 (N_4708,N_3055,N_3824);
nand U4709 (N_4709,N_3750,N_3807);
or U4710 (N_4710,N_3170,N_3462);
or U4711 (N_4711,N_3894,N_3653);
nor U4712 (N_4712,N_3263,N_3511);
nand U4713 (N_4713,N_3988,N_3660);
or U4714 (N_4714,N_3428,N_3101);
nor U4715 (N_4715,N_3311,N_3728);
or U4716 (N_4716,N_3159,N_3547);
xor U4717 (N_4717,N_3316,N_3085);
and U4718 (N_4718,N_3773,N_3762);
or U4719 (N_4719,N_3153,N_3464);
and U4720 (N_4720,N_3980,N_3869);
and U4721 (N_4721,N_3933,N_3546);
nor U4722 (N_4722,N_3461,N_3105);
and U4723 (N_4723,N_3076,N_3009);
xnor U4724 (N_4724,N_3989,N_3144);
nor U4725 (N_4725,N_3514,N_3051);
nor U4726 (N_4726,N_3882,N_3940);
or U4727 (N_4727,N_3618,N_3698);
and U4728 (N_4728,N_3214,N_3700);
nand U4729 (N_4729,N_3185,N_3642);
nor U4730 (N_4730,N_3982,N_3885);
nand U4731 (N_4731,N_3734,N_3059);
nand U4732 (N_4732,N_3837,N_3295);
nor U4733 (N_4733,N_3002,N_3663);
and U4734 (N_4734,N_3998,N_3516);
nor U4735 (N_4735,N_3762,N_3529);
nor U4736 (N_4736,N_3741,N_3753);
and U4737 (N_4737,N_3203,N_3609);
nor U4738 (N_4738,N_3464,N_3724);
nor U4739 (N_4739,N_3786,N_3971);
xnor U4740 (N_4740,N_3759,N_3103);
and U4741 (N_4741,N_3895,N_3309);
xor U4742 (N_4742,N_3168,N_3261);
and U4743 (N_4743,N_3630,N_3670);
nor U4744 (N_4744,N_3315,N_3801);
and U4745 (N_4745,N_3910,N_3003);
nor U4746 (N_4746,N_3476,N_3782);
nor U4747 (N_4747,N_3584,N_3491);
and U4748 (N_4748,N_3301,N_3246);
nand U4749 (N_4749,N_3327,N_3261);
nor U4750 (N_4750,N_3312,N_3084);
nand U4751 (N_4751,N_3587,N_3229);
or U4752 (N_4752,N_3383,N_3322);
and U4753 (N_4753,N_3819,N_3620);
nor U4754 (N_4754,N_3879,N_3882);
and U4755 (N_4755,N_3800,N_3436);
nand U4756 (N_4756,N_3659,N_3027);
and U4757 (N_4757,N_3265,N_3119);
nor U4758 (N_4758,N_3903,N_3862);
or U4759 (N_4759,N_3764,N_3997);
nand U4760 (N_4760,N_3030,N_3698);
or U4761 (N_4761,N_3268,N_3284);
nand U4762 (N_4762,N_3473,N_3725);
nor U4763 (N_4763,N_3352,N_3129);
or U4764 (N_4764,N_3350,N_3494);
nor U4765 (N_4765,N_3759,N_3871);
nand U4766 (N_4766,N_3203,N_3603);
nand U4767 (N_4767,N_3241,N_3760);
and U4768 (N_4768,N_3287,N_3135);
nand U4769 (N_4769,N_3321,N_3017);
nor U4770 (N_4770,N_3854,N_3415);
xnor U4771 (N_4771,N_3028,N_3808);
and U4772 (N_4772,N_3929,N_3999);
nor U4773 (N_4773,N_3352,N_3619);
and U4774 (N_4774,N_3507,N_3855);
nor U4775 (N_4775,N_3675,N_3901);
or U4776 (N_4776,N_3869,N_3224);
or U4777 (N_4777,N_3483,N_3777);
nor U4778 (N_4778,N_3316,N_3960);
nand U4779 (N_4779,N_3215,N_3217);
or U4780 (N_4780,N_3400,N_3606);
or U4781 (N_4781,N_3869,N_3360);
and U4782 (N_4782,N_3283,N_3780);
or U4783 (N_4783,N_3699,N_3494);
nor U4784 (N_4784,N_3843,N_3498);
or U4785 (N_4785,N_3925,N_3646);
or U4786 (N_4786,N_3235,N_3812);
nor U4787 (N_4787,N_3945,N_3994);
nand U4788 (N_4788,N_3529,N_3861);
nor U4789 (N_4789,N_3221,N_3118);
nor U4790 (N_4790,N_3700,N_3906);
nand U4791 (N_4791,N_3172,N_3436);
nor U4792 (N_4792,N_3317,N_3975);
and U4793 (N_4793,N_3037,N_3926);
and U4794 (N_4794,N_3239,N_3144);
nor U4795 (N_4795,N_3906,N_3124);
nor U4796 (N_4796,N_3993,N_3671);
or U4797 (N_4797,N_3284,N_3317);
or U4798 (N_4798,N_3388,N_3526);
nor U4799 (N_4799,N_3671,N_3099);
nor U4800 (N_4800,N_3433,N_3280);
and U4801 (N_4801,N_3753,N_3469);
nor U4802 (N_4802,N_3775,N_3104);
or U4803 (N_4803,N_3791,N_3153);
nor U4804 (N_4804,N_3691,N_3794);
and U4805 (N_4805,N_3617,N_3800);
or U4806 (N_4806,N_3592,N_3953);
or U4807 (N_4807,N_3221,N_3282);
nand U4808 (N_4808,N_3033,N_3934);
or U4809 (N_4809,N_3556,N_3587);
and U4810 (N_4810,N_3314,N_3369);
and U4811 (N_4811,N_3677,N_3054);
nor U4812 (N_4812,N_3742,N_3337);
and U4813 (N_4813,N_3523,N_3550);
or U4814 (N_4814,N_3043,N_3681);
and U4815 (N_4815,N_3579,N_3296);
or U4816 (N_4816,N_3302,N_3321);
nor U4817 (N_4817,N_3583,N_3107);
nor U4818 (N_4818,N_3442,N_3910);
nor U4819 (N_4819,N_3294,N_3339);
and U4820 (N_4820,N_3702,N_3584);
nor U4821 (N_4821,N_3540,N_3446);
nand U4822 (N_4822,N_3256,N_3447);
and U4823 (N_4823,N_3771,N_3260);
nor U4824 (N_4824,N_3445,N_3972);
or U4825 (N_4825,N_3517,N_3865);
or U4826 (N_4826,N_3044,N_3780);
xnor U4827 (N_4827,N_3227,N_3840);
or U4828 (N_4828,N_3760,N_3254);
and U4829 (N_4829,N_3857,N_3852);
or U4830 (N_4830,N_3289,N_3888);
or U4831 (N_4831,N_3434,N_3474);
nand U4832 (N_4832,N_3572,N_3270);
nand U4833 (N_4833,N_3571,N_3687);
nor U4834 (N_4834,N_3538,N_3045);
or U4835 (N_4835,N_3877,N_3202);
or U4836 (N_4836,N_3385,N_3438);
nand U4837 (N_4837,N_3631,N_3358);
and U4838 (N_4838,N_3924,N_3371);
nor U4839 (N_4839,N_3817,N_3197);
or U4840 (N_4840,N_3201,N_3928);
nand U4841 (N_4841,N_3707,N_3329);
nor U4842 (N_4842,N_3170,N_3106);
nor U4843 (N_4843,N_3383,N_3321);
nor U4844 (N_4844,N_3343,N_3097);
nor U4845 (N_4845,N_3475,N_3039);
nor U4846 (N_4846,N_3534,N_3557);
and U4847 (N_4847,N_3877,N_3768);
xor U4848 (N_4848,N_3812,N_3809);
nor U4849 (N_4849,N_3233,N_3529);
nor U4850 (N_4850,N_3747,N_3507);
or U4851 (N_4851,N_3419,N_3955);
nand U4852 (N_4852,N_3353,N_3578);
nor U4853 (N_4853,N_3626,N_3095);
or U4854 (N_4854,N_3399,N_3991);
and U4855 (N_4855,N_3691,N_3554);
and U4856 (N_4856,N_3850,N_3624);
nor U4857 (N_4857,N_3218,N_3134);
and U4858 (N_4858,N_3647,N_3888);
or U4859 (N_4859,N_3027,N_3896);
nor U4860 (N_4860,N_3593,N_3148);
or U4861 (N_4861,N_3133,N_3961);
and U4862 (N_4862,N_3029,N_3594);
and U4863 (N_4863,N_3636,N_3972);
nand U4864 (N_4864,N_3568,N_3635);
nand U4865 (N_4865,N_3202,N_3730);
xnor U4866 (N_4866,N_3988,N_3731);
or U4867 (N_4867,N_3380,N_3296);
or U4868 (N_4868,N_3228,N_3754);
nand U4869 (N_4869,N_3045,N_3610);
nand U4870 (N_4870,N_3917,N_3996);
nor U4871 (N_4871,N_3800,N_3199);
and U4872 (N_4872,N_3625,N_3759);
and U4873 (N_4873,N_3976,N_3559);
nand U4874 (N_4874,N_3220,N_3961);
nand U4875 (N_4875,N_3257,N_3273);
nand U4876 (N_4876,N_3152,N_3412);
and U4877 (N_4877,N_3230,N_3551);
nand U4878 (N_4878,N_3590,N_3611);
nor U4879 (N_4879,N_3584,N_3047);
or U4880 (N_4880,N_3131,N_3786);
nor U4881 (N_4881,N_3307,N_3704);
and U4882 (N_4882,N_3774,N_3163);
nor U4883 (N_4883,N_3540,N_3408);
nand U4884 (N_4884,N_3063,N_3246);
and U4885 (N_4885,N_3789,N_3425);
and U4886 (N_4886,N_3836,N_3837);
or U4887 (N_4887,N_3268,N_3394);
or U4888 (N_4888,N_3887,N_3224);
and U4889 (N_4889,N_3070,N_3905);
or U4890 (N_4890,N_3247,N_3176);
and U4891 (N_4891,N_3968,N_3553);
nor U4892 (N_4892,N_3285,N_3775);
nand U4893 (N_4893,N_3084,N_3430);
nor U4894 (N_4894,N_3264,N_3461);
nor U4895 (N_4895,N_3107,N_3958);
nand U4896 (N_4896,N_3930,N_3002);
and U4897 (N_4897,N_3879,N_3517);
nor U4898 (N_4898,N_3059,N_3369);
and U4899 (N_4899,N_3412,N_3542);
or U4900 (N_4900,N_3900,N_3725);
and U4901 (N_4901,N_3782,N_3982);
or U4902 (N_4902,N_3076,N_3491);
and U4903 (N_4903,N_3801,N_3514);
nand U4904 (N_4904,N_3794,N_3470);
or U4905 (N_4905,N_3538,N_3931);
or U4906 (N_4906,N_3736,N_3396);
nor U4907 (N_4907,N_3594,N_3658);
and U4908 (N_4908,N_3994,N_3918);
and U4909 (N_4909,N_3635,N_3002);
nor U4910 (N_4910,N_3066,N_3089);
or U4911 (N_4911,N_3951,N_3121);
nand U4912 (N_4912,N_3294,N_3999);
nand U4913 (N_4913,N_3184,N_3399);
nand U4914 (N_4914,N_3008,N_3017);
nor U4915 (N_4915,N_3490,N_3310);
and U4916 (N_4916,N_3663,N_3219);
or U4917 (N_4917,N_3267,N_3098);
nand U4918 (N_4918,N_3154,N_3266);
nand U4919 (N_4919,N_3001,N_3537);
and U4920 (N_4920,N_3712,N_3720);
and U4921 (N_4921,N_3833,N_3160);
or U4922 (N_4922,N_3303,N_3105);
and U4923 (N_4923,N_3115,N_3717);
nand U4924 (N_4924,N_3271,N_3757);
and U4925 (N_4925,N_3448,N_3393);
nand U4926 (N_4926,N_3847,N_3316);
or U4927 (N_4927,N_3653,N_3146);
nand U4928 (N_4928,N_3928,N_3510);
or U4929 (N_4929,N_3646,N_3335);
nand U4930 (N_4930,N_3841,N_3134);
nand U4931 (N_4931,N_3950,N_3646);
or U4932 (N_4932,N_3626,N_3860);
and U4933 (N_4933,N_3257,N_3758);
or U4934 (N_4934,N_3316,N_3835);
and U4935 (N_4935,N_3659,N_3447);
or U4936 (N_4936,N_3919,N_3170);
or U4937 (N_4937,N_3780,N_3167);
and U4938 (N_4938,N_3583,N_3286);
nand U4939 (N_4939,N_3925,N_3546);
or U4940 (N_4940,N_3232,N_3983);
nor U4941 (N_4941,N_3135,N_3146);
or U4942 (N_4942,N_3632,N_3813);
or U4943 (N_4943,N_3951,N_3393);
nand U4944 (N_4944,N_3625,N_3546);
nor U4945 (N_4945,N_3772,N_3503);
xor U4946 (N_4946,N_3961,N_3019);
nand U4947 (N_4947,N_3227,N_3907);
nand U4948 (N_4948,N_3886,N_3668);
or U4949 (N_4949,N_3390,N_3029);
or U4950 (N_4950,N_3552,N_3749);
nor U4951 (N_4951,N_3605,N_3904);
nand U4952 (N_4952,N_3968,N_3628);
or U4953 (N_4953,N_3816,N_3350);
nor U4954 (N_4954,N_3790,N_3996);
and U4955 (N_4955,N_3887,N_3479);
nor U4956 (N_4956,N_3828,N_3005);
nand U4957 (N_4957,N_3531,N_3631);
nor U4958 (N_4958,N_3851,N_3675);
xnor U4959 (N_4959,N_3130,N_3923);
nor U4960 (N_4960,N_3837,N_3155);
nand U4961 (N_4961,N_3112,N_3259);
nor U4962 (N_4962,N_3355,N_3899);
or U4963 (N_4963,N_3673,N_3041);
or U4964 (N_4964,N_3245,N_3113);
nand U4965 (N_4965,N_3094,N_3841);
and U4966 (N_4966,N_3035,N_3685);
nor U4967 (N_4967,N_3674,N_3748);
and U4968 (N_4968,N_3955,N_3135);
nand U4969 (N_4969,N_3109,N_3562);
or U4970 (N_4970,N_3132,N_3988);
nor U4971 (N_4971,N_3376,N_3709);
nand U4972 (N_4972,N_3357,N_3556);
nand U4973 (N_4973,N_3341,N_3356);
or U4974 (N_4974,N_3757,N_3572);
or U4975 (N_4975,N_3264,N_3898);
or U4976 (N_4976,N_3350,N_3906);
nor U4977 (N_4977,N_3363,N_3726);
nor U4978 (N_4978,N_3764,N_3827);
and U4979 (N_4979,N_3015,N_3329);
nor U4980 (N_4980,N_3220,N_3082);
or U4981 (N_4981,N_3988,N_3561);
and U4982 (N_4982,N_3148,N_3587);
nor U4983 (N_4983,N_3094,N_3248);
nand U4984 (N_4984,N_3405,N_3788);
and U4985 (N_4985,N_3335,N_3316);
nor U4986 (N_4986,N_3479,N_3758);
and U4987 (N_4987,N_3953,N_3893);
or U4988 (N_4988,N_3118,N_3316);
or U4989 (N_4989,N_3108,N_3376);
and U4990 (N_4990,N_3756,N_3217);
or U4991 (N_4991,N_3422,N_3216);
nor U4992 (N_4992,N_3421,N_3325);
or U4993 (N_4993,N_3338,N_3206);
nor U4994 (N_4994,N_3248,N_3193);
and U4995 (N_4995,N_3045,N_3895);
or U4996 (N_4996,N_3557,N_3981);
and U4997 (N_4997,N_3420,N_3537);
or U4998 (N_4998,N_3947,N_3141);
nand U4999 (N_4999,N_3009,N_3781);
or U5000 (N_5000,N_4032,N_4875);
nor U5001 (N_5001,N_4444,N_4918);
or U5002 (N_5002,N_4248,N_4895);
nor U5003 (N_5003,N_4637,N_4643);
nor U5004 (N_5004,N_4971,N_4791);
nor U5005 (N_5005,N_4126,N_4221);
or U5006 (N_5006,N_4404,N_4225);
or U5007 (N_5007,N_4164,N_4828);
and U5008 (N_5008,N_4131,N_4217);
nand U5009 (N_5009,N_4072,N_4878);
nor U5010 (N_5010,N_4325,N_4832);
nor U5011 (N_5011,N_4201,N_4142);
or U5012 (N_5012,N_4863,N_4845);
and U5013 (N_5013,N_4240,N_4665);
and U5014 (N_5014,N_4502,N_4384);
nor U5015 (N_5015,N_4298,N_4912);
nor U5016 (N_5016,N_4563,N_4631);
or U5017 (N_5017,N_4544,N_4997);
and U5018 (N_5018,N_4046,N_4380);
and U5019 (N_5019,N_4901,N_4717);
and U5020 (N_5020,N_4408,N_4242);
nand U5021 (N_5021,N_4497,N_4396);
nand U5022 (N_5022,N_4690,N_4733);
or U5023 (N_5023,N_4926,N_4840);
nor U5024 (N_5024,N_4587,N_4740);
nor U5025 (N_5025,N_4282,N_4602);
and U5026 (N_5026,N_4769,N_4513);
nand U5027 (N_5027,N_4180,N_4522);
and U5028 (N_5028,N_4102,N_4741);
or U5029 (N_5029,N_4434,N_4146);
and U5030 (N_5030,N_4361,N_4367);
nand U5031 (N_5031,N_4711,N_4600);
nor U5032 (N_5032,N_4705,N_4662);
and U5033 (N_5033,N_4684,N_4827);
nor U5034 (N_5034,N_4567,N_4512);
or U5035 (N_5035,N_4830,N_4945);
or U5036 (N_5036,N_4871,N_4825);
nor U5037 (N_5037,N_4556,N_4419);
nand U5038 (N_5038,N_4105,N_4610);
or U5039 (N_5039,N_4036,N_4682);
nand U5040 (N_5040,N_4211,N_4215);
nand U5041 (N_5041,N_4383,N_4999);
nand U5042 (N_5042,N_4039,N_4420);
nor U5043 (N_5043,N_4286,N_4317);
nand U5044 (N_5044,N_4862,N_4781);
nand U5045 (N_5045,N_4532,N_4223);
nor U5046 (N_5046,N_4641,N_4509);
nand U5047 (N_5047,N_4961,N_4341);
and U5048 (N_5048,N_4043,N_4307);
nand U5049 (N_5049,N_4392,N_4692);
nor U5050 (N_5050,N_4698,N_4375);
and U5051 (N_5051,N_4757,N_4937);
and U5052 (N_5052,N_4776,N_4707);
nand U5053 (N_5053,N_4730,N_4909);
or U5054 (N_5054,N_4951,N_4274);
and U5055 (N_5055,N_4054,N_4089);
or U5056 (N_5056,N_4818,N_4988);
nor U5057 (N_5057,N_4887,N_4750);
nor U5058 (N_5058,N_4449,N_4321);
nand U5059 (N_5059,N_4800,N_4172);
nand U5060 (N_5060,N_4499,N_4721);
and U5061 (N_5061,N_4447,N_4680);
nand U5062 (N_5062,N_4629,N_4122);
nand U5063 (N_5063,N_4946,N_4084);
or U5064 (N_5064,N_4272,N_4255);
nand U5065 (N_5065,N_4473,N_4922);
or U5066 (N_5066,N_4930,N_4134);
xnor U5067 (N_5067,N_4468,N_4273);
or U5068 (N_5068,N_4149,N_4914);
and U5069 (N_5069,N_4552,N_4656);
xnor U5070 (N_5070,N_4899,N_4026);
nand U5071 (N_5071,N_4749,N_4715);
or U5072 (N_5072,N_4919,N_4572);
and U5073 (N_5073,N_4984,N_4271);
nor U5074 (N_5074,N_4695,N_4894);
and U5075 (N_5075,N_4127,N_4132);
nor U5076 (N_5076,N_4306,N_4472);
nand U5077 (N_5077,N_4068,N_4344);
nor U5078 (N_5078,N_4836,N_4826);
or U5079 (N_5079,N_4435,N_4837);
nand U5080 (N_5080,N_4718,N_4940);
or U5081 (N_5081,N_4753,N_4652);
nand U5082 (N_5082,N_4374,N_4927);
or U5083 (N_5083,N_4719,N_4989);
and U5084 (N_5084,N_4446,N_4051);
and U5085 (N_5085,N_4152,N_4070);
nor U5086 (N_5086,N_4017,N_4167);
or U5087 (N_5087,N_4429,N_4492);
nand U5088 (N_5088,N_4364,N_4906);
and U5089 (N_5089,N_4183,N_4520);
nand U5090 (N_5090,N_4693,N_4474);
and U5091 (N_5091,N_4237,N_4409);
nand U5092 (N_5092,N_4751,N_4424);
nor U5093 (N_5093,N_4639,N_4041);
or U5094 (N_5094,N_4091,N_4100);
nand U5095 (N_5095,N_4397,N_4066);
nor U5096 (N_5096,N_4571,N_4580);
nor U5097 (N_5097,N_4523,N_4574);
nor U5098 (N_5098,N_4959,N_4583);
and U5099 (N_5099,N_4978,N_4780);
nand U5100 (N_5100,N_4075,N_4889);
or U5101 (N_5101,N_4943,N_4853);
or U5102 (N_5102,N_4345,N_4597);
nand U5103 (N_5103,N_4599,N_4977);
and U5104 (N_5104,N_4963,N_4213);
nand U5105 (N_5105,N_4592,N_4713);
or U5106 (N_5106,N_4209,N_4170);
nor U5107 (N_5107,N_4445,N_4924);
nor U5108 (N_5108,N_4014,N_4994);
or U5109 (N_5109,N_4003,N_4353);
nor U5110 (N_5110,N_4253,N_4803);
xor U5111 (N_5111,N_4260,N_4030);
or U5112 (N_5112,N_4726,N_4033);
nand U5113 (N_5113,N_4355,N_4337);
nor U5114 (N_5114,N_4107,N_4722);
or U5115 (N_5115,N_4542,N_4136);
nand U5116 (N_5116,N_4839,N_4621);
and U5117 (N_5117,N_4179,N_4056);
nand U5118 (N_5118,N_4627,N_4254);
or U5119 (N_5119,N_4511,N_4328);
nor U5120 (N_5120,N_4302,N_4773);
or U5121 (N_5121,N_4723,N_4967);
nand U5122 (N_5122,N_4159,N_4354);
or U5123 (N_5123,N_4866,N_4276);
nor U5124 (N_5124,N_4885,N_4049);
nor U5125 (N_5125,N_4890,N_4139);
and U5126 (N_5126,N_4288,N_4615);
nor U5127 (N_5127,N_4299,N_4281);
nand U5128 (N_5128,N_4864,N_4881);
nand U5129 (N_5129,N_4547,N_4261);
or U5130 (N_5130,N_4078,N_4736);
nand U5131 (N_5131,N_4086,N_4324);
or U5132 (N_5132,N_4934,N_4188);
nand U5133 (N_5133,N_4311,N_4764);
and U5134 (N_5134,N_4475,N_4203);
nor U5135 (N_5135,N_4913,N_4809);
or U5136 (N_5136,N_4193,N_4888);
nor U5137 (N_5137,N_4331,N_4505);
and U5138 (N_5138,N_4731,N_4168);
nor U5139 (N_5139,N_4326,N_4679);
nor U5140 (N_5140,N_4413,N_4130);
and U5141 (N_5141,N_4290,N_4148);
nor U5142 (N_5142,N_4504,N_4605);
nand U5143 (N_5143,N_4280,N_4391);
nor U5144 (N_5144,N_4891,N_4099);
nor U5145 (N_5145,N_4467,N_4378);
or U5146 (N_5146,N_4027,N_4441);
nand U5147 (N_5147,N_4759,N_4227);
and U5148 (N_5148,N_4442,N_4111);
and U5149 (N_5149,N_4038,N_4287);
or U5150 (N_5150,N_4647,N_4606);
nand U5151 (N_5151,N_4969,N_4297);
or U5152 (N_5152,N_4974,N_4857);
or U5153 (N_5153,N_4941,N_4028);
nand U5154 (N_5154,N_4990,N_4716);
or U5155 (N_5155,N_4305,N_4524);
or U5156 (N_5156,N_4729,N_4438);
or U5157 (N_5157,N_4867,N_4493);
nand U5158 (N_5158,N_4477,N_4192);
nand U5159 (N_5159,N_4898,N_4085);
nor U5160 (N_5160,N_4976,N_4601);
or U5161 (N_5161,N_4060,N_4938);
nor U5162 (N_5162,N_4115,N_4576);
or U5163 (N_5163,N_4902,N_4772);
and U5164 (N_5164,N_4655,N_4121);
and U5165 (N_5165,N_4246,N_4229);
or U5166 (N_5166,N_4171,N_4588);
nand U5167 (N_5167,N_4784,N_4048);
nor U5168 (N_5168,N_4155,N_4425);
nand U5169 (N_5169,N_4980,N_4573);
or U5170 (N_5170,N_4158,N_4151);
nand U5171 (N_5171,N_4598,N_4373);
nor U5172 (N_5172,N_4376,N_4120);
and U5173 (N_5173,N_4019,N_4702);
nor U5174 (N_5174,N_4470,N_4917);
nand U5175 (N_5175,N_4503,N_4205);
or U5176 (N_5176,N_4042,N_4029);
nor U5177 (N_5177,N_4135,N_4212);
or U5178 (N_5178,N_4521,N_4338);
nor U5179 (N_5179,N_4559,N_4986);
nor U5180 (N_5180,N_4362,N_4834);
nor U5181 (N_5181,N_4628,N_4219);
and U5182 (N_5182,N_4058,N_4916);
or U5183 (N_5183,N_4765,N_4357);
and U5184 (N_5184,N_4400,N_4358);
and U5185 (N_5185,N_4284,N_4744);
nor U5186 (N_5186,N_4880,N_4451);
nor U5187 (N_5187,N_4103,N_4322);
or U5188 (N_5188,N_4265,N_4398);
or U5189 (N_5189,N_4390,N_4972);
nor U5190 (N_5190,N_4023,N_4402);
nand U5191 (N_5191,N_4195,N_4300);
nor U5192 (N_5192,N_4482,N_4113);
or U5193 (N_5193,N_4316,N_4549);
nor U5194 (N_5194,N_4208,N_4604);
nor U5195 (N_5195,N_4868,N_4092);
nand U5196 (N_5196,N_4896,N_4388);
nand U5197 (N_5197,N_4098,N_4104);
and U5198 (N_5198,N_4275,N_4418);
nor U5199 (N_5199,N_4983,N_4040);
nor U5200 (N_5200,N_4794,N_4793);
and U5201 (N_5201,N_4329,N_4238);
or U5202 (N_5202,N_4557,N_4256);
nor U5203 (N_5203,N_4385,N_4709);
or U5204 (N_5204,N_4622,N_4579);
or U5205 (N_5205,N_4489,N_4634);
nor U5206 (N_5206,N_4071,N_4452);
and U5207 (N_5207,N_4423,N_4401);
nand U5208 (N_5208,N_4194,N_4775);
or U5209 (N_5209,N_4654,N_4844);
nand U5210 (N_5210,N_4154,N_4987);
nand U5211 (N_5211,N_4998,N_4675);
and U5212 (N_5212,N_4389,N_4935);
nor U5213 (N_5213,N_4703,N_4620);
and U5214 (N_5214,N_4739,N_4228);
nand U5215 (N_5215,N_4767,N_4245);
and U5216 (N_5216,N_4189,N_4525);
and U5217 (N_5217,N_4727,N_4301);
nor U5218 (N_5218,N_4488,N_4143);
or U5219 (N_5219,N_4197,N_4437);
nor U5220 (N_5220,N_4309,N_4796);
and U5221 (N_5221,N_4562,N_4187);
and U5222 (N_5222,N_4607,N_4979);
and U5223 (N_5223,N_4578,N_4960);
nor U5224 (N_5224,N_4821,N_4348);
and U5225 (N_5225,N_4096,N_4267);
or U5226 (N_5226,N_4176,N_4507);
nor U5227 (N_5227,N_4965,N_4632);
or U5228 (N_5228,N_4911,N_4701);
and U5229 (N_5229,N_4589,N_4625);
or U5230 (N_5230,N_4145,N_4169);
and U5231 (N_5231,N_4982,N_4590);
and U5232 (N_5232,N_4585,N_4529);
nor U5233 (N_5233,N_4216,N_4761);
or U5234 (N_5234,N_4732,N_4500);
nand U5235 (N_5235,N_4519,N_4285);
nor U5236 (N_5236,N_4514,N_4182);
nand U5237 (N_5237,N_4231,N_4462);
nor U5238 (N_5238,N_4820,N_4101);
nor U5239 (N_5239,N_4683,N_4806);
and U5240 (N_5240,N_4932,N_4005);
nand U5241 (N_5241,N_4463,N_4431);
and U5242 (N_5242,N_4414,N_4697);
nand U5243 (N_5243,N_4185,N_4200);
nor U5244 (N_5244,N_4907,N_4584);
nor U5245 (N_5245,N_4365,N_4668);
and U5246 (N_5246,N_4735,N_4886);
xnor U5247 (N_5247,N_4905,N_4903);
nand U5248 (N_5248,N_4882,N_4289);
or U5249 (N_5249,N_4291,N_4710);
and U5250 (N_5250,N_4817,N_4777);
nand U5251 (N_5251,N_4560,N_4128);
or U5252 (N_5252,N_4129,N_4498);
nand U5253 (N_5253,N_4947,N_4696);
and U5254 (N_5254,N_4214,N_4320);
nand U5255 (N_5255,N_4869,N_4861);
or U5256 (N_5256,N_4411,N_4024);
nor U5257 (N_5257,N_4269,N_4531);
or U5258 (N_5258,N_4277,N_4177);
xnor U5259 (N_5259,N_4161,N_4993);
and U5260 (N_5260,N_4457,N_4884);
or U5261 (N_5261,N_4966,N_4190);
nand U5262 (N_5262,N_4856,N_4671);
nand U5263 (N_5263,N_4021,N_4802);
nand U5264 (N_5264,N_4700,N_4065);
or U5265 (N_5265,N_4008,N_4184);
and U5266 (N_5266,N_4007,N_4748);
and U5267 (N_5267,N_4642,N_4659);
and U5268 (N_5268,N_4530,N_4422);
and U5269 (N_5269,N_4816,N_4236);
nor U5270 (N_5270,N_4268,N_4510);
xnor U5271 (N_5271,N_4546,N_4336);
nand U5272 (N_5272,N_4714,N_4553);
and U5273 (N_5273,N_4681,N_4343);
nor U5274 (N_5274,N_4224,N_4165);
or U5275 (N_5275,N_4076,N_4063);
or U5276 (N_5276,N_4910,N_4543);
nor U5277 (N_5277,N_4819,N_4855);
nand U5278 (N_5278,N_4694,N_4724);
and U5279 (N_5279,N_4258,N_4677);
nor U5280 (N_5280,N_4031,N_4985);
and U5281 (N_5281,N_4279,N_4570);
nor U5282 (N_5282,N_4555,N_4953);
and U5283 (N_5283,N_4371,N_4596);
or U5284 (N_5284,N_4412,N_4178);
or U5285 (N_5285,N_4110,N_4015);
or U5286 (N_5286,N_4252,N_4807);
nor U5287 (N_5287,N_4251,N_4518);
nor U5288 (N_5288,N_4421,N_4929);
nor U5289 (N_5289,N_4323,N_4097);
nor U5290 (N_5290,N_4480,N_4439);
nor U5291 (N_5291,N_4673,N_4053);
or U5292 (N_5292,N_4814,N_4846);
or U5293 (N_5293,N_4250,N_4619);
or U5294 (N_5294,N_4395,N_4350);
or U5295 (N_5295,N_4339,N_4900);
or U5296 (N_5296,N_4405,N_4244);
or U5297 (N_5297,N_4202,N_4624);
or U5298 (N_5298,N_4931,N_4204);
or U5299 (N_5299,N_4756,N_4897);
nor U5300 (N_5300,N_4270,N_4633);
or U5301 (N_5301,N_4372,N_4550);
nand U5302 (N_5302,N_4640,N_4535);
and U5303 (N_5303,N_4018,N_4226);
nor U5304 (N_5304,N_4013,N_4332);
nand U5305 (N_5305,N_4537,N_4783);
nor U5306 (N_5306,N_4181,N_4660);
nand U5307 (N_5307,N_4688,N_4558);
or U5308 (N_5308,N_4786,N_4370);
nor U5309 (N_5309,N_4992,N_4737);
or U5310 (N_5310,N_4536,N_4568);
xor U5311 (N_5311,N_4137,N_4407);
or U5312 (N_5312,N_4991,N_4594);
nand U5313 (N_5313,N_4812,N_4908);
and U5314 (N_5314,N_4108,N_4808);
nor U5315 (N_5315,N_4936,N_4118);
nand U5316 (N_5316,N_4327,N_4533);
nand U5317 (N_5317,N_4426,N_4232);
nor U5318 (N_5318,N_4958,N_4798);
or U5319 (N_5319,N_4645,N_4491);
xor U5320 (N_5320,N_4481,N_4319);
nor U5321 (N_5321,N_4174,N_4062);
nor U5322 (N_5322,N_4487,N_4415);
nand U5323 (N_5323,N_4312,N_4849);
or U5324 (N_5324,N_4883,N_4460);
or U5325 (N_5325,N_4313,N_4548);
nand U5326 (N_5326,N_4506,N_4790);
nor U5327 (N_5327,N_4904,N_4626);
or U5328 (N_5328,N_4870,N_4330);
nor U5329 (N_5329,N_4768,N_4554);
xor U5330 (N_5330,N_4801,N_4067);
or U5331 (N_5331,N_4581,N_4459);
nor U5332 (N_5332,N_4792,N_4090);
or U5333 (N_5333,N_4484,N_4379);
nand U5334 (N_5334,N_4293,N_4386);
and U5335 (N_5335,N_4725,N_4047);
nand U5336 (N_5336,N_4476,N_4050);
or U5337 (N_5337,N_4608,N_4763);
and U5338 (N_5338,N_4670,N_4206);
or U5339 (N_5339,N_4124,N_4925);
nor U5340 (N_5340,N_4455,N_4387);
nand U5341 (N_5341,N_4356,N_4686);
nor U5342 (N_5342,N_4012,N_4859);
nor U5343 (N_5343,N_4464,N_4000);
and U5344 (N_5344,N_4950,N_4962);
xor U5345 (N_5345,N_4340,N_4813);
xnor U5346 (N_5346,N_4416,N_4644);
nand U5347 (N_5347,N_4045,N_4347);
or U5348 (N_5348,N_4616,N_4087);
and U5349 (N_5349,N_4303,N_4382);
nor U5350 (N_5350,N_4586,N_4191);
or U5351 (N_5351,N_4496,N_4754);
and U5352 (N_5352,N_4842,N_4877);
or U5353 (N_5353,N_4479,N_4708);
or U5354 (N_5354,N_4004,N_4335);
or U5355 (N_5355,N_4264,N_4630);
and U5356 (N_5356,N_4157,N_4996);
and U5357 (N_5357,N_4403,N_4551);
or U5358 (N_5358,N_4646,N_4283);
or U5359 (N_5359,N_4234,N_4636);
nor U5360 (N_5360,N_4949,N_4678);
or U5361 (N_5361,N_4366,N_4222);
nand U5362 (N_5362,N_4406,N_4981);
nor U5363 (N_5363,N_4658,N_4501);
nor U5364 (N_5364,N_4687,N_4975);
or U5365 (N_5365,N_4743,N_4093);
and U5366 (N_5366,N_4095,N_4198);
nand U5367 (N_5367,N_4249,N_4617);
and U5368 (N_5368,N_4851,N_4841);
nor U5369 (N_5369,N_4788,N_4766);
or U5370 (N_5370,N_4314,N_4799);
or U5371 (N_5371,N_4349,N_4294);
or U5372 (N_5372,N_4112,N_4346);
and U5373 (N_5373,N_4823,N_4651);
nor U5374 (N_5374,N_4123,N_4114);
xor U5375 (N_5375,N_4002,N_4352);
or U5376 (N_5376,N_4241,N_4676);
nand U5377 (N_5377,N_4210,N_4239);
or U5378 (N_5378,N_4672,N_4057);
or U5379 (N_5379,N_4163,N_4565);
nor U5380 (N_5380,N_4109,N_4508);
nand U5381 (N_5381,N_4230,N_4025);
nor U5382 (N_5382,N_4485,N_4942);
and U5383 (N_5383,N_4360,N_4612);
nand U5384 (N_5384,N_4561,N_4649);
or U5385 (N_5385,N_4674,N_4666);
and U5386 (N_5386,N_4923,N_4199);
nand U5387 (N_5387,N_4699,N_4745);
and U5388 (N_5388,N_4009,N_4296);
nand U5389 (N_5389,N_4117,N_4611);
and U5390 (N_5390,N_4059,N_4436);
and U5391 (N_5391,N_4534,N_4865);
and U5392 (N_5392,N_4689,N_4428);
or U5393 (N_5393,N_4074,N_4016);
nand U5394 (N_5394,N_4448,N_4838);
nand U5395 (N_5395,N_4342,N_4495);
nand U5396 (N_5396,N_4712,N_4133);
and U5397 (N_5397,N_4787,N_4939);
nor U5398 (N_5398,N_4450,N_4593);
nor U5399 (N_5399,N_4540,N_4779);
nand U5400 (N_5400,N_4797,N_4609);
or U5401 (N_5401,N_4247,N_4262);
nor U5402 (N_5402,N_4860,N_4119);
nand U5403 (N_5403,N_4852,N_4259);
or U5404 (N_5404,N_4055,N_4833);
or U5405 (N_5405,N_4044,N_4022);
and U5406 (N_5406,N_4006,N_4359);
and U5407 (N_5407,N_4334,N_4077);
nand U5408 (N_5408,N_4207,N_4758);
nand U5409 (N_5409,N_4618,N_4278);
nand U5410 (N_5410,N_4664,N_4011);
or U5411 (N_5411,N_4140,N_4125);
nand U5412 (N_5412,N_4661,N_4892);
nor U5413 (N_5413,N_4368,N_4874);
or U5414 (N_5414,N_4399,N_4545);
or U5415 (N_5415,N_4738,N_4156);
or U5416 (N_5416,N_4295,N_4527);
and U5417 (N_5417,N_4876,N_4653);
nor U5418 (N_5418,N_4762,N_4410);
or U5419 (N_5419,N_4691,N_4263);
nand U5420 (N_5420,N_4381,N_4954);
or U5421 (N_5421,N_4582,N_4315);
and U5422 (N_5422,N_4094,N_4995);
nand U5423 (N_5423,N_4915,N_4657);
and U5424 (N_5424,N_4854,N_4517);
xnor U5425 (N_5425,N_4569,N_4144);
and U5426 (N_5426,N_4465,N_4037);
or U5427 (N_5427,N_4635,N_4486);
and U5428 (N_5428,N_4153,N_4957);
nand U5429 (N_5429,N_4061,N_4218);
nor U5430 (N_5430,N_4704,N_4685);
and U5431 (N_5431,N_4638,N_4526);
nor U5432 (N_5432,N_4515,N_4955);
and U5433 (N_5433,N_4669,N_4815);
and U5434 (N_5434,N_4483,N_4591);
or U5435 (N_5435,N_4811,N_4528);
nor U5436 (N_5436,N_4752,N_4432);
and U5437 (N_5437,N_4850,N_4478);
nor U5438 (N_5438,N_4564,N_4079);
nor U5439 (N_5439,N_4603,N_4734);
nand U5440 (N_5440,N_4968,N_4795);
or U5441 (N_5441,N_4956,N_4020);
nor U5442 (N_5442,N_4948,N_4706);
nand U5443 (N_5443,N_4829,N_4292);
nand U5444 (N_5444,N_4427,N_4970);
nor U5445 (N_5445,N_4010,N_4150);
nand U5446 (N_5446,N_4848,N_4538);
and U5447 (N_5447,N_4541,N_4082);
nand U5448 (N_5448,N_4663,N_4810);
or U5449 (N_5449,N_4566,N_4393);
and U5450 (N_5450,N_4872,N_4220);
nand U5451 (N_5451,N_4433,N_4873);
or U5452 (N_5452,N_4822,N_4835);
nand U5453 (N_5453,N_4667,N_4141);
and U5454 (N_5454,N_4944,N_4196);
nor U5455 (N_5455,N_4494,N_4742);
nand U5456 (N_5456,N_4377,N_4081);
nor U5457 (N_5457,N_4928,N_4824);
nand U5458 (N_5458,N_4443,N_4964);
and U5459 (N_5459,N_4920,N_4369);
xor U5460 (N_5460,N_4720,N_4166);
nand U5461 (N_5461,N_4138,N_4243);
nor U5462 (N_5462,N_4147,N_4539);
nand U5463 (N_5463,N_4052,N_4847);
nand U5464 (N_5464,N_4162,N_4035);
or U5465 (N_5465,N_4774,N_4471);
and U5466 (N_5466,N_4073,N_4778);
or U5467 (N_5467,N_4308,N_4760);
nor U5468 (N_5468,N_4333,N_4235);
or U5469 (N_5469,N_4175,N_4458);
or U5470 (N_5470,N_4804,N_4080);
nor U5471 (N_5471,N_4831,N_4575);
nand U5472 (N_5472,N_4614,N_4577);
and U5473 (N_5473,N_4440,N_4516);
or U5474 (N_5474,N_4613,N_4933);
nand U5475 (N_5475,N_4363,N_4843);
nor U5476 (N_5476,N_4973,N_4893);
nand U5477 (N_5477,N_4595,N_4116);
and U5478 (N_5478,N_4623,N_4728);
xor U5479 (N_5479,N_4747,N_4310);
xnor U5480 (N_5480,N_4069,N_4921);
nand U5481 (N_5481,N_4417,N_4466);
or U5482 (N_5482,N_4805,N_4266);
nand U5483 (N_5483,N_4453,N_4858);
or U5484 (N_5484,N_4770,N_4233);
nand U5485 (N_5485,N_4785,N_4304);
nand U5486 (N_5486,N_4430,N_4351);
or U5487 (N_5487,N_4186,N_4469);
and U5488 (N_5488,N_4771,N_4257);
nand U5489 (N_5489,N_4456,N_4454);
nor U5490 (N_5490,N_4160,N_4106);
nor U5491 (N_5491,N_4490,N_4650);
nand U5492 (N_5492,N_4173,N_4083);
or U5493 (N_5493,N_4755,N_4001);
nand U5494 (N_5494,N_4952,N_4746);
nand U5495 (N_5495,N_4789,N_4461);
or U5496 (N_5496,N_4394,N_4879);
or U5497 (N_5497,N_4088,N_4064);
nor U5498 (N_5498,N_4648,N_4782);
and U5499 (N_5499,N_4318,N_4034);
and U5500 (N_5500,N_4492,N_4956);
nand U5501 (N_5501,N_4111,N_4358);
and U5502 (N_5502,N_4152,N_4291);
nor U5503 (N_5503,N_4903,N_4118);
nor U5504 (N_5504,N_4784,N_4776);
xor U5505 (N_5505,N_4709,N_4082);
nor U5506 (N_5506,N_4845,N_4732);
nor U5507 (N_5507,N_4653,N_4688);
and U5508 (N_5508,N_4439,N_4834);
or U5509 (N_5509,N_4362,N_4719);
and U5510 (N_5510,N_4573,N_4436);
and U5511 (N_5511,N_4715,N_4063);
nand U5512 (N_5512,N_4270,N_4005);
nand U5513 (N_5513,N_4315,N_4252);
nand U5514 (N_5514,N_4985,N_4722);
xnor U5515 (N_5515,N_4866,N_4028);
nand U5516 (N_5516,N_4848,N_4473);
or U5517 (N_5517,N_4302,N_4878);
nor U5518 (N_5518,N_4050,N_4905);
nor U5519 (N_5519,N_4036,N_4584);
or U5520 (N_5520,N_4796,N_4095);
or U5521 (N_5521,N_4540,N_4744);
or U5522 (N_5522,N_4800,N_4004);
xnor U5523 (N_5523,N_4491,N_4806);
or U5524 (N_5524,N_4794,N_4792);
or U5525 (N_5525,N_4304,N_4634);
and U5526 (N_5526,N_4340,N_4537);
nor U5527 (N_5527,N_4626,N_4780);
xor U5528 (N_5528,N_4437,N_4913);
and U5529 (N_5529,N_4150,N_4919);
nor U5530 (N_5530,N_4370,N_4399);
nor U5531 (N_5531,N_4034,N_4437);
nor U5532 (N_5532,N_4296,N_4888);
nand U5533 (N_5533,N_4440,N_4284);
and U5534 (N_5534,N_4461,N_4574);
nor U5535 (N_5535,N_4605,N_4023);
nor U5536 (N_5536,N_4430,N_4120);
and U5537 (N_5537,N_4426,N_4513);
and U5538 (N_5538,N_4597,N_4290);
or U5539 (N_5539,N_4565,N_4343);
and U5540 (N_5540,N_4192,N_4029);
nor U5541 (N_5541,N_4946,N_4101);
or U5542 (N_5542,N_4029,N_4022);
nor U5543 (N_5543,N_4572,N_4119);
nor U5544 (N_5544,N_4874,N_4605);
and U5545 (N_5545,N_4290,N_4102);
or U5546 (N_5546,N_4018,N_4928);
nand U5547 (N_5547,N_4194,N_4459);
nor U5548 (N_5548,N_4486,N_4224);
nor U5549 (N_5549,N_4261,N_4967);
and U5550 (N_5550,N_4454,N_4760);
and U5551 (N_5551,N_4982,N_4835);
nand U5552 (N_5552,N_4864,N_4179);
nor U5553 (N_5553,N_4198,N_4758);
and U5554 (N_5554,N_4027,N_4853);
nand U5555 (N_5555,N_4350,N_4937);
nor U5556 (N_5556,N_4160,N_4617);
and U5557 (N_5557,N_4587,N_4219);
or U5558 (N_5558,N_4508,N_4516);
and U5559 (N_5559,N_4546,N_4646);
nand U5560 (N_5560,N_4240,N_4659);
or U5561 (N_5561,N_4961,N_4998);
or U5562 (N_5562,N_4062,N_4263);
nand U5563 (N_5563,N_4355,N_4068);
and U5564 (N_5564,N_4280,N_4675);
nand U5565 (N_5565,N_4462,N_4926);
nor U5566 (N_5566,N_4854,N_4615);
or U5567 (N_5567,N_4350,N_4790);
or U5568 (N_5568,N_4317,N_4179);
or U5569 (N_5569,N_4729,N_4183);
and U5570 (N_5570,N_4613,N_4280);
xor U5571 (N_5571,N_4690,N_4859);
or U5572 (N_5572,N_4714,N_4865);
nor U5573 (N_5573,N_4971,N_4373);
or U5574 (N_5574,N_4928,N_4712);
nand U5575 (N_5575,N_4580,N_4487);
nand U5576 (N_5576,N_4656,N_4762);
nor U5577 (N_5577,N_4325,N_4780);
nor U5578 (N_5578,N_4067,N_4123);
or U5579 (N_5579,N_4535,N_4511);
and U5580 (N_5580,N_4299,N_4025);
nand U5581 (N_5581,N_4289,N_4061);
or U5582 (N_5582,N_4149,N_4050);
or U5583 (N_5583,N_4744,N_4026);
and U5584 (N_5584,N_4954,N_4848);
nor U5585 (N_5585,N_4361,N_4148);
nand U5586 (N_5586,N_4635,N_4791);
or U5587 (N_5587,N_4983,N_4893);
nor U5588 (N_5588,N_4333,N_4852);
nor U5589 (N_5589,N_4070,N_4643);
and U5590 (N_5590,N_4822,N_4463);
or U5591 (N_5591,N_4730,N_4764);
nand U5592 (N_5592,N_4672,N_4536);
nor U5593 (N_5593,N_4835,N_4292);
nand U5594 (N_5594,N_4469,N_4038);
nand U5595 (N_5595,N_4944,N_4702);
and U5596 (N_5596,N_4774,N_4339);
nor U5597 (N_5597,N_4520,N_4114);
nor U5598 (N_5598,N_4614,N_4948);
nand U5599 (N_5599,N_4601,N_4870);
and U5600 (N_5600,N_4456,N_4581);
and U5601 (N_5601,N_4287,N_4479);
or U5602 (N_5602,N_4720,N_4780);
and U5603 (N_5603,N_4754,N_4618);
xor U5604 (N_5604,N_4769,N_4357);
and U5605 (N_5605,N_4628,N_4204);
nor U5606 (N_5606,N_4566,N_4691);
and U5607 (N_5607,N_4464,N_4228);
or U5608 (N_5608,N_4987,N_4506);
and U5609 (N_5609,N_4384,N_4380);
nor U5610 (N_5610,N_4594,N_4713);
nand U5611 (N_5611,N_4340,N_4268);
nor U5612 (N_5612,N_4572,N_4220);
nor U5613 (N_5613,N_4471,N_4702);
and U5614 (N_5614,N_4393,N_4872);
or U5615 (N_5615,N_4338,N_4609);
nand U5616 (N_5616,N_4608,N_4633);
or U5617 (N_5617,N_4614,N_4669);
nand U5618 (N_5618,N_4638,N_4601);
nor U5619 (N_5619,N_4660,N_4454);
nand U5620 (N_5620,N_4629,N_4231);
and U5621 (N_5621,N_4029,N_4212);
nand U5622 (N_5622,N_4084,N_4089);
and U5623 (N_5623,N_4483,N_4410);
nor U5624 (N_5624,N_4063,N_4433);
and U5625 (N_5625,N_4951,N_4447);
xor U5626 (N_5626,N_4257,N_4794);
or U5627 (N_5627,N_4967,N_4192);
nand U5628 (N_5628,N_4803,N_4846);
nand U5629 (N_5629,N_4860,N_4457);
and U5630 (N_5630,N_4075,N_4800);
nor U5631 (N_5631,N_4253,N_4349);
nand U5632 (N_5632,N_4547,N_4601);
or U5633 (N_5633,N_4624,N_4808);
nand U5634 (N_5634,N_4726,N_4312);
or U5635 (N_5635,N_4904,N_4908);
or U5636 (N_5636,N_4170,N_4539);
nor U5637 (N_5637,N_4478,N_4070);
nor U5638 (N_5638,N_4696,N_4411);
nand U5639 (N_5639,N_4778,N_4182);
xnor U5640 (N_5640,N_4618,N_4076);
nor U5641 (N_5641,N_4877,N_4636);
nand U5642 (N_5642,N_4121,N_4300);
or U5643 (N_5643,N_4385,N_4148);
nor U5644 (N_5644,N_4553,N_4649);
nor U5645 (N_5645,N_4463,N_4107);
xnor U5646 (N_5646,N_4951,N_4560);
nand U5647 (N_5647,N_4136,N_4994);
or U5648 (N_5648,N_4335,N_4832);
and U5649 (N_5649,N_4163,N_4016);
nor U5650 (N_5650,N_4718,N_4678);
or U5651 (N_5651,N_4156,N_4174);
and U5652 (N_5652,N_4138,N_4568);
or U5653 (N_5653,N_4686,N_4398);
or U5654 (N_5654,N_4160,N_4537);
nor U5655 (N_5655,N_4788,N_4920);
or U5656 (N_5656,N_4067,N_4485);
or U5657 (N_5657,N_4050,N_4343);
nor U5658 (N_5658,N_4780,N_4743);
nand U5659 (N_5659,N_4893,N_4588);
nand U5660 (N_5660,N_4403,N_4570);
nand U5661 (N_5661,N_4405,N_4000);
and U5662 (N_5662,N_4834,N_4848);
or U5663 (N_5663,N_4824,N_4166);
nand U5664 (N_5664,N_4628,N_4425);
nor U5665 (N_5665,N_4304,N_4225);
nand U5666 (N_5666,N_4441,N_4976);
nor U5667 (N_5667,N_4871,N_4394);
and U5668 (N_5668,N_4361,N_4513);
nand U5669 (N_5669,N_4264,N_4052);
nor U5670 (N_5670,N_4505,N_4802);
xnor U5671 (N_5671,N_4912,N_4919);
nand U5672 (N_5672,N_4698,N_4704);
or U5673 (N_5673,N_4811,N_4416);
nand U5674 (N_5674,N_4211,N_4003);
nand U5675 (N_5675,N_4724,N_4267);
and U5676 (N_5676,N_4815,N_4184);
nor U5677 (N_5677,N_4763,N_4448);
nor U5678 (N_5678,N_4450,N_4680);
and U5679 (N_5679,N_4333,N_4783);
nand U5680 (N_5680,N_4531,N_4601);
or U5681 (N_5681,N_4316,N_4912);
nor U5682 (N_5682,N_4395,N_4978);
nand U5683 (N_5683,N_4320,N_4370);
nand U5684 (N_5684,N_4614,N_4237);
and U5685 (N_5685,N_4958,N_4480);
or U5686 (N_5686,N_4813,N_4869);
nand U5687 (N_5687,N_4569,N_4285);
or U5688 (N_5688,N_4997,N_4128);
nor U5689 (N_5689,N_4270,N_4555);
or U5690 (N_5690,N_4303,N_4162);
nor U5691 (N_5691,N_4842,N_4555);
or U5692 (N_5692,N_4757,N_4216);
nor U5693 (N_5693,N_4370,N_4650);
nor U5694 (N_5694,N_4867,N_4084);
nand U5695 (N_5695,N_4503,N_4973);
nor U5696 (N_5696,N_4299,N_4312);
nand U5697 (N_5697,N_4712,N_4878);
and U5698 (N_5698,N_4138,N_4678);
nor U5699 (N_5699,N_4560,N_4424);
nand U5700 (N_5700,N_4588,N_4205);
nand U5701 (N_5701,N_4605,N_4084);
nor U5702 (N_5702,N_4436,N_4745);
nand U5703 (N_5703,N_4045,N_4168);
nand U5704 (N_5704,N_4698,N_4859);
or U5705 (N_5705,N_4557,N_4653);
or U5706 (N_5706,N_4051,N_4408);
and U5707 (N_5707,N_4081,N_4638);
nor U5708 (N_5708,N_4032,N_4955);
nand U5709 (N_5709,N_4880,N_4395);
nor U5710 (N_5710,N_4482,N_4108);
and U5711 (N_5711,N_4511,N_4172);
and U5712 (N_5712,N_4085,N_4980);
nand U5713 (N_5713,N_4757,N_4548);
and U5714 (N_5714,N_4925,N_4220);
or U5715 (N_5715,N_4763,N_4142);
or U5716 (N_5716,N_4911,N_4126);
nor U5717 (N_5717,N_4509,N_4630);
nor U5718 (N_5718,N_4298,N_4624);
or U5719 (N_5719,N_4230,N_4871);
and U5720 (N_5720,N_4358,N_4120);
nor U5721 (N_5721,N_4283,N_4917);
and U5722 (N_5722,N_4316,N_4343);
or U5723 (N_5723,N_4783,N_4174);
and U5724 (N_5724,N_4044,N_4646);
xnor U5725 (N_5725,N_4941,N_4678);
or U5726 (N_5726,N_4520,N_4585);
or U5727 (N_5727,N_4945,N_4020);
and U5728 (N_5728,N_4426,N_4907);
nor U5729 (N_5729,N_4047,N_4860);
nor U5730 (N_5730,N_4893,N_4431);
or U5731 (N_5731,N_4636,N_4946);
and U5732 (N_5732,N_4660,N_4091);
or U5733 (N_5733,N_4702,N_4443);
or U5734 (N_5734,N_4945,N_4327);
nand U5735 (N_5735,N_4364,N_4386);
nor U5736 (N_5736,N_4186,N_4192);
and U5737 (N_5737,N_4014,N_4732);
xor U5738 (N_5738,N_4007,N_4698);
nand U5739 (N_5739,N_4796,N_4160);
nor U5740 (N_5740,N_4210,N_4686);
or U5741 (N_5741,N_4817,N_4058);
nor U5742 (N_5742,N_4169,N_4578);
or U5743 (N_5743,N_4691,N_4756);
and U5744 (N_5744,N_4635,N_4394);
nand U5745 (N_5745,N_4154,N_4619);
nand U5746 (N_5746,N_4766,N_4139);
nor U5747 (N_5747,N_4983,N_4531);
and U5748 (N_5748,N_4557,N_4102);
or U5749 (N_5749,N_4141,N_4351);
or U5750 (N_5750,N_4803,N_4326);
xor U5751 (N_5751,N_4899,N_4613);
and U5752 (N_5752,N_4582,N_4260);
nand U5753 (N_5753,N_4948,N_4881);
nor U5754 (N_5754,N_4272,N_4711);
nor U5755 (N_5755,N_4556,N_4477);
nor U5756 (N_5756,N_4291,N_4251);
or U5757 (N_5757,N_4251,N_4944);
nor U5758 (N_5758,N_4760,N_4260);
and U5759 (N_5759,N_4732,N_4922);
nand U5760 (N_5760,N_4952,N_4628);
nor U5761 (N_5761,N_4139,N_4839);
or U5762 (N_5762,N_4394,N_4281);
or U5763 (N_5763,N_4894,N_4549);
or U5764 (N_5764,N_4732,N_4837);
nor U5765 (N_5765,N_4813,N_4310);
or U5766 (N_5766,N_4596,N_4510);
and U5767 (N_5767,N_4888,N_4534);
nor U5768 (N_5768,N_4006,N_4573);
nor U5769 (N_5769,N_4319,N_4001);
and U5770 (N_5770,N_4366,N_4135);
and U5771 (N_5771,N_4229,N_4550);
nand U5772 (N_5772,N_4385,N_4945);
and U5773 (N_5773,N_4612,N_4338);
nand U5774 (N_5774,N_4779,N_4006);
or U5775 (N_5775,N_4535,N_4619);
and U5776 (N_5776,N_4051,N_4996);
and U5777 (N_5777,N_4948,N_4784);
nand U5778 (N_5778,N_4016,N_4246);
or U5779 (N_5779,N_4095,N_4851);
nor U5780 (N_5780,N_4033,N_4601);
or U5781 (N_5781,N_4949,N_4743);
nand U5782 (N_5782,N_4959,N_4543);
or U5783 (N_5783,N_4795,N_4007);
and U5784 (N_5784,N_4589,N_4518);
nand U5785 (N_5785,N_4738,N_4296);
nand U5786 (N_5786,N_4244,N_4560);
and U5787 (N_5787,N_4478,N_4060);
and U5788 (N_5788,N_4497,N_4972);
and U5789 (N_5789,N_4742,N_4409);
nor U5790 (N_5790,N_4336,N_4034);
or U5791 (N_5791,N_4659,N_4979);
nand U5792 (N_5792,N_4452,N_4338);
and U5793 (N_5793,N_4089,N_4092);
nor U5794 (N_5794,N_4177,N_4554);
nor U5795 (N_5795,N_4379,N_4998);
or U5796 (N_5796,N_4707,N_4294);
or U5797 (N_5797,N_4886,N_4089);
nor U5798 (N_5798,N_4288,N_4879);
or U5799 (N_5799,N_4250,N_4830);
xor U5800 (N_5800,N_4078,N_4930);
nand U5801 (N_5801,N_4960,N_4666);
nor U5802 (N_5802,N_4070,N_4147);
nand U5803 (N_5803,N_4799,N_4244);
and U5804 (N_5804,N_4675,N_4143);
nand U5805 (N_5805,N_4472,N_4283);
and U5806 (N_5806,N_4291,N_4588);
nand U5807 (N_5807,N_4918,N_4060);
or U5808 (N_5808,N_4980,N_4519);
and U5809 (N_5809,N_4324,N_4881);
nand U5810 (N_5810,N_4395,N_4859);
nor U5811 (N_5811,N_4465,N_4820);
nor U5812 (N_5812,N_4634,N_4715);
or U5813 (N_5813,N_4329,N_4593);
or U5814 (N_5814,N_4966,N_4761);
or U5815 (N_5815,N_4798,N_4745);
and U5816 (N_5816,N_4360,N_4860);
and U5817 (N_5817,N_4518,N_4657);
or U5818 (N_5818,N_4951,N_4643);
nor U5819 (N_5819,N_4178,N_4374);
or U5820 (N_5820,N_4956,N_4075);
and U5821 (N_5821,N_4632,N_4549);
or U5822 (N_5822,N_4687,N_4245);
xnor U5823 (N_5823,N_4695,N_4705);
xnor U5824 (N_5824,N_4542,N_4017);
nand U5825 (N_5825,N_4326,N_4331);
nand U5826 (N_5826,N_4391,N_4513);
nand U5827 (N_5827,N_4250,N_4526);
and U5828 (N_5828,N_4508,N_4351);
nand U5829 (N_5829,N_4539,N_4380);
nand U5830 (N_5830,N_4967,N_4352);
xnor U5831 (N_5831,N_4520,N_4380);
nor U5832 (N_5832,N_4696,N_4966);
nor U5833 (N_5833,N_4269,N_4292);
and U5834 (N_5834,N_4113,N_4179);
or U5835 (N_5835,N_4067,N_4419);
nand U5836 (N_5836,N_4659,N_4367);
or U5837 (N_5837,N_4067,N_4898);
and U5838 (N_5838,N_4118,N_4781);
nor U5839 (N_5839,N_4287,N_4807);
nand U5840 (N_5840,N_4483,N_4317);
nand U5841 (N_5841,N_4012,N_4272);
or U5842 (N_5842,N_4457,N_4915);
and U5843 (N_5843,N_4740,N_4894);
nor U5844 (N_5844,N_4583,N_4907);
and U5845 (N_5845,N_4363,N_4857);
and U5846 (N_5846,N_4373,N_4360);
and U5847 (N_5847,N_4705,N_4366);
and U5848 (N_5848,N_4971,N_4965);
or U5849 (N_5849,N_4896,N_4053);
nand U5850 (N_5850,N_4890,N_4627);
or U5851 (N_5851,N_4961,N_4050);
and U5852 (N_5852,N_4345,N_4993);
and U5853 (N_5853,N_4299,N_4376);
nor U5854 (N_5854,N_4763,N_4929);
nor U5855 (N_5855,N_4028,N_4962);
or U5856 (N_5856,N_4684,N_4963);
and U5857 (N_5857,N_4764,N_4956);
or U5858 (N_5858,N_4372,N_4464);
nor U5859 (N_5859,N_4324,N_4889);
xnor U5860 (N_5860,N_4891,N_4938);
and U5861 (N_5861,N_4539,N_4258);
or U5862 (N_5862,N_4463,N_4482);
xor U5863 (N_5863,N_4441,N_4967);
nor U5864 (N_5864,N_4068,N_4036);
nor U5865 (N_5865,N_4926,N_4099);
and U5866 (N_5866,N_4094,N_4924);
nor U5867 (N_5867,N_4980,N_4849);
nand U5868 (N_5868,N_4156,N_4325);
xnor U5869 (N_5869,N_4041,N_4189);
and U5870 (N_5870,N_4883,N_4401);
or U5871 (N_5871,N_4300,N_4243);
nor U5872 (N_5872,N_4044,N_4318);
or U5873 (N_5873,N_4645,N_4710);
and U5874 (N_5874,N_4094,N_4807);
or U5875 (N_5875,N_4902,N_4451);
nor U5876 (N_5876,N_4052,N_4595);
nor U5877 (N_5877,N_4704,N_4062);
nor U5878 (N_5878,N_4445,N_4903);
and U5879 (N_5879,N_4563,N_4489);
nor U5880 (N_5880,N_4047,N_4537);
nor U5881 (N_5881,N_4750,N_4262);
or U5882 (N_5882,N_4542,N_4553);
nand U5883 (N_5883,N_4927,N_4991);
nor U5884 (N_5884,N_4397,N_4235);
or U5885 (N_5885,N_4356,N_4391);
or U5886 (N_5886,N_4765,N_4148);
nor U5887 (N_5887,N_4921,N_4623);
and U5888 (N_5888,N_4205,N_4610);
nand U5889 (N_5889,N_4896,N_4497);
nor U5890 (N_5890,N_4701,N_4714);
and U5891 (N_5891,N_4689,N_4840);
nand U5892 (N_5892,N_4043,N_4445);
and U5893 (N_5893,N_4575,N_4003);
or U5894 (N_5894,N_4587,N_4033);
nand U5895 (N_5895,N_4060,N_4538);
nand U5896 (N_5896,N_4280,N_4136);
or U5897 (N_5897,N_4321,N_4024);
or U5898 (N_5898,N_4934,N_4511);
and U5899 (N_5899,N_4094,N_4551);
nor U5900 (N_5900,N_4069,N_4075);
or U5901 (N_5901,N_4227,N_4612);
nand U5902 (N_5902,N_4580,N_4151);
and U5903 (N_5903,N_4229,N_4855);
or U5904 (N_5904,N_4923,N_4338);
nand U5905 (N_5905,N_4230,N_4081);
nand U5906 (N_5906,N_4243,N_4681);
or U5907 (N_5907,N_4521,N_4752);
nand U5908 (N_5908,N_4356,N_4558);
or U5909 (N_5909,N_4190,N_4742);
nand U5910 (N_5910,N_4630,N_4113);
or U5911 (N_5911,N_4325,N_4388);
and U5912 (N_5912,N_4117,N_4783);
and U5913 (N_5913,N_4543,N_4277);
nor U5914 (N_5914,N_4365,N_4212);
and U5915 (N_5915,N_4062,N_4281);
nand U5916 (N_5916,N_4089,N_4598);
or U5917 (N_5917,N_4124,N_4730);
nand U5918 (N_5918,N_4305,N_4617);
and U5919 (N_5919,N_4156,N_4839);
nor U5920 (N_5920,N_4755,N_4686);
or U5921 (N_5921,N_4992,N_4353);
nand U5922 (N_5922,N_4295,N_4693);
nand U5923 (N_5923,N_4107,N_4093);
nand U5924 (N_5924,N_4470,N_4307);
nand U5925 (N_5925,N_4903,N_4917);
and U5926 (N_5926,N_4529,N_4110);
nor U5927 (N_5927,N_4674,N_4550);
nor U5928 (N_5928,N_4445,N_4414);
nor U5929 (N_5929,N_4670,N_4013);
and U5930 (N_5930,N_4095,N_4018);
or U5931 (N_5931,N_4938,N_4042);
nand U5932 (N_5932,N_4702,N_4194);
and U5933 (N_5933,N_4889,N_4595);
nand U5934 (N_5934,N_4075,N_4945);
nor U5935 (N_5935,N_4330,N_4486);
nor U5936 (N_5936,N_4399,N_4146);
nand U5937 (N_5937,N_4793,N_4225);
nand U5938 (N_5938,N_4786,N_4361);
nor U5939 (N_5939,N_4500,N_4675);
nand U5940 (N_5940,N_4736,N_4996);
nand U5941 (N_5941,N_4356,N_4370);
nand U5942 (N_5942,N_4712,N_4033);
nand U5943 (N_5943,N_4577,N_4112);
and U5944 (N_5944,N_4012,N_4173);
and U5945 (N_5945,N_4821,N_4793);
or U5946 (N_5946,N_4348,N_4480);
nand U5947 (N_5947,N_4216,N_4163);
or U5948 (N_5948,N_4851,N_4709);
nor U5949 (N_5949,N_4488,N_4659);
nor U5950 (N_5950,N_4048,N_4538);
nand U5951 (N_5951,N_4835,N_4750);
nor U5952 (N_5952,N_4532,N_4732);
or U5953 (N_5953,N_4064,N_4727);
nor U5954 (N_5954,N_4370,N_4698);
or U5955 (N_5955,N_4432,N_4783);
nor U5956 (N_5956,N_4248,N_4780);
nor U5957 (N_5957,N_4561,N_4248);
nor U5958 (N_5958,N_4043,N_4787);
and U5959 (N_5959,N_4037,N_4804);
and U5960 (N_5960,N_4011,N_4939);
and U5961 (N_5961,N_4060,N_4472);
nor U5962 (N_5962,N_4953,N_4245);
nor U5963 (N_5963,N_4790,N_4426);
and U5964 (N_5964,N_4105,N_4141);
nor U5965 (N_5965,N_4558,N_4209);
nor U5966 (N_5966,N_4619,N_4504);
and U5967 (N_5967,N_4802,N_4893);
nand U5968 (N_5968,N_4660,N_4170);
nor U5969 (N_5969,N_4088,N_4705);
nand U5970 (N_5970,N_4777,N_4791);
and U5971 (N_5971,N_4558,N_4461);
nor U5972 (N_5972,N_4765,N_4401);
nor U5973 (N_5973,N_4989,N_4273);
nor U5974 (N_5974,N_4115,N_4059);
nor U5975 (N_5975,N_4035,N_4116);
or U5976 (N_5976,N_4431,N_4347);
nand U5977 (N_5977,N_4671,N_4391);
nand U5978 (N_5978,N_4236,N_4703);
nor U5979 (N_5979,N_4780,N_4981);
and U5980 (N_5980,N_4078,N_4151);
nand U5981 (N_5981,N_4651,N_4166);
and U5982 (N_5982,N_4220,N_4569);
or U5983 (N_5983,N_4765,N_4843);
and U5984 (N_5984,N_4243,N_4494);
nand U5985 (N_5985,N_4046,N_4108);
and U5986 (N_5986,N_4567,N_4292);
or U5987 (N_5987,N_4329,N_4939);
nand U5988 (N_5988,N_4452,N_4089);
nor U5989 (N_5989,N_4451,N_4755);
xor U5990 (N_5990,N_4309,N_4487);
and U5991 (N_5991,N_4276,N_4343);
nor U5992 (N_5992,N_4752,N_4456);
nand U5993 (N_5993,N_4388,N_4683);
and U5994 (N_5994,N_4290,N_4837);
nor U5995 (N_5995,N_4768,N_4563);
or U5996 (N_5996,N_4560,N_4641);
nand U5997 (N_5997,N_4139,N_4875);
nand U5998 (N_5998,N_4645,N_4944);
xor U5999 (N_5999,N_4366,N_4937);
or U6000 (N_6000,N_5585,N_5659);
nand U6001 (N_6001,N_5580,N_5940);
or U6002 (N_6002,N_5710,N_5217);
and U6003 (N_6003,N_5104,N_5187);
xor U6004 (N_6004,N_5903,N_5501);
xnor U6005 (N_6005,N_5427,N_5166);
nor U6006 (N_6006,N_5488,N_5632);
nand U6007 (N_6007,N_5938,N_5729);
nor U6008 (N_6008,N_5790,N_5958);
or U6009 (N_6009,N_5907,N_5440);
or U6010 (N_6010,N_5119,N_5718);
and U6011 (N_6011,N_5540,N_5816);
or U6012 (N_6012,N_5994,N_5365);
nor U6013 (N_6013,N_5570,N_5114);
nor U6014 (N_6014,N_5830,N_5693);
and U6015 (N_6015,N_5058,N_5189);
and U6016 (N_6016,N_5424,N_5688);
nand U6017 (N_6017,N_5452,N_5256);
nand U6018 (N_6018,N_5476,N_5571);
nor U6019 (N_6019,N_5920,N_5285);
and U6020 (N_6020,N_5018,N_5557);
nor U6021 (N_6021,N_5368,N_5526);
nor U6022 (N_6022,N_5982,N_5354);
nor U6023 (N_6023,N_5727,N_5981);
nand U6024 (N_6024,N_5579,N_5504);
or U6025 (N_6025,N_5653,N_5845);
nor U6026 (N_6026,N_5881,N_5431);
and U6027 (N_6027,N_5265,N_5900);
nand U6028 (N_6028,N_5877,N_5208);
nand U6029 (N_6029,N_5963,N_5181);
or U6030 (N_6030,N_5482,N_5893);
and U6031 (N_6031,N_5038,N_5964);
and U6032 (N_6032,N_5142,N_5651);
or U6033 (N_6033,N_5264,N_5303);
and U6034 (N_6034,N_5233,N_5660);
and U6035 (N_6035,N_5478,N_5875);
and U6036 (N_6036,N_5808,N_5274);
and U6037 (N_6037,N_5528,N_5458);
nor U6038 (N_6038,N_5453,N_5983);
and U6039 (N_6039,N_5369,N_5402);
and U6040 (N_6040,N_5507,N_5882);
or U6041 (N_6041,N_5673,N_5449);
nor U6042 (N_6042,N_5690,N_5908);
nor U6043 (N_6043,N_5569,N_5413);
and U6044 (N_6044,N_5681,N_5305);
nor U6045 (N_6045,N_5692,N_5203);
or U6046 (N_6046,N_5812,N_5025);
or U6047 (N_6047,N_5950,N_5205);
nand U6048 (N_6048,N_5778,N_5193);
nor U6049 (N_6049,N_5694,N_5498);
nor U6050 (N_6050,N_5664,N_5514);
nand U6051 (N_6051,N_5253,N_5210);
or U6052 (N_6052,N_5002,N_5192);
or U6053 (N_6053,N_5496,N_5966);
nor U6054 (N_6054,N_5141,N_5717);
and U6055 (N_6055,N_5311,N_5574);
and U6056 (N_6056,N_5480,N_5202);
nor U6057 (N_6057,N_5495,N_5149);
and U6058 (N_6058,N_5095,N_5280);
or U6059 (N_6059,N_5392,N_5765);
nand U6060 (N_6060,N_5968,N_5323);
nor U6061 (N_6061,N_5014,N_5521);
nor U6062 (N_6062,N_5857,N_5872);
and U6063 (N_6063,N_5417,N_5602);
nor U6064 (N_6064,N_5869,N_5609);
and U6065 (N_6065,N_5039,N_5566);
xor U6066 (N_6066,N_5426,N_5530);
or U6067 (N_6067,N_5022,N_5735);
nand U6068 (N_6068,N_5590,N_5071);
nand U6069 (N_6069,N_5858,N_5337);
and U6070 (N_6070,N_5593,N_5827);
nor U6071 (N_6071,N_5883,N_5581);
or U6072 (N_6072,N_5661,N_5257);
nand U6073 (N_6073,N_5955,N_5545);
or U6074 (N_6074,N_5578,N_5915);
and U6075 (N_6075,N_5315,N_5596);
and U6076 (N_6076,N_5251,N_5298);
and U6077 (N_6077,N_5377,N_5836);
and U6078 (N_6078,N_5299,N_5644);
or U6079 (N_6079,N_5465,N_5942);
nor U6080 (N_6080,N_5922,N_5435);
nor U6081 (N_6081,N_5512,N_5373);
nand U6082 (N_6082,N_5446,N_5469);
nor U6083 (N_6083,N_5577,N_5375);
nor U6084 (N_6084,N_5143,N_5973);
nand U6085 (N_6085,N_5050,N_5949);
nand U6086 (N_6086,N_5161,N_5916);
nor U6087 (N_6087,N_5394,N_5185);
or U6088 (N_6088,N_5783,N_5627);
nor U6089 (N_6089,N_5535,N_5636);
and U6090 (N_6090,N_5500,N_5333);
xnor U6091 (N_6091,N_5975,N_5352);
nand U6092 (N_6092,N_5689,N_5183);
or U6093 (N_6093,N_5764,N_5445);
or U6094 (N_6094,N_5906,N_5065);
and U6095 (N_6095,N_5246,N_5312);
nor U6096 (N_6096,N_5471,N_5291);
and U6097 (N_6097,N_5033,N_5235);
and U6098 (N_6098,N_5163,N_5697);
or U6099 (N_6099,N_5854,N_5505);
and U6100 (N_6100,N_5616,N_5948);
nand U6101 (N_6101,N_5999,N_5112);
nor U6102 (N_6102,N_5592,N_5603);
nor U6103 (N_6103,N_5666,N_5206);
or U6104 (N_6104,N_5489,N_5629);
and U6105 (N_6105,N_5158,N_5788);
and U6106 (N_6106,N_5013,N_5294);
or U6107 (N_6107,N_5364,N_5840);
and U6108 (N_6108,N_5306,N_5277);
nor U6109 (N_6109,N_5642,N_5699);
or U6110 (N_6110,N_5726,N_5792);
or U6111 (N_6111,N_5110,N_5209);
nand U6112 (N_6112,N_5643,N_5069);
and U6113 (N_6113,N_5288,N_5194);
nand U6114 (N_6114,N_5125,N_5524);
and U6115 (N_6115,N_5782,N_5750);
nor U6116 (N_6116,N_5229,N_5184);
nand U6117 (N_6117,N_5484,N_5584);
nand U6118 (N_6118,N_5096,N_5587);
or U6119 (N_6119,N_5000,N_5770);
or U6120 (N_6120,N_5946,N_5292);
nor U6121 (N_6121,N_5687,N_5224);
and U6122 (N_6122,N_5696,N_5672);
or U6123 (N_6123,N_5595,N_5116);
and U6124 (N_6124,N_5541,N_5680);
nor U6125 (N_6125,N_5047,N_5046);
or U6126 (N_6126,N_5434,N_5554);
nor U6127 (N_6127,N_5519,N_5391);
nand U6128 (N_6128,N_5227,N_5492);
or U6129 (N_6129,N_5138,N_5561);
nand U6130 (N_6130,N_5057,N_5043);
and U6131 (N_6131,N_5275,N_5068);
nand U6132 (N_6132,N_5721,N_5175);
or U6133 (N_6133,N_5834,N_5040);
and U6134 (N_6134,N_5191,N_5021);
or U6135 (N_6135,N_5977,N_5508);
or U6136 (N_6136,N_5272,N_5268);
nand U6137 (N_6137,N_5219,N_5657);
nor U6138 (N_6138,N_5873,N_5329);
and U6139 (N_6139,N_5620,N_5885);
and U6140 (N_6140,N_5326,N_5487);
or U6141 (N_6141,N_5506,N_5685);
nand U6142 (N_6142,N_5943,N_5742);
nor U6143 (N_6143,N_5670,N_5316);
nand U6144 (N_6144,N_5317,N_5167);
nand U6145 (N_6145,N_5608,N_5220);
and U6146 (N_6146,N_5925,N_5150);
or U6147 (N_6147,N_5748,N_5513);
and U6148 (N_6148,N_5041,N_5995);
nor U6149 (N_6149,N_5042,N_5543);
nand U6150 (N_6150,N_5361,N_5271);
or U6151 (N_6151,N_5803,N_5542);
or U6152 (N_6152,N_5518,N_5850);
or U6153 (N_6153,N_5769,N_5852);
nor U6154 (N_6154,N_5991,N_5090);
or U6155 (N_6155,N_5768,N_5357);
nand U6156 (N_6156,N_5197,N_5060);
and U6157 (N_6157,N_5867,N_5130);
nor U6158 (N_6158,N_5663,N_5447);
or U6159 (N_6159,N_5386,N_5266);
or U6160 (N_6160,N_5855,N_5888);
or U6161 (N_6161,N_5332,N_5558);
or U6162 (N_6162,N_5555,N_5878);
nor U6163 (N_6163,N_5250,N_5811);
and U6164 (N_6164,N_5509,N_5847);
nand U6165 (N_6165,N_5752,N_5556);
nand U6166 (N_6166,N_5610,N_5404);
or U6167 (N_6167,N_5347,N_5957);
nand U6168 (N_6168,N_5012,N_5269);
nand U6169 (N_6169,N_5630,N_5705);
or U6170 (N_6170,N_5416,N_5846);
nor U6171 (N_6171,N_5213,N_5247);
nand U6172 (N_6172,N_5457,N_5635);
and U6173 (N_6173,N_5407,N_5573);
or U6174 (N_6174,N_5722,N_5563);
nor U6175 (N_6175,N_5342,N_5686);
or U6176 (N_6176,N_5639,N_5338);
or U6177 (N_6177,N_5460,N_5700);
nand U6178 (N_6178,N_5385,N_5007);
nand U6179 (N_6179,N_5100,N_5249);
and U6180 (N_6180,N_5199,N_5665);
nand U6181 (N_6181,N_5165,N_5132);
nor U6182 (N_6182,N_5243,N_5522);
or U6183 (N_6183,N_5862,N_5910);
and U6184 (N_6184,N_5698,N_5860);
nor U6185 (N_6185,N_5024,N_5422);
nor U6186 (N_6186,N_5497,N_5008);
nand U6187 (N_6187,N_5137,N_5919);
nor U6188 (N_6188,N_5456,N_5151);
nand U6189 (N_6189,N_5234,N_5108);
and U6190 (N_6190,N_5675,N_5641);
nand U6191 (N_6191,N_5281,N_5472);
nor U6192 (N_6192,N_5241,N_5182);
nand U6193 (N_6193,N_5201,N_5147);
and U6194 (N_6194,N_5087,N_5853);
nor U6195 (N_6195,N_5083,N_5470);
nand U6196 (N_6196,N_5838,N_5795);
and U6197 (N_6197,N_5668,N_5564);
and U6198 (N_6198,N_5738,N_5913);
or U6199 (N_6199,N_5619,N_5604);
and U6200 (N_6200,N_5929,N_5839);
nand U6201 (N_6201,N_5437,N_5451);
and U6202 (N_6202,N_5905,N_5985);
nand U6203 (N_6203,N_5390,N_5844);
nor U6204 (N_6204,N_5055,N_5341);
nor U6205 (N_6205,N_5749,N_5646);
xor U6206 (N_6206,N_5328,N_5180);
nand U6207 (N_6207,N_5831,N_5576);
or U6208 (N_6208,N_5794,N_5898);
nand U6209 (N_6209,N_5010,N_5403);
and U6210 (N_6210,N_5529,N_5466);
nand U6211 (N_6211,N_5947,N_5760);
nor U6212 (N_6212,N_5345,N_5767);
nor U6213 (N_6213,N_5992,N_5015);
nand U6214 (N_6214,N_5463,N_5829);
and U6215 (N_6215,N_5918,N_5911);
and U6216 (N_6216,N_5682,N_5841);
or U6217 (N_6217,N_5837,N_5117);
and U6218 (N_6218,N_5037,N_5493);
and U6219 (N_6219,N_5876,N_5168);
or U6220 (N_6220,N_5155,N_5886);
or U6221 (N_6221,N_5684,N_5173);
or U6222 (N_6222,N_5270,N_5066);
nor U6223 (N_6223,N_5936,N_5436);
and U6224 (N_6224,N_5605,N_5360);
and U6225 (N_6225,N_5023,N_5061);
nor U6226 (N_6226,N_5399,N_5070);
nor U6227 (N_6227,N_5945,N_5239);
nand U6228 (N_6228,N_5828,N_5704);
nand U6229 (N_6229,N_5230,N_5473);
nand U6230 (N_6230,N_5093,N_5804);
nor U6231 (N_6231,N_5927,N_5640);
and U6232 (N_6232,N_5589,N_5546);
nor U6233 (N_6233,N_5186,N_5412);
and U6234 (N_6234,N_5433,N_5088);
and U6235 (N_6235,N_5279,N_5379);
nand U6236 (N_6236,N_5931,N_5309);
nor U6237 (N_6237,N_5154,N_5724);
nand U6238 (N_6238,N_5725,N_5099);
xor U6239 (N_6239,N_5313,N_5094);
and U6240 (N_6240,N_5153,N_5990);
nor U6241 (N_6241,N_5773,N_5459);
or U6242 (N_6242,N_5741,N_5565);
or U6243 (N_6243,N_5959,N_5650);
or U6244 (N_6244,N_5516,N_5005);
and U6245 (N_6245,N_5889,N_5824);
and U6246 (N_6246,N_5172,N_5145);
nor U6247 (N_6247,N_5904,N_5708);
nand U6248 (N_6248,N_5932,N_5358);
xor U6249 (N_6249,N_5989,N_5009);
nor U6250 (N_6250,N_5089,N_5113);
and U6251 (N_6251,N_5396,N_5638);
nand U6252 (N_6252,N_5737,N_5380);
nor U6253 (N_6253,N_5398,N_5606);
nor U6254 (N_6254,N_5429,N_5510);
or U6255 (N_6255,N_5215,N_5988);
and U6256 (N_6256,N_5971,N_5625);
and U6257 (N_6257,N_5884,N_5863);
or U6258 (N_6258,N_5411,N_5754);
and U6259 (N_6259,N_5074,N_5715);
nand U6260 (N_6260,N_5683,N_5819);
nor U6261 (N_6261,N_5679,N_5621);
nand U6262 (N_6262,N_5133,N_5842);
nand U6263 (N_6263,N_5986,N_5410);
and U6264 (N_6264,N_5937,N_5597);
xor U6265 (N_6265,N_5822,N_5740);
nand U6266 (N_6266,N_5418,N_5136);
and U6267 (N_6267,N_5295,N_5691);
nand U6268 (N_6268,N_5996,N_5951);
nand U6269 (N_6269,N_5965,N_5178);
and U6270 (N_6270,N_5674,N_5924);
nor U6271 (N_6271,N_5871,N_5314);
or U6272 (N_6272,N_5382,N_5772);
or U6273 (N_6273,N_5258,N_5102);
or U6274 (N_6274,N_5118,N_5400);
or U6275 (N_6275,N_5899,N_5601);
xor U6276 (N_6276,N_5960,N_5775);
nand U6277 (N_6277,N_5408,N_5798);
or U6278 (N_6278,N_5976,N_5286);
nand U6279 (N_6279,N_5053,N_5739);
or U6280 (N_6280,N_5421,N_5438);
nand U6281 (N_6281,N_5188,N_5962);
and U6282 (N_6282,N_5054,N_5912);
and U6283 (N_6283,N_5503,N_5848);
nor U6284 (N_6284,N_5260,N_5146);
or U6285 (N_6285,N_5720,N_5887);
nor U6286 (N_6286,N_5802,N_5226);
and U6287 (N_6287,N_5044,N_5395);
nand U6288 (N_6288,N_5917,N_5953);
and U6289 (N_6289,N_5654,N_5441);
and U6290 (N_6290,N_5159,N_5036);
xor U6291 (N_6291,N_5124,N_5761);
or U6292 (N_6292,N_5961,N_5901);
and U6293 (N_6293,N_5835,N_5228);
nor U6294 (N_6294,N_5276,N_5216);
and U6295 (N_6295,N_5020,N_5970);
nor U6296 (N_6296,N_5304,N_5211);
nor U6297 (N_6297,N_5063,N_5111);
nor U6298 (N_6298,N_5709,N_5198);
nor U6299 (N_6299,N_5598,N_5520);
nor U6300 (N_6300,N_5784,N_5359);
nor U6301 (N_6301,N_5204,N_5669);
nor U6302 (N_6302,N_5252,N_5930);
nand U6303 (N_6303,N_5527,N_5032);
and U6304 (N_6304,N_5353,N_5174);
nand U6305 (N_6305,N_5567,N_5572);
nor U6306 (N_6306,N_5156,N_5736);
xor U6307 (N_6307,N_5339,N_5894);
and U6308 (N_6308,N_5370,N_5979);
nor U6309 (N_6309,N_5348,N_5397);
and U6310 (N_6310,N_5231,N_5085);
and U6311 (N_6311,N_5468,N_5956);
nor U6312 (N_6312,N_5310,N_5122);
nand U6313 (N_6313,N_5092,N_5006);
or U6314 (N_6314,N_5637,N_5030);
and U6315 (N_6315,N_5611,N_5287);
xor U6316 (N_6316,N_5677,N_5515);
and U6317 (N_6317,N_5594,N_5049);
or U6318 (N_6318,N_5072,N_5475);
and U6319 (N_6319,N_5479,N_5805);
and U6320 (N_6320,N_5890,N_5731);
nand U6321 (N_6321,N_5103,N_5486);
nand U6322 (N_6322,N_5952,N_5714);
and U6323 (N_6323,N_5381,N_5483);
and U6324 (N_6324,N_5052,N_5222);
nand U6325 (N_6325,N_5255,N_5363);
or U6326 (N_6326,N_5248,N_5330);
nand U6327 (N_6327,N_5533,N_5549);
and U6328 (N_6328,N_5236,N_5001);
nor U6329 (N_6329,N_5467,N_5097);
xnor U6330 (N_6330,N_5485,N_5716);
and U6331 (N_6331,N_5575,N_5356);
or U6332 (N_6332,N_5212,N_5162);
nor U6333 (N_6333,N_5176,N_5179);
nor U6334 (N_6334,N_5393,N_5107);
xor U6335 (N_6335,N_5517,N_5327);
or U6336 (N_6336,N_5810,N_5780);
nand U6337 (N_6337,N_5712,N_5879);
nand U6338 (N_6338,N_5695,N_5164);
nor U6339 (N_6339,N_5336,N_5101);
and U6340 (N_6340,N_5613,N_5634);
nand U6341 (N_6341,N_5225,N_5238);
nor U6342 (N_6342,N_5531,N_5652);
nand U6343 (N_6343,N_5614,N_5711);
nor U6344 (N_6344,N_5762,N_5091);
nor U6345 (N_6345,N_5997,N_5617);
nor U6346 (N_6346,N_5800,N_5797);
nor U6347 (N_6347,N_5171,N_5388);
nor U6348 (N_6348,N_5321,N_5713);
and U6349 (N_6349,N_5031,N_5322);
or U6350 (N_6350,N_5851,N_5525);
nor U6351 (N_6351,N_5387,N_5600);
nor U6352 (N_6352,N_5254,N_5921);
or U6353 (N_6353,N_5335,N_5443);
and U6354 (N_6354,N_5523,N_5734);
nor U6355 (N_6355,N_5261,N_5823);
xnor U6356 (N_6356,N_5073,N_5745);
nand U6357 (N_6357,N_5035,N_5537);
or U6358 (N_6358,N_5926,N_5384);
xnor U6359 (N_6359,N_5892,N_5051);
or U6360 (N_6360,N_5914,N_5121);
or U6361 (N_6361,N_5993,N_5730);
nor U6362 (N_6362,N_5732,N_5334);
and U6363 (N_6363,N_5372,N_5552);
and U6364 (N_6364,N_5389,N_5454);
and U6365 (N_6365,N_5719,N_5371);
and U6366 (N_6366,N_5902,N_5987);
and U6367 (N_6367,N_5706,N_5405);
nand U6368 (N_6368,N_5733,N_5702);
nor U6369 (N_6369,N_5755,N_5771);
nand U6370 (N_6370,N_5293,N_5980);
nand U6371 (N_6371,N_5544,N_5870);
nand U6372 (N_6372,N_5079,N_5757);
or U6373 (N_6373,N_5756,N_5029);
and U6374 (N_6374,N_5809,N_5591);
nand U6375 (N_6375,N_5599,N_5307);
or U6376 (N_6376,N_5200,N_5701);
nand U6377 (N_6377,N_5290,N_5267);
nor U6378 (N_6378,N_5656,N_5195);
nand U6379 (N_6379,N_5273,N_5568);
nor U6380 (N_6380,N_5813,N_5297);
and U6381 (N_6381,N_5821,N_5753);
or U6382 (N_6382,N_5350,N_5779);
and U6383 (N_6383,N_5607,N_5814);
nor U6384 (N_6384,N_5758,N_5144);
nand U6385 (N_6385,N_5196,N_5263);
nand U6386 (N_6386,N_5978,N_5115);
or U6387 (N_6387,N_5425,N_5550);
or U6388 (N_6388,N_5056,N_5160);
nand U6389 (N_6389,N_5909,N_5207);
nor U6390 (N_6390,N_5623,N_5865);
nor U6391 (N_6391,N_5658,N_5494);
and U6392 (N_6392,N_5628,N_5744);
nand U6393 (N_6393,N_5786,N_5242);
nand U6394 (N_6394,N_5671,N_5944);
and U6395 (N_6395,N_5301,N_5874);
or U6396 (N_6396,N_5098,N_5707);
nand U6397 (N_6397,N_5461,N_5170);
or U6398 (N_6398,N_5633,N_5895);
nand U6399 (N_6399,N_5868,N_5583);
or U6400 (N_6400,N_5622,N_5678);
nor U6401 (N_6401,N_5262,N_5536);
xnor U6402 (N_6402,N_5462,N_5084);
or U6403 (N_6403,N_5064,N_5237);
nand U6404 (N_6404,N_5320,N_5562);
nand U6405 (N_6405,N_5477,N_5300);
or U6406 (N_6406,N_5880,N_5324);
nor U6407 (N_6407,N_5776,N_5777);
nor U6408 (N_6408,N_5662,N_5134);
or U6409 (N_6409,N_5420,N_5131);
and U6410 (N_6410,N_5016,N_5126);
nand U6411 (N_6411,N_5011,N_5820);
nor U6412 (N_6412,N_5864,N_5296);
nor U6413 (N_6413,N_5340,N_5972);
and U6414 (N_6414,N_5284,N_5082);
and U6415 (N_6415,N_5817,N_5774);
and U6416 (N_6416,N_5763,N_5086);
nor U6417 (N_6417,N_5409,N_5490);
nand U6418 (N_6418,N_5645,N_5941);
or U6419 (N_6419,N_5406,N_5442);
nand U6420 (N_6420,N_5048,N_5259);
or U6421 (N_6421,N_5366,N_5140);
or U6422 (N_6422,N_5746,N_5157);
nand U6423 (N_6423,N_5430,N_5548);
nand U6424 (N_6424,N_5080,N_5933);
nor U6425 (N_6425,N_5464,N_5378);
nor U6426 (N_6426,N_5766,N_5723);
or U6427 (N_6427,N_5428,N_5139);
and U6428 (N_6428,N_5969,N_5935);
and U6429 (N_6429,N_5190,N_5826);
and U6430 (N_6430,N_5649,N_5667);
or U6431 (N_6431,N_5081,N_5825);
nor U6432 (N_6432,N_5148,N_5123);
nand U6433 (N_6433,N_5415,N_5588);
or U6434 (N_6434,N_5027,N_5967);
or U6435 (N_6435,N_5807,N_5376);
nand U6436 (N_6436,N_5401,N_5034);
and U6437 (N_6437,N_5560,N_5367);
nand U6438 (N_6438,N_5538,N_5221);
nor U6439 (N_6439,N_5998,N_5059);
or U6440 (N_6440,N_5344,N_5278);
xnor U6441 (N_6441,N_5129,N_5244);
or U6442 (N_6442,N_5747,N_5491);
or U6443 (N_6443,N_5106,N_5120);
nand U6444 (N_6444,N_5896,N_5539);
or U6445 (N_6445,N_5728,N_5283);
and U6446 (N_6446,N_5559,N_5078);
or U6447 (N_6447,N_5152,N_5939);
nand U6448 (N_6448,N_5308,N_5781);
and U6449 (N_6449,N_5109,N_5815);
nand U6450 (N_6450,N_5240,N_5432);
or U6451 (N_6451,N_5759,N_5003);
and U6452 (N_6452,N_5631,N_5004);
and U6453 (N_6453,N_5789,N_5612);
nor U6454 (N_6454,N_5444,N_5105);
or U6455 (N_6455,N_5128,N_5026);
or U6456 (N_6456,N_5624,N_5843);
nand U6457 (N_6457,N_5511,N_5076);
nor U6458 (N_6458,N_5954,N_5223);
and U6459 (N_6459,N_5859,N_5891);
nor U6460 (N_6460,N_5502,N_5618);
and U6461 (N_6461,N_5374,N_5615);
nor U6462 (N_6462,N_5077,N_5806);
and U6463 (N_6463,N_5801,N_5028);
and U6464 (N_6464,N_5289,N_5832);
and U6465 (N_6465,N_5177,N_5703);
or U6466 (N_6466,N_5383,N_5343);
or U6467 (N_6467,N_5450,N_5553);
nor U6468 (N_6468,N_5648,N_5743);
or U6469 (N_6469,N_5551,N_5799);
or U6470 (N_6470,N_5833,N_5934);
or U6471 (N_6471,N_5302,N_5785);
or U6472 (N_6472,N_5818,N_5325);
nand U6473 (N_6473,N_5861,N_5582);
nand U6474 (N_6474,N_5751,N_5355);
nor U6475 (N_6475,N_5547,N_5984);
and U6476 (N_6476,N_5351,N_5218);
and U6477 (N_6477,N_5232,N_5017);
or U6478 (N_6478,N_5974,N_5423);
nor U6479 (N_6479,N_5793,N_5647);
or U6480 (N_6480,N_5897,N_5019);
and U6481 (N_6481,N_5135,N_5455);
and U6482 (N_6482,N_5532,N_5319);
or U6483 (N_6483,N_5349,N_5075);
nor U6484 (N_6484,N_5481,N_5127);
nor U6485 (N_6485,N_5067,N_5923);
or U6486 (N_6486,N_5346,N_5439);
nand U6487 (N_6487,N_5499,N_5419);
and U6488 (N_6488,N_5849,N_5626);
xnor U6489 (N_6489,N_5586,N_5474);
nand U6490 (N_6490,N_5414,N_5796);
or U6491 (N_6491,N_5245,N_5856);
nor U6492 (N_6492,N_5169,N_5214);
nor U6493 (N_6493,N_5787,N_5362);
and U6494 (N_6494,N_5866,N_5448);
and U6495 (N_6495,N_5331,N_5676);
and U6496 (N_6496,N_5534,N_5045);
nand U6497 (N_6497,N_5318,N_5928);
nor U6498 (N_6498,N_5062,N_5791);
or U6499 (N_6499,N_5282,N_5655);
and U6500 (N_6500,N_5937,N_5052);
nor U6501 (N_6501,N_5349,N_5694);
nor U6502 (N_6502,N_5641,N_5049);
and U6503 (N_6503,N_5842,N_5409);
or U6504 (N_6504,N_5267,N_5230);
and U6505 (N_6505,N_5205,N_5167);
and U6506 (N_6506,N_5069,N_5858);
or U6507 (N_6507,N_5395,N_5708);
nor U6508 (N_6508,N_5478,N_5147);
or U6509 (N_6509,N_5168,N_5575);
nor U6510 (N_6510,N_5011,N_5777);
nand U6511 (N_6511,N_5380,N_5001);
and U6512 (N_6512,N_5898,N_5602);
nand U6513 (N_6513,N_5230,N_5234);
nand U6514 (N_6514,N_5474,N_5812);
and U6515 (N_6515,N_5568,N_5683);
nand U6516 (N_6516,N_5952,N_5214);
nor U6517 (N_6517,N_5857,N_5986);
and U6518 (N_6518,N_5332,N_5733);
nand U6519 (N_6519,N_5053,N_5190);
or U6520 (N_6520,N_5568,N_5541);
and U6521 (N_6521,N_5771,N_5944);
nor U6522 (N_6522,N_5143,N_5676);
nand U6523 (N_6523,N_5700,N_5668);
nor U6524 (N_6524,N_5949,N_5089);
nand U6525 (N_6525,N_5985,N_5960);
nor U6526 (N_6526,N_5364,N_5097);
xor U6527 (N_6527,N_5930,N_5168);
or U6528 (N_6528,N_5339,N_5478);
nor U6529 (N_6529,N_5187,N_5510);
or U6530 (N_6530,N_5103,N_5609);
xnor U6531 (N_6531,N_5563,N_5499);
nor U6532 (N_6532,N_5670,N_5206);
nor U6533 (N_6533,N_5180,N_5368);
nand U6534 (N_6534,N_5043,N_5499);
nand U6535 (N_6535,N_5917,N_5592);
nor U6536 (N_6536,N_5271,N_5000);
and U6537 (N_6537,N_5869,N_5891);
nand U6538 (N_6538,N_5597,N_5496);
nand U6539 (N_6539,N_5229,N_5118);
or U6540 (N_6540,N_5790,N_5430);
nor U6541 (N_6541,N_5064,N_5173);
and U6542 (N_6542,N_5179,N_5937);
nor U6543 (N_6543,N_5676,N_5742);
and U6544 (N_6544,N_5247,N_5686);
and U6545 (N_6545,N_5423,N_5228);
nand U6546 (N_6546,N_5310,N_5258);
and U6547 (N_6547,N_5096,N_5629);
or U6548 (N_6548,N_5156,N_5089);
nor U6549 (N_6549,N_5916,N_5859);
or U6550 (N_6550,N_5245,N_5805);
nor U6551 (N_6551,N_5863,N_5958);
nor U6552 (N_6552,N_5711,N_5139);
and U6553 (N_6553,N_5802,N_5243);
and U6554 (N_6554,N_5759,N_5851);
nor U6555 (N_6555,N_5458,N_5397);
xor U6556 (N_6556,N_5719,N_5860);
or U6557 (N_6557,N_5098,N_5260);
and U6558 (N_6558,N_5067,N_5256);
nor U6559 (N_6559,N_5650,N_5671);
and U6560 (N_6560,N_5572,N_5952);
nor U6561 (N_6561,N_5270,N_5807);
nor U6562 (N_6562,N_5580,N_5199);
or U6563 (N_6563,N_5384,N_5259);
nor U6564 (N_6564,N_5155,N_5942);
and U6565 (N_6565,N_5304,N_5656);
and U6566 (N_6566,N_5940,N_5240);
or U6567 (N_6567,N_5119,N_5245);
nand U6568 (N_6568,N_5270,N_5028);
nor U6569 (N_6569,N_5934,N_5810);
or U6570 (N_6570,N_5631,N_5229);
or U6571 (N_6571,N_5953,N_5306);
nor U6572 (N_6572,N_5054,N_5252);
and U6573 (N_6573,N_5185,N_5202);
nor U6574 (N_6574,N_5370,N_5642);
nor U6575 (N_6575,N_5204,N_5063);
nor U6576 (N_6576,N_5188,N_5748);
nor U6577 (N_6577,N_5414,N_5188);
nand U6578 (N_6578,N_5749,N_5952);
and U6579 (N_6579,N_5061,N_5543);
or U6580 (N_6580,N_5036,N_5635);
xnor U6581 (N_6581,N_5789,N_5082);
or U6582 (N_6582,N_5804,N_5778);
and U6583 (N_6583,N_5864,N_5538);
or U6584 (N_6584,N_5189,N_5900);
nand U6585 (N_6585,N_5963,N_5001);
or U6586 (N_6586,N_5569,N_5878);
and U6587 (N_6587,N_5287,N_5756);
nand U6588 (N_6588,N_5056,N_5459);
nor U6589 (N_6589,N_5546,N_5225);
or U6590 (N_6590,N_5600,N_5471);
and U6591 (N_6591,N_5766,N_5847);
nor U6592 (N_6592,N_5236,N_5298);
nand U6593 (N_6593,N_5410,N_5386);
nand U6594 (N_6594,N_5270,N_5078);
or U6595 (N_6595,N_5393,N_5466);
and U6596 (N_6596,N_5008,N_5930);
nor U6597 (N_6597,N_5409,N_5064);
or U6598 (N_6598,N_5675,N_5063);
and U6599 (N_6599,N_5520,N_5371);
nor U6600 (N_6600,N_5002,N_5954);
nor U6601 (N_6601,N_5302,N_5508);
nor U6602 (N_6602,N_5400,N_5766);
or U6603 (N_6603,N_5314,N_5831);
or U6604 (N_6604,N_5493,N_5444);
or U6605 (N_6605,N_5932,N_5146);
nand U6606 (N_6606,N_5514,N_5647);
nor U6607 (N_6607,N_5810,N_5906);
or U6608 (N_6608,N_5122,N_5716);
nor U6609 (N_6609,N_5605,N_5776);
nand U6610 (N_6610,N_5234,N_5280);
nand U6611 (N_6611,N_5063,N_5859);
nand U6612 (N_6612,N_5954,N_5744);
and U6613 (N_6613,N_5844,N_5203);
and U6614 (N_6614,N_5079,N_5675);
nor U6615 (N_6615,N_5516,N_5549);
and U6616 (N_6616,N_5021,N_5029);
or U6617 (N_6617,N_5663,N_5338);
or U6618 (N_6618,N_5837,N_5788);
nor U6619 (N_6619,N_5814,N_5764);
and U6620 (N_6620,N_5245,N_5520);
or U6621 (N_6621,N_5441,N_5704);
and U6622 (N_6622,N_5881,N_5841);
and U6623 (N_6623,N_5843,N_5577);
nor U6624 (N_6624,N_5751,N_5612);
nand U6625 (N_6625,N_5577,N_5344);
nor U6626 (N_6626,N_5706,N_5849);
and U6627 (N_6627,N_5904,N_5993);
and U6628 (N_6628,N_5203,N_5615);
nand U6629 (N_6629,N_5683,N_5720);
nor U6630 (N_6630,N_5885,N_5978);
and U6631 (N_6631,N_5909,N_5688);
or U6632 (N_6632,N_5531,N_5279);
nand U6633 (N_6633,N_5607,N_5638);
and U6634 (N_6634,N_5656,N_5260);
and U6635 (N_6635,N_5311,N_5486);
nand U6636 (N_6636,N_5017,N_5452);
and U6637 (N_6637,N_5000,N_5254);
nand U6638 (N_6638,N_5906,N_5070);
or U6639 (N_6639,N_5988,N_5639);
or U6640 (N_6640,N_5558,N_5064);
nor U6641 (N_6641,N_5972,N_5069);
nor U6642 (N_6642,N_5709,N_5293);
or U6643 (N_6643,N_5805,N_5888);
and U6644 (N_6644,N_5782,N_5356);
or U6645 (N_6645,N_5021,N_5018);
nor U6646 (N_6646,N_5003,N_5382);
nand U6647 (N_6647,N_5284,N_5460);
nor U6648 (N_6648,N_5731,N_5865);
and U6649 (N_6649,N_5946,N_5999);
and U6650 (N_6650,N_5682,N_5655);
or U6651 (N_6651,N_5181,N_5590);
and U6652 (N_6652,N_5576,N_5324);
nor U6653 (N_6653,N_5240,N_5176);
nor U6654 (N_6654,N_5705,N_5669);
and U6655 (N_6655,N_5851,N_5027);
nand U6656 (N_6656,N_5521,N_5081);
nor U6657 (N_6657,N_5777,N_5882);
nor U6658 (N_6658,N_5017,N_5994);
and U6659 (N_6659,N_5113,N_5598);
or U6660 (N_6660,N_5626,N_5168);
nor U6661 (N_6661,N_5280,N_5794);
and U6662 (N_6662,N_5933,N_5587);
nor U6663 (N_6663,N_5585,N_5571);
or U6664 (N_6664,N_5196,N_5406);
and U6665 (N_6665,N_5162,N_5364);
and U6666 (N_6666,N_5394,N_5670);
and U6667 (N_6667,N_5752,N_5801);
and U6668 (N_6668,N_5720,N_5307);
nand U6669 (N_6669,N_5480,N_5443);
and U6670 (N_6670,N_5910,N_5453);
nor U6671 (N_6671,N_5946,N_5777);
nor U6672 (N_6672,N_5820,N_5430);
nor U6673 (N_6673,N_5262,N_5294);
nand U6674 (N_6674,N_5963,N_5264);
and U6675 (N_6675,N_5083,N_5618);
nand U6676 (N_6676,N_5416,N_5086);
nor U6677 (N_6677,N_5387,N_5493);
and U6678 (N_6678,N_5039,N_5127);
nand U6679 (N_6679,N_5418,N_5715);
or U6680 (N_6680,N_5633,N_5147);
or U6681 (N_6681,N_5834,N_5642);
or U6682 (N_6682,N_5030,N_5533);
xnor U6683 (N_6683,N_5465,N_5967);
or U6684 (N_6684,N_5655,N_5896);
or U6685 (N_6685,N_5397,N_5676);
nor U6686 (N_6686,N_5540,N_5638);
nand U6687 (N_6687,N_5823,N_5877);
and U6688 (N_6688,N_5375,N_5327);
nor U6689 (N_6689,N_5468,N_5250);
nand U6690 (N_6690,N_5155,N_5085);
and U6691 (N_6691,N_5538,N_5244);
nand U6692 (N_6692,N_5733,N_5308);
or U6693 (N_6693,N_5755,N_5243);
and U6694 (N_6694,N_5766,N_5240);
or U6695 (N_6695,N_5538,N_5423);
nand U6696 (N_6696,N_5048,N_5645);
or U6697 (N_6697,N_5429,N_5686);
nor U6698 (N_6698,N_5494,N_5123);
nand U6699 (N_6699,N_5681,N_5831);
nand U6700 (N_6700,N_5577,N_5115);
nor U6701 (N_6701,N_5778,N_5450);
nand U6702 (N_6702,N_5854,N_5569);
nand U6703 (N_6703,N_5808,N_5885);
nor U6704 (N_6704,N_5292,N_5645);
or U6705 (N_6705,N_5429,N_5319);
nand U6706 (N_6706,N_5966,N_5886);
nor U6707 (N_6707,N_5806,N_5501);
or U6708 (N_6708,N_5771,N_5891);
nand U6709 (N_6709,N_5182,N_5348);
and U6710 (N_6710,N_5766,N_5326);
xor U6711 (N_6711,N_5095,N_5324);
nor U6712 (N_6712,N_5372,N_5450);
or U6713 (N_6713,N_5706,N_5285);
or U6714 (N_6714,N_5562,N_5731);
nand U6715 (N_6715,N_5439,N_5545);
and U6716 (N_6716,N_5393,N_5523);
nor U6717 (N_6717,N_5277,N_5073);
nor U6718 (N_6718,N_5162,N_5134);
or U6719 (N_6719,N_5358,N_5396);
or U6720 (N_6720,N_5235,N_5853);
and U6721 (N_6721,N_5532,N_5173);
and U6722 (N_6722,N_5276,N_5641);
and U6723 (N_6723,N_5363,N_5711);
nand U6724 (N_6724,N_5416,N_5801);
nand U6725 (N_6725,N_5126,N_5989);
nand U6726 (N_6726,N_5277,N_5760);
and U6727 (N_6727,N_5049,N_5095);
or U6728 (N_6728,N_5584,N_5764);
and U6729 (N_6729,N_5323,N_5114);
nand U6730 (N_6730,N_5795,N_5181);
nor U6731 (N_6731,N_5584,N_5085);
or U6732 (N_6732,N_5520,N_5774);
and U6733 (N_6733,N_5666,N_5712);
and U6734 (N_6734,N_5111,N_5492);
nor U6735 (N_6735,N_5824,N_5944);
nand U6736 (N_6736,N_5842,N_5440);
and U6737 (N_6737,N_5689,N_5344);
nand U6738 (N_6738,N_5229,N_5589);
and U6739 (N_6739,N_5947,N_5730);
nor U6740 (N_6740,N_5599,N_5068);
nand U6741 (N_6741,N_5349,N_5571);
or U6742 (N_6742,N_5381,N_5595);
and U6743 (N_6743,N_5172,N_5405);
nor U6744 (N_6744,N_5335,N_5623);
and U6745 (N_6745,N_5288,N_5970);
or U6746 (N_6746,N_5695,N_5381);
nand U6747 (N_6747,N_5755,N_5800);
nor U6748 (N_6748,N_5369,N_5173);
nor U6749 (N_6749,N_5129,N_5285);
and U6750 (N_6750,N_5637,N_5831);
nor U6751 (N_6751,N_5082,N_5881);
xnor U6752 (N_6752,N_5413,N_5828);
nor U6753 (N_6753,N_5503,N_5539);
or U6754 (N_6754,N_5398,N_5333);
and U6755 (N_6755,N_5417,N_5207);
or U6756 (N_6756,N_5349,N_5631);
or U6757 (N_6757,N_5086,N_5124);
and U6758 (N_6758,N_5647,N_5581);
nand U6759 (N_6759,N_5766,N_5246);
and U6760 (N_6760,N_5710,N_5882);
and U6761 (N_6761,N_5809,N_5878);
or U6762 (N_6762,N_5436,N_5162);
xnor U6763 (N_6763,N_5715,N_5294);
nor U6764 (N_6764,N_5340,N_5485);
and U6765 (N_6765,N_5626,N_5550);
nand U6766 (N_6766,N_5638,N_5117);
and U6767 (N_6767,N_5742,N_5260);
or U6768 (N_6768,N_5354,N_5630);
or U6769 (N_6769,N_5364,N_5813);
nand U6770 (N_6770,N_5865,N_5321);
nor U6771 (N_6771,N_5174,N_5410);
nor U6772 (N_6772,N_5979,N_5201);
and U6773 (N_6773,N_5259,N_5233);
nor U6774 (N_6774,N_5154,N_5096);
xor U6775 (N_6775,N_5663,N_5372);
or U6776 (N_6776,N_5611,N_5260);
or U6777 (N_6777,N_5636,N_5600);
nor U6778 (N_6778,N_5993,N_5317);
and U6779 (N_6779,N_5738,N_5051);
or U6780 (N_6780,N_5914,N_5701);
and U6781 (N_6781,N_5095,N_5931);
nor U6782 (N_6782,N_5271,N_5641);
or U6783 (N_6783,N_5478,N_5331);
and U6784 (N_6784,N_5410,N_5809);
nand U6785 (N_6785,N_5933,N_5678);
nand U6786 (N_6786,N_5539,N_5676);
and U6787 (N_6787,N_5718,N_5641);
nand U6788 (N_6788,N_5810,N_5957);
and U6789 (N_6789,N_5625,N_5611);
and U6790 (N_6790,N_5628,N_5528);
or U6791 (N_6791,N_5109,N_5313);
or U6792 (N_6792,N_5755,N_5973);
or U6793 (N_6793,N_5023,N_5132);
and U6794 (N_6794,N_5781,N_5389);
or U6795 (N_6795,N_5124,N_5788);
and U6796 (N_6796,N_5586,N_5351);
nor U6797 (N_6797,N_5843,N_5773);
and U6798 (N_6798,N_5050,N_5007);
nor U6799 (N_6799,N_5128,N_5970);
or U6800 (N_6800,N_5827,N_5500);
nor U6801 (N_6801,N_5793,N_5896);
nand U6802 (N_6802,N_5457,N_5364);
and U6803 (N_6803,N_5733,N_5451);
nor U6804 (N_6804,N_5080,N_5402);
and U6805 (N_6805,N_5963,N_5584);
and U6806 (N_6806,N_5921,N_5401);
and U6807 (N_6807,N_5597,N_5703);
and U6808 (N_6808,N_5072,N_5070);
and U6809 (N_6809,N_5906,N_5356);
nor U6810 (N_6810,N_5016,N_5393);
and U6811 (N_6811,N_5845,N_5097);
or U6812 (N_6812,N_5018,N_5870);
or U6813 (N_6813,N_5463,N_5913);
nor U6814 (N_6814,N_5673,N_5101);
nor U6815 (N_6815,N_5724,N_5282);
and U6816 (N_6816,N_5215,N_5009);
or U6817 (N_6817,N_5969,N_5560);
and U6818 (N_6818,N_5283,N_5635);
nand U6819 (N_6819,N_5356,N_5968);
xnor U6820 (N_6820,N_5627,N_5370);
nand U6821 (N_6821,N_5862,N_5132);
nor U6822 (N_6822,N_5835,N_5356);
nor U6823 (N_6823,N_5087,N_5467);
or U6824 (N_6824,N_5513,N_5022);
nor U6825 (N_6825,N_5379,N_5641);
and U6826 (N_6826,N_5039,N_5245);
and U6827 (N_6827,N_5328,N_5084);
and U6828 (N_6828,N_5091,N_5419);
nor U6829 (N_6829,N_5899,N_5719);
nand U6830 (N_6830,N_5564,N_5296);
and U6831 (N_6831,N_5441,N_5615);
nand U6832 (N_6832,N_5481,N_5980);
or U6833 (N_6833,N_5539,N_5406);
nand U6834 (N_6834,N_5854,N_5923);
nand U6835 (N_6835,N_5263,N_5916);
nand U6836 (N_6836,N_5446,N_5363);
or U6837 (N_6837,N_5326,N_5960);
or U6838 (N_6838,N_5235,N_5880);
or U6839 (N_6839,N_5176,N_5553);
nor U6840 (N_6840,N_5207,N_5996);
nand U6841 (N_6841,N_5045,N_5103);
nand U6842 (N_6842,N_5161,N_5830);
or U6843 (N_6843,N_5775,N_5450);
xor U6844 (N_6844,N_5629,N_5842);
and U6845 (N_6845,N_5585,N_5150);
nand U6846 (N_6846,N_5717,N_5715);
nor U6847 (N_6847,N_5282,N_5441);
nand U6848 (N_6848,N_5710,N_5211);
nand U6849 (N_6849,N_5541,N_5095);
nor U6850 (N_6850,N_5932,N_5377);
nor U6851 (N_6851,N_5160,N_5625);
nand U6852 (N_6852,N_5433,N_5870);
nor U6853 (N_6853,N_5586,N_5279);
nor U6854 (N_6854,N_5106,N_5771);
nand U6855 (N_6855,N_5853,N_5188);
nor U6856 (N_6856,N_5695,N_5698);
nand U6857 (N_6857,N_5423,N_5408);
and U6858 (N_6858,N_5578,N_5755);
or U6859 (N_6859,N_5686,N_5713);
nor U6860 (N_6860,N_5946,N_5695);
nand U6861 (N_6861,N_5506,N_5456);
nand U6862 (N_6862,N_5217,N_5102);
nor U6863 (N_6863,N_5090,N_5433);
nor U6864 (N_6864,N_5785,N_5209);
or U6865 (N_6865,N_5992,N_5670);
and U6866 (N_6866,N_5473,N_5121);
nand U6867 (N_6867,N_5697,N_5396);
and U6868 (N_6868,N_5576,N_5777);
or U6869 (N_6869,N_5537,N_5805);
and U6870 (N_6870,N_5492,N_5902);
or U6871 (N_6871,N_5300,N_5892);
and U6872 (N_6872,N_5169,N_5277);
and U6873 (N_6873,N_5749,N_5469);
and U6874 (N_6874,N_5492,N_5681);
and U6875 (N_6875,N_5603,N_5263);
or U6876 (N_6876,N_5745,N_5389);
nor U6877 (N_6877,N_5762,N_5765);
and U6878 (N_6878,N_5083,N_5600);
nand U6879 (N_6879,N_5107,N_5244);
or U6880 (N_6880,N_5795,N_5810);
or U6881 (N_6881,N_5194,N_5770);
and U6882 (N_6882,N_5999,N_5874);
and U6883 (N_6883,N_5354,N_5492);
nor U6884 (N_6884,N_5478,N_5355);
or U6885 (N_6885,N_5281,N_5094);
nand U6886 (N_6886,N_5423,N_5762);
nor U6887 (N_6887,N_5413,N_5541);
nand U6888 (N_6888,N_5989,N_5400);
and U6889 (N_6889,N_5828,N_5886);
nand U6890 (N_6890,N_5001,N_5363);
nor U6891 (N_6891,N_5389,N_5247);
nor U6892 (N_6892,N_5263,N_5443);
and U6893 (N_6893,N_5112,N_5381);
and U6894 (N_6894,N_5079,N_5151);
nand U6895 (N_6895,N_5129,N_5571);
or U6896 (N_6896,N_5866,N_5019);
nor U6897 (N_6897,N_5719,N_5465);
nand U6898 (N_6898,N_5449,N_5588);
or U6899 (N_6899,N_5577,N_5398);
and U6900 (N_6900,N_5819,N_5632);
and U6901 (N_6901,N_5037,N_5665);
or U6902 (N_6902,N_5616,N_5829);
nand U6903 (N_6903,N_5970,N_5258);
nand U6904 (N_6904,N_5132,N_5935);
nor U6905 (N_6905,N_5402,N_5421);
and U6906 (N_6906,N_5068,N_5931);
nor U6907 (N_6907,N_5401,N_5722);
and U6908 (N_6908,N_5516,N_5220);
nand U6909 (N_6909,N_5262,N_5617);
nor U6910 (N_6910,N_5605,N_5172);
and U6911 (N_6911,N_5051,N_5197);
nor U6912 (N_6912,N_5782,N_5105);
or U6913 (N_6913,N_5705,N_5415);
and U6914 (N_6914,N_5136,N_5007);
or U6915 (N_6915,N_5918,N_5825);
or U6916 (N_6916,N_5294,N_5047);
and U6917 (N_6917,N_5177,N_5372);
nor U6918 (N_6918,N_5769,N_5694);
nor U6919 (N_6919,N_5226,N_5597);
nor U6920 (N_6920,N_5448,N_5059);
nand U6921 (N_6921,N_5971,N_5043);
and U6922 (N_6922,N_5367,N_5176);
nand U6923 (N_6923,N_5612,N_5998);
or U6924 (N_6924,N_5328,N_5057);
nand U6925 (N_6925,N_5089,N_5846);
nand U6926 (N_6926,N_5460,N_5644);
or U6927 (N_6927,N_5866,N_5718);
or U6928 (N_6928,N_5571,N_5111);
or U6929 (N_6929,N_5130,N_5768);
nand U6930 (N_6930,N_5700,N_5305);
nand U6931 (N_6931,N_5930,N_5389);
nand U6932 (N_6932,N_5248,N_5317);
or U6933 (N_6933,N_5659,N_5540);
or U6934 (N_6934,N_5722,N_5063);
nand U6935 (N_6935,N_5623,N_5032);
or U6936 (N_6936,N_5022,N_5999);
and U6937 (N_6937,N_5356,N_5311);
and U6938 (N_6938,N_5384,N_5717);
nor U6939 (N_6939,N_5181,N_5115);
nor U6940 (N_6940,N_5676,N_5528);
nor U6941 (N_6941,N_5313,N_5461);
or U6942 (N_6942,N_5563,N_5946);
and U6943 (N_6943,N_5039,N_5784);
or U6944 (N_6944,N_5716,N_5217);
or U6945 (N_6945,N_5665,N_5485);
and U6946 (N_6946,N_5683,N_5184);
nor U6947 (N_6947,N_5005,N_5749);
and U6948 (N_6948,N_5092,N_5049);
xnor U6949 (N_6949,N_5749,N_5720);
and U6950 (N_6950,N_5227,N_5679);
and U6951 (N_6951,N_5673,N_5136);
or U6952 (N_6952,N_5287,N_5129);
nor U6953 (N_6953,N_5687,N_5035);
nand U6954 (N_6954,N_5893,N_5708);
nand U6955 (N_6955,N_5752,N_5159);
nand U6956 (N_6956,N_5500,N_5774);
nand U6957 (N_6957,N_5867,N_5651);
nor U6958 (N_6958,N_5465,N_5836);
and U6959 (N_6959,N_5757,N_5975);
nor U6960 (N_6960,N_5260,N_5225);
nor U6961 (N_6961,N_5723,N_5852);
xnor U6962 (N_6962,N_5513,N_5351);
nand U6963 (N_6963,N_5887,N_5338);
nor U6964 (N_6964,N_5901,N_5350);
nor U6965 (N_6965,N_5816,N_5673);
nor U6966 (N_6966,N_5594,N_5476);
nor U6967 (N_6967,N_5112,N_5949);
and U6968 (N_6968,N_5668,N_5958);
and U6969 (N_6969,N_5440,N_5547);
and U6970 (N_6970,N_5055,N_5276);
or U6971 (N_6971,N_5247,N_5562);
nor U6972 (N_6972,N_5343,N_5160);
nand U6973 (N_6973,N_5259,N_5226);
and U6974 (N_6974,N_5686,N_5423);
nand U6975 (N_6975,N_5394,N_5509);
nor U6976 (N_6976,N_5391,N_5877);
nor U6977 (N_6977,N_5735,N_5501);
nand U6978 (N_6978,N_5095,N_5397);
nor U6979 (N_6979,N_5033,N_5149);
or U6980 (N_6980,N_5638,N_5094);
and U6981 (N_6981,N_5559,N_5940);
and U6982 (N_6982,N_5563,N_5117);
and U6983 (N_6983,N_5444,N_5396);
nand U6984 (N_6984,N_5184,N_5575);
nor U6985 (N_6985,N_5708,N_5644);
and U6986 (N_6986,N_5194,N_5957);
or U6987 (N_6987,N_5337,N_5687);
and U6988 (N_6988,N_5534,N_5646);
or U6989 (N_6989,N_5735,N_5328);
xnor U6990 (N_6990,N_5790,N_5673);
xor U6991 (N_6991,N_5922,N_5083);
nor U6992 (N_6992,N_5313,N_5698);
or U6993 (N_6993,N_5375,N_5334);
nor U6994 (N_6994,N_5242,N_5798);
and U6995 (N_6995,N_5525,N_5056);
nand U6996 (N_6996,N_5996,N_5915);
nor U6997 (N_6997,N_5819,N_5072);
nand U6998 (N_6998,N_5887,N_5364);
nand U6999 (N_6999,N_5937,N_5320);
nand U7000 (N_7000,N_6140,N_6189);
and U7001 (N_7001,N_6495,N_6577);
nor U7002 (N_7002,N_6070,N_6408);
or U7003 (N_7003,N_6736,N_6347);
or U7004 (N_7004,N_6034,N_6953);
nor U7005 (N_7005,N_6267,N_6298);
nor U7006 (N_7006,N_6066,N_6321);
or U7007 (N_7007,N_6925,N_6669);
nand U7008 (N_7008,N_6633,N_6843);
and U7009 (N_7009,N_6053,N_6875);
nand U7010 (N_7010,N_6046,N_6162);
and U7011 (N_7011,N_6338,N_6793);
or U7012 (N_7012,N_6651,N_6294);
or U7013 (N_7013,N_6429,N_6625);
nor U7014 (N_7014,N_6454,N_6261);
and U7015 (N_7015,N_6404,N_6750);
or U7016 (N_7016,N_6753,N_6616);
and U7017 (N_7017,N_6782,N_6710);
nor U7018 (N_7018,N_6342,N_6693);
nor U7019 (N_7019,N_6412,N_6075);
nor U7020 (N_7020,N_6500,N_6292);
or U7021 (N_7021,N_6557,N_6738);
or U7022 (N_7022,N_6808,N_6584);
or U7023 (N_7023,N_6526,N_6993);
and U7024 (N_7024,N_6688,N_6135);
or U7025 (N_7025,N_6871,N_6825);
xor U7026 (N_7026,N_6927,N_6932);
nor U7027 (N_7027,N_6388,N_6835);
or U7028 (N_7028,N_6546,N_6804);
xor U7029 (N_7029,N_6987,N_6494);
nand U7030 (N_7030,N_6097,N_6703);
nor U7031 (N_7031,N_6837,N_6992);
and U7032 (N_7032,N_6854,N_6354);
and U7033 (N_7033,N_6439,N_6905);
and U7034 (N_7034,N_6886,N_6205);
nor U7035 (N_7035,N_6620,N_6493);
and U7036 (N_7036,N_6296,N_6801);
and U7037 (N_7037,N_6374,N_6184);
or U7038 (N_7038,N_6779,N_6107);
nor U7039 (N_7039,N_6085,N_6402);
nor U7040 (N_7040,N_6972,N_6483);
nand U7041 (N_7041,N_6155,N_6446);
or U7042 (N_7042,N_6605,N_6131);
nor U7043 (N_7043,N_6502,N_6910);
and U7044 (N_7044,N_6436,N_6885);
nand U7045 (N_7045,N_6365,N_6626);
nand U7046 (N_7046,N_6563,N_6776);
and U7047 (N_7047,N_6799,N_6040);
nor U7048 (N_7048,N_6105,N_6924);
or U7049 (N_7049,N_6274,N_6441);
nand U7050 (N_7050,N_6806,N_6028);
nand U7051 (N_7051,N_6878,N_6552);
nor U7052 (N_7052,N_6132,N_6055);
nor U7053 (N_7053,N_6550,N_6985);
or U7054 (N_7054,N_6676,N_6218);
nor U7055 (N_7055,N_6424,N_6283);
and U7056 (N_7056,N_6571,N_6369);
nand U7057 (N_7057,N_6008,N_6513);
or U7058 (N_7058,N_6694,N_6948);
or U7059 (N_7059,N_6265,N_6718);
or U7060 (N_7060,N_6371,N_6826);
nor U7061 (N_7061,N_6101,N_6514);
nor U7062 (N_7062,N_6348,N_6252);
nor U7063 (N_7063,N_6963,N_6504);
and U7064 (N_7064,N_6401,N_6870);
and U7065 (N_7065,N_6095,N_6790);
and U7066 (N_7066,N_6057,N_6848);
and U7067 (N_7067,N_6312,N_6244);
or U7068 (N_7068,N_6376,N_6734);
or U7069 (N_7069,N_6512,N_6645);
nand U7070 (N_7070,N_6813,N_6456);
or U7071 (N_7071,N_6364,N_6974);
xnor U7072 (N_7072,N_6938,N_6781);
and U7073 (N_7073,N_6959,N_6181);
nand U7074 (N_7074,N_6355,N_6481);
or U7075 (N_7075,N_6982,N_6224);
nor U7076 (N_7076,N_6907,N_6467);
or U7077 (N_7077,N_6064,N_6275);
or U7078 (N_7078,N_6197,N_6295);
xor U7079 (N_7079,N_6358,N_6247);
or U7080 (N_7080,N_6145,N_6153);
and U7081 (N_7081,N_6964,N_6702);
nor U7082 (N_7082,N_6035,N_6920);
nor U7083 (N_7083,N_6524,N_6721);
and U7084 (N_7084,N_6683,N_6003);
nand U7085 (N_7085,N_6262,N_6660);
nand U7086 (N_7086,N_6742,N_6989);
nor U7087 (N_7087,N_6233,N_6478);
and U7088 (N_7088,N_6036,N_6735);
nand U7089 (N_7089,N_6328,N_6484);
xor U7090 (N_7090,N_6007,N_6450);
or U7091 (N_7091,N_6919,N_6444);
or U7092 (N_7092,N_6531,N_6600);
and U7093 (N_7093,N_6780,N_6178);
or U7094 (N_7094,N_6293,N_6892);
and U7095 (N_7095,N_6316,N_6027);
or U7096 (N_7096,N_6350,N_6739);
and U7097 (N_7097,N_6990,N_6640);
xor U7098 (N_7098,N_6148,N_6667);
and U7099 (N_7099,N_6241,N_6186);
and U7100 (N_7100,N_6277,N_6949);
or U7101 (N_7101,N_6713,N_6593);
nor U7102 (N_7102,N_6379,N_6157);
and U7103 (N_7103,N_6315,N_6544);
and U7104 (N_7104,N_6111,N_6980);
or U7105 (N_7105,N_6006,N_6209);
nor U7106 (N_7106,N_6333,N_6406);
or U7107 (N_7107,N_6706,N_6015);
and U7108 (N_7108,N_6290,N_6849);
or U7109 (N_7109,N_6615,N_6921);
or U7110 (N_7110,N_6319,N_6193);
nand U7111 (N_7111,N_6324,N_6161);
nor U7112 (N_7112,N_6856,N_6462);
nor U7113 (N_7113,N_6597,N_6395);
or U7114 (N_7114,N_6682,N_6226);
nand U7115 (N_7115,N_6438,N_6941);
or U7116 (N_7116,N_6672,N_6863);
nor U7117 (N_7117,N_6448,N_6955);
nor U7118 (N_7118,N_6665,N_6582);
nand U7119 (N_7119,N_6847,N_6983);
nor U7120 (N_7120,N_6872,N_6175);
nand U7121 (N_7121,N_6213,N_6929);
nor U7122 (N_7122,N_6271,N_6398);
or U7123 (N_7123,N_6819,N_6426);
nor U7124 (N_7124,N_6033,N_6889);
or U7125 (N_7125,N_6332,N_6092);
nand U7126 (N_7126,N_6908,N_6760);
and U7127 (N_7127,N_6463,N_6177);
nor U7128 (N_7128,N_6857,N_6881);
nand U7129 (N_7129,N_6081,N_6420);
or U7130 (N_7130,N_6530,N_6630);
or U7131 (N_7131,N_6746,N_6657);
or U7132 (N_7132,N_6010,N_6896);
nand U7133 (N_7133,N_6535,N_6000);
or U7134 (N_7134,N_6748,N_6063);
nor U7135 (N_7135,N_6270,N_6216);
nand U7136 (N_7136,N_6134,N_6680);
and U7137 (N_7137,N_6701,N_6268);
nand U7138 (N_7138,N_6491,N_6390);
or U7139 (N_7139,N_6166,N_6897);
nor U7140 (N_7140,N_6805,N_6545);
nand U7141 (N_7141,N_6926,N_6138);
and U7142 (N_7142,N_6818,N_6062);
and U7143 (N_7143,N_6414,N_6147);
and U7144 (N_7144,N_6740,N_6477);
nor U7145 (N_7145,N_6343,N_6789);
and U7146 (N_7146,N_6698,N_6384);
and U7147 (N_7147,N_6664,N_6998);
or U7148 (N_7148,N_6098,N_6048);
and U7149 (N_7149,N_6588,N_6565);
nor U7150 (N_7150,N_6966,N_6188);
or U7151 (N_7151,N_6995,N_6278);
nand U7152 (N_7152,N_6018,N_6853);
or U7153 (N_7153,N_6637,N_6418);
or U7154 (N_7154,N_6641,N_6833);
and U7155 (N_7155,N_6410,N_6173);
and U7156 (N_7156,N_6263,N_6564);
nor U7157 (N_7157,N_6204,N_6472);
nand U7158 (N_7158,N_6014,N_6044);
or U7159 (N_7159,N_6662,N_6093);
nor U7160 (N_7160,N_6827,N_6538);
nand U7161 (N_7161,N_6215,N_6503);
nand U7162 (N_7162,N_6747,N_6023);
and U7163 (N_7163,N_6841,N_6944);
or U7164 (N_7164,N_6834,N_6203);
nand U7165 (N_7165,N_6668,N_6936);
nand U7166 (N_7166,N_6136,N_6970);
and U7167 (N_7167,N_6457,N_6126);
nor U7168 (N_7168,N_6214,N_6560);
nand U7169 (N_7169,N_6422,N_6671);
nor U7170 (N_7170,N_6225,N_6172);
nor U7171 (N_7171,N_6150,N_6898);
nand U7172 (N_7172,N_6783,N_6470);
nand U7173 (N_7173,N_6729,N_6069);
nor U7174 (N_7174,N_6976,N_6345);
nor U7175 (N_7175,N_6182,N_6221);
or U7176 (N_7176,N_6466,N_6967);
nand U7177 (N_7177,N_6796,N_6077);
nand U7178 (N_7178,N_6143,N_6643);
and U7179 (N_7179,N_6187,N_6639);
and U7180 (N_7180,N_6961,N_6471);
nor U7181 (N_7181,N_6958,N_6823);
or U7182 (N_7182,N_6285,N_6373);
nand U7183 (N_7183,N_6722,N_6541);
nor U7184 (N_7184,N_6720,N_6845);
or U7185 (N_7185,N_6874,N_6752);
nor U7186 (N_7186,N_6501,N_6918);
nand U7187 (N_7187,N_6956,N_6527);
nand U7188 (N_7188,N_6393,N_6231);
or U7189 (N_7189,N_6579,N_6762);
nor U7190 (N_7190,N_6540,N_6712);
and U7191 (N_7191,N_6968,N_6297);
nand U7192 (N_7192,N_6844,N_6674);
nand U7193 (N_7193,N_6673,N_6542);
or U7194 (N_7194,N_6442,N_6201);
xor U7195 (N_7195,N_6074,N_6902);
nand U7196 (N_7196,N_6239,N_6330);
and U7197 (N_7197,N_6962,N_6122);
and U7198 (N_7198,N_6852,N_6585);
nand U7199 (N_7199,N_6128,N_6230);
and U7200 (N_7200,N_6289,N_6159);
or U7201 (N_7201,N_6287,N_6777);
and U7202 (N_7202,N_6026,N_6476);
and U7203 (N_7203,N_6340,N_6228);
nor U7204 (N_7204,N_6096,N_6891);
or U7205 (N_7205,N_6025,N_6430);
and U7206 (N_7206,N_6427,N_6211);
nand U7207 (N_7207,N_6650,N_6496);
nand U7208 (N_7208,N_6490,N_6409);
and U7209 (N_7209,N_6709,N_6334);
or U7210 (N_7210,N_6784,N_6519);
nor U7211 (N_7211,N_6733,N_6183);
nand U7212 (N_7212,N_6125,N_6685);
nor U7213 (N_7213,N_6679,N_6573);
xor U7214 (N_7214,N_6191,N_6217);
nor U7215 (N_7215,N_6914,N_6807);
nor U7216 (N_7216,N_6730,N_6952);
nand U7217 (N_7217,N_6696,N_6254);
nand U7218 (N_7218,N_6774,N_6016);
and U7219 (N_7219,N_6725,N_6004);
nand U7220 (N_7220,N_6031,N_6485);
nand U7221 (N_7221,N_6200,N_6618);
nand U7222 (N_7222,N_6836,N_6264);
nor U7223 (N_7223,N_6583,N_6802);
nor U7224 (N_7224,N_6558,N_6407);
or U7225 (N_7225,N_6460,N_6829);
and U7226 (N_7226,N_6115,N_6121);
nand U7227 (N_7227,N_6094,N_6243);
and U7228 (N_7228,N_6634,N_6359);
or U7229 (N_7229,N_6242,N_6435);
nand U7230 (N_7230,N_6341,N_6307);
nor U7231 (N_7231,N_6220,N_6603);
or U7232 (N_7232,N_6509,N_6876);
nor U7233 (N_7233,N_6492,N_6366);
or U7234 (N_7234,N_6386,N_6144);
nor U7235 (N_7235,N_6459,N_6598);
and U7236 (N_7236,N_6475,N_6771);
nand U7237 (N_7237,N_6912,N_6595);
xnor U7238 (N_7238,N_6656,N_6528);
or U7239 (N_7239,N_6288,N_6377);
nand U7240 (N_7240,N_6991,N_6440);
nand U7241 (N_7241,N_6786,N_6934);
nor U7242 (N_7242,N_6068,N_6576);
nand U7243 (N_7243,N_6689,N_6434);
nand U7244 (N_7244,N_6282,N_6346);
or U7245 (N_7245,N_6511,N_6417);
nand U7246 (N_7246,N_6488,N_6971);
and U7247 (N_7247,N_6447,N_6482);
and U7248 (N_7248,N_6001,N_6719);
nand U7249 (N_7249,N_6102,N_6078);
nand U7250 (N_7250,N_6864,N_6516);
and U7251 (N_7251,N_6916,N_6553);
nand U7252 (N_7252,N_6965,N_6562);
nand U7253 (N_7253,N_6032,N_6272);
nor U7254 (N_7254,N_6794,N_6723);
xor U7255 (N_7255,N_6761,N_6058);
and U7256 (N_7256,N_6380,N_6325);
nand U7257 (N_7257,N_6899,N_6116);
and U7258 (N_7258,N_6627,N_6104);
and U7259 (N_7259,N_6568,N_6318);
and U7260 (N_7260,N_6717,N_6691);
nand U7261 (N_7261,N_6362,N_6869);
or U7262 (N_7262,N_6399,N_6291);
or U7263 (N_7263,N_6950,N_6590);
nor U7264 (N_7264,N_6419,N_6704);
and U7265 (N_7265,N_6745,N_6821);
or U7266 (N_7266,N_6711,N_6151);
nor U7267 (N_7267,N_6253,N_6146);
nand U7268 (N_7268,N_6310,N_6969);
or U7269 (N_7269,N_6909,N_6561);
or U7270 (N_7270,N_6529,N_6397);
or U7271 (N_7271,N_6309,N_6769);
nand U7272 (N_7272,N_6049,N_6798);
and U7273 (N_7273,N_6403,N_6154);
xnor U7274 (N_7274,N_6273,N_6065);
and U7275 (N_7275,N_6222,N_6108);
xor U7276 (N_7276,N_6613,N_6185);
nor U7277 (N_7277,N_6661,N_6533);
nand U7278 (N_7278,N_6587,N_6363);
and U7279 (N_7279,N_6946,N_6707);
and U7280 (N_7280,N_6867,N_6570);
and U7281 (N_7281,N_6644,N_6269);
or U7282 (N_7282,N_6522,N_6208);
and U7283 (N_7283,N_6601,N_6594);
nand U7284 (N_7284,N_6756,N_6778);
nor U7285 (N_7285,N_6659,N_6280);
and U7286 (N_7286,N_6022,N_6973);
nand U7287 (N_7287,N_6368,N_6009);
or U7288 (N_7288,N_6002,N_6432);
nand U7289 (N_7289,N_6019,N_6056);
nor U7290 (N_7290,N_6817,N_6050);
nand U7291 (N_7291,N_6168,N_6591);
and U7292 (N_7292,N_6250,N_6809);
nor U7293 (N_7293,N_6089,N_6631);
nand U7294 (N_7294,N_6619,N_6517);
nor U7295 (N_7295,N_6917,N_6716);
or U7296 (N_7296,N_6383,N_6795);
or U7297 (N_7297,N_6549,N_6286);
nor U7298 (N_7298,N_6830,N_6678);
nand U7299 (N_7299,N_6327,N_6556);
nand U7300 (N_7300,N_6791,N_6523);
or U7301 (N_7301,N_6532,N_6339);
or U7302 (N_7302,N_6862,N_6389);
and U7303 (N_7303,N_6411,N_6083);
or U7304 (N_7304,N_6127,N_6797);
nor U7305 (N_7305,N_6114,N_6884);
and U7306 (N_7306,N_6306,N_6329);
nor U7307 (N_7307,N_6978,N_6913);
nor U7308 (N_7308,N_6012,N_6951);
or U7309 (N_7309,N_6349,N_6117);
nor U7310 (N_7310,N_6646,N_6464);
nor U7311 (N_7311,N_6937,N_6113);
nand U7312 (N_7312,N_6455,N_6106);
and U7313 (N_7313,N_6163,N_6405);
nand U7314 (N_7314,N_6248,N_6653);
nor U7315 (N_7315,N_6041,N_6785);
nand U7316 (N_7316,N_6842,N_6604);
or U7317 (N_7317,N_6638,N_6473);
nor U7318 (N_7318,N_6690,N_6137);
nor U7319 (N_7319,N_6882,N_6303);
nor U7320 (N_7320,N_6566,N_6822);
nand U7321 (N_7321,N_6624,N_6623);
nor U7322 (N_7322,N_6816,N_6235);
and U7323 (N_7323,N_6589,N_6534);
and U7324 (N_7324,N_6751,N_6947);
or U7325 (N_7325,N_6569,N_6423);
or U7326 (N_7326,N_6812,N_6815);
and U7327 (N_7327,N_6728,N_6610);
nor U7328 (N_7328,N_6787,N_6652);
and U7329 (N_7329,N_6520,N_6317);
and U7330 (N_7330,N_6120,N_6505);
or U7331 (N_7331,N_6479,N_6960);
nor U7332 (N_7332,N_6675,N_6536);
or U7333 (N_7333,N_6042,N_6428);
or U7334 (N_7334,N_6764,N_6635);
and U7335 (N_7335,N_6110,N_6606);
nand U7336 (N_7336,N_6090,N_6803);
or U7337 (N_7337,N_6773,N_6465);
or U7338 (N_7338,N_6452,N_6086);
nand U7339 (N_7339,N_6612,N_6957);
nor U7340 (N_7340,N_6547,N_6893);
nor U7341 (N_7341,N_6904,N_6212);
or U7342 (N_7342,N_6883,N_6586);
nor U7343 (N_7343,N_6737,N_6416);
nor U7344 (N_7344,N_6999,N_6234);
nor U7345 (N_7345,N_6431,N_6109);
nand U7346 (N_7346,N_6614,N_6301);
nand U7347 (N_7347,N_6846,N_6394);
and U7348 (N_7348,N_6194,N_6602);
and U7349 (N_7349,N_6940,N_6179);
and U7350 (N_7350,N_6988,N_6986);
or U7351 (N_7351,N_6979,N_6020);
nand U7352 (N_7352,N_6381,N_6017);
and U7353 (N_7353,N_6352,N_6119);
or U7354 (N_7354,N_6013,N_6831);
nor U7355 (N_7355,N_6578,N_6572);
nor U7356 (N_7356,N_6498,N_6305);
or U7357 (N_7357,N_6887,N_6130);
and U7358 (N_7358,N_6326,N_6024);
xor U7359 (N_7359,N_6911,N_6581);
and U7360 (N_7360,N_6385,N_6543);
and U7361 (N_7361,N_6903,N_6219);
and U7362 (N_7362,N_6039,N_6284);
or U7363 (N_7363,N_6067,N_6169);
nor U7364 (N_7364,N_6072,N_6029);
or U7365 (N_7365,N_6888,N_6087);
and U7366 (N_7366,N_6890,N_6480);
nor U7367 (N_7367,N_6344,N_6060);
nand U7368 (N_7368,N_6198,N_6915);
and U7369 (N_7369,N_6684,N_6775);
and U7370 (N_7370,N_6567,N_6859);
nor U7371 (N_7371,N_6866,N_6763);
or U7372 (N_7372,N_6508,N_6715);
nand U7373 (N_7373,N_6458,N_6839);
or U7374 (N_7374,N_6400,N_6199);
nand U7375 (N_7375,N_6592,N_6256);
or U7376 (N_7376,N_6596,N_6170);
nor U7377 (N_7377,N_6861,N_6037);
or U7378 (N_7378,N_6375,N_6206);
nand U7379 (N_7379,N_6084,N_6336);
nor U7380 (N_7380,N_6099,N_6810);
nor U7381 (N_7381,N_6320,N_6335);
and U7382 (N_7382,N_6433,N_6621);
or U7383 (N_7383,N_6900,N_6071);
xor U7384 (N_7384,N_6202,N_6337);
nor U7385 (N_7385,N_6415,N_6164);
nor U7386 (N_7386,N_6840,N_6832);
nand U7387 (N_7387,N_6931,N_6190);
nor U7388 (N_7388,N_6323,N_6061);
nor U7389 (N_7389,N_6757,N_6497);
nor U7390 (N_7390,N_6895,N_6539);
nand U7391 (N_7391,N_6311,N_6677);
or U7392 (N_7392,N_6873,N_6636);
or U7393 (N_7393,N_6628,N_6043);
nand U7394 (N_7394,N_6518,N_6954);
nand U7395 (N_7395,N_6192,N_6975);
nand U7396 (N_7396,N_6575,N_6554);
nor U7397 (N_7397,N_6894,N_6227);
nor U7398 (N_7398,N_6741,N_6788);
nor U7399 (N_7399,N_6647,N_6824);
or U7400 (N_7400,N_6977,N_6744);
nor U7401 (N_7401,N_6580,N_6331);
or U7402 (N_7402,N_6814,N_6489);
and U7403 (N_7403,N_6877,N_6850);
nor U7404 (N_7404,N_6160,N_6445);
or U7405 (N_7405,N_6670,N_6207);
xnor U7406 (N_7406,N_6129,N_6302);
or U7407 (N_7407,N_6149,N_6076);
or U7408 (N_7408,N_6724,N_6167);
or U7409 (N_7409,N_6632,N_6743);
and U7410 (N_7410,N_6054,N_6361);
or U7411 (N_7411,N_6642,N_6906);
nand U7412 (N_7412,N_6051,N_6353);
or U7413 (N_7413,N_6142,N_6767);
or U7414 (N_7414,N_6755,N_6382);
nand U7415 (N_7415,N_6052,N_6073);
and U7416 (N_7416,N_6608,N_6141);
and U7417 (N_7417,N_6158,N_6469);
nor U7418 (N_7418,N_6663,N_6091);
or U7419 (N_7419,N_6981,N_6468);
or U7420 (N_7420,N_6727,N_6708);
or U7421 (N_7421,N_6654,N_6360);
nand U7422 (N_7422,N_6240,N_6259);
nor U7423 (N_7423,N_6487,N_6139);
nor U7424 (N_7424,N_6928,N_6768);
xnor U7425 (N_7425,N_6506,N_6515);
and U7426 (N_7426,N_6123,N_6370);
nor U7427 (N_7427,N_6387,N_6666);
and U7428 (N_7428,N_6997,N_6421);
nor U7429 (N_7429,N_6372,N_6011);
nor U7430 (N_7430,N_6942,N_6700);
nor U7431 (N_7431,N_6555,N_6599);
nand U7432 (N_7432,N_6299,N_6437);
or U7433 (N_7433,N_6443,N_6021);
and U7434 (N_7434,N_6658,N_6229);
and U7435 (N_7435,N_6695,N_6266);
or U7436 (N_7436,N_6521,N_6629);
nand U7437 (N_7437,N_6223,N_6461);
or U7438 (N_7438,N_6935,N_6367);
nor U7439 (N_7439,N_6868,N_6322);
xor U7440 (N_7440,N_6655,N_6766);
or U7441 (N_7441,N_6171,N_6257);
nor U7442 (N_7442,N_6574,N_6922);
and U7443 (N_7443,N_6196,N_6314);
nand U7444 (N_7444,N_6103,N_6047);
nand U7445 (N_7445,N_6237,N_6260);
nand U7446 (N_7446,N_6609,N_6879);
and U7447 (N_7447,N_6697,N_6537);
or U7448 (N_7448,N_6249,N_6548);
and U7449 (N_7449,N_6943,N_6692);
nand U7450 (N_7450,N_6300,N_6617);
or U7451 (N_7451,N_6754,N_6939);
nand U7452 (N_7452,N_6732,N_6276);
or U7453 (N_7453,N_6686,N_6770);
or U7454 (N_7454,N_6118,N_6486);
or U7455 (N_7455,N_6232,N_6152);
nor U7456 (N_7456,N_6313,N_6030);
and U7457 (N_7457,N_6923,N_6758);
and U7458 (N_7458,N_6174,N_6378);
nor U7459 (N_7459,N_6392,N_6238);
and U7460 (N_7460,N_6251,N_6765);
nand U7461 (N_7461,N_6124,N_6525);
or U7462 (N_7462,N_6945,N_6100);
or U7463 (N_7463,N_6156,N_6996);
nor U7464 (N_7464,N_6255,N_6855);
and U7465 (N_7465,N_6681,N_6749);
nor U7466 (N_7466,N_6792,N_6507);
nor U7467 (N_7467,N_6699,N_6731);
nor U7468 (N_7468,N_6357,N_6279);
or U7469 (N_7469,N_6082,N_6930);
and U7470 (N_7470,N_6112,N_6451);
or U7471 (N_7471,N_6246,N_6611);
nand U7472 (N_7472,N_6705,N_6005);
and U7473 (N_7473,N_6391,N_6258);
nand U7474 (N_7474,N_6648,N_6649);
and U7475 (N_7475,N_6281,N_6820);
and U7476 (N_7476,N_6133,N_6180);
or U7477 (N_7477,N_6045,N_6838);
and U7478 (N_7478,N_6860,N_6811);
and U7479 (N_7479,N_6088,N_6994);
nor U7480 (N_7480,N_6851,N_6080);
or U7481 (N_7481,N_6499,N_6059);
and U7482 (N_7482,N_6984,N_6165);
or U7483 (N_7483,N_6714,N_6356);
and U7484 (N_7484,N_6474,N_6236);
nor U7485 (N_7485,N_6726,N_6622);
nor U7486 (N_7486,N_6828,N_6304);
or U7487 (N_7487,N_6858,N_6901);
and U7488 (N_7488,N_6510,N_6800);
nor U7489 (N_7489,N_6351,N_6425);
nand U7490 (N_7490,N_6687,N_6079);
nand U7491 (N_7491,N_6210,N_6759);
xnor U7492 (N_7492,N_6453,N_6880);
or U7493 (N_7493,N_6772,N_6038);
nand U7494 (N_7494,N_6308,N_6865);
or U7495 (N_7495,N_6413,N_6176);
nand U7496 (N_7496,N_6195,N_6551);
or U7497 (N_7497,N_6396,N_6245);
and U7498 (N_7498,N_6559,N_6607);
and U7499 (N_7499,N_6933,N_6449);
or U7500 (N_7500,N_6446,N_6923);
or U7501 (N_7501,N_6818,N_6884);
or U7502 (N_7502,N_6745,N_6716);
nor U7503 (N_7503,N_6677,N_6672);
and U7504 (N_7504,N_6833,N_6119);
nor U7505 (N_7505,N_6719,N_6503);
nand U7506 (N_7506,N_6936,N_6401);
or U7507 (N_7507,N_6622,N_6578);
nand U7508 (N_7508,N_6354,N_6667);
or U7509 (N_7509,N_6303,N_6633);
nor U7510 (N_7510,N_6183,N_6141);
nand U7511 (N_7511,N_6475,N_6911);
nand U7512 (N_7512,N_6718,N_6362);
or U7513 (N_7513,N_6671,N_6057);
and U7514 (N_7514,N_6715,N_6994);
and U7515 (N_7515,N_6139,N_6914);
and U7516 (N_7516,N_6786,N_6308);
and U7517 (N_7517,N_6008,N_6389);
and U7518 (N_7518,N_6400,N_6244);
and U7519 (N_7519,N_6362,N_6903);
xor U7520 (N_7520,N_6756,N_6456);
and U7521 (N_7521,N_6180,N_6933);
and U7522 (N_7522,N_6228,N_6519);
nor U7523 (N_7523,N_6076,N_6300);
and U7524 (N_7524,N_6920,N_6936);
nor U7525 (N_7525,N_6759,N_6489);
or U7526 (N_7526,N_6336,N_6315);
xnor U7527 (N_7527,N_6821,N_6807);
or U7528 (N_7528,N_6788,N_6014);
and U7529 (N_7529,N_6571,N_6893);
nand U7530 (N_7530,N_6906,N_6483);
nand U7531 (N_7531,N_6301,N_6744);
nor U7532 (N_7532,N_6791,N_6046);
or U7533 (N_7533,N_6112,N_6407);
nor U7534 (N_7534,N_6903,N_6200);
xnor U7535 (N_7535,N_6530,N_6112);
nor U7536 (N_7536,N_6857,N_6913);
and U7537 (N_7537,N_6494,N_6400);
nand U7538 (N_7538,N_6793,N_6365);
nor U7539 (N_7539,N_6068,N_6042);
nor U7540 (N_7540,N_6329,N_6583);
or U7541 (N_7541,N_6881,N_6799);
nor U7542 (N_7542,N_6056,N_6101);
or U7543 (N_7543,N_6531,N_6556);
and U7544 (N_7544,N_6997,N_6871);
nor U7545 (N_7545,N_6760,N_6384);
nor U7546 (N_7546,N_6265,N_6138);
nand U7547 (N_7547,N_6516,N_6973);
nand U7548 (N_7548,N_6264,N_6017);
and U7549 (N_7549,N_6467,N_6185);
nand U7550 (N_7550,N_6935,N_6652);
nor U7551 (N_7551,N_6990,N_6652);
and U7552 (N_7552,N_6751,N_6096);
and U7553 (N_7553,N_6071,N_6881);
nor U7554 (N_7554,N_6157,N_6845);
or U7555 (N_7555,N_6044,N_6108);
or U7556 (N_7556,N_6874,N_6889);
and U7557 (N_7557,N_6548,N_6765);
or U7558 (N_7558,N_6444,N_6280);
xor U7559 (N_7559,N_6996,N_6885);
nor U7560 (N_7560,N_6155,N_6844);
or U7561 (N_7561,N_6715,N_6396);
nor U7562 (N_7562,N_6744,N_6591);
and U7563 (N_7563,N_6044,N_6133);
and U7564 (N_7564,N_6327,N_6356);
and U7565 (N_7565,N_6899,N_6055);
or U7566 (N_7566,N_6904,N_6187);
nand U7567 (N_7567,N_6340,N_6195);
or U7568 (N_7568,N_6743,N_6633);
or U7569 (N_7569,N_6233,N_6838);
nor U7570 (N_7570,N_6627,N_6076);
nand U7571 (N_7571,N_6406,N_6359);
nor U7572 (N_7572,N_6237,N_6520);
nor U7573 (N_7573,N_6834,N_6986);
nand U7574 (N_7574,N_6452,N_6171);
or U7575 (N_7575,N_6819,N_6022);
or U7576 (N_7576,N_6331,N_6884);
nand U7577 (N_7577,N_6670,N_6027);
or U7578 (N_7578,N_6108,N_6121);
or U7579 (N_7579,N_6690,N_6446);
nor U7580 (N_7580,N_6668,N_6005);
or U7581 (N_7581,N_6473,N_6499);
nand U7582 (N_7582,N_6431,N_6335);
or U7583 (N_7583,N_6856,N_6409);
or U7584 (N_7584,N_6206,N_6662);
nor U7585 (N_7585,N_6071,N_6396);
and U7586 (N_7586,N_6621,N_6179);
nor U7587 (N_7587,N_6324,N_6228);
or U7588 (N_7588,N_6472,N_6099);
nand U7589 (N_7589,N_6460,N_6572);
nand U7590 (N_7590,N_6650,N_6304);
and U7591 (N_7591,N_6467,N_6406);
or U7592 (N_7592,N_6003,N_6800);
or U7593 (N_7593,N_6821,N_6473);
or U7594 (N_7594,N_6730,N_6663);
nand U7595 (N_7595,N_6939,N_6533);
and U7596 (N_7596,N_6781,N_6970);
and U7597 (N_7597,N_6649,N_6178);
nor U7598 (N_7598,N_6057,N_6268);
nand U7599 (N_7599,N_6483,N_6708);
nor U7600 (N_7600,N_6325,N_6211);
nor U7601 (N_7601,N_6103,N_6867);
and U7602 (N_7602,N_6221,N_6850);
nor U7603 (N_7603,N_6060,N_6353);
or U7604 (N_7604,N_6441,N_6032);
or U7605 (N_7605,N_6740,N_6770);
nor U7606 (N_7606,N_6509,N_6944);
or U7607 (N_7607,N_6645,N_6332);
nor U7608 (N_7608,N_6334,N_6885);
and U7609 (N_7609,N_6676,N_6827);
nor U7610 (N_7610,N_6387,N_6435);
nor U7611 (N_7611,N_6076,N_6139);
or U7612 (N_7612,N_6410,N_6230);
or U7613 (N_7613,N_6734,N_6924);
and U7614 (N_7614,N_6494,N_6150);
nand U7615 (N_7615,N_6484,N_6619);
nor U7616 (N_7616,N_6455,N_6632);
or U7617 (N_7617,N_6330,N_6282);
nand U7618 (N_7618,N_6865,N_6614);
and U7619 (N_7619,N_6223,N_6280);
or U7620 (N_7620,N_6566,N_6710);
and U7621 (N_7621,N_6916,N_6920);
and U7622 (N_7622,N_6861,N_6503);
and U7623 (N_7623,N_6195,N_6666);
and U7624 (N_7624,N_6921,N_6889);
or U7625 (N_7625,N_6297,N_6494);
or U7626 (N_7626,N_6445,N_6714);
nand U7627 (N_7627,N_6751,N_6026);
nor U7628 (N_7628,N_6293,N_6044);
or U7629 (N_7629,N_6704,N_6577);
and U7630 (N_7630,N_6138,N_6611);
nand U7631 (N_7631,N_6992,N_6731);
or U7632 (N_7632,N_6523,N_6230);
or U7633 (N_7633,N_6003,N_6116);
or U7634 (N_7634,N_6396,N_6525);
or U7635 (N_7635,N_6434,N_6578);
nor U7636 (N_7636,N_6752,N_6141);
and U7637 (N_7637,N_6654,N_6106);
or U7638 (N_7638,N_6765,N_6135);
nor U7639 (N_7639,N_6120,N_6497);
nor U7640 (N_7640,N_6730,N_6495);
xor U7641 (N_7641,N_6506,N_6954);
and U7642 (N_7642,N_6073,N_6800);
and U7643 (N_7643,N_6544,N_6495);
and U7644 (N_7644,N_6021,N_6181);
nand U7645 (N_7645,N_6393,N_6838);
nor U7646 (N_7646,N_6348,N_6150);
or U7647 (N_7647,N_6090,N_6045);
nor U7648 (N_7648,N_6454,N_6485);
nor U7649 (N_7649,N_6140,N_6273);
or U7650 (N_7650,N_6008,N_6442);
or U7651 (N_7651,N_6172,N_6375);
nand U7652 (N_7652,N_6865,N_6228);
or U7653 (N_7653,N_6747,N_6933);
or U7654 (N_7654,N_6798,N_6145);
or U7655 (N_7655,N_6343,N_6276);
and U7656 (N_7656,N_6574,N_6549);
nor U7657 (N_7657,N_6950,N_6969);
nor U7658 (N_7658,N_6282,N_6892);
and U7659 (N_7659,N_6503,N_6207);
and U7660 (N_7660,N_6209,N_6964);
nor U7661 (N_7661,N_6129,N_6601);
or U7662 (N_7662,N_6850,N_6384);
or U7663 (N_7663,N_6724,N_6133);
nor U7664 (N_7664,N_6019,N_6043);
nand U7665 (N_7665,N_6265,N_6522);
nor U7666 (N_7666,N_6669,N_6810);
nor U7667 (N_7667,N_6414,N_6619);
nand U7668 (N_7668,N_6478,N_6089);
and U7669 (N_7669,N_6691,N_6617);
nand U7670 (N_7670,N_6623,N_6491);
nand U7671 (N_7671,N_6826,N_6866);
and U7672 (N_7672,N_6246,N_6991);
and U7673 (N_7673,N_6777,N_6954);
or U7674 (N_7674,N_6368,N_6246);
or U7675 (N_7675,N_6733,N_6738);
nor U7676 (N_7676,N_6132,N_6959);
or U7677 (N_7677,N_6997,N_6310);
nand U7678 (N_7678,N_6382,N_6038);
nand U7679 (N_7679,N_6963,N_6772);
nand U7680 (N_7680,N_6291,N_6258);
or U7681 (N_7681,N_6703,N_6463);
xor U7682 (N_7682,N_6777,N_6263);
and U7683 (N_7683,N_6614,N_6789);
or U7684 (N_7684,N_6544,N_6175);
and U7685 (N_7685,N_6855,N_6336);
nor U7686 (N_7686,N_6147,N_6437);
nor U7687 (N_7687,N_6232,N_6079);
and U7688 (N_7688,N_6408,N_6934);
nand U7689 (N_7689,N_6316,N_6783);
nor U7690 (N_7690,N_6179,N_6642);
and U7691 (N_7691,N_6362,N_6366);
nand U7692 (N_7692,N_6670,N_6558);
nand U7693 (N_7693,N_6120,N_6314);
or U7694 (N_7694,N_6045,N_6753);
nand U7695 (N_7695,N_6043,N_6434);
xnor U7696 (N_7696,N_6171,N_6172);
nand U7697 (N_7697,N_6977,N_6878);
nor U7698 (N_7698,N_6994,N_6893);
and U7699 (N_7699,N_6639,N_6274);
nor U7700 (N_7700,N_6710,N_6605);
or U7701 (N_7701,N_6745,N_6196);
nand U7702 (N_7702,N_6373,N_6234);
or U7703 (N_7703,N_6672,N_6970);
or U7704 (N_7704,N_6229,N_6003);
and U7705 (N_7705,N_6464,N_6708);
and U7706 (N_7706,N_6713,N_6782);
or U7707 (N_7707,N_6509,N_6239);
nor U7708 (N_7708,N_6001,N_6872);
and U7709 (N_7709,N_6644,N_6946);
nor U7710 (N_7710,N_6837,N_6450);
and U7711 (N_7711,N_6338,N_6671);
and U7712 (N_7712,N_6696,N_6873);
or U7713 (N_7713,N_6240,N_6635);
nor U7714 (N_7714,N_6073,N_6938);
or U7715 (N_7715,N_6251,N_6125);
and U7716 (N_7716,N_6817,N_6445);
or U7717 (N_7717,N_6900,N_6572);
nor U7718 (N_7718,N_6008,N_6487);
and U7719 (N_7719,N_6143,N_6617);
nor U7720 (N_7720,N_6525,N_6131);
nand U7721 (N_7721,N_6274,N_6938);
and U7722 (N_7722,N_6681,N_6172);
or U7723 (N_7723,N_6352,N_6011);
or U7724 (N_7724,N_6122,N_6449);
or U7725 (N_7725,N_6058,N_6369);
xor U7726 (N_7726,N_6306,N_6210);
nand U7727 (N_7727,N_6008,N_6402);
or U7728 (N_7728,N_6749,N_6739);
nor U7729 (N_7729,N_6326,N_6987);
nand U7730 (N_7730,N_6499,N_6963);
and U7731 (N_7731,N_6631,N_6650);
nor U7732 (N_7732,N_6348,N_6513);
or U7733 (N_7733,N_6171,N_6805);
or U7734 (N_7734,N_6007,N_6366);
nor U7735 (N_7735,N_6479,N_6863);
nor U7736 (N_7736,N_6360,N_6148);
or U7737 (N_7737,N_6643,N_6108);
nand U7738 (N_7738,N_6581,N_6728);
nor U7739 (N_7739,N_6303,N_6626);
nor U7740 (N_7740,N_6121,N_6787);
nor U7741 (N_7741,N_6717,N_6201);
or U7742 (N_7742,N_6169,N_6163);
nand U7743 (N_7743,N_6305,N_6192);
nor U7744 (N_7744,N_6288,N_6018);
nor U7745 (N_7745,N_6912,N_6332);
nor U7746 (N_7746,N_6964,N_6948);
nand U7747 (N_7747,N_6704,N_6283);
xnor U7748 (N_7748,N_6352,N_6250);
nand U7749 (N_7749,N_6032,N_6415);
nor U7750 (N_7750,N_6583,N_6730);
nor U7751 (N_7751,N_6613,N_6506);
nor U7752 (N_7752,N_6139,N_6755);
and U7753 (N_7753,N_6841,N_6377);
nor U7754 (N_7754,N_6167,N_6291);
or U7755 (N_7755,N_6551,N_6077);
nor U7756 (N_7756,N_6764,N_6328);
nand U7757 (N_7757,N_6816,N_6593);
nor U7758 (N_7758,N_6090,N_6564);
and U7759 (N_7759,N_6875,N_6427);
and U7760 (N_7760,N_6208,N_6201);
and U7761 (N_7761,N_6572,N_6186);
nand U7762 (N_7762,N_6744,N_6407);
nor U7763 (N_7763,N_6922,N_6689);
nand U7764 (N_7764,N_6216,N_6609);
and U7765 (N_7765,N_6108,N_6861);
and U7766 (N_7766,N_6858,N_6656);
or U7767 (N_7767,N_6626,N_6262);
and U7768 (N_7768,N_6198,N_6021);
and U7769 (N_7769,N_6697,N_6807);
nor U7770 (N_7770,N_6030,N_6434);
and U7771 (N_7771,N_6530,N_6015);
xor U7772 (N_7772,N_6329,N_6767);
or U7773 (N_7773,N_6224,N_6464);
or U7774 (N_7774,N_6360,N_6128);
nor U7775 (N_7775,N_6497,N_6486);
nand U7776 (N_7776,N_6659,N_6221);
nand U7777 (N_7777,N_6480,N_6428);
nand U7778 (N_7778,N_6261,N_6587);
nor U7779 (N_7779,N_6488,N_6363);
nand U7780 (N_7780,N_6286,N_6729);
and U7781 (N_7781,N_6571,N_6406);
nor U7782 (N_7782,N_6312,N_6298);
nor U7783 (N_7783,N_6958,N_6321);
nor U7784 (N_7784,N_6982,N_6583);
nor U7785 (N_7785,N_6905,N_6514);
and U7786 (N_7786,N_6405,N_6343);
nand U7787 (N_7787,N_6593,N_6654);
nor U7788 (N_7788,N_6827,N_6241);
nand U7789 (N_7789,N_6335,N_6832);
nand U7790 (N_7790,N_6232,N_6199);
nor U7791 (N_7791,N_6650,N_6011);
nor U7792 (N_7792,N_6261,N_6325);
nand U7793 (N_7793,N_6287,N_6759);
and U7794 (N_7794,N_6687,N_6645);
or U7795 (N_7795,N_6161,N_6050);
nand U7796 (N_7796,N_6838,N_6153);
and U7797 (N_7797,N_6619,N_6042);
or U7798 (N_7798,N_6733,N_6576);
nor U7799 (N_7799,N_6214,N_6407);
and U7800 (N_7800,N_6042,N_6525);
or U7801 (N_7801,N_6376,N_6118);
or U7802 (N_7802,N_6787,N_6041);
and U7803 (N_7803,N_6974,N_6390);
nor U7804 (N_7804,N_6976,N_6689);
nand U7805 (N_7805,N_6459,N_6296);
or U7806 (N_7806,N_6715,N_6286);
or U7807 (N_7807,N_6001,N_6490);
or U7808 (N_7808,N_6127,N_6182);
nand U7809 (N_7809,N_6349,N_6303);
or U7810 (N_7810,N_6056,N_6989);
and U7811 (N_7811,N_6741,N_6431);
and U7812 (N_7812,N_6872,N_6756);
or U7813 (N_7813,N_6215,N_6905);
or U7814 (N_7814,N_6449,N_6955);
and U7815 (N_7815,N_6193,N_6291);
nand U7816 (N_7816,N_6071,N_6184);
and U7817 (N_7817,N_6931,N_6916);
nor U7818 (N_7818,N_6205,N_6617);
nand U7819 (N_7819,N_6799,N_6899);
nor U7820 (N_7820,N_6002,N_6417);
nand U7821 (N_7821,N_6302,N_6660);
xnor U7822 (N_7822,N_6805,N_6277);
and U7823 (N_7823,N_6550,N_6459);
and U7824 (N_7824,N_6397,N_6316);
and U7825 (N_7825,N_6214,N_6087);
nor U7826 (N_7826,N_6932,N_6730);
and U7827 (N_7827,N_6339,N_6619);
nor U7828 (N_7828,N_6869,N_6879);
nor U7829 (N_7829,N_6169,N_6679);
and U7830 (N_7830,N_6552,N_6514);
or U7831 (N_7831,N_6822,N_6248);
nor U7832 (N_7832,N_6611,N_6604);
or U7833 (N_7833,N_6250,N_6578);
nand U7834 (N_7834,N_6351,N_6519);
nor U7835 (N_7835,N_6752,N_6719);
or U7836 (N_7836,N_6714,N_6094);
nor U7837 (N_7837,N_6367,N_6825);
or U7838 (N_7838,N_6606,N_6117);
or U7839 (N_7839,N_6431,N_6273);
or U7840 (N_7840,N_6779,N_6140);
nor U7841 (N_7841,N_6286,N_6637);
xor U7842 (N_7842,N_6405,N_6832);
nand U7843 (N_7843,N_6562,N_6167);
or U7844 (N_7844,N_6067,N_6001);
nand U7845 (N_7845,N_6767,N_6392);
or U7846 (N_7846,N_6640,N_6875);
and U7847 (N_7847,N_6491,N_6665);
nor U7848 (N_7848,N_6909,N_6800);
and U7849 (N_7849,N_6914,N_6800);
and U7850 (N_7850,N_6530,N_6912);
xnor U7851 (N_7851,N_6558,N_6772);
nor U7852 (N_7852,N_6929,N_6994);
and U7853 (N_7853,N_6092,N_6163);
and U7854 (N_7854,N_6057,N_6335);
nand U7855 (N_7855,N_6909,N_6189);
nand U7856 (N_7856,N_6631,N_6598);
and U7857 (N_7857,N_6881,N_6889);
or U7858 (N_7858,N_6674,N_6308);
nor U7859 (N_7859,N_6295,N_6704);
and U7860 (N_7860,N_6336,N_6106);
nand U7861 (N_7861,N_6497,N_6790);
nor U7862 (N_7862,N_6335,N_6412);
and U7863 (N_7863,N_6024,N_6751);
xor U7864 (N_7864,N_6344,N_6238);
and U7865 (N_7865,N_6311,N_6034);
xor U7866 (N_7866,N_6772,N_6094);
or U7867 (N_7867,N_6194,N_6181);
nor U7868 (N_7868,N_6531,N_6807);
or U7869 (N_7869,N_6017,N_6673);
and U7870 (N_7870,N_6836,N_6749);
or U7871 (N_7871,N_6506,N_6162);
nand U7872 (N_7872,N_6541,N_6286);
nand U7873 (N_7873,N_6527,N_6048);
and U7874 (N_7874,N_6252,N_6880);
and U7875 (N_7875,N_6065,N_6998);
or U7876 (N_7876,N_6297,N_6392);
or U7877 (N_7877,N_6860,N_6529);
nand U7878 (N_7878,N_6724,N_6172);
nand U7879 (N_7879,N_6638,N_6354);
nand U7880 (N_7880,N_6884,N_6752);
nand U7881 (N_7881,N_6591,N_6586);
nand U7882 (N_7882,N_6208,N_6247);
nor U7883 (N_7883,N_6242,N_6737);
or U7884 (N_7884,N_6232,N_6640);
and U7885 (N_7885,N_6827,N_6829);
and U7886 (N_7886,N_6993,N_6936);
nand U7887 (N_7887,N_6814,N_6709);
nor U7888 (N_7888,N_6379,N_6898);
nor U7889 (N_7889,N_6428,N_6288);
and U7890 (N_7890,N_6658,N_6892);
or U7891 (N_7891,N_6607,N_6771);
and U7892 (N_7892,N_6816,N_6218);
nor U7893 (N_7893,N_6346,N_6383);
nor U7894 (N_7894,N_6113,N_6944);
nor U7895 (N_7895,N_6864,N_6857);
nor U7896 (N_7896,N_6547,N_6619);
nor U7897 (N_7897,N_6816,N_6048);
and U7898 (N_7898,N_6687,N_6304);
nor U7899 (N_7899,N_6832,N_6750);
nand U7900 (N_7900,N_6907,N_6116);
nor U7901 (N_7901,N_6429,N_6210);
nand U7902 (N_7902,N_6074,N_6678);
or U7903 (N_7903,N_6501,N_6970);
nor U7904 (N_7904,N_6981,N_6056);
and U7905 (N_7905,N_6490,N_6971);
or U7906 (N_7906,N_6930,N_6835);
nor U7907 (N_7907,N_6801,N_6493);
nand U7908 (N_7908,N_6403,N_6902);
nand U7909 (N_7909,N_6439,N_6111);
and U7910 (N_7910,N_6241,N_6035);
nand U7911 (N_7911,N_6835,N_6112);
nand U7912 (N_7912,N_6579,N_6388);
nand U7913 (N_7913,N_6362,N_6948);
nor U7914 (N_7914,N_6209,N_6420);
or U7915 (N_7915,N_6758,N_6565);
nand U7916 (N_7916,N_6131,N_6096);
nor U7917 (N_7917,N_6862,N_6839);
nor U7918 (N_7918,N_6933,N_6639);
and U7919 (N_7919,N_6563,N_6554);
and U7920 (N_7920,N_6541,N_6333);
nand U7921 (N_7921,N_6850,N_6130);
nor U7922 (N_7922,N_6530,N_6633);
nand U7923 (N_7923,N_6603,N_6293);
and U7924 (N_7924,N_6061,N_6766);
and U7925 (N_7925,N_6408,N_6364);
and U7926 (N_7926,N_6785,N_6675);
and U7927 (N_7927,N_6283,N_6337);
xor U7928 (N_7928,N_6961,N_6868);
or U7929 (N_7929,N_6937,N_6133);
nand U7930 (N_7930,N_6593,N_6805);
nor U7931 (N_7931,N_6847,N_6984);
and U7932 (N_7932,N_6012,N_6385);
nand U7933 (N_7933,N_6858,N_6741);
nor U7934 (N_7934,N_6064,N_6567);
or U7935 (N_7935,N_6047,N_6319);
and U7936 (N_7936,N_6320,N_6364);
and U7937 (N_7937,N_6310,N_6895);
nand U7938 (N_7938,N_6312,N_6762);
or U7939 (N_7939,N_6343,N_6132);
nand U7940 (N_7940,N_6261,N_6125);
or U7941 (N_7941,N_6101,N_6815);
or U7942 (N_7942,N_6926,N_6607);
nor U7943 (N_7943,N_6080,N_6769);
nor U7944 (N_7944,N_6426,N_6211);
nor U7945 (N_7945,N_6225,N_6820);
nand U7946 (N_7946,N_6751,N_6682);
nor U7947 (N_7947,N_6459,N_6718);
and U7948 (N_7948,N_6934,N_6137);
or U7949 (N_7949,N_6915,N_6811);
or U7950 (N_7950,N_6391,N_6329);
nor U7951 (N_7951,N_6991,N_6467);
and U7952 (N_7952,N_6541,N_6947);
nand U7953 (N_7953,N_6207,N_6196);
nand U7954 (N_7954,N_6526,N_6508);
and U7955 (N_7955,N_6098,N_6282);
nand U7956 (N_7956,N_6269,N_6838);
xnor U7957 (N_7957,N_6602,N_6314);
nor U7958 (N_7958,N_6534,N_6211);
nand U7959 (N_7959,N_6651,N_6776);
nor U7960 (N_7960,N_6820,N_6571);
nor U7961 (N_7961,N_6111,N_6712);
xor U7962 (N_7962,N_6024,N_6489);
and U7963 (N_7963,N_6243,N_6642);
or U7964 (N_7964,N_6423,N_6071);
nand U7965 (N_7965,N_6516,N_6459);
and U7966 (N_7966,N_6345,N_6149);
and U7967 (N_7967,N_6105,N_6352);
or U7968 (N_7968,N_6697,N_6468);
nand U7969 (N_7969,N_6380,N_6071);
or U7970 (N_7970,N_6843,N_6493);
or U7971 (N_7971,N_6623,N_6916);
nand U7972 (N_7972,N_6366,N_6385);
and U7973 (N_7973,N_6714,N_6893);
nand U7974 (N_7974,N_6663,N_6676);
xnor U7975 (N_7975,N_6177,N_6447);
nor U7976 (N_7976,N_6254,N_6302);
nand U7977 (N_7977,N_6382,N_6337);
nor U7978 (N_7978,N_6216,N_6655);
nor U7979 (N_7979,N_6805,N_6926);
or U7980 (N_7980,N_6525,N_6931);
nor U7981 (N_7981,N_6031,N_6695);
or U7982 (N_7982,N_6413,N_6010);
nor U7983 (N_7983,N_6207,N_6040);
and U7984 (N_7984,N_6487,N_6196);
and U7985 (N_7985,N_6741,N_6146);
and U7986 (N_7986,N_6604,N_6660);
or U7987 (N_7987,N_6503,N_6738);
and U7988 (N_7988,N_6203,N_6145);
and U7989 (N_7989,N_6221,N_6127);
or U7990 (N_7990,N_6939,N_6620);
or U7991 (N_7991,N_6015,N_6354);
or U7992 (N_7992,N_6744,N_6057);
nor U7993 (N_7993,N_6815,N_6885);
nor U7994 (N_7994,N_6062,N_6018);
nor U7995 (N_7995,N_6061,N_6011);
or U7996 (N_7996,N_6440,N_6751);
nor U7997 (N_7997,N_6321,N_6892);
nor U7998 (N_7998,N_6888,N_6200);
or U7999 (N_7999,N_6029,N_6248);
nor U8000 (N_8000,N_7168,N_7174);
or U8001 (N_8001,N_7010,N_7428);
or U8002 (N_8002,N_7240,N_7455);
and U8003 (N_8003,N_7535,N_7638);
nand U8004 (N_8004,N_7761,N_7381);
and U8005 (N_8005,N_7923,N_7832);
or U8006 (N_8006,N_7324,N_7201);
nand U8007 (N_8007,N_7263,N_7417);
and U8008 (N_8008,N_7975,N_7176);
nand U8009 (N_8009,N_7237,N_7561);
nor U8010 (N_8010,N_7164,N_7096);
nor U8011 (N_8011,N_7342,N_7668);
and U8012 (N_8012,N_7114,N_7976);
or U8013 (N_8013,N_7597,N_7525);
nor U8014 (N_8014,N_7770,N_7574);
or U8015 (N_8015,N_7282,N_7393);
or U8016 (N_8016,N_7407,N_7548);
xor U8017 (N_8017,N_7704,N_7048);
nor U8018 (N_8018,N_7618,N_7585);
nor U8019 (N_8019,N_7427,N_7065);
and U8020 (N_8020,N_7945,N_7312);
or U8021 (N_8021,N_7150,N_7703);
nor U8022 (N_8022,N_7152,N_7082);
nand U8023 (N_8023,N_7510,N_7496);
nor U8024 (N_8024,N_7038,N_7803);
and U8025 (N_8025,N_7280,N_7452);
nor U8026 (N_8026,N_7921,N_7582);
and U8027 (N_8027,N_7523,N_7659);
and U8028 (N_8028,N_7666,N_7292);
nor U8029 (N_8029,N_7589,N_7112);
and U8030 (N_8030,N_7678,N_7692);
nor U8031 (N_8031,N_7441,N_7362);
or U8032 (N_8032,N_7738,N_7556);
nand U8033 (N_8033,N_7911,N_7485);
xnor U8034 (N_8034,N_7872,N_7575);
or U8035 (N_8035,N_7186,N_7071);
and U8036 (N_8036,N_7093,N_7996);
or U8037 (N_8037,N_7415,N_7330);
nand U8038 (N_8038,N_7265,N_7951);
nor U8039 (N_8039,N_7504,N_7273);
or U8040 (N_8040,N_7306,N_7771);
nor U8041 (N_8041,N_7453,N_7365);
and U8042 (N_8042,N_7805,N_7867);
and U8043 (N_8043,N_7420,N_7933);
nand U8044 (N_8044,N_7645,N_7020);
and U8045 (N_8045,N_7220,N_7818);
or U8046 (N_8046,N_7607,N_7717);
nor U8047 (N_8047,N_7664,N_7379);
and U8048 (N_8048,N_7806,N_7327);
nand U8049 (N_8049,N_7260,N_7444);
nand U8050 (N_8050,N_7231,N_7235);
nand U8051 (N_8051,N_7521,N_7336);
and U8052 (N_8052,N_7744,N_7920);
nor U8053 (N_8053,N_7963,N_7013);
nor U8054 (N_8054,N_7889,N_7087);
or U8055 (N_8055,N_7021,N_7387);
nor U8056 (N_8056,N_7541,N_7028);
nand U8057 (N_8057,N_7464,N_7497);
or U8058 (N_8058,N_7786,N_7003);
nand U8059 (N_8059,N_7739,N_7917);
or U8060 (N_8060,N_7191,N_7898);
nor U8061 (N_8061,N_7211,N_7881);
xor U8062 (N_8062,N_7080,N_7034);
or U8063 (N_8063,N_7622,N_7536);
nand U8064 (N_8064,N_7859,N_7103);
or U8065 (N_8065,N_7627,N_7180);
and U8066 (N_8066,N_7479,N_7059);
nor U8067 (N_8067,N_7251,N_7555);
or U8068 (N_8068,N_7126,N_7932);
nand U8069 (N_8069,N_7751,N_7367);
or U8070 (N_8070,N_7915,N_7785);
nand U8071 (N_8071,N_7446,N_7939);
or U8072 (N_8072,N_7526,N_7499);
or U8073 (N_8073,N_7721,N_7577);
or U8074 (N_8074,N_7671,N_7188);
xnor U8075 (N_8075,N_7078,N_7460);
nand U8076 (N_8076,N_7935,N_7552);
nand U8077 (N_8077,N_7062,N_7027);
xnor U8078 (N_8078,N_7605,N_7790);
and U8079 (N_8079,N_7438,N_7686);
nand U8080 (N_8080,N_7902,N_7547);
nand U8081 (N_8081,N_7084,N_7736);
nand U8082 (N_8082,N_7008,N_7965);
nand U8083 (N_8083,N_7085,N_7846);
or U8084 (N_8084,N_7383,N_7352);
and U8085 (N_8085,N_7852,N_7332);
or U8086 (N_8086,N_7505,N_7366);
and U8087 (N_8087,N_7328,N_7716);
nand U8088 (N_8088,N_7373,N_7562);
nor U8089 (N_8089,N_7097,N_7899);
and U8090 (N_8090,N_7787,N_7949);
nand U8091 (N_8091,N_7701,N_7817);
or U8092 (N_8092,N_7626,N_7691);
xor U8093 (N_8093,N_7601,N_7323);
nor U8094 (N_8094,N_7494,N_7754);
nor U8095 (N_8095,N_7539,N_7912);
nand U8096 (N_8096,N_7603,N_7179);
or U8097 (N_8097,N_7349,N_7000);
and U8098 (N_8098,N_7128,N_7928);
nor U8099 (N_8099,N_7882,N_7683);
nand U8100 (N_8100,N_7811,N_7989);
nor U8101 (N_8101,N_7388,N_7372);
and U8102 (N_8102,N_7752,N_7623);
and U8103 (N_8103,N_7143,N_7064);
and U8104 (N_8104,N_7224,N_7631);
and U8105 (N_8105,N_7586,N_7782);
and U8106 (N_8106,N_7836,N_7741);
nor U8107 (N_8107,N_7293,N_7764);
or U8108 (N_8108,N_7490,N_7987);
or U8109 (N_8109,N_7432,N_7285);
nand U8110 (N_8110,N_7212,N_7540);
nor U8111 (N_8111,N_7252,N_7133);
and U8112 (N_8112,N_7045,N_7542);
or U8113 (N_8113,N_7317,N_7392);
nand U8114 (N_8114,N_7066,N_7072);
or U8115 (N_8115,N_7054,N_7750);
nor U8116 (N_8116,N_7959,N_7967);
or U8117 (N_8117,N_7147,N_7728);
or U8118 (N_8118,N_7070,N_7962);
or U8119 (N_8119,N_7157,N_7579);
nand U8120 (N_8120,N_7647,N_7216);
or U8121 (N_8121,N_7635,N_7927);
and U8122 (N_8122,N_7783,N_7758);
nor U8123 (N_8123,N_7981,N_7644);
nor U8124 (N_8124,N_7808,N_7980);
or U8125 (N_8125,N_7069,N_7047);
or U8126 (N_8126,N_7591,N_7827);
nand U8127 (N_8127,N_7459,N_7232);
or U8128 (N_8128,N_7410,N_7759);
nand U8129 (N_8129,N_7290,N_7534);
nand U8130 (N_8130,N_7409,N_7506);
nand U8131 (N_8131,N_7462,N_7977);
nor U8132 (N_8132,N_7086,N_7897);
and U8133 (N_8133,N_7310,N_7138);
nand U8134 (N_8134,N_7606,N_7361);
nor U8135 (N_8135,N_7974,N_7705);
nor U8136 (N_8136,N_7257,N_7258);
and U8137 (N_8137,N_7612,N_7926);
xnor U8138 (N_8138,N_7681,N_7311);
nand U8139 (N_8139,N_7480,N_7887);
nor U8140 (N_8140,N_7694,N_7457);
nand U8141 (N_8141,N_7522,N_7725);
or U8142 (N_8142,N_7798,N_7091);
and U8143 (N_8143,N_7884,N_7160);
nand U8144 (N_8144,N_7471,N_7304);
nand U8145 (N_8145,N_7492,N_7356);
or U8146 (N_8146,N_7210,N_7637);
and U8147 (N_8147,N_7394,N_7531);
or U8148 (N_8148,N_7727,N_7609);
nor U8149 (N_8149,N_7360,N_7203);
or U8150 (N_8150,N_7537,N_7847);
nor U8151 (N_8151,N_7776,N_7733);
and U8152 (N_8152,N_7735,N_7227);
and U8153 (N_8153,N_7804,N_7826);
nand U8154 (N_8154,N_7063,N_7919);
nand U8155 (N_8155,N_7335,N_7320);
and U8156 (N_8156,N_7760,N_7192);
nand U8157 (N_8157,N_7406,N_7560);
nand U8158 (N_8158,N_7600,N_7171);
nor U8159 (N_8159,N_7057,N_7667);
nor U8160 (N_8160,N_7954,N_7971);
and U8161 (N_8161,N_7610,N_7014);
or U8162 (N_8162,N_7763,N_7820);
nor U8163 (N_8163,N_7824,N_7223);
and U8164 (N_8164,N_7132,N_7665);
nand U8165 (N_8165,N_7937,N_7891);
nor U8166 (N_8166,N_7994,N_7982);
and U8167 (N_8167,N_7658,N_7706);
or U8168 (N_8168,N_7075,N_7398);
and U8169 (N_8169,N_7343,N_7295);
nor U8170 (N_8170,N_7866,N_7219);
nor U8171 (N_8171,N_7158,N_7823);
and U8172 (N_8172,N_7868,N_7777);
and U8173 (N_8173,N_7153,N_7834);
or U8174 (N_8174,N_7642,N_7938);
or U8175 (N_8175,N_7390,N_7837);
and U8176 (N_8176,N_7643,N_7943);
nor U8177 (N_8177,N_7207,N_7594);
nand U8178 (N_8178,N_7794,N_7397);
or U8179 (N_8179,N_7012,N_7255);
and U8180 (N_8180,N_7876,N_7419);
nor U8181 (N_8181,N_7857,N_7156);
nor U8182 (N_8182,N_7461,N_7493);
nand U8183 (N_8183,N_7083,N_7656);
nand U8184 (N_8184,N_7380,N_7913);
or U8185 (N_8185,N_7119,N_7142);
and U8186 (N_8186,N_7375,N_7289);
or U8187 (N_8187,N_7007,N_7468);
nand U8188 (N_8188,N_7433,N_7151);
nand U8189 (N_8189,N_7925,N_7067);
nor U8190 (N_8190,N_7746,N_7473);
and U8191 (N_8191,N_7726,N_7743);
nand U8192 (N_8192,N_7508,N_7140);
xor U8193 (N_8193,N_7630,N_7968);
nand U8194 (N_8194,N_7720,N_7831);
nor U8195 (N_8195,N_7756,N_7329);
nor U8196 (N_8196,N_7570,N_7347);
nor U8197 (N_8197,N_7718,N_7524);
nand U8198 (N_8198,N_7970,N_7769);
and U8199 (N_8199,N_7737,N_7841);
or U8200 (N_8200,N_7044,N_7858);
and U8201 (N_8201,N_7426,N_7340);
nor U8202 (N_8202,N_7037,N_7530);
nand U8203 (N_8203,N_7074,N_7043);
and U8204 (N_8204,N_7039,N_7214);
or U8205 (N_8205,N_7113,N_7303);
xnor U8206 (N_8206,N_7567,N_7500);
or U8207 (N_8207,N_7414,N_7789);
and U8208 (N_8208,N_7979,N_7175);
nor U8209 (N_8209,N_7529,N_7946);
and U8210 (N_8210,N_7877,N_7477);
and U8211 (N_8211,N_7424,N_7543);
nor U8212 (N_8212,N_7809,N_7550);
nand U8213 (N_8213,N_7930,N_7402);
or U8214 (N_8214,N_7162,N_7275);
or U8215 (N_8215,N_7125,N_7382);
nand U8216 (N_8216,N_7272,N_7922);
xor U8217 (N_8217,N_7041,N_7100);
nand U8218 (N_8218,N_7730,N_7319);
and U8219 (N_8219,N_7217,N_7001);
nand U8220 (N_8220,N_7613,N_7641);
or U8221 (N_8221,N_7908,N_7910);
nor U8222 (N_8222,N_7370,N_7476);
or U8223 (N_8223,N_7081,N_7840);
nor U8224 (N_8224,N_7848,N_7440);
nor U8225 (N_8225,N_7105,N_7774);
nor U8226 (N_8226,N_7307,N_7115);
or U8227 (N_8227,N_7545,N_7914);
or U8228 (N_8228,N_7262,N_7895);
nor U8229 (N_8229,N_7302,N_7639);
nor U8230 (N_8230,N_7936,N_7901);
and U8231 (N_8231,N_7401,N_7269);
xnor U8232 (N_8232,N_7052,N_7715);
and U8233 (N_8233,N_7792,N_7321);
nand U8234 (N_8234,N_7843,N_7511);
or U8235 (N_8235,N_7183,N_7042);
nand U8236 (N_8236,N_7791,N_7270);
or U8237 (N_8237,N_7177,N_7907);
nand U8238 (N_8238,N_7345,N_7766);
nor U8239 (N_8239,N_7838,N_7009);
nand U8240 (N_8240,N_7624,N_7842);
or U8241 (N_8241,N_7181,N_7314);
nand U8242 (N_8242,N_7608,N_7137);
and U8243 (N_8243,N_7695,N_7924);
nand U8244 (N_8244,N_7076,N_7679);
or U8245 (N_8245,N_7865,N_7346);
and U8246 (N_8246,N_7972,N_7299);
nor U8247 (N_8247,N_7055,N_7870);
nand U8248 (N_8248,N_7144,N_7532);
nand U8249 (N_8249,N_7748,N_7713);
and U8250 (N_8250,N_7677,N_7620);
nand U8251 (N_8251,N_7032,N_7807);
and U8252 (N_8252,N_7249,N_7578);
and U8253 (N_8253,N_7145,N_7101);
nand U8254 (N_8254,N_7619,N_7948);
nor U8255 (N_8255,N_7829,N_7458);
and U8256 (N_8256,N_7376,N_7491);
nand U8257 (N_8257,N_7454,N_7830);
nand U8258 (N_8258,N_7173,N_7256);
nor U8259 (N_8259,N_7628,N_7474);
and U8260 (N_8260,N_7185,N_7833);
nand U8261 (N_8261,N_7206,N_7230);
xor U8262 (N_8262,N_7657,N_7193);
and U8263 (N_8263,N_7466,N_7095);
or U8264 (N_8264,N_7149,N_7035);
and U8265 (N_8265,N_7931,N_7029);
nor U8266 (N_8266,N_7617,N_7326);
xnor U8267 (N_8267,N_7159,N_7200);
nand U8268 (N_8268,N_7779,N_7309);
nand U8269 (N_8269,N_7709,N_7077);
or U8270 (N_8270,N_7333,N_7538);
nand U8271 (N_8271,N_7958,N_7519);
or U8272 (N_8272,N_7104,N_7563);
and U8273 (N_8273,N_7633,N_7773);
and U8274 (N_8274,N_7729,N_7015);
or U8275 (N_8275,N_7942,N_7405);
nand U8276 (N_8276,N_7364,N_7139);
and U8277 (N_8277,N_7278,N_7799);
nor U8278 (N_8278,N_7892,N_7950);
nand U8279 (N_8279,N_7576,N_7780);
nand U8280 (N_8280,N_7880,N_7018);
nor U8281 (N_8281,N_7845,N_7022);
or U8282 (N_8282,N_7225,N_7463);
and U8283 (N_8283,N_7221,N_7855);
nand U8284 (N_8284,N_7983,N_7821);
nor U8285 (N_8285,N_7348,N_7384);
and U8286 (N_8286,N_7050,N_7565);
or U8287 (N_8287,N_7445,N_7587);
nor U8288 (N_8288,N_7969,N_7089);
nor U8289 (N_8289,N_7973,N_7734);
and U8290 (N_8290,N_7564,N_7676);
or U8291 (N_8291,N_7353,N_7484);
or U8292 (N_8292,N_7288,N_7488);
nor U8293 (N_8293,N_7684,N_7862);
xnor U8294 (N_8294,N_7673,N_7204);
nor U8295 (N_8295,N_7056,N_7629);
or U8296 (N_8296,N_7250,N_7451);
and U8297 (N_8297,N_7616,N_7988);
nand U8298 (N_8298,N_7742,N_7111);
nor U8299 (N_8299,N_7590,N_7351);
nor U8300 (N_8300,N_7284,N_7634);
and U8301 (N_8301,N_7513,N_7190);
and U8302 (N_8302,N_7481,N_7599);
or U8303 (N_8303,N_7130,N_7672);
nor U8304 (N_8304,N_7124,N_7423);
nor U8305 (N_8305,N_7819,N_7412);
nand U8306 (N_8306,N_7966,N_7236);
or U8307 (N_8307,N_7244,N_7984);
or U8308 (N_8308,N_7448,N_7693);
and U8309 (N_8309,N_7017,N_7723);
or U8310 (N_8310,N_7313,N_7437);
nor U8311 (N_8311,N_7267,N_7429);
and U8312 (N_8312,N_7102,N_7205);
nand U8313 (N_8313,N_7688,N_7395);
nand U8314 (N_8314,N_7116,N_7430);
or U8315 (N_8315,N_7696,N_7184);
nor U8316 (N_8316,N_7470,N_7245);
or U8317 (N_8317,N_7719,N_7369);
or U8318 (N_8318,N_7886,N_7800);
xor U8319 (N_8319,N_7990,N_7435);
nor U8320 (N_8320,N_7136,N_7873);
nand U8321 (N_8321,N_7960,N_7992);
or U8322 (N_8322,N_7334,N_7215);
nor U8323 (N_8323,N_7797,N_7991);
nand U8324 (N_8324,N_7172,N_7649);
nand U8325 (N_8325,N_7894,N_7088);
nand U8326 (N_8326,N_7812,N_7690);
and U8327 (N_8327,N_7952,N_7229);
nand U8328 (N_8328,N_7110,N_7934);
nor U8329 (N_8329,N_7604,N_7653);
nand U8330 (N_8330,N_7486,N_7197);
or U8331 (N_8331,N_7456,N_7167);
xnor U8332 (N_8332,N_7724,N_7903);
nand U8333 (N_8333,N_7815,N_7469);
or U8334 (N_8334,N_7465,N_7707);
or U8335 (N_8335,N_7993,N_7222);
nand U8336 (N_8336,N_7700,N_7109);
or U8337 (N_8337,N_7788,N_7861);
and U8338 (N_8338,N_7941,N_7520);
nand U8339 (N_8339,N_7650,N_7025);
nor U8340 (N_8340,N_7450,N_7431);
or U8341 (N_8341,N_7006,N_7940);
nand U8342 (N_8342,N_7853,N_7860);
nor U8343 (N_8343,N_7475,N_7554);
or U8344 (N_8344,N_7999,N_7711);
and U8345 (N_8345,N_7553,N_7300);
nor U8346 (N_8346,N_7305,N_7259);
or U8347 (N_8347,N_7793,N_7745);
nand U8348 (N_8348,N_7411,N_7166);
nor U8349 (N_8349,N_7418,N_7287);
nand U8350 (N_8350,N_7439,N_7238);
nor U8351 (N_8351,N_7512,N_7024);
and U8352 (N_8352,N_7325,N_7614);
or U8353 (N_8353,N_7318,N_7663);
or U8354 (N_8354,N_7883,N_7233);
nor U8355 (N_8355,N_7828,N_7680);
or U8356 (N_8356,N_7344,N_7698);
or U8357 (N_8357,N_7875,N_7801);
nand U8358 (N_8358,N_7098,N_7169);
and U8359 (N_8359,N_7122,N_7094);
nand U8360 (N_8360,N_7957,N_7961);
nor U8361 (N_8361,N_7655,N_7885);
nand U8362 (N_8362,N_7516,N_7294);
and U8363 (N_8363,N_7955,N_7675);
nand U8364 (N_8364,N_7596,N_7117);
nand U8365 (N_8365,N_7482,N_7929);
or U8366 (N_8366,N_7503,N_7363);
or U8367 (N_8367,N_7757,N_7593);
and U8368 (N_8368,N_7092,N_7854);
nor U8369 (N_8369,N_7507,N_7781);
and U8370 (N_8370,N_7755,N_7198);
and U8371 (N_8371,N_7864,N_7031);
or U8372 (N_8372,N_7813,N_7583);
nand U8373 (N_8373,N_7953,N_7163);
nor U8374 (N_8374,N_7850,N_7396);
nor U8375 (N_8375,N_7796,N_7909);
nand U8376 (N_8376,N_7544,N_7732);
nand U8377 (N_8377,N_7918,N_7712);
nand U8378 (N_8378,N_7165,N_7515);
nor U8379 (N_8379,N_7368,N_7443);
and U8380 (N_8380,N_7199,N_7403);
and U8381 (N_8381,N_7566,N_7154);
nand U8382 (N_8382,N_7572,N_7291);
and U8383 (N_8383,N_7208,N_7023);
nor U8384 (N_8384,N_7339,N_7660);
nand U8385 (N_8385,N_7266,N_7749);
nor U8386 (N_8386,N_7767,N_7986);
nand U8387 (N_8387,N_7890,N_7598);
or U8388 (N_8388,N_7584,N_7355);
nor U8389 (N_8389,N_7371,N_7646);
nor U8390 (N_8390,N_7322,N_7196);
or U8391 (N_8391,N_7416,N_7514);
nand U8392 (N_8392,N_7073,N_7674);
or U8393 (N_8393,N_7337,N_7839);
nand U8394 (N_8394,N_7995,N_7436);
and U8395 (N_8395,N_7549,N_7241);
or U8396 (N_8396,N_7871,N_7533);
nor U8397 (N_8397,N_7408,N_7682);
and U8398 (N_8398,N_7625,N_7107);
nor U8399 (N_8399,N_7271,N_7498);
nand U8400 (N_8400,N_7517,N_7651);
or U8401 (N_8401,N_7816,N_7648);
and U8402 (N_8402,N_7518,N_7869);
and U8403 (N_8403,N_7026,N_7315);
and U8404 (N_8404,N_7226,N_7276);
nand U8405 (N_8405,N_7004,N_7264);
or U8406 (N_8406,N_7784,N_7106);
or U8407 (N_8407,N_7472,N_7243);
and U8408 (N_8408,N_7279,N_7856);
nand U8409 (N_8409,N_7509,N_7722);
and U8410 (N_8410,N_7033,N_7247);
or U8411 (N_8411,N_7557,N_7049);
or U8412 (N_8412,N_7246,N_7385);
nor U8413 (N_8413,N_7146,N_7254);
or U8414 (N_8414,N_7558,N_7134);
or U8415 (N_8415,N_7099,N_7581);
or U8416 (N_8416,N_7277,N_7449);
nor U8417 (N_8417,N_7195,N_7316);
nand U8418 (N_8418,N_7580,N_7611);
and U8419 (N_8419,N_7374,N_7068);
nand U8420 (N_8420,N_7708,N_7689);
nand U8421 (N_8421,N_7849,N_7768);
nand U8422 (N_8422,N_7778,N_7141);
and U8423 (N_8423,N_7242,N_7358);
xnor U8424 (N_8424,N_7825,N_7810);
nand U8425 (N_8425,N_7592,N_7389);
and U8426 (N_8426,N_7005,N_7011);
nor U8427 (N_8427,N_7019,N_7404);
nand U8428 (N_8428,N_7661,N_7239);
or U8429 (N_8429,N_7030,N_7985);
nand U8430 (N_8430,N_7187,N_7501);
and U8431 (N_8431,N_7123,N_7747);
nand U8432 (N_8432,N_7685,N_7051);
or U8433 (N_8433,N_7844,N_7573);
or U8434 (N_8434,N_7568,N_7447);
or U8435 (N_8435,N_7234,N_7377);
nor U8436 (N_8436,N_7127,N_7061);
or U8437 (N_8437,N_7878,N_7527);
nor U8438 (N_8438,N_7546,N_7662);
nor U8439 (N_8439,N_7253,N_7189);
nand U8440 (N_8440,N_7400,N_7331);
xnor U8441 (N_8441,N_7148,N_7298);
nand U8442 (N_8442,N_7079,N_7060);
or U8443 (N_8443,N_7155,N_7194);
nor U8444 (N_8444,N_7286,N_7851);
nor U8445 (N_8445,N_7697,N_7670);
and U8446 (N_8446,N_7893,N_7731);
or U8447 (N_8447,N_7559,N_7178);
and U8448 (N_8448,N_7202,N_7467);
nor U8449 (N_8449,N_7964,N_7425);
and U8450 (N_8450,N_7274,N_7386);
nor U8451 (N_8451,N_7775,N_7998);
nor U8452 (N_8452,N_7121,N_7636);
nand U8453 (N_8453,N_7874,N_7338);
nand U8454 (N_8454,N_7978,N_7301);
and U8455 (N_8455,N_7218,N_7569);
nand U8456 (N_8456,N_7359,N_7652);
and U8457 (N_8457,N_7997,N_7740);
nor U8458 (N_8458,N_7905,N_7956);
or U8459 (N_8459,N_7090,N_7213);
and U8460 (N_8460,N_7710,N_7422);
and U8461 (N_8461,N_7640,N_7487);
nor U8462 (N_8462,N_7354,N_7046);
or U8463 (N_8463,N_7297,N_7296);
or U8464 (N_8464,N_7350,N_7765);
nor U8465 (N_8465,N_7551,N_7916);
or U8466 (N_8466,N_7906,N_7129);
nand U8467 (N_8467,N_7528,N_7378);
and U8468 (N_8468,N_7131,N_7483);
and U8469 (N_8469,N_7002,N_7879);
nand U8470 (N_8470,N_7268,N_7621);
nand U8471 (N_8471,N_7161,N_7357);
nor U8472 (N_8472,N_7900,N_7413);
nand U8473 (N_8473,N_7714,N_7228);
nand U8474 (N_8474,N_7261,N_7863);
nand U8475 (N_8475,N_7135,N_7036);
nor U8476 (N_8476,N_7795,N_7421);
and U8477 (N_8477,N_7308,N_7814);
nor U8478 (N_8478,N_7595,N_7904);
or U8479 (N_8479,N_7108,N_7442);
nand U8480 (N_8480,N_7753,N_7654);
nand U8481 (N_8481,N_7615,N_7478);
and U8482 (N_8482,N_7762,N_7120);
nor U8483 (N_8483,N_7699,N_7209);
nor U8484 (N_8484,N_7669,N_7053);
nand U8485 (N_8485,N_7896,N_7632);
or U8486 (N_8486,N_7341,N_7944);
nor U8487 (N_8487,N_7571,N_7702);
nand U8488 (N_8488,N_7040,N_7118);
or U8489 (N_8489,N_7602,N_7772);
nand U8490 (N_8490,N_7399,N_7888);
or U8491 (N_8491,N_7502,N_7248);
or U8492 (N_8492,N_7802,N_7588);
or U8493 (N_8493,N_7495,N_7182);
nor U8494 (N_8494,N_7835,N_7170);
or U8495 (N_8495,N_7016,N_7822);
nor U8496 (N_8496,N_7391,N_7947);
nand U8497 (N_8497,N_7687,N_7283);
nand U8498 (N_8498,N_7281,N_7489);
and U8499 (N_8499,N_7058,N_7434);
nand U8500 (N_8500,N_7969,N_7974);
and U8501 (N_8501,N_7050,N_7476);
and U8502 (N_8502,N_7121,N_7683);
nand U8503 (N_8503,N_7810,N_7323);
and U8504 (N_8504,N_7047,N_7443);
and U8505 (N_8505,N_7743,N_7723);
and U8506 (N_8506,N_7658,N_7953);
nand U8507 (N_8507,N_7569,N_7835);
or U8508 (N_8508,N_7771,N_7544);
nor U8509 (N_8509,N_7925,N_7172);
nand U8510 (N_8510,N_7666,N_7344);
nand U8511 (N_8511,N_7777,N_7001);
and U8512 (N_8512,N_7717,N_7316);
nor U8513 (N_8513,N_7929,N_7564);
or U8514 (N_8514,N_7563,N_7535);
and U8515 (N_8515,N_7091,N_7517);
nor U8516 (N_8516,N_7287,N_7253);
nor U8517 (N_8517,N_7625,N_7109);
nand U8518 (N_8518,N_7041,N_7422);
or U8519 (N_8519,N_7422,N_7186);
nand U8520 (N_8520,N_7914,N_7973);
or U8521 (N_8521,N_7898,N_7792);
xnor U8522 (N_8522,N_7881,N_7635);
or U8523 (N_8523,N_7841,N_7554);
nor U8524 (N_8524,N_7376,N_7654);
nand U8525 (N_8525,N_7832,N_7124);
nor U8526 (N_8526,N_7367,N_7459);
nor U8527 (N_8527,N_7182,N_7382);
nor U8528 (N_8528,N_7492,N_7061);
and U8529 (N_8529,N_7168,N_7785);
xor U8530 (N_8530,N_7782,N_7254);
nor U8531 (N_8531,N_7850,N_7051);
xor U8532 (N_8532,N_7798,N_7002);
or U8533 (N_8533,N_7739,N_7945);
nand U8534 (N_8534,N_7695,N_7631);
nand U8535 (N_8535,N_7502,N_7669);
or U8536 (N_8536,N_7889,N_7154);
and U8537 (N_8537,N_7445,N_7712);
nand U8538 (N_8538,N_7787,N_7150);
nand U8539 (N_8539,N_7198,N_7092);
nand U8540 (N_8540,N_7967,N_7463);
or U8541 (N_8541,N_7212,N_7484);
nor U8542 (N_8542,N_7880,N_7316);
or U8543 (N_8543,N_7452,N_7230);
nand U8544 (N_8544,N_7234,N_7549);
nand U8545 (N_8545,N_7368,N_7619);
nand U8546 (N_8546,N_7407,N_7266);
or U8547 (N_8547,N_7107,N_7615);
nor U8548 (N_8548,N_7200,N_7823);
nor U8549 (N_8549,N_7612,N_7768);
nor U8550 (N_8550,N_7204,N_7278);
nor U8551 (N_8551,N_7046,N_7964);
nand U8552 (N_8552,N_7536,N_7943);
xnor U8553 (N_8553,N_7062,N_7107);
or U8554 (N_8554,N_7487,N_7908);
nor U8555 (N_8555,N_7799,N_7989);
nand U8556 (N_8556,N_7837,N_7284);
or U8557 (N_8557,N_7756,N_7530);
nor U8558 (N_8558,N_7477,N_7736);
or U8559 (N_8559,N_7897,N_7816);
nand U8560 (N_8560,N_7753,N_7652);
or U8561 (N_8561,N_7015,N_7646);
or U8562 (N_8562,N_7902,N_7671);
nor U8563 (N_8563,N_7169,N_7064);
nor U8564 (N_8564,N_7016,N_7705);
and U8565 (N_8565,N_7939,N_7457);
nand U8566 (N_8566,N_7669,N_7660);
nand U8567 (N_8567,N_7603,N_7353);
nor U8568 (N_8568,N_7888,N_7200);
xor U8569 (N_8569,N_7592,N_7017);
nor U8570 (N_8570,N_7295,N_7589);
and U8571 (N_8571,N_7419,N_7904);
and U8572 (N_8572,N_7573,N_7371);
nand U8573 (N_8573,N_7293,N_7725);
or U8574 (N_8574,N_7217,N_7496);
nand U8575 (N_8575,N_7861,N_7254);
nand U8576 (N_8576,N_7613,N_7007);
or U8577 (N_8577,N_7794,N_7324);
nand U8578 (N_8578,N_7074,N_7989);
and U8579 (N_8579,N_7556,N_7739);
nand U8580 (N_8580,N_7613,N_7289);
and U8581 (N_8581,N_7433,N_7489);
nor U8582 (N_8582,N_7992,N_7705);
nor U8583 (N_8583,N_7847,N_7055);
nor U8584 (N_8584,N_7554,N_7601);
nor U8585 (N_8585,N_7790,N_7492);
nand U8586 (N_8586,N_7673,N_7669);
nand U8587 (N_8587,N_7485,N_7608);
nand U8588 (N_8588,N_7337,N_7626);
nand U8589 (N_8589,N_7998,N_7643);
or U8590 (N_8590,N_7043,N_7513);
nand U8591 (N_8591,N_7981,N_7247);
or U8592 (N_8592,N_7282,N_7685);
and U8593 (N_8593,N_7547,N_7546);
nand U8594 (N_8594,N_7544,N_7772);
and U8595 (N_8595,N_7190,N_7919);
nand U8596 (N_8596,N_7561,N_7734);
xnor U8597 (N_8597,N_7991,N_7964);
nor U8598 (N_8598,N_7073,N_7718);
or U8599 (N_8599,N_7874,N_7240);
nor U8600 (N_8600,N_7763,N_7054);
nor U8601 (N_8601,N_7694,N_7091);
nand U8602 (N_8602,N_7486,N_7128);
or U8603 (N_8603,N_7434,N_7843);
nor U8604 (N_8604,N_7904,N_7478);
nor U8605 (N_8605,N_7515,N_7427);
nand U8606 (N_8606,N_7038,N_7460);
and U8607 (N_8607,N_7293,N_7974);
nand U8608 (N_8608,N_7391,N_7835);
nand U8609 (N_8609,N_7503,N_7333);
and U8610 (N_8610,N_7716,N_7620);
and U8611 (N_8611,N_7209,N_7051);
or U8612 (N_8612,N_7814,N_7274);
nand U8613 (N_8613,N_7969,N_7097);
nor U8614 (N_8614,N_7016,N_7375);
nand U8615 (N_8615,N_7348,N_7017);
xor U8616 (N_8616,N_7662,N_7161);
or U8617 (N_8617,N_7992,N_7610);
xor U8618 (N_8618,N_7383,N_7105);
nor U8619 (N_8619,N_7218,N_7787);
nor U8620 (N_8620,N_7033,N_7732);
xor U8621 (N_8621,N_7500,N_7064);
nor U8622 (N_8622,N_7373,N_7447);
and U8623 (N_8623,N_7026,N_7928);
nor U8624 (N_8624,N_7652,N_7253);
nor U8625 (N_8625,N_7174,N_7684);
nand U8626 (N_8626,N_7684,N_7154);
nor U8627 (N_8627,N_7734,N_7638);
nand U8628 (N_8628,N_7033,N_7436);
nand U8629 (N_8629,N_7901,N_7507);
or U8630 (N_8630,N_7942,N_7823);
nand U8631 (N_8631,N_7780,N_7510);
nand U8632 (N_8632,N_7677,N_7597);
nand U8633 (N_8633,N_7421,N_7747);
and U8634 (N_8634,N_7387,N_7107);
and U8635 (N_8635,N_7053,N_7452);
nor U8636 (N_8636,N_7548,N_7747);
or U8637 (N_8637,N_7998,N_7407);
nor U8638 (N_8638,N_7287,N_7473);
nand U8639 (N_8639,N_7345,N_7901);
or U8640 (N_8640,N_7218,N_7636);
and U8641 (N_8641,N_7154,N_7428);
or U8642 (N_8642,N_7433,N_7545);
nor U8643 (N_8643,N_7174,N_7301);
or U8644 (N_8644,N_7070,N_7310);
or U8645 (N_8645,N_7088,N_7494);
and U8646 (N_8646,N_7557,N_7480);
and U8647 (N_8647,N_7252,N_7713);
or U8648 (N_8648,N_7193,N_7011);
nor U8649 (N_8649,N_7683,N_7198);
nand U8650 (N_8650,N_7350,N_7700);
or U8651 (N_8651,N_7763,N_7470);
nand U8652 (N_8652,N_7133,N_7009);
or U8653 (N_8653,N_7173,N_7599);
and U8654 (N_8654,N_7216,N_7214);
nor U8655 (N_8655,N_7264,N_7575);
and U8656 (N_8656,N_7897,N_7602);
and U8657 (N_8657,N_7156,N_7082);
nor U8658 (N_8658,N_7723,N_7023);
nor U8659 (N_8659,N_7990,N_7870);
xor U8660 (N_8660,N_7065,N_7324);
nor U8661 (N_8661,N_7285,N_7734);
nand U8662 (N_8662,N_7873,N_7860);
nand U8663 (N_8663,N_7560,N_7377);
and U8664 (N_8664,N_7245,N_7820);
and U8665 (N_8665,N_7510,N_7449);
or U8666 (N_8666,N_7039,N_7463);
or U8667 (N_8667,N_7711,N_7934);
nor U8668 (N_8668,N_7171,N_7379);
and U8669 (N_8669,N_7702,N_7144);
nand U8670 (N_8670,N_7078,N_7360);
nand U8671 (N_8671,N_7971,N_7443);
and U8672 (N_8672,N_7833,N_7798);
or U8673 (N_8673,N_7796,N_7339);
nor U8674 (N_8674,N_7563,N_7737);
nand U8675 (N_8675,N_7601,N_7830);
xnor U8676 (N_8676,N_7614,N_7589);
or U8677 (N_8677,N_7250,N_7722);
nor U8678 (N_8678,N_7468,N_7892);
nor U8679 (N_8679,N_7909,N_7957);
nand U8680 (N_8680,N_7845,N_7344);
and U8681 (N_8681,N_7388,N_7421);
nand U8682 (N_8682,N_7017,N_7258);
nor U8683 (N_8683,N_7436,N_7342);
or U8684 (N_8684,N_7602,N_7866);
or U8685 (N_8685,N_7843,N_7697);
and U8686 (N_8686,N_7140,N_7622);
and U8687 (N_8687,N_7651,N_7274);
and U8688 (N_8688,N_7231,N_7899);
nor U8689 (N_8689,N_7298,N_7456);
and U8690 (N_8690,N_7284,N_7304);
nand U8691 (N_8691,N_7618,N_7745);
nand U8692 (N_8692,N_7683,N_7378);
and U8693 (N_8693,N_7483,N_7336);
nand U8694 (N_8694,N_7602,N_7178);
or U8695 (N_8695,N_7595,N_7666);
nand U8696 (N_8696,N_7560,N_7767);
and U8697 (N_8697,N_7627,N_7963);
nor U8698 (N_8698,N_7697,N_7411);
nor U8699 (N_8699,N_7292,N_7803);
and U8700 (N_8700,N_7231,N_7738);
nand U8701 (N_8701,N_7141,N_7392);
nand U8702 (N_8702,N_7681,N_7048);
and U8703 (N_8703,N_7183,N_7041);
nor U8704 (N_8704,N_7478,N_7345);
nand U8705 (N_8705,N_7815,N_7148);
xnor U8706 (N_8706,N_7372,N_7554);
or U8707 (N_8707,N_7801,N_7994);
nor U8708 (N_8708,N_7448,N_7646);
nor U8709 (N_8709,N_7808,N_7128);
nand U8710 (N_8710,N_7053,N_7697);
nand U8711 (N_8711,N_7349,N_7377);
nand U8712 (N_8712,N_7498,N_7904);
nand U8713 (N_8713,N_7510,N_7227);
nand U8714 (N_8714,N_7028,N_7870);
nand U8715 (N_8715,N_7639,N_7088);
nand U8716 (N_8716,N_7835,N_7123);
and U8717 (N_8717,N_7503,N_7685);
and U8718 (N_8718,N_7096,N_7823);
xnor U8719 (N_8719,N_7869,N_7061);
nor U8720 (N_8720,N_7814,N_7181);
nand U8721 (N_8721,N_7025,N_7016);
or U8722 (N_8722,N_7178,N_7617);
nor U8723 (N_8723,N_7566,N_7840);
or U8724 (N_8724,N_7567,N_7907);
nand U8725 (N_8725,N_7861,N_7944);
nor U8726 (N_8726,N_7960,N_7970);
and U8727 (N_8727,N_7872,N_7990);
or U8728 (N_8728,N_7592,N_7825);
or U8729 (N_8729,N_7311,N_7687);
and U8730 (N_8730,N_7708,N_7548);
nor U8731 (N_8731,N_7115,N_7025);
nor U8732 (N_8732,N_7766,N_7339);
nand U8733 (N_8733,N_7247,N_7969);
nor U8734 (N_8734,N_7432,N_7120);
and U8735 (N_8735,N_7000,N_7382);
and U8736 (N_8736,N_7630,N_7048);
or U8737 (N_8737,N_7191,N_7381);
nor U8738 (N_8738,N_7842,N_7398);
or U8739 (N_8739,N_7748,N_7901);
nor U8740 (N_8740,N_7581,N_7967);
nor U8741 (N_8741,N_7690,N_7495);
and U8742 (N_8742,N_7956,N_7032);
nor U8743 (N_8743,N_7701,N_7469);
and U8744 (N_8744,N_7142,N_7580);
and U8745 (N_8745,N_7553,N_7086);
and U8746 (N_8746,N_7593,N_7711);
nor U8747 (N_8747,N_7715,N_7540);
nor U8748 (N_8748,N_7316,N_7113);
or U8749 (N_8749,N_7665,N_7898);
and U8750 (N_8750,N_7996,N_7585);
and U8751 (N_8751,N_7119,N_7757);
nand U8752 (N_8752,N_7957,N_7056);
nand U8753 (N_8753,N_7214,N_7678);
and U8754 (N_8754,N_7194,N_7929);
nor U8755 (N_8755,N_7051,N_7557);
nand U8756 (N_8756,N_7772,N_7030);
and U8757 (N_8757,N_7959,N_7633);
and U8758 (N_8758,N_7227,N_7609);
nor U8759 (N_8759,N_7836,N_7053);
nand U8760 (N_8760,N_7352,N_7498);
nor U8761 (N_8761,N_7159,N_7862);
nand U8762 (N_8762,N_7819,N_7991);
nand U8763 (N_8763,N_7229,N_7456);
xor U8764 (N_8764,N_7867,N_7017);
nor U8765 (N_8765,N_7540,N_7910);
and U8766 (N_8766,N_7738,N_7331);
nor U8767 (N_8767,N_7571,N_7936);
or U8768 (N_8768,N_7785,N_7106);
and U8769 (N_8769,N_7246,N_7059);
nand U8770 (N_8770,N_7290,N_7618);
nand U8771 (N_8771,N_7748,N_7334);
and U8772 (N_8772,N_7992,N_7529);
nand U8773 (N_8773,N_7130,N_7204);
or U8774 (N_8774,N_7721,N_7500);
and U8775 (N_8775,N_7483,N_7789);
xnor U8776 (N_8776,N_7636,N_7504);
nand U8777 (N_8777,N_7706,N_7454);
and U8778 (N_8778,N_7281,N_7120);
or U8779 (N_8779,N_7373,N_7825);
and U8780 (N_8780,N_7072,N_7098);
and U8781 (N_8781,N_7285,N_7759);
and U8782 (N_8782,N_7265,N_7232);
and U8783 (N_8783,N_7531,N_7582);
or U8784 (N_8784,N_7940,N_7521);
or U8785 (N_8785,N_7729,N_7200);
nand U8786 (N_8786,N_7641,N_7563);
or U8787 (N_8787,N_7915,N_7495);
xor U8788 (N_8788,N_7169,N_7649);
and U8789 (N_8789,N_7837,N_7188);
and U8790 (N_8790,N_7051,N_7082);
nor U8791 (N_8791,N_7296,N_7762);
nand U8792 (N_8792,N_7293,N_7818);
and U8793 (N_8793,N_7250,N_7934);
nand U8794 (N_8794,N_7678,N_7632);
or U8795 (N_8795,N_7252,N_7882);
or U8796 (N_8796,N_7902,N_7338);
nand U8797 (N_8797,N_7622,N_7174);
nand U8798 (N_8798,N_7790,N_7228);
nor U8799 (N_8799,N_7368,N_7009);
nor U8800 (N_8800,N_7106,N_7924);
or U8801 (N_8801,N_7476,N_7504);
and U8802 (N_8802,N_7867,N_7197);
or U8803 (N_8803,N_7396,N_7166);
nand U8804 (N_8804,N_7219,N_7566);
nand U8805 (N_8805,N_7243,N_7656);
and U8806 (N_8806,N_7852,N_7293);
and U8807 (N_8807,N_7647,N_7721);
nor U8808 (N_8808,N_7291,N_7510);
or U8809 (N_8809,N_7279,N_7275);
and U8810 (N_8810,N_7126,N_7698);
nor U8811 (N_8811,N_7195,N_7984);
and U8812 (N_8812,N_7985,N_7306);
and U8813 (N_8813,N_7960,N_7075);
and U8814 (N_8814,N_7491,N_7395);
or U8815 (N_8815,N_7331,N_7782);
nor U8816 (N_8816,N_7582,N_7429);
and U8817 (N_8817,N_7022,N_7378);
or U8818 (N_8818,N_7955,N_7731);
nand U8819 (N_8819,N_7124,N_7394);
nand U8820 (N_8820,N_7243,N_7056);
and U8821 (N_8821,N_7358,N_7005);
or U8822 (N_8822,N_7686,N_7569);
and U8823 (N_8823,N_7717,N_7104);
nor U8824 (N_8824,N_7509,N_7476);
nor U8825 (N_8825,N_7878,N_7152);
and U8826 (N_8826,N_7477,N_7221);
and U8827 (N_8827,N_7896,N_7709);
and U8828 (N_8828,N_7500,N_7950);
nand U8829 (N_8829,N_7099,N_7031);
nor U8830 (N_8830,N_7692,N_7213);
or U8831 (N_8831,N_7550,N_7534);
nand U8832 (N_8832,N_7348,N_7462);
or U8833 (N_8833,N_7356,N_7756);
nor U8834 (N_8834,N_7098,N_7291);
nor U8835 (N_8835,N_7303,N_7326);
or U8836 (N_8836,N_7980,N_7285);
and U8837 (N_8837,N_7163,N_7354);
or U8838 (N_8838,N_7352,N_7394);
nand U8839 (N_8839,N_7750,N_7577);
or U8840 (N_8840,N_7123,N_7286);
or U8841 (N_8841,N_7123,N_7500);
or U8842 (N_8842,N_7926,N_7040);
or U8843 (N_8843,N_7515,N_7690);
and U8844 (N_8844,N_7515,N_7733);
nand U8845 (N_8845,N_7843,N_7681);
nand U8846 (N_8846,N_7241,N_7830);
and U8847 (N_8847,N_7474,N_7253);
nor U8848 (N_8848,N_7155,N_7087);
nand U8849 (N_8849,N_7528,N_7097);
nand U8850 (N_8850,N_7793,N_7257);
nand U8851 (N_8851,N_7102,N_7169);
or U8852 (N_8852,N_7389,N_7348);
nand U8853 (N_8853,N_7662,N_7286);
and U8854 (N_8854,N_7985,N_7775);
nor U8855 (N_8855,N_7302,N_7137);
nand U8856 (N_8856,N_7918,N_7145);
and U8857 (N_8857,N_7275,N_7055);
nor U8858 (N_8858,N_7026,N_7646);
nand U8859 (N_8859,N_7625,N_7831);
or U8860 (N_8860,N_7011,N_7054);
nor U8861 (N_8861,N_7308,N_7392);
nor U8862 (N_8862,N_7234,N_7655);
or U8863 (N_8863,N_7343,N_7315);
and U8864 (N_8864,N_7696,N_7318);
or U8865 (N_8865,N_7512,N_7649);
nand U8866 (N_8866,N_7009,N_7990);
nand U8867 (N_8867,N_7024,N_7285);
or U8868 (N_8868,N_7011,N_7677);
or U8869 (N_8869,N_7653,N_7294);
nand U8870 (N_8870,N_7118,N_7324);
nand U8871 (N_8871,N_7553,N_7208);
nor U8872 (N_8872,N_7737,N_7905);
nand U8873 (N_8873,N_7723,N_7718);
and U8874 (N_8874,N_7882,N_7510);
and U8875 (N_8875,N_7457,N_7131);
nor U8876 (N_8876,N_7757,N_7653);
nor U8877 (N_8877,N_7898,N_7375);
or U8878 (N_8878,N_7694,N_7258);
and U8879 (N_8879,N_7208,N_7697);
or U8880 (N_8880,N_7864,N_7539);
nor U8881 (N_8881,N_7111,N_7183);
and U8882 (N_8882,N_7435,N_7556);
nand U8883 (N_8883,N_7863,N_7955);
and U8884 (N_8884,N_7429,N_7876);
nand U8885 (N_8885,N_7783,N_7401);
and U8886 (N_8886,N_7994,N_7121);
and U8887 (N_8887,N_7289,N_7055);
or U8888 (N_8888,N_7087,N_7648);
nand U8889 (N_8889,N_7282,N_7284);
nand U8890 (N_8890,N_7181,N_7075);
or U8891 (N_8891,N_7610,N_7457);
nor U8892 (N_8892,N_7680,N_7594);
nor U8893 (N_8893,N_7877,N_7128);
or U8894 (N_8894,N_7836,N_7300);
or U8895 (N_8895,N_7932,N_7994);
nor U8896 (N_8896,N_7110,N_7719);
nor U8897 (N_8897,N_7437,N_7796);
and U8898 (N_8898,N_7152,N_7034);
nor U8899 (N_8899,N_7109,N_7287);
nand U8900 (N_8900,N_7507,N_7945);
or U8901 (N_8901,N_7626,N_7504);
nor U8902 (N_8902,N_7609,N_7620);
nand U8903 (N_8903,N_7462,N_7587);
nand U8904 (N_8904,N_7072,N_7658);
or U8905 (N_8905,N_7228,N_7598);
or U8906 (N_8906,N_7907,N_7022);
nand U8907 (N_8907,N_7403,N_7669);
and U8908 (N_8908,N_7319,N_7134);
and U8909 (N_8909,N_7166,N_7039);
or U8910 (N_8910,N_7531,N_7375);
and U8911 (N_8911,N_7008,N_7815);
nand U8912 (N_8912,N_7096,N_7378);
nor U8913 (N_8913,N_7954,N_7285);
nor U8914 (N_8914,N_7397,N_7859);
xnor U8915 (N_8915,N_7305,N_7554);
or U8916 (N_8916,N_7457,N_7254);
xor U8917 (N_8917,N_7959,N_7113);
or U8918 (N_8918,N_7709,N_7373);
nand U8919 (N_8919,N_7805,N_7956);
and U8920 (N_8920,N_7805,N_7687);
nand U8921 (N_8921,N_7197,N_7370);
or U8922 (N_8922,N_7520,N_7821);
and U8923 (N_8923,N_7329,N_7292);
nor U8924 (N_8924,N_7562,N_7595);
nor U8925 (N_8925,N_7295,N_7967);
nor U8926 (N_8926,N_7958,N_7010);
and U8927 (N_8927,N_7355,N_7052);
or U8928 (N_8928,N_7818,N_7755);
or U8929 (N_8929,N_7310,N_7386);
or U8930 (N_8930,N_7258,N_7570);
nand U8931 (N_8931,N_7702,N_7617);
or U8932 (N_8932,N_7947,N_7913);
nor U8933 (N_8933,N_7641,N_7123);
xnor U8934 (N_8934,N_7442,N_7899);
nor U8935 (N_8935,N_7429,N_7041);
or U8936 (N_8936,N_7379,N_7359);
nand U8937 (N_8937,N_7899,N_7438);
nand U8938 (N_8938,N_7079,N_7941);
or U8939 (N_8939,N_7121,N_7077);
or U8940 (N_8940,N_7952,N_7434);
or U8941 (N_8941,N_7975,N_7570);
xor U8942 (N_8942,N_7788,N_7135);
or U8943 (N_8943,N_7387,N_7856);
and U8944 (N_8944,N_7850,N_7540);
nor U8945 (N_8945,N_7041,N_7058);
and U8946 (N_8946,N_7024,N_7219);
nand U8947 (N_8947,N_7619,N_7764);
and U8948 (N_8948,N_7194,N_7786);
nand U8949 (N_8949,N_7787,N_7147);
and U8950 (N_8950,N_7135,N_7595);
and U8951 (N_8951,N_7100,N_7278);
nor U8952 (N_8952,N_7700,N_7589);
or U8953 (N_8953,N_7272,N_7142);
or U8954 (N_8954,N_7996,N_7257);
and U8955 (N_8955,N_7267,N_7828);
nor U8956 (N_8956,N_7981,N_7002);
and U8957 (N_8957,N_7396,N_7622);
nor U8958 (N_8958,N_7219,N_7015);
nor U8959 (N_8959,N_7675,N_7983);
nor U8960 (N_8960,N_7086,N_7978);
nand U8961 (N_8961,N_7021,N_7968);
nand U8962 (N_8962,N_7102,N_7149);
or U8963 (N_8963,N_7449,N_7168);
and U8964 (N_8964,N_7065,N_7030);
nand U8965 (N_8965,N_7268,N_7535);
nand U8966 (N_8966,N_7619,N_7268);
nand U8967 (N_8967,N_7394,N_7463);
or U8968 (N_8968,N_7658,N_7319);
nor U8969 (N_8969,N_7173,N_7819);
or U8970 (N_8970,N_7451,N_7513);
nor U8971 (N_8971,N_7950,N_7526);
or U8972 (N_8972,N_7290,N_7903);
nor U8973 (N_8973,N_7202,N_7680);
nand U8974 (N_8974,N_7341,N_7800);
and U8975 (N_8975,N_7483,N_7695);
and U8976 (N_8976,N_7814,N_7862);
and U8977 (N_8977,N_7051,N_7016);
nand U8978 (N_8978,N_7826,N_7676);
and U8979 (N_8979,N_7976,N_7904);
and U8980 (N_8980,N_7813,N_7965);
nor U8981 (N_8981,N_7131,N_7535);
or U8982 (N_8982,N_7211,N_7633);
nor U8983 (N_8983,N_7011,N_7262);
and U8984 (N_8984,N_7358,N_7879);
nand U8985 (N_8985,N_7237,N_7659);
or U8986 (N_8986,N_7861,N_7052);
and U8987 (N_8987,N_7192,N_7009);
nor U8988 (N_8988,N_7497,N_7329);
nor U8989 (N_8989,N_7174,N_7906);
nand U8990 (N_8990,N_7432,N_7321);
or U8991 (N_8991,N_7545,N_7685);
nor U8992 (N_8992,N_7022,N_7918);
or U8993 (N_8993,N_7064,N_7227);
nand U8994 (N_8994,N_7699,N_7730);
and U8995 (N_8995,N_7131,N_7493);
xnor U8996 (N_8996,N_7310,N_7520);
nor U8997 (N_8997,N_7770,N_7227);
nor U8998 (N_8998,N_7842,N_7486);
nor U8999 (N_8999,N_7578,N_7430);
and U9000 (N_9000,N_8245,N_8713);
nor U9001 (N_9001,N_8434,N_8096);
or U9002 (N_9002,N_8221,N_8488);
or U9003 (N_9003,N_8115,N_8742);
nand U9004 (N_9004,N_8171,N_8048);
or U9005 (N_9005,N_8251,N_8888);
nor U9006 (N_9006,N_8200,N_8003);
and U9007 (N_9007,N_8635,N_8816);
and U9008 (N_9008,N_8284,N_8930);
nand U9009 (N_9009,N_8750,N_8006);
nand U9010 (N_9010,N_8908,N_8521);
nor U9011 (N_9011,N_8013,N_8380);
nor U9012 (N_9012,N_8509,N_8177);
or U9013 (N_9013,N_8698,N_8960);
or U9014 (N_9014,N_8611,N_8173);
nand U9015 (N_9015,N_8243,N_8957);
and U9016 (N_9016,N_8996,N_8703);
or U9017 (N_9017,N_8364,N_8322);
or U9018 (N_9018,N_8358,N_8621);
and U9019 (N_9019,N_8104,N_8819);
or U9020 (N_9020,N_8292,N_8300);
and U9021 (N_9021,N_8791,N_8682);
or U9022 (N_9022,N_8023,N_8343);
nand U9023 (N_9023,N_8568,N_8369);
or U9024 (N_9024,N_8922,N_8301);
or U9025 (N_9025,N_8591,N_8867);
nor U9026 (N_9026,N_8349,N_8271);
or U9027 (N_9027,N_8734,N_8550);
nor U9028 (N_9028,N_8407,N_8099);
nand U9029 (N_9029,N_8864,N_8092);
xnor U9030 (N_9030,N_8031,N_8589);
nand U9031 (N_9031,N_8726,N_8356);
nor U9032 (N_9032,N_8983,N_8004);
nand U9033 (N_9033,N_8144,N_8677);
or U9034 (N_9034,N_8291,N_8946);
and U9035 (N_9035,N_8925,N_8389);
nor U9036 (N_9036,N_8508,N_8386);
nand U9037 (N_9037,N_8669,N_8972);
or U9038 (N_9038,N_8774,N_8307);
and U9039 (N_9039,N_8075,N_8184);
nand U9040 (N_9040,N_8757,N_8978);
and U9041 (N_9041,N_8047,N_8648);
nor U9042 (N_9042,N_8627,N_8687);
nand U9043 (N_9043,N_8760,N_8602);
xnor U9044 (N_9044,N_8168,N_8487);
nor U9045 (N_9045,N_8007,N_8994);
nand U9046 (N_9046,N_8321,N_8704);
nor U9047 (N_9047,N_8026,N_8676);
nor U9048 (N_9048,N_8832,N_8605);
nand U9049 (N_9049,N_8989,N_8257);
or U9050 (N_9050,N_8691,N_8163);
nand U9051 (N_9051,N_8986,N_8016);
nor U9052 (N_9052,N_8896,N_8014);
and U9053 (N_9053,N_8593,N_8671);
nor U9054 (N_9054,N_8727,N_8039);
nand U9055 (N_9055,N_8862,N_8125);
nand U9056 (N_9056,N_8638,N_8143);
and U9057 (N_9057,N_8641,N_8134);
and U9058 (N_9058,N_8378,N_8265);
nand U9059 (N_9059,N_8650,N_8797);
or U9060 (N_9060,N_8890,N_8062);
and U9061 (N_9061,N_8656,N_8792);
nor U9062 (N_9062,N_8324,N_8736);
and U9063 (N_9063,N_8154,N_8326);
nand U9064 (N_9064,N_8151,N_8808);
and U9065 (N_9065,N_8082,N_8640);
nand U9066 (N_9066,N_8519,N_8230);
nand U9067 (N_9067,N_8950,N_8021);
nand U9068 (N_9068,N_8795,N_8875);
or U9069 (N_9069,N_8212,N_8601);
nand U9070 (N_9070,N_8854,N_8877);
or U9071 (N_9071,N_8217,N_8309);
and U9072 (N_9072,N_8468,N_8432);
or U9073 (N_9073,N_8274,N_8109);
nand U9074 (N_9074,N_8534,N_8639);
or U9075 (N_9075,N_8775,N_8603);
nand U9076 (N_9076,N_8566,N_8279);
and U9077 (N_9077,N_8270,N_8447);
nor U9078 (N_9078,N_8554,N_8341);
or U9079 (N_9079,N_8680,N_8830);
nand U9080 (N_9080,N_8673,N_8111);
nand U9081 (N_9081,N_8945,N_8114);
nand U9082 (N_9082,N_8751,N_8348);
or U9083 (N_9083,N_8852,N_8954);
and U9084 (N_9084,N_8281,N_8740);
and U9085 (N_9085,N_8215,N_8707);
nand U9086 (N_9086,N_8132,N_8318);
nor U9087 (N_9087,N_8231,N_8112);
or U9088 (N_9088,N_8197,N_8624);
nor U9089 (N_9089,N_8761,N_8219);
nor U9090 (N_9090,N_8347,N_8926);
nor U9091 (N_9091,N_8804,N_8339);
nand U9092 (N_9092,N_8123,N_8174);
or U9093 (N_9093,N_8008,N_8465);
nor U9094 (N_9094,N_8204,N_8699);
or U9095 (N_9095,N_8503,N_8009);
nand U9096 (N_9096,N_8258,N_8452);
nand U9097 (N_9097,N_8192,N_8117);
or U9098 (N_9098,N_8497,N_8352);
xnor U9099 (N_9099,N_8442,N_8787);
nor U9100 (N_9100,N_8187,N_8728);
and U9101 (N_9101,N_8501,N_8553);
nor U9102 (N_9102,N_8098,N_8581);
nand U9103 (N_9103,N_8619,N_8579);
and U9104 (N_9104,N_8773,N_8165);
nand U9105 (N_9105,N_8222,N_8238);
nor U9106 (N_9106,N_8911,N_8990);
nand U9107 (N_9107,N_8664,N_8116);
or U9108 (N_9108,N_8555,N_8871);
nand U9109 (N_9109,N_8236,N_8695);
nor U9110 (N_9110,N_8282,N_8651);
nand U9111 (N_9111,N_8355,N_8528);
nor U9112 (N_9112,N_8334,N_8275);
or U9113 (N_9113,N_8044,N_8580);
and U9114 (N_9114,N_8499,N_8036);
or U9115 (N_9115,N_8859,N_8588);
or U9116 (N_9116,N_8128,N_8817);
and U9117 (N_9117,N_8303,N_8252);
nor U9118 (N_9118,N_8066,N_8971);
or U9119 (N_9119,N_8645,N_8456);
and U9120 (N_9120,N_8467,N_8879);
and U9121 (N_9121,N_8480,N_8183);
nor U9122 (N_9122,N_8460,N_8053);
and U9123 (N_9123,N_8675,N_8045);
or U9124 (N_9124,N_8312,N_8224);
nor U9125 (N_9125,N_8313,N_8970);
and U9126 (N_9126,N_8567,N_8402);
nand U9127 (N_9127,N_8725,N_8840);
nand U9128 (N_9128,N_8213,N_8608);
nor U9129 (N_9129,N_8845,N_8518);
or U9130 (N_9130,N_8121,N_8873);
and U9131 (N_9131,N_8074,N_8371);
or U9132 (N_9132,N_8195,N_8674);
and U9133 (N_9133,N_8937,N_8548);
and U9134 (N_9134,N_8935,N_8110);
nor U9135 (N_9135,N_8190,N_8874);
nor U9136 (N_9136,N_8866,N_8562);
or U9137 (N_9137,N_8798,N_8511);
nor U9138 (N_9138,N_8240,N_8210);
and U9139 (N_9139,N_8781,N_8712);
and U9140 (N_9140,N_8137,N_8136);
nor U9141 (N_9141,N_8785,N_8564);
or U9142 (N_9142,N_8885,N_8998);
and U9143 (N_9143,N_8860,N_8666);
or U9144 (N_9144,N_8153,N_8801);
or U9145 (N_9145,N_8827,N_8084);
or U9146 (N_9146,N_8440,N_8470);
nand U9147 (N_9147,N_8061,N_8614);
nand U9148 (N_9148,N_8055,N_8850);
or U9149 (N_9149,N_8103,N_8232);
nor U9150 (N_9150,N_8410,N_8118);
or U9151 (N_9151,N_8020,N_8451);
nand U9152 (N_9152,N_8108,N_8536);
and U9153 (N_9153,N_8182,N_8382);
nand U9154 (N_9154,N_8472,N_8263);
nor U9155 (N_9155,N_8444,N_8510);
and U9156 (N_9156,N_8283,N_8379);
nor U9157 (N_9157,N_8863,N_8482);
nand U9158 (N_9158,N_8513,N_8040);
nor U9159 (N_9159,N_8540,N_8932);
nor U9160 (N_9160,N_8626,N_8526);
and U9161 (N_9161,N_8572,N_8005);
or U9162 (N_9162,N_8720,N_8001);
or U9163 (N_9163,N_8158,N_8933);
nand U9164 (N_9164,N_8576,N_8431);
nand U9165 (N_9165,N_8962,N_8135);
and U9166 (N_9166,N_8944,N_8196);
and U9167 (N_9167,N_8476,N_8119);
and U9168 (N_9168,N_8966,N_8354);
nand U9169 (N_9169,N_8067,N_8705);
and U9170 (N_9170,N_8984,N_8749);
or U9171 (N_9171,N_8256,N_8636);
and U9172 (N_9172,N_8401,N_8069);
and U9173 (N_9173,N_8934,N_8592);
nor U9174 (N_9174,N_8900,N_8964);
xor U9175 (N_9175,N_8170,N_8500);
nand U9176 (N_9176,N_8027,N_8063);
or U9177 (N_9177,N_8314,N_8746);
or U9178 (N_9178,N_8708,N_8894);
and U9179 (N_9179,N_8072,N_8530);
or U9180 (N_9180,N_8527,N_8895);
or U9181 (N_9181,N_8419,N_8331);
and U9182 (N_9182,N_8290,N_8433);
and U9183 (N_9183,N_8756,N_8686);
nand U9184 (N_9184,N_8856,N_8679);
nand U9185 (N_9185,N_8541,N_8768);
or U9186 (N_9186,N_8024,N_8305);
xor U9187 (N_9187,N_8122,N_8623);
nand U9188 (N_9188,N_8818,N_8461);
and U9189 (N_9189,N_8872,N_8884);
and U9190 (N_9190,N_8525,N_8459);
or U9191 (N_9191,N_8507,N_8247);
nand U9192 (N_9192,N_8223,N_8942);
and U9193 (N_9193,N_8571,N_8975);
nand U9194 (N_9194,N_8824,N_8924);
nor U9195 (N_9195,N_8046,N_8308);
nor U9196 (N_9196,N_8344,N_8437);
nand U9197 (N_9197,N_8429,N_8965);
nand U9198 (N_9198,N_8094,N_8724);
or U9199 (N_9199,N_8847,N_8963);
nor U9200 (N_9200,N_8477,N_8454);
nor U9201 (N_9201,N_8237,N_8029);
or U9202 (N_9202,N_8939,N_8478);
and U9203 (N_9203,N_8051,N_8778);
nand U9204 (N_9204,N_8901,N_8865);
xor U9205 (N_9205,N_8398,N_8628);
xor U9206 (N_9206,N_8770,N_8523);
or U9207 (N_9207,N_8428,N_8587);
and U9208 (N_9208,N_8915,N_8464);
nand U9209 (N_9209,N_8595,N_8524);
and U9210 (N_9210,N_8769,N_8837);
or U9211 (N_9211,N_8552,N_8169);
nand U9212 (N_9212,N_8397,N_8194);
nor U9213 (N_9213,N_8413,N_8388);
nor U9214 (N_9214,N_8604,N_8898);
and U9215 (N_9215,N_8373,N_8362);
and U9216 (N_9216,N_8064,N_8022);
nand U9217 (N_9217,N_8383,N_8302);
nand U9218 (N_9218,N_8269,N_8150);
and U9219 (N_9219,N_8202,N_8181);
or U9220 (N_9220,N_8738,N_8372);
or U9221 (N_9221,N_8948,N_8325);
nor U9222 (N_9222,N_8779,N_8130);
and U9223 (N_9223,N_8390,N_8149);
and U9224 (N_9224,N_8980,N_8920);
and U9225 (N_9225,N_8462,N_8829);
nand U9226 (N_9226,N_8492,N_8618);
and U9227 (N_9227,N_8392,N_8156);
nor U9228 (N_9228,N_8903,N_8229);
or U9229 (N_9229,N_8748,N_8657);
nand U9230 (N_9230,N_8559,N_8883);
or U9231 (N_9231,N_8491,N_8083);
or U9232 (N_9232,N_8600,N_8216);
nor U9233 (N_9233,N_8556,N_8665);
nand U9234 (N_9234,N_8346,N_8041);
or U9235 (N_9235,N_8340,N_8709);
nor U9236 (N_9236,N_8849,N_8489);
nor U9237 (N_9237,N_8812,N_8424);
and U9238 (N_9238,N_8512,N_8805);
nor U9239 (N_9239,N_8304,N_8205);
and U9240 (N_9240,N_8266,N_8767);
nor U9241 (N_9241,N_8228,N_8642);
and U9242 (N_9242,N_8320,N_8765);
and U9243 (N_9243,N_8474,N_8949);
and U9244 (N_9244,N_8124,N_8723);
nand U9245 (N_9245,N_8690,N_8549);
nor U9246 (N_9246,N_8159,N_8080);
or U9247 (N_9247,N_8280,N_8696);
or U9248 (N_9248,N_8073,N_8869);
and U9249 (N_9249,N_8741,N_8057);
or U9250 (N_9250,N_8880,N_8764);
nand U9251 (N_9251,N_8891,N_8947);
and U9252 (N_9252,N_8446,N_8995);
nand U9253 (N_9253,N_8661,N_8493);
or U9254 (N_9254,N_8471,N_8246);
nor U9255 (N_9255,N_8090,N_8670);
and U9256 (N_9256,N_8427,N_8976);
xnor U9257 (N_9257,N_8351,N_8718);
nand U9258 (N_9258,N_8175,N_8662);
xor U9259 (N_9259,N_8913,N_8833);
xor U9260 (N_9260,N_8365,N_8453);
nand U9261 (N_9261,N_8058,N_8370);
nand U9262 (N_9262,N_8188,N_8846);
and U9263 (N_9263,N_8793,N_8086);
or U9264 (N_9264,N_8311,N_8537);
and U9265 (N_9265,N_8828,N_8059);
nor U9266 (N_9266,N_8146,N_8583);
and U9267 (N_9267,N_8927,N_8218);
nand U9268 (N_9268,N_8414,N_8233);
nor U9269 (N_9269,N_8702,N_8178);
and U9270 (N_9270,N_8733,N_8455);
nor U9271 (N_9271,N_8254,N_8490);
nor U9272 (N_9272,N_8531,N_8140);
nand U9273 (N_9273,N_8028,N_8485);
nand U9274 (N_9274,N_8813,N_8532);
and U9275 (N_9275,N_8186,N_8198);
nor U9276 (N_9276,N_8923,N_8577);
nand U9277 (N_9277,N_8988,N_8220);
and U9278 (N_9278,N_8585,N_8789);
or U9279 (N_9279,N_8054,N_8782);
and U9280 (N_9280,N_8836,N_8479);
or U9281 (N_9281,N_8701,N_8406);
or U9282 (N_9282,N_8719,N_8466);
and U9283 (N_9283,N_8113,N_8739);
and U9284 (N_9284,N_8597,N_8070);
nor U9285 (N_9285,N_8166,N_8495);
or U9286 (N_9286,N_8226,N_8209);
nor U9287 (N_9287,N_8043,N_8077);
or U9288 (N_9288,N_8260,N_8276);
nor U9289 (N_9289,N_8992,N_8071);
and U9290 (N_9290,N_8042,N_8449);
and U9291 (N_9291,N_8337,N_8502);
and U9292 (N_9292,N_8496,N_8288);
or U9293 (N_9293,N_8842,N_8936);
nor U9294 (N_9294,N_8561,N_8185);
and U9295 (N_9295,N_8049,N_8285);
nor U9296 (N_9296,N_8810,N_8943);
or U9297 (N_9297,N_8558,N_8332);
or U9298 (N_9298,N_8338,N_8542);
and U9299 (N_9299,N_8716,N_8107);
or U9300 (N_9300,N_8881,N_8617);
nand U9301 (N_9301,N_8018,N_8814);
nor U9302 (N_9302,N_8363,N_8417);
or U9303 (N_9303,N_8921,N_8399);
or U9304 (N_9304,N_8844,N_8835);
or U9305 (N_9305,N_8786,N_8010);
or U9306 (N_9306,N_8323,N_8752);
nor U9307 (N_9307,N_8203,N_8899);
nor U9308 (N_9308,N_8375,N_8823);
nor U9309 (N_9309,N_8918,N_8529);
and U9310 (N_9310,N_8999,N_8299);
or U9311 (N_9311,N_8578,N_8784);
nand U9312 (N_9312,N_8711,N_8715);
nor U9313 (N_9313,N_8929,N_8298);
or U9314 (N_9314,N_8412,N_8147);
nand U9315 (N_9315,N_8076,N_8653);
nand U9316 (N_9316,N_8145,N_8085);
xnor U9317 (N_9317,N_8295,N_8404);
and U9318 (N_9318,N_8958,N_8423);
or U9319 (N_9319,N_8977,N_8902);
and U9320 (N_9320,N_8876,N_8025);
or U9321 (N_9321,N_8357,N_8969);
nor U9322 (N_9322,N_8762,N_8056);
nand U9323 (N_9323,N_8878,N_8296);
nor U9324 (N_9324,N_8825,N_8289);
or U9325 (N_9325,N_8790,N_8486);
or U9326 (N_9326,N_8450,N_8931);
nand U9327 (N_9327,N_8234,N_8050);
xnor U9328 (N_9328,N_8294,N_8148);
nor U9329 (N_9329,N_8904,N_8857);
and U9330 (N_9330,N_8646,N_8264);
nor U9331 (N_9331,N_8387,N_8776);
nand U9332 (N_9332,N_8633,N_8938);
or U9333 (N_9333,N_8991,N_8505);
and U9334 (N_9334,N_8342,N_8967);
or U9335 (N_9335,N_8017,N_8851);
or U9336 (N_9336,N_8244,N_8102);
nor U9337 (N_9337,N_8262,N_8133);
or U9338 (N_9338,N_8415,N_8685);
nor U9339 (N_9339,N_8772,N_8754);
nor U9340 (N_9340,N_8612,N_8584);
xnor U9341 (N_9341,N_8997,N_8443);
or U9342 (N_9342,N_8138,N_8586);
nand U9343 (N_9343,N_8538,N_8652);
and U9344 (N_9344,N_8838,N_8655);
nand U9345 (N_9345,N_8737,N_8139);
and U9346 (N_9346,N_8065,N_8097);
or U9347 (N_9347,N_8317,N_8350);
and U9348 (N_9348,N_8011,N_8081);
nand U9349 (N_9349,N_8206,N_8167);
nor U9350 (N_9350,N_8853,N_8516);
nor U9351 (N_9351,N_8193,N_8408);
nor U9352 (N_9352,N_8570,N_8335);
nand U9353 (N_9353,N_8126,N_8870);
nor U9354 (N_9354,N_8806,N_8469);
or U9355 (N_9355,N_8800,N_8887);
nand U9356 (N_9356,N_8032,N_8546);
or U9357 (N_9357,N_8643,N_8882);
xor U9358 (N_9358,N_8157,N_8253);
nor U9359 (N_9359,N_8328,N_8594);
or U9360 (N_9360,N_8473,N_8214);
nor U9361 (N_9361,N_8543,N_8091);
nor U9362 (N_9362,N_8979,N_8631);
nor U9363 (N_9363,N_8393,N_8239);
or U9364 (N_9364,N_8809,N_8038);
or U9365 (N_9365,N_8384,N_8688);
or U9366 (N_9366,N_8089,N_8129);
nor U9367 (N_9367,N_8242,N_8160);
or U9368 (N_9368,N_8095,N_8327);
or U9369 (N_9369,N_8227,N_8127);
nand U9370 (N_9370,N_8141,N_8483);
and U9371 (N_9371,N_8692,N_8191);
nand U9372 (N_9372,N_8951,N_8919);
and U9373 (N_9373,N_8161,N_8912);
nor U9374 (N_9374,N_8609,N_8426);
and U9375 (N_9375,N_8396,N_8034);
or U9376 (N_9376,N_8259,N_8211);
nor U9377 (N_9377,N_8506,N_8015);
nor U9378 (N_9378,N_8649,N_8416);
nand U9379 (N_9379,N_8498,N_8573);
or U9380 (N_9380,N_8697,N_8436);
nand U9381 (N_9381,N_8208,N_8441);
nand U9382 (N_9382,N_8400,N_8164);
nor U9383 (N_9383,N_8272,N_8457);
nor U9384 (N_9384,N_8861,N_8616);
or U9385 (N_9385,N_8235,N_8316);
or U9386 (N_9386,N_8753,N_8367);
nand U9387 (N_9387,N_8799,N_8207);
nor U9388 (N_9388,N_8162,N_8336);
nand U9389 (N_9389,N_8820,N_8831);
or U9390 (N_9390,N_8729,N_8391);
and U9391 (N_9391,N_8681,N_8142);
nand U9392 (N_9392,N_8179,N_8261);
nor U9393 (N_9393,N_8421,N_8189);
nor U9394 (N_9394,N_8155,N_8255);
nor U9395 (N_9395,N_8731,N_8700);
nand U9396 (N_9396,N_8668,N_8632);
xor U9397 (N_9397,N_8458,N_8897);
nor U9398 (N_9398,N_8815,N_8771);
or U9399 (N_9399,N_8973,N_8405);
nand U9400 (N_9400,N_8788,N_8395);
or U9401 (N_9401,N_8659,N_8093);
nor U9402 (N_9402,N_8745,N_8019);
and U9403 (N_9403,N_8180,N_8598);
nor U9404 (N_9404,N_8484,N_8959);
and U9405 (N_9405,N_8359,N_8802);
or U9406 (N_9406,N_8744,N_8613);
or U9407 (N_9407,N_8078,N_8514);
or U9408 (N_9408,N_8868,N_8941);
and U9409 (N_9409,N_8940,N_8625);
or U9410 (N_9410,N_8893,N_8855);
nor U9411 (N_9411,N_8360,N_8286);
nor U9412 (N_9412,N_8435,N_8361);
nor U9413 (N_9413,N_8035,N_8647);
nor U9414 (N_9414,N_8068,N_8610);
and U9415 (N_9415,N_8105,N_8520);
nand U9416 (N_9416,N_8858,N_8374);
nor U9417 (N_9417,N_8545,N_8630);
or U9418 (N_9418,N_8310,N_8088);
nor U9419 (N_9419,N_8743,N_8678);
nor U9420 (N_9420,N_8841,N_8796);
nor U9421 (N_9421,N_8907,N_8917);
nand U9422 (N_9422,N_8599,N_8225);
nor U9423 (N_9423,N_8268,N_8582);
nand U9424 (N_9424,N_8710,N_8777);
nand U9425 (N_9425,N_8315,N_8366);
nor U9426 (N_9426,N_8293,N_8544);
nor U9427 (N_9427,N_8481,N_8394);
nor U9428 (N_9428,N_8910,N_8590);
nand U9429 (N_9429,N_8974,N_8714);
and U9430 (N_9430,N_8607,N_8445);
nand U9431 (N_9431,N_8560,N_8152);
nand U9432 (N_9432,N_8834,N_8535);
nand U9433 (N_9433,N_8886,N_8241);
nand U9434 (N_9434,N_8333,N_8377);
and U9435 (N_9435,N_8663,N_8732);
nand U9436 (N_9436,N_8418,N_8249);
and U9437 (N_9437,N_8987,N_8176);
nor U9438 (N_9438,N_8199,N_8803);
and U9439 (N_9439,N_8667,N_8329);
nand U9440 (N_9440,N_8287,N_8422);
and U9441 (N_9441,N_8672,N_8660);
or U9442 (N_9442,N_8250,N_8248);
nand U9443 (N_9443,N_8131,N_8952);
and U9444 (N_9444,N_8345,N_8905);
nor U9445 (N_9445,N_8968,N_8848);
nor U9446 (N_9446,N_8683,N_8030);
nand U9447 (N_9447,N_8615,N_8759);
or U9448 (N_9448,N_8892,N_8551);
nor U9449 (N_9449,N_8722,N_8906);
nand U9450 (N_9450,N_8330,N_8430);
and U9451 (N_9451,N_8494,N_8758);
or U9452 (N_9452,N_8569,N_8689);
and U9453 (N_9453,N_8953,N_8563);
or U9454 (N_9454,N_8634,N_8620);
and U9455 (N_9455,N_8278,N_8353);
or U9456 (N_9456,N_8574,N_8985);
nor U9457 (N_9457,N_8409,N_8012);
nand U9458 (N_9458,N_8201,N_8783);
and U9459 (N_9459,N_8956,N_8811);
nand U9460 (N_9460,N_8843,N_8439);
xor U9461 (N_9461,N_8822,N_8807);
or U9462 (N_9462,N_8981,N_8596);
or U9463 (N_9463,N_8684,N_8087);
and U9464 (N_9464,N_8504,N_8267);
and U9465 (N_9465,N_8694,N_8993);
or U9466 (N_9466,N_8794,N_8622);
nor U9467 (N_9467,N_8839,N_8575);
or U9468 (N_9468,N_8916,N_8914);
xor U9469 (N_9469,N_8730,N_8448);
or U9470 (N_9470,N_8368,N_8079);
and U9471 (N_9471,N_8106,N_8376);
and U9472 (N_9472,N_8306,N_8766);
and U9473 (N_9473,N_8780,N_8381);
nor U9474 (N_9474,N_8637,N_8000);
or U9475 (N_9475,N_8120,N_8297);
or U9476 (N_9476,N_8539,N_8475);
nor U9477 (N_9477,N_8721,N_8717);
nor U9478 (N_9478,N_8273,N_8517);
or U9479 (N_9479,N_8658,N_8002);
nand U9480 (N_9480,N_8928,N_8629);
nor U9481 (N_9481,N_8557,N_8982);
and U9482 (N_9482,N_8961,N_8955);
nand U9483 (N_9483,N_8654,N_8889);
nand U9484 (N_9484,N_8826,N_8755);
nor U9485 (N_9485,N_8606,N_8909);
or U9486 (N_9486,N_8420,N_8052);
nand U9487 (N_9487,N_8277,N_8735);
nand U9488 (N_9488,N_8385,N_8101);
or U9489 (N_9489,N_8747,N_8425);
nor U9490 (N_9490,N_8693,N_8763);
or U9491 (N_9491,N_8533,N_8172);
and U9492 (N_9492,N_8547,N_8463);
and U9493 (N_9493,N_8100,N_8060);
and U9494 (N_9494,N_8037,N_8438);
nand U9495 (N_9495,N_8515,N_8706);
and U9496 (N_9496,N_8403,N_8411);
nor U9497 (N_9497,N_8319,N_8033);
or U9498 (N_9498,N_8565,N_8644);
or U9499 (N_9499,N_8522,N_8821);
or U9500 (N_9500,N_8474,N_8237);
nor U9501 (N_9501,N_8558,N_8288);
nor U9502 (N_9502,N_8125,N_8459);
nor U9503 (N_9503,N_8808,N_8937);
and U9504 (N_9504,N_8084,N_8007);
or U9505 (N_9505,N_8813,N_8327);
or U9506 (N_9506,N_8112,N_8158);
or U9507 (N_9507,N_8706,N_8534);
or U9508 (N_9508,N_8862,N_8542);
and U9509 (N_9509,N_8726,N_8171);
nor U9510 (N_9510,N_8567,N_8347);
and U9511 (N_9511,N_8303,N_8969);
nand U9512 (N_9512,N_8422,N_8047);
or U9513 (N_9513,N_8339,N_8235);
or U9514 (N_9514,N_8452,N_8946);
nand U9515 (N_9515,N_8300,N_8704);
or U9516 (N_9516,N_8861,N_8963);
nor U9517 (N_9517,N_8165,N_8399);
nand U9518 (N_9518,N_8765,N_8821);
nor U9519 (N_9519,N_8969,N_8099);
and U9520 (N_9520,N_8736,N_8019);
nor U9521 (N_9521,N_8149,N_8338);
and U9522 (N_9522,N_8388,N_8019);
and U9523 (N_9523,N_8269,N_8997);
nand U9524 (N_9524,N_8380,N_8674);
and U9525 (N_9525,N_8611,N_8551);
nand U9526 (N_9526,N_8368,N_8461);
and U9527 (N_9527,N_8582,N_8883);
nor U9528 (N_9528,N_8579,N_8570);
nand U9529 (N_9529,N_8022,N_8622);
nor U9530 (N_9530,N_8289,N_8267);
or U9531 (N_9531,N_8958,N_8775);
nand U9532 (N_9532,N_8007,N_8204);
nand U9533 (N_9533,N_8498,N_8786);
or U9534 (N_9534,N_8319,N_8304);
nor U9535 (N_9535,N_8591,N_8602);
or U9536 (N_9536,N_8022,N_8357);
nand U9537 (N_9537,N_8065,N_8336);
and U9538 (N_9538,N_8863,N_8014);
nand U9539 (N_9539,N_8187,N_8012);
nand U9540 (N_9540,N_8546,N_8699);
or U9541 (N_9541,N_8940,N_8358);
nor U9542 (N_9542,N_8387,N_8714);
and U9543 (N_9543,N_8689,N_8624);
and U9544 (N_9544,N_8832,N_8328);
and U9545 (N_9545,N_8584,N_8452);
and U9546 (N_9546,N_8854,N_8979);
or U9547 (N_9547,N_8990,N_8732);
or U9548 (N_9548,N_8403,N_8494);
or U9549 (N_9549,N_8783,N_8080);
nor U9550 (N_9550,N_8076,N_8722);
nand U9551 (N_9551,N_8223,N_8756);
or U9552 (N_9552,N_8272,N_8685);
and U9553 (N_9553,N_8267,N_8439);
or U9554 (N_9554,N_8138,N_8038);
or U9555 (N_9555,N_8613,N_8171);
nand U9556 (N_9556,N_8026,N_8454);
nor U9557 (N_9557,N_8225,N_8436);
nand U9558 (N_9558,N_8125,N_8281);
nor U9559 (N_9559,N_8606,N_8582);
nand U9560 (N_9560,N_8071,N_8432);
xor U9561 (N_9561,N_8899,N_8270);
and U9562 (N_9562,N_8421,N_8781);
and U9563 (N_9563,N_8691,N_8226);
nand U9564 (N_9564,N_8141,N_8430);
nor U9565 (N_9565,N_8766,N_8488);
and U9566 (N_9566,N_8140,N_8069);
nand U9567 (N_9567,N_8863,N_8431);
nor U9568 (N_9568,N_8455,N_8574);
nand U9569 (N_9569,N_8840,N_8858);
nor U9570 (N_9570,N_8479,N_8808);
nor U9571 (N_9571,N_8247,N_8025);
or U9572 (N_9572,N_8409,N_8593);
nand U9573 (N_9573,N_8331,N_8082);
nand U9574 (N_9574,N_8724,N_8250);
nand U9575 (N_9575,N_8963,N_8178);
nor U9576 (N_9576,N_8184,N_8498);
nand U9577 (N_9577,N_8214,N_8893);
nand U9578 (N_9578,N_8469,N_8880);
or U9579 (N_9579,N_8596,N_8518);
and U9580 (N_9580,N_8930,N_8859);
and U9581 (N_9581,N_8151,N_8462);
nor U9582 (N_9582,N_8024,N_8504);
and U9583 (N_9583,N_8506,N_8226);
nor U9584 (N_9584,N_8076,N_8015);
or U9585 (N_9585,N_8356,N_8170);
and U9586 (N_9586,N_8905,N_8915);
nand U9587 (N_9587,N_8987,N_8565);
xnor U9588 (N_9588,N_8899,N_8051);
or U9589 (N_9589,N_8750,N_8682);
nor U9590 (N_9590,N_8372,N_8504);
nor U9591 (N_9591,N_8745,N_8282);
nor U9592 (N_9592,N_8012,N_8046);
and U9593 (N_9593,N_8078,N_8327);
nor U9594 (N_9594,N_8645,N_8879);
nand U9595 (N_9595,N_8701,N_8809);
nor U9596 (N_9596,N_8839,N_8480);
and U9597 (N_9597,N_8097,N_8693);
nand U9598 (N_9598,N_8533,N_8659);
and U9599 (N_9599,N_8516,N_8011);
nand U9600 (N_9600,N_8333,N_8887);
nor U9601 (N_9601,N_8971,N_8546);
nand U9602 (N_9602,N_8331,N_8605);
and U9603 (N_9603,N_8890,N_8608);
and U9604 (N_9604,N_8997,N_8032);
xnor U9605 (N_9605,N_8663,N_8712);
nor U9606 (N_9606,N_8530,N_8796);
or U9607 (N_9607,N_8044,N_8924);
nand U9608 (N_9608,N_8201,N_8769);
nor U9609 (N_9609,N_8855,N_8123);
nor U9610 (N_9610,N_8461,N_8372);
and U9611 (N_9611,N_8839,N_8634);
nor U9612 (N_9612,N_8953,N_8084);
or U9613 (N_9613,N_8616,N_8615);
or U9614 (N_9614,N_8413,N_8045);
nand U9615 (N_9615,N_8788,N_8718);
nand U9616 (N_9616,N_8411,N_8237);
nor U9617 (N_9617,N_8931,N_8659);
nand U9618 (N_9618,N_8781,N_8429);
nor U9619 (N_9619,N_8867,N_8430);
nand U9620 (N_9620,N_8888,N_8156);
and U9621 (N_9621,N_8382,N_8332);
and U9622 (N_9622,N_8662,N_8540);
nand U9623 (N_9623,N_8390,N_8981);
and U9624 (N_9624,N_8283,N_8394);
nand U9625 (N_9625,N_8940,N_8863);
nor U9626 (N_9626,N_8065,N_8367);
nor U9627 (N_9627,N_8684,N_8321);
or U9628 (N_9628,N_8018,N_8860);
and U9629 (N_9629,N_8912,N_8943);
nor U9630 (N_9630,N_8106,N_8444);
and U9631 (N_9631,N_8066,N_8097);
or U9632 (N_9632,N_8058,N_8791);
nand U9633 (N_9633,N_8841,N_8107);
nor U9634 (N_9634,N_8822,N_8595);
nand U9635 (N_9635,N_8598,N_8030);
and U9636 (N_9636,N_8109,N_8198);
or U9637 (N_9637,N_8896,N_8523);
nand U9638 (N_9638,N_8635,N_8403);
or U9639 (N_9639,N_8097,N_8098);
and U9640 (N_9640,N_8914,N_8618);
and U9641 (N_9641,N_8529,N_8293);
or U9642 (N_9642,N_8877,N_8702);
and U9643 (N_9643,N_8188,N_8585);
and U9644 (N_9644,N_8545,N_8888);
or U9645 (N_9645,N_8010,N_8089);
nand U9646 (N_9646,N_8737,N_8158);
and U9647 (N_9647,N_8474,N_8293);
nor U9648 (N_9648,N_8714,N_8135);
and U9649 (N_9649,N_8566,N_8584);
or U9650 (N_9650,N_8099,N_8458);
nor U9651 (N_9651,N_8373,N_8229);
or U9652 (N_9652,N_8593,N_8762);
or U9653 (N_9653,N_8747,N_8006);
and U9654 (N_9654,N_8458,N_8609);
nor U9655 (N_9655,N_8758,N_8304);
nor U9656 (N_9656,N_8719,N_8039);
nor U9657 (N_9657,N_8024,N_8271);
and U9658 (N_9658,N_8413,N_8443);
or U9659 (N_9659,N_8253,N_8175);
nand U9660 (N_9660,N_8127,N_8507);
nand U9661 (N_9661,N_8830,N_8941);
nor U9662 (N_9662,N_8789,N_8413);
xnor U9663 (N_9663,N_8382,N_8540);
nand U9664 (N_9664,N_8012,N_8486);
or U9665 (N_9665,N_8278,N_8492);
or U9666 (N_9666,N_8903,N_8025);
nor U9667 (N_9667,N_8099,N_8689);
nand U9668 (N_9668,N_8280,N_8222);
nand U9669 (N_9669,N_8586,N_8099);
xnor U9670 (N_9670,N_8831,N_8350);
and U9671 (N_9671,N_8443,N_8441);
nand U9672 (N_9672,N_8940,N_8363);
nand U9673 (N_9673,N_8543,N_8523);
nor U9674 (N_9674,N_8721,N_8756);
nand U9675 (N_9675,N_8686,N_8938);
nor U9676 (N_9676,N_8939,N_8209);
nor U9677 (N_9677,N_8298,N_8958);
or U9678 (N_9678,N_8949,N_8521);
or U9679 (N_9679,N_8859,N_8061);
nor U9680 (N_9680,N_8090,N_8543);
and U9681 (N_9681,N_8030,N_8705);
nand U9682 (N_9682,N_8209,N_8483);
or U9683 (N_9683,N_8205,N_8889);
or U9684 (N_9684,N_8313,N_8575);
and U9685 (N_9685,N_8459,N_8668);
xor U9686 (N_9686,N_8629,N_8954);
nand U9687 (N_9687,N_8805,N_8622);
or U9688 (N_9688,N_8155,N_8829);
nor U9689 (N_9689,N_8324,N_8955);
and U9690 (N_9690,N_8739,N_8875);
nor U9691 (N_9691,N_8613,N_8969);
xor U9692 (N_9692,N_8300,N_8854);
xor U9693 (N_9693,N_8830,N_8998);
nor U9694 (N_9694,N_8657,N_8251);
or U9695 (N_9695,N_8932,N_8777);
nor U9696 (N_9696,N_8281,N_8602);
nor U9697 (N_9697,N_8479,N_8249);
nand U9698 (N_9698,N_8695,N_8605);
nor U9699 (N_9699,N_8913,N_8889);
or U9700 (N_9700,N_8058,N_8943);
nor U9701 (N_9701,N_8859,N_8595);
nor U9702 (N_9702,N_8088,N_8309);
nor U9703 (N_9703,N_8241,N_8809);
and U9704 (N_9704,N_8613,N_8695);
nand U9705 (N_9705,N_8451,N_8388);
and U9706 (N_9706,N_8980,N_8473);
nand U9707 (N_9707,N_8461,N_8578);
nor U9708 (N_9708,N_8627,N_8559);
nand U9709 (N_9709,N_8641,N_8581);
or U9710 (N_9710,N_8169,N_8216);
or U9711 (N_9711,N_8015,N_8311);
nor U9712 (N_9712,N_8822,N_8476);
and U9713 (N_9713,N_8877,N_8546);
nand U9714 (N_9714,N_8251,N_8828);
nand U9715 (N_9715,N_8530,N_8688);
and U9716 (N_9716,N_8271,N_8681);
or U9717 (N_9717,N_8050,N_8963);
nand U9718 (N_9718,N_8000,N_8527);
nand U9719 (N_9719,N_8588,N_8241);
nor U9720 (N_9720,N_8991,N_8397);
nand U9721 (N_9721,N_8175,N_8219);
and U9722 (N_9722,N_8788,N_8117);
and U9723 (N_9723,N_8165,N_8253);
and U9724 (N_9724,N_8365,N_8118);
nand U9725 (N_9725,N_8216,N_8651);
nor U9726 (N_9726,N_8978,N_8336);
or U9727 (N_9727,N_8377,N_8973);
or U9728 (N_9728,N_8868,N_8437);
nand U9729 (N_9729,N_8733,N_8017);
nor U9730 (N_9730,N_8088,N_8078);
or U9731 (N_9731,N_8844,N_8424);
or U9732 (N_9732,N_8560,N_8549);
nor U9733 (N_9733,N_8769,N_8991);
nand U9734 (N_9734,N_8386,N_8760);
nor U9735 (N_9735,N_8553,N_8861);
or U9736 (N_9736,N_8124,N_8395);
nand U9737 (N_9737,N_8108,N_8359);
and U9738 (N_9738,N_8061,N_8337);
nand U9739 (N_9739,N_8530,N_8851);
nor U9740 (N_9740,N_8813,N_8107);
nor U9741 (N_9741,N_8186,N_8004);
and U9742 (N_9742,N_8591,N_8234);
nand U9743 (N_9743,N_8822,N_8389);
or U9744 (N_9744,N_8612,N_8531);
and U9745 (N_9745,N_8036,N_8977);
nand U9746 (N_9746,N_8139,N_8118);
nand U9747 (N_9747,N_8798,N_8632);
and U9748 (N_9748,N_8105,N_8288);
nand U9749 (N_9749,N_8861,N_8278);
and U9750 (N_9750,N_8543,N_8172);
or U9751 (N_9751,N_8533,N_8614);
or U9752 (N_9752,N_8497,N_8133);
and U9753 (N_9753,N_8667,N_8962);
nand U9754 (N_9754,N_8661,N_8503);
nand U9755 (N_9755,N_8531,N_8904);
and U9756 (N_9756,N_8972,N_8125);
nand U9757 (N_9757,N_8377,N_8028);
and U9758 (N_9758,N_8508,N_8897);
and U9759 (N_9759,N_8394,N_8463);
nor U9760 (N_9760,N_8767,N_8290);
nand U9761 (N_9761,N_8602,N_8492);
nand U9762 (N_9762,N_8206,N_8037);
and U9763 (N_9763,N_8859,N_8419);
and U9764 (N_9764,N_8880,N_8638);
nor U9765 (N_9765,N_8751,N_8532);
nor U9766 (N_9766,N_8284,N_8984);
and U9767 (N_9767,N_8586,N_8881);
nand U9768 (N_9768,N_8583,N_8386);
nand U9769 (N_9769,N_8395,N_8753);
nor U9770 (N_9770,N_8675,N_8950);
or U9771 (N_9771,N_8914,N_8624);
and U9772 (N_9772,N_8265,N_8966);
xnor U9773 (N_9773,N_8321,N_8669);
or U9774 (N_9774,N_8417,N_8029);
nand U9775 (N_9775,N_8336,N_8472);
nor U9776 (N_9776,N_8699,N_8649);
and U9777 (N_9777,N_8031,N_8060);
nand U9778 (N_9778,N_8109,N_8795);
nand U9779 (N_9779,N_8372,N_8071);
and U9780 (N_9780,N_8416,N_8351);
nor U9781 (N_9781,N_8292,N_8083);
nor U9782 (N_9782,N_8679,N_8091);
nand U9783 (N_9783,N_8066,N_8268);
and U9784 (N_9784,N_8107,N_8428);
and U9785 (N_9785,N_8975,N_8040);
or U9786 (N_9786,N_8011,N_8067);
nand U9787 (N_9787,N_8197,N_8314);
nor U9788 (N_9788,N_8233,N_8505);
nor U9789 (N_9789,N_8609,N_8158);
nand U9790 (N_9790,N_8108,N_8624);
or U9791 (N_9791,N_8337,N_8806);
nor U9792 (N_9792,N_8744,N_8628);
and U9793 (N_9793,N_8927,N_8673);
nand U9794 (N_9794,N_8110,N_8514);
and U9795 (N_9795,N_8245,N_8048);
and U9796 (N_9796,N_8189,N_8989);
nand U9797 (N_9797,N_8113,N_8450);
or U9798 (N_9798,N_8472,N_8602);
nor U9799 (N_9799,N_8402,N_8042);
and U9800 (N_9800,N_8499,N_8570);
nor U9801 (N_9801,N_8622,N_8877);
nand U9802 (N_9802,N_8968,N_8429);
and U9803 (N_9803,N_8768,N_8866);
or U9804 (N_9804,N_8306,N_8664);
nand U9805 (N_9805,N_8450,N_8455);
nand U9806 (N_9806,N_8865,N_8635);
nand U9807 (N_9807,N_8425,N_8794);
nand U9808 (N_9808,N_8400,N_8944);
or U9809 (N_9809,N_8077,N_8144);
nand U9810 (N_9810,N_8205,N_8427);
or U9811 (N_9811,N_8615,N_8007);
nor U9812 (N_9812,N_8747,N_8761);
or U9813 (N_9813,N_8586,N_8342);
nor U9814 (N_9814,N_8694,N_8733);
nand U9815 (N_9815,N_8806,N_8995);
and U9816 (N_9816,N_8429,N_8796);
nor U9817 (N_9817,N_8811,N_8905);
xnor U9818 (N_9818,N_8866,N_8223);
or U9819 (N_9819,N_8464,N_8697);
or U9820 (N_9820,N_8264,N_8568);
nor U9821 (N_9821,N_8974,N_8878);
nand U9822 (N_9822,N_8255,N_8942);
and U9823 (N_9823,N_8962,N_8380);
nor U9824 (N_9824,N_8091,N_8278);
nor U9825 (N_9825,N_8964,N_8369);
nor U9826 (N_9826,N_8793,N_8029);
and U9827 (N_9827,N_8304,N_8847);
or U9828 (N_9828,N_8763,N_8448);
or U9829 (N_9829,N_8099,N_8250);
nand U9830 (N_9830,N_8306,N_8809);
nor U9831 (N_9831,N_8917,N_8490);
or U9832 (N_9832,N_8735,N_8615);
nor U9833 (N_9833,N_8659,N_8007);
and U9834 (N_9834,N_8100,N_8936);
or U9835 (N_9835,N_8711,N_8468);
nor U9836 (N_9836,N_8605,N_8806);
nand U9837 (N_9837,N_8805,N_8795);
nor U9838 (N_9838,N_8471,N_8328);
and U9839 (N_9839,N_8691,N_8734);
nand U9840 (N_9840,N_8682,N_8378);
nand U9841 (N_9841,N_8671,N_8977);
and U9842 (N_9842,N_8077,N_8896);
or U9843 (N_9843,N_8138,N_8666);
nand U9844 (N_9844,N_8448,N_8160);
nor U9845 (N_9845,N_8028,N_8900);
nand U9846 (N_9846,N_8225,N_8536);
nand U9847 (N_9847,N_8928,N_8547);
or U9848 (N_9848,N_8758,N_8520);
or U9849 (N_9849,N_8301,N_8104);
nand U9850 (N_9850,N_8192,N_8824);
nor U9851 (N_9851,N_8746,N_8303);
nor U9852 (N_9852,N_8993,N_8410);
and U9853 (N_9853,N_8464,N_8980);
or U9854 (N_9854,N_8028,N_8670);
or U9855 (N_9855,N_8207,N_8874);
nor U9856 (N_9856,N_8803,N_8914);
nor U9857 (N_9857,N_8190,N_8616);
xor U9858 (N_9858,N_8015,N_8765);
and U9859 (N_9859,N_8652,N_8333);
or U9860 (N_9860,N_8092,N_8211);
nor U9861 (N_9861,N_8010,N_8923);
nand U9862 (N_9862,N_8954,N_8076);
and U9863 (N_9863,N_8853,N_8375);
and U9864 (N_9864,N_8527,N_8027);
and U9865 (N_9865,N_8730,N_8177);
or U9866 (N_9866,N_8229,N_8574);
and U9867 (N_9867,N_8499,N_8823);
nand U9868 (N_9868,N_8886,N_8852);
nor U9869 (N_9869,N_8773,N_8319);
and U9870 (N_9870,N_8627,N_8038);
nand U9871 (N_9871,N_8457,N_8687);
and U9872 (N_9872,N_8381,N_8360);
and U9873 (N_9873,N_8806,N_8905);
xnor U9874 (N_9874,N_8092,N_8146);
nor U9875 (N_9875,N_8991,N_8004);
or U9876 (N_9876,N_8949,N_8490);
or U9877 (N_9877,N_8843,N_8876);
nand U9878 (N_9878,N_8148,N_8136);
nor U9879 (N_9879,N_8209,N_8770);
and U9880 (N_9880,N_8332,N_8321);
nand U9881 (N_9881,N_8273,N_8039);
nand U9882 (N_9882,N_8352,N_8981);
or U9883 (N_9883,N_8579,N_8704);
nand U9884 (N_9884,N_8151,N_8137);
nor U9885 (N_9885,N_8551,N_8940);
or U9886 (N_9886,N_8612,N_8763);
nand U9887 (N_9887,N_8202,N_8294);
nand U9888 (N_9888,N_8715,N_8502);
or U9889 (N_9889,N_8091,N_8467);
or U9890 (N_9890,N_8881,N_8754);
nor U9891 (N_9891,N_8679,N_8904);
nor U9892 (N_9892,N_8953,N_8044);
nand U9893 (N_9893,N_8695,N_8462);
and U9894 (N_9894,N_8920,N_8323);
and U9895 (N_9895,N_8923,N_8517);
nor U9896 (N_9896,N_8700,N_8615);
nand U9897 (N_9897,N_8704,N_8721);
or U9898 (N_9898,N_8816,N_8805);
nor U9899 (N_9899,N_8965,N_8763);
and U9900 (N_9900,N_8818,N_8843);
or U9901 (N_9901,N_8277,N_8791);
or U9902 (N_9902,N_8503,N_8933);
nand U9903 (N_9903,N_8812,N_8466);
and U9904 (N_9904,N_8383,N_8330);
nand U9905 (N_9905,N_8251,N_8150);
or U9906 (N_9906,N_8812,N_8116);
and U9907 (N_9907,N_8464,N_8223);
nor U9908 (N_9908,N_8670,N_8371);
nand U9909 (N_9909,N_8597,N_8007);
or U9910 (N_9910,N_8427,N_8288);
and U9911 (N_9911,N_8563,N_8669);
nand U9912 (N_9912,N_8888,N_8082);
and U9913 (N_9913,N_8389,N_8835);
nand U9914 (N_9914,N_8468,N_8032);
or U9915 (N_9915,N_8565,N_8754);
xnor U9916 (N_9916,N_8009,N_8287);
or U9917 (N_9917,N_8244,N_8727);
nand U9918 (N_9918,N_8847,N_8047);
and U9919 (N_9919,N_8460,N_8862);
and U9920 (N_9920,N_8204,N_8575);
nor U9921 (N_9921,N_8773,N_8191);
nor U9922 (N_9922,N_8055,N_8281);
or U9923 (N_9923,N_8954,N_8223);
nand U9924 (N_9924,N_8439,N_8867);
or U9925 (N_9925,N_8807,N_8522);
or U9926 (N_9926,N_8562,N_8812);
nand U9927 (N_9927,N_8227,N_8135);
and U9928 (N_9928,N_8219,N_8315);
nor U9929 (N_9929,N_8682,N_8611);
or U9930 (N_9930,N_8142,N_8108);
and U9931 (N_9931,N_8720,N_8544);
and U9932 (N_9932,N_8803,N_8164);
and U9933 (N_9933,N_8963,N_8600);
nor U9934 (N_9934,N_8209,N_8980);
xor U9935 (N_9935,N_8975,N_8904);
and U9936 (N_9936,N_8767,N_8403);
nor U9937 (N_9937,N_8634,N_8998);
and U9938 (N_9938,N_8342,N_8267);
and U9939 (N_9939,N_8880,N_8218);
xnor U9940 (N_9940,N_8144,N_8948);
or U9941 (N_9941,N_8942,N_8461);
and U9942 (N_9942,N_8450,N_8987);
nor U9943 (N_9943,N_8056,N_8428);
and U9944 (N_9944,N_8064,N_8456);
or U9945 (N_9945,N_8544,N_8687);
nor U9946 (N_9946,N_8981,N_8770);
nand U9947 (N_9947,N_8779,N_8108);
and U9948 (N_9948,N_8354,N_8685);
nand U9949 (N_9949,N_8015,N_8949);
and U9950 (N_9950,N_8110,N_8334);
nor U9951 (N_9951,N_8467,N_8226);
and U9952 (N_9952,N_8538,N_8073);
or U9953 (N_9953,N_8668,N_8663);
nand U9954 (N_9954,N_8907,N_8904);
nor U9955 (N_9955,N_8817,N_8565);
or U9956 (N_9956,N_8335,N_8680);
nand U9957 (N_9957,N_8351,N_8991);
nor U9958 (N_9958,N_8737,N_8299);
and U9959 (N_9959,N_8003,N_8780);
nand U9960 (N_9960,N_8728,N_8428);
nand U9961 (N_9961,N_8499,N_8373);
nor U9962 (N_9962,N_8891,N_8771);
and U9963 (N_9963,N_8105,N_8820);
nand U9964 (N_9964,N_8231,N_8664);
or U9965 (N_9965,N_8110,N_8402);
and U9966 (N_9966,N_8197,N_8882);
nand U9967 (N_9967,N_8115,N_8582);
or U9968 (N_9968,N_8212,N_8927);
and U9969 (N_9969,N_8160,N_8592);
or U9970 (N_9970,N_8066,N_8509);
nor U9971 (N_9971,N_8604,N_8603);
or U9972 (N_9972,N_8196,N_8723);
and U9973 (N_9973,N_8654,N_8779);
nand U9974 (N_9974,N_8684,N_8213);
or U9975 (N_9975,N_8128,N_8640);
nand U9976 (N_9976,N_8105,N_8851);
xor U9977 (N_9977,N_8928,N_8692);
and U9978 (N_9978,N_8143,N_8255);
xor U9979 (N_9979,N_8745,N_8184);
nand U9980 (N_9980,N_8572,N_8089);
or U9981 (N_9981,N_8939,N_8299);
nor U9982 (N_9982,N_8759,N_8314);
and U9983 (N_9983,N_8448,N_8787);
nand U9984 (N_9984,N_8358,N_8293);
nand U9985 (N_9985,N_8847,N_8088);
and U9986 (N_9986,N_8685,N_8710);
or U9987 (N_9987,N_8135,N_8553);
nand U9988 (N_9988,N_8176,N_8523);
or U9989 (N_9989,N_8005,N_8223);
nor U9990 (N_9990,N_8060,N_8705);
nor U9991 (N_9991,N_8733,N_8842);
or U9992 (N_9992,N_8773,N_8430);
and U9993 (N_9993,N_8779,N_8377);
nand U9994 (N_9994,N_8644,N_8770);
nand U9995 (N_9995,N_8547,N_8379);
or U9996 (N_9996,N_8302,N_8101);
nand U9997 (N_9997,N_8137,N_8261);
and U9998 (N_9998,N_8736,N_8404);
nand U9999 (N_9999,N_8905,N_8489);
and UO_0 (O_0,N_9625,N_9669);
and UO_1 (O_1,N_9379,N_9296);
and UO_2 (O_2,N_9491,N_9744);
or UO_3 (O_3,N_9888,N_9824);
nand UO_4 (O_4,N_9701,N_9801);
nor UO_5 (O_5,N_9278,N_9402);
and UO_6 (O_6,N_9364,N_9469);
or UO_7 (O_7,N_9093,N_9566);
nor UO_8 (O_8,N_9401,N_9212);
nor UO_9 (O_9,N_9443,N_9041);
and UO_10 (O_10,N_9799,N_9941);
nand UO_11 (O_11,N_9440,N_9189);
nor UO_12 (O_12,N_9028,N_9785);
nor UO_13 (O_13,N_9319,N_9829);
nor UO_14 (O_14,N_9606,N_9490);
and UO_15 (O_15,N_9851,N_9155);
nand UO_16 (O_16,N_9183,N_9609);
and UO_17 (O_17,N_9315,N_9865);
nor UO_18 (O_18,N_9232,N_9917);
or UO_19 (O_19,N_9772,N_9036);
nand UO_20 (O_20,N_9235,N_9707);
and UO_21 (O_21,N_9570,N_9731);
nand UO_22 (O_22,N_9321,N_9124);
or UO_23 (O_23,N_9020,N_9494);
or UO_24 (O_24,N_9386,N_9287);
and UO_25 (O_25,N_9295,N_9162);
and UO_26 (O_26,N_9030,N_9144);
or UO_27 (O_27,N_9070,N_9456);
nand UO_28 (O_28,N_9485,N_9417);
nor UO_29 (O_29,N_9045,N_9457);
nor UO_30 (O_30,N_9782,N_9989);
and UO_31 (O_31,N_9329,N_9381);
or UO_32 (O_32,N_9695,N_9786);
nor UO_33 (O_33,N_9397,N_9895);
nor UO_34 (O_34,N_9460,N_9657);
and UO_35 (O_35,N_9811,N_9013);
nand UO_36 (O_36,N_9913,N_9780);
nor UO_37 (O_37,N_9055,N_9825);
and UO_38 (O_38,N_9252,N_9520);
nor UO_39 (O_39,N_9065,N_9451);
or UO_40 (O_40,N_9131,N_9970);
and UO_41 (O_41,N_9798,N_9638);
nand UO_42 (O_42,N_9269,N_9437);
nand UO_43 (O_43,N_9057,N_9463);
nor UO_44 (O_44,N_9756,N_9213);
xor UO_45 (O_45,N_9271,N_9699);
nor UO_46 (O_46,N_9503,N_9170);
nor UO_47 (O_47,N_9080,N_9412);
or UO_48 (O_48,N_9858,N_9420);
and UO_49 (O_49,N_9653,N_9072);
or UO_50 (O_50,N_9433,N_9807);
nor UO_51 (O_51,N_9445,N_9083);
nand UO_52 (O_52,N_9975,N_9671);
nand UO_53 (O_53,N_9761,N_9035);
nand UO_54 (O_54,N_9769,N_9151);
nand UO_55 (O_55,N_9593,N_9636);
nor UO_56 (O_56,N_9371,N_9733);
nand UO_57 (O_57,N_9037,N_9675);
nor UO_58 (O_58,N_9794,N_9471);
nor UO_59 (O_59,N_9129,N_9889);
or UO_60 (O_60,N_9748,N_9499);
nor UO_61 (O_61,N_9366,N_9353);
or UO_62 (O_62,N_9834,N_9474);
nor UO_63 (O_63,N_9727,N_9288);
or UO_64 (O_64,N_9309,N_9899);
nand UO_65 (O_65,N_9481,N_9467);
and UO_66 (O_66,N_9119,N_9776);
or UO_67 (O_67,N_9758,N_9926);
and UO_68 (O_68,N_9512,N_9539);
nand UO_69 (O_69,N_9425,N_9850);
and UO_70 (O_70,N_9424,N_9197);
nand UO_71 (O_71,N_9831,N_9588);
nand UO_72 (O_72,N_9432,N_9999);
nor UO_73 (O_73,N_9614,N_9584);
and UO_74 (O_74,N_9549,N_9613);
or UO_75 (O_75,N_9002,N_9979);
nor UO_76 (O_76,N_9383,N_9971);
or UO_77 (O_77,N_9160,N_9308);
and UO_78 (O_78,N_9513,N_9479);
nand UO_79 (O_79,N_9202,N_9001);
nand UO_80 (O_80,N_9942,N_9578);
nand UO_81 (O_81,N_9016,N_9908);
nor UO_82 (O_82,N_9249,N_9310);
nor UO_83 (O_83,N_9947,N_9459);
or UO_84 (O_84,N_9873,N_9784);
or UO_85 (O_85,N_9668,N_9869);
and UO_86 (O_86,N_9262,N_9218);
or UO_87 (O_87,N_9062,N_9079);
nand UO_88 (O_88,N_9587,N_9767);
nand UO_89 (O_89,N_9883,N_9209);
xor UO_90 (O_90,N_9964,N_9838);
or UO_91 (O_91,N_9012,N_9900);
and UO_92 (O_92,N_9489,N_9418);
nand UO_93 (O_93,N_9763,N_9674);
or UO_94 (O_94,N_9981,N_9577);
or UO_95 (O_95,N_9090,N_9227);
or UO_96 (O_96,N_9203,N_9049);
nor UO_97 (O_97,N_9709,N_9690);
and UO_98 (O_98,N_9634,N_9648);
and UO_99 (O_99,N_9832,N_9069);
and UO_100 (O_100,N_9804,N_9642);
and UO_101 (O_101,N_9809,N_9810);
nor UO_102 (O_102,N_9454,N_9447);
and UO_103 (O_103,N_9497,N_9714);
nor UO_104 (O_104,N_9562,N_9555);
nor UO_105 (O_105,N_9931,N_9560);
and UO_106 (O_106,N_9132,N_9268);
nor UO_107 (O_107,N_9641,N_9110);
or UO_108 (O_108,N_9253,N_9184);
nand UO_109 (O_109,N_9328,N_9396);
or UO_110 (O_110,N_9033,N_9403);
and UO_111 (O_111,N_9984,N_9747);
xnor UO_112 (O_112,N_9439,N_9177);
or UO_113 (O_113,N_9201,N_9726);
or UO_114 (O_114,N_9380,N_9478);
or UO_115 (O_115,N_9219,N_9918);
or UO_116 (O_116,N_9392,N_9568);
nand UO_117 (O_117,N_9795,N_9639);
nor UO_118 (O_118,N_9333,N_9152);
and UO_119 (O_119,N_9879,N_9708);
nand UO_120 (O_120,N_9534,N_9571);
and UO_121 (O_121,N_9482,N_9522);
nor UO_122 (O_122,N_9140,N_9157);
nand UO_123 (O_123,N_9629,N_9221);
nand UO_124 (O_124,N_9250,N_9382);
nand UO_125 (O_125,N_9737,N_9870);
nor UO_126 (O_126,N_9738,N_9398);
and UO_127 (O_127,N_9764,N_9027);
or UO_128 (O_128,N_9265,N_9349);
and UO_129 (O_129,N_9821,N_9969);
and UO_130 (O_130,N_9043,N_9082);
nor UO_131 (O_131,N_9640,N_9556);
xnor UO_132 (O_132,N_9230,N_9031);
nor UO_133 (O_133,N_9951,N_9682);
nand UO_134 (O_134,N_9646,N_9912);
xnor UO_135 (O_135,N_9150,N_9360);
and UO_136 (O_136,N_9506,N_9040);
and UO_137 (O_137,N_9102,N_9073);
nand UO_138 (O_138,N_9061,N_9192);
and UO_139 (O_139,N_9359,N_9188);
xor UO_140 (O_140,N_9435,N_9346);
nor UO_141 (O_141,N_9470,N_9475);
nor UO_142 (O_142,N_9289,N_9930);
nor UO_143 (O_143,N_9210,N_9370);
nand UO_144 (O_144,N_9903,N_9029);
nand UO_145 (O_145,N_9298,N_9117);
nor UO_146 (O_146,N_9906,N_9014);
or UO_147 (O_147,N_9176,N_9751);
and UO_148 (O_148,N_9750,N_9796);
nand UO_149 (O_149,N_9994,N_9270);
nand UO_150 (O_150,N_9987,N_9755);
nor UO_151 (O_151,N_9676,N_9967);
and UO_152 (O_152,N_9797,N_9258);
or UO_153 (O_153,N_9960,N_9948);
nand UO_154 (O_154,N_9423,N_9363);
and UO_155 (O_155,N_9523,N_9441);
and UO_156 (O_156,N_9427,N_9728);
and UO_157 (O_157,N_9004,N_9876);
or UO_158 (O_158,N_9881,N_9193);
nor UO_159 (O_159,N_9458,N_9226);
nand UO_160 (O_160,N_9774,N_9856);
xnor UO_161 (O_161,N_9374,N_9276);
nor UO_162 (O_162,N_9871,N_9718);
nand UO_163 (O_163,N_9125,N_9375);
nand UO_164 (O_164,N_9692,N_9200);
nor UO_165 (O_165,N_9112,N_9108);
nor UO_166 (O_166,N_9091,N_9605);
and UO_167 (O_167,N_9990,N_9376);
nand UO_168 (O_168,N_9581,N_9312);
xnor UO_169 (O_169,N_9836,N_9863);
nor UO_170 (O_170,N_9317,N_9206);
or UO_171 (O_171,N_9995,N_9938);
or UO_172 (O_172,N_9179,N_9934);
nor UO_173 (O_173,N_9904,N_9135);
and UO_174 (O_174,N_9922,N_9067);
or UO_175 (O_175,N_9923,N_9944);
or UO_176 (O_176,N_9963,N_9788);
nand UO_177 (O_177,N_9837,N_9126);
nand UO_178 (O_178,N_9596,N_9046);
nand UO_179 (O_179,N_9414,N_9666);
and UO_180 (O_180,N_9436,N_9518);
or UO_181 (O_181,N_9515,N_9600);
nor UO_182 (O_182,N_9717,N_9525);
nor UO_183 (O_183,N_9473,N_9945);
nor UO_184 (O_184,N_9331,N_9540);
and UO_185 (O_185,N_9064,N_9721);
nor UO_186 (O_186,N_9056,N_9407);
nor UO_187 (O_187,N_9186,N_9204);
nor UO_188 (O_188,N_9385,N_9257);
xor UO_189 (O_189,N_9632,N_9338);
xor UO_190 (O_190,N_9365,N_9053);
and UO_191 (O_191,N_9263,N_9530);
nor UO_192 (O_192,N_9452,N_9734);
and UO_193 (O_193,N_9134,N_9318);
and UO_194 (O_194,N_9448,N_9618);
or UO_195 (O_195,N_9130,N_9431);
nor UO_196 (O_196,N_9563,N_9006);
or UO_197 (O_197,N_9567,N_9988);
nand UO_198 (O_198,N_9216,N_9575);
nand UO_199 (O_199,N_9136,N_9116);
or UO_200 (O_200,N_9720,N_9591);
nor UO_201 (O_201,N_9991,N_9369);
nand UO_202 (O_202,N_9616,N_9624);
nand UO_203 (O_203,N_9211,N_9167);
nand UO_204 (O_204,N_9389,N_9550);
and UO_205 (O_205,N_9815,N_9816);
and UO_206 (O_206,N_9808,N_9827);
and UO_207 (O_207,N_9351,N_9509);
or UO_208 (O_208,N_9408,N_9345);
nand UO_209 (O_209,N_9251,N_9196);
xor UO_210 (O_210,N_9855,N_9956);
nor UO_211 (O_211,N_9996,N_9238);
nor UO_212 (O_212,N_9933,N_9878);
nand UO_213 (O_213,N_9792,N_9754);
or UO_214 (O_214,N_9628,N_9156);
or UO_215 (O_215,N_9356,N_9667);
nand UO_216 (O_216,N_9762,N_9773);
nand UO_217 (O_217,N_9533,N_9521);
and UO_218 (O_218,N_9388,N_9501);
and UO_219 (O_219,N_9915,N_9283);
nor UO_220 (O_220,N_9145,N_9677);
nor UO_221 (O_221,N_9602,N_9921);
nand UO_222 (O_222,N_9358,N_9480);
or UO_223 (O_223,N_9670,N_9580);
or UO_224 (O_224,N_9248,N_9927);
and UO_225 (O_225,N_9940,N_9281);
and UO_226 (O_226,N_9617,N_9565);
or UO_227 (O_227,N_9847,N_9254);
or UO_228 (O_228,N_9696,N_9866);
nand UO_229 (O_229,N_9384,N_9620);
and UO_230 (O_230,N_9531,N_9925);
nand UO_231 (O_231,N_9510,N_9954);
nand UO_232 (O_232,N_9495,N_9259);
xor UO_233 (O_233,N_9965,N_9553);
and UO_234 (O_234,N_9172,N_9500);
nand UO_235 (O_235,N_9305,N_9654);
and UO_236 (O_236,N_9099,N_9453);
nand UO_237 (O_237,N_9656,N_9461);
and UO_238 (O_238,N_9504,N_9687);
or UO_239 (O_239,N_9400,N_9542);
and UO_240 (O_240,N_9973,N_9817);
or UO_241 (O_241,N_9139,N_9178);
or UO_242 (O_242,N_9180,N_9141);
nor UO_243 (O_243,N_9828,N_9455);
or UO_244 (O_244,N_9688,N_9887);
and UO_245 (O_245,N_9896,N_9122);
nand UO_246 (O_246,N_9548,N_9980);
nor UO_247 (O_247,N_9631,N_9611);
or UO_248 (O_248,N_9972,N_9468);
and UO_249 (O_249,N_9929,N_9303);
nand UO_250 (O_250,N_9875,N_9355);
and UO_251 (O_251,N_9823,N_9864);
and UO_252 (O_252,N_9789,N_9127);
and UO_253 (O_253,N_9739,N_9937);
and UO_254 (O_254,N_9077,N_9604);
or UO_255 (O_255,N_9819,N_9324);
nand UO_256 (O_256,N_9010,N_9505);
nand UO_257 (O_257,N_9021,N_9208);
nand UO_258 (O_258,N_9089,N_9757);
and UO_259 (O_259,N_9939,N_9284);
nand UO_260 (O_260,N_9777,N_9068);
and UO_261 (O_261,N_9015,N_9672);
and UO_262 (O_262,N_9241,N_9868);
or UO_263 (O_263,N_9813,N_9377);
nor UO_264 (O_264,N_9048,N_9543);
nand UO_265 (O_265,N_9217,N_9835);
nand UO_266 (O_266,N_9233,N_9623);
xnor UO_267 (O_267,N_9582,N_9422);
nor UO_268 (O_268,N_9507,N_9859);
or UO_269 (O_269,N_9545,N_9341);
nand UO_270 (O_270,N_9861,N_9662);
nor UO_271 (O_271,N_9541,N_9845);
nor UO_272 (O_272,N_9256,N_9450);
nand UO_273 (O_273,N_9434,N_9898);
nand UO_274 (O_274,N_9000,N_9168);
nor UO_275 (O_275,N_9337,N_9444);
or UO_276 (O_276,N_9322,N_9891);
or UO_277 (O_277,N_9092,N_9771);
or UO_278 (O_278,N_9063,N_9853);
nor UO_279 (O_279,N_9818,N_9966);
nor UO_280 (O_280,N_9590,N_9703);
nor UO_281 (O_281,N_9462,N_9914);
nor UO_282 (O_282,N_9350,N_9952);
or UO_283 (O_283,N_9017,N_9985);
and UO_284 (O_284,N_9274,N_9830);
nand UO_285 (O_285,N_9694,N_9084);
or UO_286 (O_286,N_9411,N_9658);
nor UO_287 (O_287,N_9689,N_9008);
or UO_288 (O_288,N_9273,N_9222);
or UO_289 (O_289,N_9992,N_9279);
nor UO_290 (O_290,N_9702,N_9399);
and UO_291 (O_291,N_9215,N_9742);
or UO_292 (O_292,N_9320,N_9595);
or UO_293 (O_293,N_9993,N_9982);
and UO_294 (O_294,N_9569,N_9877);
and UO_295 (O_295,N_9950,N_9519);
and UO_296 (O_296,N_9007,N_9621);
nor UO_297 (O_297,N_9104,N_9759);
nor UO_298 (O_298,N_9340,N_9404);
nor UO_299 (O_299,N_9449,N_9723);
nor UO_300 (O_300,N_9722,N_9928);
nor UO_301 (O_301,N_9693,N_9299);
nor UO_302 (O_302,N_9220,N_9109);
and UO_303 (O_303,N_9793,N_9790);
nor UO_304 (O_304,N_9976,N_9619);
and UO_305 (O_305,N_9214,N_9526);
and UO_306 (O_306,N_9103,N_9493);
nand UO_307 (O_307,N_9231,N_9100);
nand UO_308 (O_308,N_9111,N_9304);
and UO_309 (O_309,N_9022,N_9935);
nand UO_310 (O_310,N_9867,N_9635);
xor UO_311 (O_311,N_9466,N_9026);
and UO_312 (O_312,N_9032,N_9781);
or UO_313 (O_313,N_9622,N_9812);
nand UO_314 (O_314,N_9246,N_9054);
and UO_315 (O_315,N_9266,N_9332);
nor UO_316 (O_316,N_9665,N_9237);
and UO_317 (O_317,N_9649,N_9415);
nand UO_318 (O_318,N_9391,N_9292);
and UO_319 (O_319,N_9872,N_9806);
or UO_320 (O_320,N_9559,N_9775);
and UO_321 (O_321,N_9612,N_9583);
nand UO_322 (O_322,N_9038,N_9302);
nor UO_323 (O_323,N_9586,N_9874);
or UO_324 (O_324,N_9752,N_9442);
nor UO_325 (O_325,N_9405,N_9538);
nand UO_326 (O_326,N_9770,N_9347);
nand UO_327 (O_327,N_9713,N_9114);
nor UO_328 (O_328,N_9023,N_9882);
nor UO_329 (O_329,N_9892,N_9557);
and UO_330 (O_330,N_9191,N_9229);
and UO_331 (O_331,N_9361,N_9050);
nand UO_332 (O_332,N_9660,N_9949);
nor UO_333 (O_333,N_9961,N_9730);
nor UO_334 (O_334,N_9148,N_9743);
nor UO_335 (O_335,N_9146,N_9760);
or UO_336 (O_336,N_9516,N_9011);
nor UO_337 (O_337,N_9678,N_9164);
nand UO_338 (O_338,N_9496,N_9833);
nand UO_339 (O_339,N_9367,N_9686);
nand UO_340 (O_340,N_9645,N_9698);
and UO_341 (O_341,N_9153,N_9768);
and UO_342 (O_342,N_9143,N_9528);
or UO_343 (O_343,N_9920,N_9326);
nor UO_344 (O_344,N_9607,N_9650);
or UO_345 (O_345,N_9066,N_9290);
and UO_346 (O_346,N_9060,N_9169);
and UO_347 (O_347,N_9857,N_9907);
or UO_348 (O_348,N_9805,N_9511);
or UO_349 (O_349,N_9860,N_9524);
and UO_350 (O_350,N_9018,N_9814);
or UO_351 (O_351,N_9198,N_9843);
nor UO_352 (O_352,N_9339,N_9552);
or UO_353 (O_353,N_9615,N_9300);
and UO_354 (O_354,N_9745,N_9428);
and UO_355 (O_355,N_9862,N_9225);
or UO_356 (O_356,N_9142,N_9240);
nand UO_357 (O_357,N_9659,N_9476);
or UO_358 (O_358,N_9932,N_9086);
nor UO_359 (O_359,N_9390,N_9732);
nand UO_360 (O_360,N_9047,N_9009);
nor UO_361 (O_361,N_9044,N_9572);
and UO_362 (O_362,N_9651,N_9242);
and UO_363 (O_363,N_9924,N_9330);
or UO_364 (O_364,N_9003,N_9573);
nand UO_365 (O_365,N_9098,N_9753);
nand UO_366 (O_366,N_9313,N_9663);
nor UO_367 (O_367,N_9343,N_9729);
nor UO_368 (O_368,N_9826,N_9592);
or UO_369 (O_369,N_9911,N_9081);
nand UO_370 (O_370,N_9704,N_9395);
xnor UO_371 (O_371,N_9741,N_9630);
or UO_372 (O_372,N_9589,N_9679);
nor UO_373 (O_373,N_9438,N_9311);
or UO_374 (O_374,N_9844,N_9419);
nor UO_375 (O_375,N_9267,N_9165);
and UO_376 (O_376,N_9087,N_9239);
and UO_377 (O_377,N_9558,N_9706);
nand UO_378 (O_378,N_9071,N_9885);
nand UO_379 (O_379,N_9532,N_9551);
nor UO_380 (O_380,N_9195,N_9800);
and UO_381 (O_381,N_9194,N_9643);
xor UO_382 (O_382,N_9681,N_9464);
nor UO_383 (O_383,N_9357,N_9477);
or UO_384 (O_384,N_9137,N_9373);
or UO_385 (O_385,N_9546,N_9897);
nand UO_386 (O_386,N_9223,N_9652);
nor UO_387 (O_387,N_9159,N_9094);
nor UO_388 (O_388,N_9998,N_9352);
and UO_389 (O_389,N_9413,N_9410);
or UO_390 (O_390,N_9955,N_9393);
nand UO_391 (O_391,N_9166,N_9421);
xnor UO_392 (O_392,N_9749,N_9429);
or UO_393 (O_393,N_9236,N_9058);
and UO_394 (O_394,N_9585,N_9426);
and UO_395 (O_395,N_9502,N_9307);
nor UO_396 (O_396,N_9901,N_9154);
or UO_397 (O_397,N_9626,N_9536);
nor UO_398 (O_398,N_9247,N_9336);
and UO_399 (O_399,N_9959,N_9255);
and UO_400 (O_400,N_9051,N_9486);
or UO_401 (O_401,N_9601,N_9133);
or UO_402 (O_402,N_9115,N_9644);
and UO_403 (O_403,N_9842,N_9661);
nor UO_404 (O_404,N_9746,N_9547);
or UO_405 (O_405,N_9342,N_9783);
or UO_406 (O_406,N_9492,N_9088);
or UO_407 (O_407,N_9664,N_9803);
or UO_408 (O_408,N_9149,N_9778);
and UO_409 (O_409,N_9121,N_9095);
and UO_410 (O_410,N_9905,N_9181);
nor UO_411 (O_411,N_9936,N_9711);
or UO_412 (O_412,N_9498,N_9561);
and UO_413 (O_413,N_9120,N_9986);
nand UO_414 (O_414,N_9647,N_9085);
or UO_415 (O_415,N_9446,N_9291);
or UO_416 (O_416,N_9128,N_9724);
nor UO_417 (O_417,N_9323,N_9282);
nor UO_418 (O_418,N_9185,N_9484);
xor UO_419 (O_419,N_9406,N_9138);
or UO_420 (O_420,N_9544,N_9603);
or UO_421 (O_421,N_9107,N_9627);
nor UO_422 (O_422,N_9535,N_9019);
or UO_423 (O_423,N_9902,N_9576);
nand UO_424 (O_424,N_9234,N_9161);
nand UO_425 (O_425,N_9052,N_9372);
nor UO_426 (O_426,N_9113,N_9465);
and UO_427 (O_427,N_9285,N_9683);
nand UO_428 (O_428,N_9118,N_9537);
and UO_429 (O_429,N_9314,N_9554);
and UO_430 (O_430,N_9106,N_9884);
and UO_431 (O_431,N_9264,N_9190);
nand UO_432 (O_432,N_9894,N_9527);
nor UO_433 (O_433,N_9039,N_9916);
nor UO_434 (O_434,N_9316,N_9243);
nand UO_435 (O_435,N_9074,N_9637);
nor UO_436 (O_436,N_9260,N_9655);
and UO_437 (O_437,N_9684,N_9791);
nor UO_438 (O_438,N_9597,N_9354);
nand UO_439 (O_439,N_9293,N_9059);
nor UO_440 (O_440,N_9978,N_9890);
xnor UO_441 (O_441,N_9096,N_9598);
xor UO_442 (O_442,N_9919,N_9943);
and UO_443 (O_443,N_9173,N_9297);
or UO_444 (O_444,N_9705,N_9294);
nor UO_445 (O_445,N_9691,N_9075);
or UO_446 (O_446,N_9387,N_9005);
and UO_447 (O_447,N_9910,N_9710);
or UO_448 (O_448,N_9719,N_9725);
xnor UO_449 (O_449,N_9848,N_9378);
or UO_450 (O_450,N_9224,N_9430);
nor UO_451 (O_451,N_9362,N_9680);
nand UO_452 (O_452,N_9610,N_9529);
nand UO_453 (O_453,N_9025,N_9301);
nand UO_454 (O_454,N_9997,N_9205);
nor UO_455 (O_455,N_9974,N_9736);
nand UO_456 (O_456,N_9483,N_9101);
and UO_457 (O_457,N_9277,N_9840);
nand UO_458 (O_458,N_9034,N_9822);
nand UO_459 (O_459,N_9275,N_9787);
nor UO_460 (O_460,N_9508,N_9097);
nand UO_461 (O_461,N_9174,N_9594);
or UO_462 (O_462,N_9261,N_9517);
nand UO_463 (O_463,N_9171,N_9344);
nand UO_464 (O_464,N_9849,N_9368);
nand UO_465 (O_465,N_9909,N_9716);
or UO_466 (O_466,N_9574,N_9712);
or UO_467 (O_467,N_9740,N_9272);
nor UO_468 (O_468,N_9187,N_9608);
nor UO_469 (O_469,N_9766,N_9487);
nand UO_470 (O_470,N_9633,N_9685);
nand UO_471 (O_471,N_9946,N_9042);
and UO_472 (O_472,N_9673,N_9962);
xnor UO_473 (O_473,N_9244,N_9182);
nand UO_474 (O_474,N_9779,N_9306);
or UO_475 (O_475,N_9957,N_9697);
and UO_476 (O_476,N_9841,N_9765);
nor UO_477 (O_477,N_9854,N_9280);
nand UO_478 (O_478,N_9199,N_9880);
nor UO_479 (O_479,N_9958,N_9207);
or UO_480 (O_480,N_9078,N_9886);
and UO_481 (O_481,N_9286,N_9599);
and UO_482 (O_482,N_9105,N_9327);
nand UO_483 (O_483,N_9564,N_9968);
nor UO_484 (O_484,N_9735,N_9076);
nor UO_485 (O_485,N_9245,N_9175);
or UO_486 (O_486,N_9977,N_9416);
and UO_487 (O_487,N_9893,N_9123);
nand UO_488 (O_488,N_9953,N_9348);
nor UO_489 (O_489,N_9983,N_9334);
nand UO_490 (O_490,N_9163,N_9472);
nand UO_491 (O_491,N_9839,N_9147);
or UO_492 (O_492,N_9715,N_9700);
or UO_493 (O_493,N_9335,N_9846);
nor UO_494 (O_494,N_9852,N_9488);
or UO_495 (O_495,N_9394,N_9820);
nand UO_496 (O_496,N_9228,N_9579);
nand UO_497 (O_497,N_9409,N_9802);
and UO_498 (O_498,N_9024,N_9514);
nor UO_499 (O_499,N_9325,N_9158);
nor UO_500 (O_500,N_9039,N_9844);
nand UO_501 (O_501,N_9461,N_9757);
nand UO_502 (O_502,N_9943,N_9318);
nand UO_503 (O_503,N_9246,N_9414);
and UO_504 (O_504,N_9969,N_9028);
nand UO_505 (O_505,N_9390,N_9316);
nor UO_506 (O_506,N_9118,N_9631);
and UO_507 (O_507,N_9955,N_9755);
nand UO_508 (O_508,N_9991,N_9081);
nor UO_509 (O_509,N_9614,N_9599);
nand UO_510 (O_510,N_9344,N_9767);
or UO_511 (O_511,N_9936,N_9140);
or UO_512 (O_512,N_9607,N_9015);
nor UO_513 (O_513,N_9962,N_9108);
or UO_514 (O_514,N_9796,N_9986);
and UO_515 (O_515,N_9302,N_9459);
nor UO_516 (O_516,N_9920,N_9588);
nor UO_517 (O_517,N_9362,N_9457);
or UO_518 (O_518,N_9266,N_9555);
or UO_519 (O_519,N_9519,N_9571);
nor UO_520 (O_520,N_9011,N_9122);
nand UO_521 (O_521,N_9886,N_9141);
nand UO_522 (O_522,N_9747,N_9175);
nor UO_523 (O_523,N_9873,N_9574);
nor UO_524 (O_524,N_9267,N_9746);
and UO_525 (O_525,N_9687,N_9860);
and UO_526 (O_526,N_9213,N_9222);
and UO_527 (O_527,N_9384,N_9941);
or UO_528 (O_528,N_9706,N_9497);
or UO_529 (O_529,N_9418,N_9416);
and UO_530 (O_530,N_9037,N_9489);
nand UO_531 (O_531,N_9795,N_9843);
nor UO_532 (O_532,N_9954,N_9769);
xnor UO_533 (O_533,N_9503,N_9016);
nand UO_534 (O_534,N_9227,N_9988);
nand UO_535 (O_535,N_9824,N_9728);
nor UO_536 (O_536,N_9075,N_9014);
nand UO_537 (O_537,N_9894,N_9515);
and UO_538 (O_538,N_9350,N_9998);
nand UO_539 (O_539,N_9453,N_9224);
nor UO_540 (O_540,N_9073,N_9185);
nand UO_541 (O_541,N_9130,N_9404);
and UO_542 (O_542,N_9329,N_9503);
nor UO_543 (O_543,N_9914,N_9703);
nand UO_544 (O_544,N_9168,N_9812);
or UO_545 (O_545,N_9646,N_9516);
and UO_546 (O_546,N_9590,N_9347);
nand UO_547 (O_547,N_9624,N_9307);
or UO_548 (O_548,N_9962,N_9425);
nor UO_549 (O_549,N_9585,N_9293);
nor UO_550 (O_550,N_9821,N_9688);
and UO_551 (O_551,N_9308,N_9447);
or UO_552 (O_552,N_9765,N_9378);
nand UO_553 (O_553,N_9948,N_9868);
or UO_554 (O_554,N_9657,N_9498);
and UO_555 (O_555,N_9706,N_9816);
nor UO_556 (O_556,N_9968,N_9018);
nor UO_557 (O_557,N_9328,N_9978);
and UO_558 (O_558,N_9800,N_9351);
nor UO_559 (O_559,N_9802,N_9064);
nor UO_560 (O_560,N_9872,N_9339);
and UO_561 (O_561,N_9308,N_9467);
and UO_562 (O_562,N_9861,N_9269);
nor UO_563 (O_563,N_9808,N_9091);
nor UO_564 (O_564,N_9247,N_9360);
and UO_565 (O_565,N_9017,N_9320);
nand UO_566 (O_566,N_9010,N_9728);
or UO_567 (O_567,N_9673,N_9575);
nor UO_568 (O_568,N_9082,N_9690);
nor UO_569 (O_569,N_9212,N_9976);
nand UO_570 (O_570,N_9045,N_9387);
nand UO_571 (O_571,N_9910,N_9807);
nand UO_572 (O_572,N_9292,N_9701);
nand UO_573 (O_573,N_9818,N_9118);
nand UO_574 (O_574,N_9704,N_9618);
or UO_575 (O_575,N_9141,N_9178);
nand UO_576 (O_576,N_9544,N_9446);
or UO_577 (O_577,N_9461,N_9947);
nand UO_578 (O_578,N_9752,N_9556);
or UO_579 (O_579,N_9753,N_9082);
nor UO_580 (O_580,N_9098,N_9121);
nor UO_581 (O_581,N_9593,N_9909);
nand UO_582 (O_582,N_9683,N_9707);
or UO_583 (O_583,N_9970,N_9734);
or UO_584 (O_584,N_9292,N_9576);
nand UO_585 (O_585,N_9339,N_9831);
xnor UO_586 (O_586,N_9319,N_9823);
and UO_587 (O_587,N_9288,N_9403);
and UO_588 (O_588,N_9894,N_9606);
and UO_589 (O_589,N_9583,N_9693);
or UO_590 (O_590,N_9401,N_9237);
nor UO_591 (O_591,N_9227,N_9200);
nand UO_592 (O_592,N_9242,N_9130);
and UO_593 (O_593,N_9891,N_9054);
xor UO_594 (O_594,N_9187,N_9217);
nor UO_595 (O_595,N_9123,N_9027);
nand UO_596 (O_596,N_9213,N_9503);
nand UO_597 (O_597,N_9416,N_9733);
or UO_598 (O_598,N_9980,N_9974);
nor UO_599 (O_599,N_9827,N_9833);
nand UO_600 (O_600,N_9878,N_9097);
nand UO_601 (O_601,N_9994,N_9100);
nor UO_602 (O_602,N_9896,N_9018);
or UO_603 (O_603,N_9475,N_9823);
or UO_604 (O_604,N_9406,N_9411);
nand UO_605 (O_605,N_9683,N_9007);
nand UO_606 (O_606,N_9026,N_9410);
and UO_607 (O_607,N_9842,N_9945);
nand UO_608 (O_608,N_9407,N_9175);
nand UO_609 (O_609,N_9684,N_9194);
nor UO_610 (O_610,N_9455,N_9096);
or UO_611 (O_611,N_9167,N_9539);
nand UO_612 (O_612,N_9245,N_9789);
and UO_613 (O_613,N_9217,N_9874);
or UO_614 (O_614,N_9612,N_9326);
and UO_615 (O_615,N_9447,N_9809);
nor UO_616 (O_616,N_9851,N_9987);
nor UO_617 (O_617,N_9709,N_9970);
nand UO_618 (O_618,N_9793,N_9400);
or UO_619 (O_619,N_9867,N_9724);
nor UO_620 (O_620,N_9614,N_9513);
and UO_621 (O_621,N_9735,N_9266);
nor UO_622 (O_622,N_9577,N_9282);
and UO_623 (O_623,N_9730,N_9975);
nor UO_624 (O_624,N_9921,N_9154);
nor UO_625 (O_625,N_9308,N_9584);
nand UO_626 (O_626,N_9363,N_9111);
nand UO_627 (O_627,N_9663,N_9564);
nor UO_628 (O_628,N_9938,N_9834);
or UO_629 (O_629,N_9556,N_9376);
nand UO_630 (O_630,N_9482,N_9266);
nor UO_631 (O_631,N_9130,N_9223);
or UO_632 (O_632,N_9300,N_9940);
nor UO_633 (O_633,N_9259,N_9596);
or UO_634 (O_634,N_9315,N_9063);
and UO_635 (O_635,N_9747,N_9485);
or UO_636 (O_636,N_9537,N_9535);
nand UO_637 (O_637,N_9882,N_9960);
nor UO_638 (O_638,N_9346,N_9215);
nor UO_639 (O_639,N_9229,N_9415);
or UO_640 (O_640,N_9320,N_9677);
nor UO_641 (O_641,N_9909,N_9267);
or UO_642 (O_642,N_9787,N_9806);
or UO_643 (O_643,N_9798,N_9261);
nor UO_644 (O_644,N_9086,N_9921);
nor UO_645 (O_645,N_9036,N_9944);
and UO_646 (O_646,N_9327,N_9548);
or UO_647 (O_647,N_9118,N_9942);
nor UO_648 (O_648,N_9327,N_9907);
nand UO_649 (O_649,N_9812,N_9704);
and UO_650 (O_650,N_9376,N_9090);
nand UO_651 (O_651,N_9364,N_9884);
or UO_652 (O_652,N_9803,N_9342);
nor UO_653 (O_653,N_9767,N_9722);
or UO_654 (O_654,N_9172,N_9895);
nor UO_655 (O_655,N_9093,N_9060);
nand UO_656 (O_656,N_9639,N_9306);
nand UO_657 (O_657,N_9854,N_9799);
nor UO_658 (O_658,N_9586,N_9951);
or UO_659 (O_659,N_9670,N_9772);
and UO_660 (O_660,N_9899,N_9759);
nor UO_661 (O_661,N_9333,N_9631);
and UO_662 (O_662,N_9827,N_9768);
nand UO_663 (O_663,N_9377,N_9392);
nor UO_664 (O_664,N_9660,N_9007);
or UO_665 (O_665,N_9833,N_9034);
nor UO_666 (O_666,N_9236,N_9776);
or UO_667 (O_667,N_9136,N_9485);
or UO_668 (O_668,N_9044,N_9006);
nand UO_669 (O_669,N_9107,N_9439);
and UO_670 (O_670,N_9738,N_9406);
nor UO_671 (O_671,N_9122,N_9927);
and UO_672 (O_672,N_9641,N_9028);
and UO_673 (O_673,N_9743,N_9911);
and UO_674 (O_674,N_9905,N_9877);
nand UO_675 (O_675,N_9239,N_9546);
nand UO_676 (O_676,N_9047,N_9871);
and UO_677 (O_677,N_9104,N_9721);
and UO_678 (O_678,N_9364,N_9679);
or UO_679 (O_679,N_9363,N_9596);
or UO_680 (O_680,N_9210,N_9998);
and UO_681 (O_681,N_9801,N_9778);
or UO_682 (O_682,N_9077,N_9541);
xor UO_683 (O_683,N_9842,N_9889);
nor UO_684 (O_684,N_9620,N_9142);
and UO_685 (O_685,N_9656,N_9617);
nor UO_686 (O_686,N_9144,N_9873);
nor UO_687 (O_687,N_9136,N_9421);
nor UO_688 (O_688,N_9471,N_9392);
or UO_689 (O_689,N_9264,N_9181);
nor UO_690 (O_690,N_9837,N_9364);
and UO_691 (O_691,N_9326,N_9749);
and UO_692 (O_692,N_9495,N_9564);
nor UO_693 (O_693,N_9714,N_9414);
nor UO_694 (O_694,N_9367,N_9385);
and UO_695 (O_695,N_9885,N_9224);
and UO_696 (O_696,N_9656,N_9355);
or UO_697 (O_697,N_9024,N_9169);
or UO_698 (O_698,N_9888,N_9738);
and UO_699 (O_699,N_9753,N_9503);
xnor UO_700 (O_700,N_9004,N_9575);
and UO_701 (O_701,N_9176,N_9810);
and UO_702 (O_702,N_9433,N_9679);
or UO_703 (O_703,N_9393,N_9570);
or UO_704 (O_704,N_9287,N_9390);
or UO_705 (O_705,N_9021,N_9266);
nor UO_706 (O_706,N_9293,N_9368);
nand UO_707 (O_707,N_9434,N_9272);
nand UO_708 (O_708,N_9782,N_9640);
and UO_709 (O_709,N_9169,N_9293);
nor UO_710 (O_710,N_9204,N_9022);
and UO_711 (O_711,N_9907,N_9919);
nand UO_712 (O_712,N_9205,N_9602);
and UO_713 (O_713,N_9850,N_9010);
and UO_714 (O_714,N_9896,N_9526);
nor UO_715 (O_715,N_9846,N_9002);
nor UO_716 (O_716,N_9493,N_9677);
and UO_717 (O_717,N_9841,N_9626);
and UO_718 (O_718,N_9172,N_9676);
nor UO_719 (O_719,N_9768,N_9817);
nor UO_720 (O_720,N_9412,N_9655);
and UO_721 (O_721,N_9914,N_9155);
nand UO_722 (O_722,N_9244,N_9218);
nand UO_723 (O_723,N_9511,N_9976);
or UO_724 (O_724,N_9574,N_9577);
nor UO_725 (O_725,N_9481,N_9378);
nand UO_726 (O_726,N_9285,N_9377);
or UO_727 (O_727,N_9697,N_9943);
nand UO_728 (O_728,N_9780,N_9834);
and UO_729 (O_729,N_9664,N_9688);
nand UO_730 (O_730,N_9660,N_9820);
and UO_731 (O_731,N_9144,N_9966);
or UO_732 (O_732,N_9355,N_9713);
nand UO_733 (O_733,N_9186,N_9142);
or UO_734 (O_734,N_9385,N_9400);
nor UO_735 (O_735,N_9580,N_9775);
nor UO_736 (O_736,N_9256,N_9979);
nor UO_737 (O_737,N_9955,N_9170);
nand UO_738 (O_738,N_9649,N_9928);
nand UO_739 (O_739,N_9066,N_9593);
and UO_740 (O_740,N_9662,N_9039);
and UO_741 (O_741,N_9576,N_9816);
nand UO_742 (O_742,N_9363,N_9792);
nor UO_743 (O_743,N_9977,N_9370);
and UO_744 (O_744,N_9507,N_9737);
nand UO_745 (O_745,N_9975,N_9448);
or UO_746 (O_746,N_9965,N_9103);
and UO_747 (O_747,N_9338,N_9162);
nand UO_748 (O_748,N_9379,N_9785);
nand UO_749 (O_749,N_9310,N_9794);
and UO_750 (O_750,N_9824,N_9109);
nor UO_751 (O_751,N_9159,N_9002);
or UO_752 (O_752,N_9322,N_9908);
and UO_753 (O_753,N_9040,N_9930);
or UO_754 (O_754,N_9141,N_9953);
nand UO_755 (O_755,N_9541,N_9578);
nor UO_756 (O_756,N_9938,N_9080);
nor UO_757 (O_757,N_9471,N_9686);
and UO_758 (O_758,N_9870,N_9957);
nor UO_759 (O_759,N_9672,N_9883);
nor UO_760 (O_760,N_9605,N_9755);
nor UO_761 (O_761,N_9700,N_9264);
or UO_762 (O_762,N_9044,N_9463);
and UO_763 (O_763,N_9501,N_9868);
nor UO_764 (O_764,N_9892,N_9518);
nor UO_765 (O_765,N_9667,N_9010);
or UO_766 (O_766,N_9382,N_9860);
and UO_767 (O_767,N_9204,N_9823);
and UO_768 (O_768,N_9471,N_9331);
nor UO_769 (O_769,N_9936,N_9143);
or UO_770 (O_770,N_9859,N_9572);
and UO_771 (O_771,N_9304,N_9347);
nand UO_772 (O_772,N_9367,N_9549);
nand UO_773 (O_773,N_9319,N_9119);
or UO_774 (O_774,N_9812,N_9926);
or UO_775 (O_775,N_9974,N_9234);
and UO_776 (O_776,N_9121,N_9633);
and UO_777 (O_777,N_9513,N_9713);
or UO_778 (O_778,N_9392,N_9213);
nand UO_779 (O_779,N_9246,N_9766);
nor UO_780 (O_780,N_9162,N_9017);
or UO_781 (O_781,N_9483,N_9428);
or UO_782 (O_782,N_9698,N_9872);
or UO_783 (O_783,N_9162,N_9738);
nor UO_784 (O_784,N_9851,N_9319);
nand UO_785 (O_785,N_9437,N_9876);
xor UO_786 (O_786,N_9295,N_9776);
and UO_787 (O_787,N_9926,N_9798);
or UO_788 (O_788,N_9027,N_9060);
nand UO_789 (O_789,N_9900,N_9621);
or UO_790 (O_790,N_9473,N_9573);
nand UO_791 (O_791,N_9849,N_9113);
or UO_792 (O_792,N_9667,N_9953);
and UO_793 (O_793,N_9874,N_9046);
nand UO_794 (O_794,N_9835,N_9624);
and UO_795 (O_795,N_9951,N_9422);
and UO_796 (O_796,N_9336,N_9257);
nor UO_797 (O_797,N_9522,N_9132);
and UO_798 (O_798,N_9973,N_9249);
nor UO_799 (O_799,N_9427,N_9043);
nand UO_800 (O_800,N_9378,N_9836);
or UO_801 (O_801,N_9465,N_9472);
and UO_802 (O_802,N_9656,N_9665);
or UO_803 (O_803,N_9180,N_9800);
or UO_804 (O_804,N_9430,N_9102);
nor UO_805 (O_805,N_9748,N_9059);
nor UO_806 (O_806,N_9580,N_9503);
nand UO_807 (O_807,N_9172,N_9529);
or UO_808 (O_808,N_9525,N_9519);
nand UO_809 (O_809,N_9709,N_9134);
or UO_810 (O_810,N_9739,N_9359);
and UO_811 (O_811,N_9053,N_9839);
and UO_812 (O_812,N_9336,N_9176);
nand UO_813 (O_813,N_9534,N_9163);
nor UO_814 (O_814,N_9970,N_9342);
nand UO_815 (O_815,N_9513,N_9702);
nand UO_816 (O_816,N_9330,N_9644);
or UO_817 (O_817,N_9506,N_9999);
or UO_818 (O_818,N_9388,N_9331);
nand UO_819 (O_819,N_9423,N_9715);
nor UO_820 (O_820,N_9148,N_9793);
or UO_821 (O_821,N_9400,N_9743);
nor UO_822 (O_822,N_9995,N_9715);
or UO_823 (O_823,N_9297,N_9990);
nor UO_824 (O_824,N_9740,N_9422);
xnor UO_825 (O_825,N_9123,N_9283);
nand UO_826 (O_826,N_9477,N_9252);
nor UO_827 (O_827,N_9748,N_9110);
or UO_828 (O_828,N_9251,N_9500);
nand UO_829 (O_829,N_9892,N_9217);
or UO_830 (O_830,N_9591,N_9041);
nand UO_831 (O_831,N_9868,N_9076);
or UO_832 (O_832,N_9208,N_9241);
and UO_833 (O_833,N_9030,N_9888);
or UO_834 (O_834,N_9122,N_9616);
and UO_835 (O_835,N_9285,N_9599);
and UO_836 (O_836,N_9304,N_9267);
or UO_837 (O_837,N_9168,N_9427);
nand UO_838 (O_838,N_9839,N_9133);
or UO_839 (O_839,N_9700,N_9677);
nor UO_840 (O_840,N_9094,N_9670);
and UO_841 (O_841,N_9778,N_9137);
nand UO_842 (O_842,N_9937,N_9629);
nor UO_843 (O_843,N_9615,N_9131);
nand UO_844 (O_844,N_9886,N_9233);
and UO_845 (O_845,N_9188,N_9091);
nand UO_846 (O_846,N_9075,N_9817);
or UO_847 (O_847,N_9396,N_9559);
or UO_848 (O_848,N_9500,N_9524);
nand UO_849 (O_849,N_9291,N_9741);
nor UO_850 (O_850,N_9362,N_9330);
or UO_851 (O_851,N_9690,N_9835);
and UO_852 (O_852,N_9368,N_9760);
and UO_853 (O_853,N_9577,N_9814);
nor UO_854 (O_854,N_9975,N_9745);
and UO_855 (O_855,N_9298,N_9640);
nor UO_856 (O_856,N_9134,N_9285);
and UO_857 (O_857,N_9971,N_9503);
or UO_858 (O_858,N_9320,N_9780);
or UO_859 (O_859,N_9994,N_9977);
nand UO_860 (O_860,N_9235,N_9319);
nand UO_861 (O_861,N_9473,N_9312);
and UO_862 (O_862,N_9076,N_9704);
or UO_863 (O_863,N_9552,N_9714);
nand UO_864 (O_864,N_9733,N_9920);
nand UO_865 (O_865,N_9820,N_9726);
nand UO_866 (O_866,N_9997,N_9326);
nor UO_867 (O_867,N_9433,N_9766);
nor UO_868 (O_868,N_9243,N_9963);
or UO_869 (O_869,N_9805,N_9211);
or UO_870 (O_870,N_9739,N_9883);
and UO_871 (O_871,N_9416,N_9057);
and UO_872 (O_872,N_9328,N_9469);
nor UO_873 (O_873,N_9158,N_9935);
or UO_874 (O_874,N_9081,N_9147);
and UO_875 (O_875,N_9234,N_9039);
nand UO_876 (O_876,N_9461,N_9466);
nand UO_877 (O_877,N_9623,N_9754);
and UO_878 (O_878,N_9363,N_9659);
and UO_879 (O_879,N_9387,N_9493);
and UO_880 (O_880,N_9419,N_9200);
nand UO_881 (O_881,N_9160,N_9065);
or UO_882 (O_882,N_9601,N_9073);
nand UO_883 (O_883,N_9428,N_9891);
nand UO_884 (O_884,N_9468,N_9616);
nand UO_885 (O_885,N_9691,N_9148);
nand UO_886 (O_886,N_9791,N_9288);
nand UO_887 (O_887,N_9372,N_9685);
or UO_888 (O_888,N_9690,N_9681);
and UO_889 (O_889,N_9634,N_9113);
nand UO_890 (O_890,N_9589,N_9635);
or UO_891 (O_891,N_9960,N_9872);
nor UO_892 (O_892,N_9304,N_9121);
and UO_893 (O_893,N_9168,N_9809);
nor UO_894 (O_894,N_9273,N_9101);
or UO_895 (O_895,N_9717,N_9551);
nor UO_896 (O_896,N_9197,N_9811);
and UO_897 (O_897,N_9488,N_9791);
nand UO_898 (O_898,N_9312,N_9842);
nor UO_899 (O_899,N_9287,N_9406);
nor UO_900 (O_900,N_9372,N_9578);
or UO_901 (O_901,N_9457,N_9706);
and UO_902 (O_902,N_9385,N_9981);
and UO_903 (O_903,N_9895,N_9287);
nand UO_904 (O_904,N_9199,N_9200);
nor UO_905 (O_905,N_9072,N_9472);
or UO_906 (O_906,N_9076,N_9685);
nand UO_907 (O_907,N_9518,N_9261);
or UO_908 (O_908,N_9027,N_9959);
nor UO_909 (O_909,N_9861,N_9070);
or UO_910 (O_910,N_9456,N_9437);
or UO_911 (O_911,N_9686,N_9701);
nor UO_912 (O_912,N_9861,N_9766);
or UO_913 (O_913,N_9079,N_9220);
and UO_914 (O_914,N_9575,N_9298);
or UO_915 (O_915,N_9837,N_9980);
nand UO_916 (O_916,N_9176,N_9760);
or UO_917 (O_917,N_9545,N_9158);
nand UO_918 (O_918,N_9194,N_9143);
nor UO_919 (O_919,N_9761,N_9090);
and UO_920 (O_920,N_9646,N_9503);
and UO_921 (O_921,N_9574,N_9023);
nand UO_922 (O_922,N_9985,N_9126);
and UO_923 (O_923,N_9585,N_9370);
nand UO_924 (O_924,N_9534,N_9222);
and UO_925 (O_925,N_9978,N_9733);
nand UO_926 (O_926,N_9920,N_9229);
nand UO_927 (O_927,N_9976,N_9844);
nor UO_928 (O_928,N_9912,N_9315);
nor UO_929 (O_929,N_9877,N_9164);
nand UO_930 (O_930,N_9840,N_9285);
nand UO_931 (O_931,N_9216,N_9754);
nor UO_932 (O_932,N_9786,N_9199);
nor UO_933 (O_933,N_9088,N_9655);
nand UO_934 (O_934,N_9505,N_9640);
nor UO_935 (O_935,N_9763,N_9203);
nor UO_936 (O_936,N_9172,N_9137);
or UO_937 (O_937,N_9140,N_9255);
or UO_938 (O_938,N_9476,N_9589);
or UO_939 (O_939,N_9626,N_9649);
nor UO_940 (O_940,N_9893,N_9311);
or UO_941 (O_941,N_9187,N_9142);
or UO_942 (O_942,N_9762,N_9709);
and UO_943 (O_943,N_9469,N_9591);
nor UO_944 (O_944,N_9749,N_9793);
nor UO_945 (O_945,N_9557,N_9967);
or UO_946 (O_946,N_9168,N_9788);
nand UO_947 (O_947,N_9717,N_9454);
nand UO_948 (O_948,N_9402,N_9583);
nand UO_949 (O_949,N_9795,N_9390);
xor UO_950 (O_950,N_9283,N_9728);
nor UO_951 (O_951,N_9782,N_9005);
nand UO_952 (O_952,N_9892,N_9977);
nand UO_953 (O_953,N_9400,N_9628);
or UO_954 (O_954,N_9519,N_9147);
nor UO_955 (O_955,N_9093,N_9946);
xnor UO_956 (O_956,N_9208,N_9419);
or UO_957 (O_957,N_9054,N_9043);
or UO_958 (O_958,N_9552,N_9623);
nor UO_959 (O_959,N_9224,N_9150);
and UO_960 (O_960,N_9059,N_9377);
and UO_961 (O_961,N_9964,N_9370);
nand UO_962 (O_962,N_9512,N_9060);
or UO_963 (O_963,N_9225,N_9777);
nor UO_964 (O_964,N_9576,N_9934);
nand UO_965 (O_965,N_9839,N_9007);
nand UO_966 (O_966,N_9150,N_9223);
nand UO_967 (O_967,N_9298,N_9104);
or UO_968 (O_968,N_9980,N_9014);
nand UO_969 (O_969,N_9049,N_9489);
or UO_970 (O_970,N_9667,N_9269);
or UO_971 (O_971,N_9878,N_9210);
and UO_972 (O_972,N_9408,N_9410);
nand UO_973 (O_973,N_9848,N_9717);
nand UO_974 (O_974,N_9237,N_9671);
and UO_975 (O_975,N_9565,N_9200);
nor UO_976 (O_976,N_9179,N_9625);
and UO_977 (O_977,N_9883,N_9977);
and UO_978 (O_978,N_9357,N_9793);
or UO_979 (O_979,N_9818,N_9392);
nor UO_980 (O_980,N_9372,N_9199);
nor UO_981 (O_981,N_9435,N_9573);
and UO_982 (O_982,N_9671,N_9494);
nand UO_983 (O_983,N_9147,N_9824);
and UO_984 (O_984,N_9830,N_9679);
and UO_985 (O_985,N_9781,N_9469);
and UO_986 (O_986,N_9784,N_9534);
nor UO_987 (O_987,N_9907,N_9943);
nor UO_988 (O_988,N_9157,N_9680);
or UO_989 (O_989,N_9663,N_9271);
or UO_990 (O_990,N_9360,N_9237);
xor UO_991 (O_991,N_9247,N_9216);
or UO_992 (O_992,N_9617,N_9863);
and UO_993 (O_993,N_9406,N_9383);
and UO_994 (O_994,N_9365,N_9560);
or UO_995 (O_995,N_9438,N_9037);
nand UO_996 (O_996,N_9458,N_9423);
and UO_997 (O_997,N_9382,N_9704);
nor UO_998 (O_998,N_9471,N_9234);
nor UO_999 (O_999,N_9916,N_9976);
nor UO_1000 (O_1000,N_9277,N_9068);
nor UO_1001 (O_1001,N_9727,N_9378);
and UO_1002 (O_1002,N_9061,N_9134);
nor UO_1003 (O_1003,N_9565,N_9047);
nand UO_1004 (O_1004,N_9900,N_9441);
nand UO_1005 (O_1005,N_9827,N_9851);
and UO_1006 (O_1006,N_9220,N_9188);
and UO_1007 (O_1007,N_9978,N_9996);
nor UO_1008 (O_1008,N_9105,N_9793);
and UO_1009 (O_1009,N_9141,N_9749);
and UO_1010 (O_1010,N_9931,N_9092);
nor UO_1011 (O_1011,N_9081,N_9537);
and UO_1012 (O_1012,N_9466,N_9627);
and UO_1013 (O_1013,N_9234,N_9141);
nor UO_1014 (O_1014,N_9670,N_9689);
or UO_1015 (O_1015,N_9947,N_9283);
nor UO_1016 (O_1016,N_9628,N_9908);
and UO_1017 (O_1017,N_9848,N_9183);
nor UO_1018 (O_1018,N_9685,N_9968);
and UO_1019 (O_1019,N_9771,N_9270);
nand UO_1020 (O_1020,N_9988,N_9778);
or UO_1021 (O_1021,N_9085,N_9357);
nand UO_1022 (O_1022,N_9691,N_9568);
or UO_1023 (O_1023,N_9141,N_9622);
nor UO_1024 (O_1024,N_9113,N_9782);
nand UO_1025 (O_1025,N_9041,N_9723);
and UO_1026 (O_1026,N_9046,N_9310);
or UO_1027 (O_1027,N_9235,N_9586);
and UO_1028 (O_1028,N_9579,N_9201);
nor UO_1029 (O_1029,N_9892,N_9955);
or UO_1030 (O_1030,N_9695,N_9194);
and UO_1031 (O_1031,N_9893,N_9809);
nand UO_1032 (O_1032,N_9074,N_9187);
nand UO_1033 (O_1033,N_9566,N_9191);
nand UO_1034 (O_1034,N_9339,N_9928);
and UO_1035 (O_1035,N_9195,N_9942);
or UO_1036 (O_1036,N_9298,N_9509);
and UO_1037 (O_1037,N_9526,N_9061);
nor UO_1038 (O_1038,N_9140,N_9350);
and UO_1039 (O_1039,N_9688,N_9592);
or UO_1040 (O_1040,N_9461,N_9033);
nor UO_1041 (O_1041,N_9183,N_9095);
and UO_1042 (O_1042,N_9217,N_9124);
nand UO_1043 (O_1043,N_9199,N_9339);
nor UO_1044 (O_1044,N_9172,N_9581);
nor UO_1045 (O_1045,N_9804,N_9887);
nor UO_1046 (O_1046,N_9010,N_9362);
and UO_1047 (O_1047,N_9790,N_9504);
or UO_1048 (O_1048,N_9562,N_9671);
nor UO_1049 (O_1049,N_9647,N_9030);
and UO_1050 (O_1050,N_9526,N_9396);
or UO_1051 (O_1051,N_9763,N_9014);
or UO_1052 (O_1052,N_9092,N_9867);
nor UO_1053 (O_1053,N_9061,N_9850);
and UO_1054 (O_1054,N_9916,N_9256);
nor UO_1055 (O_1055,N_9212,N_9814);
or UO_1056 (O_1056,N_9153,N_9521);
nor UO_1057 (O_1057,N_9001,N_9696);
nand UO_1058 (O_1058,N_9908,N_9914);
nor UO_1059 (O_1059,N_9044,N_9254);
nand UO_1060 (O_1060,N_9099,N_9160);
nand UO_1061 (O_1061,N_9575,N_9846);
nand UO_1062 (O_1062,N_9753,N_9832);
nand UO_1063 (O_1063,N_9943,N_9544);
nor UO_1064 (O_1064,N_9408,N_9777);
nand UO_1065 (O_1065,N_9150,N_9795);
nor UO_1066 (O_1066,N_9749,N_9766);
nand UO_1067 (O_1067,N_9012,N_9104);
nand UO_1068 (O_1068,N_9183,N_9708);
nor UO_1069 (O_1069,N_9115,N_9749);
nor UO_1070 (O_1070,N_9644,N_9654);
nand UO_1071 (O_1071,N_9264,N_9940);
or UO_1072 (O_1072,N_9795,N_9439);
or UO_1073 (O_1073,N_9604,N_9193);
and UO_1074 (O_1074,N_9377,N_9526);
nor UO_1075 (O_1075,N_9005,N_9473);
and UO_1076 (O_1076,N_9600,N_9031);
or UO_1077 (O_1077,N_9047,N_9279);
nand UO_1078 (O_1078,N_9943,N_9866);
or UO_1079 (O_1079,N_9243,N_9988);
nand UO_1080 (O_1080,N_9183,N_9280);
nor UO_1081 (O_1081,N_9348,N_9075);
and UO_1082 (O_1082,N_9821,N_9714);
or UO_1083 (O_1083,N_9971,N_9729);
nor UO_1084 (O_1084,N_9367,N_9137);
xnor UO_1085 (O_1085,N_9609,N_9687);
or UO_1086 (O_1086,N_9294,N_9034);
xnor UO_1087 (O_1087,N_9656,N_9381);
nand UO_1088 (O_1088,N_9129,N_9955);
or UO_1089 (O_1089,N_9821,N_9120);
and UO_1090 (O_1090,N_9541,N_9926);
nand UO_1091 (O_1091,N_9076,N_9845);
and UO_1092 (O_1092,N_9001,N_9570);
nor UO_1093 (O_1093,N_9766,N_9761);
nand UO_1094 (O_1094,N_9097,N_9010);
or UO_1095 (O_1095,N_9043,N_9585);
or UO_1096 (O_1096,N_9813,N_9038);
and UO_1097 (O_1097,N_9410,N_9447);
and UO_1098 (O_1098,N_9304,N_9981);
and UO_1099 (O_1099,N_9028,N_9633);
nand UO_1100 (O_1100,N_9923,N_9940);
and UO_1101 (O_1101,N_9907,N_9872);
nand UO_1102 (O_1102,N_9938,N_9619);
nand UO_1103 (O_1103,N_9860,N_9406);
nor UO_1104 (O_1104,N_9297,N_9122);
nor UO_1105 (O_1105,N_9059,N_9722);
xor UO_1106 (O_1106,N_9674,N_9510);
or UO_1107 (O_1107,N_9015,N_9517);
or UO_1108 (O_1108,N_9217,N_9108);
nand UO_1109 (O_1109,N_9935,N_9941);
xnor UO_1110 (O_1110,N_9191,N_9944);
or UO_1111 (O_1111,N_9042,N_9472);
and UO_1112 (O_1112,N_9332,N_9286);
and UO_1113 (O_1113,N_9992,N_9525);
and UO_1114 (O_1114,N_9299,N_9712);
nand UO_1115 (O_1115,N_9625,N_9161);
nand UO_1116 (O_1116,N_9766,N_9970);
and UO_1117 (O_1117,N_9771,N_9107);
nand UO_1118 (O_1118,N_9375,N_9007);
nor UO_1119 (O_1119,N_9499,N_9707);
or UO_1120 (O_1120,N_9848,N_9780);
nor UO_1121 (O_1121,N_9706,N_9440);
or UO_1122 (O_1122,N_9145,N_9402);
and UO_1123 (O_1123,N_9566,N_9765);
or UO_1124 (O_1124,N_9568,N_9989);
or UO_1125 (O_1125,N_9608,N_9010);
or UO_1126 (O_1126,N_9091,N_9813);
nand UO_1127 (O_1127,N_9595,N_9511);
or UO_1128 (O_1128,N_9044,N_9643);
and UO_1129 (O_1129,N_9127,N_9558);
and UO_1130 (O_1130,N_9467,N_9311);
or UO_1131 (O_1131,N_9162,N_9744);
and UO_1132 (O_1132,N_9563,N_9600);
or UO_1133 (O_1133,N_9239,N_9843);
and UO_1134 (O_1134,N_9877,N_9889);
and UO_1135 (O_1135,N_9455,N_9623);
nor UO_1136 (O_1136,N_9180,N_9267);
and UO_1137 (O_1137,N_9389,N_9170);
or UO_1138 (O_1138,N_9082,N_9699);
or UO_1139 (O_1139,N_9162,N_9532);
nor UO_1140 (O_1140,N_9866,N_9872);
and UO_1141 (O_1141,N_9245,N_9918);
and UO_1142 (O_1142,N_9322,N_9306);
and UO_1143 (O_1143,N_9686,N_9870);
or UO_1144 (O_1144,N_9488,N_9221);
nand UO_1145 (O_1145,N_9779,N_9398);
and UO_1146 (O_1146,N_9595,N_9637);
nor UO_1147 (O_1147,N_9358,N_9100);
xor UO_1148 (O_1148,N_9175,N_9189);
or UO_1149 (O_1149,N_9036,N_9750);
or UO_1150 (O_1150,N_9415,N_9351);
nand UO_1151 (O_1151,N_9303,N_9825);
nor UO_1152 (O_1152,N_9094,N_9472);
nor UO_1153 (O_1153,N_9399,N_9357);
nor UO_1154 (O_1154,N_9888,N_9808);
and UO_1155 (O_1155,N_9765,N_9657);
or UO_1156 (O_1156,N_9946,N_9468);
nand UO_1157 (O_1157,N_9509,N_9530);
nand UO_1158 (O_1158,N_9275,N_9778);
and UO_1159 (O_1159,N_9653,N_9045);
and UO_1160 (O_1160,N_9848,N_9316);
or UO_1161 (O_1161,N_9911,N_9549);
and UO_1162 (O_1162,N_9649,N_9127);
and UO_1163 (O_1163,N_9243,N_9856);
xnor UO_1164 (O_1164,N_9115,N_9198);
and UO_1165 (O_1165,N_9092,N_9066);
nor UO_1166 (O_1166,N_9633,N_9812);
and UO_1167 (O_1167,N_9941,N_9566);
or UO_1168 (O_1168,N_9163,N_9130);
nand UO_1169 (O_1169,N_9095,N_9442);
and UO_1170 (O_1170,N_9617,N_9639);
or UO_1171 (O_1171,N_9141,N_9954);
nand UO_1172 (O_1172,N_9975,N_9737);
nand UO_1173 (O_1173,N_9239,N_9972);
or UO_1174 (O_1174,N_9022,N_9836);
nand UO_1175 (O_1175,N_9947,N_9824);
nand UO_1176 (O_1176,N_9779,N_9404);
nor UO_1177 (O_1177,N_9044,N_9720);
or UO_1178 (O_1178,N_9772,N_9357);
nor UO_1179 (O_1179,N_9889,N_9316);
nor UO_1180 (O_1180,N_9924,N_9094);
nor UO_1181 (O_1181,N_9652,N_9388);
nand UO_1182 (O_1182,N_9127,N_9381);
and UO_1183 (O_1183,N_9186,N_9911);
nor UO_1184 (O_1184,N_9194,N_9391);
and UO_1185 (O_1185,N_9187,N_9178);
and UO_1186 (O_1186,N_9553,N_9311);
and UO_1187 (O_1187,N_9309,N_9150);
nor UO_1188 (O_1188,N_9661,N_9635);
or UO_1189 (O_1189,N_9817,N_9979);
nor UO_1190 (O_1190,N_9621,N_9542);
nand UO_1191 (O_1191,N_9600,N_9847);
nor UO_1192 (O_1192,N_9865,N_9409);
and UO_1193 (O_1193,N_9639,N_9528);
and UO_1194 (O_1194,N_9031,N_9487);
nand UO_1195 (O_1195,N_9609,N_9299);
nand UO_1196 (O_1196,N_9794,N_9398);
nand UO_1197 (O_1197,N_9285,N_9854);
or UO_1198 (O_1198,N_9831,N_9290);
nor UO_1199 (O_1199,N_9608,N_9216);
nand UO_1200 (O_1200,N_9024,N_9736);
nand UO_1201 (O_1201,N_9380,N_9233);
nand UO_1202 (O_1202,N_9530,N_9775);
and UO_1203 (O_1203,N_9177,N_9664);
or UO_1204 (O_1204,N_9400,N_9411);
or UO_1205 (O_1205,N_9528,N_9873);
nor UO_1206 (O_1206,N_9265,N_9047);
nand UO_1207 (O_1207,N_9692,N_9767);
nand UO_1208 (O_1208,N_9136,N_9275);
nor UO_1209 (O_1209,N_9398,N_9835);
nand UO_1210 (O_1210,N_9596,N_9197);
and UO_1211 (O_1211,N_9585,N_9382);
and UO_1212 (O_1212,N_9279,N_9176);
nor UO_1213 (O_1213,N_9072,N_9233);
and UO_1214 (O_1214,N_9132,N_9158);
and UO_1215 (O_1215,N_9686,N_9943);
nor UO_1216 (O_1216,N_9758,N_9508);
nand UO_1217 (O_1217,N_9320,N_9503);
or UO_1218 (O_1218,N_9221,N_9983);
and UO_1219 (O_1219,N_9030,N_9662);
nand UO_1220 (O_1220,N_9086,N_9865);
and UO_1221 (O_1221,N_9901,N_9921);
and UO_1222 (O_1222,N_9413,N_9912);
and UO_1223 (O_1223,N_9946,N_9395);
nor UO_1224 (O_1224,N_9998,N_9988);
nor UO_1225 (O_1225,N_9173,N_9292);
nor UO_1226 (O_1226,N_9484,N_9092);
and UO_1227 (O_1227,N_9575,N_9798);
and UO_1228 (O_1228,N_9224,N_9531);
or UO_1229 (O_1229,N_9558,N_9718);
nor UO_1230 (O_1230,N_9498,N_9169);
nor UO_1231 (O_1231,N_9803,N_9750);
and UO_1232 (O_1232,N_9075,N_9764);
or UO_1233 (O_1233,N_9093,N_9463);
or UO_1234 (O_1234,N_9583,N_9186);
and UO_1235 (O_1235,N_9082,N_9201);
and UO_1236 (O_1236,N_9932,N_9139);
nand UO_1237 (O_1237,N_9787,N_9790);
or UO_1238 (O_1238,N_9655,N_9326);
nor UO_1239 (O_1239,N_9575,N_9720);
and UO_1240 (O_1240,N_9600,N_9272);
nand UO_1241 (O_1241,N_9019,N_9248);
nand UO_1242 (O_1242,N_9773,N_9475);
nand UO_1243 (O_1243,N_9025,N_9060);
or UO_1244 (O_1244,N_9856,N_9094);
nor UO_1245 (O_1245,N_9691,N_9146);
nand UO_1246 (O_1246,N_9363,N_9724);
and UO_1247 (O_1247,N_9575,N_9333);
or UO_1248 (O_1248,N_9414,N_9241);
nor UO_1249 (O_1249,N_9181,N_9071);
and UO_1250 (O_1250,N_9365,N_9441);
nand UO_1251 (O_1251,N_9346,N_9944);
nand UO_1252 (O_1252,N_9112,N_9994);
nand UO_1253 (O_1253,N_9676,N_9373);
nor UO_1254 (O_1254,N_9680,N_9649);
nand UO_1255 (O_1255,N_9538,N_9176);
nor UO_1256 (O_1256,N_9550,N_9614);
nor UO_1257 (O_1257,N_9563,N_9735);
and UO_1258 (O_1258,N_9277,N_9805);
or UO_1259 (O_1259,N_9360,N_9458);
nor UO_1260 (O_1260,N_9113,N_9567);
or UO_1261 (O_1261,N_9767,N_9531);
or UO_1262 (O_1262,N_9175,N_9517);
nor UO_1263 (O_1263,N_9657,N_9832);
nor UO_1264 (O_1264,N_9758,N_9424);
nand UO_1265 (O_1265,N_9981,N_9059);
nor UO_1266 (O_1266,N_9735,N_9673);
or UO_1267 (O_1267,N_9577,N_9381);
nor UO_1268 (O_1268,N_9624,N_9033);
or UO_1269 (O_1269,N_9261,N_9940);
nand UO_1270 (O_1270,N_9547,N_9381);
nand UO_1271 (O_1271,N_9686,N_9066);
or UO_1272 (O_1272,N_9083,N_9360);
nand UO_1273 (O_1273,N_9738,N_9349);
and UO_1274 (O_1274,N_9077,N_9479);
nor UO_1275 (O_1275,N_9653,N_9565);
xnor UO_1276 (O_1276,N_9537,N_9479);
nor UO_1277 (O_1277,N_9790,N_9526);
nor UO_1278 (O_1278,N_9310,N_9934);
nor UO_1279 (O_1279,N_9362,N_9228);
nand UO_1280 (O_1280,N_9354,N_9826);
xor UO_1281 (O_1281,N_9333,N_9630);
nor UO_1282 (O_1282,N_9560,N_9669);
xor UO_1283 (O_1283,N_9813,N_9110);
or UO_1284 (O_1284,N_9535,N_9919);
and UO_1285 (O_1285,N_9808,N_9131);
or UO_1286 (O_1286,N_9905,N_9037);
nand UO_1287 (O_1287,N_9046,N_9568);
nand UO_1288 (O_1288,N_9542,N_9128);
and UO_1289 (O_1289,N_9581,N_9173);
and UO_1290 (O_1290,N_9868,N_9571);
and UO_1291 (O_1291,N_9344,N_9312);
nor UO_1292 (O_1292,N_9326,N_9356);
nand UO_1293 (O_1293,N_9585,N_9605);
nand UO_1294 (O_1294,N_9022,N_9635);
and UO_1295 (O_1295,N_9179,N_9082);
nor UO_1296 (O_1296,N_9839,N_9639);
nor UO_1297 (O_1297,N_9680,N_9286);
and UO_1298 (O_1298,N_9301,N_9164);
nor UO_1299 (O_1299,N_9385,N_9287);
or UO_1300 (O_1300,N_9753,N_9293);
and UO_1301 (O_1301,N_9831,N_9825);
or UO_1302 (O_1302,N_9522,N_9449);
nand UO_1303 (O_1303,N_9962,N_9584);
nand UO_1304 (O_1304,N_9866,N_9595);
nor UO_1305 (O_1305,N_9344,N_9291);
nand UO_1306 (O_1306,N_9008,N_9195);
and UO_1307 (O_1307,N_9125,N_9704);
and UO_1308 (O_1308,N_9351,N_9948);
nor UO_1309 (O_1309,N_9044,N_9519);
nand UO_1310 (O_1310,N_9172,N_9965);
nand UO_1311 (O_1311,N_9678,N_9141);
and UO_1312 (O_1312,N_9165,N_9552);
nand UO_1313 (O_1313,N_9795,N_9743);
nand UO_1314 (O_1314,N_9767,N_9519);
nand UO_1315 (O_1315,N_9059,N_9158);
or UO_1316 (O_1316,N_9051,N_9018);
xor UO_1317 (O_1317,N_9063,N_9501);
and UO_1318 (O_1318,N_9648,N_9216);
and UO_1319 (O_1319,N_9573,N_9922);
nand UO_1320 (O_1320,N_9892,N_9438);
nand UO_1321 (O_1321,N_9641,N_9709);
nand UO_1322 (O_1322,N_9520,N_9510);
or UO_1323 (O_1323,N_9821,N_9415);
nand UO_1324 (O_1324,N_9733,N_9743);
and UO_1325 (O_1325,N_9202,N_9189);
nand UO_1326 (O_1326,N_9823,N_9725);
nand UO_1327 (O_1327,N_9358,N_9120);
and UO_1328 (O_1328,N_9286,N_9267);
and UO_1329 (O_1329,N_9809,N_9137);
or UO_1330 (O_1330,N_9896,N_9086);
nand UO_1331 (O_1331,N_9216,N_9115);
and UO_1332 (O_1332,N_9372,N_9831);
or UO_1333 (O_1333,N_9365,N_9722);
nor UO_1334 (O_1334,N_9842,N_9322);
nor UO_1335 (O_1335,N_9027,N_9954);
nand UO_1336 (O_1336,N_9297,N_9032);
nand UO_1337 (O_1337,N_9363,N_9133);
and UO_1338 (O_1338,N_9417,N_9717);
nand UO_1339 (O_1339,N_9395,N_9818);
nor UO_1340 (O_1340,N_9309,N_9910);
and UO_1341 (O_1341,N_9652,N_9872);
and UO_1342 (O_1342,N_9563,N_9453);
nor UO_1343 (O_1343,N_9510,N_9185);
nor UO_1344 (O_1344,N_9537,N_9349);
nand UO_1345 (O_1345,N_9239,N_9952);
and UO_1346 (O_1346,N_9473,N_9427);
nor UO_1347 (O_1347,N_9385,N_9992);
or UO_1348 (O_1348,N_9223,N_9744);
nor UO_1349 (O_1349,N_9947,N_9660);
xnor UO_1350 (O_1350,N_9132,N_9285);
nor UO_1351 (O_1351,N_9116,N_9839);
nor UO_1352 (O_1352,N_9353,N_9301);
or UO_1353 (O_1353,N_9104,N_9269);
or UO_1354 (O_1354,N_9460,N_9954);
nand UO_1355 (O_1355,N_9430,N_9388);
and UO_1356 (O_1356,N_9804,N_9412);
nor UO_1357 (O_1357,N_9398,N_9564);
nor UO_1358 (O_1358,N_9127,N_9082);
nor UO_1359 (O_1359,N_9685,N_9957);
nor UO_1360 (O_1360,N_9712,N_9393);
nand UO_1361 (O_1361,N_9497,N_9835);
and UO_1362 (O_1362,N_9969,N_9648);
nor UO_1363 (O_1363,N_9463,N_9058);
and UO_1364 (O_1364,N_9489,N_9378);
nand UO_1365 (O_1365,N_9888,N_9116);
or UO_1366 (O_1366,N_9334,N_9728);
nand UO_1367 (O_1367,N_9467,N_9774);
nand UO_1368 (O_1368,N_9045,N_9982);
nand UO_1369 (O_1369,N_9253,N_9159);
or UO_1370 (O_1370,N_9846,N_9300);
and UO_1371 (O_1371,N_9791,N_9674);
nand UO_1372 (O_1372,N_9471,N_9980);
nor UO_1373 (O_1373,N_9811,N_9349);
and UO_1374 (O_1374,N_9755,N_9890);
xnor UO_1375 (O_1375,N_9524,N_9236);
and UO_1376 (O_1376,N_9935,N_9114);
xnor UO_1377 (O_1377,N_9484,N_9548);
nor UO_1378 (O_1378,N_9928,N_9605);
or UO_1379 (O_1379,N_9877,N_9571);
and UO_1380 (O_1380,N_9805,N_9849);
and UO_1381 (O_1381,N_9609,N_9374);
nor UO_1382 (O_1382,N_9733,N_9181);
nor UO_1383 (O_1383,N_9113,N_9649);
nor UO_1384 (O_1384,N_9813,N_9929);
nand UO_1385 (O_1385,N_9701,N_9764);
xnor UO_1386 (O_1386,N_9416,N_9492);
and UO_1387 (O_1387,N_9143,N_9934);
and UO_1388 (O_1388,N_9766,N_9620);
and UO_1389 (O_1389,N_9050,N_9854);
nor UO_1390 (O_1390,N_9537,N_9588);
nand UO_1391 (O_1391,N_9324,N_9961);
or UO_1392 (O_1392,N_9900,N_9842);
or UO_1393 (O_1393,N_9286,N_9915);
or UO_1394 (O_1394,N_9427,N_9347);
or UO_1395 (O_1395,N_9029,N_9476);
or UO_1396 (O_1396,N_9294,N_9398);
or UO_1397 (O_1397,N_9830,N_9084);
and UO_1398 (O_1398,N_9980,N_9741);
nand UO_1399 (O_1399,N_9451,N_9664);
and UO_1400 (O_1400,N_9050,N_9557);
nand UO_1401 (O_1401,N_9492,N_9017);
xnor UO_1402 (O_1402,N_9671,N_9849);
and UO_1403 (O_1403,N_9379,N_9255);
or UO_1404 (O_1404,N_9073,N_9274);
nor UO_1405 (O_1405,N_9144,N_9750);
nor UO_1406 (O_1406,N_9353,N_9554);
or UO_1407 (O_1407,N_9226,N_9902);
nor UO_1408 (O_1408,N_9816,N_9525);
or UO_1409 (O_1409,N_9695,N_9924);
and UO_1410 (O_1410,N_9946,N_9991);
and UO_1411 (O_1411,N_9565,N_9606);
and UO_1412 (O_1412,N_9202,N_9993);
or UO_1413 (O_1413,N_9225,N_9514);
and UO_1414 (O_1414,N_9242,N_9334);
nand UO_1415 (O_1415,N_9920,N_9048);
or UO_1416 (O_1416,N_9791,N_9924);
nand UO_1417 (O_1417,N_9523,N_9457);
nor UO_1418 (O_1418,N_9694,N_9082);
nand UO_1419 (O_1419,N_9313,N_9624);
or UO_1420 (O_1420,N_9936,N_9915);
or UO_1421 (O_1421,N_9455,N_9687);
nor UO_1422 (O_1422,N_9834,N_9712);
nor UO_1423 (O_1423,N_9554,N_9738);
or UO_1424 (O_1424,N_9262,N_9110);
nand UO_1425 (O_1425,N_9498,N_9428);
and UO_1426 (O_1426,N_9195,N_9643);
nand UO_1427 (O_1427,N_9705,N_9195);
nor UO_1428 (O_1428,N_9618,N_9757);
or UO_1429 (O_1429,N_9682,N_9891);
and UO_1430 (O_1430,N_9426,N_9577);
nand UO_1431 (O_1431,N_9323,N_9421);
and UO_1432 (O_1432,N_9073,N_9963);
or UO_1433 (O_1433,N_9954,N_9052);
or UO_1434 (O_1434,N_9202,N_9293);
nor UO_1435 (O_1435,N_9430,N_9092);
nor UO_1436 (O_1436,N_9134,N_9065);
nand UO_1437 (O_1437,N_9170,N_9944);
nor UO_1438 (O_1438,N_9205,N_9781);
nand UO_1439 (O_1439,N_9031,N_9370);
and UO_1440 (O_1440,N_9459,N_9192);
nor UO_1441 (O_1441,N_9151,N_9641);
or UO_1442 (O_1442,N_9918,N_9835);
nor UO_1443 (O_1443,N_9546,N_9247);
or UO_1444 (O_1444,N_9293,N_9016);
nand UO_1445 (O_1445,N_9283,N_9376);
nor UO_1446 (O_1446,N_9451,N_9592);
or UO_1447 (O_1447,N_9146,N_9690);
nor UO_1448 (O_1448,N_9548,N_9277);
or UO_1449 (O_1449,N_9140,N_9607);
nor UO_1450 (O_1450,N_9972,N_9849);
or UO_1451 (O_1451,N_9423,N_9279);
nor UO_1452 (O_1452,N_9190,N_9315);
or UO_1453 (O_1453,N_9655,N_9557);
or UO_1454 (O_1454,N_9730,N_9212);
xnor UO_1455 (O_1455,N_9565,N_9469);
nand UO_1456 (O_1456,N_9701,N_9006);
nor UO_1457 (O_1457,N_9257,N_9077);
or UO_1458 (O_1458,N_9213,N_9830);
nand UO_1459 (O_1459,N_9428,N_9806);
nor UO_1460 (O_1460,N_9722,N_9841);
or UO_1461 (O_1461,N_9645,N_9898);
or UO_1462 (O_1462,N_9582,N_9789);
and UO_1463 (O_1463,N_9639,N_9449);
and UO_1464 (O_1464,N_9060,N_9833);
and UO_1465 (O_1465,N_9749,N_9395);
nor UO_1466 (O_1466,N_9200,N_9176);
nor UO_1467 (O_1467,N_9004,N_9201);
nor UO_1468 (O_1468,N_9444,N_9738);
and UO_1469 (O_1469,N_9538,N_9998);
nand UO_1470 (O_1470,N_9714,N_9075);
and UO_1471 (O_1471,N_9629,N_9260);
and UO_1472 (O_1472,N_9546,N_9272);
nor UO_1473 (O_1473,N_9785,N_9088);
nor UO_1474 (O_1474,N_9838,N_9117);
xnor UO_1475 (O_1475,N_9312,N_9599);
nor UO_1476 (O_1476,N_9729,N_9473);
nand UO_1477 (O_1477,N_9685,N_9859);
and UO_1478 (O_1478,N_9469,N_9344);
or UO_1479 (O_1479,N_9508,N_9161);
and UO_1480 (O_1480,N_9940,N_9823);
and UO_1481 (O_1481,N_9573,N_9130);
nand UO_1482 (O_1482,N_9594,N_9271);
or UO_1483 (O_1483,N_9931,N_9450);
or UO_1484 (O_1484,N_9892,N_9450);
and UO_1485 (O_1485,N_9655,N_9242);
nor UO_1486 (O_1486,N_9845,N_9609);
and UO_1487 (O_1487,N_9722,N_9015);
and UO_1488 (O_1488,N_9448,N_9582);
nand UO_1489 (O_1489,N_9846,N_9246);
or UO_1490 (O_1490,N_9244,N_9037);
nor UO_1491 (O_1491,N_9221,N_9707);
nor UO_1492 (O_1492,N_9332,N_9182);
nor UO_1493 (O_1493,N_9639,N_9921);
or UO_1494 (O_1494,N_9640,N_9476);
and UO_1495 (O_1495,N_9223,N_9449);
nand UO_1496 (O_1496,N_9675,N_9654);
nor UO_1497 (O_1497,N_9895,N_9499);
or UO_1498 (O_1498,N_9730,N_9924);
and UO_1499 (O_1499,N_9803,N_9952);
endmodule