module basic_3000_30000_3500_20_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nor U0 (N_0,In_1358,In_909);
nor U1 (N_1,In_1759,In_1210);
xor U2 (N_2,In_1754,In_261);
xnor U3 (N_3,In_2727,In_2957);
xnor U4 (N_4,In_981,In_345);
or U5 (N_5,In_2080,In_392);
nand U6 (N_6,In_993,In_2443);
nor U7 (N_7,In_654,In_34);
xnor U8 (N_8,In_1721,In_1971);
and U9 (N_9,In_1417,In_484);
and U10 (N_10,In_1433,In_2208);
and U11 (N_11,In_529,In_1834);
or U12 (N_12,In_92,In_459);
nand U13 (N_13,In_2608,In_1154);
nand U14 (N_14,In_2797,In_2534);
xnor U15 (N_15,In_89,In_729);
xnor U16 (N_16,In_2870,In_1114);
nand U17 (N_17,In_2025,In_2967);
nand U18 (N_18,In_1564,In_2357);
nand U19 (N_19,In_867,In_977);
xnor U20 (N_20,In_814,In_887);
nand U21 (N_21,In_2193,In_1791);
xor U22 (N_22,In_1609,In_255);
nor U23 (N_23,In_7,In_2773);
or U24 (N_24,In_1751,In_1265);
nand U25 (N_25,In_2513,In_690);
xor U26 (N_26,In_2987,In_1818);
nor U27 (N_27,In_1195,In_970);
and U28 (N_28,In_1938,In_640);
and U29 (N_29,In_296,In_2110);
or U30 (N_30,In_28,In_2878);
and U31 (N_31,In_1365,In_660);
and U32 (N_32,In_2910,In_1402);
nor U33 (N_33,In_2285,In_363);
nand U34 (N_34,In_2273,In_1764);
xnor U35 (N_35,In_2129,In_2146);
xnor U36 (N_36,In_903,In_4);
or U37 (N_37,In_2504,In_830);
or U38 (N_38,In_451,In_643);
nand U39 (N_39,In_986,In_2127);
and U40 (N_40,In_1549,In_2275);
xor U41 (N_41,In_2834,In_1303);
nor U42 (N_42,In_450,In_2259);
and U43 (N_43,In_330,In_305);
xor U44 (N_44,In_2133,In_2658);
nor U45 (N_45,In_989,In_2798);
and U46 (N_46,In_2388,In_143);
nor U47 (N_47,In_1249,In_1837);
nor U48 (N_48,In_2576,In_2912);
and U49 (N_49,In_2941,In_1251);
and U50 (N_50,In_1998,In_2569);
and U51 (N_51,In_2663,In_418);
and U52 (N_52,In_793,In_2284);
and U53 (N_53,In_403,In_2488);
and U54 (N_54,In_2360,In_2184);
nand U55 (N_55,In_120,In_2947);
and U56 (N_56,In_966,In_1250);
and U57 (N_57,In_2304,In_1792);
xnor U58 (N_58,In_838,In_1723);
nor U59 (N_59,In_2254,In_247);
or U60 (N_60,In_727,In_1187);
or U61 (N_61,In_127,In_937);
nor U62 (N_62,In_2832,In_2078);
xor U63 (N_63,In_806,In_269);
nor U64 (N_64,In_2328,In_1228);
nand U65 (N_65,In_709,In_782);
or U66 (N_66,In_338,In_2567);
nand U67 (N_67,In_1184,In_2483);
nand U68 (N_68,In_1127,In_647);
nor U69 (N_69,In_1933,In_41);
or U70 (N_70,In_949,In_1682);
nor U71 (N_71,In_693,In_1934);
xor U72 (N_72,In_1239,In_2082);
or U73 (N_73,In_2026,In_1599);
or U74 (N_74,In_2010,In_552);
nand U75 (N_75,In_1364,In_286);
nor U76 (N_76,In_2351,In_776);
and U77 (N_77,In_2323,In_2937);
and U78 (N_78,In_1438,In_2035);
nand U79 (N_79,In_2215,In_539);
nor U80 (N_80,In_1879,In_1530);
nor U81 (N_81,In_1805,In_388);
nor U82 (N_82,In_657,In_868);
nor U83 (N_83,In_2991,In_1084);
nand U84 (N_84,In_1427,In_1204);
nor U85 (N_85,In_118,In_2940);
nand U86 (N_86,In_2480,In_195);
and U87 (N_87,In_465,In_2506);
xnor U88 (N_88,In_2349,In_2058);
nand U89 (N_89,In_2620,In_275);
and U90 (N_90,In_163,In_2482);
and U91 (N_91,In_2337,In_580);
and U92 (N_92,In_2116,In_891);
xnor U93 (N_93,In_2302,In_2740);
nand U94 (N_94,In_1973,In_568);
xor U95 (N_95,In_495,In_2801);
and U96 (N_96,In_1028,In_1581);
or U97 (N_97,In_417,In_760);
nand U98 (N_98,In_1103,In_1387);
or U99 (N_99,In_601,In_2889);
xnor U100 (N_100,In_1651,In_1768);
nor U101 (N_101,In_2770,In_954);
xor U102 (N_102,In_1489,In_1864);
xor U103 (N_103,In_1355,In_2476);
xnor U104 (N_104,In_1687,In_503);
nand U105 (N_105,In_1146,In_979);
xnor U106 (N_106,In_2516,In_1869);
nor U107 (N_107,In_1806,In_2712);
or U108 (N_108,In_2134,In_1141);
xnor U109 (N_109,In_2697,In_245);
nor U110 (N_110,In_1510,In_1883);
xnor U111 (N_111,In_2097,In_570);
xnor U112 (N_112,In_2218,In_2996);
and U113 (N_113,In_1529,In_2120);
xnor U114 (N_114,In_2494,In_871);
and U115 (N_115,In_2682,In_1590);
nand U116 (N_116,In_2175,In_1331);
nor U117 (N_117,In_1371,In_1099);
nand U118 (N_118,In_694,In_75);
and U119 (N_119,In_683,In_2156);
or U120 (N_120,In_1043,In_447);
nand U121 (N_121,In_1385,In_859);
xor U122 (N_122,In_946,In_1380);
and U123 (N_123,In_577,In_2990);
nand U124 (N_124,In_1755,In_209);
nor U125 (N_125,In_1793,In_721);
nor U126 (N_126,In_825,In_1812);
nor U127 (N_127,In_2203,In_2370);
and U128 (N_128,In_49,In_1006);
or U129 (N_129,In_2105,In_1844);
nand U130 (N_130,In_742,In_2547);
and U131 (N_131,In_186,In_1594);
nand U132 (N_132,In_565,In_1205);
xnor U133 (N_133,In_182,In_944);
nand U134 (N_134,In_1736,In_1875);
or U135 (N_135,In_1074,In_2316);
xnor U136 (N_136,In_1993,In_1577);
nand U137 (N_137,In_708,In_1895);
and U138 (N_138,In_2309,In_1740);
and U139 (N_139,In_2319,In_254);
or U140 (N_140,In_2719,In_393);
and U141 (N_141,In_2264,In_2391);
nor U142 (N_142,In_1468,In_2907);
nor U143 (N_143,In_2693,In_2439);
xor U144 (N_144,In_1002,In_1904);
nand U145 (N_145,In_1802,In_2074);
xor U146 (N_146,In_386,In_2123);
and U147 (N_147,In_822,In_1817);
nor U148 (N_148,In_1928,In_1282);
xor U149 (N_149,In_1729,In_2999);
nor U150 (N_150,In_688,In_215);
nand U151 (N_151,In_2161,In_2532);
xnor U152 (N_152,In_1992,In_2292);
or U153 (N_153,In_159,In_1444);
and U154 (N_154,In_546,In_2242);
and U155 (N_155,In_2921,In_1559);
and U156 (N_156,In_1674,In_1872);
or U157 (N_157,In_131,In_119);
nand U158 (N_158,In_2070,In_2462);
xor U159 (N_159,In_1470,In_508);
xnor U160 (N_160,In_2998,In_288);
or U161 (N_161,In_1953,In_627);
or U162 (N_162,In_2306,In_1563);
nor U163 (N_163,In_905,In_950);
or U164 (N_164,In_1156,In_609);
or U165 (N_165,In_30,In_2627);
nor U166 (N_166,In_2826,In_2326);
xnor U167 (N_167,In_274,In_784);
xor U168 (N_168,In_2185,In_860);
and U169 (N_169,In_2952,In_1369);
nor U170 (N_170,In_2313,In_2979);
or U171 (N_171,In_2509,In_1996);
nand U172 (N_172,In_1461,In_2631);
xnor U173 (N_173,In_2041,In_2964);
or U174 (N_174,In_6,In_1349);
xor U175 (N_175,In_2278,In_679);
or U176 (N_176,In_1691,In_2322);
and U177 (N_177,In_479,In_1541);
nand U178 (N_178,In_723,In_2290);
or U179 (N_179,In_1741,In_169);
nand U180 (N_180,In_472,In_1058);
nand U181 (N_181,In_2841,In_302);
or U182 (N_182,In_464,In_545);
xnor U183 (N_183,In_732,In_2380);
nor U184 (N_184,In_337,In_2039);
or U185 (N_185,In_2427,In_1675);
and U186 (N_186,In_1334,In_2831);
and U187 (N_187,In_2455,In_1714);
nand U188 (N_188,In_1424,In_551);
nor U189 (N_189,In_278,In_843);
nor U190 (N_190,In_1843,In_1177);
and U191 (N_191,In_2685,In_2481);
nand U192 (N_192,In_1273,In_1968);
xnor U193 (N_193,In_1857,In_1639);
nor U194 (N_194,In_2020,In_2873);
nor U195 (N_195,In_2965,In_1051);
and U196 (N_196,In_1743,In_2782);
or U197 (N_197,In_2104,In_1964);
xnor U198 (N_198,In_139,In_817);
nand U199 (N_199,In_942,In_1285);
or U200 (N_200,In_1218,In_1931);
xnor U201 (N_201,In_2823,In_1652);
nand U202 (N_202,In_921,In_1025);
nor U203 (N_203,In_2007,In_2718);
xor U204 (N_204,In_1499,In_325);
and U205 (N_205,In_2840,In_629);
nand U206 (N_206,In_2670,In_2706);
nor U207 (N_207,In_344,In_1143);
and U208 (N_208,In_51,In_1272);
nand U209 (N_209,In_1975,In_757);
xnor U210 (N_210,In_2407,In_1897);
or U211 (N_211,In_107,In_291);
nor U212 (N_212,In_1955,In_1268);
nand U213 (N_213,In_415,In_1160);
or U214 (N_214,In_2400,In_1023);
and U215 (N_215,In_1752,In_831);
nor U216 (N_216,In_470,In_1894);
nand U217 (N_217,In_2027,In_2923);
xnor U218 (N_218,In_2002,In_2543);
xor U219 (N_219,In_481,In_399);
and U220 (N_220,In_1466,In_54);
nand U221 (N_221,In_2913,In_2593);
and U222 (N_222,In_967,In_1400);
xor U223 (N_223,In_1874,In_411);
and U224 (N_224,In_395,In_2283);
and U225 (N_225,In_1799,In_2880);
nor U226 (N_226,In_533,In_1645);
nor U227 (N_227,In_2938,In_492);
nand U228 (N_228,In_1207,In_2363);
xor U229 (N_229,In_2911,In_743);
nand U230 (N_230,In_733,In_2997);
xnor U231 (N_231,In_1881,In_1685);
nor U232 (N_232,In_112,In_2949);
and U233 (N_233,In_2881,In_982);
nor U234 (N_234,In_372,In_1474);
nor U235 (N_235,In_1479,In_1698);
or U236 (N_236,In_1570,In_243);
nor U237 (N_237,In_2368,In_2687);
nand U238 (N_238,In_162,In_2066);
xnor U239 (N_239,In_2850,In_586);
and U240 (N_240,In_1157,In_1943);
nor U241 (N_241,In_359,In_68);
and U242 (N_242,In_1488,In_2032);
nor U243 (N_243,In_2886,In_1608);
nand U244 (N_244,In_611,In_2711);
nand U245 (N_245,In_483,In_358);
xnor U246 (N_246,In_1319,In_452);
nor U247 (N_247,In_2595,In_2386);
nand U248 (N_248,In_383,In_1071);
xnor U249 (N_249,In_656,In_960);
xor U250 (N_250,In_2471,In_2836);
and U251 (N_251,In_796,In_246);
nand U252 (N_252,In_886,In_360);
nor U253 (N_253,In_1647,In_1936);
xor U254 (N_254,In_1669,In_2746);
or U255 (N_255,In_1356,In_649);
or U256 (N_256,In_2170,In_2311);
xnor U257 (N_257,In_1450,In_2924);
nand U258 (N_258,In_2508,In_1505);
and U259 (N_259,In_252,In_1136);
nor U260 (N_260,In_1761,In_841);
xor U261 (N_261,In_914,In_2069);
nor U262 (N_262,In_1109,In_1448);
nand U263 (N_263,In_2046,In_2882);
nor U264 (N_264,In_2745,In_501);
or U265 (N_265,In_1506,In_715);
nand U266 (N_266,In_1306,In_2568);
or U267 (N_267,In_64,In_1354);
xnor U268 (N_268,In_2668,In_477);
xor U269 (N_269,In_2592,In_1014);
xnor U270 (N_270,In_1893,In_1392);
and U271 (N_271,In_1262,In_1101);
and U272 (N_272,In_521,In_2022);
or U273 (N_273,In_1924,In_998);
nor U274 (N_274,In_2475,In_1738);
and U275 (N_275,In_2739,In_1560);
nand U276 (N_276,In_1889,In_1910);
or U277 (N_277,In_2255,In_384);
or U278 (N_278,In_926,In_198);
or U279 (N_279,In_579,In_2409);
or U280 (N_280,In_2993,In_136);
xnor U281 (N_281,In_1223,In_2174);
and U282 (N_282,In_2209,In_2945);
nand U283 (N_283,In_1460,In_351);
nand U284 (N_284,In_1199,In_2616);
nor U285 (N_285,In_2399,In_1970);
xor U286 (N_286,In_1001,In_1307);
xnor U287 (N_287,In_414,In_1870);
and U288 (N_288,In_2795,In_1238);
xor U289 (N_289,In_596,In_73);
nor U290 (N_290,In_1604,In_560);
nand U291 (N_291,In_756,In_2604);
and U292 (N_292,In_267,In_1010);
nor U293 (N_293,In_204,In_1850);
nor U294 (N_294,In_2437,In_129);
xnor U295 (N_295,In_170,In_2893);
nand U296 (N_296,In_1467,In_1062);
xor U297 (N_297,In_572,In_865);
and U298 (N_298,In_513,In_2454);
xnor U299 (N_299,In_1007,In_2198);
or U300 (N_300,In_2503,In_558);
and U301 (N_301,In_1048,In_193);
or U302 (N_302,In_592,In_2294);
xor U303 (N_303,In_2920,In_1416);
and U304 (N_304,In_2050,In_105);
nand U305 (N_305,In_1018,In_1659);
nor U306 (N_306,In_1591,In_2853);
nand U307 (N_307,In_697,In_2601);
or U308 (N_308,In_922,In_2270);
xnor U309 (N_309,In_2724,In_199);
or U310 (N_310,In_2710,In_2220);
nor U311 (N_311,In_740,In_2771);
nor U312 (N_312,In_2436,In_1453);
nand U313 (N_313,In_2819,In_826);
nand U314 (N_314,In_1965,In_1621);
and U315 (N_315,In_1983,In_1600);
nand U316 (N_316,In_851,In_2111);
and U317 (N_317,In_778,In_583);
nand U318 (N_318,In_2644,In_2128);
and U319 (N_319,In_2461,In_2808);
or U320 (N_320,In_2582,In_1497);
and U321 (N_321,In_2365,In_1767);
or U322 (N_322,In_175,In_316);
xor U323 (N_323,In_2154,In_1397);
xor U324 (N_324,In_295,In_1341);
and U325 (N_325,In_2778,In_2969);
or U326 (N_326,In_2056,In_1734);
and U327 (N_327,In_2546,In_2694);
xnor U328 (N_328,In_1871,In_1391);
or U329 (N_329,In_2757,In_430);
or U330 (N_330,In_1289,In_226);
xnor U331 (N_331,In_2879,In_206);
or U332 (N_332,In_675,In_2239);
nor U333 (N_333,In_2837,In_2384);
xor U334 (N_334,In_1633,In_2062);
and U335 (N_335,In_1966,In_2825);
nand U336 (N_336,In_355,In_1327);
and U337 (N_337,In_714,In_2344);
and U338 (N_338,In_728,In_2635);
xor U339 (N_339,In_2673,In_1293);
nand U340 (N_340,In_1941,In_233);
or U341 (N_341,In_2667,In_900);
and U342 (N_342,In_700,In_2354);
and U343 (N_343,In_47,In_549);
xnor U344 (N_344,In_379,In_1286);
or U345 (N_345,In_842,In_1537);
nand U346 (N_346,In_534,In_84);
xnor U347 (N_347,In_2652,In_951);
xnor U348 (N_348,In_1437,In_1381);
or U349 (N_349,In_1361,In_229);
and U350 (N_350,In_2009,In_1902);
xnor U351 (N_351,In_1649,In_1192);
or U352 (N_352,In_745,In_1994);
nor U353 (N_353,In_2452,In_2001);
or U354 (N_354,In_1015,In_189);
nand U355 (N_355,In_1059,In_478);
nand U356 (N_356,In_1935,In_624);
xnor U357 (N_357,In_1828,In_2347);
xor U358 (N_358,In_2160,In_293);
nor U359 (N_359,In_468,In_837);
and U360 (N_360,In_1022,In_1235);
and U361 (N_361,In_1884,In_2570);
and U362 (N_362,In_1906,In_1840);
xnor U363 (N_363,In_1706,In_60);
and U364 (N_364,In_2390,In_2141);
xnor U365 (N_365,In_443,In_666);
xnor U366 (N_366,In_2647,In_561);
xnor U367 (N_367,In_1950,In_2519);
nand U368 (N_368,In_783,In_724);
or U369 (N_369,In_2251,In_1703);
nand U370 (N_370,In_781,In_2792);
xor U371 (N_371,In_1072,In_1209);
or U372 (N_372,In_2079,In_1390);
and U373 (N_373,In_2816,In_767);
nor U374 (N_374,In_1471,In_108);
nor U375 (N_375,In_347,In_2325);
or U376 (N_376,In_2790,In_2854);
nand U377 (N_377,In_2226,In_2342);
xnor U378 (N_378,In_987,In_1571);
xnor U379 (N_379,In_1915,In_1255);
nor U380 (N_380,In_1845,In_397);
or U381 (N_381,In_2491,In_766);
xnor U382 (N_382,In_805,In_436);
or U383 (N_383,In_2700,In_2151);
nand U384 (N_384,In_2406,In_1670);
xnor U385 (N_385,In_735,In_913);
nand U386 (N_386,In_336,In_90);
nand U387 (N_387,In_1627,In_2868);
and U388 (N_388,In_150,In_2828);
or U389 (N_389,In_190,In_439);
nand U390 (N_390,In_1495,In_357);
nand U391 (N_391,In_227,In_98);
nand U392 (N_392,In_1795,In_2232);
or U393 (N_393,In_378,In_884);
xnor U394 (N_394,In_2250,In_1082);
nand U395 (N_395,In_1820,In_497);
and U396 (N_396,In_1532,In_2199);
xor U397 (N_397,In_1287,In_301);
nor U398 (N_398,In_2684,In_2733);
xor U399 (N_399,In_1991,In_976);
and U400 (N_400,In_2762,In_815);
nor U401 (N_401,In_2691,In_40);
xnor U402 (N_402,In_1725,In_2340);
or U403 (N_403,In_1317,In_582);
nand U404 (N_404,In_2061,In_848);
nor U405 (N_405,In_795,In_2467);
nor U406 (N_406,In_2662,In_466);
nor U407 (N_407,In_234,In_1350);
nor U408 (N_408,In_1690,In_2445);
and U409 (N_409,In_2432,In_1498);
nand U410 (N_410,In_2403,In_2899);
xor U411 (N_411,In_2064,In_114);
nand U412 (N_412,In_346,In_863);
or U413 (N_413,In_2268,In_1584);
xnor U414 (N_414,In_2925,In_2367);
nand U415 (N_415,In_1203,In_1961);
xnor U416 (N_416,In_2810,In_791);
xor U417 (N_417,In_2555,In_2666);
nand U418 (N_418,In_2962,In_297);
nand U419 (N_419,In_854,In_2291);
nand U420 (N_420,In_2152,In_134);
nand U421 (N_421,In_1019,In_111);
xnor U422 (N_422,In_1900,In_404);
xor U423 (N_423,In_875,In_705);
and U424 (N_424,In_2522,In_1665);
nor U425 (N_425,In_1044,In_1395);
or U426 (N_426,In_540,In_1679);
or U427 (N_427,In_232,In_2971);
nand U428 (N_428,In_824,In_1359);
and U429 (N_429,In_2638,In_1513);
and U430 (N_430,In_1054,In_1715);
or U431 (N_431,In_2589,In_2888);
nand U432 (N_432,In_1052,In_1903);
xor U433 (N_433,In_165,In_1447);
and U434 (N_434,In_803,In_1423);
or U435 (N_435,In_2672,In_974);
and U436 (N_436,In_2614,In_2789);
xor U437 (N_437,In_125,In_527);
and U438 (N_438,In_2791,In_1403);
and U439 (N_439,In_1543,In_1113);
and U440 (N_440,In_489,In_659);
nor U441 (N_441,In_1110,In_2732);
xor U442 (N_442,In_1276,In_2645);
and U443 (N_443,In_1511,In_1295);
or U444 (N_444,In_1353,In_928);
nand U445 (N_445,In_1108,In_1663);
xnor U446 (N_446,In_419,In_1986);
nor U447 (N_447,In_1727,In_941);
and U448 (N_448,In_1678,In_520);
or U449 (N_449,In_1462,In_2894);
and U450 (N_450,In_829,In_260);
nand U451 (N_451,In_1237,In_2261);
nand U452 (N_452,In_2600,In_181);
or U453 (N_453,In_1758,In_2521);
nand U454 (N_454,In_2258,In_1275);
nand U455 (N_455,In_608,In_562);
xor U456 (N_456,In_1509,In_2550);
nand U457 (N_457,In_259,In_1032);
nand U458 (N_458,In_630,In_2813);
xor U459 (N_459,In_2702,In_2995);
xor U460 (N_460,In_29,In_1115);
or U461 (N_461,In_2037,In_599);
and U462 (N_462,In_2845,In_2588);
and U463 (N_463,In_1765,In_2728);
and U464 (N_464,In_716,In_1455);
xnor U465 (N_465,In_1990,In_573);
nand U466 (N_466,In_2247,In_1882);
nor U467 (N_467,In_1069,In_703);
or U468 (N_468,In_2905,In_1603);
nor U469 (N_469,In_2043,In_2063);
nand U470 (N_470,In_606,In_486);
and U471 (N_471,In_591,In_2787);
nand U472 (N_472,In_2851,In_1167);
xor U473 (N_473,In_948,In_1330);
nand U474 (N_474,In_2090,In_2927);
nand U475 (N_475,In_2866,In_1719);
nor U476 (N_476,In_2219,In_2742);
nand U477 (N_477,In_2353,In_1304);
and U478 (N_478,In_2736,In_1957);
nor U479 (N_479,In_1568,In_2763);
nor U480 (N_480,In_2747,In_1042);
nand U481 (N_481,In_203,In_930);
nor U482 (N_482,In_2210,In_1551);
nand U483 (N_483,In_855,In_853);
nor U484 (N_484,In_634,In_564);
and U485 (N_485,In_1085,In_2159);
nor U486 (N_486,In_1456,In_1097);
and U487 (N_487,In_1852,In_1756);
or U488 (N_488,In_626,In_2171);
or U489 (N_489,In_1086,In_1034);
or U490 (N_490,In_1625,In_2619);
and U491 (N_491,In_1024,In_1368);
nand U492 (N_492,In_2815,In_2562);
or U493 (N_493,In_1717,In_2656);
nand U494 (N_494,In_1526,In_2574);
xnor U495 (N_495,In_1377,In_2341);
or U496 (N_496,In_1841,In_2520);
nor U497 (N_497,In_2705,In_2817);
and U498 (N_498,In_23,In_1213);
nor U499 (N_499,In_754,In_1219);
xnor U500 (N_500,In_895,In_958);
nor U501 (N_501,In_927,In_2238);
nor U502 (N_502,In_1348,In_401);
nand U503 (N_503,In_2005,In_1280);
nand U504 (N_504,In_216,In_2122);
and U505 (N_505,In_687,In_1650);
or U506 (N_506,In_2654,In_1801);
nor U507 (N_507,In_2846,In_2484);
nand U508 (N_508,In_819,In_1742);
nor U509 (N_509,In_2256,In_2413);
nand U510 (N_510,In_2699,In_1020);
xor U511 (N_511,In_1261,In_102);
xor U512 (N_512,In_2678,In_1716);
nor U513 (N_513,In_42,In_1798);
xnor U514 (N_514,In_2463,In_1995);
nor U515 (N_515,In_67,In_771);
nand U516 (N_516,In_437,In_2003);
xor U517 (N_517,In_510,In_1472);
and U518 (N_518,In_2676,In_1561);
or U519 (N_519,In_2603,In_2206);
or U520 (N_520,In_2777,In_1038);
nand U521 (N_521,In_441,In_664);
and U522 (N_522,In_2892,In_711);
nand U523 (N_523,In_176,In_1270);
xnor U524 (N_524,In_2982,In_205);
xor U525 (N_525,In_1345,In_1155);
nand U526 (N_526,In_61,In_1425);
xnor U527 (N_527,In_1822,In_2717);
and U528 (N_528,In_786,In_1284);
and U529 (N_529,In_2628,In_1313);
nand U530 (N_530,In_390,In_2495);
and U531 (N_531,In_2060,In_1899);
xor U532 (N_532,In_335,In_1533);
nand U533 (N_533,In_2338,In_2269);
nor U534 (N_534,In_96,In_622);
nand U535 (N_535,In_738,In_1245);
nor U536 (N_536,In_898,In_2867);
nand U537 (N_537,In_371,In_1831);
or U538 (N_538,In_53,In_2946);
xnor U539 (N_539,In_2350,In_343);
xor U540 (N_540,In_2561,In_1748);
xor U541 (N_541,In_1972,In_1139);
nor U542 (N_542,In_1839,In_2753);
xnor U543 (N_543,In_2478,In_1713);
and U544 (N_544,In_2468,In_2646);
xor U545 (N_545,In_2180,In_1605);
nand U546 (N_546,In_1301,In_179);
nand U547 (N_547,In_1016,In_1636);
xor U548 (N_548,In_2440,In_1865);
xor U549 (N_549,In_811,In_78);
or U550 (N_550,In_1333,In_33);
and U551 (N_551,In_1316,In_1112);
nor U552 (N_552,In_444,In_1773);
xor U553 (N_553,In_122,In_2890);
nand U554 (N_554,In_172,In_2012);
or U555 (N_555,In_1763,In_1266);
and U556 (N_556,In_631,In_2359);
nor U557 (N_557,In_1393,In_1693);
nand U558 (N_558,In_1324,In_2597);
nor U559 (N_559,In_2143,In_2930);
and U560 (N_560,In_1528,In_2108);
xor U561 (N_561,In_21,In_2540);
nand U562 (N_562,In_487,In_166);
or U563 (N_563,In_1244,In_2785);
and U564 (N_564,In_1892,In_1554);
and U565 (N_565,In_1208,In_1696);
nand U566 (N_566,In_66,In_1866);
or U567 (N_567,In_2166,In_1332);
nor U568 (N_568,In_1206,In_1782);
nor U569 (N_569,In_1579,In_1216);
or U570 (N_570,In_2249,In_1976);
xnor U571 (N_571,In_1057,In_1070);
nand U572 (N_572,In_2263,In_910);
or U573 (N_573,In_1544,In_1578);
xnor U574 (N_574,In_2759,In_423);
nor U575 (N_575,In_2827,In_2373);
and U576 (N_576,In_2411,In_957);
xor U577 (N_577,In_2805,In_85);
nand U578 (N_578,In_1312,In_2665);
nand U579 (N_579,In_2486,In_1386);
or U580 (N_580,In_780,In_2767);
and U581 (N_581,In_2501,In_1618);
nand U582 (N_582,In_2293,In_965);
nand U583 (N_583,In_576,In_2430);
or U584 (N_584,In_2928,In_2076);
and U585 (N_585,In_1056,In_178);
and U586 (N_586,In_1648,In_2541);
nand U587 (N_587,In_2877,In_224);
xnor U588 (N_588,In_408,In_2240);
xor U589 (N_589,In_787,In_2094);
nand U590 (N_590,In_1624,In_448);
nand U591 (N_591,In_453,In_1811);
or U592 (N_592,In_1325,In_469);
nand U593 (N_593,In_1490,In_2267);
nor U594 (N_594,In_1181,In_1012);
xor U595 (N_595,In_1919,In_2958);
nor U596 (N_596,In_59,In_171);
xnor U597 (N_597,In_2017,In_113);
xnor U598 (N_598,In_2343,In_2824);
xnor U599 (N_599,In_1419,In_902);
xor U600 (N_600,In_1642,In_2650);
and U601 (N_601,In_2004,In_731);
or U602 (N_602,In_2119,In_1458);
nor U603 (N_603,In_1179,In_1477);
nand U604 (N_604,In_2132,In_1920);
or U605 (N_605,In_416,In_197);
and U606 (N_606,In_2554,In_307);
or U607 (N_607,In_2307,In_554);
nor U608 (N_608,In_2202,In_2956);
or U609 (N_609,In_1226,In_1299);
and U610 (N_610,In_1493,In_2751);
or U611 (N_611,In_929,In_2548);
nor U612 (N_612,In_2028,In_241);
nand U613 (N_613,In_1794,In_1073);
nor U614 (N_614,In_1566,In_2934);
and U615 (N_615,In_2289,In_1783);
xor U616 (N_616,In_621,In_1407);
nor U617 (N_617,In_633,In_480);
nand U618 (N_618,In_1138,In_542);
or U619 (N_619,In_2788,In_2221);
xnor U620 (N_620,In_1657,In_314);
nand U621 (N_621,In_2317,In_1008);
xor U622 (N_622,In_712,In_1434);
nand U623 (N_623,In_685,In_2149);
or U624 (N_624,In_2101,In_1017);
nor U625 (N_625,In_1100,In_1093);
xor U626 (N_626,In_559,In_1277);
nor U627 (N_627,In_1375,In_1514);
and U628 (N_628,In_1984,In_739);
xnor U629 (N_629,In_673,In_475);
or U630 (N_630,In_434,In_1290);
xor U631 (N_631,In_123,In_2228);
nand U632 (N_632,In_270,In_1147);
nand U633 (N_633,In_2774,In_106);
nor U634 (N_634,In_1372,In_2015);
xor U635 (N_635,In_2818,In_2915);
xnor U636 (N_636,In_2262,In_1501);
xnor U637 (N_637,In_2299,In_2738);
nor U638 (N_638,In_2081,In_1807);
xor U639 (N_639,In_361,In_2114);
xnor U640 (N_640,In_333,In_1516);
xnor U641 (N_641,In_924,In_1248);
nor U642 (N_642,In_2490,In_334);
and U643 (N_643,In_2944,In_2985);
xnor U644 (N_644,In_1810,In_605);
nand U645 (N_645,In_256,In_1766);
and U646 (N_646,In_1105,In_485);
nor U647 (N_647,In_1135,In_230);
and U648 (N_648,In_2809,In_846);
or U649 (N_649,In_2405,In_2287);
or U650 (N_650,In_968,In_590);
nor U651 (N_651,In_1930,In_320);
or U652 (N_652,In_2625,In_496);
nor U653 (N_653,In_1021,In_713);
or U654 (N_654,In_904,In_2820);
and U655 (N_655,In_222,In_258);
nand U656 (N_656,In_571,In_2075);
xor U657 (N_657,In_1692,In_665);
xnor U658 (N_658,In_1033,In_2356);
and U659 (N_659,In_1847,In_1853);
xor U660 (N_660,In_1730,In_460);
nor U661 (N_661,In_223,In_1412);
nand U662 (N_662,In_200,In_158);
and U663 (N_663,In_116,In_2917);
nand U664 (N_664,In_720,In_1712);
xor U665 (N_665,In_1908,In_1629);
nor U666 (N_666,In_1030,In_828);
or U667 (N_667,In_2843,In_1126);
xnor U668 (N_668,In_1263,In_2444);
or U669 (N_669,In_318,In_177);
or U670 (N_670,In_1267,In_1762);
xor U671 (N_671,In_1538,In_2583);
and U672 (N_672,In_1329,In_2086);
nand U673 (N_673,In_1620,In_1484);
and U674 (N_674,In_1066,In_512);
nand U675 (N_675,In_2044,In_706);
nand U676 (N_676,In_2634,In_1821);
or U677 (N_677,In_128,In_263);
xnor U678 (N_678,In_2000,In_2376);
nand U679 (N_679,In_272,In_519);
nor U680 (N_680,In_82,In_276);
nor U681 (N_681,In_313,In_628);
xnor U682 (N_682,In_862,In_975);
xor U683 (N_683,In_916,In_2321);
nand U684 (N_684,In_1457,In_1227);
nor U685 (N_685,In_1431,In_168);
nand U686 (N_686,In_777,In_1116);
nor U687 (N_687,In_95,In_461);
nor U688 (N_688,In_2435,In_2803);
nand U689 (N_689,In_1378,In_997);
nand U690 (N_690,In_1653,In_65);
nand U691 (N_691,In_668,In_2098);
and U692 (N_692,In_455,In_1880);
nor U693 (N_693,In_994,In_812);
nand U694 (N_694,In_422,In_2176);
and U695 (N_695,In_1132,In_1664);
xnor U696 (N_696,In_1088,In_2052);
or U697 (N_697,In_2655,In_2187);
or U698 (N_698,In_20,In_1589);
nor U699 (N_699,In_2661,In_1318);
nor U700 (N_700,In_2914,In_1320);
and U701 (N_701,In_1917,In_2204);
and U702 (N_702,In_1172,In_2113);
nor U703 (N_703,In_567,In_2192);
and U704 (N_704,In_1547,In_2327);
nand U705 (N_705,In_1186,In_421);
nor U706 (N_706,In_2355,In_615);
and U707 (N_707,In_1940,In_1118);
and U708 (N_708,In_242,In_1164);
xor U709 (N_709,In_1323,In_872);
nand U710 (N_710,In_2095,In_569);
nor U711 (N_711,In_2806,In_341);
and U712 (N_712,In_1326,In_1482);
nand U713 (N_713,In_912,In_890);
xor U714 (N_714,In_1414,In_446);
nor U715 (N_715,In_1449,In_2931);
nand U716 (N_716,In_310,In_217);
xnor U717 (N_717,In_614,In_225);
and U718 (N_718,In_160,In_2720);
nor U719 (N_719,In_2053,In_1830);
xor U720 (N_720,In_69,In_1827);
and U721 (N_721,In_2244,In_1258);
xnor U722 (N_722,In_1373,In_774);
nor U723 (N_723,In_2364,In_790);
nor U724 (N_724,In_280,In_137);
or U725 (N_725,In_598,In_1780);
or U726 (N_726,In_2714,In_50);
and U727 (N_727,In_1300,In_488);
xor U728 (N_728,In_1531,In_2531);
nand U729 (N_729,In_1366,In_431);
nor U730 (N_730,In_1520,In_2395);
xnor U731 (N_731,In_2681,In_2722);
xnor U732 (N_732,In_377,In_2392);
nor U733 (N_733,In_2756,In_1796);
nand U734 (N_734,In_1596,In_482);
nand U735 (N_735,In_1481,In_1169);
nor U736 (N_736,In_1357,In_1129);
xnor U737 (N_737,In_147,In_1668);
nor U738 (N_738,In_2799,In_2707);
or U739 (N_739,In_1724,In_196);
nand U740 (N_740,In_1336,In_1120);
or U741 (N_741,In_2847,In_2420);
and U742 (N_742,In_321,In_2498);
nor U743 (N_743,In_1635,In_1540);
nand U744 (N_744,In_1704,In_2303);
or U745 (N_745,In_555,In_595);
and U746 (N_746,In_1896,In_1886);
nor U747 (N_747,In_2216,In_2779);
xor U748 (N_748,In_722,In_1310);
nand U749 (N_749,In_1646,In_328);
nand U750 (N_750,In_2425,In_309);
xnor U751 (N_751,In_1439,In_880);
xnor U752 (N_752,In_1684,In_2951);
xor U753 (N_753,In_827,In_1662);
nand U754 (N_754,In_719,In_1952);
nor U755 (N_755,In_1410,In_103);
nor U756 (N_756,In_257,In_2992);
or U757 (N_757,In_279,In_2051);
nand U758 (N_758,In_1785,In_2901);
and U759 (N_759,In_1429,In_2535);
nand U760 (N_760,In_2874,In_1912);
nor U761 (N_761,In_1885,In_273);
or U762 (N_762,In_2458,In_1230);
nor U763 (N_763,In_834,In_409);
xnor U764 (N_764,In_1779,In_1194);
xnor U765 (N_765,In_1980,In_2112);
nand U766 (N_766,In_2415,In_109);
or U767 (N_767,In_2217,In_566);
or U768 (N_768,In_237,In_1096);
xor U769 (N_769,In_772,In_2281);
xnor U770 (N_770,In_2396,In_88);
nor U771 (N_771,In_1573,In_684);
nand U772 (N_772,In_25,In_769);
or U773 (N_773,In_636,In_2980);
or U774 (N_774,In_18,In_2473);
xor U775 (N_775,In_1451,In_2158);
nand U776 (N_776,In_2330,In_816);
nor U777 (N_777,In_1702,In_725);
nor U778 (N_778,In_1374,In_208);
nor U779 (N_779,In_2253,In_945);
nor U780 (N_780,In_2741,In_511);
nand U781 (N_781,In_2515,In_741);
and U782 (N_782,In_70,In_1111);
xnor U783 (N_783,In_1686,In_2919);
nand U784 (N_784,In_1747,In_476);
or U785 (N_785,In_284,In_2528);
nand U786 (N_786,In_2248,In_1677);
or U787 (N_787,In_952,In_1225);
nand U788 (N_788,In_1588,In_2649);
xor U789 (N_789,In_584,In_369);
nor U790 (N_790,In_2153,In_1150);
nand U791 (N_791,In_936,In_1697);
or U792 (N_792,In_1958,In_1065);
nand U793 (N_793,In_2013,In_1095);
nor U794 (N_794,In_138,In_1718);
nand U795 (N_795,In_1388,In_2752);
xor U796 (N_796,In_2607,In_1089);
nor U797 (N_797,In_290,In_1305);
and U798 (N_798,In_1776,In_1676);
xor U799 (N_799,In_2296,In_702);
xor U800 (N_800,In_1708,In_2781);
nor U801 (N_801,In_2096,In_2117);
xor U802 (N_802,In_135,In_13);
nor U803 (N_803,In_917,In_1149);
xor U804 (N_804,In_1929,In_2018);
xnor U805 (N_805,In_1029,In_2089);
xor U806 (N_806,In_710,In_2716);
xor U807 (N_807,In_1582,In_471);
or U808 (N_808,In_2383,In_2366);
nand U809 (N_809,In_541,In_943);
and U810 (N_810,In_121,In_2348);
nand U811 (N_811,In_2358,In_2812);
and U812 (N_812,In_428,In_406);
xnor U813 (N_813,In_885,In_1311);
and U814 (N_814,In_518,In_2130);
nand U815 (N_815,In_2511,In_2872);
and U816 (N_816,In_2523,In_1188);
or U817 (N_817,In_364,In_612);
nor U818 (N_818,In_311,In_370);
xnor U819 (N_819,In_2412,In_2300);
xnor U820 (N_820,In_157,In_2895);
nor U821 (N_821,In_2936,In_494);
nand U822 (N_822,In_1671,In_2698);
nand U823 (N_823,In_2648,In_2235);
nand U824 (N_824,In_1587,In_2518);
xnor U825 (N_825,In_2643,In_1891);
or U826 (N_826,In_400,In_2047);
or U827 (N_827,In_2974,In_2929);
nor U828 (N_828,In_2918,In_2594);
and U829 (N_829,In_1695,In_1454);
and U830 (N_830,In_350,In_1370);
xor U831 (N_831,In_1816,In_2038);
and U832 (N_832,In_154,In_600);
nand U833 (N_833,In_536,In_2138);
or U834 (N_834,In_2900,In_670);
nand U835 (N_835,In_1446,In_2286);
xnor U836 (N_836,In_2865,In_616);
nor U837 (N_837,In_2282,In_1868);
and U838 (N_838,In_1985,In_1175);
xnor U839 (N_839,In_1634,In_212);
nor U840 (N_840,In_381,In_463);
or U841 (N_841,In_2073,In_2416);
xor U842 (N_842,In_1083,In_1503);
and U843 (N_843,In_2237,In_58);
or U844 (N_844,In_955,In_644);
nor U845 (N_845,In_947,In_1432);
and U846 (N_846,In_1825,In_617);
and U847 (N_847,In_185,In_973);
or U848 (N_848,In_1193,In_1978);
and U849 (N_849,In_1254,In_1315);
nand U850 (N_850,In_1328,In_759);
xnor U851 (N_851,In_1347,In_2769);
nand U852 (N_852,In_1606,In_788);
or U853 (N_853,In_1638,In_117);
and U854 (N_854,In_180,In_1185);
nor U855 (N_855,In_2324,In_1487);
and U856 (N_856,In_1005,In_1576);
and U857 (N_857,In_2887,In_523);
xor U858 (N_858,In_1296,In_2765);
xnor U859 (N_859,In_2137,In_2057);
nand U860 (N_860,In_773,In_845);
nor U861 (N_861,In_2169,In_142);
nand U862 (N_862,In_2660,In_2784);
and U863 (N_863,In_1035,In_2297);
nor U864 (N_864,In_2657,In_1848);
xor U865 (N_865,In_1279,In_15);
nand U866 (N_866,In_2214,In_1463);
nand U867 (N_867,In_1384,In_799);
nand U868 (N_868,In_2933,In_2492);
xnor U869 (N_869,In_2794,In_1486);
xor U870 (N_870,In_1851,In_1527);
or U871 (N_871,In_1824,In_2860);
nand U872 (N_872,In_44,In_2960);
nand U873 (N_873,In_1483,In_1626);
nand U874 (N_874,In_2,In_2188);
nor U875 (N_875,In_1637,In_2804);
nand U876 (N_876,In_695,In_2689);
nor U877 (N_877,In_2241,In_1863);
nor U878 (N_878,In_2761,In_707);
or U879 (N_879,In_2581,In_1294);
nand U880 (N_880,In_1283,In_319);
nand U881 (N_881,In_2932,In_133);
xor U882 (N_882,In_1104,In_1632);
or U883 (N_883,In_1611,In_613);
xnor U884 (N_884,In_304,In_2451);
and U885 (N_885,In_1944,In_1404);
nor U886 (N_886,In_1688,In_2606);
nand U887 (N_887,In_2776,In_2618);
and U888 (N_888,In_2864,In_1426);
and U889 (N_889,In_2453,In_2155);
nand U890 (N_890,In_1163,In_2131);
or U891 (N_891,In_1198,In_2164);
xnor U892 (N_892,In_1585,In_1809);
nor U893 (N_893,In_2084,In_1142);
nor U894 (N_894,In_607,In_2822);
or U895 (N_895,In_3,In_2861);
nor U896 (N_896,In_1161,In_2916);
and U897 (N_897,In_1623,In_1079);
xnor U898 (N_898,In_2279,In_0);
and U899 (N_899,In_1615,In_1475);
xor U900 (N_900,In_1041,In_515);
xnor U901 (N_901,In_2590,In_2981);
xnor U902 (N_902,In_2871,In_2100);
and U903 (N_903,In_2524,In_852);
nand U904 (N_904,In_939,In_1888);
xnor U905 (N_905,In_268,In_2207);
nor U906 (N_906,In_849,In_2371);
and U907 (N_907,In_2793,In_1145);
nor U908 (N_908,In_658,In_1926);
nor U909 (N_909,In_2196,In_2586);
nand U910 (N_910,In_2796,In_2260);
and U911 (N_911,In_2102,In_1178);
nor U912 (N_912,In_1124,In_1542);
and U913 (N_913,In_2460,In_2257);
xnor U914 (N_914,In_2200,In_1221);
or U915 (N_915,In_1011,In_543);
nand U916 (N_916,In_2749,In_1856);
or U917 (N_917,In_83,In_505);
xor U918 (N_918,In_474,In_2536);
nand U919 (N_919,In_2560,In_2737);
or U920 (N_920,In_1586,In_992);
nand U921 (N_921,In_126,In_2201);
nor U922 (N_922,In_2599,In_672);
xor U923 (N_923,In_1003,In_1628);
nand U924 (N_924,In_911,In_581);
nor U925 (N_925,In_730,In_1119);
and U926 (N_926,In_2145,In_2527);
nor U927 (N_927,In_1037,In_1091);
xnor U928 (N_928,In_1389,In_271);
nor U929 (N_929,In_641,In_646);
and U930 (N_930,In_1246,In_2637);
xnor U931 (N_931,In_1131,In_2487);
nand U932 (N_932,In_785,In_1873);
nor U933 (N_933,In_1061,In_980);
nor U934 (N_934,In_597,In_2664);
xnor U935 (N_935,In_1288,In_2623);
and U936 (N_936,In_1949,In_413);
and U937 (N_937,In_315,In_1987);
and U938 (N_938,In_2071,In_1200);
nand U939 (N_939,In_1257,In_2450);
nand U940 (N_940,In_931,In_2563);
or U941 (N_941,In_2529,In_1534);
or U942 (N_942,In_1480,In_2065);
nand U943 (N_943,In_1854,In_2723);
nand U944 (N_944,In_861,In_1413);
or U945 (N_945,In_1405,In_2404);
nor U946 (N_946,In_2572,In_144);
or U947 (N_947,In_925,In_883);
and U948 (N_948,In_2397,In_2953);
xor U949 (N_949,In_1644,In_2271);
and U950 (N_950,In_1860,In_1643);
nand U951 (N_951,In_167,In_2469);
nand U952 (N_952,In_2126,In_342);
nand U953 (N_953,In_1739,In_1180);
nand U954 (N_954,In_1379,In_1435);
nor U955 (N_955,In_426,In_1580);
or U956 (N_956,In_1689,In_219);
and U957 (N_957,In_1815,In_1982);
nor U958 (N_958,In_2224,In_2630);
and U959 (N_959,In_820,In_2639);
nand U960 (N_960,In_1500,In_2230);
or U961 (N_961,In_1445,In_317);
nand U962 (N_962,In_14,In_1190);
and U963 (N_963,In_101,In_438);
xnor U964 (N_964,In_650,In_1087);
xor U965 (N_965,In_1409,In_462);
xor U966 (N_966,In_354,In_1641);
nand U967 (N_967,In_2457,In_933);
nor U968 (N_968,In_2394,In_2510);
nand U969 (N_969,In_2566,In_2335);
xor U970 (N_970,In_1826,In_2496);
xnor U971 (N_971,In_2147,In_2466);
xnor U972 (N_972,In_1781,In_547);
and U973 (N_973,In_491,In_1102);
and U974 (N_974,In_1555,In_1309);
xor U975 (N_975,In_818,In_1556);
or U976 (N_976,In_1055,In_374);
and U977 (N_977,In_300,In_251);
nand U978 (N_978,In_499,In_548);
nor U979 (N_979,In_874,In_934);
and U980 (N_980,In_1849,In_1770);
nor U981 (N_981,In_2375,In_680);
nor U982 (N_982,In_1988,In_2428);
nand U983 (N_983,In_458,In_2447);
or U984 (N_984,In_2909,In_2977);
xnor U985 (N_985,In_1064,In_1790);
nor U986 (N_986,In_2194,In_2033);
and U987 (N_987,In_2414,In_677);
and U988 (N_988,In_332,In_764);
or U989 (N_989,In_1060,In_2381);
and U990 (N_990,In_737,In_2512);
and U991 (N_991,In_1264,In_2233);
or U992 (N_992,In_866,In_1786);
xor U993 (N_993,In_2389,In_1789);
nor U994 (N_994,In_1707,In_522);
xor U995 (N_995,In_331,In_1274);
nand U996 (N_996,In_2674,In_734);
nand U997 (N_997,In_2743,In_490);
and U998 (N_998,In_1914,In_2103);
xor U999 (N_999,In_1026,In_2922);
nand U1000 (N_1000,In_1861,In_2470);
nand U1001 (N_1001,In_2030,In_1681);
nand U1002 (N_1002,In_2659,In_2398);
xor U1003 (N_1003,In_2182,In_429);
nor U1004 (N_1004,In_2963,In_398);
nor U1005 (N_1005,In_2612,In_1137);
xor U1006 (N_1006,In_183,In_1833);
or U1007 (N_1007,In_74,In_2229);
or U1008 (N_1008,In_504,In_2211);
and U1009 (N_1009,In_1932,In_789);
or U1010 (N_1010,In_52,In_686);
nand U1011 (N_1011,In_152,In_365);
nand U1012 (N_1012,In_526,In_765);
xor U1013 (N_1013,In_894,In_2856);
xnor U1014 (N_1014,In_1067,In_250);
or U1015 (N_1015,In_2613,In_906);
nor U1016 (N_1016,In_81,In_1913);
and U1017 (N_1017,In_10,In_1140);
and U1018 (N_1018,In_1963,In_2549);
xor U1019 (N_1019,In_983,In_2677);
or U1020 (N_1020,In_110,In_153);
and U1021 (N_1021,In_1292,In_2314);
and U1022 (N_1022,In_1321,In_802);
nor U1023 (N_1023,In_1673,In_1442);
nor U1024 (N_1024,In_2197,In_2298);
and U1025 (N_1025,In_963,In_692);
xnor U1026 (N_1026,In_2301,In_2449);
and U1027 (N_1027,In_420,In_2333);
xor U1028 (N_1028,In_2884,In_79);
nand U1029 (N_1029,In_396,In_1459);
xnor U1030 (N_1030,In_1631,In_807);
or U1031 (N_1031,In_804,In_873);
and U1032 (N_1032,In_1308,In_2713);
nor U1033 (N_1033,In_238,In_1660);
xor U1034 (N_1034,In_2288,In_1951);
or U1035 (N_1035,In_1602,In_473);
nand U1036 (N_1036,In_235,In_239);
nor U1037 (N_1037,In_2533,In_9);
xnor U1038 (N_1038,In_156,In_1658);
nand U1039 (N_1039,In_1162,In_1152);
nor U1040 (N_1040,In_2539,In_2849);
nand U1041 (N_1041,In_1960,In_2021);
or U1042 (N_1042,In_2760,In_2857);
and U1043 (N_1043,In_218,In_2190);
xor U1044 (N_1044,In_283,In_1918);
and U1045 (N_1045,In_1977,In_329);
or U1046 (N_1046,In_46,In_2014);
or U1047 (N_1047,In_2975,In_1133);
and U1048 (N_1048,In_1046,In_1338);
and U1049 (N_1049,In_639,In_62);
nand U1050 (N_1050,In_352,In_810);
nor U1051 (N_1051,In_969,In_2310);
nor U1052 (N_1052,In_574,In_1619);
or U1053 (N_1053,In_1722,In_1737);
and U1054 (N_1054,In_2423,In_2935);
or U1055 (N_1055,In_762,In_407);
nor U1056 (N_1056,In_93,In_2231);
and U1057 (N_1057,In_1271,In_2610);
and U1058 (N_1058,In_1494,In_2972);
xor U1059 (N_1059,In_2472,In_882);
nor U1060 (N_1060,In_899,In_678);
nor U1061 (N_1061,In_1236,In_1705);
or U1062 (N_1062,In_368,In_2485);
nor U1063 (N_1063,In_2811,In_1508);
xnor U1064 (N_1064,In_2148,In_2978);
xnor U1065 (N_1065,In_1937,In_467);
xnor U1066 (N_1066,In_2085,In_2191);
and U1067 (N_1067,In_299,In_2433);
and U1068 (N_1068,In_327,In_857);
nor U1069 (N_1069,In_2140,In_1622);
nand U1070 (N_1070,In_2750,In_2605);
nand U1071 (N_1071,In_2016,In_682);
and U1072 (N_1072,In_1049,In_1441);
and U1073 (N_1073,In_1383,In_2615);
xnor U1074 (N_1074,In_1165,In_2852);
or U1075 (N_1075,In_45,In_2234);
nor U1076 (N_1076,In_493,In_1081);
xor U1077 (N_1077,In_2088,In_2704);
xnor U1078 (N_1078,In_1524,In_149);
and U1079 (N_1079,In_2320,In_55);
and U1080 (N_1080,In_1829,In_427);
nand U1081 (N_1081,In_2829,In_858);
xnor U1082 (N_1082,In_210,In_43);
xnor U1083 (N_1083,In_1492,In_1159);
nor U1084 (N_1084,In_531,In_2408);
and U1085 (N_1085,In_57,In_151);
nand U1086 (N_1086,In_1233,In_1476);
nand U1087 (N_1087,In_2564,In_1189);
or U1088 (N_1088,In_380,In_1775);
xor U1089 (N_1089,In_27,In_2833);
nor U1090 (N_1090,In_2973,In_2352);
nand U1091 (N_1091,In_2402,In_2172);
nand U1092 (N_1092,In_1923,In_2633);
nor U1093 (N_1093,In_249,In_869);
nand U1094 (N_1094,In_2006,In_1469);
nor U1095 (N_1095,In_556,In_2212);
xnor U1096 (N_1096,In_2876,In_897);
or U1097 (N_1097,In_1640,In_2276);
or U1098 (N_1098,In_1567,In_1760);
or U1099 (N_1099,In_2640,In_2162);
or U1100 (N_1100,In_2179,In_220);
and U1101 (N_1101,In_1572,In_1176);
or U1102 (N_1102,In_667,In_1418);
xor U1103 (N_1103,In_1430,In_642);
and U1104 (N_1104,In_1774,In_2731);
nand U1105 (N_1105,In_2124,In_1344);
or U1106 (N_1106,In_2587,In_587);
xnor U1107 (N_1107,In_26,In_2434);
xnor U1108 (N_1108,In_632,In_971);
or U1109 (N_1109,In_896,In_2859);
nand U1110 (N_1110,In_751,In_308);
or U1111 (N_1111,In_2031,In_1728);
or U1112 (N_1112,In_2265,In_2545);
nand U1113 (N_1113,In_1898,In_578);
and U1114 (N_1114,In_292,In_194);
nand U1115 (N_1115,In_1027,In_1855);
nor U1116 (N_1116,In_888,In_132);
or U1117 (N_1117,In_375,In_2272);
xor U1118 (N_1118,In_1683,In_1045);
or U1119 (N_1119,In_2692,In_2479);
and U1120 (N_1120,In_294,In_2274);
nor U1121 (N_1121,In_821,In_1981);
nand U1122 (N_1122,In_2167,In_1772);
and U1123 (N_1123,In_588,In_532);
nand U1124 (N_1124,In_1168,In_1502);
or U1125 (N_1125,In_1342,In_1558);
and U1126 (N_1126,In_1473,In_1788);
nand U1127 (N_1127,In_1959,In_86);
nand U1128 (N_1128,In_1539,In_2308);
and U1129 (N_1129,In_277,In_2744);
and U1130 (N_1130,In_187,In_2959);
or U1131 (N_1131,In_2382,In_262);
xnor U1132 (N_1132,In_978,In_2195);
xor U1133 (N_1133,In_2701,In_174);
xnor U1134 (N_1134,In_1630,In_1744);
nand U1135 (N_1135,In_908,In_620);
nor U1136 (N_1136,In_2024,In_1260);
nor U1137 (N_1137,In_840,In_164);
nor U1138 (N_1138,In_1945,In_2984);
and U1139 (N_1139,In_2556,In_2459);
or U1140 (N_1140,In_1921,In_221);
nand U1141 (N_1141,In_323,In_1040);
or U1142 (N_1142,In_2983,In_1166);
and U1143 (N_1143,In_1797,In_2093);
nor U1144 (N_1144,In_990,In_2734);
nand U1145 (N_1145,In_456,In_1859);
xor U1146 (N_1146,In_2072,In_1507);
and U1147 (N_1147,In_1050,In_326);
or U1148 (N_1148,In_2903,In_1130);
and U1149 (N_1149,In_1803,In_1117);
nor U1150 (N_1150,In_752,In_823);
or U1151 (N_1151,In_1813,In_1878);
and U1152 (N_1152,In_537,In_2994);
nand U1153 (N_1153,In_2429,In_71);
xor U1154 (N_1154,In_1999,In_1222);
nor U1155 (N_1155,In_602,In_813);
nand U1156 (N_1156,In_870,In_1077);
nand U1157 (N_1157,In_1121,In_2227);
and U1158 (N_1158,In_1039,In_2163);
nor U1159 (N_1159,In_2855,In_405);
nor U1160 (N_1160,In_2544,In_847);
nor U1161 (N_1161,In_2708,In_1422);
or U1162 (N_1162,In_798,In_11);
nand U1163 (N_1163,In_1771,In_1214);
nor U1164 (N_1164,In_394,In_1750);
and U1165 (N_1165,In_391,In_850);
xnor U1166 (N_1166,In_2955,In_953);
or U1167 (N_1167,In_2507,In_32);
or U1168 (N_1168,In_191,In_48);
and U1169 (N_1169,In_959,In_31);
nand U1170 (N_1170,In_674,In_2858);
nand U1171 (N_1171,In_1819,In_2377);
nor U1172 (N_1172,In_1224,In_2968);
xor U1173 (N_1173,In_303,In_2598);
or U1174 (N_1174,In_671,In_662);
and U1175 (N_1175,In_228,In_348);
or U1176 (N_1176,In_1215,In_718);
and U1177 (N_1177,In_35,In_2362);
nor U1178 (N_1178,In_2976,In_184);
nand U1179 (N_1179,In_2505,In_1253);
and U1180 (N_1180,In_1107,In_530);
or U1181 (N_1181,In_2418,In_2624);
nor U1182 (N_1182,In_988,In_1597);
nor U1183 (N_1183,In_1491,In_281);
and U1184 (N_1184,In_1234,In_792);
xor U1185 (N_1185,In_748,In_1974);
nand U1186 (N_1186,In_1814,In_2641);
xor U1187 (N_1187,In_1546,In_1047);
nor U1188 (N_1188,In_1927,In_2926);
or U1189 (N_1189,In_915,In_701);
or U1190 (N_1190,In_704,In_2686);
nor U1191 (N_1191,In_161,In_699);
or U1192 (N_1192,In_2904,In_2908);
and U1193 (N_1193,In_39,In_2896);
or U1194 (N_1194,In_923,In_1916);
nor U1195 (N_1195,In_525,In_2565);
xor U1196 (N_1196,In_1080,In_881);
nand U1197 (N_1197,In_625,In_236);
xor U1198 (N_1198,In_353,In_287);
and U1199 (N_1199,In_213,In_36);
nor U1200 (N_1200,In_1867,In_1666);
xnor U1201 (N_1201,In_2551,In_1485);
or U1202 (N_1202,In_445,In_2008);
or U1203 (N_1203,In_22,In_2573);
or U1204 (N_1204,In_87,In_938);
nand U1205 (N_1205,In_2780,In_1174);
nor U1206 (N_1206,In_2609,In_2361);
or U1207 (N_1207,In_1720,In_2835);
xnor U1208 (N_1208,In_148,In_2577);
or U1209 (N_1209,In_1376,In_1614);
and U1210 (N_1210,In_1519,In_2135);
or U1211 (N_1211,In_962,In_432);
or U1212 (N_1212,In_516,In_2223);
nor U1213 (N_1213,In_758,In_797);
nor U1214 (N_1214,In_2591,In_995);
or U1215 (N_1215,In_99,In_94);
nor U1216 (N_1216,In_1068,In_2989);
or U1217 (N_1217,In_2830,In_1428);
or U1218 (N_1218,In_918,In_2091);
and U1219 (N_1219,In_2121,In_2177);
and U1220 (N_1220,In_1733,In_801);
or U1221 (N_1221,In_2048,In_2517);
nor U1222 (N_1222,In_1536,In_2165);
and U1223 (N_1223,In_1247,In_2754);
nor U1224 (N_1224,In_2558,In_77);
or U1225 (N_1225,In_2106,In_1464);
xor U1226 (N_1226,In_2222,In_878);
or U1227 (N_1227,In_972,In_1905);
nand U1228 (N_1228,In_2690,In_2842);
xor U1229 (N_1229,In_19,In_1948);
nand U1230 (N_1230,In_339,In_844);
or U1231 (N_1231,In_1694,In_652);
xnor U1232 (N_1232,In_285,In_2029);
xnor U1233 (N_1233,In_1909,In_2942);
nor U1234 (N_1234,In_940,In_173);
xor U1235 (N_1235,In_1942,In_1036);
and U1236 (N_1236,In_2087,In_1823);
nor U1237 (N_1237,In_779,In_1925);
and U1238 (N_1238,In_1220,In_517);
and U1239 (N_1239,In_964,In_1610);
xnor U1240 (N_1240,In_698,In_2891);
nor U1241 (N_1241,In_2764,In_1197);
nand U1242 (N_1242,In_514,In_188);
nor U1243 (N_1243,In_1134,In_1256);
xor U1244 (N_1244,In_1700,In_248);
xor U1245 (N_1245,In_1592,In_1962);
or U1246 (N_1246,In_1512,In_1680);
and U1247 (N_1247,In_2067,In_1229);
and U1248 (N_1248,In_498,In_2553);
nor U1249 (N_1249,In_1075,In_2329);
or U1250 (N_1250,In_1574,In_2125);
and U1251 (N_1251,In_749,In_2236);
nor U1252 (N_1252,In_2579,In_839);
nand U1253 (N_1253,In_2011,In_1106);
and U1254 (N_1254,In_2446,In_535);
nand U1255 (N_1255,In_2755,In_382);
or U1256 (N_1256,In_1787,In_1436);
or U1257 (N_1257,In_1804,In_2378);
nor U1258 (N_1258,In_669,In_2502);
xor U1259 (N_1259,In_1835,In_2848);
xnor U1260 (N_1260,In_892,In_2578);
or U1261 (N_1261,In_442,In_648);
or U1262 (N_1262,In_1128,In_2213);
or U1263 (N_1263,In_1876,In_2419);
xnor U1264 (N_1264,In_2493,In_1170);
nor U1265 (N_1265,In_2772,In_2844);
or U1266 (N_1266,In_637,In_1979);
xnor U1267 (N_1267,In_1956,In_619);
xnor U1268 (N_1268,In_1367,In_2246);
nand U1269 (N_1269,In_1211,In_2189);
nor U1270 (N_1270,In_635,In_775);
nand U1271 (N_1271,In_2019,In_1553);
xnor U1272 (N_1272,In_362,In_746);
xnor U1273 (N_1273,In_2305,In_681);
xor U1274 (N_1274,In_1842,In_808);
xnor U1275 (N_1275,In_2318,In_1314);
or U1276 (N_1276,In_744,In_76);
and U1277 (N_1277,In_2768,In_1777);
nand U1278 (N_1278,In_266,In_1569);
and U1279 (N_1279,In_1420,In_1158);
nor U1280 (N_1280,In_1343,In_2083);
nand U1281 (N_1281,In_2948,In_1613);
or U1282 (N_1282,In_1522,In_676);
nand U1283 (N_1283,In_651,In_80);
nor U1284 (N_1284,In_2783,In_1201);
nor U1285 (N_1285,In_2442,In_1092);
or U1286 (N_1286,In_2045,In_2181);
xnor U1287 (N_1287,In_440,In_1153);
or U1288 (N_1288,In_2417,In_528);
and U1289 (N_1289,In_2150,In_2068);
or U1290 (N_1290,In_1518,In_1654);
nor U1291 (N_1291,In_2814,In_2243);
or U1292 (N_1292,In_835,In_2725);
nor U1293 (N_1293,In_1394,In_1382);
nor U1294 (N_1294,In_202,In_689);
or U1295 (N_1295,In_1408,In_1415);
nand U1296 (N_1296,In_544,In_2883);
xor U1297 (N_1297,In_1550,In_755);
xor U1298 (N_1298,In_2049,In_506);
nand U1299 (N_1299,In_2499,In_961);
nor U1300 (N_1300,In_661,In_996);
nor U1301 (N_1301,In_1031,In_1125);
nand U1302 (N_1302,In_2902,In_2312);
or U1303 (N_1303,In_104,In_991);
and U1304 (N_1304,In_2766,In_2115);
and U1305 (N_1305,In_2642,In_747);
xnor U1306 (N_1306,In_2186,In_2431);
and U1307 (N_1307,In_2580,In_2621);
nand U1308 (N_1308,In_2675,In_2726);
nand U1309 (N_1309,In_1778,In_1183);
nor U1310 (N_1310,In_2721,In_253);
nor U1311 (N_1311,In_207,In_2970);
xnor U1312 (N_1312,In_1954,In_1241);
nand U1313 (N_1313,In_2671,In_1832);
or U1314 (N_1314,In_2346,In_2775);
and U1315 (N_1315,In_1212,In_2077);
nor U1316 (N_1316,In_1595,In_663);
nand U1317 (N_1317,In_500,In_201);
and U1318 (N_1318,In_761,In_1411);
nand U1319 (N_1319,In_1655,In_2514);
nor U1320 (N_1320,In_2695,In_1302);
nand U1321 (N_1321,In_312,In_575);
nand U1322 (N_1322,In_2617,In_2092);
nand U1323 (N_1323,In_1575,In_1699);
or U1324 (N_1324,In_424,In_1399);
nand U1325 (N_1325,In_2107,In_2552);
and U1326 (N_1326,In_524,In_56);
and U1327 (N_1327,In_2136,In_2679);
nor U1328 (N_1328,In_1607,In_2054);
and U1329 (N_1329,In_38,In_1523);
and U1330 (N_1330,In_1242,In_63);
and U1331 (N_1331,In_2611,In_1989);
nand U1332 (N_1332,In_691,In_2800);
nor U1333 (N_1333,In_2537,In_1346);
or U1334 (N_1334,In_2950,In_1846);
and U1335 (N_1335,In_1259,In_2410);
nor U1336 (N_1336,In_2178,In_889);
or U1337 (N_1337,In_2142,In_1947);
or U1338 (N_1338,In_1616,In_2906);
nand U1339 (N_1339,In_17,In_2636);
nor U1340 (N_1340,In_920,In_2602);
nor U1341 (N_1341,In_594,In_2489);
nor U1342 (N_1342,In_2575,In_832);
or U1343 (N_1343,In_1726,In_2622);
xor U1344 (N_1344,In_1800,In_2786);
xnor U1345 (N_1345,In_2374,In_833);
nor U1346 (N_1346,In_1243,In_1887);
xnor U1347 (N_1347,In_2526,In_1396);
xnor U1348 (N_1348,In_856,In_1352);
and U1349 (N_1349,In_2748,In_1337);
nor U1350 (N_1350,In_1322,In_750);
nor U1351 (N_1351,In_509,In_1478);
or U1352 (N_1352,In_2474,In_1545);
nor U1353 (N_1353,In_2525,In_1009);
and U1354 (N_1354,In_402,In_1298);
and U1355 (N_1355,In_1601,In_2055);
nor U1356 (N_1356,In_1291,In_2988);
nand U1357 (N_1357,In_1901,In_984);
or U1358 (N_1358,In_932,In_585);
nor U1359 (N_1359,In_2683,In_2875);
or U1360 (N_1360,In_655,In_1911);
xnor U1361 (N_1361,In_2339,In_2986);
nand U1362 (N_1362,In_100,In_1053);
nand U1363 (N_1363,In_2557,In_1753);
nand U1364 (N_1364,In_5,In_2118);
or U1365 (N_1365,In_2042,In_553);
or U1366 (N_1366,In_211,In_1746);
nand U1367 (N_1367,In_2807,In_425);
or U1368 (N_1368,In_373,In_2040);
nor U1369 (N_1369,In_8,In_1144);
and U1370 (N_1370,In_507,In_1340);
nand U1371 (N_1371,In_2332,In_1552);
nand U1372 (N_1372,In_2424,In_603);
or U1373 (N_1373,In_16,In_1997);
and U1374 (N_1374,In_324,In_214);
xor U1375 (N_1375,In_1231,In_2168);
xnor U1376 (N_1376,In_264,In_2266);
nand U1377 (N_1377,In_2571,In_563);
or U1378 (N_1378,In_145,In_146);
nand U1379 (N_1379,In_91,In_2954);
and U1380 (N_1380,In_1557,In_1656);
nand U1381 (N_1381,In_1701,In_2315);
or U1382 (N_1382,In_2885,In_155);
or U1383 (N_1383,In_794,In_389);
nor U1384 (N_1384,In_2530,In_2372);
nand U1385 (N_1385,In_2651,In_726);
xnor U1386 (N_1386,In_2393,In_864);
or U1387 (N_1387,In_877,In_231);
nor U1388 (N_1388,In_1013,In_2802);
xnor U1389 (N_1389,In_876,In_2629);
or U1390 (N_1390,In_1517,In_1907);
or U1391 (N_1391,In_140,In_24);
xor U1392 (N_1392,In_2331,In_1004);
nor U1393 (N_1393,In_1171,In_638);
and U1394 (N_1394,In_1667,In_2729);
nor U1395 (N_1395,In_2500,In_1612);
nand U1396 (N_1396,In_2245,In_1297);
xor U1397 (N_1397,In_763,In_618);
nand U1398 (N_1398,In_1240,In_2696);
and U1399 (N_1399,In_97,In_768);
nand U1400 (N_1400,In_2730,In_433);
nand U1401 (N_1401,In_240,In_2538);
nor U1402 (N_1402,In_1452,In_124);
or U1403 (N_1403,In_1521,In_1836);
xor U1404 (N_1404,In_2205,In_919);
nor U1405 (N_1405,In_2144,In_879);
or U1406 (N_1406,In_2379,In_1);
and U1407 (N_1407,In_1939,In_2838);
and U1408 (N_1408,In_2426,In_385);
or U1409 (N_1409,In_1922,In_2277);
nor U1410 (N_1410,In_2626,In_1063);
xor U1411 (N_1411,In_244,In_1278);
xnor U1412 (N_1412,In_985,In_893);
nor U1413 (N_1413,In_935,In_1094);
xnor U1414 (N_1414,In_2173,In_1749);
and U1415 (N_1415,In_340,In_2034);
or U1416 (N_1416,In_130,In_2703);
and U1417 (N_1417,In_593,In_2477);
and U1418 (N_1418,In_72,In_1757);
nor U1419 (N_1419,In_1076,In_2497);
nand U1420 (N_1420,In_2559,In_435);
and U1421 (N_1421,In_1862,In_736);
or U1422 (N_1422,In_2441,In_306);
xnor U1423 (N_1423,In_753,In_907);
xnor U1424 (N_1424,In_2839,In_2542);
xnor U1425 (N_1425,In_1351,In_610);
and U1426 (N_1426,In_1732,In_2465);
nor U1427 (N_1427,In_2036,In_1535);
nor U1428 (N_1428,In_2939,In_1784);
and U1429 (N_1429,In_2456,In_604);
xor U1430 (N_1430,In_1098,In_1148);
nand U1431 (N_1431,In_1122,In_2897);
or U1432 (N_1432,In_2688,In_1173);
or U1433 (N_1433,In_2225,In_1548);
or U1434 (N_1434,In_1335,In_367);
nand U1435 (N_1435,In_2345,In_1731);
xnor U1436 (N_1436,In_1078,In_37);
xor U1437 (N_1437,In_1525,In_1182);
nor U1438 (N_1438,In_410,In_538);
xor U1439 (N_1439,In_1583,In_1360);
nor U1440 (N_1440,In_2862,In_141);
nand U1441 (N_1441,In_1967,In_2252);
or U1442 (N_1442,In_1090,In_2369);
nand U1443 (N_1443,In_2898,In_2422);
and U1444 (N_1444,In_2653,In_454);
nand U1445 (N_1445,In_2334,In_1593);
xnor U1446 (N_1446,In_387,In_1562);
nand U1447 (N_1447,In_956,In_356);
nor U1448 (N_1448,In_1440,In_115);
or U1449 (N_1449,In_2295,In_1269);
xor U1450 (N_1450,In_1946,In_2183);
or U1451 (N_1451,In_2821,In_376);
nor U1452 (N_1452,In_449,In_1232);
nor U1453 (N_1453,In_1745,In_1000);
and U1454 (N_1454,In_1890,In_412);
or U1455 (N_1455,In_2869,In_1877);
nand U1456 (N_1456,In_2632,In_2385);
xnor U1457 (N_1457,In_2157,In_2059);
nor U1458 (N_1458,In_289,In_2280);
and U1459 (N_1459,In_1709,In_1661);
nor U1460 (N_1460,In_1191,In_696);
or U1461 (N_1461,In_2966,In_1406);
xor U1462 (N_1462,In_1808,In_1363);
or U1463 (N_1463,In_1711,In_1969);
xnor U1464 (N_1464,In_557,In_1465);
nor U1465 (N_1465,In_2943,In_282);
and U1466 (N_1466,In_2669,In_1202);
nand U1467 (N_1467,In_1858,In_1421);
xor U1468 (N_1468,In_322,In_457);
nor U1469 (N_1469,In_2438,In_2401);
nor U1470 (N_1470,In_717,In_2863);
xor U1471 (N_1471,In_2099,In_589);
nand U1472 (N_1472,In_366,In_1565);
or U1473 (N_1473,In_1769,In_502);
and U1474 (N_1474,In_2448,In_192);
xnor U1475 (N_1475,In_550,In_2584);
nor U1476 (N_1476,In_2387,In_1398);
and U1477 (N_1477,In_645,In_999);
and U1478 (N_1478,In_623,In_1401);
nand U1479 (N_1479,In_1339,In_2109);
nand U1480 (N_1480,In_1196,In_836);
and U1481 (N_1481,In_12,In_1252);
xor U1482 (N_1482,In_1443,In_2758);
or U1483 (N_1483,In_770,In_1515);
nand U1484 (N_1484,In_1496,In_1672);
nand U1485 (N_1485,In_2680,In_1362);
nand U1486 (N_1486,In_2139,In_1123);
or U1487 (N_1487,In_1151,In_809);
xnor U1488 (N_1488,In_1598,In_2585);
nand U1489 (N_1489,In_1217,In_1281);
nand U1490 (N_1490,In_1710,In_2709);
nand U1491 (N_1491,In_2464,In_2961);
and U1492 (N_1492,In_2336,In_1617);
and U1493 (N_1493,In_800,In_901);
or U1494 (N_1494,In_653,In_265);
and U1495 (N_1495,In_298,In_2735);
xor U1496 (N_1496,In_2596,In_2715);
nor U1497 (N_1497,In_1838,In_349);
xnor U1498 (N_1498,In_2421,In_1735);
nor U1499 (N_1499,In_1504,In_2023);
nor U1500 (N_1500,N_241,N_118);
and U1501 (N_1501,N_1317,N_542);
or U1502 (N_1502,N_753,N_1030);
nor U1503 (N_1503,N_535,N_874);
nand U1504 (N_1504,N_1250,N_1394);
nor U1505 (N_1505,N_253,N_928);
nor U1506 (N_1506,N_77,N_713);
nand U1507 (N_1507,N_1094,N_1184);
and U1508 (N_1508,N_1160,N_60);
or U1509 (N_1509,N_975,N_992);
or U1510 (N_1510,N_955,N_1011);
xnor U1511 (N_1511,N_1022,N_1149);
or U1512 (N_1512,N_762,N_1358);
and U1513 (N_1513,N_613,N_426);
and U1514 (N_1514,N_1173,N_967);
or U1515 (N_1515,N_1348,N_476);
and U1516 (N_1516,N_312,N_1225);
and U1517 (N_1517,N_353,N_729);
or U1518 (N_1518,N_1479,N_177);
xor U1519 (N_1519,N_149,N_335);
and U1520 (N_1520,N_1486,N_1470);
or U1521 (N_1521,N_442,N_66);
xnor U1522 (N_1522,N_75,N_1362);
nor U1523 (N_1523,N_1034,N_1241);
nand U1524 (N_1524,N_594,N_1027);
or U1525 (N_1525,N_395,N_945);
and U1526 (N_1526,N_962,N_522);
and U1527 (N_1527,N_293,N_1489);
and U1528 (N_1528,N_574,N_742);
nand U1529 (N_1529,N_101,N_1006);
xor U1530 (N_1530,N_1251,N_1180);
nand U1531 (N_1531,N_496,N_1273);
xor U1532 (N_1532,N_451,N_879);
nand U1533 (N_1533,N_1240,N_707);
nor U1534 (N_1534,N_1104,N_1238);
and U1535 (N_1535,N_259,N_1301);
xnor U1536 (N_1536,N_1287,N_759);
nor U1537 (N_1537,N_815,N_144);
or U1538 (N_1538,N_204,N_425);
and U1539 (N_1539,N_1298,N_172);
nor U1540 (N_1540,N_1329,N_937);
nand U1541 (N_1541,N_986,N_1260);
xnor U1542 (N_1542,N_786,N_864);
or U1543 (N_1543,N_927,N_748);
or U1544 (N_1544,N_1336,N_701);
nand U1545 (N_1545,N_637,N_607);
or U1546 (N_1546,N_1320,N_1335);
nand U1547 (N_1547,N_656,N_740);
nand U1548 (N_1548,N_447,N_1477);
nor U1549 (N_1549,N_1130,N_1097);
xor U1550 (N_1550,N_1378,N_1126);
nor U1551 (N_1551,N_205,N_57);
nand U1552 (N_1552,N_325,N_524);
nor U1553 (N_1553,N_378,N_1115);
nor U1554 (N_1554,N_1436,N_723);
nor U1555 (N_1555,N_616,N_124);
xnor U1556 (N_1556,N_208,N_1039);
xnor U1557 (N_1557,N_1171,N_248);
xnor U1558 (N_1558,N_1476,N_844);
nor U1559 (N_1559,N_16,N_1013);
nor U1560 (N_1560,N_1310,N_155);
xor U1561 (N_1561,N_145,N_48);
xnor U1562 (N_1562,N_1031,N_317);
nand U1563 (N_1563,N_941,N_649);
or U1564 (N_1564,N_427,N_338);
xor U1565 (N_1565,N_531,N_1349);
or U1566 (N_1566,N_418,N_318);
nor U1567 (N_1567,N_942,N_777);
nand U1568 (N_1568,N_1129,N_153);
nand U1569 (N_1569,N_190,N_188);
nor U1570 (N_1570,N_421,N_978);
xor U1571 (N_1571,N_345,N_1140);
and U1572 (N_1572,N_509,N_646);
or U1573 (N_1573,N_1437,N_1357);
nor U1574 (N_1574,N_126,N_1272);
or U1575 (N_1575,N_543,N_1478);
xnor U1576 (N_1576,N_904,N_581);
nand U1577 (N_1577,N_552,N_525);
nor U1578 (N_1578,N_1463,N_1131);
nor U1579 (N_1579,N_1262,N_894);
and U1580 (N_1580,N_582,N_1277);
xnor U1581 (N_1581,N_728,N_930);
or U1582 (N_1582,N_592,N_209);
nand U1583 (N_1583,N_40,N_672);
and U1584 (N_1584,N_896,N_1105);
xor U1585 (N_1585,N_946,N_29);
or U1586 (N_1586,N_834,N_1066);
and U1587 (N_1587,N_968,N_1109);
or U1588 (N_1588,N_107,N_796);
nor U1589 (N_1589,N_849,N_749);
and U1590 (N_1590,N_1367,N_1368);
or U1591 (N_1591,N_62,N_711);
or U1592 (N_1592,N_812,N_781);
or U1593 (N_1593,N_1164,N_89);
nor U1594 (N_1594,N_918,N_1050);
and U1595 (N_1595,N_617,N_1435);
xnor U1596 (N_1596,N_985,N_676);
xor U1597 (N_1597,N_1258,N_682);
and U1598 (N_1598,N_1366,N_1386);
nor U1599 (N_1599,N_20,N_726);
xor U1600 (N_1600,N_533,N_792);
nand U1601 (N_1601,N_140,N_595);
and U1602 (N_1602,N_34,N_703);
or U1603 (N_1603,N_498,N_561);
xor U1604 (N_1604,N_911,N_814);
xnor U1605 (N_1605,N_310,N_1061);
nor U1606 (N_1606,N_423,N_1043);
and U1607 (N_1607,N_1497,N_443);
or U1608 (N_1608,N_207,N_169);
nand U1609 (N_1609,N_1350,N_1138);
and U1610 (N_1610,N_1462,N_689);
nand U1611 (N_1611,N_411,N_1452);
nor U1612 (N_1612,N_512,N_341);
or U1613 (N_1613,N_623,N_1237);
xnor U1614 (N_1614,N_388,N_55);
or U1615 (N_1615,N_113,N_1247);
xnor U1616 (N_1616,N_1148,N_1450);
and U1617 (N_1617,N_712,N_836);
xor U1618 (N_1618,N_120,N_1003);
xor U1619 (N_1619,N_467,N_458);
xnor U1620 (N_1620,N_1025,N_1100);
and U1621 (N_1621,N_1224,N_908);
xor U1622 (N_1622,N_839,N_990);
nor U1623 (N_1623,N_575,N_1356);
or U1624 (N_1624,N_755,N_1255);
or U1625 (N_1625,N_269,N_1267);
nand U1626 (N_1626,N_1363,N_56);
xor U1627 (N_1627,N_529,N_1079);
xnor U1628 (N_1628,N_700,N_1323);
and U1629 (N_1629,N_1412,N_1125);
nand U1630 (N_1630,N_604,N_240);
nand U1631 (N_1631,N_731,N_737);
and U1632 (N_1632,N_608,N_891);
nand U1633 (N_1633,N_486,N_1374);
and U1634 (N_1634,N_1454,N_1198);
and U1635 (N_1635,N_1249,N_286);
or U1636 (N_1636,N_494,N_297);
nand U1637 (N_1637,N_1114,N_995);
or U1638 (N_1638,N_1334,N_2);
nand U1639 (N_1639,N_610,N_308);
and U1640 (N_1640,N_633,N_95);
xor U1641 (N_1641,N_501,N_644);
nand U1642 (N_1642,N_1215,N_788);
nor U1643 (N_1643,N_348,N_1226);
or U1644 (N_1644,N_1113,N_1112);
or U1645 (N_1645,N_571,N_1279);
xor U1646 (N_1646,N_1353,N_505);
and U1647 (N_1647,N_733,N_285);
and U1648 (N_1648,N_444,N_277);
nor U1649 (N_1649,N_175,N_1218);
and U1650 (N_1650,N_1417,N_976);
or U1651 (N_1651,N_160,N_958);
or U1652 (N_1652,N_632,N_429);
nand U1653 (N_1653,N_1385,N_5);
or U1654 (N_1654,N_1339,N_117);
nor U1655 (N_1655,N_827,N_994);
nand U1656 (N_1656,N_799,N_299);
nor U1657 (N_1657,N_1341,N_898);
nor U1658 (N_1658,N_566,N_1455);
and U1659 (N_1659,N_1415,N_1338);
xnor U1660 (N_1660,N_944,N_300);
nand U1661 (N_1661,N_634,N_539);
nor U1662 (N_1662,N_273,N_32);
nor U1663 (N_1663,N_9,N_1332);
nor U1664 (N_1664,N_939,N_1046);
nand U1665 (N_1665,N_254,N_226);
nor U1666 (N_1666,N_243,N_1048);
nor U1667 (N_1667,N_1480,N_428);
nor U1668 (N_1668,N_119,N_472);
and U1669 (N_1669,N_282,N_773);
nand U1670 (N_1670,N_1185,N_600);
xnor U1671 (N_1671,N_970,N_1191);
and U1672 (N_1672,N_1005,N_513);
nor U1673 (N_1673,N_885,N_1360);
xor U1674 (N_1674,N_201,N_289);
nand U1675 (N_1675,N_1167,N_1281);
nand U1676 (N_1676,N_1453,N_1364);
nor U1677 (N_1677,N_598,N_123);
nand U1678 (N_1678,N_70,N_459);
and U1679 (N_1679,N_1206,N_1018);
nor U1680 (N_1680,N_1248,N_210);
nor U1681 (N_1681,N_752,N_206);
xnor U1682 (N_1682,N_316,N_841);
nor U1683 (N_1683,N_1159,N_1244);
nor U1684 (N_1684,N_650,N_593);
xor U1685 (N_1685,N_1060,N_1442);
xor U1686 (N_1686,N_18,N_25);
xor U1687 (N_1687,N_1089,N_453);
xor U1688 (N_1688,N_1064,N_419);
nor U1689 (N_1689,N_347,N_1192);
xor U1690 (N_1690,N_806,N_1481);
or U1691 (N_1691,N_1351,N_79);
xor U1692 (N_1692,N_867,N_791);
xnor U1693 (N_1693,N_1395,N_838);
xnor U1694 (N_1694,N_863,N_167);
or U1695 (N_1695,N_1404,N_384);
and U1696 (N_1696,N_342,N_195);
and U1697 (N_1697,N_988,N_1372);
nand U1698 (N_1698,N_1231,N_1441);
and U1699 (N_1699,N_1128,N_197);
and U1700 (N_1700,N_1433,N_407);
and U1701 (N_1701,N_485,N_1195);
nand U1702 (N_1702,N_354,N_1181);
and U1703 (N_1703,N_690,N_191);
and U1704 (N_1704,N_1314,N_871);
nor U1705 (N_1705,N_916,N_949);
and U1706 (N_1706,N_1033,N_1049);
nand U1707 (N_1707,N_54,N_580);
xor U1708 (N_1708,N_638,N_971);
or U1709 (N_1709,N_471,N_1042);
nor U1710 (N_1710,N_374,N_223);
and U1711 (N_1711,N_1299,N_432);
xnor U1712 (N_1712,N_38,N_1228);
and U1713 (N_1713,N_440,N_591);
and U1714 (N_1714,N_1135,N_74);
nor U1715 (N_1715,N_528,N_301);
xnor U1716 (N_1716,N_1210,N_1145);
xor U1717 (N_1717,N_103,N_776);
and U1718 (N_1718,N_653,N_363);
and U1719 (N_1719,N_369,N_902);
nand U1720 (N_1720,N_719,N_1387);
xnor U1721 (N_1721,N_4,N_292);
nor U1722 (N_1722,N_150,N_965);
or U1723 (N_1723,N_115,N_563);
nand U1724 (N_1724,N_10,N_1127);
xor U1725 (N_1725,N_856,N_376);
and U1726 (N_1726,N_540,N_1292);
nand U1727 (N_1727,N_185,N_966);
nand U1728 (N_1728,N_1074,N_1090);
xnor U1729 (N_1729,N_230,N_1254);
and U1730 (N_1730,N_1012,N_659);
nor U1731 (N_1731,N_769,N_714);
or U1732 (N_1732,N_473,N_1425);
and U1733 (N_1733,N_1146,N_387);
and U1734 (N_1734,N_1391,N_502);
nor U1735 (N_1735,N_200,N_1214);
nand U1736 (N_1736,N_417,N_914);
nor U1737 (N_1737,N_640,N_860);
and U1738 (N_1738,N_64,N_1352);
nor U1739 (N_1739,N_984,N_164);
and U1740 (N_1740,N_692,N_431);
nand U1741 (N_1741,N_1133,N_287);
nor U1742 (N_1742,N_1384,N_655);
or U1743 (N_1743,N_1291,N_837);
nand U1744 (N_1744,N_1078,N_754);
nand U1745 (N_1745,N_1439,N_1174);
and U1746 (N_1746,N_961,N_1370);
and U1747 (N_1747,N_42,N_1222);
xor U1748 (N_1748,N_463,N_1359);
xnor U1749 (N_1749,N_702,N_1445);
nand U1750 (N_1750,N_578,N_192);
nor U1751 (N_1751,N_1054,N_324);
or U1752 (N_1752,N_1449,N_541);
nand U1753 (N_1753,N_979,N_379);
or U1754 (N_1754,N_832,N_361);
nand U1755 (N_1755,N_156,N_220);
and U1756 (N_1756,N_104,N_802);
and U1757 (N_1757,N_266,N_323);
nor U1758 (N_1758,N_86,N_59);
or U1759 (N_1759,N_319,N_818);
and U1760 (N_1760,N_1202,N_905);
xnor U1761 (N_1761,N_1156,N_820);
and U1762 (N_1762,N_138,N_861);
xnor U1763 (N_1763,N_482,N_275);
nand U1764 (N_1764,N_1165,N_932);
nand U1765 (N_1765,N_370,N_315);
nor U1766 (N_1766,N_202,N_480);
xor U1767 (N_1767,N_1219,N_217);
nand U1768 (N_1768,N_367,N_1151);
and U1769 (N_1769,N_1408,N_1058);
nor U1770 (N_1770,N_1411,N_1383);
nand U1771 (N_1771,N_495,N_99);
or U1772 (N_1772,N_1253,N_910);
nor U1773 (N_1773,N_267,N_436);
nor U1774 (N_1774,N_35,N_642);
or U1775 (N_1775,N_1398,N_148);
xor U1776 (N_1776,N_404,N_196);
or U1777 (N_1777,N_734,N_412);
nand U1778 (N_1778,N_981,N_461);
and U1779 (N_1779,N_772,N_1313);
xnor U1780 (N_1780,N_356,N_165);
nand U1781 (N_1781,N_565,N_309);
or U1782 (N_1782,N_507,N_105);
nand U1783 (N_1783,N_987,N_1328);
nand U1784 (N_1784,N_194,N_1178);
nand U1785 (N_1785,N_1380,N_621);
and U1786 (N_1786,N_96,N_334);
and U1787 (N_1787,N_390,N_602);
or U1788 (N_1788,N_178,N_705);
and U1789 (N_1789,N_132,N_516);
nor U1790 (N_1790,N_314,N_1234);
and U1791 (N_1791,N_1209,N_199);
or U1792 (N_1792,N_887,N_556);
or U1793 (N_1793,N_61,N_213);
nand U1794 (N_1794,N_147,N_500);
or U1795 (N_1795,N_330,N_1397);
nand U1796 (N_1796,N_569,N_557);
xnor U1797 (N_1797,N_215,N_1289);
and U1798 (N_1798,N_398,N_969);
and U1799 (N_1799,N_1008,N_1492);
xnor U1800 (N_1800,N_784,N_294);
and U1801 (N_1801,N_562,N_506);
nor U1802 (N_1802,N_1403,N_758);
and U1803 (N_1803,N_1423,N_280);
nor U1804 (N_1804,N_1170,N_295);
nand U1805 (N_1805,N_1306,N_605);
nor U1806 (N_1806,N_250,N_527);
or U1807 (N_1807,N_1426,N_953);
or U1808 (N_1808,N_1321,N_738);
nor U1809 (N_1809,N_1242,N_1302);
and U1810 (N_1810,N_373,N_44);
nand U1811 (N_1811,N_1396,N_1278);
nor U1812 (N_1812,N_892,N_1296);
or U1813 (N_1813,N_679,N_1169);
nor U1814 (N_1814,N_671,N_1459);
or U1815 (N_1815,N_337,N_151);
nand U1816 (N_1816,N_1498,N_249);
nand U1817 (N_1817,N_15,N_350);
nor U1818 (N_1818,N_234,N_1246);
or U1819 (N_1819,N_1261,N_17);
or U1820 (N_1820,N_783,N_1312);
nor U1821 (N_1821,N_380,N_1045);
or U1822 (N_1822,N_183,N_232);
nand U1823 (N_1823,N_227,N_365);
or U1824 (N_1824,N_1158,N_1051);
nand U1825 (N_1825,N_851,N_678);
xnor U1826 (N_1826,N_710,N_597);
nor U1827 (N_1827,N_478,N_1154);
xor U1828 (N_1828,N_1065,N_554);
xnor U1829 (N_1829,N_1482,N_998);
nor U1830 (N_1830,N_52,N_116);
nand U1831 (N_1831,N_1085,N_1121);
or U1832 (N_1832,N_1490,N_567);
or U1833 (N_1833,N_816,N_750);
nand U1834 (N_1834,N_1020,N_639);
nand U1835 (N_1835,N_222,N_745);
and U1836 (N_1836,N_635,N_619);
nand U1837 (N_1837,N_1091,N_782);
or U1838 (N_1838,N_715,N_828);
xor U1839 (N_1839,N_1457,N_601);
nor U1840 (N_1840,N_789,N_694);
and U1841 (N_1841,N_6,N_654);
and U1842 (N_1842,N_1239,N_1421);
nand U1843 (N_1843,N_238,N_304);
nor U1844 (N_1844,N_1168,N_1438);
nor U1845 (N_1845,N_1132,N_19);
xor U1846 (N_1846,N_811,N_1311);
nor U1847 (N_1847,N_848,N_795);
and U1848 (N_1848,N_677,N_893);
nand U1849 (N_1849,N_1179,N_1389);
nor U1850 (N_1850,N_808,N_1252);
or U1851 (N_1851,N_1266,N_801);
xor U1852 (N_1852,N_357,N_673);
xnor U1853 (N_1853,N_331,N_550);
or U1854 (N_1854,N_835,N_1354);
nor U1855 (N_1855,N_258,N_947);
nand U1856 (N_1856,N_903,N_184);
xor U1857 (N_1857,N_876,N_27);
and U1858 (N_1858,N_276,N_1136);
xor U1859 (N_1859,N_143,N_1371);
or U1860 (N_1860,N_1276,N_724);
or U1861 (N_1861,N_1137,N_1208);
and U1862 (N_1862,N_1496,N_313);
nand U1863 (N_1863,N_1203,N_173);
or U1864 (N_1864,N_433,N_765);
nand U1865 (N_1865,N_1468,N_161);
and U1866 (N_1866,N_957,N_408);
nor U1867 (N_1867,N_1036,N_950);
and U1868 (N_1868,N_687,N_880);
and U1869 (N_1869,N_780,N_465);
or U1870 (N_1870,N_667,N_492);
xnor U1871 (N_1871,N_198,N_171);
and U1872 (N_1872,N_1162,N_68);
nand U1873 (N_1873,N_1422,N_1183);
and U1874 (N_1874,N_954,N_993);
nand U1875 (N_1875,N_1243,N_850);
or U1876 (N_1876,N_1193,N_570);
nor U1877 (N_1877,N_127,N_274);
nor U1878 (N_1878,N_1429,N_503);
xor U1879 (N_1879,N_1080,N_133);
or U1880 (N_1880,N_872,N_328);
nor U1881 (N_1881,N_706,N_430);
xor U1882 (N_1882,N_870,N_611);
xor U1883 (N_1883,N_446,N_1283);
xnor U1884 (N_1884,N_1344,N_1333);
nand U1885 (N_1885,N_721,N_1432);
nand U1886 (N_1886,N_1297,N_383);
nand U1887 (N_1887,N_920,N_479);
nor U1888 (N_1888,N_926,N_1274);
xor U1889 (N_1889,N_1290,N_154);
or U1890 (N_1890,N_997,N_1014);
or U1891 (N_1891,N_1393,N_329);
xor U1892 (N_1892,N_278,N_1245);
xnor U1893 (N_1893,N_1414,N_523);
nand U1894 (N_1894,N_1001,N_1176);
and U1895 (N_1895,N_858,N_100);
nor U1896 (N_1896,N_1285,N_493);
nand U1897 (N_1897,N_1155,N_1);
nand U1898 (N_1898,N_0,N_3);
xnor U1899 (N_1899,N_1232,N_84);
or U1900 (N_1900,N_521,N_270);
nand U1901 (N_1901,N_810,N_1229);
nand U1902 (N_1902,N_691,N_321);
or U1903 (N_1903,N_544,N_1216);
and U1904 (N_1904,N_49,N_257);
nand U1905 (N_1905,N_1392,N_53);
and U1906 (N_1906,N_51,N_1293);
xnor U1907 (N_1907,N_1377,N_1163);
nand U1908 (N_1908,N_628,N_80);
xor U1909 (N_1909,N_71,N_1032);
and U1910 (N_1910,N_1139,N_1120);
nor U1911 (N_1911,N_651,N_76);
nand U1912 (N_1912,N_389,N_1053);
and U1913 (N_1913,N_1002,N_1447);
nand U1914 (N_1914,N_555,N_170);
xor U1915 (N_1915,N_211,N_716);
xor U1916 (N_1916,N_262,N_730);
nor U1917 (N_1917,N_1147,N_212);
and U1918 (N_1918,N_1217,N_739);
and U1919 (N_1919,N_125,N_663);
or U1920 (N_1920,N_193,N_1373);
xor U1921 (N_1921,N_1300,N_406);
nor U1922 (N_1922,N_375,N_751);
and U1923 (N_1923,N_332,N_807);
nand U1924 (N_1924,N_797,N_1271);
nor U1925 (N_1925,N_265,N_233);
nand U1926 (N_1926,N_1111,N_366);
nor U1927 (N_1927,N_1092,N_372);
xnor U1928 (N_1928,N_1021,N_824);
and U1929 (N_1929,N_1355,N_746);
nor U1930 (N_1930,N_551,N_973);
nor U1931 (N_1931,N_481,N_470);
nand U1932 (N_1932,N_1223,N_821);
nand U1933 (N_1933,N_307,N_359);
xnor U1934 (N_1934,N_1399,N_1375);
and U1935 (N_1935,N_514,N_1390);
or U1936 (N_1936,N_888,N_627);
xor U1937 (N_1937,N_587,N_386);
nand U1938 (N_1938,N_362,N_1213);
nor U1939 (N_1939,N_1081,N_434);
and U1940 (N_1940,N_722,N_1010);
or U1941 (N_1941,N_1177,N_727);
or U1942 (N_1942,N_1117,N_1190);
and U1943 (N_1943,N_1466,N_237);
nor U1944 (N_1944,N_596,N_1052);
and U1945 (N_1945,N_163,N_272);
or U1946 (N_1946,N_1007,N_1026);
nor U1947 (N_1947,N_424,N_519);
xor U1948 (N_1948,N_239,N_686);
and U1949 (N_1949,N_474,N_940);
and U1950 (N_1950,N_1485,N_878);
nor U1951 (N_1951,N_203,N_588);
xnor U1952 (N_1952,N_92,N_320);
xnor U1953 (N_1953,N_983,N_515);
nor U1954 (N_1954,N_186,N_800);
nor U1955 (N_1955,N_1294,N_684);
and U1956 (N_1956,N_558,N_311);
and U1957 (N_1957,N_283,N_112);
xor U1958 (N_1958,N_688,N_1096);
nand U1959 (N_1959,N_1047,N_1221);
nand U1960 (N_1960,N_1345,N_852);
xnor U1961 (N_1961,N_111,N_744);
nand U1962 (N_1962,N_1326,N_162);
and U1963 (N_1963,N_825,N_895);
or U1964 (N_1964,N_182,N_302);
xor U1965 (N_1965,N_402,N_549);
or U1966 (N_1966,N_1077,N_831);
nor U1967 (N_1967,N_798,N_405);
and U1968 (N_1968,N_1400,N_819);
or U1969 (N_1969,N_959,N_271);
and U1970 (N_1970,N_855,N_674);
nor U1971 (N_1971,N_1330,N_108);
or U1972 (N_1972,N_1166,N_483);
nand U1973 (N_1973,N_26,N_382);
nor U1974 (N_1974,N_564,N_648);
nand U1975 (N_1975,N_1465,N_268);
and U1976 (N_1976,N_909,N_131);
and U1977 (N_1977,N_935,N_951);
xnor U1978 (N_1978,N_1424,N_1016);
xor U1979 (N_1979,N_747,N_787);
xor U1980 (N_1980,N_464,N_736);
and U1981 (N_1981,N_83,N_245);
or U1982 (N_1982,N_768,N_845);
nand U1983 (N_1983,N_881,N_397);
nor U1984 (N_1984,N_39,N_33);
or U1985 (N_1985,N_1172,N_1444);
nand U1986 (N_1986,N_1056,N_360);
or U1987 (N_1987,N_1134,N_774);
nor U1988 (N_1988,N_189,N_1106);
nor U1989 (N_1989,N_877,N_530);
xor U1990 (N_1990,N_1309,N_1388);
nand U1991 (N_1991,N_82,N_1075);
and U1992 (N_1992,N_899,N_862);
nor U1993 (N_1993,N_847,N_794);
and U1994 (N_1994,N_1458,N_288);
nand U1995 (N_1995,N_1153,N_214);
or U1996 (N_1996,N_460,N_1263);
xnor U1997 (N_1997,N_1495,N_518);
nand U1998 (N_1998,N_1024,N_1028);
nor U1999 (N_1999,N_583,N_1009);
or U2000 (N_2000,N_1443,N_1175);
or U2001 (N_2001,N_445,N_261);
or U2002 (N_2002,N_437,N_603);
and U2003 (N_2003,N_683,N_146);
nand U2004 (N_2004,N_449,N_438);
and U2005 (N_2005,N_1446,N_826);
and U2006 (N_2006,N_526,N_219);
xor U2007 (N_2007,N_469,N_906);
nor U2008 (N_2008,N_883,N_303);
and U2009 (N_2009,N_1275,N_1376);
or U2010 (N_2010,N_14,N_882);
and U2011 (N_2011,N_129,N_696);
or U2012 (N_2012,N_590,N_1324);
and U2013 (N_2013,N_1083,N_181);
and U2014 (N_2014,N_47,N_1406);
and U2015 (N_2015,N_1227,N_1282);
nor U2016 (N_2016,N_252,N_1337);
and U2017 (N_2017,N_1040,N_924);
xnor U2018 (N_2018,N_484,N_913);
or U2019 (N_2019,N_1063,N_218);
nand U2020 (N_2020,N_1123,N_999);
or U2021 (N_2021,N_804,N_128);
nor U2022 (N_2022,N_65,N_381);
and U2023 (N_2023,N_1088,N_657);
nor U2024 (N_2024,N_612,N_1035);
nand U2025 (N_2025,N_573,N_536);
xor U2026 (N_2026,N_1304,N_58);
and U2027 (N_2027,N_718,N_1110);
xnor U2028 (N_2028,N_658,N_1315);
and U2029 (N_2029,N_1182,N_532);
and U2030 (N_2030,N_391,N_73);
and U2031 (N_2031,N_256,N_560);
and U2032 (N_2032,N_615,N_1460);
nand U2033 (N_2033,N_790,N_956);
nand U2034 (N_2034,N_842,N_1379);
and U2035 (N_2035,N_698,N_624);
xor U2036 (N_2036,N_93,N_545);
nor U2037 (N_2037,N_306,N_487);
and U2038 (N_2038,N_251,N_1087);
or U2039 (N_2039,N_1144,N_422);
or U2040 (N_2040,N_1093,N_629);
or U2041 (N_2041,N_1331,N_1086);
xor U2042 (N_2042,N_901,N_385);
nor U2043 (N_2043,N_1044,N_697);
nand U2044 (N_2044,N_1230,N_168);
nand U2045 (N_2045,N_989,N_344);
nor U2046 (N_2046,N_43,N_22);
or U2047 (N_2047,N_670,N_546);
and U2048 (N_2048,N_1196,N_1409);
and U2049 (N_2049,N_122,N_255);
or U2050 (N_2050,N_537,N_1322);
nor U2051 (N_2051,N_817,N_187);
nor U2052 (N_2052,N_139,N_85);
or U2053 (N_2053,N_1142,N_645);
nor U2054 (N_2054,N_685,N_890);
nand U2055 (N_2055,N_1098,N_853);
nor U2056 (N_2056,N_933,N_392);
xnor U2057 (N_2057,N_606,N_977);
nor U2058 (N_2058,N_599,N_441);
and U2059 (N_2059,N_641,N_110);
xnor U2060 (N_2060,N_72,N_1431);
xnor U2061 (N_2061,N_900,N_456);
xnor U2062 (N_2062,N_450,N_1471);
nor U2063 (N_2063,N_36,N_912);
and U2064 (N_2064,N_1286,N_1019);
xnor U2065 (N_2065,N_1101,N_489);
nor U2066 (N_2066,N_964,N_413);
nand U2067 (N_2067,N_517,N_1316);
nor U2068 (N_2068,N_1150,N_829);
xor U2069 (N_2069,N_343,N_349);
or U2070 (N_2070,N_1259,N_336);
or U2071 (N_2071,N_1430,N_371);
nand U2072 (N_2072,N_1119,N_1467);
xnor U2073 (N_2073,N_520,N_1082);
xnor U2074 (N_2074,N_1070,N_875);
nand U2075 (N_2075,N_1197,N_873);
nor U2076 (N_2076,N_1122,N_1141);
xor U2077 (N_2077,N_410,N_771);
or U2078 (N_2078,N_843,N_298);
or U2079 (N_2079,N_180,N_630);
and U2080 (N_2080,N_106,N_680);
and U2081 (N_2081,N_1186,N_7);
xnor U2082 (N_2082,N_1475,N_770);
and U2083 (N_2083,N_1211,N_457);
or U2084 (N_2084,N_510,N_1201);
and U2085 (N_2085,N_377,N_823);
or U2086 (N_2086,N_63,N_1000);
nand U2087 (N_2087,N_358,N_1493);
xnor U2088 (N_2088,N_246,N_720);
and U2089 (N_2089,N_1418,N_717);
nand U2090 (N_2090,N_403,N_236);
and U2091 (N_2091,N_866,N_704);
xor U2092 (N_2092,N_466,N_547);
and U2093 (N_2093,N_1451,N_228);
nor U2094 (N_2094,N_247,N_693);
nand U2095 (N_2095,N_1305,N_568);
xor U2096 (N_2096,N_936,N_622);
or U2097 (N_2097,N_631,N_1095);
nor U2098 (N_2098,N_1108,N_1303);
nand U2099 (N_2099,N_109,N_1199);
and U2100 (N_2100,N_416,N_1401);
nand U2101 (N_2101,N_1416,N_1038);
nand U2102 (N_2102,N_1057,N_508);
xor U2103 (N_2103,N_1143,N_1469);
xor U2104 (N_2104,N_1084,N_1188);
nand U2105 (N_2105,N_1235,N_263);
or U2106 (N_2106,N_454,N_589);
xnor U2107 (N_2107,N_553,N_1236);
xor U2108 (N_2108,N_559,N_1340);
and U2109 (N_2109,N_869,N_1161);
nor U2110 (N_2110,N_1488,N_91);
nand U2111 (N_2111,N_69,N_322);
or U2112 (N_2112,N_1308,N_1073);
nor U2113 (N_2113,N_158,N_668);
xnor U2114 (N_2114,N_468,N_760);
or U2115 (N_2115,N_1346,N_577);
and U2116 (N_2116,N_1410,N_757);
and U2117 (N_2117,N_785,N_934);
and U2118 (N_2118,N_333,N_735);
or U2119 (N_2119,N_1365,N_114);
nand U2120 (N_2120,N_1343,N_579);
nor U2121 (N_2121,N_1076,N_1037);
xor U2122 (N_2122,N_778,N_216);
xnor U2123 (N_2123,N_538,N_121);
and U2124 (N_2124,N_339,N_1212);
and U2125 (N_2125,N_1270,N_488);
and U2126 (N_2126,N_660,N_960);
xnor U2127 (N_2127,N_709,N_399);
nor U2128 (N_2128,N_1288,N_290);
nand U2129 (N_2129,N_625,N_1280);
and U2130 (N_2130,N_779,N_50);
xor U2131 (N_2131,N_766,N_665);
nand U2132 (N_2132,N_1407,N_974);
nand U2133 (N_2133,N_435,N_1023);
nor U2134 (N_2134,N_857,N_346);
nor U2135 (N_2135,N_504,N_1307);
nand U2136 (N_2136,N_452,N_647);
or U2137 (N_2137,N_166,N_279);
or U2138 (N_2138,N_732,N_938);
nand U2139 (N_2139,N_1472,N_401);
nand U2140 (N_2140,N_499,N_1420);
or U2141 (N_2141,N_221,N_41);
nand U2142 (N_2142,N_865,N_136);
nor U2143 (N_2143,N_1062,N_284);
xnor U2144 (N_2144,N_699,N_1059);
or U2145 (N_2145,N_364,N_1072);
xor U2146 (N_2146,N_1152,N_305);
or U2147 (N_2147,N_925,N_982);
nor U2148 (N_2148,N_907,N_97);
and U2149 (N_2149,N_130,N_1405);
or U2150 (N_2150,N_1067,N_142);
xor U2151 (N_2151,N_840,N_393);
nor U2152 (N_2152,N_917,N_420);
xnor U2153 (N_2153,N_805,N_1499);
nor U2154 (N_2154,N_152,N_490);
xnor U2155 (N_2155,N_37,N_1069);
or U2156 (N_2156,N_1118,N_1456);
nor U2157 (N_2157,N_1194,N_475);
xor U2158 (N_2158,N_681,N_244);
nor U2159 (N_2159,N_134,N_1318);
xor U2160 (N_2160,N_756,N_643);
nand U2161 (N_2161,N_830,N_11);
xnor U2162 (N_2162,N_8,N_1204);
and U2163 (N_2163,N_963,N_1464);
xnor U2164 (N_2164,N_548,N_1256);
xnor U2165 (N_2165,N_235,N_919);
xnor U2166 (N_2166,N_921,N_922);
nand U2167 (N_2167,N_368,N_30);
nor U2168 (N_2168,N_67,N_224);
nor U2169 (N_2169,N_854,N_929);
nand U2170 (N_2170,N_396,N_260);
or U2171 (N_2171,N_1448,N_1319);
or U2172 (N_2172,N_1071,N_1369);
xor U2173 (N_2173,N_135,N_897);
and U2174 (N_2174,N_620,N_31);
nand U2175 (N_2175,N_1284,N_1015);
or U2176 (N_2176,N_618,N_491);
nand U2177 (N_2177,N_1116,N_1347);
nor U2178 (N_2178,N_415,N_586);
nand U2179 (N_2179,N_1428,N_179);
or U2180 (N_2180,N_1157,N_943);
nand U2181 (N_2181,N_102,N_94);
nor U2182 (N_2182,N_1107,N_439);
or U2183 (N_2183,N_242,N_455);
xor U2184 (N_2184,N_28,N_23);
and U2185 (N_2185,N_340,N_229);
and U2186 (N_2186,N_813,N_1402);
or U2187 (N_2187,N_1200,N_352);
and U2188 (N_2188,N_88,N_1427);
xnor U2189 (N_2189,N_1483,N_803);
nor U2190 (N_2190,N_174,N_1189);
xor U2191 (N_2191,N_394,N_1434);
nand U2192 (N_2192,N_1041,N_980);
xor U2193 (N_2193,N_355,N_81);
nand U2194 (N_2194,N_1102,N_675);
xnor U2195 (N_2195,N_666,N_972);
nor U2196 (N_2196,N_763,N_326);
nor U2197 (N_2197,N_1327,N_1361);
nand U2198 (N_2198,N_327,N_351);
nand U2199 (N_2199,N_846,N_477);
and U2200 (N_2200,N_1207,N_626);
nand U2201 (N_2201,N_1461,N_884);
and U2202 (N_2202,N_609,N_511);
or U2203 (N_2203,N_996,N_725);
and U2204 (N_2204,N_78,N_761);
or U2205 (N_2205,N_793,N_1068);
nor U2206 (N_2206,N_1491,N_90);
xor U2207 (N_2207,N_1325,N_1103);
or U2208 (N_2208,N_1268,N_572);
xor U2209 (N_2209,N_176,N_1265);
and U2210 (N_2210,N_661,N_1099);
xor U2211 (N_2211,N_1381,N_1473);
xnor U2212 (N_2212,N_889,N_931);
xnor U2213 (N_2213,N_87,N_886);
nand U2214 (N_2214,N_296,N_1124);
nor U2215 (N_2215,N_157,N_822);
nor U2216 (N_2216,N_1257,N_24);
nand U2217 (N_2217,N_585,N_915);
xnor U2218 (N_2218,N_1295,N_1187);
xnor U2219 (N_2219,N_409,N_98);
xor U2220 (N_2220,N_1494,N_1220);
nand U2221 (N_2221,N_833,N_1029);
nor U2222 (N_2222,N_137,N_448);
and U2223 (N_2223,N_534,N_497);
nor U2224 (N_2224,N_614,N_1004);
and U2225 (N_2225,N_809,N_1264);
xnor U2226 (N_2226,N_400,N_743);
and U2227 (N_2227,N_1413,N_708);
xnor U2228 (N_2228,N_281,N_12);
and U2229 (N_2229,N_576,N_1055);
and U2230 (N_2230,N_664,N_991);
or U2231 (N_2231,N_231,N_1484);
nor U2232 (N_2232,N_1342,N_948);
and U2233 (N_2233,N_1474,N_868);
xnor U2234 (N_2234,N_159,N_952);
and U2235 (N_2235,N_767,N_462);
and U2236 (N_2236,N_1487,N_45);
and U2237 (N_2237,N_264,N_1382);
nor U2238 (N_2238,N_141,N_584);
nand U2239 (N_2239,N_21,N_652);
nor U2240 (N_2240,N_13,N_225);
and U2241 (N_2241,N_669,N_1419);
xor U2242 (N_2242,N_695,N_741);
xnor U2243 (N_2243,N_923,N_859);
nor U2244 (N_2244,N_764,N_1440);
and U2245 (N_2245,N_1017,N_662);
nor U2246 (N_2246,N_291,N_775);
nor U2247 (N_2247,N_46,N_1205);
xnor U2248 (N_2248,N_1269,N_414);
xnor U2249 (N_2249,N_636,N_1233);
and U2250 (N_2250,N_462,N_958);
and U2251 (N_2251,N_1160,N_730);
or U2252 (N_2252,N_1165,N_558);
and U2253 (N_2253,N_1143,N_361);
nor U2254 (N_2254,N_726,N_305);
nor U2255 (N_2255,N_529,N_111);
xor U2256 (N_2256,N_243,N_1392);
nand U2257 (N_2257,N_396,N_471);
nor U2258 (N_2258,N_505,N_121);
or U2259 (N_2259,N_1400,N_1168);
or U2260 (N_2260,N_918,N_419);
xor U2261 (N_2261,N_1075,N_305);
nand U2262 (N_2262,N_261,N_806);
xor U2263 (N_2263,N_97,N_879);
and U2264 (N_2264,N_1010,N_479);
and U2265 (N_2265,N_210,N_332);
or U2266 (N_2266,N_524,N_1119);
nand U2267 (N_2267,N_467,N_79);
xor U2268 (N_2268,N_1494,N_1332);
nand U2269 (N_2269,N_1419,N_1220);
and U2270 (N_2270,N_269,N_540);
nor U2271 (N_2271,N_529,N_1186);
and U2272 (N_2272,N_335,N_915);
nor U2273 (N_2273,N_1266,N_1288);
or U2274 (N_2274,N_21,N_687);
nor U2275 (N_2275,N_415,N_1049);
and U2276 (N_2276,N_520,N_929);
xor U2277 (N_2277,N_1074,N_1108);
nand U2278 (N_2278,N_1213,N_769);
xor U2279 (N_2279,N_1290,N_1379);
and U2280 (N_2280,N_287,N_282);
and U2281 (N_2281,N_797,N_293);
nand U2282 (N_2282,N_716,N_1359);
nor U2283 (N_2283,N_612,N_327);
nand U2284 (N_2284,N_1469,N_1061);
nand U2285 (N_2285,N_580,N_921);
nor U2286 (N_2286,N_1480,N_567);
and U2287 (N_2287,N_228,N_1379);
nor U2288 (N_2288,N_1044,N_141);
xor U2289 (N_2289,N_213,N_719);
xor U2290 (N_2290,N_1000,N_673);
nor U2291 (N_2291,N_1421,N_680);
or U2292 (N_2292,N_581,N_1140);
xor U2293 (N_2293,N_616,N_805);
nand U2294 (N_2294,N_177,N_831);
nand U2295 (N_2295,N_247,N_1284);
nor U2296 (N_2296,N_386,N_243);
nand U2297 (N_2297,N_131,N_161);
or U2298 (N_2298,N_1310,N_474);
nand U2299 (N_2299,N_1040,N_472);
xor U2300 (N_2300,N_1117,N_526);
nand U2301 (N_2301,N_1450,N_228);
nor U2302 (N_2302,N_827,N_655);
nor U2303 (N_2303,N_309,N_885);
nand U2304 (N_2304,N_1100,N_1283);
and U2305 (N_2305,N_1298,N_58);
or U2306 (N_2306,N_511,N_658);
or U2307 (N_2307,N_343,N_539);
and U2308 (N_2308,N_149,N_1428);
and U2309 (N_2309,N_744,N_97);
xnor U2310 (N_2310,N_699,N_705);
nand U2311 (N_2311,N_104,N_501);
or U2312 (N_2312,N_377,N_1280);
nor U2313 (N_2313,N_1087,N_764);
nand U2314 (N_2314,N_817,N_945);
nand U2315 (N_2315,N_644,N_972);
or U2316 (N_2316,N_1372,N_1128);
nor U2317 (N_2317,N_707,N_1004);
or U2318 (N_2318,N_732,N_1339);
nor U2319 (N_2319,N_405,N_568);
xnor U2320 (N_2320,N_1072,N_718);
nand U2321 (N_2321,N_1183,N_1280);
nor U2322 (N_2322,N_10,N_1448);
and U2323 (N_2323,N_9,N_278);
or U2324 (N_2324,N_643,N_895);
nor U2325 (N_2325,N_447,N_829);
nand U2326 (N_2326,N_34,N_692);
and U2327 (N_2327,N_349,N_18);
xor U2328 (N_2328,N_1299,N_910);
and U2329 (N_2329,N_611,N_1405);
or U2330 (N_2330,N_1159,N_122);
nand U2331 (N_2331,N_2,N_1320);
or U2332 (N_2332,N_1345,N_1399);
nand U2333 (N_2333,N_707,N_52);
nor U2334 (N_2334,N_1491,N_181);
nor U2335 (N_2335,N_1399,N_1);
nand U2336 (N_2336,N_600,N_1420);
nor U2337 (N_2337,N_1432,N_1282);
and U2338 (N_2338,N_718,N_617);
and U2339 (N_2339,N_401,N_271);
nand U2340 (N_2340,N_1220,N_942);
or U2341 (N_2341,N_1497,N_57);
and U2342 (N_2342,N_1312,N_849);
nand U2343 (N_2343,N_1036,N_108);
nand U2344 (N_2344,N_180,N_354);
and U2345 (N_2345,N_1237,N_1358);
nor U2346 (N_2346,N_76,N_1210);
nor U2347 (N_2347,N_330,N_485);
and U2348 (N_2348,N_576,N_1370);
and U2349 (N_2349,N_1279,N_1085);
and U2350 (N_2350,N_1208,N_535);
nand U2351 (N_2351,N_173,N_263);
or U2352 (N_2352,N_137,N_1387);
nor U2353 (N_2353,N_1481,N_77);
or U2354 (N_2354,N_1400,N_35);
and U2355 (N_2355,N_1381,N_206);
and U2356 (N_2356,N_137,N_558);
nand U2357 (N_2357,N_27,N_1111);
xor U2358 (N_2358,N_357,N_891);
nand U2359 (N_2359,N_1227,N_1344);
nand U2360 (N_2360,N_798,N_521);
xnor U2361 (N_2361,N_1459,N_1260);
nor U2362 (N_2362,N_254,N_1472);
and U2363 (N_2363,N_981,N_1032);
xor U2364 (N_2364,N_1319,N_1085);
xor U2365 (N_2365,N_904,N_1205);
nand U2366 (N_2366,N_523,N_342);
nor U2367 (N_2367,N_1462,N_916);
or U2368 (N_2368,N_1412,N_1189);
nand U2369 (N_2369,N_742,N_1256);
xor U2370 (N_2370,N_744,N_1387);
and U2371 (N_2371,N_1263,N_624);
xnor U2372 (N_2372,N_967,N_355);
or U2373 (N_2373,N_872,N_1237);
nand U2374 (N_2374,N_328,N_443);
nand U2375 (N_2375,N_569,N_1464);
and U2376 (N_2376,N_1183,N_949);
nand U2377 (N_2377,N_329,N_87);
or U2378 (N_2378,N_466,N_639);
nor U2379 (N_2379,N_224,N_294);
and U2380 (N_2380,N_1220,N_634);
xor U2381 (N_2381,N_1445,N_860);
or U2382 (N_2382,N_1197,N_339);
xor U2383 (N_2383,N_964,N_496);
nand U2384 (N_2384,N_1474,N_1450);
and U2385 (N_2385,N_439,N_290);
nand U2386 (N_2386,N_687,N_387);
or U2387 (N_2387,N_1194,N_705);
nor U2388 (N_2388,N_411,N_988);
or U2389 (N_2389,N_841,N_1138);
xnor U2390 (N_2390,N_991,N_510);
xor U2391 (N_2391,N_1101,N_668);
or U2392 (N_2392,N_1009,N_915);
xor U2393 (N_2393,N_1116,N_1284);
nor U2394 (N_2394,N_156,N_207);
and U2395 (N_2395,N_1336,N_653);
xnor U2396 (N_2396,N_1183,N_860);
nor U2397 (N_2397,N_183,N_777);
nor U2398 (N_2398,N_1373,N_101);
or U2399 (N_2399,N_1341,N_1133);
xnor U2400 (N_2400,N_1333,N_1289);
and U2401 (N_2401,N_157,N_1223);
and U2402 (N_2402,N_1310,N_197);
xnor U2403 (N_2403,N_1318,N_471);
nor U2404 (N_2404,N_1450,N_1132);
nand U2405 (N_2405,N_87,N_1224);
and U2406 (N_2406,N_1402,N_829);
xnor U2407 (N_2407,N_1130,N_1312);
xnor U2408 (N_2408,N_1434,N_108);
nand U2409 (N_2409,N_246,N_1287);
and U2410 (N_2410,N_306,N_80);
nor U2411 (N_2411,N_59,N_204);
xnor U2412 (N_2412,N_795,N_435);
nor U2413 (N_2413,N_290,N_970);
or U2414 (N_2414,N_446,N_1154);
xnor U2415 (N_2415,N_1101,N_294);
nor U2416 (N_2416,N_647,N_507);
nand U2417 (N_2417,N_472,N_1454);
or U2418 (N_2418,N_41,N_1026);
xor U2419 (N_2419,N_1111,N_272);
xor U2420 (N_2420,N_1269,N_1175);
and U2421 (N_2421,N_1410,N_269);
nor U2422 (N_2422,N_1284,N_1039);
or U2423 (N_2423,N_1353,N_78);
and U2424 (N_2424,N_747,N_1027);
or U2425 (N_2425,N_946,N_1482);
nor U2426 (N_2426,N_752,N_1303);
or U2427 (N_2427,N_1113,N_228);
nor U2428 (N_2428,N_92,N_1496);
nor U2429 (N_2429,N_613,N_120);
or U2430 (N_2430,N_1208,N_868);
and U2431 (N_2431,N_501,N_1234);
and U2432 (N_2432,N_234,N_738);
xor U2433 (N_2433,N_705,N_66);
xor U2434 (N_2434,N_589,N_476);
nand U2435 (N_2435,N_277,N_536);
and U2436 (N_2436,N_1118,N_201);
xor U2437 (N_2437,N_1067,N_1288);
and U2438 (N_2438,N_935,N_767);
nor U2439 (N_2439,N_1248,N_485);
and U2440 (N_2440,N_1274,N_901);
nor U2441 (N_2441,N_60,N_1139);
nand U2442 (N_2442,N_1357,N_212);
and U2443 (N_2443,N_975,N_476);
nand U2444 (N_2444,N_671,N_808);
nor U2445 (N_2445,N_988,N_727);
nor U2446 (N_2446,N_185,N_1038);
xnor U2447 (N_2447,N_338,N_1420);
or U2448 (N_2448,N_1419,N_1125);
nor U2449 (N_2449,N_640,N_678);
and U2450 (N_2450,N_1113,N_759);
nand U2451 (N_2451,N_889,N_605);
xor U2452 (N_2452,N_1081,N_1304);
nor U2453 (N_2453,N_863,N_585);
nand U2454 (N_2454,N_927,N_988);
xor U2455 (N_2455,N_875,N_1225);
or U2456 (N_2456,N_627,N_596);
and U2457 (N_2457,N_1162,N_212);
nor U2458 (N_2458,N_722,N_362);
or U2459 (N_2459,N_796,N_88);
nand U2460 (N_2460,N_861,N_1131);
or U2461 (N_2461,N_1058,N_1327);
or U2462 (N_2462,N_71,N_1198);
and U2463 (N_2463,N_142,N_71);
nand U2464 (N_2464,N_273,N_292);
and U2465 (N_2465,N_1009,N_75);
xor U2466 (N_2466,N_261,N_177);
xnor U2467 (N_2467,N_884,N_1127);
and U2468 (N_2468,N_23,N_140);
or U2469 (N_2469,N_69,N_1271);
nor U2470 (N_2470,N_162,N_580);
nor U2471 (N_2471,N_464,N_350);
xnor U2472 (N_2472,N_977,N_204);
and U2473 (N_2473,N_254,N_1371);
or U2474 (N_2474,N_572,N_1429);
nor U2475 (N_2475,N_1100,N_783);
or U2476 (N_2476,N_1241,N_1300);
nand U2477 (N_2477,N_702,N_658);
or U2478 (N_2478,N_267,N_516);
nand U2479 (N_2479,N_951,N_1304);
nand U2480 (N_2480,N_820,N_947);
xor U2481 (N_2481,N_525,N_1385);
nor U2482 (N_2482,N_878,N_475);
or U2483 (N_2483,N_1168,N_267);
nand U2484 (N_2484,N_1471,N_1039);
nor U2485 (N_2485,N_1311,N_1392);
xor U2486 (N_2486,N_1177,N_869);
xor U2487 (N_2487,N_1231,N_1470);
nor U2488 (N_2488,N_1417,N_258);
xor U2489 (N_2489,N_1144,N_973);
and U2490 (N_2490,N_1239,N_524);
or U2491 (N_2491,N_1047,N_842);
or U2492 (N_2492,N_1222,N_1459);
and U2493 (N_2493,N_221,N_1445);
and U2494 (N_2494,N_456,N_731);
xnor U2495 (N_2495,N_1118,N_386);
and U2496 (N_2496,N_1061,N_948);
or U2497 (N_2497,N_940,N_760);
and U2498 (N_2498,N_805,N_410);
or U2499 (N_2499,N_467,N_1056);
and U2500 (N_2500,N_127,N_1319);
or U2501 (N_2501,N_1221,N_884);
xnor U2502 (N_2502,N_747,N_1442);
nand U2503 (N_2503,N_1424,N_640);
nor U2504 (N_2504,N_236,N_510);
or U2505 (N_2505,N_989,N_1090);
or U2506 (N_2506,N_35,N_376);
and U2507 (N_2507,N_588,N_1018);
nor U2508 (N_2508,N_142,N_1121);
and U2509 (N_2509,N_1316,N_728);
or U2510 (N_2510,N_1426,N_127);
nand U2511 (N_2511,N_445,N_921);
xor U2512 (N_2512,N_373,N_722);
nor U2513 (N_2513,N_129,N_870);
xor U2514 (N_2514,N_328,N_807);
nor U2515 (N_2515,N_376,N_668);
and U2516 (N_2516,N_770,N_781);
nand U2517 (N_2517,N_573,N_219);
nand U2518 (N_2518,N_754,N_541);
xor U2519 (N_2519,N_816,N_291);
nor U2520 (N_2520,N_1270,N_106);
nand U2521 (N_2521,N_1118,N_1077);
or U2522 (N_2522,N_287,N_554);
and U2523 (N_2523,N_1279,N_850);
nand U2524 (N_2524,N_889,N_62);
nand U2525 (N_2525,N_898,N_604);
xor U2526 (N_2526,N_466,N_836);
and U2527 (N_2527,N_155,N_859);
nand U2528 (N_2528,N_561,N_283);
xnor U2529 (N_2529,N_1386,N_960);
or U2530 (N_2530,N_22,N_72);
or U2531 (N_2531,N_277,N_1003);
xnor U2532 (N_2532,N_758,N_914);
xor U2533 (N_2533,N_43,N_375);
or U2534 (N_2534,N_298,N_1318);
and U2535 (N_2535,N_1017,N_1182);
nand U2536 (N_2536,N_1336,N_1209);
or U2537 (N_2537,N_1471,N_1282);
nand U2538 (N_2538,N_1015,N_1);
and U2539 (N_2539,N_139,N_1047);
or U2540 (N_2540,N_1275,N_464);
and U2541 (N_2541,N_943,N_115);
and U2542 (N_2542,N_453,N_1154);
and U2543 (N_2543,N_133,N_1215);
nand U2544 (N_2544,N_527,N_603);
nor U2545 (N_2545,N_1052,N_1453);
nand U2546 (N_2546,N_529,N_721);
and U2547 (N_2547,N_1457,N_549);
and U2548 (N_2548,N_1141,N_1420);
and U2549 (N_2549,N_831,N_842);
nor U2550 (N_2550,N_828,N_1028);
nand U2551 (N_2551,N_1330,N_1313);
nand U2552 (N_2552,N_1385,N_53);
nor U2553 (N_2553,N_1334,N_358);
nor U2554 (N_2554,N_1462,N_175);
or U2555 (N_2555,N_1174,N_1138);
nand U2556 (N_2556,N_391,N_105);
or U2557 (N_2557,N_640,N_527);
and U2558 (N_2558,N_1359,N_386);
and U2559 (N_2559,N_1117,N_11);
nor U2560 (N_2560,N_948,N_1382);
nor U2561 (N_2561,N_282,N_322);
nand U2562 (N_2562,N_1102,N_1459);
and U2563 (N_2563,N_529,N_1060);
nor U2564 (N_2564,N_374,N_1250);
nor U2565 (N_2565,N_760,N_847);
nor U2566 (N_2566,N_876,N_1195);
and U2567 (N_2567,N_705,N_782);
or U2568 (N_2568,N_1104,N_599);
or U2569 (N_2569,N_989,N_748);
or U2570 (N_2570,N_1475,N_72);
nor U2571 (N_2571,N_1203,N_1135);
nand U2572 (N_2572,N_1094,N_1290);
or U2573 (N_2573,N_501,N_536);
or U2574 (N_2574,N_968,N_47);
and U2575 (N_2575,N_1412,N_524);
and U2576 (N_2576,N_969,N_1060);
and U2577 (N_2577,N_1055,N_629);
xnor U2578 (N_2578,N_1270,N_187);
nor U2579 (N_2579,N_742,N_1115);
nor U2580 (N_2580,N_310,N_868);
and U2581 (N_2581,N_808,N_938);
or U2582 (N_2582,N_910,N_890);
nor U2583 (N_2583,N_150,N_226);
nor U2584 (N_2584,N_352,N_0);
or U2585 (N_2585,N_1322,N_611);
nand U2586 (N_2586,N_1052,N_744);
nand U2587 (N_2587,N_821,N_1304);
nor U2588 (N_2588,N_1125,N_1338);
nor U2589 (N_2589,N_299,N_232);
and U2590 (N_2590,N_1281,N_1138);
nand U2591 (N_2591,N_1263,N_478);
xnor U2592 (N_2592,N_1361,N_566);
and U2593 (N_2593,N_1460,N_429);
nor U2594 (N_2594,N_1263,N_559);
or U2595 (N_2595,N_1466,N_34);
and U2596 (N_2596,N_760,N_569);
nor U2597 (N_2597,N_1198,N_888);
or U2598 (N_2598,N_948,N_548);
or U2599 (N_2599,N_1381,N_733);
nand U2600 (N_2600,N_629,N_1491);
nand U2601 (N_2601,N_1426,N_838);
and U2602 (N_2602,N_1404,N_1364);
nor U2603 (N_2603,N_1277,N_1233);
nand U2604 (N_2604,N_838,N_88);
and U2605 (N_2605,N_1368,N_971);
nand U2606 (N_2606,N_1356,N_538);
nand U2607 (N_2607,N_1221,N_27);
or U2608 (N_2608,N_864,N_1245);
or U2609 (N_2609,N_125,N_1141);
or U2610 (N_2610,N_5,N_336);
nand U2611 (N_2611,N_1055,N_624);
or U2612 (N_2612,N_263,N_217);
or U2613 (N_2613,N_22,N_941);
xor U2614 (N_2614,N_1198,N_430);
and U2615 (N_2615,N_38,N_541);
nand U2616 (N_2616,N_1174,N_932);
nand U2617 (N_2617,N_1399,N_529);
nor U2618 (N_2618,N_741,N_1258);
nand U2619 (N_2619,N_1058,N_155);
and U2620 (N_2620,N_365,N_1284);
nand U2621 (N_2621,N_466,N_1429);
or U2622 (N_2622,N_431,N_881);
nor U2623 (N_2623,N_1037,N_953);
and U2624 (N_2624,N_1448,N_585);
and U2625 (N_2625,N_151,N_1046);
nor U2626 (N_2626,N_1488,N_1172);
xor U2627 (N_2627,N_398,N_123);
xnor U2628 (N_2628,N_502,N_895);
nor U2629 (N_2629,N_375,N_454);
or U2630 (N_2630,N_1182,N_1400);
and U2631 (N_2631,N_794,N_1456);
or U2632 (N_2632,N_714,N_59);
and U2633 (N_2633,N_904,N_795);
xor U2634 (N_2634,N_739,N_1454);
nand U2635 (N_2635,N_195,N_773);
nor U2636 (N_2636,N_720,N_775);
and U2637 (N_2637,N_79,N_1336);
nor U2638 (N_2638,N_19,N_1274);
or U2639 (N_2639,N_1284,N_525);
or U2640 (N_2640,N_104,N_202);
or U2641 (N_2641,N_886,N_1347);
nor U2642 (N_2642,N_1152,N_661);
nor U2643 (N_2643,N_1442,N_346);
and U2644 (N_2644,N_1452,N_1080);
or U2645 (N_2645,N_1483,N_40);
and U2646 (N_2646,N_831,N_61);
and U2647 (N_2647,N_318,N_591);
xor U2648 (N_2648,N_103,N_803);
nor U2649 (N_2649,N_1237,N_1019);
or U2650 (N_2650,N_1039,N_975);
nand U2651 (N_2651,N_386,N_865);
xor U2652 (N_2652,N_1000,N_1010);
or U2653 (N_2653,N_725,N_493);
or U2654 (N_2654,N_780,N_594);
nand U2655 (N_2655,N_378,N_1483);
nor U2656 (N_2656,N_1207,N_1169);
xnor U2657 (N_2657,N_747,N_758);
nand U2658 (N_2658,N_492,N_1219);
nor U2659 (N_2659,N_365,N_805);
nand U2660 (N_2660,N_640,N_1261);
nand U2661 (N_2661,N_912,N_623);
or U2662 (N_2662,N_1032,N_213);
nor U2663 (N_2663,N_1438,N_843);
nand U2664 (N_2664,N_1229,N_1465);
xor U2665 (N_2665,N_757,N_224);
nor U2666 (N_2666,N_521,N_1028);
nand U2667 (N_2667,N_1321,N_249);
nor U2668 (N_2668,N_113,N_283);
and U2669 (N_2669,N_240,N_1392);
xor U2670 (N_2670,N_1359,N_702);
or U2671 (N_2671,N_1240,N_1480);
nor U2672 (N_2672,N_584,N_753);
and U2673 (N_2673,N_378,N_1206);
and U2674 (N_2674,N_57,N_453);
or U2675 (N_2675,N_492,N_1105);
nor U2676 (N_2676,N_807,N_225);
and U2677 (N_2677,N_909,N_1144);
xor U2678 (N_2678,N_669,N_5);
and U2679 (N_2679,N_536,N_1362);
xnor U2680 (N_2680,N_247,N_422);
nor U2681 (N_2681,N_545,N_920);
xnor U2682 (N_2682,N_1182,N_1415);
nand U2683 (N_2683,N_405,N_1192);
nor U2684 (N_2684,N_1396,N_1191);
and U2685 (N_2685,N_982,N_182);
nand U2686 (N_2686,N_1027,N_66);
nand U2687 (N_2687,N_21,N_1042);
nor U2688 (N_2688,N_1004,N_577);
xor U2689 (N_2689,N_1119,N_203);
or U2690 (N_2690,N_1358,N_278);
nor U2691 (N_2691,N_366,N_1067);
or U2692 (N_2692,N_1032,N_452);
nand U2693 (N_2693,N_773,N_166);
nand U2694 (N_2694,N_1336,N_771);
nor U2695 (N_2695,N_1268,N_946);
and U2696 (N_2696,N_750,N_1451);
nor U2697 (N_2697,N_215,N_764);
nor U2698 (N_2698,N_307,N_1414);
and U2699 (N_2699,N_1394,N_1042);
or U2700 (N_2700,N_510,N_813);
nand U2701 (N_2701,N_658,N_505);
or U2702 (N_2702,N_412,N_1247);
nor U2703 (N_2703,N_1135,N_866);
nand U2704 (N_2704,N_1127,N_1187);
nor U2705 (N_2705,N_1384,N_529);
and U2706 (N_2706,N_440,N_249);
or U2707 (N_2707,N_1207,N_1264);
nor U2708 (N_2708,N_402,N_972);
and U2709 (N_2709,N_576,N_1173);
or U2710 (N_2710,N_1214,N_697);
or U2711 (N_2711,N_1073,N_391);
and U2712 (N_2712,N_518,N_979);
nand U2713 (N_2713,N_899,N_898);
nor U2714 (N_2714,N_1269,N_1023);
and U2715 (N_2715,N_1318,N_1213);
nor U2716 (N_2716,N_28,N_846);
nand U2717 (N_2717,N_1196,N_970);
nand U2718 (N_2718,N_1389,N_720);
nand U2719 (N_2719,N_1017,N_428);
nand U2720 (N_2720,N_1182,N_915);
and U2721 (N_2721,N_360,N_280);
and U2722 (N_2722,N_707,N_300);
xor U2723 (N_2723,N_947,N_299);
xor U2724 (N_2724,N_931,N_1480);
or U2725 (N_2725,N_1121,N_1285);
nand U2726 (N_2726,N_496,N_641);
and U2727 (N_2727,N_398,N_587);
xor U2728 (N_2728,N_128,N_419);
nand U2729 (N_2729,N_22,N_135);
xor U2730 (N_2730,N_261,N_915);
xnor U2731 (N_2731,N_673,N_108);
or U2732 (N_2732,N_852,N_669);
nand U2733 (N_2733,N_548,N_702);
nand U2734 (N_2734,N_1436,N_1483);
nand U2735 (N_2735,N_900,N_299);
nor U2736 (N_2736,N_1216,N_1334);
or U2737 (N_2737,N_1206,N_181);
xor U2738 (N_2738,N_1369,N_508);
nor U2739 (N_2739,N_623,N_821);
xor U2740 (N_2740,N_561,N_584);
xnor U2741 (N_2741,N_1432,N_1116);
and U2742 (N_2742,N_1387,N_392);
nor U2743 (N_2743,N_301,N_1401);
xnor U2744 (N_2744,N_1403,N_241);
nor U2745 (N_2745,N_527,N_738);
and U2746 (N_2746,N_1214,N_1077);
and U2747 (N_2747,N_477,N_435);
nor U2748 (N_2748,N_1078,N_708);
nand U2749 (N_2749,N_30,N_1434);
nor U2750 (N_2750,N_1267,N_1055);
xor U2751 (N_2751,N_892,N_834);
nor U2752 (N_2752,N_931,N_1183);
nor U2753 (N_2753,N_962,N_625);
nor U2754 (N_2754,N_1466,N_802);
nor U2755 (N_2755,N_1358,N_440);
or U2756 (N_2756,N_787,N_1308);
nor U2757 (N_2757,N_372,N_826);
xor U2758 (N_2758,N_1343,N_1165);
nand U2759 (N_2759,N_1267,N_581);
or U2760 (N_2760,N_846,N_472);
and U2761 (N_2761,N_940,N_813);
nand U2762 (N_2762,N_231,N_1458);
xnor U2763 (N_2763,N_132,N_1081);
or U2764 (N_2764,N_154,N_394);
and U2765 (N_2765,N_1149,N_1477);
and U2766 (N_2766,N_670,N_1166);
nor U2767 (N_2767,N_1122,N_521);
nor U2768 (N_2768,N_79,N_1139);
xnor U2769 (N_2769,N_343,N_1100);
xnor U2770 (N_2770,N_1430,N_1243);
nor U2771 (N_2771,N_1102,N_1020);
xor U2772 (N_2772,N_1354,N_1318);
or U2773 (N_2773,N_99,N_1189);
nor U2774 (N_2774,N_1351,N_290);
nor U2775 (N_2775,N_925,N_619);
nand U2776 (N_2776,N_1247,N_1303);
or U2777 (N_2777,N_1185,N_257);
nor U2778 (N_2778,N_1343,N_1366);
xnor U2779 (N_2779,N_621,N_1070);
xnor U2780 (N_2780,N_954,N_958);
nand U2781 (N_2781,N_267,N_284);
xor U2782 (N_2782,N_291,N_104);
or U2783 (N_2783,N_321,N_639);
or U2784 (N_2784,N_1078,N_283);
and U2785 (N_2785,N_38,N_914);
nand U2786 (N_2786,N_156,N_841);
nor U2787 (N_2787,N_393,N_1098);
or U2788 (N_2788,N_938,N_1222);
nor U2789 (N_2789,N_815,N_1293);
or U2790 (N_2790,N_1285,N_1333);
nor U2791 (N_2791,N_829,N_963);
or U2792 (N_2792,N_1162,N_208);
xnor U2793 (N_2793,N_803,N_1149);
xor U2794 (N_2794,N_1399,N_841);
and U2795 (N_2795,N_873,N_1416);
xnor U2796 (N_2796,N_372,N_183);
xor U2797 (N_2797,N_1334,N_1355);
nor U2798 (N_2798,N_165,N_777);
nor U2799 (N_2799,N_1063,N_780);
and U2800 (N_2800,N_1132,N_1479);
xor U2801 (N_2801,N_858,N_1152);
and U2802 (N_2802,N_1035,N_867);
xnor U2803 (N_2803,N_57,N_68);
and U2804 (N_2804,N_5,N_367);
xor U2805 (N_2805,N_706,N_296);
or U2806 (N_2806,N_870,N_1397);
and U2807 (N_2807,N_560,N_946);
nand U2808 (N_2808,N_1008,N_370);
xor U2809 (N_2809,N_443,N_706);
nor U2810 (N_2810,N_1161,N_47);
nor U2811 (N_2811,N_902,N_852);
xor U2812 (N_2812,N_89,N_463);
or U2813 (N_2813,N_928,N_759);
nor U2814 (N_2814,N_1450,N_616);
and U2815 (N_2815,N_183,N_219);
or U2816 (N_2816,N_367,N_1035);
and U2817 (N_2817,N_734,N_1106);
nand U2818 (N_2818,N_920,N_1086);
nor U2819 (N_2819,N_819,N_157);
nand U2820 (N_2820,N_853,N_1194);
or U2821 (N_2821,N_835,N_1160);
xnor U2822 (N_2822,N_930,N_1230);
nor U2823 (N_2823,N_1388,N_586);
and U2824 (N_2824,N_68,N_849);
or U2825 (N_2825,N_655,N_1251);
nand U2826 (N_2826,N_1338,N_301);
or U2827 (N_2827,N_713,N_1337);
or U2828 (N_2828,N_1182,N_465);
nor U2829 (N_2829,N_1452,N_372);
xor U2830 (N_2830,N_1161,N_314);
and U2831 (N_2831,N_1458,N_657);
nor U2832 (N_2832,N_33,N_1337);
and U2833 (N_2833,N_872,N_616);
nand U2834 (N_2834,N_1254,N_770);
or U2835 (N_2835,N_1215,N_708);
and U2836 (N_2836,N_561,N_658);
nor U2837 (N_2837,N_935,N_401);
and U2838 (N_2838,N_1117,N_1332);
and U2839 (N_2839,N_1316,N_534);
and U2840 (N_2840,N_493,N_850);
nand U2841 (N_2841,N_146,N_1382);
nand U2842 (N_2842,N_42,N_1038);
nand U2843 (N_2843,N_1069,N_28);
xor U2844 (N_2844,N_1344,N_821);
and U2845 (N_2845,N_751,N_129);
and U2846 (N_2846,N_234,N_1099);
and U2847 (N_2847,N_1492,N_224);
xnor U2848 (N_2848,N_1454,N_1029);
xnor U2849 (N_2849,N_1144,N_656);
nor U2850 (N_2850,N_777,N_337);
nor U2851 (N_2851,N_1382,N_827);
nor U2852 (N_2852,N_53,N_655);
and U2853 (N_2853,N_567,N_1023);
nor U2854 (N_2854,N_816,N_1258);
xnor U2855 (N_2855,N_968,N_18);
or U2856 (N_2856,N_595,N_593);
or U2857 (N_2857,N_263,N_378);
nand U2858 (N_2858,N_403,N_165);
nand U2859 (N_2859,N_657,N_1014);
and U2860 (N_2860,N_873,N_798);
or U2861 (N_2861,N_556,N_309);
and U2862 (N_2862,N_202,N_374);
and U2863 (N_2863,N_874,N_1234);
or U2864 (N_2864,N_1191,N_603);
or U2865 (N_2865,N_1246,N_1142);
nor U2866 (N_2866,N_375,N_69);
nand U2867 (N_2867,N_809,N_389);
and U2868 (N_2868,N_62,N_1023);
and U2869 (N_2869,N_478,N_368);
or U2870 (N_2870,N_747,N_1318);
and U2871 (N_2871,N_110,N_1288);
xnor U2872 (N_2872,N_762,N_1495);
xnor U2873 (N_2873,N_397,N_889);
and U2874 (N_2874,N_793,N_1486);
nand U2875 (N_2875,N_404,N_498);
and U2876 (N_2876,N_1450,N_538);
xnor U2877 (N_2877,N_908,N_525);
nor U2878 (N_2878,N_1483,N_546);
and U2879 (N_2879,N_369,N_667);
nor U2880 (N_2880,N_467,N_190);
and U2881 (N_2881,N_135,N_1382);
and U2882 (N_2882,N_726,N_146);
nor U2883 (N_2883,N_1097,N_401);
xnor U2884 (N_2884,N_193,N_1258);
nor U2885 (N_2885,N_363,N_100);
or U2886 (N_2886,N_298,N_230);
nor U2887 (N_2887,N_898,N_1199);
nand U2888 (N_2888,N_189,N_71);
nor U2889 (N_2889,N_1069,N_1097);
nand U2890 (N_2890,N_1017,N_210);
or U2891 (N_2891,N_1460,N_495);
nand U2892 (N_2892,N_203,N_633);
xor U2893 (N_2893,N_132,N_651);
and U2894 (N_2894,N_710,N_857);
and U2895 (N_2895,N_1292,N_1181);
xor U2896 (N_2896,N_749,N_14);
nor U2897 (N_2897,N_1072,N_1160);
nand U2898 (N_2898,N_1411,N_247);
nand U2899 (N_2899,N_1056,N_950);
nand U2900 (N_2900,N_1289,N_445);
xnor U2901 (N_2901,N_156,N_353);
or U2902 (N_2902,N_254,N_816);
or U2903 (N_2903,N_182,N_1001);
nor U2904 (N_2904,N_772,N_654);
xor U2905 (N_2905,N_1158,N_36);
nor U2906 (N_2906,N_1482,N_1037);
nor U2907 (N_2907,N_383,N_61);
or U2908 (N_2908,N_770,N_272);
or U2909 (N_2909,N_243,N_1059);
and U2910 (N_2910,N_329,N_952);
nand U2911 (N_2911,N_464,N_864);
nand U2912 (N_2912,N_956,N_1361);
or U2913 (N_2913,N_1098,N_1416);
xor U2914 (N_2914,N_1283,N_263);
xnor U2915 (N_2915,N_267,N_1420);
nor U2916 (N_2916,N_475,N_487);
nor U2917 (N_2917,N_278,N_1417);
nand U2918 (N_2918,N_949,N_1415);
xor U2919 (N_2919,N_881,N_1488);
nand U2920 (N_2920,N_200,N_1495);
nor U2921 (N_2921,N_423,N_685);
nor U2922 (N_2922,N_241,N_852);
or U2923 (N_2923,N_966,N_220);
and U2924 (N_2924,N_1279,N_917);
or U2925 (N_2925,N_1348,N_528);
nand U2926 (N_2926,N_67,N_312);
or U2927 (N_2927,N_410,N_1024);
nand U2928 (N_2928,N_1285,N_560);
or U2929 (N_2929,N_839,N_1274);
nand U2930 (N_2930,N_1219,N_818);
xnor U2931 (N_2931,N_77,N_1178);
xnor U2932 (N_2932,N_531,N_964);
or U2933 (N_2933,N_1271,N_1083);
nand U2934 (N_2934,N_1251,N_922);
xnor U2935 (N_2935,N_569,N_70);
or U2936 (N_2936,N_1336,N_1000);
nor U2937 (N_2937,N_666,N_1422);
nor U2938 (N_2938,N_392,N_394);
or U2939 (N_2939,N_55,N_374);
nand U2940 (N_2940,N_879,N_1254);
xnor U2941 (N_2941,N_474,N_1160);
xor U2942 (N_2942,N_474,N_1120);
or U2943 (N_2943,N_877,N_371);
xor U2944 (N_2944,N_785,N_345);
or U2945 (N_2945,N_370,N_56);
and U2946 (N_2946,N_599,N_857);
or U2947 (N_2947,N_971,N_482);
xor U2948 (N_2948,N_134,N_903);
nor U2949 (N_2949,N_557,N_881);
nand U2950 (N_2950,N_191,N_628);
and U2951 (N_2951,N_1453,N_1232);
nor U2952 (N_2952,N_722,N_196);
nand U2953 (N_2953,N_949,N_548);
and U2954 (N_2954,N_429,N_1345);
or U2955 (N_2955,N_1160,N_419);
or U2956 (N_2956,N_829,N_962);
xnor U2957 (N_2957,N_615,N_717);
nand U2958 (N_2958,N_408,N_30);
nor U2959 (N_2959,N_498,N_1400);
and U2960 (N_2960,N_465,N_316);
and U2961 (N_2961,N_471,N_807);
and U2962 (N_2962,N_1090,N_52);
or U2963 (N_2963,N_465,N_987);
nor U2964 (N_2964,N_1316,N_1454);
nand U2965 (N_2965,N_1299,N_1362);
xnor U2966 (N_2966,N_1111,N_282);
and U2967 (N_2967,N_1163,N_444);
nand U2968 (N_2968,N_1302,N_1225);
and U2969 (N_2969,N_579,N_590);
nand U2970 (N_2970,N_1490,N_876);
xnor U2971 (N_2971,N_596,N_536);
or U2972 (N_2972,N_883,N_649);
or U2973 (N_2973,N_1412,N_687);
xor U2974 (N_2974,N_1323,N_1116);
and U2975 (N_2975,N_1403,N_523);
and U2976 (N_2976,N_66,N_1457);
or U2977 (N_2977,N_557,N_843);
and U2978 (N_2978,N_874,N_21);
nand U2979 (N_2979,N_780,N_38);
nand U2980 (N_2980,N_627,N_54);
or U2981 (N_2981,N_1028,N_600);
nand U2982 (N_2982,N_661,N_309);
nor U2983 (N_2983,N_1021,N_1197);
and U2984 (N_2984,N_1278,N_1320);
nand U2985 (N_2985,N_39,N_416);
nand U2986 (N_2986,N_1180,N_682);
and U2987 (N_2987,N_1229,N_356);
nor U2988 (N_2988,N_336,N_1052);
or U2989 (N_2989,N_425,N_349);
nand U2990 (N_2990,N_402,N_104);
xnor U2991 (N_2991,N_1043,N_313);
xor U2992 (N_2992,N_1009,N_1281);
or U2993 (N_2993,N_1479,N_764);
nand U2994 (N_2994,N_281,N_646);
nand U2995 (N_2995,N_763,N_640);
and U2996 (N_2996,N_1312,N_744);
nor U2997 (N_2997,N_1073,N_812);
and U2998 (N_2998,N_233,N_381);
nor U2999 (N_2999,N_1319,N_53);
nor U3000 (N_3000,N_2052,N_1727);
nor U3001 (N_3001,N_2720,N_1530);
or U3002 (N_3002,N_2976,N_1837);
xor U3003 (N_3003,N_2311,N_2135);
xnor U3004 (N_3004,N_2159,N_2436);
or U3005 (N_3005,N_1806,N_2300);
nand U3006 (N_3006,N_2476,N_2348);
nor U3007 (N_3007,N_2938,N_2801);
and U3008 (N_3008,N_1804,N_1868);
nand U3009 (N_3009,N_1945,N_1904);
nor U3010 (N_3010,N_2776,N_1696);
nor U3011 (N_3011,N_1703,N_1722);
and U3012 (N_3012,N_2027,N_2502);
nor U3013 (N_3013,N_2811,N_1520);
and U3014 (N_3014,N_2802,N_1562);
or U3015 (N_3015,N_1902,N_1524);
xnor U3016 (N_3016,N_2378,N_1645);
and U3017 (N_3017,N_2550,N_1617);
xor U3018 (N_3018,N_1823,N_1847);
nand U3019 (N_3019,N_2767,N_2968);
xnor U3020 (N_3020,N_2765,N_2702);
or U3021 (N_3021,N_2483,N_2501);
nand U3022 (N_3022,N_2030,N_2608);
nand U3023 (N_3023,N_2790,N_2784);
nand U3024 (N_3024,N_1824,N_2783);
xnor U3025 (N_3025,N_1856,N_2373);
or U3026 (N_3026,N_2077,N_2506);
and U3027 (N_3027,N_2635,N_2128);
nor U3028 (N_3028,N_1719,N_1517);
xor U3029 (N_3029,N_2655,N_1564);
nor U3030 (N_3030,N_1712,N_2902);
and U3031 (N_3031,N_2724,N_2481);
or U3032 (N_3032,N_1798,N_2888);
or U3033 (N_3033,N_2672,N_1637);
xnor U3034 (N_3034,N_2002,N_2020);
nor U3035 (N_3035,N_1888,N_2915);
xnor U3036 (N_3036,N_1605,N_2858);
or U3037 (N_3037,N_1646,N_2990);
nor U3038 (N_3038,N_2369,N_2735);
nor U3039 (N_3039,N_2880,N_1958);
nand U3040 (N_3040,N_2038,N_2165);
nor U3041 (N_3041,N_1840,N_2531);
nor U3042 (N_3042,N_1933,N_2952);
or U3043 (N_3043,N_2541,N_1778);
nor U3044 (N_3044,N_2658,N_2979);
nor U3045 (N_3045,N_2828,N_1923);
nand U3046 (N_3046,N_2549,N_2386);
xnor U3047 (N_3047,N_2132,N_2357);
and U3048 (N_3048,N_2682,N_2005);
and U3049 (N_3049,N_1539,N_1615);
nand U3050 (N_3050,N_2423,N_2071);
nand U3051 (N_3051,N_2210,N_1952);
or U3052 (N_3052,N_2670,N_2257);
or U3053 (N_3053,N_1619,N_2393);
nor U3054 (N_3054,N_2881,N_1765);
and U3055 (N_3055,N_2972,N_1805);
xor U3056 (N_3056,N_1582,N_1982);
or U3057 (N_3057,N_2362,N_2420);
nor U3058 (N_3058,N_2583,N_2461);
nand U3059 (N_3059,N_2248,N_2993);
xnor U3060 (N_3060,N_1946,N_2891);
nor U3061 (N_3061,N_2459,N_1748);
nor U3062 (N_3062,N_2325,N_1760);
nor U3063 (N_3063,N_1649,N_1786);
or U3064 (N_3064,N_2074,N_2309);
xor U3065 (N_3065,N_1764,N_2199);
nor U3066 (N_3066,N_2305,N_1504);
or U3067 (N_3067,N_2691,N_2176);
or U3068 (N_3068,N_2463,N_1964);
nor U3069 (N_3069,N_1828,N_2050);
and U3070 (N_3070,N_2152,N_2588);
nand U3071 (N_3071,N_1870,N_1818);
and U3072 (N_3072,N_1578,N_2901);
xnor U3073 (N_3073,N_2557,N_2838);
or U3074 (N_3074,N_2752,N_2668);
or U3075 (N_3075,N_2139,N_1745);
or U3076 (N_3076,N_1723,N_1730);
nor U3077 (N_3077,N_1788,N_2489);
or U3078 (N_3078,N_2546,N_2690);
and U3079 (N_3079,N_2145,N_2162);
nor U3080 (N_3080,N_2742,N_2841);
or U3081 (N_3081,N_2298,N_2101);
or U3082 (N_3082,N_1709,N_2948);
nor U3083 (N_3083,N_1717,N_1859);
xor U3084 (N_3084,N_2236,N_2195);
nand U3085 (N_3085,N_1598,N_2959);
xnor U3086 (N_3086,N_1893,N_2033);
nor U3087 (N_3087,N_2158,N_2708);
xnor U3088 (N_3088,N_2225,N_2409);
xor U3089 (N_3089,N_2653,N_2478);
and U3090 (N_3090,N_2065,N_2839);
and U3091 (N_3091,N_2267,N_1927);
or U3092 (N_3092,N_1607,N_2333);
nand U3093 (N_3093,N_1855,N_1987);
and U3094 (N_3094,N_2835,N_2249);
xor U3095 (N_3095,N_1542,N_1635);
nor U3096 (N_3096,N_2810,N_1708);
or U3097 (N_3097,N_2946,N_1548);
or U3098 (N_3098,N_1971,N_1928);
xnor U3099 (N_3099,N_2494,N_2751);
nand U3100 (N_3100,N_2078,N_2469);
nand U3101 (N_3101,N_2407,N_2713);
nand U3102 (N_3102,N_2542,N_2062);
nand U3103 (N_3103,N_2777,N_2485);
or U3104 (N_3104,N_2214,N_2610);
nand U3105 (N_3105,N_2491,N_2171);
or U3106 (N_3106,N_1892,N_2906);
or U3107 (N_3107,N_1606,N_2007);
nand U3108 (N_3108,N_1726,N_2253);
nor U3109 (N_3109,N_2592,N_2831);
or U3110 (N_3110,N_2336,N_2000);
or U3111 (N_3111,N_2875,N_2524);
nor U3112 (N_3112,N_2846,N_2046);
nand U3113 (N_3113,N_2163,N_2315);
or U3114 (N_3114,N_2111,N_1999);
xnor U3115 (N_3115,N_1960,N_1947);
nand U3116 (N_3116,N_2868,N_2757);
or U3117 (N_3117,N_1616,N_1560);
or U3118 (N_3118,N_2486,N_2568);
xor U3119 (N_3119,N_1643,N_2345);
xor U3120 (N_3120,N_2351,N_2642);
or U3121 (N_3121,N_1853,N_1647);
and U3122 (N_3122,N_2308,N_1629);
nand U3123 (N_3123,N_2109,N_2271);
and U3124 (N_3124,N_2723,N_2657);
xnor U3125 (N_3125,N_1826,N_2645);
nand U3126 (N_3126,N_1846,N_2866);
xnor U3127 (N_3127,N_2072,N_2701);
xnor U3128 (N_3128,N_2457,N_2586);
nor U3129 (N_3129,N_2445,N_2400);
and U3130 (N_3130,N_1660,N_2056);
nand U3131 (N_3131,N_2410,N_2837);
and U3132 (N_3132,N_2477,N_2370);
nor U3133 (N_3133,N_2185,N_2661);
nor U3134 (N_3134,N_2646,N_2431);
or U3135 (N_3135,N_1995,N_2045);
and U3136 (N_3136,N_1869,N_2180);
xor U3137 (N_3137,N_2355,N_2081);
and U3138 (N_3138,N_1527,N_2890);
nand U3139 (N_3139,N_1711,N_1608);
nor U3140 (N_3140,N_2048,N_2090);
nor U3141 (N_3141,N_2965,N_2201);
or U3142 (N_3142,N_2977,N_2051);
nand U3143 (N_3143,N_2921,N_2272);
and U3144 (N_3144,N_2747,N_1916);
and U3145 (N_3145,N_2627,N_2403);
nand U3146 (N_3146,N_1781,N_2037);
or U3147 (N_3147,N_2907,N_2816);
and U3148 (N_3148,N_1566,N_2834);
nor U3149 (N_3149,N_2986,N_2064);
or U3150 (N_3150,N_2874,N_1509);
or U3151 (N_3151,N_2454,N_2399);
or U3152 (N_3152,N_1599,N_2694);
xnor U3153 (N_3153,N_1561,N_1796);
nor U3154 (N_3154,N_2900,N_2745);
xor U3155 (N_3155,N_1570,N_2832);
and U3156 (N_3156,N_1501,N_1985);
nor U3157 (N_3157,N_2628,N_1890);
or U3158 (N_3158,N_2482,N_1515);
and U3159 (N_3159,N_2367,N_2060);
xnor U3160 (N_3160,N_2252,N_2748);
nor U3161 (N_3161,N_2458,N_2607);
and U3162 (N_3162,N_2974,N_2865);
nand U3163 (N_3163,N_2329,N_1986);
xor U3164 (N_3164,N_2093,N_2406);
xor U3165 (N_3165,N_2232,N_2994);
nand U3166 (N_3166,N_2640,N_1678);
or U3167 (N_3167,N_1857,N_2989);
xor U3168 (N_3168,N_2917,N_2619);
nor U3169 (N_3169,N_2818,N_2840);
nor U3170 (N_3170,N_2326,N_2677);
or U3171 (N_3171,N_2319,N_2995);
nand U3172 (N_3172,N_2911,N_2168);
or U3173 (N_3173,N_1767,N_1731);
nor U3174 (N_3174,N_2036,N_2375);
and U3175 (N_3175,N_2953,N_2039);
nand U3176 (N_3176,N_2435,N_2470);
xor U3177 (N_3177,N_1636,N_2753);
or U3178 (N_3178,N_2983,N_2923);
nor U3179 (N_3179,N_2722,N_1741);
and U3180 (N_3180,N_2258,N_1942);
xnor U3181 (N_3181,N_1791,N_2872);
or U3182 (N_3182,N_2604,N_1925);
nand U3183 (N_3183,N_1962,N_2277);
or U3184 (N_3184,N_1692,N_1753);
nand U3185 (N_3185,N_2746,N_1743);
or U3186 (N_3186,N_2088,N_2630);
nand U3187 (N_3187,N_2716,N_2584);
and U3188 (N_3188,N_2766,N_2026);
and U3189 (N_3189,N_2732,N_2867);
nand U3190 (N_3190,N_2164,N_1513);
nand U3191 (N_3191,N_2161,N_1655);
or U3192 (N_3192,N_2927,N_2744);
nor U3193 (N_3193,N_1961,N_2573);
nand U3194 (N_3194,N_1894,N_2131);
or U3195 (N_3195,N_2594,N_2652);
xnor U3196 (N_3196,N_2044,N_2443);
and U3197 (N_3197,N_1871,N_2103);
nand U3198 (N_3198,N_2422,N_1863);
and U3199 (N_3199,N_2439,N_2073);
nor U3200 (N_3200,N_1911,N_2061);
nor U3201 (N_3201,N_2449,N_1734);
or U3202 (N_3202,N_2089,N_2666);
or U3203 (N_3203,N_2869,N_2565);
nand U3204 (N_3204,N_2845,N_2692);
nor U3205 (N_3205,N_2391,N_1750);
and U3206 (N_3206,N_2206,N_2421);
and U3207 (N_3207,N_1864,N_2532);
nor U3208 (N_3208,N_1662,N_1682);
nand U3209 (N_3209,N_1541,N_2432);
xnor U3210 (N_3210,N_2616,N_1814);
and U3211 (N_3211,N_2467,N_1590);
nor U3212 (N_3212,N_2499,N_2197);
xor U3213 (N_3213,N_2262,N_2817);
and U3214 (N_3214,N_2942,N_2969);
xor U3215 (N_3215,N_2040,N_1833);
xor U3216 (N_3216,N_2173,N_2762);
nand U3217 (N_3217,N_1956,N_1758);
xnor U3218 (N_3218,N_2374,N_1808);
nor U3219 (N_3219,N_2970,N_2123);
or U3220 (N_3220,N_1525,N_2255);
nand U3221 (N_3221,N_2384,N_2263);
or U3222 (N_3222,N_2562,N_2782);
or U3223 (N_3223,N_1867,N_2772);
nand U3224 (N_3224,N_2122,N_2612);
or U3225 (N_3225,N_2515,N_2428);
or U3226 (N_3226,N_2426,N_2718);
xor U3227 (N_3227,N_2217,N_2053);
nor U3228 (N_3228,N_1913,N_2058);
nand U3229 (N_3229,N_1984,N_1609);
and U3230 (N_3230,N_2287,N_2887);
or U3231 (N_3231,N_2087,N_1991);
nand U3232 (N_3232,N_2773,N_2647);
xnor U3233 (N_3233,N_1702,N_2864);
nor U3234 (N_3234,N_2219,N_2849);
nand U3235 (N_3235,N_2699,N_1792);
xor U3236 (N_3236,N_1969,N_1965);
nand U3237 (N_3237,N_1751,N_2031);
xor U3238 (N_3238,N_2117,N_2352);
nand U3239 (N_3239,N_2679,N_2144);
nand U3240 (N_3240,N_1897,N_2689);
or U3241 (N_3241,N_1966,N_1924);
xor U3242 (N_3242,N_2274,N_1533);
and U3243 (N_3243,N_2803,N_2106);
nand U3244 (N_3244,N_2843,N_1754);
and U3245 (N_3245,N_2855,N_1879);
or U3246 (N_3246,N_1790,N_2259);
xor U3247 (N_3247,N_2341,N_2205);
xnor U3248 (N_3248,N_1626,N_2231);
or U3249 (N_3249,N_2737,N_1983);
nand U3250 (N_3250,N_2022,N_2987);
and U3251 (N_3251,N_1832,N_2365);
and U3252 (N_3252,N_2364,N_2908);
and U3253 (N_3253,N_2430,N_2024);
nand U3254 (N_3254,N_2581,N_2247);
nand U3255 (N_3255,N_2285,N_1794);
or U3256 (N_3256,N_2340,N_2934);
nand U3257 (N_3257,N_2954,N_2779);
nand U3258 (N_3258,N_2508,N_2631);
xnor U3259 (N_3259,N_2154,N_2929);
and U3260 (N_3260,N_2376,N_2015);
or U3261 (N_3261,N_2504,N_2394);
and U3262 (N_3262,N_2316,N_1877);
or U3263 (N_3263,N_2611,N_2202);
nor U3264 (N_3264,N_2184,N_2105);
nor U3265 (N_3265,N_2768,N_2785);
or U3266 (N_3266,N_2119,N_2805);
and U3267 (N_3267,N_2844,N_2149);
or U3268 (N_3268,N_2335,N_2726);
and U3269 (N_3269,N_1631,N_2894);
or U3270 (N_3270,N_1848,N_2648);
or U3271 (N_3271,N_2936,N_2043);
xnor U3272 (N_3272,N_2503,N_2956);
nand U3273 (N_3273,N_2032,N_2150);
or U3274 (N_3274,N_2674,N_2561);
xnor U3275 (N_3275,N_1736,N_2118);
nor U3276 (N_3276,N_2728,N_1816);
xnor U3277 (N_3277,N_2415,N_1777);
nand U3278 (N_3278,N_2480,N_2035);
or U3279 (N_3279,N_2736,N_2223);
and U3280 (N_3280,N_1595,N_2447);
nor U3281 (N_3281,N_2633,N_2448);
nor U3282 (N_3282,N_2136,N_2034);
nor U3283 (N_3283,N_2905,N_2229);
nand U3284 (N_3284,N_2730,N_2179);
xor U3285 (N_3285,N_2492,N_1632);
or U3286 (N_3286,N_2237,N_2526);
and U3287 (N_3287,N_2731,N_2893);
xnor U3288 (N_3288,N_2011,N_1621);
nand U3289 (N_3289,N_1716,N_2575);
or U3290 (N_3290,N_2517,N_2638);
nor U3291 (N_3291,N_2112,N_1644);
xnor U3292 (N_3292,N_2388,N_1679);
nand U3293 (N_3293,N_1648,N_2497);
nor U3294 (N_3294,N_2949,N_2697);
or U3295 (N_3295,N_2456,N_2127);
xnor U3296 (N_3296,N_2585,N_1953);
nor U3297 (N_3297,N_2903,N_2660);
and U3298 (N_3298,N_2787,N_1671);
or U3299 (N_3299,N_1785,N_1554);
xor U3300 (N_3300,N_1979,N_1683);
nor U3301 (N_3301,N_1576,N_2066);
nor U3302 (N_3302,N_1993,N_2462);
or U3303 (N_3303,N_2955,N_1669);
xnor U3304 (N_3304,N_2387,N_2487);
nor U3305 (N_3305,N_2589,N_2595);
and U3306 (N_3306,N_1774,N_2650);
xor U3307 (N_3307,N_2290,N_2010);
nor U3308 (N_3308,N_1591,N_1914);
or U3309 (N_3309,N_2804,N_2576);
nand U3310 (N_3310,N_1883,N_1603);
or U3311 (N_3311,N_2615,N_1843);
nand U3312 (N_3312,N_2978,N_2626);
nor U3313 (N_3313,N_2068,N_2922);
and U3314 (N_3314,N_1976,N_2649);
nand U3315 (N_3315,N_1875,N_2244);
or U3316 (N_3316,N_2299,N_1663);
xor U3317 (N_3317,N_1784,N_1728);
nor U3318 (N_3318,N_2795,N_2157);
nor U3319 (N_3319,N_2166,N_1813);
and U3320 (N_3320,N_2466,N_1587);
nor U3321 (N_3321,N_1614,N_2284);
and U3322 (N_3322,N_2143,N_2475);
xor U3323 (N_3323,N_2600,N_2055);
nor U3324 (N_3324,N_2641,N_2813);
or U3325 (N_3325,N_2383,N_2438);
xnor U3326 (N_3326,N_1651,N_2572);
nor U3327 (N_3327,N_1756,N_2663);
xnor U3328 (N_3328,N_2991,N_1811);
or U3329 (N_3329,N_2707,N_2529);
nand U3330 (N_3330,N_1620,N_2347);
xor U3331 (N_3331,N_2268,N_2304);
or U3332 (N_3332,N_1740,N_2873);
or U3333 (N_3333,N_2819,N_1691);
xor U3334 (N_3334,N_1665,N_2192);
xnor U3335 (N_3335,N_2537,N_2181);
xor U3336 (N_3336,N_2187,N_1768);
nand U3337 (N_3337,N_2919,N_2273);
nand U3338 (N_3338,N_2230,N_2774);
nor U3339 (N_3339,N_2850,N_1565);
nand U3340 (N_3340,N_2870,N_1771);
nor U3341 (N_3341,N_2239,N_1543);
nand U3342 (N_3342,N_2014,N_1831);
or U3343 (N_3343,N_2148,N_2629);
nor U3344 (N_3344,N_2009,N_2320);
nand U3345 (N_3345,N_1625,N_2433);
and U3346 (N_3346,N_2241,N_2621);
or U3347 (N_3347,N_1820,N_1989);
xor U3348 (N_3348,N_2985,N_2964);
nor U3349 (N_3349,N_2349,N_1738);
xnor U3350 (N_3350,N_2429,N_2997);
and U3351 (N_3351,N_2590,N_1687);
xor U3352 (N_3352,N_2973,N_2301);
nor U3353 (N_3353,N_1623,N_1929);
xor U3354 (N_3354,N_1567,N_2548);
xnor U3355 (N_3355,N_1807,N_2528);
nor U3356 (N_3356,N_2509,N_1749);
nand U3357 (N_3357,N_1659,N_1638);
and U3358 (N_3358,N_1546,N_2396);
nand U3359 (N_3359,N_2013,N_2861);
nand U3360 (N_3360,N_1729,N_1675);
xor U3361 (N_3361,N_2847,N_1510);
nor U3362 (N_3362,N_2084,N_2366);
nand U3363 (N_3363,N_1575,N_1656);
and U3364 (N_3364,N_1944,N_1650);
nand U3365 (N_3365,N_2593,N_2750);
and U3366 (N_3366,N_1940,N_1919);
or U3367 (N_3367,N_2306,N_1742);
xnor U3368 (N_3368,N_1770,N_2878);
nand U3369 (N_3369,N_2980,N_1994);
nor U3370 (N_3370,N_1528,N_2727);
nand U3371 (N_3371,N_2534,N_2564);
xor U3372 (N_3372,N_2076,N_2662);
or U3373 (N_3373,N_2740,N_1630);
nor U3374 (N_3374,N_2715,N_2587);
or U3375 (N_3375,N_2703,N_2233);
nor U3376 (N_3376,N_2389,N_2883);
xnor U3377 (N_3377,N_2178,N_2709);
or U3378 (N_3378,N_2981,N_1556);
nor U3379 (N_3379,N_2170,N_2042);
nor U3380 (N_3380,N_2222,N_2684);
nor U3381 (N_3381,N_1674,N_2198);
nand U3382 (N_3382,N_2472,N_2829);
nand U3383 (N_3383,N_2780,N_2656);
or U3384 (N_3384,N_1755,N_1901);
and U3385 (N_3385,N_1553,N_1512);
or U3386 (N_3386,N_2121,N_2892);
nor U3387 (N_3387,N_2967,N_2518);
nor U3388 (N_3388,N_1930,N_2473);
xnor U3389 (N_3389,N_1747,N_1628);
or U3390 (N_3390,N_2282,N_2675);
and U3391 (N_3391,N_2687,N_2857);
nor U3392 (N_3392,N_2108,N_2097);
and U3393 (N_3393,N_1865,N_1851);
xor U3394 (N_3394,N_1910,N_2380);
nand U3395 (N_3395,N_1761,N_2332);
nand U3396 (N_3396,N_2533,N_2328);
and U3397 (N_3397,N_2634,N_1954);
or U3398 (N_3398,N_2414,N_2183);
nor U3399 (N_3399,N_1695,N_2514);
nor U3400 (N_3400,N_1589,N_2558);
or U3401 (N_3401,N_2113,N_2789);
nor U3402 (N_3402,N_2465,N_2944);
or U3403 (N_3403,N_2279,N_2717);
xnor U3404 (N_3404,N_2155,N_2212);
nor U3405 (N_3405,N_1858,N_2698);
nand U3406 (N_3406,N_2297,N_2075);
xor U3407 (N_3407,N_2413,N_2931);
xor U3408 (N_3408,N_2190,N_2791);
and U3409 (N_3409,N_1921,N_2398);
nand U3410 (N_3410,N_1834,N_1523);
nand U3411 (N_3411,N_1508,N_2153);
or U3412 (N_3412,N_1992,N_1502);
xor U3413 (N_3413,N_1941,N_2729);
and U3414 (N_3414,N_1900,N_1949);
nor U3415 (N_3415,N_2004,N_2028);
and U3416 (N_3416,N_2963,N_2360);
nand U3417 (N_3417,N_1948,N_2254);
nand U3418 (N_3418,N_2063,N_2047);
or U3419 (N_3419,N_1693,N_2137);
and U3420 (N_3420,N_1839,N_2574);
nor U3421 (N_3421,N_1592,N_1641);
nand U3422 (N_3422,N_2226,N_2317);
or U3423 (N_3423,N_2437,N_2852);
or U3424 (N_3424,N_1822,N_1699);
nand U3425 (N_3425,N_2871,N_2371);
xnor U3426 (N_3426,N_2884,N_2704);
nor U3427 (N_3427,N_2734,N_2275);
or U3428 (N_3428,N_2823,N_2826);
nand U3429 (N_3429,N_1787,N_2256);
nor U3430 (N_3430,N_2292,N_2937);
and U3431 (N_3431,N_1852,N_2250);
and U3432 (N_3432,N_2833,N_2895);
or U3433 (N_3433,N_2142,N_2602);
and U3434 (N_3434,N_2909,N_2115);
and U3435 (N_3435,N_2029,N_2951);
or U3436 (N_3436,N_1835,N_2368);
nor U3437 (N_3437,N_1588,N_1872);
nor U3438 (N_3438,N_1559,N_2182);
xnor U3439 (N_3439,N_1684,N_2654);
nor U3440 (N_3440,N_2941,N_1988);
nor U3441 (N_3441,N_2344,N_2207);
nor U3442 (N_3442,N_2786,N_1757);
nor U3443 (N_3443,N_2688,N_2186);
xnor U3444 (N_3444,N_2283,N_1574);
or U3445 (N_3445,N_1762,N_1676);
xor U3446 (N_3446,N_1874,N_2536);
and U3447 (N_3447,N_1547,N_1664);
and U3448 (N_3448,N_2450,N_2008);
xnor U3449 (N_3449,N_2114,N_1780);
nor U3450 (N_3450,N_2769,N_2792);
nor U3451 (N_3451,N_1766,N_2552);
or U3452 (N_3452,N_2651,N_1885);
or U3453 (N_3453,N_2664,N_2996);
nor U3454 (N_3454,N_1604,N_2982);
nor U3455 (N_3455,N_1521,N_2778);
nand U3456 (N_3456,N_1795,N_2382);
nand U3457 (N_3457,N_2234,N_2617);
nor U3458 (N_3458,N_2401,N_2966);
or U3459 (N_3459,N_2270,N_1600);
nand U3460 (N_3460,N_2577,N_2825);
xor U3461 (N_3461,N_2681,N_2411);
xor U3462 (N_3462,N_2912,N_1680);
xor U3463 (N_3463,N_1772,N_1585);
nand U3464 (N_3464,N_1531,N_2719);
nor U3465 (N_3465,N_2337,N_1866);
nor U3466 (N_3466,N_2194,N_1549);
and U3467 (N_3467,N_2019,N_1861);
nand U3468 (N_3468,N_2538,N_2754);
nand U3469 (N_3469,N_2644,N_1596);
xnor U3470 (N_3470,N_1555,N_2307);
nor U3471 (N_3471,N_1661,N_1815);
or U3472 (N_3472,N_2579,N_1918);
or U3473 (N_3473,N_1640,N_2067);
and U3474 (N_3474,N_1704,N_2224);
nor U3475 (N_3475,N_1746,N_1972);
nand U3476 (N_3476,N_1819,N_2356);
xor U3477 (N_3477,N_2624,N_1580);
nand U3478 (N_3478,N_2312,N_2877);
nor U3479 (N_3479,N_2842,N_2759);
xnor U3480 (N_3480,N_2797,N_1903);
and U3481 (N_3481,N_1597,N_1882);
or U3482 (N_3482,N_2025,N_1579);
nor U3483 (N_3483,N_2623,N_2943);
xnor U3484 (N_3484,N_2221,N_2334);
and U3485 (N_3485,N_2721,N_1797);
nand U3486 (N_3486,N_2147,N_2243);
nor U3487 (N_3487,N_1516,N_1799);
nor U3488 (N_3488,N_2808,N_2156);
nor U3489 (N_3489,N_2208,N_2683);
nor U3490 (N_3490,N_2488,N_2601);
or U3491 (N_3491,N_2310,N_2510);
nor U3492 (N_3492,N_2196,N_1666);
or U3493 (N_3493,N_1688,N_1936);
xor U3494 (N_3494,N_2296,N_2434);
or U3495 (N_3495,N_2669,N_2338);
and U3496 (N_3496,N_2827,N_2330);
and U3497 (N_3497,N_1563,N_2417);
and U3498 (N_3498,N_1889,N_2507);
xor U3499 (N_3499,N_2738,N_2960);
nor U3500 (N_3500,N_2100,N_2559);
and U3501 (N_3501,N_2676,N_2814);
xor U3502 (N_3502,N_1633,N_1594);
and U3503 (N_3503,N_2442,N_2853);
nand U3504 (N_3504,N_1895,N_2527);
xnor U3505 (N_3505,N_2696,N_2342);
or U3506 (N_3506,N_1724,N_2695);
xor U3507 (N_3507,N_2775,N_2924);
or U3508 (N_3508,N_2516,N_1763);
xnor U3509 (N_3509,N_2464,N_2609);
xnor U3510 (N_3510,N_2291,N_1963);
or U3511 (N_3511,N_2522,N_1612);
xor U3512 (N_3512,N_1618,N_1891);
xor U3513 (N_3513,N_1844,N_2597);
and U3514 (N_3514,N_2092,N_2193);
xnor U3515 (N_3515,N_1909,N_2714);
nand U3516 (N_3516,N_1970,N_2018);
xor U3517 (N_3517,N_2798,N_2896);
nand U3518 (N_3518,N_2395,N_1627);
nand U3519 (N_3519,N_2511,N_2054);
xor U3520 (N_3520,N_2331,N_2686);
nor U3521 (N_3521,N_2918,N_2794);
nand U3522 (N_3522,N_2961,N_2935);
nand U3523 (N_3523,N_1568,N_2266);
nor U3524 (N_3524,N_2578,N_1668);
xnor U3525 (N_3525,N_1686,N_1583);
or U3526 (N_3526,N_2620,N_1978);
nand U3527 (N_3527,N_2830,N_1540);
nand U3528 (N_3528,N_1672,N_2260);
nand U3529 (N_3529,N_2760,N_1873);
nand U3530 (N_3530,N_2678,N_2016);
nor U3531 (N_3531,N_2130,N_2567);
or U3532 (N_3532,N_2639,N_1845);
nand U3533 (N_3533,N_2749,N_1737);
and U3534 (N_3534,N_2474,N_1690);
and U3535 (N_3535,N_1534,N_2566);
nand U3536 (N_3536,N_1912,N_2859);
xnor U3537 (N_3537,N_2441,N_2812);
or U3538 (N_3538,N_1526,N_2886);
or U3539 (N_3539,N_2671,N_2898);
nor U3540 (N_3540,N_2003,N_1908);
nor U3541 (N_3541,N_2339,N_1550);
or U3542 (N_3542,N_2926,N_1642);
nand U3543 (N_3543,N_2096,N_1522);
nand U3544 (N_3544,N_1810,N_1573);
or U3545 (N_3545,N_1571,N_1507);
nand U3546 (N_3546,N_2126,N_1829);
and U3547 (N_3547,N_2560,N_2800);
nor U3548 (N_3548,N_1500,N_2021);
or U3549 (N_3549,N_2110,N_2006);
or U3550 (N_3550,N_2544,N_2806);
or U3551 (N_3551,N_2167,N_2390);
nor U3552 (N_3552,N_1943,N_2091);
nand U3553 (N_3553,N_1981,N_1937);
xnor U3554 (N_3554,N_2519,N_2302);
xor U3555 (N_3555,N_1634,N_1658);
and U3556 (N_3556,N_1569,N_2796);
and U3557 (N_3557,N_1572,N_1593);
or U3558 (N_3558,N_2361,N_1652);
nor U3559 (N_3559,N_1884,N_2525);
xnor U3560 (N_3560,N_2083,N_2856);
or U3561 (N_3561,N_2405,N_1939);
or U3562 (N_3562,N_2318,N_2932);
and U3563 (N_3563,N_2693,N_2294);
xnor U3564 (N_3564,N_2613,N_2363);
nand U3565 (N_3565,N_2385,N_1698);
or U3566 (N_3566,N_1782,N_1535);
xnor U3567 (N_3567,N_2209,N_2490);
nor U3568 (N_3568,N_2240,N_2359);
xnor U3569 (N_3569,N_2799,N_1906);
xor U3570 (N_3570,N_1779,N_2582);
nor U3571 (N_3571,N_1701,N_2712);
or U3572 (N_3572,N_2771,N_2764);
or U3573 (N_3573,N_2739,N_2521);
or U3574 (N_3574,N_1959,N_2512);
nand U3575 (N_3575,N_2440,N_2321);
xor U3576 (N_3576,N_1803,N_2451);
nor U3577 (N_3577,N_2276,N_2700);
xor U3578 (N_3578,N_2637,N_2295);
xnor U3579 (N_3579,N_2041,N_2346);
nand U3580 (N_3580,N_2603,N_2314);
nand U3581 (N_3581,N_2453,N_1557);
xor U3582 (N_3582,N_2822,N_2599);
nand U3583 (N_3583,N_2904,N_1821);
nor U3584 (N_3584,N_2377,N_2910);
xor U3585 (N_3585,N_2605,N_1714);
nor U3586 (N_3586,N_2945,N_1881);
or U3587 (N_3587,N_2913,N_2992);
and U3588 (N_3588,N_2513,N_2471);
nor U3589 (N_3589,N_1558,N_1720);
nor U3590 (N_3590,N_2824,N_1586);
or U3591 (N_3591,N_1990,N_1536);
nor U3592 (N_3592,N_2099,N_2444);
or U3593 (N_3593,N_1759,N_1705);
nand U3594 (N_3594,N_2151,N_2104);
nor U3595 (N_3595,N_1935,N_2755);
nand U3596 (N_3596,N_2281,N_2547);
xnor U3597 (N_3597,N_1769,N_1957);
nand U3598 (N_3598,N_1685,N_2882);
xor U3599 (N_3599,N_2733,N_2288);
nor U3600 (N_3600,N_2012,N_1801);
nor U3601 (N_3601,N_2228,N_1951);
xnor U3602 (N_3602,N_1545,N_1673);
nor U3603 (N_3603,N_1610,N_2925);
and U3604 (N_3604,N_2069,N_1725);
nand U3605 (N_3605,N_2085,N_2758);
nand U3606 (N_3606,N_2098,N_1973);
xnor U3607 (N_3607,N_1950,N_2323);
or U3608 (N_3608,N_2998,N_2238);
nor U3609 (N_3609,N_1505,N_2261);
or U3610 (N_3610,N_2618,N_2402);
xor U3611 (N_3611,N_1529,N_1689);
nor U3612 (N_3612,N_2914,N_2821);
xnor U3613 (N_3613,N_1532,N_2191);
or U3614 (N_3614,N_1955,N_2289);
nand U3615 (N_3615,N_1776,N_1789);
and U3616 (N_3616,N_2452,N_2962);
nor U3617 (N_3617,N_2353,N_2418);
nor U3618 (N_3618,N_2269,N_2070);
nand U3619 (N_3619,N_2140,N_1713);
nand U3620 (N_3620,N_1817,N_1657);
and U3621 (N_3621,N_2815,N_2141);
and U3622 (N_3622,N_2569,N_2424);
nand U3623 (N_3623,N_2479,N_1602);
nor U3624 (N_3624,N_2553,N_1653);
nor U3625 (N_3625,N_2235,N_2889);
nand U3626 (N_3626,N_2807,N_1880);
nor U3627 (N_3627,N_1639,N_2876);
and U3628 (N_3628,N_2079,N_2498);
or U3629 (N_3629,N_1739,N_2227);
and U3630 (N_3630,N_2950,N_2788);
xor U3631 (N_3631,N_2189,N_2591);
and U3632 (N_3632,N_2200,N_2947);
or U3633 (N_3633,N_1967,N_2120);
nor U3634 (N_3634,N_1654,N_2350);
nand U3635 (N_3635,N_2220,N_2975);
xnor U3636 (N_3636,N_1998,N_2493);
nor U3637 (N_3637,N_1744,N_2933);
nor U3638 (N_3638,N_2408,N_2523);
xnor U3639 (N_3639,N_2636,N_2863);
nand U3640 (N_3640,N_2756,N_2211);
nor U3641 (N_3641,N_1932,N_2862);
or U3642 (N_3642,N_2322,N_2885);
nand U3643 (N_3643,N_2133,N_2930);
xnor U3644 (N_3644,N_1551,N_1700);
nor U3645 (N_3645,N_1718,N_1899);
nand U3646 (N_3646,N_2530,N_2836);
xor U3647 (N_3647,N_1670,N_2286);
or U3648 (N_3648,N_2124,N_2425);
or U3649 (N_3649,N_2851,N_2082);
and U3650 (N_3650,N_1775,N_1887);
or U3651 (N_3651,N_2354,N_2665);
xnor U3652 (N_3652,N_2412,N_2685);
and U3653 (N_3653,N_2484,N_2107);
nand U3654 (N_3654,N_1537,N_2134);
or U3655 (N_3655,N_1862,N_2245);
nand U3656 (N_3656,N_1710,N_1854);
nor U3657 (N_3657,N_2632,N_2392);
nor U3658 (N_3658,N_2023,N_2957);
xor U3659 (N_3659,N_2057,N_1922);
nand U3660 (N_3660,N_1926,N_2673);
nor U3661 (N_3661,N_1827,N_2899);
and U3662 (N_3662,N_2781,N_1907);
nand U3663 (N_3663,N_1842,N_2264);
and U3664 (N_3664,N_2659,N_2265);
nand U3665 (N_3665,N_1735,N_2455);
and U3666 (N_3666,N_2280,N_2102);
nor U3667 (N_3667,N_2358,N_1707);
nor U3668 (N_3668,N_2086,N_2419);
and U3669 (N_3669,N_2049,N_1624);
or U3670 (N_3670,N_1850,N_2203);
or U3671 (N_3671,N_1996,N_2213);
nand U3672 (N_3672,N_2059,N_1800);
nand U3673 (N_3673,N_2381,N_2460);
nand U3674 (N_3674,N_1538,N_2770);
nor U3675 (N_3675,N_2860,N_2500);
nor U3676 (N_3676,N_2563,N_1802);
and U3677 (N_3677,N_2251,N_2324);
nor U3678 (N_3678,N_2556,N_2711);
and U3679 (N_3679,N_2246,N_1622);
or U3680 (N_3680,N_1876,N_2741);
or U3681 (N_3681,N_2129,N_2706);
nand U3682 (N_3682,N_2879,N_2095);
xnor U3683 (N_3683,N_2545,N_2303);
nand U3684 (N_3684,N_2172,N_1733);
or U3685 (N_3685,N_2372,N_1825);
nand U3686 (N_3686,N_2188,N_1849);
nand U3687 (N_3687,N_2146,N_2763);
xor U3688 (N_3688,N_2218,N_1732);
or U3689 (N_3689,N_2598,N_2174);
nand U3690 (N_3690,N_1934,N_1506);
nand U3691 (N_3691,N_1878,N_2278);
and U3692 (N_3692,N_2705,N_2999);
xnor U3693 (N_3693,N_1841,N_2643);
nor U3694 (N_3694,N_2554,N_2916);
nand U3695 (N_3695,N_2177,N_2327);
nand U3696 (N_3696,N_2551,N_2571);
nor U3697 (N_3697,N_2495,N_2138);
or U3698 (N_3698,N_1681,N_2001);
xnor U3699 (N_3699,N_2468,N_2984);
xnor U3700 (N_3700,N_1896,N_1809);
nand U3701 (N_3701,N_1584,N_2540);
or U3702 (N_3702,N_2928,N_1898);
nor U3703 (N_3703,N_1715,N_2570);
xnor U3704 (N_3704,N_2496,N_2204);
or U3705 (N_3705,N_1601,N_2293);
nor U3706 (N_3706,N_2427,N_2543);
xnor U3707 (N_3707,N_2809,N_1721);
nand U3708 (N_3708,N_1694,N_2580);
nand U3709 (N_3709,N_2397,N_2242);
and U3710 (N_3710,N_2505,N_1886);
and U3711 (N_3711,N_2080,N_1838);
or U3712 (N_3712,N_2940,N_2175);
and U3713 (N_3713,N_1974,N_1552);
xor U3714 (N_3714,N_2725,N_2555);
or U3715 (N_3715,N_2622,N_2988);
nor U3716 (N_3716,N_2614,N_1830);
and U3717 (N_3717,N_1544,N_1667);
nor U3718 (N_3718,N_2897,N_1773);
or U3719 (N_3719,N_1519,N_1917);
and U3720 (N_3720,N_1860,N_2313);
and U3721 (N_3721,N_2379,N_1518);
nand U3722 (N_3722,N_2920,N_2520);
and U3723 (N_3723,N_2539,N_1752);
or U3724 (N_3724,N_1503,N_1931);
or U3725 (N_3725,N_2169,N_2094);
and U3726 (N_3726,N_2958,N_2820);
xnor U3727 (N_3727,N_1980,N_1812);
nand U3728 (N_3728,N_1706,N_2761);
nor U3729 (N_3729,N_1975,N_2596);
and U3730 (N_3730,N_2216,N_2606);
nor U3731 (N_3731,N_1997,N_1905);
nor U3732 (N_3732,N_2017,N_1577);
and U3733 (N_3733,N_2667,N_2404);
and U3734 (N_3734,N_2939,N_2215);
xnor U3735 (N_3735,N_1611,N_1783);
or U3736 (N_3736,N_2848,N_1938);
or U3737 (N_3737,N_2535,N_2854);
or U3738 (N_3738,N_2793,N_1793);
or U3739 (N_3739,N_1677,N_1915);
and U3740 (N_3740,N_2416,N_2446);
xnor U3741 (N_3741,N_1836,N_2971);
nor U3742 (N_3742,N_2116,N_1697);
or U3743 (N_3743,N_1968,N_2680);
nor U3744 (N_3744,N_2710,N_1613);
nand U3745 (N_3745,N_1977,N_2343);
xor U3746 (N_3746,N_2743,N_2125);
or U3747 (N_3747,N_2160,N_1514);
xor U3748 (N_3748,N_2625,N_1511);
and U3749 (N_3749,N_1920,N_1581);
nand U3750 (N_3750,N_1737,N_2710);
nor U3751 (N_3751,N_2975,N_1677);
and U3752 (N_3752,N_2106,N_1581);
and U3753 (N_3753,N_1794,N_2094);
nand U3754 (N_3754,N_2544,N_2866);
nor U3755 (N_3755,N_2200,N_1683);
nand U3756 (N_3756,N_2442,N_2622);
nor U3757 (N_3757,N_2803,N_1645);
or U3758 (N_3758,N_2905,N_2767);
xnor U3759 (N_3759,N_2631,N_2504);
xnor U3760 (N_3760,N_2279,N_2683);
nor U3761 (N_3761,N_1693,N_2475);
and U3762 (N_3762,N_2306,N_1988);
nand U3763 (N_3763,N_1893,N_2687);
or U3764 (N_3764,N_2391,N_1706);
nor U3765 (N_3765,N_2220,N_2287);
and U3766 (N_3766,N_1865,N_1621);
nand U3767 (N_3767,N_1742,N_1837);
xnor U3768 (N_3768,N_2051,N_1906);
and U3769 (N_3769,N_2245,N_2603);
nand U3770 (N_3770,N_2784,N_2533);
xor U3771 (N_3771,N_2055,N_2842);
and U3772 (N_3772,N_1735,N_2857);
nor U3773 (N_3773,N_2714,N_2481);
and U3774 (N_3774,N_2616,N_1712);
nand U3775 (N_3775,N_2648,N_2687);
and U3776 (N_3776,N_2326,N_2299);
xnor U3777 (N_3777,N_1555,N_1698);
or U3778 (N_3778,N_1920,N_2884);
and U3779 (N_3779,N_1825,N_2709);
or U3780 (N_3780,N_2404,N_2795);
nor U3781 (N_3781,N_2155,N_1779);
or U3782 (N_3782,N_1763,N_2409);
xor U3783 (N_3783,N_1574,N_1765);
xnor U3784 (N_3784,N_2035,N_2531);
nor U3785 (N_3785,N_1724,N_2253);
and U3786 (N_3786,N_2756,N_2469);
and U3787 (N_3787,N_1860,N_1719);
nor U3788 (N_3788,N_2301,N_2501);
xnor U3789 (N_3789,N_2884,N_2516);
and U3790 (N_3790,N_1772,N_2035);
and U3791 (N_3791,N_2825,N_2151);
and U3792 (N_3792,N_2319,N_2370);
nand U3793 (N_3793,N_2765,N_2914);
nand U3794 (N_3794,N_2376,N_2750);
or U3795 (N_3795,N_1686,N_1923);
nand U3796 (N_3796,N_2451,N_1903);
nor U3797 (N_3797,N_1664,N_2206);
nor U3798 (N_3798,N_2104,N_2635);
or U3799 (N_3799,N_2466,N_1648);
or U3800 (N_3800,N_2184,N_1969);
xnor U3801 (N_3801,N_1882,N_2557);
or U3802 (N_3802,N_1871,N_1951);
nor U3803 (N_3803,N_1706,N_2976);
and U3804 (N_3804,N_1877,N_2290);
nor U3805 (N_3805,N_2620,N_1661);
and U3806 (N_3806,N_2773,N_2542);
and U3807 (N_3807,N_2384,N_1867);
or U3808 (N_3808,N_2891,N_2576);
nand U3809 (N_3809,N_2660,N_2208);
nor U3810 (N_3810,N_2227,N_2589);
or U3811 (N_3811,N_2107,N_1680);
and U3812 (N_3812,N_2900,N_1697);
xnor U3813 (N_3813,N_1889,N_2293);
xnor U3814 (N_3814,N_2800,N_1836);
or U3815 (N_3815,N_1875,N_1826);
or U3816 (N_3816,N_1536,N_2370);
nor U3817 (N_3817,N_2980,N_2355);
xor U3818 (N_3818,N_2632,N_1898);
nor U3819 (N_3819,N_1747,N_2033);
and U3820 (N_3820,N_1629,N_1594);
nor U3821 (N_3821,N_2233,N_2812);
nand U3822 (N_3822,N_2197,N_1956);
nor U3823 (N_3823,N_2133,N_1513);
nand U3824 (N_3824,N_2144,N_2050);
xnor U3825 (N_3825,N_1886,N_2058);
nand U3826 (N_3826,N_2534,N_2465);
xor U3827 (N_3827,N_2334,N_2176);
and U3828 (N_3828,N_2790,N_2803);
and U3829 (N_3829,N_1866,N_1633);
nor U3830 (N_3830,N_1741,N_1864);
or U3831 (N_3831,N_1688,N_1942);
xnor U3832 (N_3832,N_2635,N_2667);
nand U3833 (N_3833,N_2959,N_2642);
nand U3834 (N_3834,N_2995,N_2166);
nand U3835 (N_3835,N_1770,N_1968);
nor U3836 (N_3836,N_2208,N_2742);
nand U3837 (N_3837,N_2022,N_2314);
and U3838 (N_3838,N_1548,N_2411);
nand U3839 (N_3839,N_2802,N_2128);
or U3840 (N_3840,N_2254,N_2287);
and U3841 (N_3841,N_2993,N_1822);
or U3842 (N_3842,N_2018,N_1862);
xor U3843 (N_3843,N_1764,N_1931);
xor U3844 (N_3844,N_1778,N_1576);
xnor U3845 (N_3845,N_2828,N_2527);
or U3846 (N_3846,N_1609,N_2162);
nand U3847 (N_3847,N_2690,N_2550);
xor U3848 (N_3848,N_2092,N_1703);
nand U3849 (N_3849,N_2646,N_2047);
or U3850 (N_3850,N_1692,N_1561);
and U3851 (N_3851,N_1954,N_2200);
xnor U3852 (N_3852,N_2428,N_2330);
nand U3853 (N_3853,N_1863,N_2070);
and U3854 (N_3854,N_2792,N_1775);
and U3855 (N_3855,N_2878,N_2181);
and U3856 (N_3856,N_1989,N_2341);
or U3857 (N_3857,N_2023,N_2616);
and U3858 (N_3858,N_2463,N_2089);
and U3859 (N_3859,N_2776,N_2016);
nor U3860 (N_3860,N_2843,N_2082);
xor U3861 (N_3861,N_2626,N_2888);
nor U3862 (N_3862,N_2397,N_1980);
nand U3863 (N_3863,N_2781,N_1564);
and U3864 (N_3864,N_2581,N_1938);
and U3865 (N_3865,N_2187,N_1926);
nor U3866 (N_3866,N_2857,N_2222);
or U3867 (N_3867,N_2760,N_2068);
xnor U3868 (N_3868,N_2230,N_2641);
nand U3869 (N_3869,N_2363,N_2964);
and U3870 (N_3870,N_2345,N_1513);
nand U3871 (N_3871,N_2744,N_1887);
xor U3872 (N_3872,N_2061,N_2392);
xor U3873 (N_3873,N_1828,N_1772);
nand U3874 (N_3874,N_2049,N_2721);
nor U3875 (N_3875,N_1716,N_2545);
and U3876 (N_3876,N_2192,N_2694);
or U3877 (N_3877,N_2485,N_1515);
xor U3878 (N_3878,N_2526,N_2206);
nor U3879 (N_3879,N_2094,N_2250);
and U3880 (N_3880,N_2657,N_2446);
and U3881 (N_3881,N_2601,N_2231);
and U3882 (N_3882,N_2954,N_1524);
and U3883 (N_3883,N_2890,N_1771);
and U3884 (N_3884,N_1903,N_2270);
nand U3885 (N_3885,N_1966,N_2278);
and U3886 (N_3886,N_2742,N_1692);
nand U3887 (N_3887,N_2780,N_2749);
xnor U3888 (N_3888,N_1918,N_2436);
nor U3889 (N_3889,N_2636,N_2026);
xor U3890 (N_3890,N_1629,N_2192);
or U3891 (N_3891,N_2471,N_2927);
and U3892 (N_3892,N_2313,N_2269);
nor U3893 (N_3893,N_1584,N_2666);
and U3894 (N_3894,N_1940,N_2735);
nor U3895 (N_3895,N_2484,N_2494);
xnor U3896 (N_3896,N_2370,N_1770);
nor U3897 (N_3897,N_2740,N_1542);
nand U3898 (N_3898,N_2692,N_2243);
or U3899 (N_3899,N_2912,N_1514);
nor U3900 (N_3900,N_2810,N_1713);
nand U3901 (N_3901,N_1565,N_1945);
nor U3902 (N_3902,N_1669,N_1594);
nor U3903 (N_3903,N_1805,N_2594);
nand U3904 (N_3904,N_2381,N_1983);
or U3905 (N_3905,N_1721,N_2496);
or U3906 (N_3906,N_2543,N_1671);
xor U3907 (N_3907,N_1619,N_1528);
nand U3908 (N_3908,N_2270,N_2020);
or U3909 (N_3909,N_2982,N_2350);
or U3910 (N_3910,N_2781,N_1824);
and U3911 (N_3911,N_2391,N_2291);
nor U3912 (N_3912,N_2316,N_2080);
nor U3913 (N_3913,N_2885,N_2128);
xor U3914 (N_3914,N_2109,N_1875);
nand U3915 (N_3915,N_1597,N_1791);
nor U3916 (N_3916,N_2983,N_1824);
nor U3917 (N_3917,N_1678,N_2315);
nor U3918 (N_3918,N_1793,N_2645);
and U3919 (N_3919,N_1883,N_1637);
or U3920 (N_3920,N_2928,N_1990);
nor U3921 (N_3921,N_2867,N_2395);
nand U3922 (N_3922,N_2121,N_1545);
nor U3923 (N_3923,N_2275,N_2427);
or U3924 (N_3924,N_2408,N_2944);
or U3925 (N_3925,N_2511,N_1881);
or U3926 (N_3926,N_2800,N_2378);
and U3927 (N_3927,N_1978,N_2692);
nor U3928 (N_3928,N_2545,N_2423);
nand U3929 (N_3929,N_1997,N_1914);
or U3930 (N_3930,N_2877,N_2345);
nor U3931 (N_3931,N_1916,N_1668);
or U3932 (N_3932,N_1632,N_2530);
or U3933 (N_3933,N_2588,N_1947);
and U3934 (N_3934,N_2765,N_2109);
and U3935 (N_3935,N_1987,N_1727);
nand U3936 (N_3936,N_1566,N_2397);
or U3937 (N_3937,N_2169,N_2190);
nor U3938 (N_3938,N_1594,N_1969);
nand U3939 (N_3939,N_1916,N_1562);
or U3940 (N_3940,N_2283,N_2586);
and U3941 (N_3941,N_2765,N_2251);
and U3942 (N_3942,N_1610,N_2010);
nand U3943 (N_3943,N_2799,N_2472);
and U3944 (N_3944,N_1598,N_1754);
or U3945 (N_3945,N_1679,N_2666);
and U3946 (N_3946,N_2840,N_1826);
or U3947 (N_3947,N_2240,N_1850);
xnor U3948 (N_3948,N_2809,N_1515);
and U3949 (N_3949,N_2589,N_2759);
nand U3950 (N_3950,N_1546,N_2562);
nand U3951 (N_3951,N_1964,N_2695);
nand U3952 (N_3952,N_1832,N_1898);
nand U3953 (N_3953,N_1765,N_2972);
nand U3954 (N_3954,N_2293,N_2388);
and U3955 (N_3955,N_2070,N_2014);
nor U3956 (N_3956,N_2503,N_1928);
xor U3957 (N_3957,N_2480,N_2302);
nor U3958 (N_3958,N_2777,N_2144);
nand U3959 (N_3959,N_2333,N_2587);
nand U3960 (N_3960,N_2585,N_2666);
nand U3961 (N_3961,N_2778,N_2884);
xor U3962 (N_3962,N_2393,N_2640);
nand U3963 (N_3963,N_2804,N_2262);
nor U3964 (N_3964,N_1634,N_2602);
xor U3965 (N_3965,N_1741,N_2352);
nand U3966 (N_3966,N_2329,N_1649);
or U3967 (N_3967,N_1518,N_2947);
or U3968 (N_3968,N_1706,N_2196);
or U3969 (N_3969,N_2929,N_2206);
and U3970 (N_3970,N_2544,N_2205);
xor U3971 (N_3971,N_2816,N_2323);
nor U3972 (N_3972,N_1527,N_2077);
and U3973 (N_3973,N_2500,N_2026);
xnor U3974 (N_3974,N_2113,N_2774);
or U3975 (N_3975,N_2561,N_2249);
nand U3976 (N_3976,N_2628,N_2044);
nor U3977 (N_3977,N_1644,N_2128);
nand U3978 (N_3978,N_2850,N_2225);
and U3979 (N_3979,N_2184,N_1671);
xnor U3980 (N_3980,N_2204,N_2061);
nand U3981 (N_3981,N_2810,N_2433);
or U3982 (N_3982,N_2637,N_2799);
nand U3983 (N_3983,N_1830,N_2174);
nand U3984 (N_3984,N_2463,N_2261);
nor U3985 (N_3985,N_1889,N_2578);
or U3986 (N_3986,N_1811,N_2638);
and U3987 (N_3987,N_1734,N_2128);
xnor U3988 (N_3988,N_1742,N_1675);
or U3989 (N_3989,N_2185,N_2110);
and U3990 (N_3990,N_2061,N_2440);
nor U3991 (N_3991,N_2806,N_2659);
nand U3992 (N_3992,N_2052,N_1644);
and U3993 (N_3993,N_2435,N_1911);
nand U3994 (N_3994,N_1774,N_1749);
nor U3995 (N_3995,N_2202,N_1718);
xnor U3996 (N_3996,N_2018,N_2955);
nor U3997 (N_3997,N_1751,N_2660);
and U3998 (N_3998,N_2698,N_1951);
xor U3999 (N_3999,N_2191,N_2823);
nor U4000 (N_4000,N_2537,N_2917);
nor U4001 (N_4001,N_2946,N_2313);
or U4002 (N_4002,N_1976,N_2860);
and U4003 (N_4003,N_2445,N_2370);
xnor U4004 (N_4004,N_1558,N_2849);
or U4005 (N_4005,N_2066,N_2977);
nand U4006 (N_4006,N_2277,N_2666);
xnor U4007 (N_4007,N_2368,N_1931);
and U4008 (N_4008,N_1868,N_1512);
nor U4009 (N_4009,N_1507,N_2392);
xnor U4010 (N_4010,N_1959,N_2934);
nand U4011 (N_4011,N_2956,N_1614);
nor U4012 (N_4012,N_2910,N_1794);
nor U4013 (N_4013,N_2584,N_2916);
and U4014 (N_4014,N_1607,N_1699);
nor U4015 (N_4015,N_2064,N_2601);
or U4016 (N_4016,N_2257,N_2875);
nand U4017 (N_4017,N_2255,N_1679);
or U4018 (N_4018,N_2664,N_2929);
nor U4019 (N_4019,N_2669,N_2913);
and U4020 (N_4020,N_2558,N_2109);
nand U4021 (N_4021,N_2695,N_1910);
nand U4022 (N_4022,N_2828,N_2166);
xor U4023 (N_4023,N_2597,N_2948);
and U4024 (N_4024,N_1802,N_2339);
xnor U4025 (N_4025,N_1877,N_2889);
nand U4026 (N_4026,N_2495,N_2156);
nand U4027 (N_4027,N_1927,N_2482);
and U4028 (N_4028,N_2376,N_1611);
or U4029 (N_4029,N_2990,N_1513);
and U4030 (N_4030,N_2097,N_2793);
nand U4031 (N_4031,N_2379,N_2174);
or U4032 (N_4032,N_1851,N_2739);
nand U4033 (N_4033,N_1710,N_1716);
nand U4034 (N_4034,N_2393,N_2634);
and U4035 (N_4035,N_2443,N_2123);
xnor U4036 (N_4036,N_2961,N_2868);
and U4037 (N_4037,N_2036,N_2759);
xnor U4038 (N_4038,N_2153,N_1915);
and U4039 (N_4039,N_2481,N_1820);
and U4040 (N_4040,N_2301,N_2003);
and U4041 (N_4041,N_2084,N_1963);
xor U4042 (N_4042,N_1755,N_2108);
and U4043 (N_4043,N_1752,N_2285);
xnor U4044 (N_4044,N_1864,N_1711);
or U4045 (N_4045,N_2125,N_2080);
nand U4046 (N_4046,N_2099,N_2146);
or U4047 (N_4047,N_2248,N_2332);
or U4048 (N_4048,N_2986,N_2543);
nand U4049 (N_4049,N_2840,N_1718);
nor U4050 (N_4050,N_2787,N_2917);
nor U4051 (N_4051,N_2196,N_2054);
nor U4052 (N_4052,N_1941,N_2222);
nor U4053 (N_4053,N_2388,N_2358);
or U4054 (N_4054,N_2693,N_1894);
xor U4055 (N_4055,N_2312,N_2456);
nor U4056 (N_4056,N_2543,N_2237);
nor U4057 (N_4057,N_2223,N_2329);
nor U4058 (N_4058,N_1747,N_1833);
nor U4059 (N_4059,N_2857,N_1654);
and U4060 (N_4060,N_1937,N_1875);
nor U4061 (N_4061,N_2069,N_2220);
nor U4062 (N_4062,N_2214,N_2425);
nand U4063 (N_4063,N_2694,N_2505);
and U4064 (N_4064,N_1888,N_2549);
xnor U4065 (N_4065,N_2891,N_1667);
nand U4066 (N_4066,N_1588,N_2800);
nand U4067 (N_4067,N_2923,N_2890);
nand U4068 (N_4068,N_2531,N_1508);
and U4069 (N_4069,N_2262,N_2317);
xnor U4070 (N_4070,N_1640,N_2252);
or U4071 (N_4071,N_2942,N_2505);
nor U4072 (N_4072,N_1734,N_1874);
nand U4073 (N_4073,N_1955,N_2769);
nand U4074 (N_4074,N_1978,N_2393);
xor U4075 (N_4075,N_1586,N_1984);
and U4076 (N_4076,N_2881,N_2470);
or U4077 (N_4077,N_1903,N_2440);
and U4078 (N_4078,N_1599,N_2961);
nor U4079 (N_4079,N_1979,N_1587);
nand U4080 (N_4080,N_2231,N_2095);
nor U4081 (N_4081,N_2753,N_2632);
or U4082 (N_4082,N_2849,N_2962);
or U4083 (N_4083,N_2718,N_2704);
or U4084 (N_4084,N_1824,N_2904);
xnor U4085 (N_4085,N_2610,N_1720);
and U4086 (N_4086,N_2728,N_2888);
nor U4087 (N_4087,N_1862,N_2165);
nand U4088 (N_4088,N_2451,N_1872);
xnor U4089 (N_4089,N_2677,N_2526);
nor U4090 (N_4090,N_2093,N_1927);
nand U4091 (N_4091,N_1863,N_1790);
or U4092 (N_4092,N_1927,N_2844);
or U4093 (N_4093,N_1830,N_2220);
or U4094 (N_4094,N_2057,N_2293);
or U4095 (N_4095,N_1678,N_2547);
xnor U4096 (N_4096,N_2613,N_2984);
or U4097 (N_4097,N_2587,N_1651);
and U4098 (N_4098,N_2346,N_2857);
nand U4099 (N_4099,N_2839,N_2964);
nand U4100 (N_4100,N_2101,N_2556);
nand U4101 (N_4101,N_2191,N_2332);
or U4102 (N_4102,N_2122,N_2604);
or U4103 (N_4103,N_1896,N_1933);
xor U4104 (N_4104,N_2269,N_1701);
or U4105 (N_4105,N_1624,N_2594);
nor U4106 (N_4106,N_1645,N_2437);
nand U4107 (N_4107,N_2193,N_1778);
or U4108 (N_4108,N_2714,N_2590);
nor U4109 (N_4109,N_2149,N_2460);
nand U4110 (N_4110,N_1590,N_2414);
nand U4111 (N_4111,N_2459,N_2595);
nand U4112 (N_4112,N_2810,N_2011);
xor U4113 (N_4113,N_2426,N_2603);
and U4114 (N_4114,N_2645,N_2395);
or U4115 (N_4115,N_2404,N_1610);
nand U4116 (N_4116,N_2339,N_1526);
and U4117 (N_4117,N_1996,N_1771);
nor U4118 (N_4118,N_2786,N_2373);
nand U4119 (N_4119,N_1622,N_2068);
nand U4120 (N_4120,N_2975,N_2775);
xor U4121 (N_4121,N_1619,N_2406);
or U4122 (N_4122,N_2745,N_2222);
nor U4123 (N_4123,N_1875,N_2138);
nor U4124 (N_4124,N_2373,N_2393);
xor U4125 (N_4125,N_2231,N_2852);
nand U4126 (N_4126,N_2005,N_2090);
xor U4127 (N_4127,N_1779,N_1953);
and U4128 (N_4128,N_1974,N_1869);
or U4129 (N_4129,N_2879,N_1586);
nor U4130 (N_4130,N_2722,N_1947);
xor U4131 (N_4131,N_2695,N_1748);
xnor U4132 (N_4132,N_1924,N_1941);
xor U4133 (N_4133,N_1695,N_2749);
nand U4134 (N_4134,N_2046,N_2118);
and U4135 (N_4135,N_1846,N_1864);
xnor U4136 (N_4136,N_2458,N_1741);
nand U4137 (N_4137,N_2191,N_2839);
and U4138 (N_4138,N_1549,N_2615);
and U4139 (N_4139,N_1621,N_1792);
nand U4140 (N_4140,N_1791,N_1811);
and U4141 (N_4141,N_2835,N_2038);
nor U4142 (N_4142,N_2451,N_2123);
nand U4143 (N_4143,N_2477,N_2936);
nand U4144 (N_4144,N_1640,N_2729);
or U4145 (N_4145,N_2089,N_2412);
and U4146 (N_4146,N_2009,N_2125);
and U4147 (N_4147,N_1873,N_2064);
and U4148 (N_4148,N_1809,N_2248);
xnor U4149 (N_4149,N_1585,N_1580);
nor U4150 (N_4150,N_2066,N_1703);
nand U4151 (N_4151,N_2399,N_2323);
nand U4152 (N_4152,N_1835,N_2836);
nand U4153 (N_4153,N_2024,N_2470);
xor U4154 (N_4154,N_2651,N_2778);
xor U4155 (N_4155,N_2706,N_2363);
xor U4156 (N_4156,N_1992,N_2203);
nand U4157 (N_4157,N_2563,N_2983);
nand U4158 (N_4158,N_1817,N_1571);
and U4159 (N_4159,N_2240,N_2975);
or U4160 (N_4160,N_1672,N_1610);
or U4161 (N_4161,N_2918,N_2171);
nor U4162 (N_4162,N_2688,N_2700);
or U4163 (N_4163,N_1600,N_2089);
nor U4164 (N_4164,N_2193,N_2263);
nand U4165 (N_4165,N_2001,N_1745);
xor U4166 (N_4166,N_2164,N_2536);
nor U4167 (N_4167,N_2363,N_2021);
nor U4168 (N_4168,N_1783,N_2640);
and U4169 (N_4169,N_2902,N_1863);
xor U4170 (N_4170,N_2844,N_1683);
nor U4171 (N_4171,N_2415,N_1551);
xor U4172 (N_4172,N_1603,N_2170);
xor U4173 (N_4173,N_2582,N_1923);
xor U4174 (N_4174,N_2753,N_2426);
or U4175 (N_4175,N_2611,N_2920);
xnor U4176 (N_4176,N_1745,N_2685);
or U4177 (N_4177,N_2339,N_2124);
nand U4178 (N_4178,N_1655,N_1596);
xor U4179 (N_4179,N_2841,N_2913);
nor U4180 (N_4180,N_1548,N_2362);
and U4181 (N_4181,N_2268,N_2783);
nand U4182 (N_4182,N_2069,N_2453);
xnor U4183 (N_4183,N_2929,N_1828);
nor U4184 (N_4184,N_1713,N_2396);
xnor U4185 (N_4185,N_2976,N_1919);
nand U4186 (N_4186,N_1559,N_2862);
nand U4187 (N_4187,N_2782,N_1601);
nor U4188 (N_4188,N_1847,N_1955);
nand U4189 (N_4189,N_1841,N_2749);
or U4190 (N_4190,N_1584,N_1950);
nand U4191 (N_4191,N_2796,N_1679);
nor U4192 (N_4192,N_2780,N_1740);
nor U4193 (N_4193,N_2281,N_2275);
nor U4194 (N_4194,N_2899,N_1623);
or U4195 (N_4195,N_1534,N_1685);
xor U4196 (N_4196,N_1548,N_1640);
nor U4197 (N_4197,N_2948,N_2637);
nand U4198 (N_4198,N_2614,N_1705);
nand U4199 (N_4199,N_2330,N_1760);
or U4200 (N_4200,N_2317,N_1941);
xor U4201 (N_4201,N_1559,N_2872);
and U4202 (N_4202,N_2319,N_2264);
nand U4203 (N_4203,N_2070,N_1843);
and U4204 (N_4204,N_2576,N_2565);
nand U4205 (N_4205,N_2626,N_2770);
nand U4206 (N_4206,N_1984,N_1818);
nor U4207 (N_4207,N_2898,N_2677);
or U4208 (N_4208,N_2192,N_2898);
and U4209 (N_4209,N_2456,N_2291);
nand U4210 (N_4210,N_2821,N_2957);
nor U4211 (N_4211,N_1839,N_1875);
nand U4212 (N_4212,N_2961,N_2907);
nor U4213 (N_4213,N_1577,N_2848);
and U4214 (N_4214,N_2921,N_2668);
xor U4215 (N_4215,N_2608,N_1676);
and U4216 (N_4216,N_2632,N_2654);
nand U4217 (N_4217,N_2516,N_2323);
nor U4218 (N_4218,N_2813,N_2211);
or U4219 (N_4219,N_2864,N_2613);
nand U4220 (N_4220,N_2170,N_1810);
xor U4221 (N_4221,N_1595,N_1743);
or U4222 (N_4222,N_2159,N_2744);
and U4223 (N_4223,N_1810,N_2260);
nand U4224 (N_4224,N_2514,N_2499);
or U4225 (N_4225,N_1583,N_2251);
and U4226 (N_4226,N_2279,N_2711);
nor U4227 (N_4227,N_2483,N_1549);
xor U4228 (N_4228,N_2034,N_2397);
or U4229 (N_4229,N_1728,N_2392);
or U4230 (N_4230,N_2508,N_2160);
and U4231 (N_4231,N_2865,N_1738);
nor U4232 (N_4232,N_1593,N_2752);
and U4233 (N_4233,N_2971,N_2859);
and U4234 (N_4234,N_2030,N_2923);
nand U4235 (N_4235,N_2431,N_2351);
or U4236 (N_4236,N_2771,N_2416);
nand U4237 (N_4237,N_2452,N_1510);
nor U4238 (N_4238,N_1581,N_2682);
and U4239 (N_4239,N_2797,N_2477);
nor U4240 (N_4240,N_2871,N_1638);
xnor U4241 (N_4241,N_1775,N_2697);
and U4242 (N_4242,N_2168,N_1628);
xnor U4243 (N_4243,N_1796,N_2669);
or U4244 (N_4244,N_2672,N_1668);
or U4245 (N_4245,N_1756,N_1955);
nor U4246 (N_4246,N_2957,N_2842);
or U4247 (N_4247,N_2124,N_1913);
xnor U4248 (N_4248,N_2770,N_1857);
nand U4249 (N_4249,N_2712,N_2820);
nand U4250 (N_4250,N_2152,N_1746);
nor U4251 (N_4251,N_1520,N_2950);
or U4252 (N_4252,N_2723,N_2264);
xor U4253 (N_4253,N_1739,N_2656);
and U4254 (N_4254,N_1513,N_2717);
and U4255 (N_4255,N_2879,N_2657);
or U4256 (N_4256,N_2736,N_2332);
and U4257 (N_4257,N_2522,N_2417);
xnor U4258 (N_4258,N_2142,N_2533);
xnor U4259 (N_4259,N_2431,N_1783);
xor U4260 (N_4260,N_2030,N_2804);
nand U4261 (N_4261,N_2380,N_2599);
nand U4262 (N_4262,N_1591,N_2471);
and U4263 (N_4263,N_1692,N_2887);
and U4264 (N_4264,N_2944,N_2009);
xor U4265 (N_4265,N_1709,N_2029);
or U4266 (N_4266,N_2744,N_1740);
and U4267 (N_4267,N_2960,N_2125);
nor U4268 (N_4268,N_2032,N_2895);
nor U4269 (N_4269,N_1703,N_2448);
or U4270 (N_4270,N_2428,N_1937);
xnor U4271 (N_4271,N_2004,N_2455);
nor U4272 (N_4272,N_2532,N_1781);
xnor U4273 (N_4273,N_2847,N_2698);
or U4274 (N_4274,N_2390,N_2491);
and U4275 (N_4275,N_1599,N_2541);
nand U4276 (N_4276,N_2215,N_2653);
xor U4277 (N_4277,N_2616,N_2568);
nand U4278 (N_4278,N_1953,N_2060);
nor U4279 (N_4279,N_2729,N_1882);
nand U4280 (N_4280,N_2086,N_2849);
xor U4281 (N_4281,N_2771,N_1706);
nand U4282 (N_4282,N_2231,N_2659);
nand U4283 (N_4283,N_1899,N_1630);
nand U4284 (N_4284,N_1699,N_2994);
and U4285 (N_4285,N_2831,N_2828);
xnor U4286 (N_4286,N_1730,N_2076);
xor U4287 (N_4287,N_2445,N_1946);
and U4288 (N_4288,N_1934,N_2189);
nor U4289 (N_4289,N_2032,N_2290);
nand U4290 (N_4290,N_2233,N_2121);
or U4291 (N_4291,N_2941,N_2980);
and U4292 (N_4292,N_1798,N_1594);
nand U4293 (N_4293,N_2539,N_2148);
nand U4294 (N_4294,N_1918,N_2690);
xnor U4295 (N_4295,N_2793,N_2707);
and U4296 (N_4296,N_2365,N_2875);
nand U4297 (N_4297,N_1671,N_2302);
and U4298 (N_4298,N_1976,N_1900);
xnor U4299 (N_4299,N_2448,N_1805);
and U4300 (N_4300,N_2295,N_1933);
nand U4301 (N_4301,N_1675,N_2856);
or U4302 (N_4302,N_2623,N_2588);
nor U4303 (N_4303,N_2740,N_2619);
nand U4304 (N_4304,N_2059,N_1823);
or U4305 (N_4305,N_2579,N_1800);
nor U4306 (N_4306,N_2112,N_1764);
and U4307 (N_4307,N_1941,N_2625);
xnor U4308 (N_4308,N_1599,N_2894);
or U4309 (N_4309,N_2008,N_2416);
nor U4310 (N_4310,N_1607,N_2882);
and U4311 (N_4311,N_2114,N_2676);
xnor U4312 (N_4312,N_2731,N_1822);
nor U4313 (N_4313,N_1649,N_1840);
nor U4314 (N_4314,N_2984,N_2447);
nand U4315 (N_4315,N_1606,N_2766);
nand U4316 (N_4316,N_2668,N_2152);
and U4317 (N_4317,N_2280,N_2618);
and U4318 (N_4318,N_2745,N_2690);
nor U4319 (N_4319,N_1662,N_2076);
nand U4320 (N_4320,N_2268,N_2623);
and U4321 (N_4321,N_2203,N_2206);
and U4322 (N_4322,N_2920,N_2479);
xor U4323 (N_4323,N_2968,N_1772);
nor U4324 (N_4324,N_1678,N_2866);
xnor U4325 (N_4325,N_2826,N_2943);
nand U4326 (N_4326,N_2439,N_1678);
nand U4327 (N_4327,N_2790,N_1629);
and U4328 (N_4328,N_2048,N_2621);
xnor U4329 (N_4329,N_2210,N_1721);
and U4330 (N_4330,N_1502,N_2956);
and U4331 (N_4331,N_1729,N_2256);
nor U4332 (N_4332,N_1523,N_2250);
and U4333 (N_4333,N_2846,N_2340);
nor U4334 (N_4334,N_2088,N_1972);
nor U4335 (N_4335,N_2132,N_2363);
nand U4336 (N_4336,N_2477,N_2004);
nor U4337 (N_4337,N_1590,N_2290);
or U4338 (N_4338,N_1879,N_2331);
nor U4339 (N_4339,N_2290,N_2475);
xnor U4340 (N_4340,N_1931,N_1522);
or U4341 (N_4341,N_2823,N_2346);
xnor U4342 (N_4342,N_2015,N_1790);
or U4343 (N_4343,N_2136,N_1735);
nor U4344 (N_4344,N_2654,N_1864);
xnor U4345 (N_4345,N_1525,N_2406);
and U4346 (N_4346,N_2459,N_2629);
nand U4347 (N_4347,N_1849,N_2464);
nor U4348 (N_4348,N_2834,N_1796);
and U4349 (N_4349,N_2074,N_2537);
or U4350 (N_4350,N_1845,N_2934);
nand U4351 (N_4351,N_2223,N_1695);
and U4352 (N_4352,N_2557,N_1597);
and U4353 (N_4353,N_2083,N_2327);
nor U4354 (N_4354,N_2283,N_1829);
xnor U4355 (N_4355,N_1755,N_2597);
xor U4356 (N_4356,N_2161,N_1555);
xnor U4357 (N_4357,N_2558,N_2628);
xor U4358 (N_4358,N_2357,N_2375);
nand U4359 (N_4359,N_2930,N_2987);
or U4360 (N_4360,N_2254,N_2120);
and U4361 (N_4361,N_2455,N_2069);
nor U4362 (N_4362,N_2717,N_2451);
and U4363 (N_4363,N_1648,N_1557);
or U4364 (N_4364,N_2360,N_1511);
xor U4365 (N_4365,N_1654,N_1664);
nand U4366 (N_4366,N_2914,N_2522);
xnor U4367 (N_4367,N_1732,N_1521);
and U4368 (N_4368,N_2649,N_2632);
nand U4369 (N_4369,N_1848,N_2421);
xnor U4370 (N_4370,N_1599,N_1500);
nand U4371 (N_4371,N_2333,N_2013);
nor U4372 (N_4372,N_1808,N_1747);
or U4373 (N_4373,N_1886,N_2643);
nand U4374 (N_4374,N_2504,N_2930);
nand U4375 (N_4375,N_2825,N_2197);
nand U4376 (N_4376,N_2781,N_2929);
xor U4377 (N_4377,N_1832,N_1985);
nor U4378 (N_4378,N_2511,N_2797);
nand U4379 (N_4379,N_2278,N_2242);
nor U4380 (N_4380,N_1554,N_2908);
nor U4381 (N_4381,N_1583,N_2731);
nor U4382 (N_4382,N_2372,N_1869);
nand U4383 (N_4383,N_2803,N_1772);
xnor U4384 (N_4384,N_2360,N_1621);
and U4385 (N_4385,N_2873,N_2598);
and U4386 (N_4386,N_2483,N_2650);
or U4387 (N_4387,N_2725,N_2798);
and U4388 (N_4388,N_2878,N_2714);
nor U4389 (N_4389,N_2206,N_1937);
and U4390 (N_4390,N_1749,N_2935);
xnor U4391 (N_4391,N_2968,N_1930);
xor U4392 (N_4392,N_1528,N_2009);
nand U4393 (N_4393,N_1951,N_1856);
or U4394 (N_4394,N_2540,N_2946);
or U4395 (N_4395,N_1782,N_1770);
or U4396 (N_4396,N_2192,N_2529);
and U4397 (N_4397,N_2181,N_2904);
and U4398 (N_4398,N_2435,N_2102);
and U4399 (N_4399,N_2274,N_1713);
and U4400 (N_4400,N_2640,N_2304);
and U4401 (N_4401,N_2627,N_1747);
nand U4402 (N_4402,N_2033,N_1514);
and U4403 (N_4403,N_1542,N_1620);
and U4404 (N_4404,N_2528,N_1868);
xnor U4405 (N_4405,N_2528,N_2062);
xnor U4406 (N_4406,N_2049,N_2291);
nand U4407 (N_4407,N_1698,N_2969);
xor U4408 (N_4408,N_2421,N_1578);
and U4409 (N_4409,N_1731,N_1738);
or U4410 (N_4410,N_2334,N_2107);
nor U4411 (N_4411,N_2626,N_2519);
xor U4412 (N_4412,N_1744,N_2001);
nand U4413 (N_4413,N_2684,N_1646);
or U4414 (N_4414,N_1978,N_2838);
or U4415 (N_4415,N_2726,N_2333);
xor U4416 (N_4416,N_2030,N_2398);
and U4417 (N_4417,N_2106,N_2906);
and U4418 (N_4418,N_1906,N_2600);
nor U4419 (N_4419,N_2655,N_2212);
or U4420 (N_4420,N_2742,N_1818);
xor U4421 (N_4421,N_2850,N_2354);
nor U4422 (N_4422,N_2967,N_1869);
xnor U4423 (N_4423,N_2325,N_2028);
nor U4424 (N_4424,N_1799,N_2488);
nor U4425 (N_4425,N_2772,N_2573);
nor U4426 (N_4426,N_2754,N_1521);
nor U4427 (N_4427,N_2079,N_2537);
xnor U4428 (N_4428,N_2635,N_2761);
nand U4429 (N_4429,N_2415,N_1754);
nand U4430 (N_4430,N_2279,N_1849);
and U4431 (N_4431,N_2907,N_1994);
or U4432 (N_4432,N_2415,N_2074);
nor U4433 (N_4433,N_1728,N_2872);
nor U4434 (N_4434,N_1968,N_2091);
nand U4435 (N_4435,N_2039,N_1573);
nor U4436 (N_4436,N_2660,N_2623);
and U4437 (N_4437,N_2346,N_1969);
nor U4438 (N_4438,N_1722,N_1762);
nor U4439 (N_4439,N_2500,N_1667);
nor U4440 (N_4440,N_2871,N_1730);
or U4441 (N_4441,N_2901,N_2539);
xor U4442 (N_4442,N_1596,N_1574);
nand U4443 (N_4443,N_1777,N_2635);
or U4444 (N_4444,N_2969,N_2996);
nand U4445 (N_4445,N_2245,N_2516);
and U4446 (N_4446,N_2288,N_2619);
nor U4447 (N_4447,N_2892,N_1830);
or U4448 (N_4448,N_2860,N_2952);
nor U4449 (N_4449,N_2111,N_1810);
nand U4450 (N_4450,N_1770,N_1534);
xnor U4451 (N_4451,N_1824,N_1852);
or U4452 (N_4452,N_2984,N_1810);
xnor U4453 (N_4453,N_1579,N_1701);
and U4454 (N_4454,N_2028,N_2550);
or U4455 (N_4455,N_1989,N_2718);
xor U4456 (N_4456,N_2524,N_2525);
and U4457 (N_4457,N_1511,N_2245);
xnor U4458 (N_4458,N_2191,N_1629);
and U4459 (N_4459,N_2587,N_1878);
and U4460 (N_4460,N_2845,N_1620);
xnor U4461 (N_4461,N_2629,N_2528);
xnor U4462 (N_4462,N_2816,N_2199);
xnor U4463 (N_4463,N_1529,N_2828);
and U4464 (N_4464,N_2187,N_2106);
nand U4465 (N_4465,N_2204,N_2149);
nor U4466 (N_4466,N_1875,N_2848);
and U4467 (N_4467,N_2313,N_2251);
or U4468 (N_4468,N_2271,N_2792);
xnor U4469 (N_4469,N_2831,N_2139);
xor U4470 (N_4470,N_2212,N_2729);
or U4471 (N_4471,N_2616,N_1931);
and U4472 (N_4472,N_2890,N_2766);
nor U4473 (N_4473,N_1589,N_2282);
nand U4474 (N_4474,N_2656,N_2907);
xnor U4475 (N_4475,N_2504,N_2490);
nor U4476 (N_4476,N_2902,N_2008);
xnor U4477 (N_4477,N_1660,N_1560);
xnor U4478 (N_4478,N_2402,N_2382);
nor U4479 (N_4479,N_1903,N_1844);
or U4480 (N_4480,N_1990,N_2475);
nor U4481 (N_4481,N_1738,N_2097);
or U4482 (N_4482,N_1976,N_2595);
nand U4483 (N_4483,N_2522,N_1706);
or U4484 (N_4484,N_2632,N_1699);
and U4485 (N_4485,N_1849,N_1952);
and U4486 (N_4486,N_2621,N_1842);
or U4487 (N_4487,N_2813,N_2100);
nand U4488 (N_4488,N_1653,N_2567);
or U4489 (N_4489,N_1791,N_2979);
or U4490 (N_4490,N_2045,N_1677);
nor U4491 (N_4491,N_1635,N_1676);
and U4492 (N_4492,N_2926,N_2700);
nor U4493 (N_4493,N_2016,N_1924);
nand U4494 (N_4494,N_2363,N_1514);
and U4495 (N_4495,N_1734,N_1589);
or U4496 (N_4496,N_1720,N_2754);
and U4497 (N_4497,N_2785,N_1989);
nand U4498 (N_4498,N_2364,N_2979);
nor U4499 (N_4499,N_1708,N_2452);
nor U4500 (N_4500,N_3061,N_3777);
xnor U4501 (N_4501,N_3045,N_3519);
nand U4502 (N_4502,N_4201,N_3356);
or U4503 (N_4503,N_3640,N_3718);
nand U4504 (N_4504,N_3047,N_4239);
nor U4505 (N_4505,N_3533,N_4160);
nor U4506 (N_4506,N_3331,N_3340);
nor U4507 (N_4507,N_3011,N_3075);
xnor U4508 (N_4508,N_3716,N_4045);
or U4509 (N_4509,N_3135,N_3231);
and U4510 (N_4510,N_3570,N_3407);
nor U4511 (N_4511,N_3031,N_3485);
nand U4512 (N_4512,N_3264,N_3470);
nor U4513 (N_4513,N_3861,N_4063);
nand U4514 (N_4514,N_4169,N_3541);
and U4515 (N_4515,N_3741,N_3580);
and U4516 (N_4516,N_3935,N_4479);
xor U4517 (N_4517,N_4498,N_3621);
or U4518 (N_4518,N_3902,N_3066);
or U4519 (N_4519,N_4228,N_3128);
nor U4520 (N_4520,N_3280,N_3478);
and U4521 (N_4521,N_4319,N_3414);
xnor U4522 (N_4522,N_3582,N_4387);
nand U4523 (N_4523,N_3295,N_3753);
nand U4524 (N_4524,N_3700,N_4062);
or U4525 (N_4525,N_3729,N_3086);
and U4526 (N_4526,N_3088,N_3446);
or U4527 (N_4527,N_4263,N_4171);
xor U4528 (N_4528,N_3991,N_3392);
xor U4529 (N_4529,N_3471,N_4165);
xnor U4530 (N_4530,N_3746,N_3337);
nand U4531 (N_4531,N_3082,N_3821);
and U4532 (N_4532,N_3444,N_4240);
nand U4533 (N_4533,N_4312,N_4475);
or U4534 (N_4534,N_3701,N_3794);
and U4535 (N_4535,N_3968,N_4452);
and U4536 (N_4536,N_4442,N_3758);
or U4537 (N_4537,N_4107,N_3002);
or U4538 (N_4538,N_3532,N_4185);
nor U4539 (N_4539,N_4279,N_4249);
xnor U4540 (N_4540,N_3297,N_3030);
nand U4541 (N_4541,N_4294,N_4035);
and U4542 (N_4542,N_4032,N_3069);
xnor U4543 (N_4543,N_4433,N_3559);
and U4544 (N_4544,N_3327,N_4087);
nand U4545 (N_4545,N_3373,N_3574);
or U4546 (N_4546,N_4235,N_3464);
or U4547 (N_4547,N_4344,N_3008);
xnor U4548 (N_4548,N_4018,N_4441);
or U4549 (N_4549,N_3497,N_3060);
and U4550 (N_4550,N_3209,N_3742);
nor U4551 (N_4551,N_4450,N_4411);
and U4552 (N_4552,N_4264,N_3428);
or U4553 (N_4553,N_3304,N_3308);
or U4554 (N_4554,N_4334,N_3397);
xnor U4555 (N_4555,N_3710,N_3143);
nand U4556 (N_4556,N_3517,N_4400);
nand U4557 (N_4557,N_4280,N_3313);
nor U4558 (N_4558,N_3423,N_4406);
or U4559 (N_4559,N_3661,N_3554);
nor U4560 (N_4560,N_3715,N_3359);
and U4561 (N_4561,N_3546,N_3665);
xnor U4562 (N_4562,N_4446,N_3711);
and U4563 (N_4563,N_3638,N_4190);
nand U4564 (N_4564,N_4285,N_4421);
xnor U4565 (N_4565,N_4218,N_4477);
or U4566 (N_4566,N_4157,N_4170);
nand U4567 (N_4567,N_4305,N_3368);
or U4568 (N_4568,N_3823,N_4156);
xor U4569 (N_4569,N_3744,N_3169);
nand U4570 (N_4570,N_3605,N_3595);
and U4571 (N_4571,N_3867,N_3402);
or U4572 (N_4572,N_3674,N_3697);
or U4573 (N_4573,N_4448,N_3856);
nand U4574 (N_4574,N_4242,N_3918);
or U4575 (N_4575,N_4260,N_3781);
xnor U4576 (N_4576,N_3599,N_3800);
and U4577 (N_4577,N_3081,N_3147);
xor U4578 (N_4578,N_4230,N_3571);
nor U4579 (N_4579,N_3680,N_3145);
xor U4580 (N_4580,N_4451,N_4435);
or U4581 (N_4581,N_4168,N_3142);
xnor U4582 (N_4582,N_4496,N_3185);
nand U4583 (N_4583,N_4091,N_3849);
nand U4584 (N_4584,N_3797,N_4426);
nor U4585 (N_4585,N_4237,N_3287);
nand U4586 (N_4586,N_4164,N_3358);
or U4587 (N_4587,N_4017,N_3321);
nor U4588 (N_4588,N_3986,N_4343);
nor U4589 (N_4589,N_3490,N_4323);
and U4590 (N_4590,N_3527,N_3853);
nor U4591 (N_4591,N_3178,N_3237);
or U4592 (N_4592,N_3537,N_3581);
xnor U4593 (N_4593,N_3730,N_3482);
nand U4594 (N_4594,N_3585,N_3854);
or U4595 (N_4595,N_3884,N_3051);
or U4596 (N_4596,N_3474,N_4487);
nor U4597 (N_4597,N_3175,N_4161);
nand U4598 (N_4598,N_4346,N_4302);
or U4599 (N_4599,N_4311,N_4256);
and U4600 (N_4600,N_3070,N_4047);
and U4601 (N_4601,N_3450,N_3090);
xor U4602 (N_4602,N_3534,N_3488);
and U4603 (N_4603,N_3468,N_4153);
or U4604 (N_4604,N_4268,N_3545);
nor U4605 (N_4605,N_3767,N_4083);
and U4606 (N_4606,N_4104,N_3977);
xnor U4607 (N_4607,N_3370,N_4076);
or U4608 (N_4608,N_3310,N_3606);
nand U4609 (N_4609,N_3187,N_3910);
and U4610 (N_4610,N_4024,N_3641);
or U4611 (N_4611,N_4174,N_3926);
or U4612 (N_4612,N_3860,N_3072);
xor U4613 (N_4613,N_3372,N_3735);
or U4614 (N_4614,N_3350,N_4310);
xor U4615 (N_4615,N_3965,N_3673);
and U4616 (N_4616,N_3939,N_3314);
nor U4617 (N_4617,N_4222,N_3834);
nor U4618 (N_4618,N_3924,N_3165);
nor U4619 (N_4619,N_3726,N_3500);
and U4620 (N_4620,N_4288,N_3333);
and U4621 (N_4621,N_3874,N_4291);
nor U4622 (N_4622,N_4490,N_3593);
or U4623 (N_4623,N_4234,N_4395);
and U4624 (N_4624,N_3908,N_4392);
nand U4625 (N_4625,N_3870,N_4281);
xor U4626 (N_4626,N_3614,N_4079);
xor U4627 (N_4627,N_3162,N_4103);
nand U4628 (N_4628,N_4040,N_3698);
nor U4629 (N_4629,N_3424,N_4245);
nor U4630 (N_4630,N_3062,N_3583);
nand U4631 (N_4631,N_3686,N_4223);
or U4632 (N_4632,N_3899,N_3651);
or U4633 (N_4633,N_3003,N_3109);
nand U4634 (N_4634,N_3415,N_3524);
xnor U4635 (N_4635,N_3666,N_3754);
nor U4636 (N_4636,N_3448,N_3938);
and U4637 (N_4637,N_4116,N_3303);
nor U4638 (N_4638,N_3477,N_4162);
nand U4639 (N_4639,N_4020,N_4105);
or U4640 (N_4640,N_3085,N_3851);
nand U4641 (N_4641,N_3877,N_3612);
nor U4642 (N_4642,N_3865,N_3630);
nor U4643 (N_4643,N_4365,N_3844);
xor U4644 (N_4644,N_3367,N_3118);
nand U4645 (N_4645,N_3930,N_3181);
or U4646 (N_4646,N_3039,N_3048);
nand U4647 (N_4647,N_4275,N_3804);
nand U4648 (N_4648,N_4422,N_3891);
nand U4649 (N_4649,N_3025,N_3852);
xor U4650 (N_4650,N_3598,N_3608);
nor U4651 (N_4651,N_4283,N_3133);
and U4652 (N_4652,N_3012,N_3094);
xnor U4653 (N_4653,N_4316,N_3915);
xnor U4654 (N_4654,N_3761,N_3171);
or U4655 (N_4655,N_3845,N_3670);
or U4656 (N_4656,N_3576,N_3602);
xor U4657 (N_4657,N_3422,N_4251);
or U4658 (N_4658,N_3139,N_3998);
nor U4659 (N_4659,N_3572,N_4243);
nand U4660 (N_4660,N_3548,N_3360);
nand U4661 (N_4661,N_3769,N_4369);
nand U4662 (N_4662,N_3243,N_4296);
xor U4663 (N_4663,N_3880,N_3179);
nor U4664 (N_4664,N_3200,N_3018);
nor U4665 (N_4665,N_4039,N_3239);
xor U4666 (N_4666,N_3273,N_3659);
and U4667 (N_4667,N_3232,N_3839);
xor U4668 (N_4668,N_3288,N_3033);
xor U4669 (N_4669,N_3398,N_3996);
nor U4670 (N_4670,N_4466,N_3087);
nor U4671 (N_4671,N_4207,N_4217);
nor U4672 (N_4672,N_3774,N_3704);
and U4673 (N_4673,N_3250,N_3929);
xor U4674 (N_4674,N_4350,N_3124);
nand U4675 (N_4675,N_3238,N_3530);
nor U4676 (N_4676,N_4413,N_4154);
and U4677 (N_4677,N_4423,N_4238);
nor U4678 (N_4678,N_3151,N_3026);
xnor U4679 (N_4679,N_4071,N_3543);
nor U4680 (N_4680,N_3125,N_3395);
nor U4681 (N_4681,N_3771,N_4183);
xnor U4682 (N_4682,N_3636,N_3654);
xnor U4683 (N_4683,N_3903,N_3084);
and U4684 (N_4684,N_3649,N_4467);
or U4685 (N_4685,N_4236,N_4147);
or U4686 (N_4686,N_3235,N_3436);
and U4687 (N_4687,N_4341,N_4026);
nand U4688 (N_4688,N_3172,N_3529);
xor U4689 (N_4689,N_3315,N_4059);
or U4690 (N_4690,N_4025,N_3432);
xor U4691 (N_4691,N_4122,N_4070);
and U4692 (N_4692,N_3551,N_4182);
xnor U4693 (N_4693,N_3343,N_3378);
nor U4694 (N_4694,N_4011,N_3967);
nor U4695 (N_4695,N_3879,N_3285);
nor U4696 (N_4696,N_4282,N_3840);
or U4697 (N_4697,N_3400,N_3078);
nand U4698 (N_4698,N_4057,N_3672);
xnor U4699 (N_4699,N_3346,N_3847);
xnor U4700 (N_4700,N_3719,N_3153);
or U4701 (N_4701,N_4353,N_3245);
nor U4702 (N_4702,N_4370,N_3311);
xnor U4703 (N_4703,N_3679,N_3341);
and U4704 (N_4704,N_3705,N_4376);
nor U4705 (N_4705,N_3951,N_4072);
nor U4706 (N_4706,N_3765,N_3740);
xnor U4707 (N_4707,N_3150,N_3755);
xor U4708 (N_4708,N_3055,N_4273);
and U4709 (N_4709,N_3380,N_4257);
xnor U4710 (N_4710,N_3878,N_3960);
and U4711 (N_4711,N_3152,N_3412);
nand U4712 (N_4712,N_3693,N_3463);
xor U4713 (N_4713,N_4480,N_3149);
nand U4714 (N_4714,N_3272,N_4187);
xor U4715 (N_4715,N_3688,N_3540);
and U4716 (N_4716,N_3105,N_3695);
nor U4717 (N_4717,N_4494,N_3509);
and U4718 (N_4718,N_3587,N_4227);
nor U4719 (N_4719,N_3566,N_3024);
nor U4720 (N_4720,N_4184,N_3071);
nor U4721 (N_4721,N_4194,N_3508);
or U4722 (N_4722,N_4219,N_3364);
nand U4723 (N_4723,N_4088,N_4068);
nor U4724 (N_4724,N_4050,N_3589);
nand U4725 (N_4725,N_4061,N_3469);
xnor U4726 (N_4726,N_3106,N_3473);
and U4727 (N_4727,N_3757,N_4358);
or U4728 (N_4728,N_3732,N_3010);
nand U4729 (N_4729,N_4377,N_3167);
nand U4730 (N_4730,N_3776,N_4014);
nand U4731 (N_4731,N_3591,N_3305);
or U4732 (N_4732,N_3057,N_3379);
and U4733 (N_4733,N_3480,N_3934);
and U4734 (N_4734,N_3338,N_3259);
or U4735 (N_4735,N_4175,N_3980);
xor U4736 (N_4736,N_4054,N_3351);
xor U4737 (N_4737,N_3345,N_3882);
or U4738 (N_4738,N_3901,N_4259);
nor U4739 (N_4739,N_4144,N_3000);
xnor U4740 (N_4740,N_3969,N_4159);
and U4741 (N_4741,N_4383,N_3644);
xor U4742 (N_4742,N_4179,N_4155);
or U4743 (N_4743,N_3743,N_3042);
xor U4744 (N_4744,N_3898,N_3846);
xor U4745 (N_4745,N_3021,N_3481);
and U4746 (N_4746,N_3933,N_3099);
and U4747 (N_4747,N_3843,N_3044);
nor U4748 (N_4748,N_3881,N_3390);
nand U4749 (N_4749,N_4007,N_4188);
xnor U4750 (N_4750,N_4108,N_4386);
nand U4751 (N_4751,N_3760,N_4030);
nor U4752 (N_4752,N_4118,N_3076);
nor U4753 (N_4753,N_3067,N_3095);
nor U4754 (N_4754,N_3535,N_3435);
nand U4755 (N_4755,N_3862,N_3332);
nor U4756 (N_4756,N_3452,N_4145);
nand U4757 (N_4757,N_3258,N_3984);
nand U4758 (N_4758,N_3749,N_3676);
and U4759 (N_4759,N_3274,N_3159);
or U4760 (N_4760,N_3586,N_4390);
nor U4761 (N_4761,N_4396,N_3208);
xor U4762 (N_4762,N_3841,N_3850);
nor U4763 (N_4763,N_3941,N_4348);
nor U4764 (N_4764,N_4093,N_3352);
and U4765 (N_4765,N_3648,N_3079);
xor U4766 (N_4766,N_3815,N_4409);
or U4767 (N_4767,N_4089,N_3093);
nand U4768 (N_4768,N_3056,N_4081);
nand U4769 (N_4769,N_4455,N_3455);
and U4770 (N_4770,N_3203,N_3063);
nor U4771 (N_4771,N_3563,N_3161);
nand U4772 (N_4772,N_3410,N_3706);
or U4773 (N_4773,N_3122,N_4364);
nand U4774 (N_4774,N_3928,N_4028);
and U4775 (N_4775,N_3652,N_4456);
nand U4776 (N_4776,N_3600,N_3868);
nand U4777 (N_4777,N_4331,N_3445);
nor U4778 (N_4778,N_3229,N_3836);
nand U4779 (N_4779,N_4199,N_3687);
or U4780 (N_4780,N_4332,N_4158);
nand U4781 (N_4781,N_3459,N_3756);
nand U4782 (N_4782,N_4382,N_4313);
xor U4783 (N_4783,N_3956,N_4482);
nor U4784 (N_4784,N_4053,N_3032);
or U4785 (N_4785,N_3073,N_3279);
or U4786 (N_4786,N_4261,N_3731);
xnor U4787 (N_4787,N_3792,N_4074);
nor U4788 (N_4788,N_4287,N_4385);
and U4789 (N_4789,N_3752,N_3819);
or U4790 (N_4790,N_3317,N_4394);
and U4791 (N_4791,N_3027,N_3855);
and U4792 (N_4792,N_4033,N_4203);
and U4793 (N_4793,N_3068,N_4241);
and U4794 (N_4794,N_3883,N_3363);
nor U4795 (N_4795,N_3344,N_3022);
xnor U4796 (N_4796,N_4135,N_3694);
xnor U4797 (N_4797,N_4330,N_3268);
nand U4798 (N_4798,N_4002,N_4212);
nor U4799 (N_4799,N_3489,N_3427);
nor U4800 (N_4800,N_3875,N_3971);
or U4801 (N_4801,N_3816,N_3290);
nor U4802 (N_4802,N_3342,N_3461);
nand U4803 (N_4803,N_3584,N_3246);
nor U4804 (N_4804,N_3919,N_4274);
nand U4805 (N_4805,N_4021,N_3049);
xor U4806 (N_4806,N_4408,N_3725);
nor U4807 (N_4807,N_3194,N_3871);
and U4808 (N_4808,N_3872,N_3275);
or U4809 (N_4809,N_4085,N_3437);
nor U4810 (N_4810,N_3552,N_4109);
and U4811 (N_4811,N_4379,N_4225);
nand U4812 (N_4812,N_3997,N_3615);
nand U4813 (N_4813,N_3449,N_3675);
nor U4814 (N_4814,N_3521,N_3727);
nor U4815 (N_4815,N_3498,N_3708);
and U4816 (N_4816,N_4173,N_3683);
nand U4817 (N_4817,N_3629,N_4078);
xor U4818 (N_4818,N_3092,N_3191);
or U4819 (N_4819,N_4058,N_3923);
and U4820 (N_4820,N_3283,N_3005);
or U4821 (N_4821,N_4129,N_3361);
or U4822 (N_4822,N_3945,N_4132);
or U4823 (N_4823,N_3828,N_3594);
nand U4824 (N_4824,N_4042,N_4397);
nor U4825 (N_4825,N_3416,N_4029);
nor U4826 (N_4826,N_4447,N_3329);
xnor U4827 (N_4827,N_4428,N_4403);
nor U4828 (N_4828,N_3177,N_4003);
xor U4829 (N_4829,N_4101,N_4134);
nand U4830 (N_4830,N_4492,N_4143);
xor U4831 (N_4831,N_4300,N_3182);
and U4832 (N_4832,N_3100,N_4196);
nand U4833 (N_4833,N_4216,N_3964);
nand U4834 (N_4834,N_4112,N_3221);
nand U4835 (N_4835,N_3322,N_3146);
nand U4836 (N_4836,N_4202,N_3038);
nor U4837 (N_4837,N_3714,N_3262);
xor U4838 (N_4838,N_4244,N_3210);
or U4839 (N_4839,N_4205,N_4363);
and U4840 (N_4840,N_4306,N_3616);
nor U4841 (N_4841,N_3399,N_4084);
and U4842 (N_4842,N_3573,N_4270);
nand U4843 (N_4843,N_3296,N_3466);
and U4844 (N_4844,N_3721,N_3016);
nor U4845 (N_4845,N_3788,N_3226);
or U4846 (N_4846,N_4056,N_3827);
and U4847 (N_4847,N_3544,N_3479);
nor U4848 (N_4848,N_3864,N_3417);
xor U4849 (N_4849,N_4307,N_3357);
nand U4850 (N_4850,N_4473,N_3822);
or U4851 (N_4851,N_3408,N_3491);
or U4852 (N_4852,N_3431,N_4404);
xnor U4853 (N_4853,N_3190,N_4110);
or U4854 (N_4854,N_4362,N_3838);
nor U4855 (N_4855,N_3457,N_3601);
nor U4856 (N_4856,N_4258,N_3983);
nor U4857 (N_4857,N_3512,N_4317);
and U4858 (N_4858,N_4192,N_3269);
or U4859 (N_4859,N_3646,N_4342);
nor U4860 (N_4860,N_4130,N_3227);
xor U4861 (N_4861,N_3294,N_4460);
nand U4862 (N_4862,N_4303,N_4119);
or U4863 (N_4863,N_3325,N_3383);
nor U4864 (N_4864,N_3242,N_3734);
nand U4865 (N_4865,N_3801,N_3837);
xor U4866 (N_4866,N_3669,N_3204);
or U4867 (N_4867,N_3212,N_4139);
nand U4868 (N_4868,N_4338,N_3438);
or U4869 (N_4869,N_3728,N_3347);
nor U4870 (N_4870,N_3456,N_4172);
nand U4871 (N_4871,N_3810,N_4100);
xnor U4872 (N_4872,N_3957,N_4246);
nor U4873 (N_4873,N_3298,N_3324);
nor U4874 (N_4874,N_3766,N_4340);
nand U4875 (N_4875,N_3270,N_3326);
or U4876 (N_4876,N_3265,N_4361);
or U4877 (N_4877,N_3775,N_3798);
nor U4878 (N_4878,N_4027,N_4320);
nand U4879 (N_4879,N_3975,N_3739);
and U4880 (N_4880,N_4360,N_4146);
and U4881 (N_4881,N_3394,N_3107);
nand U4882 (N_4882,N_3558,N_3206);
xor U4883 (N_4883,N_3634,N_4124);
and U4884 (N_4884,N_4372,N_3216);
xor U4885 (N_4885,N_3017,N_3195);
or U4886 (N_4886,N_3240,N_3958);
nand U4887 (N_4887,N_4166,N_3434);
nand U4888 (N_4888,N_4462,N_3820);
nor U4889 (N_4889,N_3873,N_3993);
nor U4890 (N_4890,N_3130,N_3707);
nand U4891 (N_4891,N_3978,N_3131);
xnor U4892 (N_4892,N_3323,N_4200);
and U4893 (N_4893,N_3685,N_3885);
nand U4894 (N_4894,N_3318,N_3931);
nand U4895 (N_4895,N_4284,N_3230);
and U4896 (N_4896,N_3577,N_3413);
nor U4897 (N_4897,N_3132,N_4254);
xnor U4898 (N_4898,N_3531,N_4438);
and U4899 (N_4899,N_3702,N_4095);
or U4900 (N_4900,N_4314,N_4111);
nand U4901 (N_4901,N_3163,N_3103);
xor U4902 (N_4902,N_3738,N_4416);
and U4903 (N_4903,N_3371,N_3202);
nor U4904 (N_4904,N_4044,N_4125);
and U4905 (N_4905,N_3897,N_3476);
or U4906 (N_4906,N_3117,N_3029);
nand U4907 (N_4907,N_4335,N_3953);
nor U4908 (N_4908,N_3513,N_3515);
or U4909 (N_4909,N_3691,N_3014);
nand U4910 (N_4910,N_3451,N_3458);
nor U4911 (N_4911,N_4427,N_3950);
or U4912 (N_4912,N_3058,N_3336);
and U4913 (N_4913,N_3035,N_3406);
and U4914 (N_4914,N_3759,N_4276);
xor U4915 (N_4915,N_3900,N_3170);
or U4916 (N_4916,N_3557,N_3618);
or U4917 (N_4917,N_4493,N_3825);
nor U4918 (N_4918,N_3909,N_4214);
or U4919 (N_4919,N_3790,N_3401);
and U4920 (N_4920,N_4001,N_4009);
nand U4921 (N_4921,N_3981,N_3192);
nand U4922 (N_4922,N_3405,N_4272);
xnor U4923 (N_4923,N_3442,N_3927);
or U4924 (N_4924,N_4255,N_3905);
and U4925 (N_4925,N_4265,N_3144);
xnor U4926 (N_4926,N_3522,N_4469);
or U4927 (N_4927,N_3813,N_3539);
nor U4928 (N_4928,N_3604,N_3034);
xnor U4929 (N_4929,N_3526,N_3116);
or U4930 (N_4930,N_3830,N_3328);
nand U4931 (N_4931,N_3940,N_3793);
or U4932 (N_4932,N_3656,N_3462);
xnor U4933 (N_4933,N_3050,N_3660);
nand U4934 (N_4934,N_3858,N_4015);
nor U4935 (N_4935,N_4399,N_3703);
nand U4936 (N_4936,N_3538,N_4380);
nand U4937 (N_4937,N_4049,N_3579);
or U4938 (N_4938,N_4419,N_3465);
nand U4939 (N_4939,N_3440,N_3631);
nand U4940 (N_4940,N_3036,N_3890);
or U4941 (N_4941,N_4149,N_3886);
nand U4942 (N_4942,N_3712,N_3257);
nor U4943 (N_4943,N_3101,N_3963);
nand U4944 (N_4944,N_3492,N_4407);
nand U4945 (N_4945,N_3653,N_3366);
nand U4946 (N_4946,N_3300,N_3976);
and U4947 (N_4947,N_3420,N_4453);
and U4948 (N_4948,N_3484,N_4293);
nor U4949 (N_4949,N_3320,N_4191);
xor U4950 (N_4950,N_3426,N_3542);
or U4951 (N_4951,N_4444,N_4131);
nor U4952 (N_4952,N_3809,N_4333);
nor U4953 (N_4953,N_3138,N_4461);
nand U4954 (N_4954,N_3803,N_3682);
and U4955 (N_4955,N_3080,N_3013);
nand U4956 (N_4956,N_4412,N_4378);
or U4957 (N_4957,N_3511,N_4470);
and U4958 (N_4958,N_4297,N_4204);
or U4959 (N_4959,N_4048,N_3115);
and U4960 (N_4960,N_3944,N_3111);
nand U4961 (N_4961,N_3833,N_3805);
xor U4962 (N_4962,N_3421,N_4367);
nor U4963 (N_4963,N_3550,N_4292);
xor U4964 (N_4964,N_4064,N_3737);
xor U4965 (N_4965,N_4324,N_3733);
nand U4966 (N_4966,N_3388,N_3353);
xor U4967 (N_4967,N_3689,N_4349);
or U4968 (N_4968,N_4247,N_3617);
nand U4969 (N_4969,N_4253,N_4114);
and U4970 (N_4970,N_4278,N_3110);
or U4971 (N_4971,N_3525,N_3633);
or U4972 (N_4972,N_4373,N_3842);
nand U4973 (N_4973,N_3486,N_4233);
and U4974 (N_4974,N_3921,N_3988);
or U4975 (N_4975,N_4037,N_3610);
nor U4976 (N_4976,N_3425,N_4208);
nand U4977 (N_4977,N_3772,N_3947);
nand U4978 (N_4978,N_4354,N_3102);
nand U4979 (N_4979,N_4034,N_3009);
nand U4980 (N_4980,N_3176,N_3876);
nor U4981 (N_4981,N_3244,N_4420);
and U4982 (N_4982,N_3453,N_4352);
nand U4983 (N_4983,N_4000,N_3104);
and U4984 (N_4984,N_3795,N_4471);
xnor U4985 (N_4985,N_3385,N_3982);
xor U4986 (N_4986,N_3113,N_3037);
or U4987 (N_4987,N_3271,N_4478);
xnor U4988 (N_4988,N_3065,N_3384);
or U4989 (N_4989,N_4491,N_3785);
xor U4990 (N_4990,N_4266,N_3796);
xor U4991 (N_4991,N_4289,N_4468);
nor U4992 (N_4992,N_4345,N_3374);
xnor U4993 (N_4993,N_4115,N_3791);
xnor U4994 (N_4994,N_3946,N_3916);
xnor U4995 (N_4995,N_4359,N_3354);
nor U4996 (N_4996,N_3291,N_3904);
nor U4997 (N_4997,N_3677,N_3409);
or U4998 (N_4998,N_4356,N_3207);
nor U4999 (N_4999,N_3779,N_4389);
or U5000 (N_5000,N_4141,N_3657);
nand U5001 (N_5001,N_3282,N_4424);
and U5002 (N_5002,N_4454,N_3783);
nand U5003 (N_5003,N_3655,N_3504);
nand U5004 (N_5004,N_3365,N_3632);
or U5005 (N_5005,N_4436,N_3948);
nor U5006 (N_5006,N_4123,N_3808);
nand U5007 (N_5007,N_4133,N_3668);
nor U5008 (N_5008,N_3914,N_3764);
or U5009 (N_5009,N_3699,N_4295);
nand U5010 (N_5010,N_3222,N_3955);
nand U5011 (N_5011,N_3812,N_4038);
or U5012 (N_5012,N_3995,N_4195);
or U5013 (N_5013,N_4298,N_3134);
or U5014 (N_5014,N_3619,N_4121);
or U5015 (N_5015,N_3119,N_3937);
or U5016 (N_5016,N_4277,N_4004);
xor U5017 (N_5017,N_3166,N_3164);
nand U5018 (N_5018,N_3639,N_3289);
xor U5019 (N_5019,N_3089,N_3911);
nand U5020 (N_5020,N_4069,N_3198);
nor U5021 (N_5021,N_3369,N_3496);
or U5022 (N_5022,N_3319,N_3807);
xor U5023 (N_5023,N_3748,N_3802);
nor U5024 (N_5024,N_4055,N_3624);
or U5025 (N_5025,N_3989,N_3869);
nand U5026 (N_5026,N_3396,N_3174);
xnor U5027 (N_5027,N_4391,N_3555);
or U5028 (N_5028,N_4315,N_3483);
nand U5029 (N_5029,N_3778,N_3518);
or U5030 (N_5030,N_3696,N_3959);
or U5031 (N_5031,N_3768,N_4041);
and U5032 (N_5032,N_3999,N_3443);
nand U5033 (N_5033,N_4008,N_3494);
and U5034 (N_5034,N_4010,N_3472);
nor U5035 (N_5035,N_3001,N_4137);
xor U5036 (N_5036,N_3502,N_4098);
or U5037 (N_5037,N_3848,N_4464);
or U5038 (N_5038,N_3628,N_3157);
or U5039 (N_5039,N_4388,N_3381);
xnor U5040 (N_5040,N_3007,N_3786);
and U5041 (N_5041,N_3339,N_4267);
or U5042 (N_5042,N_3642,N_3441);
and U5043 (N_5043,N_3375,N_4220);
nor U5044 (N_5044,N_3403,N_4440);
nand U5045 (N_5045,N_4224,N_3233);
and U5046 (N_5046,N_3590,N_3335);
or U5047 (N_5047,N_4290,N_3309);
nand U5048 (N_5048,N_4425,N_3922);
or U5049 (N_5049,N_4019,N_4197);
and U5050 (N_5050,N_3251,N_3763);
or U5051 (N_5051,N_3355,N_3215);
nand U5052 (N_5052,N_3859,N_4304);
xor U5053 (N_5053,N_3773,N_4489);
xor U5054 (N_5054,N_4329,N_3663);
and U5055 (N_5055,N_3684,N_3199);
xnor U5056 (N_5056,N_3896,N_3787);
nand U5057 (N_5057,N_3568,N_3564);
or U5058 (N_5058,N_3780,N_3127);
xor U5059 (N_5059,N_3252,N_3316);
xnor U5060 (N_5060,N_4215,N_4077);
and U5061 (N_5061,N_3906,N_3662);
nand U5062 (N_5062,N_4262,N_3083);
or U5063 (N_5063,N_3447,N_4117);
nand U5064 (N_5064,N_4431,N_3096);
and U5065 (N_5065,N_4177,N_3499);
and U5066 (N_5066,N_3770,N_3419);
nand U5067 (N_5067,N_3724,N_3979);
and U5068 (N_5068,N_4484,N_4113);
nand U5069 (N_5069,N_3892,N_4351);
nand U5070 (N_5070,N_4250,N_3140);
or U5071 (N_5071,N_3495,N_4271);
nor U5072 (N_5072,N_3565,N_4206);
nand U5073 (N_5073,N_3330,N_3671);
xnor U5074 (N_5074,N_3218,N_3004);
or U5075 (N_5075,N_3609,N_4075);
and U5076 (N_5076,N_3936,N_3429);
or U5077 (N_5077,N_3895,N_4226);
and U5078 (N_5078,N_3286,N_4371);
xor U5079 (N_5079,N_4127,N_3818);
nand U5080 (N_5080,N_3223,N_4439);
and U5081 (N_5081,N_3196,N_3180);
or U5082 (N_5082,N_3299,N_3137);
nand U5083 (N_5083,N_4336,N_4497);
nor U5084 (N_5084,N_3006,N_3155);
and U5085 (N_5085,N_4138,N_4299);
xnor U5086 (N_5086,N_3994,N_3053);
nand U5087 (N_5087,N_3658,N_3592);
and U5088 (N_5088,N_3256,N_3992);
or U5089 (N_5089,N_3681,N_3430);
nor U5090 (N_5090,N_3120,N_4005);
nand U5091 (N_5091,N_3266,N_3217);
nor U5092 (N_5092,N_3136,N_4269);
and U5093 (N_5093,N_3241,N_3123);
xnor U5094 (N_5094,N_3201,N_4016);
nand U5095 (N_5095,N_4181,N_4046);
or U5096 (N_5096,N_4106,N_3623);
xnor U5097 (N_5097,N_3620,N_3362);
xnor U5098 (N_5098,N_3949,N_4457);
nand U5099 (N_5099,N_4023,N_3059);
nor U5100 (N_5100,N_4347,N_4309);
and U5101 (N_5101,N_4097,N_3560);
and U5102 (N_5102,N_4073,N_4437);
xnor U5103 (N_5103,N_3987,N_3857);
and U5104 (N_5104,N_3645,N_3789);
nor U5105 (N_5105,N_4325,N_4186);
xor U5106 (N_5106,N_4321,N_3647);
nand U5107 (N_5107,N_3745,N_3052);
xor U5108 (N_5108,N_3578,N_3278);
nand U5109 (N_5109,N_3528,N_4066);
or U5110 (N_5110,N_3713,N_3913);
nand U5111 (N_5111,N_3418,N_4221);
nor U5112 (N_5112,N_3306,N_4152);
and U5113 (N_5113,N_3236,N_4308);
and U5114 (N_5114,N_4368,N_3064);
nor U5115 (N_5115,N_3214,N_3129);
and U5116 (N_5116,N_3189,N_3962);
nand U5117 (N_5117,N_4458,N_3974);
or U5118 (N_5118,N_3952,N_3255);
xor U5119 (N_5119,N_3019,N_3506);
nand U5120 (N_5120,N_4476,N_3917);
or U5121 (N_5121,N_3603,N_4449);
and U5122 (N_5122,N_4384,N_4126);
xnor U5123 (N_5123,N_3722,N_3015);
nor U5124 (N_5124,N_4167,N_3467);
nand U5125 (N_5125,N_3160,N_3112);
nor U5126 (N_5126,N_4301,N_3091);
and U5127 (N_5127,N_3077,N_3205);
nand U5128 (N_5128,N_3184,N_4374);
xnor U5129 (N_5129,N_4060,N_3302);
nor U5130 (N_5130,N_3197,N_4086);
or U5131 (N_5131,N_3556,N_3188);
and U5132 (N_5132,N_3920,N_3183);
xnor U5133 (N_5133,N_4366,N_3888);
nand U5134 (N_5134,N_4094,N_3386);
nand U5135 (N_5135,N_4022,N_4180);
or U5136 (N_5136,N_3751,N_4151);
and U5137 (N_5137,N_3040,N_4459);
or U5138 (N_5138,N_4286,N_3393);
or U5139 (N_5139,N_3046,N_4210);
xnor U5140 (N_5140,N_3611,N_3023);
xnor U5141 (N_5141,N_3925,N_3650);
nand U5142 (N_5142,N_3041,N_3391);
nand U5143 (N_5143,N_3228,N_3782);
and U5144 (N_5144,N_3762,N_4211);
nand U5145 (N_5145,N_4355,N_3887);
and U5146 (N_5146,N_3943,N_3536);
and U5147 (N_5147,N_3225,N_3835);
and U5148 (N_5148,N_4142,N_3596);
nor U5149 (N_5149,N_4410,N_4463);
nor U5150 (N_5150,N_4120,N_4483);
or U5151 (N_5151,N_4051,N_4193);
nand U5152 (N_5152,N_3954,N_3348);
xnor U5153 (N_5153,N_3301,N_3520);
xor U5154 (N_5154,N_4198,N_3747);
xnor U5155 (N_5155,N_3054,N_3121);
nor U5156 (N_5156,N_3625,N_3292);
and U5157 (N_5157,N_3382,N_3097);
nand U5158 (N_5158,N_3158,N_4488);
or U5159 (N_5159,N_3678,N_4163);
and U5160 (N_5160,N_3248,N_4499);
xnor U5161 (N_5161,N_4401,N_4189);
nor U5162 (N_5162,N_4328,N_4415);
xnor U5163 (N_5163,N_4252,N_3799);
or U5164 (N_5164,N_4318,N_3889);
or U5165 (N_5165,N_3186,N_4136);
and U5166 (N_5166,N_4099,N_3547);
nor U5167 (N_5167,N_4375,N_3510);
nand U5168 (N_5168,N_3108,N_3972);
nand U5169 (N_5169,N_3866,N_3817);
xor U5170 (N_5170,N_4495,N_3020);
xnor U5171 (N_5171,N_3667,N_4398);
xor U5172 (N_5172,N_4213,N_4337);
nor U5173 (N_5173,N_3613,N_4082);
or U5174 (N_5174,N_3562,N_3173);
nand U5175 (N_5175,N_4326,N_3811);
nor U5176 (N_5176,N_3281,N_3211);
xnor U5177 (N_5177,N_3607,N_3990);
nand U5178 (N_5178,N_3114,N_4322);
nand U5179 (N_5179,N_4445,N_3043);
or U5180 (N_5180,N_3635,N_3690);
or U5181 (N_5181,N_3224,N_3692);
and U5182 (N_5182,N_3569,N_3220);
or U5183 (N_5183,N_3826,N_3293);
nand U5184 (N_5184,N_4474,N_3126);
and U5185 (N_5185,N_3454,N_4429);
and U5186 (N_5186,N_4012,N_3254);
xnor U5187 (N_5187,N_3575,N_4065);
or U5188 (N_5188,N_3709,N_4006);
nor U5189 (N_5189,N_3824,N_3312);
nor U5190 (N_5190,N_3263,N_4036);
and U5191 (N_5191,N_4418,N_3213);
and U5192 (N_5192,N_3487,N_3156);
nor U5193 (N_5193,N_4067,N_4472);
xor U5194 (N_5194,N_3567,N_4080);
or U5195 (N_5195,N_3626,N_4031);
xnor U5196 (N_5196,N_3234,N_3627);
xor U5197 (N_5197,N_4043,N_4150);
nand U5198 (N_5198,N_3247,N_3507);
xor U5199 (N_5199,N_3193,N_4393);
xor U5200 (N_5200,N_3622,N_3832);
xor U5201 (N_5201,N_4128,N_3961);
and U5202 (N_5202,N_3523,N_4486);
and U5203 (N_5203,N_3141,N_3784);
nor U5204 (N_5204,N_3460,N_3894);
nand U5205 (N_5205,N_4357,N_3349);
nor U5206 (N_5206,N_3588,N_3168);
xnor U5207 (N_5207,N_4430,N_4414);
or U5208 (N_5208,N_3549,N_3277);
nand U5209 (N_5209,N_3475,N_3377);
and U5210 (N_5210,N_3893,N_3334);
nand U5211 (N_5211,N_4231,N_3261);
nand U5212 (N_5212,N_3720,N_3912);
xnor U5213 (N_5213,N_3637,N_4052);
or U5214 (N_5214,N_3249,N_3806);
and U5215 (N_5215,N_4092,N_3561);
and U5216 (N_5216,N_3404,N_3028);
or U5217 (N_5217,N_4485,N_4432);
nor U5218 (N_5218,N_3985,N_4229);
and U5219 (N_5219,N_3148,N_3433);
or U5220 (N_5220,N_4148,N_3074);
or U5221 (N_5221,N_3723,N_4090);
nor U5222 (N_5222,N_3501,N_3597);
and U5223 (N_5223,N_3553,N_3514);
xnor U5224 (N_5224,N_3154,N_3932);
nand U5225 (N_5225,N_3717,N_3260);
and U5226 (N_5226,N_4339,N_4013);
or U5227 (N_5227,N_3831,N_3387);
xor U5228 (N_5228,N_3493,N_3503);
and U5229 (N_5229,N_4434,N_4381);
xor U5230 (N_5230,N_3973,N_4327);
or U5231 (N_5231,N_3276,N_4096);
nand U5232 (N_5232,N_4443,N_4176);
nor U5233 (N_5233,N_3376,N_4248);
nand U5234 (N_5234,N_4232,N_3284);
and U5235 (N_5235,N_4405,N_3814);
or U5236 (N_5236,N_3219,N_3253);
xor U5237 (N_5237,N_3505,N_3307);
nor U5238 (N_5238,N_3750,N_4481);
or U5239 (N_5239,N_4140,N_3966);
or U5240 (N_5240,N_3643,N_4178);
nor U5241 (N_5241,N_3516,N_3863);
nor U5242 (N_5242,N_3907,N_3736);
and U5243 (N_5243,N_3829,N_4102);
nor U5244 (N_5244,N_3439,N_3411);
nor U5245 (N_5245,N_3389,N_3942);
nor U5246 (N_5246,N_3267,N_4465);
or U5247 (N_5247,N_3664,N_4402);
and U5248 (N_5248,N_3098,N_3970);
or U5249 (N_5249,N_4417,N_4209);
xor U5250 (N_5250,N_3621,N_3591);
and U5251 (N_5251,N_3981,N_3701);
xnor U5252 (N_5252,N_3635,N_4103);
xor U5253 (N_5253,N_3699,N_4049);
nand U5254 (N_5254,N_3773,N_3674);
and U5255 (N_5255,N_3199,N_3884);
and U5256 (N_5256,N_3691,N_3785);
and U5257 (N_5257,N_3693,N_3629);
xor U5258 (N_5258,N_3335,N_3619);
nand U5259 (N_5259,N_4304,N_3723);
or U5260 (N_5260,N_4204,N_3151);
nand U5261 (N_5261,N_3940,N_3899);
and U5262 (N_5262,N_4137,N_3097);
nor U5263 (N_5263,N_3653,N_4386);
or U5264 (N_5264,N_4229,N_4148);
or U5265 (N_5265,N_3676,N_3082);
nand U5266 (N_5266,N_3064,N_4383);
nand U5267 (N_5267,N_3882,N_3177);
nand U5268 (N_5268,N_4343,N_3215);
xnor U5269 (N_5269,N_3780,N_3841);
nor U5270 (N_5270,N_3054,N_4477);
and U5271 (N_5271,N_3362,N_4157);
and U5272 (N_5272,N_3643,N_4189);
nand U5273 (N_5273,N_4049,N_3054);
or U5274 (N_5274,N_3357,N_3013);
and U5275 (N_5275,N_4203,N_3911);
nor U5276 (N_5276,N_3965,N_4298);
nand U5277 (N_5277,N_3937,N_3004);
or U5278 (N_5278,N_3947,N_3977);
and U5279 (N_5279,N_3608,N_4463);
nor U5280 (N_5280,N_3924,N_3005);
or U5281 (N_5281,N_4434,N_3114);
nand U5282 (N_5282,N_3749,N_3178);
xnor U5283 (N_5283,N_3493,N_4089);
xnor U5284 (N_5284,N_4413,N_3687);
nor U5285 (N_5285,N_3114,N_3368);
and U5286 (N_5286,N_3403,N_3357);
nor U5287 (N_5287,N_3516,N_3939);
or U5288 (N_5288,N_3135,N_3976);
and U5289 (N_5289,N_4237,N_4038);
nor U5290 (N_5290,N_3711,N_3241);
nor U5291 (N_5291,N_3432,N_3727);
xor U5292 (N_5292,N_3433,N_3210);
nand U5293 (N_5293,N_3786,N_4391);
nand U5294 (N_5294,N_3371,N_3566);
or U5295 (N_5295,N_3505,N_4273);
nor U5296 (N_5296,N_3866,N_3434);
xnor U5297 (N_5297,N_4311,N_4297);
and U5298 (N_5298,N_3636,N_3740);
xor U5299 (N_5299,N_3292,N_4351);
or U5300 (N_5300,N_3854,N_3747);
and U5301 (N_5301,N_3314,N_4348);
or U5302 (N_5302,N_3187,N_3662);
or U5303 (N_5303,N_3695,N_3634);
nor U5304 (N_5304,N_4303,N_3387);
nor U5305 (N_5305,N_3503,N_4455);
nor U5306 (N_5306,N_3659,N_4462);
and U5307 (N_5307,N_4086,N_4036);
or U5308 (N_5308,N_3203,N_3529);
xor U5309 (N_5309,N_3346,N_3617);
nor U5310 (N_5310,N_4074,N_3920);
or U5311 (N_5311,N_4364,N_3452);
xor U5312 (N_5312,N_3804,N_4164);
xor U5313 (N_5313,N_4238,N_3963);
xor U5314 (N_5314,N_3884,N_3650);
and U5315 (N_5315,N_4496,N_3661);
xnor U5316 (N_5316,N_3297,N_4164);
nand U5317 (N_5317,N_3794,N_4118);
or U5318 (N_5318,N_3516,N_3462);
and U5319 (N_5319,N_4462,N_3764);
nor U5320 (N_5320,N_3517,N_3785);
nor U5321 (N_5321,N_3560,N_4098);
xnor U5322 (N_5322,N_3669,N_4472);
xor U5323 (N_5323,N_3101,N_4124);
xnor U5324 (N_5324,N_4318,N_3601);
nand U5325 (N_5325,N_3605,N_4115);
xnor U5326 (N_5326,N_3899,N_3523);
and U5327 (N_5327,N_4080,N_3771);
or U5328 (N_5328,N_3217,N_3052);
and U5329 (N_5329,N_3333,N_3911);
nor U5330 (N_5330,N_3287,N_3176);
and U5331 (N_5331,N_3921,N_3810);
nor U5332 (N_5332,N_4429,N_3407);
nor U5333 (N_5333,N_4087,N_3335);
and U5334 (N_5334,N_3355,N_3118);
and U5335 (N_5335,N_3713,N_4231);
and U5336 (N_5336,N_4142,N_3029);
and U5337 (N_5337,N_3786,N_4195);
xor U5338 (N_5338,N_4125,N_3420);
nand U5339 (N_5339,N_3108,N_4000);
nand U5340 (N_5340,N_3676,N_3617);
nand U5341 (N_5341,N_4331,N_3338);
nor U5342 (N_5342,N_3925,N_3614);
nor U5343 (N_5343,N_3374,N_4207);
or U5344 (N_5344,N_4283,N_3458);
and U5345 (N_5345,N_3499,N_4020);
xnor U5346 (N_5346,N_3745,N_3713);
xor U5347 (N_5347,N_3850,N_3687);
xor U5348 (N_5348,N_3058,N_3768);
xnor U5349 (N_5349,N_3976,N_3416);
xnor U5350 (N_5350,N_3021,N_3230);
nand U5351 (N_5351,N_4039,N_4098);
and U5352 (N_5352,N_3663,N_4105);
and U5353 (N_5353,N_4395,N_3046);
xor U5354 (N_5354,N_3432,N_3005);
and U5355 (N_5355,N_3874,N_3651);
xor U5356 (N_5356,N_3646,N_3012);
xnor U5357 (N_5357,N_3764,N_3275);
or U5358 (N_5358,N_3640,N_3680);
xor U5359 (N_5359,N_3097,N_3698);
and U5360 (N_5360,N_4104,N_4323);
and U5361 (N_5361,N_3696,N_3040);
or U5362 (N_5362,N_4402,N_3398);
nand U5363 (N_5363,N_4310,N_3158);
and U5364 (N_5364,N_3244,N_3435);
and U5365 (N_5365,N_3219,N_4279);
nand U5366 (N_5366,N_3054,N_3194);
or U5367 (N_5367,N_3991,N_4387);
nand U5368 (N_5368,N_4037,N_4391);
nand U5369 (N_5369,N_3823,N_4272);
xor U5370 (N_5370,N_4455,N_4128);
or U5371 (N_5371,N_4029,N_3238);
or U5372 (N_5372,N_4486,N_4253);
nand U5373 (N_5373,N_4377,N_4092);
nand U5374 (N_5374,N_3578,N_3616);
nand U5375 (N_5375,N_4063,N_4044);
nand U5376 (N_5376,N_4210,N_3900);
xor U5377 (N_5377,N_3441,N_3186);
nand U5378 (N_5378,N_4090,N_3874);
or U5379 (N_5379,N_4089,N_3523);
and U5380 (N_5380,N_3073,N_3399);
or U5381 (N_5381,N_3328,N_3098);
or U5382 (N_5382,N_3154,N_3493);
xnor U5383 (N_5383,N_3507,N_3039);
or U5384 (N_5384,N_4139,N_3856);
xor U5385 (N_5385,N_4060,N_3143);
and U5386 (N_5386,N_3973,N_3110);
and U5387 (N_5387,N_3288,N_3919);
or U5388 (N_5388,N_3416,N_3454);
xor U5389 (N_5389,N_4071,N_3630);
or U5390 (N_5390,N_3995,N_3352);
xnor U5391 (N_5391,N_4130,N_3588);
nand U5392 (N_5392,N_3897,N_3148);
and U5393 (N_5393,N_3456,N_3486);
and U5394 (N_5394,N_3484,N_4072);
and U5395 (N_5395,N_3068,N_3639);
and U5396 (N_5396,N_3542,N_4017);
xnor U5397 (N_5397,N_4084,N_3219);
or U5398 (N_5398,N_3208,N_3775);
nor U5399 (N_5399,N_3038,N_3427);
nand U5400 (N_5400,N_4339,N_3530);
nor U5401 (N_5401,N_3962,N_4228);
and U5402 (N_5402,N_4472,N_4031);
nor U5403 (N_5403,N_3604,N_4488);
nor U5404 (N_5404,N_3922,N_4036);
xor U5405 (N_5405,N_4163,N_3823);
or U5406 (N_5406,N_3036,N_4104);
and U5407 (N_5407,N_3002,N_3451);
and U5408 (N_5408,N_4226,N_3940);
or U5409 (N_5409,N_4326,N_4206);
xnor U5410 (N_5410,N_4209,N_3053);
or U5411 (N_5411,N_3891,N_3180);
nor U5412 (N_5412,N_4063,N_3524);
and U5413 (N_5413,N_4124,N_4317);
xor U5414 (N_5414,N_3297,N_3313);
xnor U5415 (N_5415,N_3812,N_3090);
or U5416 (N_5416,N_3213,N_4065);
xor U5417 (N_5417,N_3265,N_3971);
nand U5418 (N_5418,N_3477,N_3667);
and U5419 (N_5419,N_3885,N_4059);
and U5420 (N_5420,N_3932,N_4070);
or U5421 (N_5421,N_3758,N_3004);
or U5422 (N_5422,N_3284,N_3591);
nor U5423 (N_5423,N_4337,N_3530);
or U5424 (N_5424,N_3716,N_4103);
or U5425 (N_5425,N_3104,N_4043);
nand U5426 (N_5426,N_3032,N_3991);
xnor U5427 (N_5427,N_3402,N_3266);
xor U5428 (N_5428,N_3096,N_3779);
xor U5429 (N_5429,N_3120,N_3097);
and U5430 (N_5430,N_3599,N_4370);
or U5431 (N_5431,N_3176,N_4081);
or U5432 (N_5432,N_3295,N_3449);
nor U5433 (N_5433,N_4196,N_3851);
and U5434 (N_5434,N_3417,N_3118);
nand U5435 (N_5435,N_3374,N_3772);
nor U5436 (N_5436,N_4382,N_3504);
nor U5437 (N_5437,N_4381,N_3112);
xnor U5438 (N_5438,N_3449,N_4126);
nand U5439 (N_5439,N_3016,N_4346);
nand U5440 (N_5440,N_3651,N_3170);
xnor U5441 (N_5441,N_3000,N_3407);
or U5442 (N_5442,N_3676,N_4140);
nand U5443 (N_5443,N_3495,N_3945);
xor U5444 (N_5444,N_3198,N_4372);
xor U5445 (N_5445,N_3070,N_3216);
nor U5446 (N_5446,N_4121,N_3464);
or U5447 (N_5447,N_4087,N_3215);
or U5448 (N_5448,N_4156,N_4106);
xnor U5449 (N_5449,N_3235,N_3659);
nor U5450 (N_5450,N_3699,N_3455);
xnor U5451 (N_5451,N_4338,N_4418);
nand U5452 (N_5452,N_3137,N_4118);
or U5453 (N_5453,N_4415,N_4098);
nand U5454 (N_5454,N_3023,N_3985);
nand U5455 (N_5455,N_3391,N_3214);
nor U5456 (N_5456,N_3360,N_4036);
or U5457 (N_5457,N_4054,N_3091);
and U5458 (N_5458,N_3360,N_3383);
nor U5459 (N_5459,N_4470,N_3666);
nor U5460 (N_5460,N_3806,N_3412);
nor U5461 (N_5461,N_3707,N_3757);
or U5462 (N_5462,N_3033,N_3766);
and U5463 (N_5463,N_4397,N_4262);
xnor U5464 (N_5464,N_3300,N_4371);
nand U5465 (N_5465,N_3734,N_4488);
and U5466 (N_5466,N_3708,N_3381);
and U5467 (N_5467,N_3618,N_3208);
nor U5468 (N_5468,N_3181,N_4189);
or U5469 (N_5469,N_3716,N_4425);
nor U5470 (N_5470,N_3780,N_4179);
nor U5471 (N_5471,N_3646,N_3972);
nor U5472 (N_5472,N_3684,N_3763);
or U5473 (N_5473,N_4410,N_3960);
nand U5474 (N_5474,N_3924,N_3795);
nand U5475 (N_5475,N_3668,N_4121);
and U5476 (N_5476,N_3054,N_3399);
and U5477 (N_5477,N_3159,N_4402);
xor U5478 (N_5478,N_3605,N_3649);
or U5479 (N_5479,N_3542,N_3387);
xor U5480 (N_5480,N_3491,N_3777);
xor U5481 (N_5481,N_3872,N_3566);
or U5482 (N_5482,N_3067,N_4460);
nor U5483 (N_5483,N_3298,N_3856);
nor U5484 (N_5484,N_3158,N_3231);
nand U5485 (N_5485,N_4447,N_4250);
and U5486 (N_5486,N_3119,N_3653);
xnor U5487 (N_5487,N_4380,N_3917);
nor U5488 (N_5488,N_3315,N_3248);
and U5489 (N_5489,N_3239,N_3199);
xnor U5490 (N_5490,N_3421,N_3725);
and U5491 (N_5491,N_3551,N_3182);
xnor U5492 (N_5492,N_3901,N_3263);
and U5493 (N_5493,N_4395,N_3079);
nor U5494 (N_5494,N_3427,N_4384);
nand U5495 (N_5495,N_3892,N_3981);
nand U5496 (N_5496,N_4157,N_3254);
and U5497 (N_5497,N_4495,N_4403);
xor U5498 (N_5498,N_3285,N_3917);
and U5499 (N_5499,N_4027,N_4245);
and U5500 (N_5500,N_3341,N_3402);
nand U5501 (N_5501,N_3205,N_4155);
and U5502 (N_5502,N_3136,N_3728);
xor U5503 (N_5503,N_3893,N_4233);
nand U5504 (N_5504,N_4453,N_3539);
or U5505 (N_5505,N_3976,N_4263);
or U5506 (N_5506,N_4356,N_3558);
xor U5507 (N_5507,N_4356,N_4011);
nand U5508 (N_5508,N_3229,N_3134);
nor U5509 (N_5509,N_3875,N_4417);
xor U5510 (N_5510,N_3029,N_3431);
xnor U5511 (N_5511,N_4037,N_4342);
nand U5512 (N_5512,N_4190,N_3728);
nor U5513 (N_5513,N_4152,N_3342);
and U5514 (N_5514,N_3957,N_3765);
nand U5515 (N_5515,N_3199,N_4130);
nand U5516 (N_5516,N_3386,N_3546);
nor U5517 (N_5517,N_4343,N_3204);
nor U5518 (N_5518,N_3607,N_3943);
nor U5519 (N_5519,N_3482,N_3400);
xor U5520 (N_5520,N_3857,N_3929);
nand U5521 (N_5521,N_4443,N_4183);
or U5522 (N_5522,N_3275,N_3862);
xor U5523 (N_5523,N_3187,N_3688);
and U5524 (N_5524,N_3617,N_4370);
xnor U5525 (N_5525,N_3538,N_4347);
nor U5526 (N_5526,N_3080,N_3314);
or U5527 (N_5527,N_3064,N_3100);
nor U5528 (N_5528,N_3444,N_4038);
xnor U5529 (N_5529,N_3525,N_3416);
xor U5530 (N_5530,N_4246,N_4034);
nand U5531 (N_5531,N_3068,N_4119);
and U5532 (N_5532,N_3563,N_3894);
nor U5533 (N_5533,N_4396,N_4389);
xor U5534 (N_5534,N_3001,N_3490);
nand U5535 (N_5535,N_3090,N_4169);
xor U5536 (N_5536,N_3814,N_4474);
or U5537 (N_5537,N_3985,N_3853);
nand U5538 (N_5538,N_3788,N_4172);
xnor U5539 (N_5539,N_3230,N_3662);
or U5540 (N_5540,N_3454,N_3331);
or U5541 (N_5541,N_3727,N_3699);
nand U5542 (N_5542,N_3062,N_4014);
xor U5543 (N_5543,N_3093,N_3205);
and U5544 (N_5544,N_3378,N_4473);
xnor U5545 (N_5545,N_4391,N_3604);
or U5546 (N_5546,N_4041,N_3746);
or U5547 (N_5547,N_3613,N_4006);
and U5548 (N_5548,N_3157,N_4161);
or U5549 (N_5549,N_3076,N_4476);
and U5550 (N_5550,N_3368,N_3987);
or U5551 (N_5551,N_3924,N_3464);
or U5552 (N_5552,N_4187,N_4179);
xnor U5553 (N_5553,N_3049,N_4457);
nor U5554 (N_5554,N_4286,N_3280);
or U5555 (N_5555,N_3691,N_3218);
or U5556 (N_5556,N_3763,N_4460);
xor U5557 (N_5557,N_3267,N_3362);
or U5558 (N_5558,N_4342,N_3590);
and U5559 (N_5559,N_3539,N_3493);
xor U5560 (N_5560,N_3880,N_4335);
nor U5561 (N_5561,N_3586,N_3663);
nor U5562 (N_5562,N_3293,N_3931);
nor U5563 (N_5563,N_3033,N_3773);
nand U5564 (N_5564,N_4018,N_3404);
xor U5565 (N_5565,N_3728,N_3768);
and U5566 (N_5566,N_3304,N_3264);
nand U5567 (N_5567,N_3800,N_3749);
and U5568 (N_5568,N_3596,N_3210);
nor U5569 (N_5569,N_4073,N_3821);
xor U5570 (N_5570,N_3366,N_4038);
nand U5571 (N_5571,N_3822,N_4315);
nor U5572 (N_5572,N_3803,N_4038);
nand U5573 (N_5573,N_4116,N_3095);
nand U5574 (N_5574,N_3037,N_4242);
and U5575 (N_5575,N_4178,N_3222);
xor U5576 (N_5576,N_3855,N_3585);
or U5577 (N_5577,N_4282,N_3082);
nor U5578 (N_5578,N_4203,N_3860);
nor U5579 (N_5579,N_3976,N_3964);
or U5580 (N_5580,N_3631,N_3636);
and U5581 (N_5581,N_3691,N_3364);
or U5582 (N_5582,N_3150,N_3384);
xor U5583 (N_5583,N_3395,N_4323);
or U5584 (N_5584,N_4045,N_3949);
nand U5585 (N_5585,N_3988,N_3661);
and U5586 (N_5586,N_4391,N_4232);
or U5587 (N_5587,N_3082,N_4379);
nand U5588 (N_5588,N_4350,N_3955);
nor U5589 (N_5589,N_4220,N_3650);
and U5590 (N_5590,N_4183,N_4426);
or U5591 (N_5591,N_4337,N_3223);
nand U5592 (N_5592,N_3052,N_3766);
or U5593 (N_5593,N_4387,N_4432);
or U5594 (N_5594,N_3230,N_3242);
nor U5595 (N_5595,N_3111,N_3679);
or U5596 (N_5596,N_3848,N_3594);
nor U5597 (N_5597,N_3473,N_3846);
nand U5598 (N_5598,N_4279,N_4023);
and U5599 (N_5599,N_3480,N_3254);
nand U5600 (N_5600,N_4211,N_3700);
nand U5601 (N_5601,N_3903,N_3695);
or U5602 (N_5602,N_3419,N_4480);
nand U5603 (N_5603,N_3597,N_3799);
xor U5604 (N_5604,N_4026,N_4075);
nor U5605 (N_5605,N_4068,N_3661);
and U5606 (N_5606,N_3459,N_3101);
xor U5607 (N_5607,N_3518,N_3679);
nor U5608 (N_5608,N_4061,N_3771);
nor U5609 (N_5609,N_4412,N_3218);
nand U5610 (N_5610,N_3985,N_4046);
nor U5611 (N_5611,N_4489,N_3627);
xor U5612 (N_5612,N_4083,N_3610);
nor U5613 (N_5613,N_4149,N_4414);
nor U5614 (N_5614,N_4256,N_3795);
and U5615 (N_5615,N_4113,N_3718);
or U5616 (N_5616,N_4463,N_4050);
or U5617 (N_5617,N_3848,N_3800);
nor U5618 (N_5618,N_3445,N_4396);
and U5619 (N_5619,N_4212,N_3686);
nand U5620 (N_5620,N_3224,N_3219);
xnor U5621 (N_5621,N_4110,N_3248);
or U5622 (N_5622,N_3186,N_3636);
xor U5623 (N_5623,N_3555,N_4010);
nand U5624 (N_5624,N_3817,N_3706);
nor U5625 (N_5625,N_4306,N_3386);
or U5626 (N_5626,N_4185,N_4072);
nand U5627 (N_5627,N_4078,N_3485);
xor U5628 (N_5628,N_4063,N_3621);
nand U5629 (N_5629,N_3439,N_3076);
xnor U5630 (N_5630,N_3786,N_3794);
or U5631 (N_5631,N_4261,N_3582);
and U5632 (N_5632,N_3785,N_4190);
nor U5633 (N_5633,N_3682,N_3119);
nor U5634 (N_5634,N_3321,N_4088);
nor U5635 (N_5635,N_4106,N_4002);
xor U5636 (N_5636,N_3714,N_3168);
xor U5637 (N_5637,N_3111,N_3840);
xor U5638 (N_5638,N_3479,N_3812);
xor U5639 (N_5639,N_4416,N_4296);
nor U5640 (N_5640,N_3546,N_3316);
nor U5641 (N_5641,N_4126,N_3665);
nand U5642 (N_5642,N_4077,N_3220);
nor U5643 (N_5643,N_4277,N_4392);
nand U5644 (N_5644,N_4275,N_3328);
or U5645 (N_5645,N_3612,N_3852);
nand U5646 (N_5646,N_4223,N_3246);
and U5647 (N_5647,N_3389,N_4434);
xor U5648 (N_5648,N_4214,N_3986);
nor U5649 (N_5649,N_3942,N_3877);
nand U5650 (N_5650,N_4054,N_3756);
or U5651 (N_5651,N_3409,N_4244);
and U5652 (N_5652,N_3134,N_3034);
or U5653 (N_5653,N_3748,N_3383);
nand U5654 (N_5654,N_3228,N_4015);
and U5655 (N_5655,N_3108,N_3966);
nor U5656 (N_5656,N_3488,N_3705);
nor U5657 (N_5657,N_4397,N_3784);
xnor U5658 (N_5658,N_4173,N_4137);
nand U5659 (N_5659,N_4136,N_3060);
or U5660 (N_5660,N_3132,N_3491);
or U5661 (N_5661,N_3303,N_3422);
nor U5662 (N_5662,N_3272,N_3443);
and U5663 (N_5663,N_3854,N_4035);
or U5664 (N_5664,N_3771,N_3784);
nor U5665 (N_5665,N_3003,N_4252);
xor U5666 (N_5666,N_3326,N_3750);
and U5667 (N_5667,N_4370,N_3365);
nand U5668 (N_5668,N_3510,N_3751);
nor U5669 (N_5669,N_3526,N_4239);
nor U5670 (N_5670,N_3101,N_3881);
xor U5671 (N_5671,N_3096,N_3673);
nand U5672 (N_5672,N_4095,N_3869);
or U5673 (N_5673,N_3897,N_3291);
and U5674 (N_5674,N_4397,N_4371);
or U5675 (N_5675,N_3277,N_3846);
or U5676 (N_5676,N_3729,N_3804);
xnor U5677 (N_5677,N_4398,N_4115);
xor U5678 (N_5678,N_3589,N_3050);
nor U5679 (N_5679,N_3808,N_3934);
and U5680 (N_5680,N_3199,N_3071);
nor U5681 (N_5681,N_4372,N_3979);
xor U5682 (N_5682,N_3229,N_3890);
xnor U5683 (N_5683,N_3286,N_4394);
nor U5684 (N_5684,N_3793,N_4097);
and U5685 (N_5685,N_3772,N_3039);
nor U5686 (N_5686,N_4426,N_3328);
xnor U5687 (N_5687,N_4333,N_4293);
and U5688 (N_5688,N_4323,N_4306);
and U5689 (N_5689,N_3254,N_3763);
or U5690 (N_5690,N_3630,N_4429);
xnor U5691 (N_5691,N_3739,N_3290);
nor U5692 (N_5692,N_3742,N_4402);
and U5693 (N_5693,N_4239,N_3516);
nand U5694 (N_5694,N_4159,N_3914);
nand U5695 (N_5695,N_3716,N_3425);
or U5696 (N_5696,N_3589,N_3657);
nand U5697 (N_5697,N_3860,N_4249);
or U5698 (N_5698,N_3087,N_3324);
nand U5699 (N_5699,N_3534,N_3668);
or U5700 (N_5700,N_4227,N_3241);
nor U5701 (N_5701,N_3268,N_3675);
nor U5702 (N_5702,N_4068,N_3951);
and U5703 (N_5703,N_4201,N_3917);
and U5704 (N_5704,N_3283,N_4193);
nor U5705 (N_5705,N_4169,N_3249);
nor U5706 (N_5706,N_4285,N_4024);
xor U5707 (N_5707,N_4360,N_3895);
or U5708 (N_5708,N_3999,N_3979);
nand U5709 (N_5709,N_4196,N_3680);
nor U5710 (N_5710,N_3545,N_4382);
or U5711 (N_5711,N_3042,N_3670);
nor U5712 (N_5712,N_3236,N_3336);
nand U5713 (N_5713,N_3449,N_3531);
and U5714 (N_5714,N_3735,N_3434);
nor U5715 (N_5715,N_3623,N_4281);
and U5716 (N_5716,N_4375,N_3275);
and U5717 (N_5717,N_3229,N_3960);
or U5718 (N_5718,N_3117,N_3718);
nand U5719 (N_5719,N_3018,N_3458);
and U5720 (N_5720,N_3610,N_3883);
xor U5721 (N_5721,N_3516,N_3637);
or U5722 (N_5722,N_4043,N_3466);
nand U5723 (N_5723,N_4369,N_3825);
and U5724 (N_5724,N_3998,N_3493);
and U5725 (N_5725,N_3395,N_4210);
nor U5726 (N_5726,N_4480,N_3327);
xor U5727 (N_5727,N_4190,N_4270);
or U5728 (N_5728,N_4416,N_3468);
nor U5729 (N_5729,N_3771,N_4043);
nand U5730 (N_5730,N_3475,N_4372);
or U5731 (N_5731,N_3973,N_3101);
nand U5732 (N_5732,N_3300,N_3916);
nor U5733 (N_5733,N_3487,N_4267);
xor U5734 (N_5734,N_4180,N_3179);
nor U5735 (N_5735,N_4157,N_4290);
nor U5736 (N_5736,N_4030,N_4136);
nand U5737 (N_5737,N_4401,N_3129);
nor U5738 (N_5738,N_3123,N_3331);
and U5739 (N_5739,N_4323,N_4314);
or U5740 (N_5740,N_4268,N_3145);
nand U5741 (N_5741,N_4104,N_3615);
and U5742 (N_5742,N_4366,N_4074);
nand U5743 (N_5743,N_3158,N_3365);
and U5744 (N_5744,N_4379,N_4052);
and U5745 (N_5745,N_3345,N_3801);
and U5746 (N_5746,N_3001,N_3062);
nor U5747 (N_5747,N_3590,N_3390);
and U5748 (N_5748,N_3426,N_3705);
nor U5749 (N_5749,N_3918,N_3330);
xor U5750 (N_5750,N_3055,N_4198);
xnor U5751 (N_5751,N_3023,N_3330);
xor U5752 (N_5752,N_4256,N_3832);
xnor U5753 (N_5753,N_4402,N_3994);
xnor U5754 (N_5754,N_3350,N_3894);
nor U5755 (N_5755,N_4353,N_3764);
nor U5756 (N_5756,N_4440,N_3932);
nor U5757 (N_5757,N_3720,N_3350);
or U5758 (N_5758,N_4204,N_3609);
and U5759 (N_5759,N_4135,N_3803);
xnor U5760 (N_5760,N_4106,N_4425);
nor U5761 (N_5761,N_3221,N_4029);
nand U5762 (N_5762,N_3859,N_3919);
or U5763 (N_5763,N_3817,N_3257);
and U5764 (N_5764,N_3309,N_4151);
nand U5765 (N_5765,N_3443,N_4452);
nand U5766 (N_5766,N_3605,N_4375);
nand U5767 (N_5767,N_3684,N_3020);
nor U5768 (N_5768,N_4324,N_3085);
nor U5769 (N_5769,N_3930,N_4426);
or U5770 (N_5770,N_3731,N_4123);
and U5771 (N_5771,N_3206,N_3029);
nor U5772 (N_5772,N_3644,N_3908);
nor U5773 (N_5773,N_3439,N_4044);
xor U5774 (N_5774,N_4274,N_3817);
nor U5775 (N_5775,N_3638,N_3670);
or U5776 (N_5776,N_3229,N_3853);
xor U5777 (N_5777,N_3725,N_3672);
and U5778 (N_5778,N_4488,N_3405);
and U5779 (N_5779,N_3435,N_3025);
xnor U5780 (N_5780,N_3204,N_3540);
xnor U5781 (N_5781,N_3501,N_3826);
nor U5782 (N_5782,N_3520,N_3653);
or U5783 (N_5783,N_4334,N_3254);
and U5784 (N_5784,N_3251,N_4418);
nand U5785 (N_5785,N_4034,N_3683);
nand U5786 (N_5786,N_4393,N_3772);
nand U5787 (N_5787,N_4104,N_3042);
xnor U5788 (N_5788,N_3706,N_4184);
nor U5789 (N_5789,N_4257,N_4435);
nor U5790 (N_5790,N_3632,N_3292);
or U5791 (N_5791,N_3284,N_3512);
and U5792 (N_5792,N_3209,N_3014);
and U5793 (N_5793,N_4297,N_3841);
and U5794 (N_5794,N_4452,N_3930);
and U5795 (N_5795,N_4349,N_3352);
nand U5796 (N_5796,N_3313,N_3696);
nand U5797 (N_5797,N_4168,N_3791);
xnor U5798 (N_5798,N_3191,N_3749);
nor U5799 (N_5799,N_4230,N_3872);
xnor U5800 (N_5800,N_3027,N_3789);
xnor U5801 (N_5801,N_3223,N_3759);
and U5802 (N_5802,N_3330,N_3439);
nand U5803 (N_5803,N_3284,N_3899);
and U5804 (N_5804,N_4001,N_4297);
and U5805 (N_5805,N_3143,N_3351);
and U5806 (N_5806,N_3014,N_3344);
xor U5807 (N_5807,N_3909,N_3454);
nor U5808 (N_5808,N_4438,N_4310);
nor U5809 (N_5809,N_3219,N_3114);
and U5810 (N_5810,N_3970,N_3854);
nand U5811 (N_5811,N_4368,N_3762);
and U5812 (N_5812,N_3779,N_3835);
and U5813 (N_5813,N_4486,N_3752);
and U5814 (N_5814,N_3303,N_4288);
nand U5815 (N_5815,N_4172,N_3989);
or U5816 (N_5816,N_4304,N_3753);
or U5817 (N_5817,N_3141,N_3802);
or U5818 (N_5818,N_3427,N_4338);
xor U5819 (N_5819,N_3945,N_3337);
or U5820 (N_5820,N_4004,N_3719);
nor U5821 (N_5821,N_4018,N_4317);
xnor U5822 (N_5822,N_4437,N_4270);
nor U5823 (N_5823,N_3994,N_3057);
nor U5824 (N_5824,N_4325,N_3265);
nor U5825 (N_5825,N_3798,N_3515);
and U5826 (N_5826,N_3037,N_4413);
nand U5827 (N_5827,N_4226,N_3063);
xor U5828 (N_5828,N_3772,N_3607);
or U5829 (N_5829,N_3822,N_3573);
nand U5830 (N_5830,N_3139,N_4044);
or U5831 (N_5831,N_3523,N_3799);
and U5832 (N_5832,N_4102,N_3350);
nand U5833 (N_5833,N_4460,N_4111);
or U5834 (N_5834,N_3641,N_3243);
nor U5835 (N_5835,N_4045,N_3802);
and U5836 (N_5836,N_3440,N_3483);
nand U5837 (N_5837,N_4404,N_4307);
and U5838 (N_5838,N_4206,N_4225);
nand U5839 (N_5839,N_3183,N_4172);
or U5840 (N_5840,N_3582,N_3061);
or U5841 (N_5841,N_4023,N_3359);
xnor U5842 (N_5842,N_3434,N_4074);
xnor U5843 (N_5843,N_4445,N_3677);
nand U5844 (N_5844,N_4299,N_3748);
and U5845 (N_5845,N_3662,N_3579);
and U5846 (N_5846,N_4345,N_3098);
and U5847 (N_5847,N_4160,N_4010);
xor U5848 (N_5848,N_3640,N_4120);
and U5849 (N_5849,N_3517,N_3956);
nor U5850 (N_5850,N_4425,N_3645);
xor U5851 (N_5851,N_4234,N_3191);
and U5852 (N_5852,N_3269,N_3096);
xor U5853 (N_5853,N_3796,N_3768);
nand U5854 (N_5854,N_3066,N_4176);
nor U5855 (N_5855,N_3116,N_3028);
xnor U5856 (N_5856,N_4356,N_4139);
nor U5857 (N_5857,N_4103,N_3780);
nor U5858 (N_5858,N_3806,N_4238);
or U5859 (N_5859,N_3296,N_3376);
xnor U5860 (N_5860,N_4241,N_4170);
or U5861 (N_5861,N_3717,N_3786);
or U5862 (N_5862,N_3099,N_3407);
or U5863 (N_5863,N_4104,N_4439);
xor U5864 (N_5864,N_4054,N_3083);
and U5865 (N_5865,N_4164,N_4206);
or U5866 (N_5866,N_3098,N_3963);
nand U5867 (N_5867,N_3327,N_4137);
nand U5868 (N_5868,N_4369,N_3071);
xnor U5869 (N_5869,N_3755,N_3877);
and U5870 (N_5870,N_3681,N_3171);
and U5871 (N_5871,N_3066,N_4181);
xnor U5872 (N_5872,N_3692,N_4100);
xor U5873 (N_5873,N_4216,N_3016);
xnor U5874 (N_5874,N_4224,N_4461);
xor U5875 (N_5875,N_3308,N_3427);
xor U5876 (N_5876,N_3816,N_4396);
or U5877 (N_5877,N_3651,N_3790);
or U5878 (N_5878,N_4386,N_4158);
nand U5879 (N_5879,N_3847,N_3834);
xor U5880 (N_5880,N_3393,N_4007);
nand U5881 (N_5881,N_4137,N_3315);
or U5882 (N_5882,N_3021,N_3125);
and U5883 (N_5883,N_3797,N_3861);
xnor U5884 (N_5884,N_3329,N_4123);
nand U5885 (N_5885,N_4263,N_3606);
or U5886 (N_5886,N_3184,N_3017);
nand U5887 (N_5887,N_4404,N_3762);
nand U5888 (N_5888,N_3728,N_3817);
and U5889 (N_5889,N_4170,N_3310);
or U5890 (N_5890,N_4013,N_4430);
nand U5891 (N_5891,N_3071,N_3040);
or U5892 (N_5892,N_4284,N_3410);
or U5893 (N_5893,N_3090,N_3241);
nor U5894 (N_5894,N_3802,N_4397);
and U5895 (N_5895,N_4316,N_4351);
xnor U5896 (N_5896,N_4289,N_4130);
nand U5897 (N_5897,N_3293,N_3047);
nor U5898 (N_5898,N_4476,N_3928);
nand U5899 (N_5899,N_3674,N_3989);
and U5900 (N_5900,N_4161,N_3708);
nor U5901 (N_5901,N_3818,N_3708);
nand U5902 (N_5902,N_4326,N_3118);
xor U5903 (N_5903,N_3687,N_4285);
or U5904 (N_5904,N_3986,N_3972);
nor U5905 (N_5905,N_4484,N_3297);
xnor U5906 (N_5906,N_3274,N_3493);
and U5907 (N_5907,N_4169,N_4162);
nor U5908 (N_5908,N_3970,N_3510);
nor U5909 (N_5909,N_4429,N_3091);
nor U5910 (N_5910,N_3947,N_3561);
nand U5911 (N_5911,N_3370,N_3863);
nand U5912 (N_5912,N_4154,N_4363);
nor U5913 (N_5913,N_4029,N_3880);
nand U5914 (N_5914,N_3827,N_4263);
nor U5915 (N_5915,N_3963,N_3822);
and U5916 (N_5916,N_3161,N_3338);
nor U5917 (N_5917,N_3551,N_4213);
nand U5918 (N_5918,N_3600,N_3562);
or U5919 (N_5919,N_4264,N_3090);
nand U5920 (N_5920,N_4373,N_4004);
and U5921 (N_5921,N_4061,N_3025);
nor U5922 (N_5922,N_3472,N_3948);
and U5923 (N_5923,N_4188,N_3628);
or U5924 (N_5924,N_3131,N_3432);
nand U5925 (N_5925,N_3556,N_4416);
nand U5926 (N_5926,N_3845,N_3887);
and U5927 (N_5927,N_4020,N_3680);
nor U5928 (N_5928,N_3642,N_3292);
nor U5929 (N_5929,N_4315,N_4465);
or U5930 (N_5930,N_3327,N_4150);
xor U5931 (N_5931,N_4141,N_4413);
and U5932 (N_5932,N_4080,N_3859);
xnor U5933 (N_5933,N_3621,N_3355);
and U5934 (N_5934,N_4295,N_3169);
nand U5935 (N_5935,N_3640,N_3188);
nand U5936 (N_5936,N_3155,N_3254);
xnor U5937 (N_5937,N_3662,N_3728);
xnor U5938 (N_5938,N_3424,N_3499);
nand U5939 (N_5939,N_3386,N_3902);
nand U5940 (N_5940,N_3791,N_3158);
nand U5941 (N_5941,N_3751,N_4094);
or U5942 (N_5942,N_3413,N_3693);
nand U5943 (N_5943,N_3516,N_3217);
nor U5944 (N_5944,N_3398,N_3066);
nor U5945 (N_5945,N_3462,N_3395);
nand U5946 (N_5946,N_3336,N_3206);
nand U5947 (N_5947,N_3482,N_3336);
or U5948 (N_5948,N_3368,N_3660);
nor U5949 (N_5949,N_3024,N_3969);
nand U5950 (N_5950,N_3861,N_4140);
and U5951 (N_5951,N_3430,N_3737);
nor U5952 (N_5952,N_3033,N_4214);
nand U5953 (N_5953,N_3798,N_4473);
and U5954 (N_5954,N_3602,N_3900);
or U5955 (N_5955,N_3330,N_3927);
nor U5956 (N_5956,N_3083,N_4401);
nor U5957 (N_5957,N_3106,N_3896);
nor U5958 (N_5958,N_3634,N_4493);
nor U5959 (N_5959,N_3075,N_3617);
and U5960 (N_5960,N_3797,N_4234);
and U5961 (N_5961,N_3216,N_3433);
and U5962 (N_5962,N_4166,N_3093);
nand U5963 (N_5963,N_4287,N_4049);
nand U5964 (N_5964,N_4092,N_4397);
and U5965 (N_5965,N_3926,N_3594);
or U5966 (N_5966,N_3192,N_3998);
nor U5967 (N_5967,N_3272,N_3477);
and U5968 (N_5968,N_4360,N_3705);
nand U5969 (N_5969,N_4352,N_3597);
nor U5970 (N_5970,N_3623,N_4452);
or U5971 (N_5971,N_3722,N_3973);
xnor U5972 (N_5972,N_3539,N_3410);
and U5973 (N_5973,N_3088,N_3221);
xor U5974 (N_5974,N_4484,N_4496);
xnor U5975 (N_5975,N_3246,N_3839);
xnor U5976 (N_5976,N_3522,N_4369);
and U5977 (N_5977,N_3494,N_4346);
nand U5978 (N_5978,N_3980,N_4176);
nor U5979 (N_5979,N_3870,N_3937);
nand U5980 (N_5980,N_4254,N_4186);
xnor U5981 (N_5981,N_3884,N_3635);
xnor U5982 (N_5982,N_4020,N_3712);
and U5983 (N_5983,N_3943,N_3818);
nor U5984 (N_5984,N_3356,N_3664);
or U5985 (N_5985,N_4239,N_4472);
nor U5986 (N_5986,N_4356,N_3918);
xor U5987 (N_5987,N_3434,N_3815);
nand U5988 (N_5988,N_4081,N_3560);
nand U5989 (N_5989,N_4318,N_4224);
xor U5990 (N_5990,N_3584,N_4332);
and U5991 (N_5991,N_3086,N_3461);
nor U5992 (N_5992,N_3396,N_4126);
xnor U5993 (N_5993,N_4173,N_3402);
nand U5994 (N_5994,N_4467,N_4211);
and U5995 (N_5995,N_4373,N_3851);
nor U5996 (N_5996,N_3781,N_4122);
xnor U5997 (N_5997,N_3930,N_3510);
nor U5998 (N_5998,N_3562,N_3577);
or U5999 (N_5999,N_3866,N_3068);
nand U6000 (N_6000,N_4737,N_4588);
xor U6001 (N_6001,N_5380,N_5734);
nand U6002 (N_6002,N_4869,N_5056);
nand U6003 (N_6003,N_4527,N_5182);
or U6004 (N_6004,N_5198,N_5565);
nor U6005 (N_6005,N_4768,N_5648);
and U6006 (N_6006,N_4924,N_5299);
or U6007 (N_6007,N_4893,N_5132);
xnor U6008 (N_6008,N_5339,N_5121);
nand U6009 (N_6009,N_4888,N_5032);
nor U6010 (N_6010,N_5956,N_4595);
and U6011 (N_6011,N_5472,N_5174);
nand U6012 (N_6012,N_4554,N_5184);
and U6013 (N_6013,N_4782,N_5438);
and U6014 (N_6014,N_4636,N_5622);
and U6015 (N_6015,N_5289,N_5509);
and U6016 (N_6016,N_5682,N_5768);
nand U6017 (N_6017,N_5569,N_4659);
or U6018 (N_6018,N_5275,N_4991);
nand U6019 (N_6019,N_4596,N_5863);
nand U6020 (N_6020,N_5270,N_5076);
and U6021 (N_6021,N_5104,N_5952);
or U6022 (N_6022,N_5852,N_4531);
nand U6023 (N_6023,N_5467,N_5235);
nor U6024 (N_6024,N_5619,N_5115);
nor U6025 (N_6025,N_5733,N_5798);
or U6026 (N_6026,N_5074,N_5628);
nor U6027 (N_6027,N_5212,N_5990);
nor U6028 (N_6028,N_5613,N_5581);
nand U6029 (N_6029,N_5240,N_4637);
or U6030 (N_6030,N_5048,N_5356);
xnor U6031 (N_6031,N_5541,N_5302);
or U6032 (N_6032,N_5858,N_4619);
and U6033 (N_6033,N_5873,N_4598);
xor U6034 (N_6034,N_5804,N_5382);
nand U6035 (N_6035,N_5111,N_4961);
nor U6036 (N_6036,N_5333,N_4909);
nor U6037 (N_6037,N_4847,N_4952);
xor U6038 (N_6038,N_5429,N_5567);
xor U6039 (N_6039,N_5582,N_5075);
nand U6040 (N_6040,N_4803,N_4901);
xor U6041 (N_6041,N_5037,N_5345);
and U6042 (N_6042,N_5757,N_4727);
xnor U6043 (N_6043,N_5815,N_5741);
xnor U6044 (N_6044,N_4953,N_5532);
and U6045 (N_6045,N_5506,N_5978);
or U6046 (N_6046,N_4826,N_5637);
or U6047 (N_6047,N_5984,N_5266);
or U6048 (N_6048,N_5829,N_4797);
xnor U6049 (N_6049,N_5477,N_5045);
xor U6050 (N_6050,N_5096,N_5624);
xnor U6051 (N_6051,N_5416,N_4730);
or U6052 (N_6052,N_5540,N_4992);
xor U6053 (N_6053,N_5727,N_5608);
nor U6054 (N_6054,N_5611,N_5267);
or U6055 (N_6055,N_5315,N_4760);
nor U6056 (N_6056,N_5676,N_5775);
xnor U6057 (N_6057,N_5888,N_5911);
and U6058 (N_6058,N_5683,N_5411);
nor U6059 (N_6059,N_4834,N_4642);
or U6060 (N_6060,N_5495,N_4950);
xor U6061 (N_6061,N_4763,N_5760);
or U6062 (N_6062,N_5549,N_5644);
nor U6063 (N_6063,N_5042,N_4646);
nor U6064 (N_6064,N_5861,N_5141);
or U6065 (N_6065,N_5112,N_5718);
nor U6066 (N_6066,N_4544,N_5072);
nor U6067 (N_6067,N_4511,N_5378);
nor U6068 (N_6068,N_5153,N_5964);
xor U6069 (N_6069,N_4623,N_5234);
nor U6070 (N_6070,N_5246,N_4603);
and U6071 (N_6071,N_4668,N_5636);
and U6072 (N_6072,N_4923,N_4703);
nand U6073 (N_6073,N_5685,N_4752);
nand U6074 (N_6074,N_4621,N_5418);
nand U6075 (N_6075,N_5519,N_4699);
and U6076 (N_6076,N_5067,N_5038);
xnor U6077 (N_6077,N_5457,N_5334);
nand U6078 (N_6078,N_5918,N_5154);
and U6079 (N_6079,N_4805,N_5763);
xnor U6080 (N_6080,N_5179,N_5460);
xor U6081 (N_6081,N_4687,N_5157);
nand U6082 (N_6082,N_5313,N_5440);
or U6083 (N_6083,N_5152,N_5951);
or U6084 (N_6084,N_4874,N_4759);
nor U6085 (N_6085,N_4656,N_5558);
nand U6086 (N_6086,N_4678,N_4962);
nand U6087 (N_6087,N_4812,N_5082);
nor U6088 (N_6088,N_4829,N_5196);
or U6089 (N_6089,N_5709,N_5747);
or U6090 (N_6090,N_4784,N_4916);
xor U6091 (N_6091,N_5982,N_5503);
xor U6092 (N_6092,N_5276,N_5372);
nand U6093 (N_6093,N_5106,N_4848);
xor U6094 (N_6094,N_5921,N_4628);
or U6095 (N_6095,N_5980,N_4648);
nand U6096 (N_6096,N_5916,N_4535);
or U6097 (N_6097,N_5499,N_5677);
nor U6098 (N_6098,N_4547,N_4618);
nor U6099 (N_6099,N_4529,N_4605);
xnor U6100 (N_6100,N_4852,N_5046);
nor U6101 (N_6101,N_4778,N_5068);
or U6102 (N_6102,N_4921,N_5263);
xor U6103 (N_6103,N_5109,N_5227);
nand U6104 (N_6104,N_5512,N_5219);
nor U6105 (N_6105,N_5208,N_5823);
or U6106 (N_6106,N_5486,N_4721);
nor U6107 (N_6107,N_5364,N_4626);
xnor U6108 (N_6108,N_5925,N_5099);
and U6109 (N_6109,N_5249,N_5343);
or U6110 (N_6110,N_5209,N_5552);
nor U6111 (N_6111,N_5946,N_5870);
nand U6112 (N_6112,N_5011,N_5363);
and U6113 (N_6113,N_4809,N_5568);
nor U6114 (N_6114,N_4503,N_5794);
and U6115 (N_6115,N_4741,N_5802);
or U6116 (N_6116,N_4692,N_5933);
nand U6117 (N_6117,N_5642,N_5094);
nor U6118 (N_6118,N_4917,N_4640);
or U6119 (N_6119,N_4689,N_5087);
nand U6120 (N_6120,N_4611,N_4684);
nor U6121 (N_6121,N_5846,N_5365);
or U6122 (N_6122,N_5195,N_4616);
or U6123 (N_6123,N_5488,N_5500);
nand U6124 (N_6124,N_5441,N_5772);
or U6125 (N_6125,N_4858,N_5756);
nor U6126 (N_6126,N_4612,N_5765);
nand U6127 (N_6127,N_4577,N_4918);
and U6128 (N_6128,N_5728,N_4823);
nand U6129 (N_6129,N_5905,N_4697);
and U6130 (N_6130,N_5721,N_4548);
nor U6131 (N_6131,N_4886,N_5653);
nand U6132 (N_6132,N_4570,N_4584);
or U6133 (N_6133,N_5556,N_5833);
nor U6134 (N_6134,N_5049,N_4824);
or U6135 (N_6135,N_5928,N_5023);
or U6136 (N_6136,N_5865,N_5373);
nand U6137 (N_6137,N_4549,N_5415);
or U6138 (N_6138,N_4690,N_5406);
and U6139 (N_6139,N_5792,N_5158);
xor U6140 (N_6140,N_4538,N_5882);
nor U6141 (N_6141,N_5239,N_4941);
nor U6142 (N_6142,N_5003,N_5137);
nor U6143 (N_6143,N_4658,N_4542);
and U6144 (N_6144,N_5024,N_5253);
xnor U6145 (N_6145,N_5889,N_5680);
or U6146 (N_6146,N_4543,N_5959);
nor U6147 (N_6147,N_4594,N_5405);
nand U6148 (N_6148,N_5831,N_4701);
nor U6149 (N_6149,N_5265,N_5183);
or U6150 (N_6150,N_5502,N_5534);
xor U6151 (N_6151,N_4682,N_5919);
xor U6152 (N_6152,N_5890,N_4739);
nor U6153 (N_6153,N_4736,N_4988);
nand U6154 (N_6154,N_5566,N_4832);
or U6155 (N_6155,N_5572,N_5430);
nand U6156 (N_6156,N_5767,N_4910);
nor U6157 (N_6157,N_5465,N_5259);
xnor U6158 (N_6158,N_4993,N_5997);
and U6159 (N_6159,N_5052,N_4558);
nand U6160 (N_6160,N_4982,N_5555);
and U6161 (N_6161,N_5230,N_5687);
or U6162 (N_6162,N_4974,N_5207);
or U6163 (N_6163,N_5017,N_4517);
and U6164 (N_6164,N_4513,N_4560);
nand U6165 (N_6165,N_4995,N_5142);
and U6166 (N_6166,N_5779,N_5001);
xnor U6167 (N_6167,N_4716,N_5362);
nor U6168 (N_6168,N_5401,N_4892);
nor U6169 (N_6169,N_5494,N_4973);
nand U6170 (N_6170,N_4674,N_5960);
xnor U6171 (N_6171,N_5523,N_5987);
xor U6172 (N_6172,N_5623,N_4706);
nand U6173 (N_6173,N_5645,N_5092);
nand U6174 (N_6174,N_5146,N_4841);
or U6175 (N_6175,N_5303,N_5497);
or U6176 (N_6176,N_5796,N_5224);
and U6177 (N_6177,N_5191,N_5963);
and U6178 (N_6178,N_5386,N_5971);
or U6179 (N_6179,N_5291,N_4860);
or U6180 (N_6180,N_5114,N_5453);
and U6181 (N_6181,N_5412,N_4602);
and U6182 (N_6182,N_4683,N_5319);
and U6183 (N_6183,N_5998,N_4694);
or U6184 (N_6184,N_4839,N_5220);
nor U6185 (N_6185,N_5290,N_5755);
xor U6186 (N_6186,N_4561,N_4601);
xor U6187 (N_6187,N_5525,N_4757);
nand U6188 (N_6188,N_4857,N_5791);
nand U6189 (N_6189,N_5696,N_5216);
or U6190 (N_6190,N_5071,N_5055);
nand U6191 (N_6191,N_5818,N_5433);
nor U6192 (N_6192,N_5520,N_5533);
nor U6193 (N_6193,N_5140,N_5836);
nand U6194 (N_6194,N_4911,N_5251);
or U6195 (N_6195,N_5922,N_4903);
xnor U6196 (N_6196,N_5716,N_5837);
xnor U6197 (N_6197,N_5012,N_4855);
xnor U6198 (N_6198,N_5840,N_4766);
nand U6199 (N_6199,N_4981,N_5394);
or U6200 (N_6200,N_5487,N_5475);
nor U6201 (N_6201,N_4740,N_4735);
and U6202 (N_6202,N_5658,N_4607);
nor U6203 (N_6203,N_5222,N_4976);
and U6204 (N_6204,N_5173,N_5670);
nand U6205 (N_6205,N_5827,N_4708);
nor U6206 (N_6206,N_4504,N_5314);
nand U6207 (N_6207,N_5039,N_5812);
and U6208 (N_6208,N_4541,N_5147);
nand U6209 (N_6209,N_5744,N_5341);
and U6210 (N_6210,N_4775,N_5879);
or U6211 (N_6211,N_4661,N_4828);
and U6212 (N_6212,N_5579,N_5213);
xor U6213 (N_6213,N_4807,N_5876);
or U6214 (N_6214,N_5553,N_5317);
nor U6215 (N_6215,N_5102,N_5590);
xnor U6216 (N_6216,N_4959,N_4927);
and U6217 (N_6217,N_4672,N_5561);
nor U6218 (N_6218,N_5193,N_5409);
or U6219 (N_6219,N_5742,N_4745);
nand U6220 (N_6220,N_5704,N_4966);
nand U6221 (N_6221,N_5088,N_4615);
or U6222 (N_6222,N_5813,N_4792);
nor U6223 (N_6223,N_4764,N_5413);
nand U6224 (N_6224,N_5217,N_4526);
nor U6225 (N_6225,N_4500,N_5535);
nand U6226 (N_6226,N_4508,N_5664);
xor U6227 (N_6227,N_4875,N_4902);
and U6228 (N_6228,N_4583,N_5439);
nand U6229 (N_6229,N_4553,N_5156);
xor U6230 (N_6230,N_5854,N_4610);
or U6231 (N_6231,N_4800,N_4505);
and U6232 (N_6232,N_5464,N_4705);
and U6233 (N_6233,N_5754,N_4691);
xnor U6234 (N_6234,N_5204,N_5910);
nand U6235 (N_6235,N_5245,N_5641);
xnor U6236 (N_6236,N_5348,N_5025);
and U6237 (N_6237,N_4753,N_5793);
and U6238 (N_6238,N_5887,N_5992);
nand U6239 (N_6239,N_5414,N_5058);
xor U6240 (N_6240,N_5404,N_4790);
nand U6241 (N_6241,N_4788,N_5949);
and U6242 (N_6242,N_4733,N_4871);
or U6243 (N_6243,N_5301,N_5857);
and U6244 (N_6244,N_5563,N_5008);
or U6245 (N_6245,N_5371,N_5178);
and U6246 (N_6246,N_5934,N_4887);
or U6247 (N_6247,N_5507,N_5399);
nand U6248 (N_6248,N_4986,N_5434);
xnor U6249 (N_6249,N_5746,N_5221);
or U6250 (N_6250,N_4806,N_4882);
nor U6251 (N_6251,N_5724,N_5458);
nand U6252 (N_6252,N_5390,N_5669);
xor U6253 (N_6253,N_5101,N_5701);
xor U6254 (N_6254,N_4681,N_5242);
and U6255 (N_6255,N_4532,N_5972);
xor U6256 (N_6256,N_5659,N_5737);
and U6257 (N_6257,N_4557,N_4710);
xnor U6258 (N_6258,N_5451,N_5929);
nand U6259 (N_6259,N_5163,N_4794);
nand U6260 (N_6260,N_4506,N_5607);
xnor U6261 (N_6261,N_4704,N_5450);
xnor U6262 (N_6262,N_5300,N_5842);
and U6263 (N_6263,N_5867,N_5410);
and U6264 (N_6264,N_5924,N_5822);
nand U6265 (N_6265,N_5395,N_5803);
or U6266 (N_6266,N_5164,N_5841);
and U6267 (N_6267,N_5376,N_5797);
nor U6268 (N_6268,N_4622,N_4914);
nand U6269 (N_6269,N_5604,N_4769);
nand U6270 (N_6270,N_4641,N_5554);
nand U6271 (N_6271,N_4589,N_4592);
nor U6272 (N_6272,N_4945,N_5626);
or U6273 (N_6273,N_5859,N_4677);
or U6274 (N_6274,N_4849,N_5279);
xor U6275 (N_6275,N_5015,N_5736);
xnor U6276 (N_6276,N_5448,N_5318);
xnor U6277 (N_6277,N_4749,N_4624);
nand U6278 (N_6278,N_5228,N_5233);
nor U6279 (N_6279,N_5599,N_5596);
xor U6280 (N_6280,N_4780,N_4669);
nand U6281 (N_6281,N_5897,N_4946);
nand U6282 (N_6282,N_5332,N_5907);
xnor U6283 (N_6283,N_4540,N_5580);
and U6284 (N_6284,N_4702,N_4937);
nand U6285 (N_6285,N_5389,N_4891);
xnor U6286 (N_6286,N_5618,N_5832);
and U6287 (N_6287,N_5965,N_5526);
nand U6288 (N_6288,N_5693,N_5155);
xor U6289 (N_6289,N_5381,N_5387);
nand U6290 (N_6290,N_5702,N_4779);
or U6291 (N_6291,N_5098,N_5469);
nor U6292 (N_6292,N_4821,N_5277);
and U6293 (N_6293,N_5546,N_4864);
and U6294 (N_6294,N_5600,N_4879);
or U6295 (N_6295,N_4578,N_5282);
xor U6296 (N_6296,N_4890,N_4932);
nand U6297 (N_6297,N_5631,N_4836);
nor U6298 (N_6298,N_5501,N_5398);
nor U6299 (N_6299,N_5684,N_5528);
and U6300 (N_6300,N_4748,N_5605);
and U6301 (N_6301,N_5481,N_4997);
nor U6302 (N_6302,N_5562,N_4719);
xor U6303 (N_6303,N_5570,N_5205);
xnor U6304 (N_6304,N_5036,N_5397);
or U6305 (N_6305,N_5914,N_5284);
nor U6306 (N_6306,N_4854,N_4666);
nand U6307 (N_6307,N_5712,N_5384);
or U6308 (N_6308,N_4808,N_5118);
nor U6309 (N_6309,N_5172,N_5128);
nor U6310 (N_6310,N_5337,N_4825);
nand U6311 (N_6311,N_4556,N_5126);
and U6312 (N_6312,N_4777,N_4660);
nand U6313 (N_6313,N_5771,N_5447);
nor U6314 (N_6314,N_5835,N_4754);
nor U6315 (N_6315,N_4522,N_5508);
and U6316 (N_6316,N_5627,N_5199);
xnor U6317 (N_6317,N_4725,N_4580);
nor U6318 (N_6318,N_4518,N_5824);
or U6319 (N_6319,N_5407,N_5969);
and U6320 (N_6320,N_5989,N_5442);
and U6321 (N_6321,N_5306,N_5085);
and U6322 (N_6322,N_4644,N_5781);
or U6323 (N_6323,N_5368,N_5629);
xnor U6324 (N_6324,N_4845,N_4655);
nand U6325 (N_6325,N_4707,N_5800);
and U6326 (N_6326,N_4520,N_5367);
or U6327 (N_6327,N_4653,N_5762);
or U6328 (N_6328,N_4731,N_5480);
and U6329 (N_6329,N_5720,N_4546);
and U6330 (N_6330,N_5238,N_5483);
or U6331 (N_6331,N_5869,N_5160);
nand U6332 (N_6332,N_5749,N_5272);
or U6333 (N_6333,N_5188,N_4843);
nand U6334 (N_6334,N_5241,N_4799);
nor U6335 (N_6335,N_4955,N_5328);
xor U6336 (N_6336,N_5961,N_5322);
nand U6337 (N_6337,N_5077,N_5258);
xnor U6338 (N_6338,N_4712,N_5493);
nand U6339 (N_6339,N_5028,N_4559);
and U6340 (N_6340,N_4604,N_5150);
xnor U6341 (N_6341,N_5811,N_5993);
and U6342 (N_6342,N_5510,N_5892);
xor U6343 (N_6343,N_5491,N_4600);
nor U6344 (N_6344,N_5575,N_5666);
or U6345 (N_6345,N_4830,N_5041);
xnor U6346 (N_6346,N_5034,N_5551);
or U6347 (N_6347,N_4724,N_5828);
nor U6348 (N_6348,N_5856,N_5923);
nor U6349 (N_6349,N_5054,N_5260);
nand U6350 (N_6350,N_4856,N_5171);
xor U6351 (N_6351,N_4969,N_5725);
xnor U6352 (N_6352,N_4726,N_4671);
nor U6353 (N_6353,N_4853,N_4850);
nor U6354 (N_6354,N_5583,N_4545);
xnor U6355 (N_6355,N_5937,N_4865);
xor U6356 (N_6356,N_4732,N_4563);
xor U6357 (N_6357,N_5005,N_5695);
xor U6358 (N_6358,N_5091,N_5672);
xnor U6359 (N_6359,N_5654,N_4873);
xor U6360 (N_6360,N_4685,N_5051);
nand U6361 (N_6361,N_5557,N_4863);
xnor U6362 (N_6362,N_5950,N_5906);
xor U6363 (N_6363,N_4620,N_5954);
xnor U6364 (N_6364,N_5388,N_5148);
and U6365 (N_6365,N_5983,N_4944);
and U6366 (N_6366,N_5930,N_5084);
xor U6367 (N_6367,N_5538,N_4512);
and U6368 (N_6368,N_4550,N_5116);
nor U6369 (N_6369,N_4936,N_4591);
and U6370 (N_6370,N_5452,N_5711);
nand U6371 (N_6371,N_5789,N_5655);
xor U6372 (N_6372,N_5252,N_5715);
xnor U6373 (N_6373,N_5123,N_5939);
xor U6374 (N_6374,N_4536,N_5675);
nor U6375 (N_6375,N_5957,N_5967);
xor U6376 (N_6376,N_5329,N_5120);
xor U6377 (N_6377,N_5283,N_5660);
and U6378 (N_6378,N_5524,N_4709);
nand U6379 (N_6379,N_5995,N_5262);
and U6380 (N_6380,N_5714,N_5776);
and U6381 (N_6381,N_5543,N_4787);
nor U6382 (N_6382,N_5625,N_5592);
nand U6383 (N_6383,N_5606,N_5639);
and U6384 (N_6384,N_4781,N_5316);
and U6385 (N_6385,N_5287,N_4625);
and U6386 (N_6386,N_5254,N_5649);
nor U6387 (N_6387,N_4978,N_5901);
nor U6388 (N_6388,N_4958,N_5635);
nand U6389 (N_6389,N_5336,N_5994);
and U6390 (N_6390,N_4811,N_5927);
nor U6391 (N_6391,N_4922,N_5587);
xnor U6392 (N_6392,N_4851,N_4816);
or U6393 (N_6393,N_4729,N_5026);
nor U6394 (N_6394,N_5559,N_5926);
nand U6395 (N_6395,N_5681,N_4817);
nand U6396 (N_6396,N_4771,N_5874);
xor U6397 (N_6397,N_5466,N_4762);
or U6398 (N_6398,N_5589,N_4534);
nor U6399 (N_6399,N_5594,N_5305);
and U6400 (N_6400,N_5866,N_4919);
nor U6401 (N_6401,N_5385,N_5663);
and U6402 (N_6402,N_4751,N_5443);
xor U6403 (N_6403,N_5062,N_5264);
nand U6404 (N_6404,N_5688,N_5795);
and U6405 (N_6405,N_5668,N_4663);
or U6406 (N_6406,N_5256,N_5880);
xnor U6407 (N_6407,N_5875,N_5144);
or U6408 (N_6408,N_4925,N_5656);
and U6409 (N_6409,N_5070,N_4931);
or U6410 (N_6410,N_5134,N_5293);
or U6411 (N_6411,N_4632,N_5877);
or U6412 (N_6412,N_5821,N_4996);
and U6413 (N_6413,N_4786,N_5029);
nor U6414 (N_6414,N_5621,N_5366);
xnor U6415 (N_6415,N_5105,N_4968);
xnor U6416 (N_6416,N_5002,N_5130);
or U6417 (N_6417,N_5324,N_5013);
and U6418 (N_6418,N_5358,N_5484);
xnor U6419 (N_6419,N_4838,N_4639);
or U6420 (N_6420,N_4539,N_4629);
or U6421 (N_6421,N_5165,N_5338);
nor U6422 (N_6422,N_5752,N_5043);
and U6423 (N_6423,N_5743,N_5027);
nor U6424 (N_6424,N_5761,N_5920);
nand U6425 (N_6425,N_5893,N_4894);
or U6426 (N_6426,N_5166,N_5177);
and U6427 (N_6427,N_5686,N_5780);
nand U6428 (N_6428,N_4552,N_4717);
nand U6429 (N_6429,N_5673,N_5269);
or U6430 (N_6430,N_4842,N_5690);
xnor U6431 (N_6431,N_5977,N_5189);
and U6432 (N_6432,N_5646,N_5312);
or U6433 (N_6433,N_5423,N_5138);
or U6434 (N_6434,N_5966,N_5202);
nand U6435 (N_6435,N_5564,N_4862);
or U6436 (N_6436,N_5192,N_5784);
nand U6437 (N_6437,N_5935,N_5853);
xor U6438 (N_6438,N_4574,N_4868);
and U6439 (N_6439,N_5975,N_4609);
and U6440 (N_6440,N_4920,N_5124);
nand U6441 (N_6441,N_5610,N_5325);
nor U6442 (N_6442,N_5110,N_5203);
nand U6443 (N_6443,N_4676,N_4840);
nor U6444 (N_6444,N_4928,N_5421);
nand U6445 (N_6445,N_5361,N_4688);
or U6446 (N_6446,N_5473,N_5307);
xor U6447 (N_6447,N_4957,N_4509);
or U6448 (N_6448,N_4964,N_5459);
nand U6449 (N_6449,N_5288,N_5790);
and U6450 (N_6450,N_5845,N_5518);
nand U6451 (N_6451,N_5243,N_5391);
nor U6452 (N_6452,N_5585,N_5229);
or U6453 (N_6453,N_5896,N_5131);
or U6454 (N_6454,N_5550,N_4715);
and U6455 (N_6455,N_5194,N_5539);
or U6456 (N_6456,N_4633,N_5446);
nor U6457 (N_6457,N_4796,N_5788);
or U6458 (N_6458,N_4835,N_4867);
nand U6459 (N_6459,N_4713,N_5197);
or U6460 (N_6460,N_5129,N_4586);
nor U6461 (N_6461,N_5425,N_4967);
nand U6462 (N_6462,N_4617,N_5516);
xor U6463 (N_6463,N_5504,N_4947);
and U6464 (N_6464,N_5090,N_4695);
xnor U6465 (N_6465,N_5586,N_5006);
xnor U6466 (N_6466,N_5424,N_5826);
and U6467 (N_6467,N_5601,N_4980);
nor U6468 (N_6468,N_4773,N_5069);
xnor U6469 (N_6469,N_5943,N_4569);
or U6470 (N_6470,N_5545,N_5047);
and U6471 (N_6471,N_5838,N_4861);
nand U6472 (N_6472,N_5855,N_5962);
and U6473 (N_6473,N_4872,N_5710);
xnor U6474 (N_6474,N_5176,N_5814);
nand U6475 (N_6475,N_5612,N_5958);
or U6476 (N_6476,N_5705,N_5825);
xor U6477 (N_6477,N_5435,N_4634);
or U6478 (N_6478,N_5170,N_5694);
xor U6479 (N_6479,N_5944,N_4744);
nor U6480 (N_6480,N_4900,N_5819);
xnor U6481 (N_6481,N_4934,N_5143);
nand U6482 (N_6482,N_5650,N_5310);
and U6483 (N_6483,N_4898,N_5432);
nand U6484 (N_6484,N_5657,N_5769);
or U6485 (N_6485,N_4951,N_4608);
and U6486 (N_6486,N_5296,N_5463);
and U6487 (N_6487,N_4822,N_5355);
and U6488 (N_6488,N_4645,N_4772);
and U6489 (N_6489,N_5326,N_4502);
or U6490 (N_6490,N_5280,N_5344);
nand U6491 (N_6491,N_5482,N_5571);
nand U6492 (N_6492,N_5089,N_5908);
xor U6493 (N_6493,N_5162,N_4567);
or U6494 (N_6494,N_5250,N_4878);
or U6495 (N_6495,N_5379,N_4804);
nand U6496 (N_6496,N_5019,N_5454);
or U6497 (N_6497,N_4614,N_5665);
nor U6498 (N_6498,N_5462,N_4907);
or U6499 (N_6499,N_5417,N_5999);
or U6500 (N_6500,N_4987,N_5139);
xor U6501 (N_6501,N_4523,N_5661);
nor U6502 (N_6502,N_4831,N_4728);
nand U6503 (N_6503,N_5375,N_4525);
or U6504 (N_6504,N_4665,N_5383);
xnor U6505 (N_6505,N_5536,N_5236);
or U6506 (N_6506,N_5020,N_5066);
or U6507 (N_6507,N_5133,N_5422);
nand U6508 (N_6508,N_5030,N_5898);
nand U6509 (N_6509,N_4747,N_4568);
nor U6510 (N_6510,N_5285,N_4994);
or U6511 (N_6511,N_4956,N_5033);
nor U6512 (N_6512,N_5374,N_4635);
xnor U6513 (N_6513,N_5360,N_5820);
nor U6514 (N_6514,N_4866,N_4643);
and U6515 (N_6515,N_5187,N_4813);
nand U6516 (N_6516,N_5717,N_4970);
and U6517 (N_6517,N_5168,N_5456);
and U6518 (N_6518,N_4696,N_4859);
nor U6519 (N_6519,N_5474,N_5151);
xor U6520 (N_6520,N_4587,N_5973);
xor U6521 (N_6521,N_4664,N_5490);
nand U6522 (N_6522,N_5547,N_4718);
nand U6523 (N_6523,N_4929,N_4515);
xor U6524 (N_6524,N_5891,N_4575);
nor U6525 (N_6525,N_4756,N_5215);
xnor U6526 (N_6526,N_5113,N_5948);
and U6527 (N_6527,N_5248,N_5774);
xnor U6528 (N_6528,N_5726,N_5231);
nand U6529 (N_6529,N_5745,N_5588);
nor U6530 (N_6530,N_5723,N_4582);
xnor U6531 (N_6531,N_4585,N_4990);
nand U6532 (N_6532,N_4983,N_5806);
or U6533 (N_6533,N_5782,N_5968);
nand U6534 (N_6534,N_5063,N_5040);
and U6535 (N_6535,N_4795,N_5022);
xor U6536 (N_6536,N_5671,N_5860);
nor U6537 (N_6537,N_5738,N_5485);
xnor U6538 (N_6538,N_4776,N_4770);
or U6539 (N_6539,N_5323,N_4734);
nor U6540 (N_6540,N_5255,N_4507);
and U6541 (N_6541,N_5640,N_5872);
and U6542 (N_6542,N_5273,N_5847);
or U6543 (N_6543,N_4758,N_4926);
xnor U6544 (N_6544,N_4579,N_5849);
and U6545 (N_6545,N_5584,N_5739);
xor U6546 (N_6546,N_5190,N_5468);
nor U6547 (N_6547,N_5830,N_5878);
xor U6548 (N_6548,N_5615,N_5713);
nor U6549 (N_6549,N_4789,N_5730);
or U6550 (N_6550,N_5009,N_5354);
xor U6551 (N_6551,N_5297,N_4963);
and U6552 (N_6552,N_5080,N_4791);
nand U6553 (N_6553,N_4652,N_4954);
or U6554 (N_6554,N_4638,N_4606);
xnor U6555 (N_6555,N_4528,N_5529);
xor U6556 (N_6556,N_5885,N_4999);
nand U6557 (N_6557,N_5991,N_4943);
nand U6558 (N_6558,N_5953,N_4884);
nor U6559 (N_6559,N_4647,N_4765);
and U6560 (N_6560,N_4649,N_5000);
xnor U6561 (N_6561,N_4514,N_5396);
nor U6562 (N_6562,N_4876,N_5359);
and U6563 (N_6563,N_4915,N_5044);
nand U6564 (N_6564,N_5909,N_5574);
xor U6565 (N_6565,N_5593,N_5595);
and U6566 (N_6566,N_5117,N_5521);
nor U6567 (N_6567,N_5785,N_5346);
nand U6568 (N_6568,N_5149,N_4593);
nor U6569 (N_6569,N_4576,N_5119);
nor U6570 (N_6570,N_5591,N_5810);
nand U6571 (N_6571,N_4870,N_4975);
nand U6572 (N_6572,N_4897,N_5634);
or U6573 (N_6573,N_5751,N_5941);
or U6574 (N_6574,N_4913,N_4698);
nand U6575 (N_6575,N_5942,N_5748);
nor U6576 (N_6576,N_4537,N_5979);
nand U6577 (N_6577,N_5308,N_5514);
or U6578 (N_6578,N_5181,N_4761);
and U6579 (N_6579,N_5232,N_4519);
nor U6580 (N_6580,N_4820,N_4572);
nand U6581 (N_6581,N_5237,N_5201);
nand U6582 (N_6582,N_5498,N_5735);
nand U6583 (N_6583,N_5577,N_5136);
and U6584 (N_6584,N_4711,N_5848);
or U6585 (N_6585,N_4679,N_5408);
or U6586 (N_6586,N_5211,N_5392);
or U6587 (N_6587,N_5335,N_5161);
xnor U6588 (N_6588,N_5548,N_4627);
nor U6589 (N_6589,N_5304,N_5834);
nor U6590 (N_6590,N_5616,N_5976);
or U6591 (N_6591,N_5729,N_5035);
or U6592 (N_6592,N_5431,N_4613);
nor U6593 (N_6593,N_5320,N_5708);
and U6594 (N_6594,N_4889,N_5899);
or U6595 (N_6595,N_5955,N_4555);
xnor U6596 (N_6596,N_5370,N_5759);
nand U6597 (N_6597,N_5352,N_4722);
xor U6598 (N_6598,N_4599,N_4979);
nand U6599 (N_6599,N_5515,N_5706);
or U6600 (N_6600,N_4720,N_5214);
and U6601 (N_6601,N_4814,N_5620);
xor U6602 (N_6602,N_5268,N_4827);
nand U6603 (N_6603,N_5478,N_4673);
xnor U6604 (N_6604,N_4533,N_5369);
xnor U6605 (N_6605,N_5881,N_5489);
and U6606 (N_6606,N_5513,N_5061);
nor U6607 (N_6607,N_5732,N_5347);
or U6608 (N_6608,N_5805,N_5786);
nor U6609 (N_6609,N_5783,N_4885);
and U6610 (N_6610,N_5200,N_4524);
nor U6611 (N_6611,N_5602,N_5932);
nor U6612 (N_6612,N_5004,N_5083);
or U6613 (N_6613,N_5479,N_5122);
nor U6614 (N_6614,N_5689,N_5281);
xnor U6615 (N_6615,N_4742,N_5614);
and U6616 (N_6616,N_4948,N_5505);
nand U6617 (N_6617,N_5135,N_5816);
nor U6618 (N_6618,N_4904,N_4895);
nor U6619 (N_6619,N_4942,N_4905);
nand U6620 (N_6620,N_5722,N_5678);
nor U6621 (N_6621,N_5206,N_4743);
or U6622 (N_6622,N_5900,N_4802);
xnor U6623 (N_6623,N_5377,N_4798);
nand U6624 (N_6624,N_5638,N_5808);
xor U6625 (N_6625,N_5517,N_4785);
or U6626 (N_6626,N_5342,N_4564);
xor U6627 (N_6627,N_5393,N_5125);
nor U6628 (N_6628,N_5773,N_5597);
and U6629 (N_6629,N_5904,N_5286);
nand U6630 (N_6630,N_4977,N_4935);
or U6631 (N_6631,N_4670,N_5850);
and U6632 (N_6632,N_5010,N_4837);
nand U6633 (N_6633,N_5309,N_5261);
xor U6634 (N_6634,N_5617,N_5471);
nor U6635 (N_6635,N_4750,N_5186);
or U6636 (N_6636,N_4662,N_5697);
nand U6637 (N_6637,N_5097,N_5330);
xor U6638 (N_6638,N_4939,N_4971);
or U6639 (N_6639,N_4844,N_5886);
xor U6640 (N_6640,N_4984,N_4818);
nand U6641 (N_6641,N_5449,N_5349);
and U6642 (N_6642,N_5169,N_5988);
nor U6643 (N_6643,N_5210,N_4846);
and U6644 (N_6644,N_4940,N_5603);
nand U6645 (N_6645,N_5014,N_5719);
and U6646 (N_6646,N_5544,N_5100);
or U6647 (N_6647,N_5257,N_5703);
or U6648 (N_6648,N_4833,N_5679);
nand U6649 (N_6649,N_5321,N_5353);
nand U6650 (N_6650,N_4998,N_5652);
xnor U6651 (N_6651,N_4675,N_5073);
nor U6652 (N_6652,N_5428,N_4521);
nor U6653 (N_6653,N_4906,N_5476);
and U6654 (N_6654,N_5103,N_5884);
nand U6655 (N_6655,N_4985,N_4930);
or U6656 (N_6656,N_4783,N_5630);
and U6657 (N_6657,N_5403,N_5651);
xnor U6658 (N_6658,N_4746,N_4571);
nand U6659 (N_6659,N_5985,N_5917);
xor U6660 (N_6660,N_4657,N_5298);
xnor U6661 (N_6661,N_5021,N_4880);
nand U6662 (N_6662,N_4899,N_4597);
nand U6663 (N_6663,N_4723,N_4877);
xnor U6664 (N_6664,N_5167,N_5492);
and U6665 (N_6665,N_4738,N_5936);
and U6666 (N_6666,N_5064,N_4516);
or U6667 (N_6667,N_5970,N_5753);
or U6668 (N_6668,N_5692,N_4651);
nor U6669 (N_6669,N_5809,N_5931);
nor U6670 (N_6670,N_4686,N_5839);
and U6671 (N_6671,N_5667,N_5981);
nor U6672 (N_6672,N_4680,N_5086);
and U6673 (N_6673,N_5894,N_4810);
and U6674 (N_6674,N_4774,N_5511);
and U6675 (N_6675,N_5292,N_5057);
nor U6676 (N_6676,N_5851,N_4510);
and U6677 (N_6677,N_5095,N_4573);
nor U6678 (N_6678,N_5461,N_5445);
nor U6679 (N_6679,N_5226,N_5400);
nand U6680 (N_6680,N_5108,N_5331);
xor U6681 (N_6681,N_5185,N_5766);
nand U6682 (N_6682,N_5127,N_5764);
nand U6683 (N_6683,N_5175,N_5145);
xnor U6684 (N_6684,N_5598,N_4933);
nor U6685 (N_6685,N_4551,N_5527);
and U6686 (N_6686,N_5159,N_4562);
xnor U6687 (N_6687,N_5311,N_5542);
or U6688 (N_6688,N_5081,N_4501);
or U6689 (N_6689,N_5895,N_5294);
nand U6690 (N_6690,N_5427,N_4530);
nand U6691 (N_6691,N_5470,N_5740);
or U6692 (N_6692,N_5986,N_5560);
xor U6693 (N_6693,N_4960,N_5940);
or U6694 (N_6694,N_5225,N_5647);
or U6695 (N_6695,N_5609,N_4793);
or U6696 (N_6696,N_4965,N_5844);
or U6697 (N_6697,N_5522,N_4755);
nor U6698 (N_6698,N_5633,N_5915);
or U6699 (N_6699,N_4819,N_5868);
or U6700 (N_6700,N_5295,N_5912);
and U6701 (N_6701,N_5357,N_5691);
nand U6702 (N_6702,N_4912,N_5496);
nor U6703 (N_6703,N_5578,N_5674);
nor U6704 (N_6704,N_5787,N_5247);
or U6705 (N_6705,N_5938,N_5437);
or U6706 (N_6706,N_5271,N_4667);
nor U6707 (N_6707,N_5698,N_5244);
or U6708 (N_6708,N_5632,N_5079);
nand U6709 (N_6709,N_5059,N_4714);
nor U6710 (N_6710,N_4908,N_5974);
nand U6711 (N_6711,N_5945,N_4654);
or U6712 (N_6712,N_4938,N_5420);
and U6713 (N_6713,N_5707,N_4581);
nor U6714 (N_6714,N_5758,N_4767);
nand U6715 (N_6715,N_4989,N_5750);
nand U6716 (N_6716,N_4590,N_4650);
xnor U6717 (N_6717,N_5947,N_5700);
xor U6718 (N_6718,N_4693,N_5699);
or U6719 (N_6719,N_5770,N_5777);
nand U6720 (N_6720,N_5426,N_5274);
or U6721 (N_6721,N_5078,N_4972);
or U6722 (N_6722,N_5065,N_5018);
nor U6723 (N_6723,N_5843,N_5913);
xor U6724 (N_6724,N_5107,N_5643);
or U6725 (N_6725,N_5807,N_5537);
or U6726 (N_6726,N_5350,N_4815);
or U6727 (N_6727,N_4630,N_5996);
nor U6728 (N_6728,N_5531,N_5218);
nor U6729 (N_6729,N_4883,N_5419);
nor U6730 (N_6730,N_5903,N_4631);
nand U6731 (N_6731,N_5278,N_5731);
nor U6732 (N_6732,N_5436,N_5180);
xor U6733 (N_6733,N_5093,N_5799);
or U6734 (N_6734,N_5530,N_5576);
nor U6735 (N_6735,N_5662,N_5864);
or U6736 (N_6736,N_4565,N_5031);
or U6737 (N_6737,N_5444,N_5327);
or U6738 (N_6738,N_5871,N_5817);
and U6739 (N_6739,N_4801,N_5050);
and U6740 (N_6740,N_5053,N_5223);
nor U6741 (N_6741,N_5883,N_5455);
xor U6742 (N_6742,N_5778,N_4700);
nand U6743 (N_6743,N_5060,N_5573);
or U6744 (N_6744,N_5340,N_5007);
xor U6745 (N_6745,N_5862,N_5402);
and U6746 (N_6746,N_4949,N_5902);
nand U6747 (N_6747,N_5016,N_4566);
and U6748 (N_6748,N_5351,N_4881);
and U6749 (N_6749,N_5801,N_4896);
nand U6750 (N_6750,N_5538,N_5747);
or U6751 (N_6751,N_5293,N_4583);
or U6752 (N_6752,N_4751,N_5539);
and U6753 (N_6753,N_4654,N_5938);
or U6754 (N_6754,N_5217,N_5014);
xor U6755 (N_6755,N_5380,N_5813);
nand U6756 (N_6756,N_4659,N_5453);
nand U6757 (N_6757,N_5338,N_5724);
nand U6758 (N_6758,N_5214,N_4687);
nor U6759 (N_6759,N_4882,N_5687);
and U6760 (N_6760,N_4734,N_5474);
nor U6761 (N_6761,N_5007,N_5429);
or U6762 (N_6762,N_4505,N_5507);
and U6763 (N_6763,N_5240,N_5784);
or U6764 (N_6764,N_5354,N_5475);
nand U6765 (N_6765,N_4769,N_4988);
and U6766 (N_6766,N_5109,N_5215);
and U6767 (N_6767,N_5029,N_4509);
nor U6768 (N_6768,N_5590,N_5929);
and U6769 (N_6769,N_5231,N_4769);
xor U6770 (N_6770,N_5816,N_5033);
nor U6771 (N_6771,N_5766,N_5782);
and U6772 (N_6772,N_4763,N_5303);
xor U6773 (N_6773,N_5897,N_5040);
xor U6774 (N_6774,N_5079,N_5180);
and U6775 (N_6775,N_5960,N_5659);
xnor U6776 (N_6776,N_5801,N_5725);
xor U6777 (N_6777,N_5463,N_5466);
nand U6778 (N_6778,N_4808,N_4767);
or U6779 (N_6779,N_5403,N_5413);
xor U6780 (N_6780,N_4796,N_5631);
xnor U6781 (N_6781,N_4643,N_5128);
nor U6782 (N_6782,N_5865,N_4981);
and U6783 (N_6783,N_4644,N_5973);
and U6784 (N_6784,N_5640,N_4601);
or U6785 (N_6785,N_5646,N_5143);
or U6786 (N_6786,N_5338,N_5880);
nor U6787 (N_6787,N_4654,N_5959);
nor U6788 (N_6788,N_5213,N_4870);
xor U6789 (N_6789,N_5179,N_5132);
nand U6790 (N_6790,N_5872,N_5771);
xnor U6791 (N_6791,N_4949,N_5600);
xnor U6792 (N_6792,N_5697,N_5691);
nor U6793 (N_6793,N_5967,N_5475);
xor U6794 (N_6794,N_4787,N_5036);
nand U6795 (N_6795,N_5571,N_5855);
nor U6796 (N_6796,N_4909,N_5419);
nor U6797 (N_6797,N_4663,N_4939);
and U6798 (N_6798,N_5702,N_4882);
nand U6799 (N_6799,N_4880,N_5487);
xnor U6800 (N_6800,N_5361,N_4517);
nand U6801 (N_6801,N_4538,N_4744);
and U6802 (N_6802,N_5447,N_5250);
or U6803 (N_6803,N_4559,N_5432);
and U6804 (N_6804,N_4960,N_4607);
nand U6805 (N_6805,N_5403,N_4618);
nand U6806 (N_6806,N_4882,N_5070);
nand U6807 (N_6807,N_5981,N_5064);
or U6808 (N_6808,N_5021,N_5326);
nand U6809 (N_6809,N_5181,N_4506);
nor U6810 (N_6810,N_5607,N_5719);
nor U6811 (N_6811,N_5501,N_4737);
nand U6812 (N_6812,N_5273,N_5578);
and U6813 (N_6813,N_4631,N_5793);
nor U6814 (N_6814,N_4813,N_4948);
and U6815 (N_6815,N_4555,N_5738);
xor U6816 (N_6816,N_5572,N_4866);
and U6817 (N_6817,N_5204,N_5337);
or U6818 (N_6818,N_5306,N_5718);
nand U6819 (N_6819,N_5432,N_5024);
xnor U6820 (N_6820,N_5246,N_5626);
and U6821 (N_6821,N_4517,N_5312);
nand U6822 (N_6822,N_4910,N_5326);
or U6823 (N_6823,N_5203,N_5470);
xnor U6824 (N_6824,N_5127,N_5601);
xnor U6825 (N_6825,N_5419,N_5957);
xnor U6826 (N_6826,N_5951,N_5776);
nor U6827 (N_6827,N_5872,N_5642);
xnor U6828 (N_6828,N_4708,N_5622);
xnor U6829 (N_6829,N_4537,N_5865);
xor U6830 (N_6830,N_5575,N_4909);
or U6831 (N_6831,N_4840,N_5476);
and U6832 (N_6832,N_5134,N_5751);
nor U6833 (N_6833,N_4872,N_5570);
nor U6834 (N_6834,N_5004,N_4975);
or U6835 (N_6835,N_4903,N_5483);
or U6836 (N_6836,N_5525,N_4667);
xor U6837 (N_6837,N_5753,N_4675);
nor U6838 (N_6838,N_5655,N_4581);
or U6839 (N_6839,N_5112,N_5869);
and U6840 (N_6840,N_5910,N_5718);
nor U6841 (N_6841,N_4817,N_5978);
xor U6842 (N_6842,N_4773,N_4988);
nor U6843 (N_6843,N_5774,N_4643);
nor U6844 (N_6844,N_5492,N_5458);
nand U6845 (N_6845,N_4977,N_4544);
and U6846 (N_6846,N_4847,N_4887);
nand U6847 (N_6847,N_5681,N_4732);
nor U6848 (N_6848,N_5558,N_4749);
xnor U6849 (N_6849,N_5765,N_5029);
or U6850 (N_6850,N_4856,N_4933);
nand U6851 (N_6851,N_4632,N_5163);
and U6852 (N_6852,N_5789,N_5165);
nor U6853 (N_6853,N_5425,N_5004);
and U6854 (N_6854,N_5292,N_5066);
nor U6855 (N_6855,N_5141,N_5098);
nand U6856 (N_6856,N_4890,N_5837);
xor U6857 (N_6857,N_5914,N_5392);
or U6858 (N_6858,N_5647,N_5106);
xnor U6859 (N_6859,N_4951,N_4553);
or U6860 (N_6860,N_5777,N_5271);
nor U6861 (N_6861,N_4672,N_5602);
nor U6862 (N_6862,N_5997,N_4954);
xor U6863 (N_6863,N_4558,N_4604);
xor U6864 (N_6864,N_5551,N_5712);
nand U6865 (N_6865,N_5433,N_5317);
xor U6866 (N_6866,N_5917,N_4671);
or U6867 (N_6867,N_5008,N_5505);
xor U6868 (N_6868,N_4794,N_5185);
or U6869 (N_6869,N_4830,N_4882);
and U6870 (N_6870,N_5302,N_5200);
nand U6871 (N_6871,N_4987,N_4552);
xor U6872 (N_6872,N_4891,N_5552);
and U6873 (N_6873,N_4645,N_5136);
or U6874 (N_6874,N_5318,N_5976);
or U6875 (N_6875,N_5348,N_5796);
and U6876 (N_6876,N_5291,N_5465);
xnor U6877 (N_6877,N_5464,N_4816);
nand U6878 (N_6878,N_4603,N_5874);
xnor U6879 (N_6879,N_4986,N_5620);
xnor U6880 (N_6880,N_4895,N_5548);
nor U6881 (N_6881,N_5364,N_4777);
and U6882 (N_6882,N_5878,N_5745);
nor U6883 (N_6883,N_4755,N_5789);
or U6884 (N_6884,N_5387,N_5145);
and U6885 (N_6885,N_5346,N_4533);
and U6886 (N_6886,N_5853,N_5741);
xor U6887 (N_6887,N_5833,N_5050);
and U6888 (N_6888,N_5516,N_5810);
or U6889 (N_6889,N_4991,N_4872);
and U6890 (N_6890,N_5064,N_5875);
nand U6891 (N_6891,N_5403,N_5511);
and U6892 (N_6892,N_4796,N_4872);
and U6893 (N_6893,N_4811,N_5295);
or U6894 (N_6894,N_5138,N_5924);
nand U6895 (N_6895,N_5953,N_5106);
nand U6896 (N_6896,N_4518,N_5911);
or U6897 (N_6897,N_5411,N_4634);
nor U6898 (N_6898,N_5960,N_5241);
or U6899 (N_6899,N_5674,N_5158);
nor U6900 (N_6900,N_5309,N_5475);
nand U6901 (N_6901,N_5928,N_5884);
xnor U6902 (N_6902,N_5410,N_5379);
and U6903 (N_6903,N_5339,N_5676);
xnor U6904 (N_6904,N_5000,N_4642);
nor U6905 (N_6905,N_4721,N_5405);
and U6906 (N_6906,N_5535,N_4968);
and U6907 (N_6907,N_4902,N_5245);
nor U6908 (N_6908,N_5587,N_5243);
xor U6909 (N_6909,N_5256,N_5433);
nor U6910 (N_6910,N_4644,N_5645);
nor U6911 (N_6911,N_4625,N_5357);
nor U6912 (N_6912,N_5122,N_5602);
nor U6913 (N_6913,N_4693,N_5301);
or U6914 (N_6914,N_5355,N_5542);
xnor U6915 (N_6915,N_5216,N_4874);
and U6916 (N_6916,N_4514,N_5263);
and U6917 (N_6917,N_5439,N_4632);
nand U6918 (N_6918,N_5043,N_4784);
and U6919 (N_6919,N_5632,N_4697);
nor U6920 (N_6920,N_5249,N_4799);
or U6921 (N_6921,N_5881,N_4905);
or U6922 (N_6922,N_5533,N_5759);
nand U6923 (N_6923,N_5113,N_5525);
nor U6924 (N_6924,N_5103,N_5440);
and U6925 (N_6925,N_5840,N_5724);
nand U6926 (N_6926,N_5576,N_5407);
nor U6927 (N_6927,N_4957,N_4896);
xor U6928 (N_6928,N_5338,N_5357);
or U6929 (N_6929,N_5989,N_5609);
nand U6930 (N_6930,N_5123,N_5356);
and U6931 (N_6931,N_5530,N_5085);
xnor U6932 (N_6932,N_5181,N_5943);
nor U6933 (N_6933,N_4704,N_4541);
nor U6934 (N_6934,N_5060,N_4708);
xnor U6935 (N_6935,N_5778,N_5268);
nor U6936 (N_6936,N_5934,N_4845);
nor U6937 (N_6937,N_4566,N_5037);
nor U6938 (N_6938,N_4871,N_5001);
and U6939 (N_6939,N_4551,N_5319);
xnor U6940 (N_6940,N_4515,N_4901);
nand U6941 (N_6941,N_5554,N_5133);
nor U6942 (N_6942,N_5759,N_5768);
xnor U6943 (N_6943,N_5372,N_5868);
and U6944 (N_6944,N_5840,N_5740);
or U6945 (N_6945,N_5417,N_4672);
and U6946 (N_6946,N_4919,N_5868);
xor U6947 (N_6947,N_5593,N_4761);
nor U6948 (N_6948,N_4758,N_4500);
or U6949 (N_6949,N_4522,N_5143);
or U6950 (N_6950,N_5788,N_5239);
nor U6951 (N_6951,N_5866,N_4526);
nand U6952 (N_6952,N_5414,N_4537);
xnor U6953 (N_6953,N_5050,N_5236);
xor U6954 (N_6954,N_5053,N_5394);
nand U6955 (N_6955,N_5623,N_4838);
nor U6956 (N_6956,N_4556,N_4985);
and U6957 (N_6957,N_4682,N_5134);
xnor U6958 (N_6958,N_4725,N_5477);
nand U6959 (N_6959,N_4690,N_4907);
or U6960 (N_6960,N_5686,N_5438);
or U6961 (N_6961,N_4506,N_4991);
nor U6962 (N_6962,N_4975,N_5803);
and U6963 (N_6963,N_5554,N_4530);
xor U6964 (N_6964,N_5161,N_5174);
nor U6965 (N_6965,N_5110,N_4726);
xnor U6966 (N_6966,N_5473,N_4582);
nor U6967 (N_6967,N_5699,N_5433);
and U6968 (N_6968,N_5751,N_4630);
nand U6969 (N_6969,N_5967,N_5623);
nand U6970 (N_6970,N_5731,N_5802);
or U6971 (N_6971,N_4763,N_5430);
and U6972 (N_6972,N_5825,N_5532);
and U6973 (N_6973,N_5688,N_5557);
and U6974 (N_6974,N_5902,N_4738);
or U6975 (N_6975,N_4593,N_5860);
xnor U6976 (N_6976,N_5927,N_5664);
xor U6977 (N_6977,N_4791,N_4547);
or U6978 (N_6978,N_4523,N_5044);
and U6979 (N_6979,N_5508,N_5637);
nand U6980 (N_6980,N_4971,N_4637);
and U6981 (N_6981,N_5493,N_5414);
xnor U6982 (N_6982,N_5572,N_4656);
nand U6983 (N_6983,N_5729,N_5920);
nor U6984 (N_6984,N_5967,N_4937);
xnor U6985 (N_6985,N_4852,N_5186);
or U6986 (N_6986,N_5420,N_5544);
and U6987 (N_6987,N_4759,N_5864);
nand U6988 (N_6988,N_5181,N_5129);
nand U6989 (N_6989,N_5465,N_5225);
and U6990 (N_6990,N_5092,N_5082);
nand U6991 (N_6991,N_4920,N_5597);
xnor U6992 (N_6992,N_5974,N_5804);
nand U6993 (N_6993,N_4763,N_5583);
or U6994 (N_6994,N_4623,N_5408);
nor U6995 (N_6995,N_5631,N_5804);
nor U6996 (N_6996,N_5816,N_5111);
xnor U6997 (N_6997,N_4830,N_4745);
nand U6998 (N_6998,N_5572,N_5160);
or U6999 (N_6999,N_5583,N_5006);
nand U7000 (N_7000,N_5124,N_5785);
xor U7001 (N_7001,N_5436,N_5880);
xnor U7002 (N_7002,N_5271,N_5844);
or U7003 (N_7003,N_4707,N_5431);
nor U7004 (N_7004,N_5164,N_5191);
nor U7005 (N_7005,N_5777,N_4674);
and U7006 (N_7006,N_5623,N_5570);
nor U7007 (N_7007,N_5299,N_5418);
nor U7008 (N_7008,N_4549,N_5483);
nand U7009 (N_7009,N_5316,N_5880);
xnor U7010 (N_7010,N_4896,N_5767);
nor U7011 (N_7011,N_4523,N_5657);
nor U7012 (N_7012,N_5591,N_5031);
nand U7013 (N_7013,N_4797,N_4838);
nor U7014 (N_7014,N_5308,N_4786);
xor U7015 (N_7015,N_5651,N_5868);
or U7016 (N_7016,N_5049,N_5102);
nor U7017 (N_7017,N_5279,N_4917);
and U7018 (N_7018,N_5228,N_5201);
xnor U7019 (N_7019,N_5011,N_5849);
nand U7020 (N_7020,N_5204,N_4970);
nand U7021 (N_7021,N_5957,N_5111);
xor U7022 (N_7022,N_5639,N_4531);
or U7023 (N_7023,N_5202,N_5853);
or U7024 (N_7024,N_4724,N_4708);
nor U7025 (N_7025,N_5695,N_5756);
nor U7026 (N_7026,N_5372,N_5933);
nand U7027 (N_7027,N_5972,N_5668);
and U7028 (N_7028,N_5247,N_5343);
xor U7029 (N_7029,N_5713,N_5744);
nand U7030 (N_7030,N_4708,N_5780);
xor U7031 (N_7031,N_4841,N_4569);
or U7032 (N_7032,N_5002,N_5905);
or U7033 (N_7033,N_4965,N_5631);
nand U7034 (N_7034,N_5442,N_5713);
and U7035 (N_7035,N_5815,N_4993);
nand U7036 (N_7036,N_5341,N_5877);
nand U7037 (N_7037,N_5627,N_5959);
nand U7038 (N_7038,N_5437,N_5366);
or U7039 (N_7039,N_4933,N_5691);
nor U7040 (N_7040,N_4965,N_5979);
and U7041 (N_7041,N_5677,N_4668);
and U7042 (N_7042,N_5363,N_4745);
nor U7043 (N_7043,N_5764,N_5370);
nand U7044 (N_7044,N_5346,N_5236);
nor U7045 (N_7045,N_5406,N_4864);
nor U7046 (N_7046,N_5527,N_4749);
xnor U7047 (N_7047,N_5669,N_5636);
nand U7048 (N_7048,N_4826,N_5265);
nor U7049 (N_7049,N_5823,N_5595);
and U7050 (N_7050,N_5711,N_5096);
xor U7051 (N_7051,N_4660,N_5584);
and U7052 (N_7052,N_5118,N_4893);
xor U7053 (N_7053,N_5635,N_4877);
xor U7054 (N_7054,N_5841,N_4749);
xnor U7055 (N_7055,N_5410,N_4600);
xnor U7056 (N_7056,N_5939,N_5737);
or U7057 (N_7057,N_5011,N_5389);
xnor U7058 (N_7058,N_5283,N_5180);
xor U7059 (N_7059,N_4553,N_4522);
nor U7060 (N_7060,N_5159,N_5583);
nand U7061 (N_7061,N_5841,N_4940);
xnor U7062 (N_7062,N_5118,N_5263);
nor U7063 (N_7063,N_5684,N_4714);
or U7064 (N_7064,N_5529,N_5759);
and U7065 (N_7065,N_5081,N_5326);
or U7066 (N_7066,N_5418,N_5629);
nor U7067 (N_7067,N_5000,N_4794);
xnor U7068 (N_7068,N_5068,N_5198);
nand U7069 (N_7069,N_5792,N_4781);
and U7070 (N_7070,N_4715,N_5603);
and U7071 (N_7071,N_5626,N_5213);
xnor U7072 (N_7072,N_4615,N_4654);
nor U7073 (N_7073,N_4848,N_5584);
xor U7074 (N_7074,N_5014,N_5957);
nor U7075 (N_7075,N_4565,N_4972);
or U7076 (N_7076,N_4954,N_5183);
nand U7077 (N_7077,N_5311,N_4540);
nor U7078 (N_7078,N_4820,N_5304);
nand U7079 (N_7079,N_4924,N_5996);
nand U7080 (N_7080,N_5623,N_4947);
nand U7081 (N_7081,N_5484,N_5491);
nor U7082 (N_7082,N_4824,N_5600);
nand U7083 (N_7083,N_4957,N_4580);
and U7084 (N_7084,N_5311,N_4515);
or U7085 (N_7085,N_5174,N_5431);
nand U7086 (N_7086,N_5788,N_5822);
or U7087 (N_7087,N_5502,N_4735);
nand U7088 (N_7088,N_4659,N_4528);
or U7089 (N_7089,N_5959,N_5682);
nor U7090 (N_7090,N_4822,N_4585);
or U7091 (N_7091,N_5462,N_4834);
or U7092 (N_7092,N_5293,N_4661);
or U7093 (N_7093,N_4567,N_4979);
nand U7094 (N_7094,N_5322,N_5743);
or U7095 (N_7095,N_4809,N_5350);
or U7096 (N_7096,N_4554,N_5455);
or U7097 (N_7097,N_4695,N_5336);
nor U7098 (N_7098,N_5228,N_4618);
or U7099 (N_7099,N_5490,N_4522);
and U7100 (N_7100,N_5996,N_4820);
and U7101 (N_7101,N_4531,N_5169);
xor U7102 (N_7102,N_5409,N_5302);
nor U7103 (N_7103,N_5819,N_5475);
xor U7104 (N_7104,N_5232,N_5270);
or U7105 (N_7105,N_5392,N_5936);
nand U7106 (N_7106,N_5023,N_5952);
nand U7107 (N_7107,N_4872,N_4522);
xnor U7108 (N_7108,N_5247,N_5878);
nor U7109 (N_7109,N_5355,N_5795);
and U7110 (N_7110,N_5795,N_5673);
nand U7111 (N_7111,N_5676,N_4937);
xnor U7112 (N_7112,N_5914,N_5265);
or U7113 (N_7113,N_5441,N_5483);
nand U7114 (N_7114,N_5617,N_4909);
nor U7115 (N_7115,N_5261,N_5071);
or U7116 (N_7116,N_5425,N_5787);
and U7117 (N_7117,N_5830,N_5274);
nor U7118 (N_7118,N_5748,N_5026);
and U7119 (N_7119,N_4944,N_4641);
and U7120 (N_7120,N_4939,N_5261);
nand U7121 (N_7121,N_4724,N_5032);
xnor U7122 (N_7122,N_5462,N_5116);
nand U7123 (N_7123,N_4693,N_5405);
and U7124 (N_7124,N_4905,N_4690);
or U7125 (N_7125,N_5401,N_5449);
and U7126 (N_7126,N_5143,N_5215);
and U7127 (N_7127,N_5887,N_4643);
nand U7128 (N_7128,N_5793,N_5856);
xor U7129 (N_7129,N_5602,N_4645);
or U7130 (N_7130,N_5919,N_5178);
xnor U7131 (N_7131,N_5309,N_5534);
nand U7132 (N_7132,N_4959,N_5884);
xor U7133 (N_7133,N_5410,N_5403);
nor U7134 (N_7134,N_5746,N_5093);
nor U7135 (N_7135,N_4918,N_5087);
and U7136 (N_7136,N_5032,N_5436);
and U7137 (N_7137,N_4502,N_4597);
or U7138 (N_7138,N_4551,N_5970);
and U7139 (N_7139,N_4808,N_5642);
xor U7140 (N_7140,N_5723,N_5052);
and U7141 (N_7141,N_5061,N_5534);
nor U7142 (N_7142,N_5916,N_4794);
and U7143 (N_7143,N_5256,N_4519);
nand U7144 (N_7144,N_5727,N_4797);
nand U7145 (N_7145,N_4737,N_5414);
and U7146 (N_7146,N_5643,N_5101);
and U7147 (N_7147,N_5304,N_4553);
or U7148 (N_7148,N_5834,N_5871);
or U7149 (N_7149,N_5513,N_5436);
or U7150 (N_7150,N_5639,N_4817);
or U7151 (N_7151,N_5546,N_4757);
or U7152 (N_7152,N_5267,N_5765);
and U7153 (N_7153,N_5709,N_5921);
nor U7154 (N_7154,N_5709,N_5431);
or U7155 (N_7155,N_5900,N_4642);
nor U7156 (N_7156,N_5210,N_4569);
and U7157 (N_7157,N_5512,N_5758);
nor U7158 (N_7158,N_5168,N_5192);
xnor U7159 (N_7159,N_5271,N_5332);
xnor U7160 (N_7160,N_5522,N_5397);
nor U7161 (N_7161,N_5025,N_5510);
xnor U7162 (N_7162,N_4570,N_5163);
nand U7163 (N_7163,N_5696,N_5057);
nand U7164 (N_7164,N_5118,N_5195);
nand U7165 (N_7165,N_5572,N_5353);
nor U7166 (N_7166,N_5393,N_4862);
xor U7167 (N_7167,N_4910,N_5654);
nand U7168 (N_7168,N_4955,N_5017);
nand U7169 (N_7169,N_5372,N_4645);
or U7170 (N_7170,N_5619,N_4693);
xor U7171 (N_7171,N_5526,N_4640);
and U7172 (N_7172,N_4541,N_5900);
or U7173 (N_7173,N_5122,N_5211);
and U7174 (N_7174,N_5523,N_5071);
xor U7175 (N_7175,N_5952,N_5633);
and U7176 (N_7176,N_4556,N_5245);
and U7177 (N_7177,N_5649,N_5424);
xor U7178 (N_7178,N_5197,N_5226);
nand U7179 (N_7179,N_5976,N_4671);
nor U7180 (N_7180,N_4859,N_4952);
and U7181 (N_7181,N_5185,N_4508);
nand U7182 (N_7182,N_4692,N_4691);
or U7183 (N_7183,N_4928,N_5904);
nand U7184 (N_7184,N_5754,N_5776);
nor U7185 (N_7185,N_5252,N_5105);
xor U7186 (N_7186,N_4921,N_5061);
nand U7187 (N_7187,N_4658,N_4912);
xnor U7188 (N_7188,N_5250,N_5256);
and U7189 (N_7189,N_5312,N_5955);
and U7190 (N_7190,N_5222,N_4834);
xor U7191 (N_7191,N_5005,N_5282);
and U7192 (N_7192,N_5795,N_5233);
nor U7193 (N_7193,N_4738,N_4898);
nand U7194 (N_7194,N_4670,N_5261);
xor U7195 (N_7195,N_5546,N_5804);
nand U7196 (N_7196,N_5115,N_5255);
nand U7197 (N_7197,N_4676,N_4753);
nor U7198 (N_7198,N_4951,N_5029);
nor U7199 (N_7199,N_5872,N_5791);
nand U7200 (N_7200,N_5063,N_5096);
or U7201 (N_7201,N_5836,N_4941);
or U7202 (N_7202,N_5634,N_5668);
nor U7203 (N_7203,N_4637,N_5174);
and U7204 (N_7204,N_4841,N_5621);
and U7205 (N_7205,N_5796,N_5950);
or U7206 (N_7206,N_5964,N_5854);
nor U7207 (N_7207,N_4662,N_5810);
nand U7208 (N_7208,N_5458,N_5528);
or U7209 (N_7209,N_5470,N_5466);
xor U7210 (N_7210,N_5990,N_5575);
nor U7211 (N_7211,N_5761,N_4733);
xor U7212 (N_7212,N_4653,N_4631);
and U7213 (N_7213,N_5732,N_5783);
nor U7214 (N_7214,N_5071,N_5756);
nor U7215 (N_7215,N_5209,N_5897);
and U7216 (N_7216,N_5282,N_4903);
and U7217 (N_7217,N_5580,N_5986);
nand U7218 (N_7218,N_5697,N_4860);
and U7219 (N_7219,N_5330,N_4599);
or U7220 (N_7220,N_5160,N_5624);
xnor U7221 (N_7221,N_5922,N_5758);
nor U7222 (N_7222,N_5289,N_4701);
or U7223 (N_7223,N_5211,N_5687);
xnor U7224 (N_7224,N_5860,N_5809);
xnor U7225 (N_7225,N_4897,N_5975);
and U7226 (N_7226,N_5250,N_5017);
nor U7227 (N_7227,N_4517,N_4837);
nand U7228 (N_7228,N_4890,N_5890);
nor U7229 (N_7229,N_5714,N_5033);
nand U7230 (N_7230,N_4714,N_4528);
nor U7231 (N_7231,N_5977,N_5319);
and U7232 (N_7232,N_5540,N_4629);
or U7233 (N_7233,N_5707,N_5247);
nand U7234 (N_7234,N_4598,N_5501);
nand U7235 (N_7235,N_4763,N_5932);
or U7236 (N_7236,N_5764,N_5075);
xnor U7237 (N_7237,N_5927,N_4554);
nor U7238 (N_7238,N_4693,N_5004);
or U7239 (N_7239,N_5562,N_5843);
nor U7240 (N_7240,N_5329,N_5281);
nor U7241 (N_7241,N_5443,N_5643);
xor U7242 (N_7242,N_5644,N_5831);
nand U7243 (N_7243,N_5088,N_4987);
xor U7244 (N_7244,N_5165,N_5479);
xor U7245 (N_7245,N_5899,N_4829);
xor U7246 (N_7246,N_4590,N_4949);
xor U7247 (N_7247,N_4877,N_5671);
xnor U7248 (N_7248,N_4611,N_5274);
and U7249 (N_7249,N_5111,N_5222);
nor U7250 (N_7250,N_5107,N_5340);
or U7251 (N_7251,N_5493,N_5175);
and U7252 (N_7252,N_4798,N_5773);
and U7253 (N_7253,N_4587,N_5889);
nand U7254 (N_7254,N_5236,N_4821);
nand U7255 (N_7255,N_5515,N_4680);
or U7256 (N_7256,N_5226,N_5073);
or U7257 (N_7257,N_5502,N_5744);
nand U7258 (N_7258,N_4921,N_5377);
nor U7259 (N_7259,N_4587,N_4786);
and U7260 (N_7260,N_5285,N_5300);
nor U7261 (N_7261,N_5918,N_5235);
nor U7262 (N_7262,N_5035,N_5470);
nand U7263 (N_7263,N_5896,N_5232);
or U7264 (N_7264,N_4857,N_5343);
nand U7265 (N_7265,N_4733,N_5693);
or U7266 (N_7266,N_5824,N_4541);
or U7267 (N_7267,N_4806,N_5375);
nor U7268 (N_7268,N_5947,N_5297);
and U7269 (N_7269,N_5816,N_5573);
nor U7270 (N_7270,N_4561,N_5473);
or U7271 (N_7271,N_5147,N_4975);
xor U7272 (N_7272,N_5241,N_5738);
or U7273 (N_7273,N_5609,N_5090);
or U7274 (N_7274,N_5058,N_5605);
nor U7275 (N_7275,N_5126,N_4635);
and U7276 (N_7276,N_4801,N_5356);
nor U7277 (N_7277,N_5113,N_5418);
xnor U7278 (N_7278,N_5499,N_5880);
xor U7279 (N_7279,N_4669,N_5787);
nand U7280 (N_7280,N_5819,N_5438);
nand U7281 (N_7281,N_4730,N_5768);
nor U7282 (N_7282,N_5773,N_4764);
and U7283 (N_7283,N_5469,N_5116);
or U7284 (N_7284,N_5489,N_4842);
xnor U7285 (N_7285,N_5874,N_4620);
and U7286 (N_7286,N_5017,N_4651);
nand U7287 (N_7287,N_5768,N_4687);
or U7288 (N_7288,N_4664,N_5400);
or U7289 (N_7289,N_5046,N_5415);
nand U7290 (N_7290,N_5275,N_5075);
nand U7291 (N_7291,N_5070,N_5689);
and U7292 (N_7292,N_5704,N_4691);
or U7293 (N_7293,N_5930,N_5643);
nand U7294 (N_7294,N_5721,N_5511);
and U7295 (N_7295,N_4948,N_5021);
or U7296 (N_7296,N_5788,N_5856);
nor U7297 (N_7297,N_5495,N_4684);
xnor U7298 (N_7298,N_4845,N_5105);
and U7299 (N_7299,N_4604,N_5121);
and U7300 (N_7300,N_5810,N_4505);
nand U7301 (N_7301,N_4602,N_5824);
nand U7302 (N_7302,N_4603,N_5833);
xnor U7303 (N_7303,N_5125,N_4554);
or U7304 (N_7304,N_4663,N_4783);
nand U7305 (N_7305,N_4566,N_5592);
and U7306 (N_7306,N_5346,N_5511);
xnor U7307 (N_7307,N_5026,N_4513);
xnor U7308 (N_7308,N_4959,N_5010);
or U7309 (N_7309,N_5256,N_4535);
and U7310 (N_7310,N_5317,N_4928);
xnor U7311 (N_7311,N_4892,N_5793);
nor U7312 (N_7312,N_5771,N_5442);
or U7313 (N_7313,N_5808,N_5090);
nand U7314 (N_7314,N_4807,N_4844);
xor U7315 (N_7315,N_5082,N_5821);
nand U7316 (N_7316,N_5464,N_4779);
and U7317 (N_7317,N_4602,N_4799);
and U7318 (N_7318,N_5610,N_5261);
and U7319 (N_7319,N_5511,N_5860);
or U7320 (N_7320,N_5048,N_5400);
xnor U7321 (N_7321,N_5222,N_5900);
xor U7322 (N_7322,N_4976,N_4669);
and U7323 (N_7323,N_4884,N_5349);
nor U7324 (N_7324,N_4748,N_5736);
or U7325 (N_7325,N_5052,N_5397);
xor U7326 (N_7326,N_4811,N_4520);
or U7327 (N_7327,N_5896,N_4555);
and U7328 (N_7328,N_4933,N_5717);
or U7329 (N_7329,N_5023,N_5950);
and U7330 (N_7330,N_5786,N_5518);
and U7331 (N_7331,N_5346,N_5621);
xor U7332 (N_7332,N_4909,N_4812);
nor U7333 (N_7333,N_4775,N_4719);
nand U7334 (N_7334,N_4516,N_4543);
and U7335 (N_7335,N_5374,N_4849);
xnor U7336 (N_7336,N_5589,N_4500);
or U7337 (N_7337,N_5081,N_5747);
nand U7338 (N_7338,N_5522,N_5819);
nor U7339 (N_7339,N_5464,N_5217);
nor U7340 (N_7340,N_5631,N_5486);
nor U7341 (N_7341,N_4700,N_5497);
nor U7342 (N_7342,N_4620,N_5985);
or U7343 (N_7343,N_4561,N_5466);
or U7344 (N_7344,N_5932,N_5519);
nand U7345 (N_7345,N_5836,N_5911);
nor U7346 (N_7346,N_5978,N_5113);
or U7347 (N_7347,N_5267,N_4940);
xor U7348 (N_7348,N_5116,N_5516);
or U7349 (N_7349,N_5095,N_4970);
and U7350 (N_7350,N_5741,N_4581);
and U7351 (N_7351,N_4648,N_5031);
and U7352 (N_7352,N_5913,N_5567);
and U7353 (N_7353,N_4548,N_4830);
and U7354 (N_7354,N_5439,N_4667);
xnor U7355 (N_7355,N_5688,N_4754);
nor U7356 (N_7356,N_5463,N_5831);
nor U7357 (N_7357,N_5964,N_5217);
xor U7358 (N_7358,N_5722,N_4565);
nand U7359 (N_7359,N_5319,N_4766);
or U7360 (N_7360,N_5008,N_4891);
nand U7361 (N_7361,N_5758,N_5491);
and U7362 (N_7362,N_4986,N_5451);
or U7363 (N_7363,N_5369,N_4913);
xor U7364 (N_7364,N_4785,N_4790);
xor U7365 (N_7365,N_5071,N_4919);
or U7366 (N_7366,N_4594,N_4962);
and U7367 (N_7367,N_5555,N_5536);
nor U7368 (N_7368,N_5073,N_5781);
xnor U7369 (N_7369,N_4795,N_5847);
nor U7370 (N_7370,N_5466,N_5261);
xor U7371 (N_7371,N_5778,N_4816);
nor U7372 (N_7372,N_4778,N_4704);
nand U7373 (N_7373,N_5226,N_5359);
xnor U7374 (N_7374,N_5437,N_5360);
nand U7375 (N_7375,N_4598,N_4798);
nor U7376 (N_7376,N_4683,N_5892);
and U7377 (N_7377,N_4979,N_5532);
nand U7378 (N_7378,N_5278,N_5937);
and U7379 (N_7379,N_5894,N_4914);
or U7380 (N_7380,N_4689,N_4961);
or U7381 (N_7381,N_4605,N_5069);
xor U7382 (N_7382,N_4982,N_4592);
nand U7383 (N_7383,N_5447,N_4659);
nand U7384 (N_7384,N_5074,N_5204);
nor U7385 (N_7385,N_4593,N_5103);
or U7386 (N_7386,N_5678,N_4919);
or U7387 (N_7387,N_4693,N_5686);
and U7388 (N_7388,N_4824,N_5324);
nand U7389 (N_7389,N_5185,N_4704);
and U7390 (N_7390,N_5057,N_5516);
nor U7391 (N_7391,N_5385,N_5424);
and U7392 (N_7392,N_4765,N_5284);
or U7393 (N_7393,N_5511,N_5484);
nor U7394 (N_7394,N_5258,N_5408);
nor U7395 (N_7395,N_4656,N_5649);
nor U7396 (N_7396,N_5930,N_5555);
and U7397 (N_7397,N_5667,N_5651);
nand U7398 (N_7398,N_5366,N_5099);
or U7399 (N_7399,N_5909,N_4945);
nor U7400 (N_7400,N_4721,N_5631);
xor U7401 (N_7401,N_4694,N_4884);
xor U7402 (N_7402,N_5636,N_5994);
or U7403 (N_7403,N_4989,N_5818);
nand U7404 (N_7404,N_4916,N_4923);
and U7405 (N_7405,N_5972,N_4905);
xor U7406 (N_7406,N_5730,N_4514);
nand U7407 (N_7407,N_5795,N_5439);
and U7408 (N_7408,N_5210,N_4761);
and U7409 (N_7409,N_4999,N_5727);
or U7410 (N_7410,N_4840,N_4556);
nand U7411 (N_7411,N_4850,N_5502);
nor U7412 (N_7412,N_5829,N_5234);
and U7413 (N_7413,N_5522,N_5161);
or U7414 (N_7414,N_5984,N_5216);
xnor U7415 (N_7415,N_5339,N_5275);
xor U7416 (N_7416,N_5851,N_5408);
nand U7417 (N_7417,N_4810,N_5800);
xnor U7418 (N_7418,N_5328,N_5230);
nand U7419 (N_7419,N_5830,N_4848);
nor U7420 (N_7420,N_5684,N_5473);
and U7421 (N_7421,N_5374,N_5975);
nand U7422 (N_7422,N_4971,N_5051);
and U7423 (N_7423,N_5324,N_5789);
nand U7424 (N_7424,N_5907,N_5301);
nand U7425 (N_7425,N_5788,N_4597);
xor U7426 (N_7426,N_5291,N_5659);
nand U7427 (N_7427,N_5932,N_5216);
nand U7428 (N_7428,N_5854,N_5119);
and U7429 (N_7429,N_4579,N_5838);
xnor U7430 (N_7430,N_5963,N_5177);
xor U7431 (N_7431,N_5529,N_5384);
or U7432 (N_7432,N_4539,N_4906);
nand U7433 (N_7433,N_5444,N_4860);
nand U7434 (N_7434,N_5320,N_5692);
or U7435 (N_7435,N_4625,N_5573);
xor U7436 (N_7436,N_4519,N_5519);
and U7437 (N_7437,N_4710,N_5394);
or U7438 (N_7438,N_5585,N_5822);
or U7439 (N_7439,N_4713,N_5766);
or U7440 (N_7440,N_5744,N_5505);
or U7441 (N_7441,N_4938,N_5084);
nand U7442 (N_7442,N_4621,N_5359);
nand U7443 (N_7443,N_5545,N_5874);
nand U7444 (N_7444,N_5889,N_4520);
and U7445 (N_7445,N_5084,N_5487);
or U7446 (N_7446,N_5230,N_5828);
nor U7447 (N_7447,N_4793,N_4852);
or U7448 (N_7448,N_5793,N_5894);
or U7449 (N_7449,N_5810,N_5938);
or U7450 (N_7450,N_5987,N_5890);
nor U7451 (N_7451,N_4839,N_5551);
and U7452 (N_7452,N_5049,N_5500);
or U7453 (N_7453,N_4696,N_5524);
or U7454 (N_7454,N_4799,N_4511);
nor U7455 (N_7455,N_5304,N_5038);
nand U7456 (N_7456,N_4544,N_4501);
nand U7457 (N_7457,N_5157,N_4746);
nor U7458 (N_7458,N_5388,N_5297);
nand U7459 (N_7459,N_4864,N_4745);
nor U7460 (N_7460,N_5433,N_5730);
or U7461 (N_7461,N_5749,N_5784);
or U7462 (N_7462,N_5949,N_5239);
and U7463 (N_7463,N_5705,N_5473);
xnor U7464 (N_7464,N_5828,N_5467);
or U7465 (N_7465,N_5752,N_4534);
xor U7466 (N_7466,N_5422,N_4599);
or U7467 (N_7467,N_5115,N_4531);
nand U7468 (N_7468,N_4524,N_4949);
and U7469 (N_7469,N_5401,N_5299);
or U7470 (N_7470,N_5954,N_5772);
nand U7471 (N_7471,N_5789,N_5976);
nor U7472 (N_7472,N_5496,N_4860);
nand U7473 (N_7473,N_4839,N_5194);
xor U7474 (N_7474,N_5448,N_4740);
nand U7475 (N_7475,N_5316,N_5683);
or U7476 (N_7476,N_5959,N_5094);
xor U7477 (N_7477,N_5767,N_4899);
and U7478 (N_7478,N_4742,N_5651);
and U7479 (N_7479,N_5911,N_5639);
or U7480 (N_7480,N_5033,N_4599);
nand U7481 (N_7481,N_5565,N_4821);
nand U7482 (N_7482,N_4894,N_5616);
nor U7483 (N_7483,N_4939,N_5011);
or U7484 (N_7484,N_4509,N_5441);
xnor U7485 (N_7485,N_5335,N_5311);
nor U7486 (N_7486,N_5879,N_4690);
and U7487 (N_7487,N_4981,N_4542);
or U7488 (N_7488,N_5858,N_4978);
and U7489 (N_7489,N_5356,N_5047);
nor U7490 (N_7490,N_5090,N_4574);
nand U7491 (N_7491,N_5215,N_5211);
and U7492 (N_7492,N_4618,N_4652);
nand U7493 (N_7493,N_4517,N_5666);
and U7494 (N_7494,N_5925,N_4606);
or U7495 (N_7495,N_5433,N_4606);
nor U7496 (N_7496,N_4691,N_5771);
nand U7497 (N_7497,N_5518,N_5877);
or U7498 (N_7498,N_5343,N_5788);
xnor U7499 (N_7499,N_5574,N_4761);
xnor U7500 (N_7500,N_7308,N_6720);
or U7501 (N_7501,N_7161,N_7395);
nor U7502 (N_7502,N_7438,N_6153);
and U7503 (N_7503,N_7276,N_7297);
nor U7504 (N_7504,N_6840,N_7182);
xnor U7505 (N_7505,N_6570,N_7199);
or U7506 (N_7506,N_6225,N_6557);
or U7507 (N_7507,N_7016,N_6715);
and U7508 (N_7508,N_6055,N_6033);
and U7509 (N_7509,N_7021,N_6109);
and U7510 (N_7510,N_7360,N_6154);
nor U7511 (N_7511,N_7142,N_6969);
nor U7512 (N_7512,N_7460,N_7196);
nand U7513 (N_7513,N_6417,N_7235);
nand U7514 (N_7514,N_7327,N_6408);
nor U7515 (N_7515,N_7126,N_6931);
nand U7516 (N_7516,N_6220,N_6922);
nand U7517 (N_7517,N_6936,N_6519);
and U7518 (N_7518,N_7148,N_7347);
nand U7519 (N_7519,N_6590,N_6444);
nor U7520 (N_7520,N_7452,N_7024);
and U7521 (N_7521,N_6729,N_7004);
or U7522 (N_7522,N_6734,N_7080);
nor U7523 (N_7523,N_6521,N_7001);
xor U7524 (N_7524,N_6064,N_6182);
nand U7525 (N_7525,N_7018,N_6008);
and U7526 (N_7526,N_6722,N_6934);
and U7527 (N_7527,N_7150,N_7417);
nand U7528 (N_7528,N_6372,N_7104);
and U7529 (N_7529,N_6569,N_6834);
nor U7530 (N_7530,N_7495,N_6295);
nor U7531 (N_7531,N_6531,N_6901);
and U7532 (N_7532,N_7408,N_6481);
nand U7533 (N_7533,N_7187,N_7087);
nand U7534 (N_7534,N_6847,N_7026);
nand U7535 (N_7535,N_6938,N_6157);
nor U7536 (N_7536,N_7449,N_6839);
or U7537 (N_7537,N_6761,N_6321);
and U7538 (N_7538,N_6887,N_6204);
and U7539 (N_7539,N_7208,N_7413);
and U7540 (N_7540,N_6130,N_7083);
and U7541 (N_7541,N_6447,N_7227);
nor U7542 (N_7542,N_7479,N_7084);
nand U7543 (N_7543,N_7487,N_6956);
nor U7544 (N_7544,N_7385,N_6616);
nand U7545 (N_7545,N_6899,N_6440);
or U7546 (N_7546,N_6341,N_6981);
nand U7547 (N_7547,N_6017,N_7473);
nor U7548 (N_7548,N_6030,N_7426);
or U7549 (N_7549,N_6515,N_7164);
or U7550 (N_7550,N_7154,N_6169);
or U7551 (N_7551,N_6076,N_6597);
xor U7552 (N_7552,N_6501,N_6875);
xnor U7553 (N_7553,N_6054,N_6402);
and U7554 (N_7554,N_6056,N_6926);
or U7555 (N_7555,N_7040,N_6268);
nand U7556 (N_7556,N_6889,N_6122);
nand U7557 (N_7557,N_7458,N_7318);
nand U7558 (N_7558,N_7422,N_7277);
nor U7559 (N_7559,N_6626,N_6797);
or U7560 (N_7560,N_6993,N_6964);
or U7561 (N_7561,N_6312,N_7488);
nand U7562 (N_7562,N_6439,N_7033);
nand U7563 (N_7563,N_6609,N_6205);
nor U7564 (N_7564,N_6283,N_6310);
xnor U7565 (N_7565,N_7482,N_6207);
xnor U7566 (N_7566,N_7129,N_6959);
xor U7567 (N_7567,N_6093,N_6504);
or U7568 (N_7568,N_6218,N_6472);
xor U7569 (N_7569,N_6343,N_6345);
nand U7570 (N_7570,N_7015,N_7117);
and U7571 (N_7571,N_6459,N_6334);
or U7572 (N_7572,N_6144,N_6335);
or U7573 (N_7573,N_7284,N_6318);
or U7574 (N_7574,N_6413,N_7287);
xnor U7575 (N_7575,N_6599,N_6682);
and U7576 (N_7576,N_6494,N_6355);
nor U7577 (N_7577,N_7290,N_6127);
and U7578 (N_7578,N_6352,N_6025);
nand U7579 (N_7579,N_7313,N_7471);
xnor U7580 (N_7580,N_6111,N_6630);
nor U7581 (N_7581,N_6082,N_7359);
nand U7582 (N_7582,N_7394,N_6685);
and U7583 (N_7583,N_7125,N_7388);
xor U7584 (N_7584,N_6702,N_6537);
nand U7585 (N_7585,N_6019,N_6420);
and U7586 (N_7586,N_6588,N_7207);
xor U7587 (N_7587,N_6237,N_7058);
xor U7588 (N_7588,N_6410,N_6112);
nor U7589 (N_7589,N_7372,N_6824);
or U7590 (N_7590,N_7094,N_6211);
nor U7591 (N_7591,N_6792,N_6699);
xor U7592 (N_7592,N_6893,N_6323);
xnor U7593 (N_7593,N_6652,N_6728);
nand U7594 (N_7594,N_7410,N_6760);
nor U7595 (N_7595,N_6966,N_7044);
nand U7596 (N_7596,N_6006,N_6480);
nand U7597 (N_7597,N_6449,N_6745);
or U7598 (N_7598,N_7442,N_6179);
or U7599 (N_7599,N_6765,N_6581);
xnor U7600 (N_7600,N_6833,N_6843);
nor U7601 (N_7601,N_7332,N_6191);
nor U7602 (N_7602,N_7115,N_7036);
or U7603 (N_7603,N_7305,N_7065);
xor U7604 (N_7604,N_7349,N_7013);
nand U7605 (N_7605,N_6433,N_6261);
xor U7606 (N_7606,N_7401,N_6479);
or U7607 (N_7607,N_6404,N_6914);
nand U7608 (N_7608,N_6687,N_7481);
nor U7609 (N_7609,N_7252,N_6585);
nor U7610 (N_7610,N_6645,N_6276);
nand U7611 (N_7611,N_6443,N_6556);
xor U7612 (N_7612,N_6490,N_6086);
or U7613 (N_7613,N_6864,N_6746);
and U7614 (N_7614,N_7257,N_6102);
xnor U7615 (N_7615,N_7456,N_6083);
and U7616 (N_7616,N_6980,N_7062);
xor U7617 (N_7617,N_6270,N_6770);
nor U7618 (N_7618,N_6520,N_6026);
nand U7619 (N_7619,N_7003,N_6841);
or U7620 (N_7620,N_6983,N_7467);
nor U7621 (N_7621,N_7234,N_7047);
nand U7622 (N_7622,N_6533,N_6041);
or U7623 (N_7623,N_7446,N_6658);
nor U7624 (N_7624,N_7213,N_7111);
nand U7625 (N_7625,N_7402,N_6393);
nor U7626 (N_7626,N_7491,N_6904);
nand U7627 (N_7627,N_6683,N_6976);
nor U7628 (N_7628,N_6452,N_7141);
and U7629 (N_7629,N_7085,N_6793);
xor U7630 (N_7630,N_6613,N_6470);
xor U7631 (N_7631,N_6669,N_6802);
nor U7632 (N_7632,N_7172,N_6484);
or U7633 (N_7633,N_7378,N_6163);
xor U7634 (N_7634,N_6328,N_7170);
nand U7635 (N_7635,N_7093,N_7181);
nor U7636 (N_7636,N_6482,N_6810);
nor U7637 (N_7637,N_7074,N_7399);
and U7638 (N_7638,N_7159,N_6339);
nor U7639 (N_7639,N_6483,N_6231);
xor U7640 (N_7640,N_6394,N_7412);
xnor U7641 (N_7641,N_6693,N_7466);
xor U7642 (N_7642,N_6743,N_6356);
nand U7643 (N_7643,N_6948,N_7464);
xnor U7644 (N_7644,N_7386,N_6527);
nand U7645 (N_7645,N_6861,N_6748);
nor U7646 (N_7646,N_6069,N_6140);
nor U7647 (N_7647,N_7192,N_7043);
nand U7648 (N_7648,N_7379,N_7498);
or U7649 (N_7649,N_6185,N_7225);
and U7650 (N_7650,N_6429,N_7333);
nor U7651 (N_7651,N_6463,N_7310);
and U7652 (N_7652,N_6880,N_7226);
xor U7653 (N_7653,N_6763,N_7162);
or U7654 (N_7654,N_6725,N_6365);
xnor U7655 (N_7655,N_7380,N_6034);
and U7656 (N_7656,N_6233,N_7215);
or U7657 (N_7657,N_6329,N_7353);
nand U7658 (N_7658,N_6274,N_6535);
and U7659 (N_7659,N_6592,N_7485);
nor U7660 (N_7660,N_6621,N_6419);
or U7661 (N_7661,N_6488,N_6364);
nand U7662 (N_7662,N_6955,N_6648);
nor U7663 (N_7663,N_7273,N_6744);
and U7664 (N_7664,N_7060,N_6657);
nor U7665 (N_7665,N_6946,N_6435);
nor U7666 (N_7666,N_6530,N_6037);
and U7667 (N_7667,N_7101,N_6507);
xor U7668 (N_7668,N_6622,N_6039);
xor U7669 (N_7669,N_7262,N_7174);
nand U7670 (N_7670,N_7269,N_6732);
xor U7671 (N_7671,N_7249,N_6892);
nor U7672 (N_7672,N_6116,N_7450);
nor U7673 (N_7673,N_6566,N_6647);
or U7674 (N_7674,N_7191,N_6513);
nor U7675 (N_7675,N_6580,N_6816);
nor U7676 (N_7676,N_6004,N_6099);
and U7677 (N_7677,N_7071,N_6397);
nand U7678 (N_7678,N_6020,N_6304);
and U7679 (N_7679,N_7280,N_6712);
xnor U7680 (N_7680,N_6717,N_6639);
or U7681 (N_7681,N_6053,N_7253);
nor U7682 (N_7682,N_6272,N_6434);
nand U7683 (N_7683,N_7447,N_6060);
nor U7684 (N_7684,N_7418,N_6092);
xnor U7685 (N_7685,N_7492,N_6865);
nor U7686 (N_7686,N_7056,N_6418);
xor U7687 (N_7687,N_6606,N_6442);
nor U7688 (N_7688,N_6921,N_6297);
and U7689 (N_7689,N_7168,N_7274);
xor U7690 (N_7690,N_6263,N_6988);
or U7691 (N_7691,N_7307,N_6758);
nor U7692 (N_7692,N_7270,N_6046);
or U7693 (N_7693,N_7184,N_6300);
or U7694 (N_7694,N_6466,N_6445);
or U7695 (N_7695,N_7392,N_7128);
nor U7696 (N_7696,N_6003,N_6045);
nand U7697 (N_7697,N_6121,N_6947);
nand U7698 (N_7698,N_7326,N_6992);
nand U7699 (N_7699,N_6990,N_6972);
nor U7700 (N_7700,N_7109,N_7254);
nor U7701 (N_7701,N_6259,N_6551);
nand U7702 (N_7702,N_7286,N_7022);
and U7703 (N_7703,N_6219,N_6094);
nand U7704 (N_7704,N_7476,N_7147);
nor U7705 (N_7705,N_6180,N_7434);
nand U7706 (N_7706,N_6097,N_6379);
and U7707 (N_7707,N_7183,N_6273);
and U7708 (N_7708,N_6845,N_6979);
or U7709 (N_7709,N_6361,N_6672);
nand U7710 (N_7710,N_7358,N_6661);
and U7711 (N_7711,N_6511,N_7139);
nand U7712 (N_7712,N_6172,N_6119);
or U7713 (N_7713,N_7362,N_6079);
nand U7714 (N_7714,N_6491,N_7311);
xnor U7715 (N_7715,N_6070,N_6548);
xnor U7716 (N_7716,N_6462,N_6857);
nor U7717 (N_7717,N_7012,N_6787);
or U7718 (N_7718,N_7312,N_6549);
nand U7719 (N_7719,N_6510,N_6898);
or U7720 (N_7720,N_6391,N_6584);
nand U7721 (N_7721,N_6349,N_6662);
or U7722 (N_7722,N_6848,N_6196);
and U7723 (N_7723,N_7376,N_6868);
nand U7724 (N_7724,N_6071,N_6516);
xor U7725 (N_7725,N_6620,N_6677);
and U7726 (N_7726,N_6291,N_6989);
xor U7727 (N_7727,N_6733,N_7251);
or U7728 (N_7728,N_7131,N_6756);
or U7729 (N_7729,N_7403,N_6108);
xor U7730 (N_7730,N_6575,N_7451);
nor U7731 (N_7731,N_7420,N_6784);
or U7732 (N_7732,N_6150,N_6450);
or U7733 (N_7733,N_6598,N_6554);
or U7734 (N_7734,N_7053,N_7266);
nand U7735 (N_7735,N_7335,N_7123);
and U7736 (N_7736,N_7160,N_6636);
or U7737 (N_7737,N_6692,N_6314);
xnor U7738 (N_7738,N_6266,N_6074);
xor U7739 (N_7739,N_6415,N_7389);
and U7740 (N_7740,N_6794,N_7247);
nor U7741 (N_7741,N_6731,N_6186);
nor U7742 (N_7742,N_6115,N_6754);
xnor U7743 (N_7743,N_6505,N_7081);
nand U7744 (N_7744,N_6928,N_6141);
and U7745 (N_7745,N_6573,N_6438);
or U7746 (N_7746,N_6177,N_6529);
xor U7747 (N_7747,N_7223,N_6736);
nand U7748 (N_7748,N_7120,N_6188);
or U7749 (N_7749,N_6867,N_7186);
and U7750 (N_7750,N_7194,N_6080);
nor U7751 (N_7751,N_6776,N_6302);
xnor U7752 (N_7752,N_6941,N_7112);
xor U7753 (N_7753,N_7090,N_6085);
and U7754 (N_7754,N_6212,N_7214);
xnor U7755 (N_7755,N_6555,N_6769);
xnor U7756 (N_7756,N_6713,N_6018);
xnor U7757 (N_7757,N_7334,N_6103);
or U7758 (N_7758,N_7052,N_6945);
or U7759 (N_7759,N_7348,N_6646);
nand U7760 (N_7760,N_6245,N_6807);
nand U7761 (N_7761,N_7441,N_6497);
or U7762 (N_7762,N_6862,N_6674);
xor U7763 (N_7763,N_6468,N_6091);
nand U7764 (N_7764,N_6113,N_7409);
xnor U7765 (N_7765,N_7116,N_7427);
and U7766 (N_7766,N_6759,N_6706);
and U7767 (N_7767,N_7124,N_7055);
xor U7768 (N_7768,N_6105,N_6615);
nand U7769 (N_7769,N_6508,N_7020);
nor U7770 (N_7770,N_6978,N_6000);
nor U7771 (N_7771,N_6721,N_6088);
xnor U7772 (N_7772,N_6289,N_7281);
and U7773 (N_7773,N_6228,N_6471);
nor U7774 (N_7774,N_7231,N_6663);
nor U7775 (N_7775,N_7075,N_6194);
nand U7776 (N_7776,N_6779,N_6160);
or U7777 (N_7777,N_6801,N_7029);
nor U7778 (N_7778,N_7285,N_7007);
or U7779 (N_7779,N_6467,N_6927);
or U7780 (N_7780,N_6458,N_7391);
and U7781 (N_7781,N_7059,N_7390);
xor U7782 (N_7782,N_6738,N_6605);
xor U7783 (N_7783,N_6709,N_6373);
nor U7784 (N_7784,N_7030,N_6991);
nor U7785 (N_7785,N_7237,N_6594);
nor U7786 (N_7786,N_7133,N_6822);
nor U7787 (N_7787,N_6856,N_7398);
nor U7788 (N_7788,N_7204,N_6900);
nand U7789 (N_7789,N_6496,N_6216);
nand U7790 (N_7790,N_7057,N_7099);
and U7791 (N_7791,N_7212,N_6799);
and U7792 (N_7792,N_6998,N_6957);
xor U7793 (N_7793,N_6528,N_6327);
or U7794 (N_7794,N_6142,N_6635);
and U7795 (N_7795,N_7278,N_6072);
xor U7796 (N_7796,N_6457,N_6846);
nor U7797 (N_7797,N_7366,N_7195);
nand U7798 (N_7798,N_7078,N_6961);
nand U7799 (N_7799,N_6021,N_6068);
xnor U7800 (N_7800,N_7175,N_6665);
and U7801 (N_7801,N_6850,N_7341);
and U7802 (N_7802,N_6775,N_7346);
and U7803 (N_7803,N_6308,N_7355);
nand U7804 (N_7804,N_7092,N_6911);
and U7805 (N_7805,N_6412,N_6742);
nand U7806 (N_7806,N_6718,N_6643);
or U7807 (N_7807,N_6971,N_7149);
or U7808 (N_7808,N_6110,N_7282);
xnor U7809 (N_7809,N_6591,N_6509);
or U7810 (N_7810,N_7203,N_7025);
nand U7811 (N_7811,N_6786,N_6939);
xor U7812 (N_7812,N_7069,N_6159);
nor U7813 (N_7813,N_7218,N_6542);
nand U7814 (N_7814,N_7086,N_7365);
nor U7815 (N_7815,N_6724,N_7437);
xnor U7816 (N_7816,N_6896,N_7381);
nand U7817 (N_7817,N_6161,N_7011);
and U7818 (N_7818,N_6705,N_6347);
nor U7819 (N_7819,N_7119,N_7445);
nor U7820 (N_7820,N_7414,N_6368);
xor U7821 (N_7821,N_7045,N_6330);
nor U7822 (N_7822,N_6062,N_7339);
or U7823 (N_7823,N_6271,N_7480);
or U7824 (N_7824,N_6366,N_7054);
nand U7825 (N_7825,N_7260,N_7406);
and U7826 (N_7826,N_6844,N_7009);
or U7827 (N_7827,N_6007,N_7006);
nand U7828 (N_7828,N_6577,N_6886);
nand U7829 (N_7829,N_7302,N_7242);
xor U7830 (N_7830,N_7490,N_6137);
nor U7831 (N_7831,N_6254,N_6132);
xnor U7832 (N_7832,N_7049,N_6708);
nand U7833 (N_7833,N_6280,N_6553);
or U7834 (N_7834,N_6578,N_6106);
xor U7835 (N_7835,N_6168,N_6309);
and U7836 (N_7836,N_6803,N_6319);
nand U7837 (N_7837,N_7136,N_6789);
nand U7838 (N_7838,N_6659,N_6853);
and U7839 (N_7839,N_6156,N_7303);
nand U7840 (N_7840,N_7041,N_7017);
or U7841 (N_7841,N_6096,N_6603);
xor U7842 (N_7842,N_7230,N_6595);
and U7843 (N_7843,N_7072,N_6388);
and U7844 (N_7844,N_6009,N_6649);
or U7845 (N_7845,N_7019,N_7165);
or U7846 (N_7846,N_6197,N_6506);
xnor U7847 (N_7847,N_6162,N_6500);
nor U7848 (N_7848,N_7163,N_6558);
nand U7849 (N_7849,N_7127,N_6485);
and U7850 (N_7850,N_6884,N_6634);
xor U7851 (N_7851,N_6690,N_6827);
nor U7852 (N_7852,N_6820,N_6707);
xor U7853 (N_7853,N_6831,N_6456);
xnor U7854 (N_7854,N_6226,N_6860);
and U7855 (N_7855,N_6910,N_6951);
nand U7856 (N_7856,N_6416,N_6935);
or U7857 (N_7857,N_7363,N_6251);
xnor U7858 (N_7858,N_7298,N_6632);
xnor U7859 (N_7859,N_6066,N_6131);
nor U7860 (N_7860,N_6241,N_6885);
or U7861 (N_7861,N_6781,N_6424);
xor U7862 (N_7862,N_7202,N_6924);
or U7863 (N_7863,N_6027,N_6011);
xor U7864 (N_7864,N_6135,N_6932);
and U7865 (N_7865,N_6664,N_6010);
or U7866 (N_7866,N_6224,N_6384);
nand U7867 (N_7867,N_6267,N_6051);
or U7868 (N_7868,N_7493,N_6158);
nor U7869 (N_7869,N_7336,N_6800);
and U7870 (N_7870,N_7245,N_6842);
and U7871 (N_7871,N_7008,N_6741);
nand U7872 (N_7872,N_7096,N_6200);
and U7873 (N_7873,N_7144,N_7352);
nor U7874 (N_7874,N_7484,N_6689);
and U7875 (N_7875,N_6042,N_7424);
xnor U7876 (N_7876,N_7419,N_6460);
and U7877 (N_7877,N_6777,N_6181);
nor U7878 (N_7878,N_6650,N_6385);
nand U7879 (N_7879,N_6136,N_6340);
xnor U7880 (N_7880,N_6336,N_6063);
and U7881 (N_7881,N_7239,N_6369);
or U7882 (N_7882,N_6532,N_7416);
nand U7883 (N_7883,N_6362,N_7475);
and U7884 (N_7884,N_6735,N_6378);
nand U7885 (N_7885,N_6107,N_7397);
and U7886 (N_7886,N_7156,N_7377);
nor U7887 (N_7887,N_6641,N_6133);
or U7888 (N_7888,N_6696,N_6812);
and U7889 (N_7889,N_7250,N_6829);
nand U7890 (N_7890,N_6453,N_7179);
and U7891 (N_7891,N_6313,N_6399);
or U7892 (N_7892,N_7108,N_6571);
xor U7893 (N_7893,N_6382,N_6075);
or U7894 (N_7894,N_6305,N_7400);
or U7895 (N_7895,N_6644,N_7210);
and U7896 (N_7896,N_7244,N_6240);
xor U7897 (N_7897,N_6975,N_6541);
or U7898 (N_7898,N_6124,N_6944);
and U7899 (N_7899,N_6499,N_6307);
and U7900 (N_7900,N_6432,N_6227);
and U7901 (N_7901,N_6441,N_6201);
and U7902 (N_7902,N_7364,N_6695);
nand U7903 (N_7903,N_7103,N_6123);
xnor U7904 (N_7904,N_6246,N_7288);
or U7905 (N_7905,N_7291,N_7338);
or U7906 (N_7906,N_7197,N_7248);
nand U7907 (N_7907,N_6214,N_6890);
nor U7908 (N_7908,N_6954,N_7264);
xnor U7909 (N_7909,N_7316,N_6286);
and U7910 (N_7910,N_6236,N_6395);
or U7911 (N_7911,N_6038,N_6147);
xor U7912 (N_7912,N_6084,N_6819);
or U7913 (N_7913,N_6611,N_7100);
and U7914 (N_7914,N_7295,N_6299);
xor U7915 (N_7915,N_6474,N_6561);
xor U7916 (N_7916,N_7224,N_6269);
xnor U7917 (N_7917,N_6563,N_6918);
nand U7918 (N_7918,N_6795,N_6916);
or U7919 (N_7919,N_6282,N_6826);
or U7920 (N_7920,N_7387,N_7423);
nor U7921 (N_7921,N_6773,N_6596);
nand U7922 (N_7922,N_7217,N_7048);
xnor U7923 (N_7923,N_6694,N_6492);
nand U7924 (N_7924,N_7206,N_6292);
nand U7925 (N_7925,N_6909,N_6583);
nand U7926 (N_7926,N_6405,N_6680);
nor U7927 (N_7927,N_7299,N_7243);
xor U7928 (N_7928,N_7265,N_7145);
or U7929 (N_7929,N_6406,N_6716);
or U7930 (N_7930,N_7146,N_6970);
nor U7931 (N_7931,N_6077,N_6782);
nor U7932 (N_7932,N_6290,N_6285);
or U7933 (N_7933,N_7216,N_7038);
nand U7934 (N_7934,N_7431,N_6950);
nor U7935 (N_7935,N_7113,N_6919);
xnor U7936 (N_7936,N_7173,N_6755);
and U7937 (N_7937,N_6997,N_6730);
or U7938 (N_7938,N_7035,N_6311);
nor U7939 (N_7939,N_6353,N_6293);
nor U7940 (N_7940,N_6184,N_7283);
or U7941 (N_7941,N_6047,N_6374);
and U7942 (N_7942,N_6170,N_6977);
xnor U7943 (N_7943,N_7494,N_7010);
or U7944 (N_7944,N_6078,N_6148);
or U7945 (N_7945,N_7039,N_6455);
and U7946 (N_7946,N_6915,N_6684);
nor U7947 (N_7947,N_6815,N_7367);
nand U7948 (N_7948,N_6711,N_6747);
nor U7949 (N_7949,N_6331,N_6982);
or U7950 (N_7950,N_6907,N_6655);
nand U7951 (N_7951,N_7324,N_6930);
or U7952 (N_7952,N_6700,N_6344);
xnor U7953 (N_7953,N_6942,N_7351);
or U7954 (N_7954,N_6818,N_7097);
and U7955 (N_7955,N_6891,N_6495);
xnor U7956 (N_7956,N_6346,N_6757);
or U7957 (N_7957,N_6866,N_7110);
nand U7958 (N_7958,N_6015,N_6888);
nor U7959 (N_7959,N_7436,N_7118);
xor U7960 (N_7960,N_6381,N_6489);
or U7961 (N_7961,N_7375,N_7404);
nor U7962 (N_7962,N_6589,N_6572);
nand U7963 (N_7963,N_6475,N_7190);
and U7964 (N_7964,N_7478,N_6849);
nor U7965 (N_7965,N_6704,N_6503);
nand U7966 (N_7966,N_7258,N_6058);
nand U7967 (N_7967,N_6653,N_6436);
nand U7968 (N_7968,N_7465,N_6545);
and U7969 (N_7969,N_6876,N_7371);
xnor U7970 (N_7970,N_7275,N_6143);
and U7971 (N_7971,N_6502,N_6421);
and U7972 (N_7972,N_6806,N_6146);
and U7973 (N_7973,N_6608,N_6973);
xor U7974 (N_7974,N_7105,N_6929);
or U7975 (N_7975,N_6044,N_6524);
and U7976 (N_7976,N_6117,N_6464);
nor U7977 (N_7977,N_6234,N_6823);
or U7978 (N_7978,N_6905,N_6255);
nand U7979 (N_7979,N_6016,N_6199);
nand U7980 (N_7980,N_6306,N_7320);
nor U7981 (N_7981,N_7301,N_7374);
nand U7982 (N_7982,N_6281,N_6768);
nand U7983 (N_7983,N_6118,N_6189);
nand U7984 (N_7984,N_6428,N_6348);
nand U7985 (N_7985,N_7198,N_7153);
and U7986 (N_7986,N_7051,N_6375);
or U7987 (N_7987,N_6873,N_6167);
nor U7988 (N_7988,N_6213,N_7428);
nor U7989 (N_7989,N_7061,N_7463);
and U7990 (N_7990,N_7430,N_6809);
nand U7991 (N_7991,N_6666,N_6656);
nor U7992 (N_7992,N_6534,N_6081);
or U7993 (N_7993,N_6040,N_6943);
nor U7994 (N_7994,N_6567,N_6155);
nor U7995 (N_7995,N_7357,N_6670);
nand U7996 (N_7996,N_7002,N_7241);
and U7997 (N_7997,N_6547,N_6798);
nor U7998 (N_7998,N_6633,N_6574);
xnor U7999 (N_7999,N_6552,N_7455);
or U8000 (N_8000,N_6223,N_6239);
or U8001 (N_8001,N_7477,N_6317);
xor U8002 (N_8002,N_6640,N_7309);
and U8003 (N_8003,N_6923,N_6874);
and U8004 (N_8004,N_7098,N_6073);
xnor U8005 (N_8005,N_6579,N_7279);
xor U8006 (N_8006,N_6012,N_6903);
nand U8007 (N_8007,N_6852,N_6883);
or U8008 (N_8008,N_6740,N_7415);
or U8009 (N_8009,N_7255,N_6427);
nor U8010 (N_8010,N_6618,N_6562);
nor U8011 (N_8011,N_6894,N_6631);
or U8012 (N_8012,N_7201,N_6090);
xor U8013 (N_8013,N_6796,N_7076);
nand U8014 (N_8014,N_6333,N_6139);
xor U8015 (N_8015,N_6023,N_7082);
or U8016 (N_8016,N_6104,N_6933);
and U8017 (N_8017,N_6902,N_7407);
and U8018 (N_8018,N_7356,N_6190);
xnor U8019 (N_8019,N_6560,N_6451);
nand U8020 (N_8020,N_6751,N_6604);
and U8021 (N_8021,N_6376,N_7068);
or U8022 (N_8022,N_7166,N_7188);
xor U8023 (N_8023,N_6908,N_6854);
and U8024 (N_8024,N_7200,N_6029);
and U8025 (N_8025,N_6913,N_7368);
and U8026 (N_8026,N_6243,N_7350);
nand U8027 (N_8027,N_7429,N_6790);
xnor U8028 (N_8028,N_6210,N_6749);
or U8029 (N_8029,N_7369,N_6476);
nand U8030 (N_8030,N_7063,N_6242);
xnor U8031 (N_8031,N_7246,N_6628);
nor U8032 (N_8032,N_7107,N_7384);
nor U8033 (N_8033,N_7178,N_6835);
or U8034 (N_8034,N_6448,N_6357);
and U8035 (N_8035,N_6493,N_6487);
xor U8036 (N_8036,N_6691,N_6454);
nor U8037 (N_8037,N_7222,N_7469);
and U8038 (N_8038,N_7405,N_7411);
nand U8039 (N_8039,N_6230,N_6617);
nor U8040 (N_8040,N_6035,N_6013);
nand U8041 (N_8041,N_6363,N_7292);
and U8042 (N_8042,N_6059,N_6920);
and U8043 (N_8043,N_6296,N_6539);
xor U8044 (N_8044,N_6586,N_6559);
or U8045 (N_8045,N_7180,N_7193);
nor U8046 (N_8046,N_6358,N_6814);
or U8047 (N_8047,N_6968,N_6209);
or U8048 (N_8048,N_6486,N_6171);
nor U8049 (N_8049,N_7177,N_6061);
nor U8050 (N_8050,N_6984,N_6870);
nand U8051 (N_8051,N_6701,N_6667);
nor U8052 (N_8052,N_6249,N_6767);
xnor U8053 (N_8053,N_6514,N_7361);
nand U8054 (N_8054,N_6031,N_7344);
nor U8055 (N_8055,N_6624,N_6838);
nor U8056 (N_8056,N_6260,N_7317);
nor U8057 (N_8057,N_6660,N_6582);
xor U8058 (N_8058,N_6774,N_6593);
nor U8059 (N_8059,N_6540,N_6726);
and U8060 (N_8060,N_6256,N_6825);
xor U8061 (N_8061,N_7483,N_6879);
nor U8062 (N_8062,N_7034,N_6377);
nand U8063 (N_8063,N_6198,N_7042);
nand U8064 (N_8064,N_6710,N_7383);
nand U8065 (N_8065,N_6149,N_6739);
nor U8066 (N_8066,N_6895,N_6791);
or U8067 (N_8067,N_6525,N_6288);
xnor U8068 (N_8068,N_6264,N_7005);
nor U8069 (N_8069,N_7337,N_6762);
nor U8070 (N_8070,N_6203,N_6469);
nand U8071 (N_8071,N_6100,N_7329);
nor U8072 (N_8072,N_6022,N_6477);
xor U8073 (N_8073,N_7102,N_6279);
nor U8074 (N_8074,N_6278,N_6817);
and U8075 (N_8075,N_7014,N_6536);
xor U8076 (N_8076,N_7114,N_6859);
or U8077 (N_8077,N_6252,N_7238);
nand U8078 (N_8078,N_6052,N_6005);
nor U8079 (N_8079,N_7176,N_6778);
or U8080 (N_8080,N_7454,N_6565);
and U8081 (N_8081,N_6937,N_7256);
and U8082 (N_8082,N_6287,N_7158);
nor U8083 (N_8083,N_6996,N_6550);
and U8084 (N_8084,N_6303,N_7468);
xnor U8085 (N_8085,N_6804,N_7421);
or U8086 (N_8086,N_7221,N_6813);
nand U8087 (N_8087,N_6960,N_7157);
nor U8088 (N_8088,N_6095,N_7137);
and U8089 (N_8089,N_6262,N_7220);
and U8090 (N_8090,N_7122,N_6325);
nor U8091 (N_8091,N_7240,N_6120);
nor U8092 (N_8092,N_6967,N_6863);
nand U8093 (N_8093,N_6320,N_6350);
or U8094 (N_8094,N_6673,N_6949);
and U8095 (N_8095,N_6002,N_6686);
nand U8096 (N_8096,N_6067,N_6430);
and U8097 (N_8097,N_6380,N_6473);
nor U8098 (N_8098,N_6805,N_7304);
nor U8099 (N_8099,N_6192,N_6940);
nand U8100 (N_8100,N_6587,N_7343);
nor U8101 (N_8101,N_7070,N_7219);
nor U8102 (N_8102,N_6265,N_6994);
nor U8103 (N_8103,N_7433,N_7228);
or U8104 (N_8104,N_6257,N_7046);
nor U8105 (N_8105,N_7095,N_6294);
or U8106 (N_8106,N_6221,N_6087);
or U8107 (N_8107,N_6342,N_6963);
nor U8108 (N_8108,N_6275,N_6881);
xnor U8109 (N_8109,N_7268,N_7314);
or U8110 (N_8110,N_6028,N_7306);
and U8111 (N_8111,N_6187,N_6411);
nand U8112 (N_8112,N_6750,N_6912);
xnor U8113 (N_8113,N_6953,N_6166);
nand U8114 (N_8114,N_6396,N_6478);
nand U8115 (N_8115,N_7031,N_7067);
nand U8116 (N_8116,N_6089,N_7342);
xor U8117 (N_8117,N_6987,N_6174);
or U8118 (N_8118,N_6877,N_6165);
nor U8119 (N_8119,N_6431,N_7461);
nand U8120 (N_8120,N_6629,N_6195);
and U8121 (N_8121,N_6414,N_7382);
and U8122 (N_8122,N_6830,N_6316);
or U8123 (N_8123,N_7396,N_7300);
and U8124 (N_8124,N_7271,N_6235);
and U8125 (N_8125,N_6858,N_6422);
nor U8126 (N_8126,N_7232,N_6101);
xnor U8127 (N_8127,N_6678,N_6371);
nor U8128 (N_8128,N_7089,N_6851);
nand U8129 (N_8129,N_6679,N_6498);
nor U8130 (N_8130,N_6871,N_6383);
and U8131 (N_8131,N_7340,N_7106);
and U8132 (N_8132,N_6049,N_6518);
and U8133 (N_8133,N_7435,N_6129);
nand U8134 (N_8134,N_7259,N_6229);
or U8135 (N_8135,N_7189,N_6952);
xnor U8136 (N_8136,N_6783,N_6248);
nor U8137 (N_8137,N_7135,N_6370);
nand U8138 (N_8138,N_6727,N_6390);
xnor U8139 (N_8139,N_6619,N_7037);
nand U8140 (N_8140,N_6523,N_6392);
or U8141 (N_8141,N_6036,N_7140);
and U8142 (N_8142,N_7079,N_7211);
or U8143 (N_8143,N_7272,N_6389);
and U8144 (N_8144,N_6753,N_7151);
or U8145 (N_8145,N_6788,N_6564);
nor U8146 (N_8146,N_7321,N_6401);
or U8147 (N_8147,N_6164,N_6176);
or U8148 (N_8148,N_6723,N_6138);
nor U8149 (N_8149,N_6151,N_7233);
nor U8150 (N_8150,N_6917,N_6232);
and U8151 (N_8151,N_7354,N_6681);
nor U8152 (N_8152,N_6050,N_6437);
xor U8153 (N_8153,N_6367,N_6752);
xnor U8154 (N_8154,N_7432,N_6821);
and U8155 (N_8155,N_7064,N_6298);
nand U8156 (N_8156,N_7294,N_6425);
xor U8157 (N_8157,N_6676,N_6697);
and U8158 (N_8158,N_6654,N_6772);
xnor U8159 (N_8159,N_7073,N_6057);
nor U8160 (N_8160,N_7066,N_6247);
or U8161 (N_8161,N_6522,N_6882);
nand U8162 (N_8162,N_7489,N_7229);
nand U8163 (N_8163,N_6222,N_7050);
nand U8164 (N_8164,N_6145,N_7132);
and U8165 (N_8165,N_6543,N_6398);
nand U8166 (N_8166,N_7143,N_7373);
or U8167 (N_8167,N_7023,N_7032);
or U8168 (N_8168,N_7263,N_7499);
nor U8169 (N_8169,N_6134,N_6600);
nand U8170 (N_8170,N_6359,N_6576);
and U8171 (N_8171,N_6301,N_6128);
and U8172 (N_8172,N_6001,N_6703);
and U8173 (N_8173,N_6627,N_7027);
and U8174 (N_8174,N_7496,N_7088);
and U8175 (N_8175,N_6360,N_6836);
nand U8176 (N_8176,N_6766,N_6958);
xor U8177 (N_8177,N_6526,N_6737);
nand U8178 (N_8178,N_7459,N_6173);
or U8179 (N_8179,N_7319,N_6183);
nor U8180 (N_8180,N_6354,N_7185);
nor U8181 (N_8181,N_6869,N_6671);
and U8182 (N_8182,N_6178,N_7443);
or U8183 (N_8183,N_6771,N_6668);
and U8184 (N_8184,N_6446,N_6546);
nor U8185 (N_8185,N_6014,N_7331);
nor U8186 (N_8186,N_7028,N_6337);
xor U8187 (N_8187,N_6811,N_7444);
or U8188 (N_8188,N_6322,N_6625);
and U8189 (N_8189,N_6675,N_6878);
and U8190 (N_8190,N_6872,N_7315);
and U8191 (N_8191,N_7289,N_6400);
or U8192 (N_8192,N_7448,N_6193);
nand U8193 (N_8193,N_7472,N_7322);
nor U8194 (N_8194,N_6065,N_6244);
nand U8195 (N_8195,N_6152,N_6785);
and U8196 (N_8196,N_7370,N_7462);
and U8197 (N_8197,N_6423,N_6607);
xor U8198 (N_8198,N_6126,N_6517);
and U8199 (N_8199,N_6217,N_7077);
nor U8200 (N_8200,N_6326,N_6828);
nand U8201 (N_8201,N_6642,N_7000);
nor U8202 (N_8202,N_6403,N_6538);
and U8203 (N_8203,N_6610,N_6215);
nor U8204 (N_8204,N_7293,N_7167);
or U8205 (N_8205,N_6461,N_6614);
xnor U8206 (N_8206,N_6208,N_7091);
xor U8207 (N_8207,N_6985,N_6258);
xnor U8208 (N_8208,N_6602,N_6999);
nor U8209 (N_8209,N_6324,N_7236);
or U8210 (N_8210,N_7209,N_7169);
xnor U8211 (N_8211,N_6426,N_6284);
nor U8212 (N_8212,N_7439,N_6043);
xnor U8213 (N_8213,N_7205,N_7393);
or U8214 (N_8214,N_6780,N_6253);
or U8215 (N_8215,N_6048,N_6544);
or U8216 (N_8216,N_6638,N_6277);
xor U8217 (N_8217,N_6568,N_6719);
nor U8218 (N_8218,N_7323,N_6986);
xnor U8219 (N_8219,N_6808,N_6925);
nor U8220 (N_8220,N_7134,N_6698);
nand U8221 (N_8221,N_6338,N_6206);
nand U8222 (N_8222,N_6837,N_6651);
and U8223 (N_8223,N_7457,N_7121);
and U8224 (N_8224,N_7296,N_6906);
or U8225 (N_8225,N_7497,N_6315);
or U8226 (N_8226,N_6688,N_6202);
nand U8227 (N_8227,N_7267,N_7152);
nor U8228 (N_8228,N_6637,N_6601);
nand U8229 (N_8229,N_6832,N_6962);
or U8230 (N_8230,N_6855,N_7138);
and U8231 (N_8231,N_7345,N_7325);
nand U8232 (N_8232,N_6114,N_6386);
or U8233 (N_8233,N_7330,N_6764);
nor U8234 (N_8234,N_6512,N_7155);
nor U8235 (N_8235,N_6332,N_6238);
and U8236 (N_8236,N_6965,N_6974);
or U8237 (N_8237,N_6387,N_7474);
and U8238 (N_8238,N_6995,N_7440);
and U8239 (N_8239,N_7171,N_6175);
nand U8240 (N_8240,N_7453,N_6351);
xor U8241 (N_8241,N_6465,N_7328);
or U8242 (N_8242,N_6024,N_6714);
or U8243 (N_8243,N_6409,N_6612);
nand U8244 (N_8244,N_6623,N_7470);
nand U8245 (N_8245,N_6125,N_7261);
nand U8246 (N_8246,N_6897,N_6098);
nor U8247 (N_8247,N_6407,N_7425);
nor U8248 (N_8248,N_6032,N_7486);
and U8249 (N_8249,N_7130,N_6250);
nor U8250 (N_8250,N_6576,N_6622);
nand U8251 (N_8251,N_6454,N_7402);
nor U8252 (N_8252,N_7455,N_7386);
and U8253 (N_8253,N_6062,N_7365);
or U8254 (N_8254,N_7323,N_7396);
nor U8255 (N_8255,N_7332,N_7273);
and U8256 (N_8256,N_6175,N_6326);
nand U8257 (N_8257,N_6716,N_6399);
xor U8258 (N_8258,N_7343,N_7311);
xnor U8259 (N_8259,N_6050,N_6252);
or U8260 (N_8260,N_7220,N_6886);
nor U8261 (N_8261,N_7467,N_6415);
nand U8262 (N_8262,N_6441,N_6394);
nand U8263 (N_8263,N_6208,N_6297);
xnor U8264 (N_8264,N_6966,N_7217);
nand U8265 (N_8265,N_6950,N_6040);
nor U8266 (N_8266,N_6120,N_7407);
nand U8267 (N_8267,N_6801,N_7489);
and U8268 (N_8268,N_7402,N_6323);
nor U8269 (N_8269,N_6347,N_6498);
nand U8270 (N_8270,N_7368,N_6753);
or U8271 (N_8271,N_6612,N_6839);
or U8272 (N_8272,N_6674,N_6555);
or U8273 (N_8273,N_6187,N_7026);
xor U8274 (N_8274,N_6949,N_6460);
xor U8275 (N_8275,N_7435,N_7402);
or U8276 (N_8276,N_6372,N_6029);
xnor U8277 (N_8277,N_6706,N_6029);
xnor U8278 (N_8278,N_7189,N_7376);
xor U8279 (N_8279,N_6743,N_6239);
xor U8280 (N_8280,N_6525,N_6939);
and U8281 (N_8281,N_6322,N_6373);
nor U8282 (N_8282,N_6336,N_7419);
xnor U8283 (N_8283,N_6182,N_6514);
or U8284 (N_8284,N_6813,N_6029);
xnor U8285 (N_8285,N_6570,N_6394);
nand U8286 (N_8286,N_7337,N_6929);
nor U8287 (N_8287,N_7232,N_6924);
or U8288 (N_8288,N_7126,N_7476);
nand U8289 (N_8289,N_6263,N_7131);
nor U8290 (N_8290,N_6150,N_7419);
nor U8291 (N_8291,N_6046,N_6368);
and U8292 (N_8292,N_6794,N_6516);
xnor U8293 (N_8293,N_6732,N_6876);
nand U8294 (N_8294,N_6100,N_6167);
xnor U8295 (N_8295,N_6038,N_6701);
nand U8296 (N_8296,N_6472,N_6795);
nand U8297 (N_8297,N_6168,N_7366);
xnor U8298 (N_8298,N_7165,N_6014);
and U8299 (N_8299,N_7076,N_7248);
nand U8300 (N_8300,N_6311,N_6074);
and U8301 (N_8301,N_7363,N_7058);
and U8302 (N_8302,N_7286,N_6619);
nor U8303 (N_8303,N_6003,N_6533);
nor U8304 (N_8304,N_6347,N_6453);
nand U8305 (N_8305,N_7165,N_6472);
and U8306 (N_8306,N_6211,N_6942);
or U8307 (N_8307,N_7047,N_6208);
nand U8308 (N_8308,N_7475,N_6257);
and U8309 (N_8309,N_6689,N_6336);
nand U8310 (N_8310,N_6698,N_6393);
nor U8311 (N_8311,N_7211,N_6460);
and U8312 (N_8312,N_6346,N_6761);
nand U8313 (N_8313,N_7430,N_7288);
or U8314 (N_8314,N_7217,N_7253);
xnor U8315 (N_8315,N_6728,N_7230);
nand U8316 (N_8316,N_6908,N_7256);
nor U8317 (N_8317,N_6190,N_7292);
and U8318 (N_8318,N_7080,N_6399);
nor U8319 (N_8319,N_6045,N_6238);
nand U8320 (N_8320,N_6327,N_6416);
nand U8321 (N_8321,N_6834,N_6590);
xnor U8322 (N_8322,N_6663,N_6701);
or U8323 (N_8323,N_6655,N_7454);
nand U8324 (N_8324,N_6890,N_6346);
nand U8325 (N_8325,N_6794,N_7470);
nand U8326 (N_8326,N_6282,N_6038);
and U8327 (N_8327,N_6538,N_6456);
xnor U8328 (N_8328,N_7142,N_6683);
or U8329 (N_8329,N_6874,N_6618);
or U8330 (N_8330,N_6692,N_6468);
nor U8331 (N_8331,N_7303,N_7295);
and U8332 (N_8332,N_6120,N_6775);
nand U8333 (N_8333,N_6442,N_6699);
nor U8334 (N_8334,N_6243,N_7302);
nand U8335 (N_8335,N_7021,N_6257);
and U8336 (N_8336,N_7464,N_7236);
nand U8337 (N_8337,N_6011,N_6720);
nand U8338 (N_8338,N_6927,N_6100);
nor U8339 (N_8339,N_6189,N_6138);
nand U8340 (N_8340,N_6917,N_6220);
xor U8341 (N_8341,N_6005,N_6354);
or U8342 (N_8342,N_6588,N_6718);
or U8343 (N_8343,N_7038,N_6317);
nand U8344 (N_8344,N_7267,N_6694);
nand U8345 (N_8345,N_6362,N_6657);
nor U8346 (N_8346,N_6736,N_6967);
nor U8347 (N_8347,N_7473,N_6443);
nand U8348 (N_8348,N_6804,N_6899);
and U8349 (N_8349,N_6145,N_6488);
and U8350 (N_8350,N_7259,N_6162);
nor U8351 (N_8351,N_6650,N_6706);
or U8352 (N_8352,N_7307,N_6225);
nand U8353 (N_8353,N_6152,N_7128);
and U8354 (N_8354,N_7045,N_6235);
or U8355 (N_8355,N_6322,N_6788);
and U8356 (N_8356,N_6719,N_6119);
xor U8357 (N_8357,N_6156,N_6074);
nor U8358 (N_8358,N_6362,N_6006);
and U8359 (N_8359,N_6017,N_6703);
and U8360 (N_8360,N_6443,N_6907);
or U8361 (N_8361,N_7253,N_6012);
nand U8362 (N_8362,N_7135,N_6737);
nor U8363 (N_8363,N_6775,N_6149);
xor U8364 (N_8364,N_6529,N_6908);
nor U8365 (N_8365,N_6299,N_6652);
and U8366 (N_8366,N_6839,N_6680);
xnor U8367 (N_8367,N_6558,N_6862);
and U8368 (N_8368,N_7079,N_7408);
nor U8369 (N_8369,N_7007,N_6046);
xnor U8370 (N_8370,N_6931,N_6614);
and U8371 (N_8371,N_7411,N_6652);
xor U8372 (N_8372,N_6552,N_6514);
nor U8373 (N_8373,N_7214,N_6709);
xor U8374 (N_8374,N_6158,N_7478);
xor U8375 (N_8375,N_6226,N_7126);
nor U8376 (N_8376,N_6246,N_7374);
xor U8377 (N_8377,N_6066,N_6054);
and U8378 (N_8378,N_6300,N_6688);
nor U8379 (N_8379,N_6511,N_6958);
nor U8380 (N_8380,N_6029,N_6340);
xor U8381 (N_8381,N_6556,N_7090);
nor U8382 (N_8382,N_6247,N_6710);
xor U8383 (N_8383,N_7480,N_6539);
xnor U8384 (N_8384,N_7283,N_6347);
nand U8385 (N_8385,N_7368,N_7152);
xor U8386 (N_8386,N_6088,N_7046);
xor U8387 (N_8387,N_7293,N_6646);
nor U8388 (N_8388,N_7293,N_7407);
xnor U8389 (N_8389,N_6052,N_6461);
nor U8390 (N_8390,N_6720,N_6123);
and U8391 (N_8391,N_7100,N_6627);
nor U8392 (N_8392,N_6599,N_7341);
nor U8393 (N_8393,N_6308,N_6987);
or U8394 (N_8394,N_6921,N_6829);
or U8395 (N_8395,N_6465,N_6994);
and U8396 (N_8396,N_6409,N_6009);
or U8397 (N_8397,N_6400,N_7361);
or U8398 (N_8398,N_7241,N_7061);
nor U8399 (N_8399,N_6293,N_7332);
nand U8400 (N_8400,N_6853,N_6924);
xnor U8401 (N_8401,N_6218,N_6383);
and U8402 (N_8402,N_6865,N_6349);
xnor U8403 (N_8403,N_7066,N_7463);
nor U8404 (N_8404,N_6497,N_7033);
or U8405 (N_8405,N_6941,N_7404);
nand U8406 (N_8406,N_6965,N_6739);
xnor U8407 (N_8407,N_6008,N_6124);
xnor U8408 (N_8408,N_6423,N_7088);
or U8409 (N_8409,N_6293,N_6284);
nor U8410 (N_8410,N_7254,N_7280);
or U8411 (N_8411,N_6084,N_6360);
xor U8412 (N_8412,N_7390,N_7222);
nand U8413 (N_8413,N_6433,N_7100);
and U8414 (N_8414,N_7029,N_6141);
xnor U8415 (N_8415,N_7254,N_6520);
nor U8416 (N_8416,N_7154,N_7062);
xor U8417 (N_8417,N_6526,N_6576);
nand U8418 (N_8418,N_7094,N_7091);
nand U8419 (N_8419,N_7257,N_6370);
nor U8420 (N_8420,N_6795,N_6419);
nand U8421 (N_8421,N_7076,N_7172);
xor U8422 (N_8422,N_6295,N_6805);
xnor U8423 (N_8423,N_6061,N_7328);
xnor U8424 (N_8424,N_6661,N_7180);
and U8425 (N_8425,N_7450,N_6427);
and U8426 (N_8426,N_6556,N_7440);
or U8427 (N_8427,N_6925,N_6930);
and U8428 (N_8428,N_7400,N_6733);
nor U8429 (N_8429,N_7360,N_7128);
and U8430 (N_8430,N_7169,N_6138);
nand U8431 (N_8431,N_7004,N_6248);
xor U8432 (N_8432,N_7395,N_7184);
or U8433 (N_8433,N_6689,N_6189);
or U8434 (N_8434,N_6154,N_6110);
or U8435 (N_8435,N_6244,N_6469);
and U8436 (N_8436,N_6457,N_6026);
and U8437 (N_8437,N_6875,N_7123);
and U8438 (N_8438,N_6730,N_7313);
nand U8439 (N_8439,N_7002,N_7174);
and U8440 (N_8440,N_6040,N_6678);
nand U8441 (N_8441,N_7175,N_7106);
or U8442 (N_8442,N_7360,N_6022);
and U8443 (N_8443,N_6872,N_7150);
xnor U8444 (N_8444,N_6336,N_6371);
and U8445 (N_8445,N_7147,N_6496);
and U8446 (N_8446,N_6276,N_6066);
xor U8447 (N_8447,N_6258,N_7031);
and U8448 (N_8448,N_6818,N_7299);
or U8449 (N_8449,N_7336,N_6924);
and U8450 (N_8450,N_7133,N_7063);
xor U8451 (N_8451,N_6440,N_7216);
or U8452 (N_8452,N_6197,N_6802);
or U8453 (N_8453,N_6683,N_6382);
and U8454 (N_8454,N_6850,N_6751);
nor U8455 (N_8455,N_6472,N_6097);
nand U8456 (N_8456,N_7401,N_7263);
nor U8457 (N_8457,N_6218,N_7182);
and U8458 (N_8458,N_6396,N_7027);
or U8459 (N_8459,N_6531,N_7371);
nor U8460 (N_8460,N_6268,N_6928);
or U8461 (N_8461,N_6889,N_6399);
nor U8462 (N_8462,N_7273,N_6156);
nor U8463 (N_8463,N_7173,N_7350);
and U8464 (N_8464,N_6380,N_6409);
nor U8465 (N_8465,N_6871,N_7414);
nand U8466 (N_8466,N_7139,N_6236);
nor U8467 (N_8467,N_6796,N_6504);
or U8468 (N_8468,N_6602,N_6659);
xnor U8469 (N_8469,N_6923,N_6527);
or U8470 (N_8470,N_6335,N_6042);
or U8471 (N_8471,N_7287,N_6352);
and U8472 (N_8472,N_6783,N_7301);
xor U8473 (N_8473,N_6541,N_6629);
xnor U8474 (N_8474,N_6788,N_7186);
and U8475 (N_8475,N_7257,N_7412);
nand U8476 (N_8476,N_6525,N_7244);
or U8477 (N_8477,N_7084,N_7331);
xor U8478 (N_8478,N_7212,N_6464);
or U8479 (N_8479,N_7112,N_6381);
nor U8480 (N_8480,N_6159,N_6266);
xnor U8481 (N_8481,N_6751,N_7151);
nand U8482 (N_8482,N_7448,N_7225);
nor U8483 (N_8483,N_6020,N_6255);
nand U8484 (N_8484,N_7342,N_6420);
nand U8485 (N_8485,N_6457,N_6005);
nand U8486 (N_8486,N_7264,N_6379);
and U8487 (N_8487,N_7057,N_7239);
or U8488 (N_8488,N_7130,N_6536);
xor U8489 (N_8489,N_6359,N_7491);
xor U8490 (N_8490,N_6300,N_6548);
or U8491 (N_8491,N_6803,N_7360);
or U8492 (N_8492,N_6098,N_7151);
nand U8493 (N_8493,N_6046,N_6167);
nor U8494 (N_8494,N_6332,N_6826);
nand U8495 (N_8495,N_6528,N_6250);
and U8496 (N_8496,N_6237,N_6074);
nor U8497 (N_8497,N_7427,N_6249);
and U8498 (N_8498,N_6169,N_6088);
nand U8499 (N_8499,N_6615,N_6833);
xnor U8500 (N_8500,N_6716,N_6664);
xnor U8501 (N_8501,N_7191,N_6784);
or U8502 (N_8502,N_7030,N_7004);
nor U8503 (N_8503,N_6910,N_7304);
nor U8504 (N_8504,N_7106,N_6689);
and U8505 (N_8505,N_6886,N_6139);
nor U8506 (N_8506,N_6417,N_7173);
xnor U8507 (N_8507,N_6503,N_6594);
or U8508 (N_8508,N_6993,N_6221);
and U8509 (N_8509,N_6606,N_6243);
xnor U8510 (N_8510,N_7292,N_7171);
nand U8511 (N_8511,N_6126,N_6661);
and U8512 (N_8512,N_6386,N_6075);
or U8513 (N_8513,N_6714,N_6368);
and U8514 (N_8514,N_6210,N_6863);
xor U8515 (N_8515,N_6383,N_6864);
and U8516 (N_8516,N_6205,N_6505);
and U8517 (N_8517,N_6554,N_6486);
nor U8518 (N_8518,N_7431,N_6417);
or U8519 (N_8519,N_7189,N_6328);
and U8520 (N_8520,N_6216,N_6954);
xor U8521 (N_8521,N_6595,N_6756);
or U8522 (N_8522,N_7000,N_7034);
nand U8523 (N_8523,N_6327,N_6760);
and U8524 (N_8524,N_6232,N_6805);
nor U8525 (N_8525,N_6028,N_6330);
xnor U8526 (N_8526,N_7430,N_7074);
nor U8527 (N_8527,N_6270,N_6338);
and U8528 (N_8528,N_7497,N_6931);
and U8529 (N_8529,N_6004,N_7420);
nand U8530 (N_8530,N_7383,N_7341);
xor U8531 (N_8531,N_7052,N_6539);
nor U8532 (N_8532,N_7448,N_6779);
or U8533 (N_8533,N_7437,N_7415);
nor U8534 (N_8534,N_6682,N_6337);
nand U8535 (N_8535,N_7413,N_7264);
nor U8536 (N_8536,N_6080,N_6046);
or U8537 (N_8537,N_7090,N_6246);
or U8538 (N_8538,N_6079,N_6851);
nand U8539 (N_8539,N_6841,N_7371);
nor U8540 (N_8540,N_6187,N_6785);
nor U8541 (N_8541,N_6537,N_6848);
xor U8542 (N_8542,N_7122,N_6928);
xor U8543 (N_8543,N_6141,N_7051);
xnor U8544 (N_8544,N_7219,N_7064);
nor U8545 (N_8545,N_6225,N_6466);
and U8546 (N_8546,N_6630,N_7143);
and U8547 (N_8547,N_6979,N_6761);
and U8548 (N_8548,N_6770,N_6034);
nand U8549 (N_8549,N_7070,N_6937);
nand U8550 (N_8550,N_6389,N_6341);
nor U8551 (N_8551,N_6043,N_6351);
nor U8552 (N_8552,N_7200,N_6230);
or U8553 (N_8553,N_6764,N_6925);
nand U8554 (N_8554,N_7075,N_7009);
nor U8555 (N_8555,N_7419,N_6419);
nand U8556 (N_8556,N_6709,N_6782);
or U8557 (N_8557,N_6017,N_6627);
nor U8558 (N_8558,N_6071,N_6419);
nor U8559 (N_8559,N_6718,N_6903);
xnor U8560 (N_8560,N_7482,N_6872);
or U8561 (N_8561,N_6050,N_6859);
nor U8562 (N_8562,N_6728,N_6861);
nor U8563 (N_8563,N_6750,N_6097);
and U8564 (N_8564,N_6498,N_6613);
xor U8565 (N_8565,N_7089,N_6384);
nor U8566 (N_8566,N_6309,N_6634);
xor U8567 (N_8567,N_6949,N_7478);
xnor U8568 (N_8568,N_6436,N_7071);
xnor U8569 (N_8569,N_6345,N_7343);
nor U8570 (N_8570,N_7246,N_6620);
nand U8571 (N_8571,N_6894,N_7028);
or U8572 (N_8572,N_6090,N_6758);
and U8573 (N_8573,N_7133,N_6682);
or U8574 (N_8574,N_6098,N_6087);
nand U8575 (N_8575,N_7043,N_6322);
nor U8576 (N_8576,N_6062,N_7399);
and U8577 (N_8577,N_6479,N_6649);
xnor U8578 (N_8578,N_7173,N_6360);
or U8579 (N_8579,N_6400,N_7155);
and U8580 (N_8580,N_7329,N_6696);
or U8581 (N_8581,N_7077,N_6767);
or U8582 (N_8582,N_6155,N_6238);
and U8583 (N_8583,N_6095,N_7273);
xnor U8584 (N_8584,N_7119,N_7474);
nor U8585 (N_8585,N_6114,N_6552);
and U8586 (N_8586,N_6380,N_6589);
xor U8587 (N_8587,N_7141,N_6577);
nand U8588 (N_8588,N_6113,N_7261);
and U8589 (N_8589,N_6839,N_6123);
or U8590 (N_8590,N_7222,N_6307);
and U8591 (N_8591,N_7252,N_6955);
or U8592 (N_8592,N_7184,N_6640);
and U8593 (N_8593,N_7329,N_6312);
nor U8594 (N_8594,N_6754,N_7386);
nor U8595 (N_8595,N_6132,N_6758);
and U8596 (N_8596,N_6096,N_6551);
nor U8597 (N_8597,N_6615,N_7092);
or U8598 (N_8598,N_7082,N_6074);
and U8599 (N_8599,N_7427,N_6463);
nand U8600 (N_8600,N_7131,N_7443);
nor U8601 (N_8601,N_6361,N_7383);
nand U8602 (N_8602,N_7354,N_7330);
nor U8603 (N_8603,N_6135,N_6737);
xor U8604 (N_8604,N_6240,N_6903);
nand U8605 (N_8605,N_7342,N_6211);
or U8606 (N_8606,N_6080,N_7345);
or U8607 (N_8607,N_6324,N_7227);
nor U8608 (N_8608,N_6095,N_6994);
and U8609 (N_8609,N_6306,N_7259);
nand U8610 (N_8610,N_6779,N_7291);
nor U8611 (N_8611,N_6442,N_6825);
nor U8612 (N_8612,N_7009,N_6611);
nor U8613 (N_8613,N_7272,N_7127);
nand U8614 (N_8614,N_6894,N_6372);
nand U8615 (N_8615,N_7295,N_6423);
nor U8616 (N_8616,N_6760,N_6787);
nor U8617 (N_8617,N_6672,N_6051);
and U8618 (N_8618,N_6257,N_6416);
nor U8619 (N_8619,N_6360,N_6092);
and U8620 (N_8620,N_6943,N_6229);
and U8621 (N_8621,N_6337,N_6717);
or U8622 (N_8622,N_6963,N_6956);
and U8623 (N_8623,N_7290,N_6490);
and U8624 (N_8624,N_7158,N_6583);
xnor U8625 (N_8625,N_6930,N_6912);
nor U8626 (N_8626,N_7227,N_6365);
or U8627 (N_8627,N_7067,N_7308);
or U8628 (N_8628,N_7211,N_7172);
nor U8629 (N_8629,N_6093,N_6646);
and U8630 (N_8630,N_7084,N_6170);
and U8631 (N_8631,N_6749,N_7172);
and U8632 (N_8632,N_7031,N_6509);
and U8633 (N_8633,N_6294,N_6981);
or U8634 (N_8634,N_7366,N_7493);
xor U8635 (N_8635,N_6041,N_6113);
and U8636 (N_8636,N_6896,N_6254);
nand U8637 (N_8637,N_6450,N_7387);
nor U8638 (N_8638,N_6238,N_6902);
or U8639 (N_8639,N_7022,N_6584);
and U8640 (N_8640,N_6576,N_6453);
xor U8641 (N_8641,N_6363,N_6045);
or U8642 (N_8642,N_6969,N_6023);
xnor U8643 (N_8643,N_7264,N_6279);
or U8644 (N_8644,N_7238,N_6311);
or U8645 (N_8645,N_6561,N_6493);
and U8646 (N_8646,N_7148,N_6280);
nor U8647 (N_8647,N_6075,N_6705);
or U8648 (N_8648,N_6245,N_7107);
and U8649 (N_8649,N_6858,N_6972);
nor U8650 (N_8650,N_6629,N_7394);
or U8651 (N_8651,N_6186,N_6778);
or U8652 (N_8652,N_6332,N_6004);
xnor U8653 (N_8653,N_6817,N_6249);
nor U8654 (N_8654,N_6565,N_6787);
or U8655 (N_8655,N_6773,N_7421);
and U8656 (N_8656,N_6913,N_6237);
nand U8657 (N_8657,N_7252,N_6954);
xnor U8658 (N_8658,N_6471,N_6231);
or U8659 (N_8659,N_6648,N_6823);
and U8660 (N_8660,N_6237,N_6504);
nand U8661 (N_8661,N_7288,N_7044);
or U8662 (N_8662,N_6721,N_6753);
nor U8663 (N_8663,N_6987,N_7445);
or U8664 (N_8664,N_6821,N_6849);
nor U8665 (N_8665,N_6076,N_6384);
nand U8666 (N_8666,N_6910,N_7483);
xor U8667 (N_8667,N_6948,N_6877);
nand U8668 (N_8668,N_6078,N_6221);
xnor U8669 (N_8669,N_7473,N_6088);
xnor U8670 (N_8670,N_7337,N_7334);
or U8671 (N_8671,N_7295,N_6760);
and U8672 (N_8672,N_6140,N_6703);
and U8673 (N_8673,N_6447,N_6854);
nand U8674 (N_8674,N_7277,N_6337);
and U8675 (N_8675,N_7356,N_7297);
or U8676 (N_8676,N_6008,N_6284);
nand U8677 (N_8677,N_7234,N_7215);
nand U8678 (N_8678,N_6359,N_6622);
nor U8679 (N_8679,N_6130,N_6524);
or U8680 (N_8680,N_6126,N_6877);
nor U8681 (N_8681,N_6629,N_7264);
xor U8682 (N_8682,N_6245,N_6024);
and U8683 (N_8683,N_6018,N_6628);
or U8684 (N_8684,N_7312,N_6165);
nor U8685 (N_8685,N_7266,N_7316);
nor U8686 (N_8686,N_6884,N_6701);
nor U8687 (N_8687,N_7346,N_6878);
nor U8688 (N_8688,N_6828,N_6624);
xnor U8689 (N_8689,N_6467,N_6625);
and U8690 (N_8690,N_6710,N_6888);
nor U8691 (N_8691,N_6946,N_6434);
nand U8692 (N_8692,N_6470,N_6822);
nand U8693 (N_8693,N_6709,N_7345);
nand U8694 (N_8694,N_6783,N_6566);
nand U8695 (N_8695,N_7300,N_6331);
nor U8696 (N_8696,N_6579,N_6666);
nand U8697 (N_8697,N_6357,N_6317);
xnor U8698 (N_8698,N_6328,N_7304);
nor U8699 (N_8699,N_7478,N_7003);
xnor U8700 (N_8700,N_6204,N_6020);
xor U8701 (N_8701,N_6996,N_6132);
nand U8702 (N_8702,N_7321,N_6980);
nor U8703 (N_8703,N_6014,N_6206);
nor U8704 (N_8704,N_7433,N_6381);
or U8705 (N_8705,N_7406,N_6924);
nor U8706 (N_8706,N_7077,N_7124);
and U8707 (N_8707,N_7017,N_7462);
nor U8708 (N_8708,N_6709,N_7045);
or U8709 (N_8709,N_6282,N_6581);
or U8710 (N_8710,N_7134,N_6090);
nand U8711 (N_8711,N_6461,N_7322);
nor U8712 (N_8712,N_6633,N_6407);
xor U8713 (N_8713,N_7405,N_6185);
and U8714 (N_8714,N_6854,N_7280);
or U8715 (N_8715,N_7086,N_7426);
nor U8716 (N_8716,N_6915,N_7443);
nand U8717 (N_8717,N_6314,N_6522);
nor U8718 (N_8718,N_6184,N_6826);
xnor U8719 (N_8719,N_7012,N_6082);
xnor U8720 (N_8720,N_6530,N_6297);
xnor U8721 (N_8721,N_6396,N_7176);
nor U8722 (N_8722,N_6826,N_6300);
and U8723 (N_8723,N_7439,N_7479);
nor U8724 (N_8724,N_7204,N_7443);
nand U8725 (N_8725,N_6714,N_6581);
and U8726 (N_8726,N_6220,N_7174);
xnor U8727 (N_8727,N_6087,N_6209);
and U8728 (N_8728,N_6050,N_6926);
nor U8729 (N_8729,N_6503,N_6513);
nor U8730 (N_8730,N_6713,N_7291);
and U8731 (N_8731,N_6454,N_6689);
nand U8732 (N_8732,N_6810,N_7298);
xnor U8733 (N_8733,N_7298,N_7064);
and U8734 (N_8734,N_7011,N_6296);
and U8735 (N_8735,N_7396,N_7315);
xnor U8736 (N_8736,N_7232,N_6723);
xnor U8737 (N_8737,N_6384,N_6757);
nand U8738 (N_8738,N_7251,N_7486);
nand U8739 (N_8739,N_6683,N_6334);
and U8740 (N_8740,N_7137,N_7470);
or U8741 (N_8741,N_6494,N_7409);
nor U8742 (N_8742,N_7187,N_6175);
nor U8743 (N_8743,N_6200,N_7435);
and U8744 (N_8744,N_6602,N_6889);
nor U8745 (N_8745,N_6266,N_6638);
and U8746 (N_8746,N_6381,N_7173);
and U8747 (N_8747,N_6494,N_6402);
and U8748 (N_8748,N_6369,N_6785);
nor U8749 (N_8749,N_6672,N_7345);
xor U8750 (N_8750,N_6628,N_7136);
nor U8751 (N_8751,N_7479,N_6141);
xor U8752 (N_8752,N_6874,N_6808);
or U8753 (N_8753,N_6223,N_7414);
nor U8754 (N_8754,N_6359,N_6853);
or U8755 (N_8755,N_6390,N_6877);
nor U8756 (N_8756,N_6953,N_6882);
or U8757 (N_8757,N_6390,N_6349);
nor U8758 (N_8758,N_6073,N_6052);
and U8759 (N_8759,N_6731,N_6068);
or U8760 (N_8760,N_6721,N_6765);
nor U8761 (N_8761,N_6474,N_6378);
and U8762 (N_8762,N_7280,N_7161);
nand U8763 (N_8763,N_6608,N_6113);
and U8764 (N_8764,N_6158,N_7154);
nand U8765 (N_8765,N_6424,N_7123);
xor U8766 (N_8766,N_7213,N_6305);
xor U8767 (N_8767,N_6716,N_6028);
and U8768 (N_8768,N_6079,N_6322);
nand U8769 (N_8769,N_7231,N_6147);
nor U8770 (N_8770,N_6447,N_7327);
nor U8771 (N_8771,N_6599,N_6568);
nand U8772 (N_8772,N_6487,N_6867);
nor U8773 (N_8773,N_6627,N_6436);
or U8774 (N_8774,N_7084,N_6075);
nand U8775 (N_8775,N_6511,N_7401);
nand U8776 (N_8776,N_6615,N_6640);
nor U8777 (N_8777,N_6656,N_6779);
xor U8778 (N_8778,N_7395,N_6612);
nor U8779 (N_8779,N_6816,N_6600);
nor U8780 (N_8780,N_6819,N_7178);
and U8781 (N_8781,N_6070,N_6622);
nor U8782 (N_8782,N_7332,N_7156);
or U8783 (N_8783,N_6517,N_7325);
or U8784 (N_8784,N_6620,N_7211);
nand U8785 (N_8785,N_6246,N_6267);
nand U8786 (N_8786,N_6789,N_6121);
xor U8787 (N_8787,N_6374,N_6969);
and U8788 (N_8788,N_6167,N_6376);
and U8789 (N_8789,N_6964,N_6206);
and U8790 (N_8790,N_6700,N_6222);
and U8791 (N_8791,N_7353,N_6414);
and U8792 (N_8792,N_7010,N_6537);
nor U8793 (N_8793,N_7105,N_6431);
xor U8794 (N_8794,N_7450,N_6262);
nand U8795 (N_8795,N_6850,N_6524);
and U8796 (N_8796,N_6225,N_6604);
nor U8797 (N_8797,N_6570,N_7348);
xnor U8798 (N_8798,N_6230,N_6148);
xnor U8799 (N_8799,N_6881,N_6555);
xor U8800 (N_8800,N_7192,N_6688);
nor U8801 (N_8801,N_6179,N_7311);
xnor U8802 (N_8802,N_6406,N_6866);
nand U8803 (N_8803,N_6809,N_7463);
and U8804 (N_8804,N_7272,N_7264);
or U8805 (N_8805,N_6898,N_6810);
xor U8806 (N_8806,N_7036,N_6427);
xnor U8807 (N_8807,N_6715,N_6431);
and U8808 (N_8808,N_6168,N_6315);
and U8809 (N_8809,N_7278,N_7256);
xnor U8810 (N_8810,N_6107,N_6590);
and U8811 (N_8811,N_6474,N_6544);
xor U8812 (N_8812,N_6760,N_6411);
or U8813 (N_8813,N_6873,N_6657);
nor U8814 (N_8814,N_7258,N_6594);
xor U8815 (N_8815,N_6007,N_6683);
nor U8816 (N_8816,N_7178,N_6846);
or U8817 (N_8817,N_6216,N_6771);
xnor U8818 (N_8818,N_6559,N_6762);
xnor U8819 (N_8819,N_6910,N_6623);
xnor U8820 (N_8820,N_7444,N_7219);
nand U8821 (N_8821,N_7094,N_6872);
nor U8822 (N_8822,N_6157,N_6834);
or U8823 (N_8823,N_7124,N_6289);
nand U8824 (N_8824,N_6926,N_7343);
nor U8825 (N_8825,N_6098,N_7149);
or U8826 (N_8826,N_6201,N_6715);
nor U8827 (N_8827,N_6251,N_6961);
or U8828 (N_8828,N_6452,N_6798);
xor U8829 (N_8829,N_7008,N_6157);
nor U8830 (N_8830,N_6030,N_6080);
nand U8831 (N_8831,N_6987,N_7227);
xor U8832 (N_8832,N_6772,N_6886);
nand U8833 (N_8833,N_7203,N_6550);
nand U8834 (N_8834,N_6543,N_7387);
xor U8835 (N_8835,N_6442,N_6288);
nand U8836 (N_8836,N_6037,N_6813);
nand U8837 (N_8837,N_7215,N_6026);
nor U8838 (N_8838,N_6025,N_6186);
nand U8839 (N_8839,N_6487,N_6402);
or U8840 (N_8840,N_7341,N_7387);
and U8841 (N_8841,N_7395,N_6423);
xnor U8842 (N_8842,N_6189,N_7273);
nor U8843 (N_8843,N_6178,N_6917);
and U8844 (N_8844,N_6763,N_6651);
or U8845 (N_8845,N_6559,N_6198);
nand U8846 (N_8846,N_6882,N_6861);
xnor U8847 (N_8847,N_6161,N_7013);
nand U8848 (N_8848,N_6054,N_7319);
or U8849 (N_8849,N_7477,N_6642);
nor U8850 (N_8850,N_7313,N_7108);
and U8851 (N_8851,N_6464,N_6560);
or U8852 (N_8852,N_6885,N_6945);
nand U8853 (N_8853,N_7162,N_6820);
nand U8854 (N_8854,N_6593,N_7253);
or U8855 (N_8855,N_6520,N_6447);
nand U8856 (N_8856,N_6507,N_6301);
or U8857 (N_8857,N_6834,N_6651);
or U8858 (N_8858,N_6716,N_7344);
nand U8859 (N_8859,N_7099,N_6350);
nand U8860 (N_8860,N_6500,N_6457);
nor U8861 (N_8861,N_6508,N_6092);
and U8862 (N_8862,N_7214,N_6928);
and U8863 (N_8863,N_7490,N_6530);
or U8864 (N_8864,N_6804,N_6118);
xnor U8865 (N_8865,N_6022,N_6743);
or U8866 (N_8866,N_6554,N_6184);
xnor U8867 (N_8867,N_6465,N_7231);
nand U8868 (N_8868,N_7110,N_7175);
nand U8869 (N_8869,N_7023,N_6397);
nor U8870 (N_8870,N_7003,N_6917);
nor U8871 (N_8871,N_7239,N_6206);
nor U8872 (N_8872,N_6990,N_7219);
or U8873 (N_8873,N_7126,N_6711);
and U8874 (N_8874,N_6324,N_7435);
and U8875 (N_8875,N_7060,N_6662);
or U8876 (N_8876,N_7036,N_6622);
or U8877 (N_8877,N_6340,N_7212);
xor U8878 (N_8878,N_6138,N_7383);
xnor U8879 (N_8879,N_7054,N_6151);
xnor U8880 (N_8880,N_6238,N_7404);
xnor U8881 (N_8881,N_6363,N_6233);
nand U8882 (N_8882,N_6176,N_6488);
or U8883 (N_8883,N_6285,N_6549);
nand U8884 (N_8884,N_6105,N_7194);
nand U8885 (N_8885,N_7040,N_6101);
xnor U8886 (N_8886,N_6372,N_7322);
or U8887 (N_8887,N_6638,N_6220);
nand U8888 (N_8888,N_6283,N_7185);
or U8889 (N_8889,N_6730,N_6163);
and U8890 (N_8890,N_6565,N_6395);
nor U8891 (N_8891,N_6395,N_7123);
nand U8892 (N_8892,N_7376,N_6478);
nand U8893 (N_8893,N_7139,N_6539);
nor U8894 (N_8894,N_7356,N_6185);
nand U8895 (N_8895,N_6081,N_7082);
or U8896 (N_8896,N_6191,N_7169);
nor U8897 (N_8897,N_6686,N_6791);
nor U8898 (N_8898,N_7027,N_6276);
nor U8899 (N_8899,N_6311,N_6289);
nand U8900 (N_8900,N_6739,N_6607);
and U8901 (N_8901,N_7401,N_6595);
xnor U8902 (N_8902,N_7426,N_6746);
and U8903 (N_8903,N_7072,N_6692);
or U8904 (N_8904,N_7076,N_6015);
xnor U8905 (N_8905,N_6095,N_6718);
nand U8906 (N_8906,N_6322,N_6560);
or U8907 (N_8907,N_6112,N_6541);
and U8908 (N_8908,N_7236,N_6387);
nand U8909 (N_8909,N_6498,N_6332);
xor U8910 (N_8910,N_7157,N_7241);
and U8911 (N_8911,N_6872,N_6100);
xnor U8912 (N_8912,N_6467,N_6850);
xnor U8913 (N_8913,N_6087,N_6489);
and U8914 (N_8914,N_7334,N_7335);
and U8915 (N_8915,N_7064,N_6387);
and U8916 (N_8916,N_6135,N_7310);
and U8917 (N_8917,N_6149,N_7287);
and U8918 (N_8918,N_6594,N_6794);
nand U8919 (N_8919,N_6864,N_6073);
and U8920 (N_8920,N_6781,N_6292);
nand U8921 (N_8921,N_6997,N_7286);
nor U8922 (N_8922,N_7432,N_6229);
xnor U8923 (N_8923,N_7054,N_7139);
xor U8924 (N_8924,N_7208,N_7294);
xnor U8925 (N_8925,N_6011,N_7473);
nor U8926 (N_8926,N_6961,N_7027);
nand U8927 (N_8927,N_6481,N_6395);
or U8928 (N_8928,N_7270,N_6625);
xor U8929 (N_8929,N_6433,N_6553);
and U8930 (N_8930,N_7084,N_6233);
and U8931 (N_8931,N_7073,N_7485);
xor U8932 (N_8932,N_6457,N_6339);
or U8933 (N_8933,N_6153,N_6504);
nor U8934 (N_8934,N_6870,N_6578);
nand U8935 (N_8935,N_6342,N_6306);
nor U8936 (N_8936,N_7292,N_6446);
nand U8937 (N_8937,N_7087,N_6035);
or U8938 (N_8938,N_7095,N_6081);
xnor U8939 (N_8939,N_7108,N_6609);
xnor U8940 (N_8940,N_6032,N_7475);
nor U8941 (N_8941,N_7496,N_7210);
or U8942 (N_8942,N_6876,N_6093);
or U8943 (N_8943,N_7246,N_6880);
nor U8944 (N_8944,N_7222,N_6294);
xor U8945 (N_8945,N_7284,N_6095);
nand U8946 (N_8946,N_7022,N_6915);
and U8947 (N_8947,N_6850,N_6721);
or U8948 (N_8948,N_6909,N_6057);
nand U8949 (N_8949,N_6204,N_6545);
and U8950 (N_8950,N_6792,N_7498);
or U8951 (N_8951,N_6196,N_6789);
nand U8952 (N_8952,N_6541,N_7378);
nand U8953 (N_8953,N_7251,N_7182);
nand U8954 (N_8954,N_6772,N_6012);
and U8955 (N_8955,N_7054,N_6906);
or U8956 (N_8956,N_6736,N_6188);
or U8957 (N_8957,N_7305,N_6997);
or U8958 (N_8958,N_6031,N_6262);
or U8959 (N_8959,N_6056,N_7039);
xnor U8960 (N_8960,N_7423,N_7098);
xor U8961 (N_8961,N_6858,N_6452);
and U8962 (N_8962,N_6025,N_7101);
nand U8963 (N_8963,N_7174,N_6467);
or U8964 (N_8964,N_6757,N_7352);
xnor U8965 (N_8965,N_6247,N_7024);
or U8966 (N_8966,N_6126,N_6244);
xnor U8967 (N_8967,N_6119,N_6945);
and U8968 (N_8968,N_7013,N_6376);
or U8969 (N_8969,N_6111,N_6415);
xnor U8970 (N_8970,N_7484,N_6107);
nand U8971 (N_8971,N_6601,N_6558);
nand U8972 (N_8972,N_7222,N_6284);
or U8973 (N_8973,N_6905,N_6792);
xnor U8974 (N_8974,N_6416,N_6365);
nor U8975 (N_8975,N_6196,N_6141);
xnor U8976 (N_8976,N_6091,N_6503);
xor U8977 (N_8977,N_6172,N_6590);
xor U8978 (N_8978,N_6868,N_7247);
nor U8979 (N_8979,N_7442,N_7406);
or U8980 (N_8980,N_6514,N_7383);
nor U8981 (N_8981,N_7144,N_6894);
nor U8982 (N_8982,N_6626,N_6887);
nor U8983 (N_8983,N_7265,N_7123);
or U8984 (N_8984,N_7000,N_7343);
and U8985 (N_8985,N_7246,N_7441);
nand U8986 (N_8986,N_6679,N_7469);
nand U8987 (N_8987,N_6540,N_6549);
and U8988 (N_8988,N_6564,N_6971);
xor U8989 (N_8989,N_6973,N_7465);
or U8990 (N_8990,N_6444,N_6609);
xnor U8991 (N_8991,N_6055,N_7027);
and U8992 (N_8992,N_7301,N_6433);
nand U8993 (N_8993,N_7334,N_6787);
and U8994 (N_8994,N_6093,N_6692);
nand U8995 (N_8995,N_7331,N_7472);
xnor U8996 (N_8996,N_7091,N_6942);
xor U8997 (N_8997,N_6992,N_6999);
nand U8998 (N_8998,N_7093,N_6644);
or U8999 (N_8999,N_6401,N_6863);
and U9000 (N_9000,N_8992,N_8674);
nand U9001 (N_9001,N_7703,N_7525);
nand U9002 (N_9002,N_7723,N_8426);
xnor U9003 (N_9003,N_8822,N_7975);
or U9004 (N_9004,N_7678,N_8051);
and U9005 (N_9005,N_8146,N_8127);
nor U9006 (N_9006,N_7559,N_7550);
nor U9007 (N_9007,N_8996,N_8695);
xor U9008 (N_9008,N_8932,N_7648);
or U9009 (N_9009,N_8858,N_8156);
and U9010 (N_9010,N_8647,N_7582);
and U9011 (N_9011,N_8696,N_8020);
and U9012 (N_9012,N_7634,N_8786);
nor U9013 (N_9013,N_8299,N_7553);
nand U9014 (N_9014,N_8045,N_7526);
and U9015 (N_9015,N_7967,N_8964);
or U9016 (N_9016,N_8735,N_8739);
nor U9017 (N_9017,N_8798,N_8547);
or U9018 (N_9018,N_7666,N_8881);
nand U9019 (N_9019,N_8869,N_7893);
xor U9020 (N_9020,N_8656,N_8870);
or U9021 (N_9021,N_7806,N_8832);
or U9022 (N_9022,N_8821,N_7583);
and U9023 (N_9023,N_8601,N_7979);
and U9024 (N_9024,N_8014,N_8662);
and U9025 (N_9025,N_7964,N_8260);
nor U9026 (N_9026,N_8002,N_8125);
and U9027 (N_9027,N_7754,N_8981);
and U9028 (N_9028,N_8036,N_8585);
and U9029 (N_9029,N_8568,N_8612);
xnor U9030 (N_9030,N_7694,N_7923);
nand U9031 (N_9031,N_8515,N_7689);
and U9032 (N_9032,N_8684,N_8635);
xor U9033 (N_9033,N_7953,N_8969);
nor U9034 (N_9034,N_7847,N_8142);
or U9035 (N_9035,N_7821,N_8683);
and U9036 (N_9036,N_8393,N_8205);
nand U9037 (N_9037,N_8615,N_8144);
xnor U9038 (N_9038,N_8166,N_8376);
and U9039 (N_9039,N_7972,N_7595);
xnor U9040 (N_9040,N_8746,N_8658);
xnor U9041 (N_9041,N_7884,N_8591);
nand U9042 (N_9042,N_7511,N_7661);
xnor U9043 (N_9043,N_8741,N_8543);
or U9044 (N_9044,N_8906,N_7504);
and U9045 (N_9045,N_7839,N_8064);
nand U9046 (N_9046,N_7643,N_7775);
xnor U9047 (N_9047,N_7992,N_7921);
nor U9048 (N_9048,N_8967,N_8318);
nor U9049 (N_9049,N_8307,N_8067);
and U9050 (N_9050,N_8015,N_8315);
xnor U9051 (N_9051,N_7960,N_8337);
nand U9052 (N_9052,N_8104,N_7716);
xor U9053 (N_9053,N_8590,N_7632);
and U9054 (N_9054,N_8183,N_7566);
nor U9055 (N_9055,N_8845,N_7513);
xnor U9056 (N_9056,N_8090,N_8617);
xor U9057 (N_9057,N_8451,N_8973);
and U9058 (N_9058,N_7853,N_8583);
nand U9059 (N_9059,N_7613,N_7672);
xnor U9060 (N_9060,N_8846,N_8633);
xor U9061 (N_9061,N_7524,N_8356);
nand U9062 (N_9062,N_8801,N_7840);
xnor U9063 (N_9063,N_7532,N_8566);
nand U9064 (N_9064,N_8797,N_7835);
nor U9065 (N_9065,N_8075,N_8332);
nor U9066 (N_9066,N_7818,N_8625);
nand U9067 (N_9067,N_8993,N_8143);
nor U9068 (N_9068,N_8302,N_8306);
or U9069 (N_9069,N_8250,N_8001);
xor U9070 (N_9070,N_8800,N_8772);
nand U9071 (N_9071,N_7955,N_7662);
or U9072 (N_9072,N_7756,N_8244);
nand U9073 (N_9073,N_8806,N_8873);
or U9074 (N_9074,N_8371,N_8502);
and U9075 (N_9075,N_8991,N_8499);
nor U9076 (N_9076,N_8460,N_7958);
nor U9077 (N_9077,N_8933,N_8910);
xor U9078 (N_9078,N_8458,N_7877);
or U9079 (N_9079,N_8366,N_8341);
nand U9080 (N_9080,N_8087,N_8079);
nor U9081 (N_9081,N_8437,N_8007);
or U9082 (N_9082,N_8101,N_7867);
nor U9083 (N_9083,N_8233,N_8638);
or U9084 (N_9084,N_8775,N_7782);
nand U9085 (N_9085,N_7738,N_8251);
nor U9086 (N_9086,N_7714,N_8455);
or U9087 (N_9087,N_7527,N_7682);
xnor U9088 (N_9088,N_7815,N_7752);
and U9089 (N_9089,N_8081,N_8164);
nor U9090 (N_9090,N_8468,N_7501);
and U9091 (N_9091,N_8073,N_7795);
or U9092 (N_9092,N_8571,N_8482);
and U9093 (N_9093,N_7909,N_8196);
xor U9094 (N_9094,N_7799,N_7858);
or U9095 (N_9095,N_7699,N_7871);
nor U9096 (N_9096,N_8833,N_8062);
xnor U9097 (N_9097,N_7649,N_8349);
or U9098 (N_9098,N_7769,N_7855);
nor U9099 (N_9099,N_8271,N_8290);
nand U9100 (N_9100,N_8540,N_8321);
and U9101 (N_9101,N_8477,N_7904);
and U9102 (N_9102,N_8363,N_7940);
nor U9103 (N_9103,N_8530,N_8140);
xnor U9104 (N_9104,N_8016,N_8569);
nand U9105 (N_9105,N_8017,N_7852);
and U9106 (N_9106,N_7599,N_8931);
xnor U9107 (N_9107,N_8918,N_7771);
or U9108 (N_9108,N_8274,N_8668);
xor U9109 (N_9109,N_8699,N_8224);
xor U9110 (N_9110,N_8550,N_7697);
xor U9111 (N_9111,N_8868,N_8747);
and U9112 (N_9112,N_7735,N_8837);
nand U9113 (N_9113,N_8680,N_8005);
nand U9114 (N_9114,N_8804,N_8395);
and U9115 (N_9115,N_7870,N_8509);
or U9116 (N_9116,N_7552,N_8094);
nand U9117 (N_9117,N_7945,N_7963);
nor U9118 (N_9118,N_7765,N_8849);
nand U9119 (N_9119,N_8528,N_8748);
xnor U9120 (N_9120,N_7618,N_8669);
xor U9121 (N_9121,N_8957,N_8961);
xnor U9122 (N_9122,N_8123,N_7936);
and U9123 (N_9123,N_8984,N_7560);
nand U9124 (N_9124,N_8847,N_8093);
xor U9125 (N_9125,N_8835,N_8080);
xor U9126 (N_9126,N_7556,N_7787);
or U9127 (N_9127,N_8154,N_7605);
or U9128 (N_9128,N_7720,N_8519);
nor U9129 (N_9129,N_7989,N_8313);
nand U9130 (N_9130,N_8273,N_8077);
xor U9131 (N_9131,N_8032,N_7897);
nor U9132 (N_9132,N_8220,N_8416);
or U9133 (N_9133,N_8374,N_8572);
and U9134 (N_9134,N_8359,N_7701);
nor U9135 (N_9135,N_8947,N_8897);
xnor U9136 (N_9136,N_8033,N_7907);
xor U9137 (N_9137,N_7746,N_8789);
or U9138 (N_9138,N_8237,N_8645);
or U9139 (N_9139,N_8796,N_8111);
and U9140 (N_9140,N_8453,N_7730);
and U9141 (N_9141,N_8657,N_8257);
and U9142 (N_9142,N_8900,N_8682);
or U9143 (N_9143,N_8926,N_7624);
or U9144 (N_9144,N_8733,N_8038);
nor U9145 (N_9145,N_8562,N_8107);
nand U9146 (N_9146,N_8608,N_8379);
nor U9147 (N_9147,N_7764,N_8238);
or U9148 (N_9148,N_8195,N_8745);
xnor U9149 (N_9149,N_7590,N_8200);
and U9150 (N_9150,N_7833,N_8281);
nand U9151 (N_9151,N_8598,N_8802);
or U9152 (N_9152,N_7538,N_8161);
and U9153 (N_9153,N_8358,N_7628);
nor U9154 (N_9154,N_7702,N_8908);
xor U9155 (N_9155,N_8278,N_8066);
nor U9156 (N_9156,N_8782,N_8893);
and U9157 (N_9157,N_8085,N_8643);
xor U9158 (N_9158,N_8115,N_8843);
and U9159 (N_9159,N_8121,N_8218);
and U9160 (N_9160,N_8539,N_8945);
nor U9161 (N_9161,N_8576,N_8095);
and U9162 (N_9162,N_8564,N_7739);
and U9163 (N_9163,N_8614,N_7652);
and U9164 (N_9164,N_8487,N_8755);
or U9165 (N_9165,N_8082,N_7760);
or U9166 (N_9166,N_8960,N_8779);
or U9167 (N_9167,N_8544,N_8605);
nor U9168 (N_9168,N_8998,N_8312);
nand U9169 (N_9169,N_8097,N_8369);
and U9170 (N_9170,N_8622,N_8185);
xor U9171 (N_9171,N_7676,N_8567);
and U9172 (N_9172,N_8227,N_7509);
and U9173 (N_9173,N_8841,N_8838);
nand U9174 (N_9174,N_7930,N_8022);
xnor U9175 (N_9175,N_8336,N_7970);
nor U9176 (N_9176,N_8357,N_8558);
nand U9177 (N_9177,N_8488,N_7996);
xnor U9178 (N_9178,N_7625,N_8179);
or U9179 (N_9179,N_8043,N_8948);
or U9180 (N_9180,N_8353,N_7601);
nand U9181 (N_9181,N_8192,N_8268);
nor U9182 (N_9182,N_7646,N_8505);
xnor U9183 (N_9183,N_7743,N_8230);
and U9184 (N_9184,N_8756,N_7696);
xnor U9185 (N_9185,N_7981,N_8974);
nand U9186 (N_9186,N_8480,N_8137);
or U9187 (N_9187,N_8814,N_8325);
nand U9188 (N_9188,N_8414,N_8108);
nand U9189 (N_9189,N_7544,N_8676);
and U9190 (N_9190,N_8848,N_7911);
and U9191 (N_9191,N_8207,N_8331);
nand U9192 (N_9192,N_8021,N_7561);
or U9193 (N_9193,N_8750,N_8825);
nand U9194 (N_9194,N_8355,N_8660);
nor U9195 (N_9195,N_8712,N_8316);
or U9196 (N_9196,N_7908,N_7914);
nor U9197 (N_9197,N_7926,N_8201);
or U9198 (N_9198,N_7660,N_8004);
or U9199 (N_9199,N_7565,N_8623);
xnor U9200 (N_9200,N_7704,N_8327);
or U9201 (N_9201,N_7905,N_7637);
nor U9202 (N_9202,N_8549,N_7857);
and U9203 (N_9203,N_8618,N_8805);
and U9204 (N_9204,N_8593,N_7917);
and U9205 (N_9205,N_7768,N_7816);
nand U9206 (N_9206,N_8134,N_7929);
nand U9207 (N_9207,N_8261,N_7830);
xor U9208 (N_9208,N_7842,N_8098);
nand U9209 (N_9209,N_8880,N_7671);
nand U9210 (N_9210,N_8370,N_8385);
or U9211 (N_9211,N_8661,N_8830);
or U9212 (N_9212,N_8913,N_7688);
and U9213 (N_9213,N_8354,N_7568);
or U9214 (N_9214,N_8026,N_8697);
nand U9215 (N_9215,N_8717,N_8646);
and U9216 (N_9216,N_8221,N_8533);
or U9217 (N_9217,N_8133,N_8124);
or U9218 (N_9218,N_8715,N_8811);
or U9219 (N_9219,N_8603,N_8091);
and U9220 (N_9220,N_7938,N_8287);
and U9221 (N_9221,N_7533,N_8512);
xor U9222 (N_9222,N_7502,N_7772);
nand U9223 (N_9223,N_7535,N_7886);
and U9224 (N_9224,N_8401,N_8874);
or U9225 (N_9225,N_7732,N_8500);
or U9226 (N_9226,N_7731,N_8671);
and U9227 (N_9227,N_8291,N_8890);
xor U9228 (N_9228,N_7635,N_8295);
or U9229 (N_9229,N_7503,N_8145);
nor U9230 (N_9230,N_8361,N_8711);
or U9231 (N_9231,N_7724,N_7757);
and U9232 (N_9232,N_7725,N_8050);
nor U9233 (N_9233,N_7789,N_8664);
or U9234 (N_9234,N_8397,N_8693);
nor U9235 (N_9235,N_8052,N_7793);
xor U9236 (N_9236,N_8044,N_8548);
or U9237 (N_9237,N_7900,N_8710);
nand U9238 (N_9238,N_7594,N_8784);
nor U9239 (N_9239,N_8765,N_8760);
or U9240 (N_9240,N_8280,N_8199);
or U9241 (N_9241,N_8485,N_8850);
nor U9242 (N_9242,N_8724,N_8348);
nor U9243 (N_9243,N_8818,N_7693);
nor U9244 (N_9244,N_8297,N_8602);
nor U9245 (N_9245,N_8186,N_7727);
and U9246 (N_9246,N_8565,N_7564);
and U9247 (N_9247,N_8616,N_8907);
nand U9248 (N_9248,N_7827,N_7781);
and U9249 (N_9249,N_7965,N_8070);
and U9250 (N_9250,N_8507,N_8628);
or U9251 (N_9251,N_7548,N_8494);
xnor U9252 (N_9252,N_7585,N_8937);
nand U9253 (N_9253,N_8063,N_7748);
nor U9254 (N_9254,N_7860,N_8673);
or U9255 (N_9255,N_7865,N_8180);
and U9256 (N_9256,N_8988,N_7747);
nor U9257 (N_9257,N_7939,N_8150);
nor U9258 (N_9258,N_7679,N_8575);
and U9259 (N_9259,N_8905,N_8110);
or U9260 (N_9260,N_7698,N_8570);
nand U9261 (N_9261,N_8398,N_8461);
nand U9262 (N_9262,N_7894,N_8057);
nor U9263 (N_9263,N_8983,N_8580);
xor U9264 (N_9264,N_7801,N_8914);
and U9265 (N_9265,N_8037,N_8761);
or U9266 (N_9266,N_8448,N_8462);
nand U9267 (N_9267,N_8940,N_7920);
and U9268 (N_9268,N_7809,N_7786);
nand U9269 (N_9269,N_8706,N_8714);
xnor U9270 (N_9270,N_7558,N_8839);
xnor U9271 (N_9271,N_8574,N_8642);
and U9272 (N_9272,N_8046,N_8729);
xnor U9273 (N_9273,N_8486,N_8386);
xor U9274 (N_9274,N_8277,N_8853);
nand U9275 (N_9275,N_7687,N_8726);
and U9276 (N_9276,N_8162,N_8351);
xor U9277 (N_9277,N_8734,N_7951);
nand U9278 (N_9278,N_8434,N_8217);
nor U9279 (N_9279,N_8989,N_8537);
nor U9280 (N_9280,N_7627,N_7977);
or U9281 (N_9281,N_7521,N_8934);
and U9282 (N_9282,N_8440,N_7633);
xor U9283 (N_9283,N_7675,N_8383);
nand U9284 (N_9284,N_8427,N_8819);
nand U9285 (N_9285,N_7997,N_8049);
or U9286 (N_9286,N_8240,N_7584);
nand U9287 (N_9287,N_7622,N_8396);
nor U9288 (N_9288,N_8152,N_7849);
nor U9289 (N_9289,N_8131,N_8688);
nor U9290 (N_9290,N_8744,N_8446);
nand U9291 (N_9291,N_7572,N_8599);
or U9292 (N_9292,N_7534,N_8381);
nand U9293 (N_9293,N_7846,N_8132);
or U9294 (N_9294,N_7978,N_8759);
or U9295 (N_9295,N_8301,N_8867);
nor U9296 (N_9296,N_7804,N_7885);
nor U9297 (N_9297,N_8826,N_8394);
or U9298 (N_9298,N_8308,N_8089);
nor U9299 (N_9299,N_8417,N_8935);
or U9300 (N_9300,N_8713,N_7986);
or U9301 (N_9301,N_7934,N_7683);
nand U9302 (N_9302,N_8971,N_8149);
nand U9303 (N_9303,N_8851,N_8820);
or U9304 (N_9304,N_7896,N_8542);
xnor U9305 (N_9305,N_7537,N_7644);
or U9306 (N_9306,N_8148,N_8269);
nand U9307 (N_9307,N_8630,N_8921);
nand U9308 (N_9308,N_8978,N_8253);
and U9309 (N_9309,N_8966,N_7792);
xor U9310 (N_9310,N_7639,N_7629);
xor U9311 (N_9311,N_8013,N_8844);
nor U9312 (N_9312,N_8343,N_7803);
nand U9313 (N_9313,N_7980,N_8326);
nor U9314 (N_9314,N_8339,N_7912);
nor U9315 (N_9315,N_8300,N_8704);
xnor U9316 (N_9316,N_7906,N_8405);
or U9317 (N_9317,N_8069,N_8008);
and U9318 (N_9318,N_8187,N_7510);
nand U9319 (N_9319,N_8247,N_8167);
xnor U9320 (N_9320,N_8632,N_7961);
or U9321 (N_9321,N_7610,N_8958);
nor U9322 (N_9322,N_8294,N_8441);
or U9323 (N_9323,N_8727,N_8424);
or U9324 (N_9324,N_7658,N_8411);
or U9325 (N_9325,N_8667,N_7657);
and U9326 (N_9326,N_8809,N_8579);
or U9327 (N_9327,N_8039,N_8454);
and U9328 (N_9328,N_8019,N_7755);
nand U9329 (N_9329,N_8743,N_7578);
or U9330 (N_9330,N_8484,N_8170);
nor U9331 (N_9331,N_8197,N_7655);
or U9332 (N_9332,N_7918,N_8223);
xnor U9333 (N_9333,N_8692,N_8871);
and U9334 (N_9334,N_7653,N_7528);
and U9335 (N_9335,N_7913,N_8293);
and U9336 (N_9336,N_8588,N_8689);
and U9337 (N_9337,N_8723,N_8634);
nand U9338 (N_9338,N_8267,N_7794);
and U9339 (N_9339,N_8229,N_8029);
nand U9340 (N_9340,N_7895,N_8286);
nor U9341 (N_9341,N_7555,N_8457);
nor U9342 (N_9342,N_7941,N_8624);
nor U9343 (N_9343,N_8687,N_7889);
and U9344 (N_9344,N_8410,N_8919);
xor U9345 (N_9345,N_7680,N_7866);
nand U9346 (N_9346,N_7623,N_7901);
nand U9347 (N_9347,N_7547,N_8065);
nor U9348 (N_9348,N_8864,N_8639);
xor U9349 (N_9349,N_7621,N_7712);
nor U9350 (N_9350,N_8000,N_8024);
nand U9351 (N_9351,N_8231,N_8136);
xor U9352 (N_9352,N_8842,N_8538);
and U9353 (N_9353,N_7545,N_7695);
or U9354 (N_9354,N_8923,N_7606);
and U9355 (N_9355,N_7935,N_8243);
nand U9356 (N_9356,N_8946,N_7761);
and U9357 (N_9357,N_7580,N_7640);
or U9358 (N_9358,N_8663,N_8053);
and U9359 (N_9359,N_8047,N_7798);
xor U9360 (N_9360,N_7593,N_8718);
xor U9361 (N_9361,N_8112,N_8606);
xor U9362 (N_9362,N_8817,N_7881);
xor U9363 (N_9363,N_7924,N_8930);
and U9364 (N_9364,N_7539,N_7665);
xnor U9365 (N_9365,N_7668,N_7726);
nand U9366 (N_9366,N_7956,N_7927);
and U9367 (N_9367,N_7514,N_8762);
and U9368 (N_9368,N_7859,N_8790);
xor U9369 (N_9369,N_8524,N_8987);
and U9370 (N_9370,N_8006,N_8768);
and U9371 (N_9371,N_8677,N_8040);
xor U9372 (N_9372,N_7834,N_7626);
nor U9373 (N_9373,N_8999,N_7691);
nor U9374 (N_9374,N_8219,N_8518);
nor U9375 (N_9375,N_8491,N_7876);
nor U9376 (N_9376,N_8702,N_8815);
xnor U9377 (N_9377,N_8577,N_7684);
nand U9378 (N_9378,N_8887,N_8432);
xnor U9379 (N_9379,N_7808,N_7734);
xnor U9380 (N_9380,N_8130,N_8780);
or U9381 (N_9381,N_8232,N_8650);
xnor U9382 (N_9382,N_8884,N_8803);
or U9383 (N_9383,N_7888,N_8228);
xor U9384 (N_9384,N_8698,N_8666);
nand U9385 (N_9385,N_8288,N_8275);
nand U9386 (N_9386,N_8452,N_8895);
and U9387 (N_9387,N_7631,N_8560);
or U9388 (N_9388,N_7844,N_7994);
and U9389 (N_9389,N_7825,N_8103);
or U9390 (N_9390,N_7600,N_8445);
nor U9391 (N_9391,N_8708,N_8912);
and U9392 (N_9392,N_8471,N_8431);
xnor U9393 (N_9393,N_8030,N_8298);
or U9394 (N_9394,N_7592,N_8404);
xnor U9395 (N_9395,N_7774,N_8292);
and U9396 (N_9396,N_8953,N_8373);
nand U9397 (N_9397,N_8936,N_8883);
and U9398 (N_9398,N_8951,N_8279);
or U9399 (N_9399,N_8686,N_8654);
and U9400 (N_9400,N_7785,N_7573);
or U9401 (N_9401,N_8909,N_7932);
xnor U9402 (N_9402,N_7674,N_7903);
xnor U9403 (N_9403,N_8866,N_7529);
nor U9404 (N_9404,N_8763,N_8060);
nor U9405 (N_9405,N_8467,N_8225);
or U9406 (N_9406,N_7673,N_7788);
nor U9407 (N_9407,N_8018,N_8831);
nor U9408 (N_9408,N_7915,N_8836);
and U9409 (N_9409,N_8465,N_8665);
nor U9410 (N_9410,N_8408,N_8757);
or U9411 (N_9411,N_8235,N_8700);
or U9412 (N_9412,N_8556,N_8545);
nand U9413 (N_9413,N_7952,N_8877);
and U9414 (N_9414,N_8776,N_8470);
xnor U9415 (N_9415,N_7990,N_8752);
nand U9416 (N_9416,N_7848,N_8248);
nand U9417 (N_9417,N_7651,N_8211);
or U9418 (N_9418,N_7557,N_7937);
xor U9419 (N_9419,N_7931,N_8425);
and U9420 (N_9420,N_8521,N_8435);
xnor U9421 (N_9421,N_7868,N_7784);
or U9422 (N_9422,N_8527,N_8319);
xor U9423 (N_9423,N_8159,N_8420);
and U9424 (N_9424,N_7591,N_8245);
or U9425 (N_9425,N_7718,N_8042);
nor U9426 (N_9426,N_8546,N_7925);
or U9427 (N_9427,N_7851,N_8289);
xnor U9428 (N_9428,N_8430,N_8754);
nand U9429 (N_9429,N_8423,N_8982);
nor U9430 (N_9430,N_7948,N_8709);
and U9431 (N_9431,N_7563,N_7959);
xnor U9432 (N_9432,N_7971,N_7777);
nand U9433 (N_9433,N_8382,N_8504);
xor U9434 (N_9434,N_8994,N_8861);
or U9435 (N_9435,N_8419,N_7619);
nor U9436 (N_9436,N_7729,N_8118);
nand U9437 (N_9437,N_8003,N_7663);
xnor U9438 (N_9438,N_7823,N_7562);
xnor U9439 (N_9439,N_8340,N_8813);
nand U9440 (N_9440,N_8116,N_7836);
or U9441 (N_9441,N_8479,N_8899);
or U9442 (N_9442,N_8514,N_8888);
xnor U9443 (N_9443,N_8557,N_7614);
nand U9444 (N_9444,N_8892,N_8249);
xor U9445 (N_9445,N_8636,N_8078);
nor U9446 (N_9446,N_8898,N_8753);
nor U9447 (N_9447,N_7811,N_7611);
nor U9448 (N_9448,N_8141,N_8190);
nor U9449 (N_9449,N_8338,N_8535);
nor U9450 (N_9450,N_8189,N_8807);
nand U9451 (N_9451,N_8429,N_8335);
nor U9452 (N_9452,N_8607,N_8594);
xor U9453 (N_9453,N_8659,N_7805);
xnor U9454 (N_9454,N_8236,N_7603);
or U9455 (N_9455,N_8113,N_8407);
or U9456 (N_9456,N_8169,N_7944);
and U9457 (N_9457,N_7711,N_7750);
or U9458 (N_9458,N_8924,N_8072);
or U9459 (N_9459,N_8592,N_8011);
xor U9460 (N_9460,N_7549,N_7783);
nor U9461 (N_9461,N_7983,N_8330);
or U9462 (N_9462,N_8391,N_7645);
or U9463 (N_9463,N_7642,N_7540);
nor U9464 (N_9464,N_8777,N_8171);
or U9465 (N_9465,N_7522,N_7519);
and U9466 (N_9466,N_8955,N_8516);
nor U9467 (N_9467,N_7576,N_8439);
and U9468 (N_9468,N_8342,N_8627);
or U9469 (N_9469,N_7737,N_8956);
and U9470 (N_9470,N_8855,N_8368);
or U9471 (N_9471,N_8239,N_7922);
xor U9472 (N_9472,N_8525,N_8498);
or U9473 (N_9473,N_8323,N_8728);
nand U9474 (N_9474,N_7837,N_7898);
or U9475 (N_9475,N_8928,N_8347);
nor U9476 (N_9476,N_8497,N_8962);
or U9477 (N_9477,N_8406,N_7700);
or U9478 (N_9478,N_8513,N_7843);
and U9479 (N_9479,N_7541,N_8959);
nand U9480 (N_9480,N_8202,N_8751);
xnor U9481 (N_9481,N_8096,N_8506);
and U9482 (N_9482,N_8573,N_8520);
and U9483 (N_9483,N_7766,N_8380);
xnor U9484 (N_9484,N_7773,N_7543);
or U9485 (N_9485,N_8725,N_8903);
nor U9486 (N_9486,N_8968,N_8027);
or U9487 (N_9487,N_8681,N_8421);
and U9488 (N_9488,N_8138,N_7790);
and U9489 (N_9489,N_8882,N_8105);
xnor U9490 (N_9490,N_8309,N_8422);
xor U9491 (N_9491,N_7797,N_8210);
and U9492 (N_9492,N_8503,N_7838);
nor U9493 (N_9493,N_8400,N_7579);
and U9494 (N_9494,N_7988,N_7767);
nor U9495 (N_9495,N_7598,N_8764);
xnor U9496 (N_9496,N_7982,N_7916);
nor U9497 (N_9497,N_8263,N_8360);
or U9498 (N_9498,N_8653,N_8773);
or U9499 (N_9499,N_8372,N_8736);
nor U9500 (N_9500,N_8977,N_8778);
and U9501 (N_9501,N_8204,N_7705);
or U9502 (N_9502,N_8889,N_8076);
nor U9503 (N_9503,N_7570,N_7589);
and U9504 (N_9504,N_7828,N_7826);
or U9505 (N_9505,N_7968,N_8995);
nor U9506 (N_9506,N_8552,N_8828);
nor U9507 (N_9507,N_8375,N_7554);
nor U9508 (N_9508,N_7681,N_8412);
or U9509 (N_9509,N_8262,N_8241);
and U9510 (N_9510,N_8466,N_8596);
and U9511 (N_9511,N_8876,N_7780);
and U9512 (N_9512,N_8084,N_8922);
nand U9513 (N_9513,N_8352,N_8810);
or U9514 (N_9514,N_7630,N_8092);
nand U9515 (N_9515,N_7740,N_7891);
nand U9516 (N_9516,N_7892,N_7506);
nor U9517 (N_9517,N_7985,N_7841);
or U9518 (N_9518,N_8365,N_8554);
nand U9519 (N_9519,N_7736,N_8917);
or U9520 (N_9520,N_8384,N_8860);
nand U9521 (N_9521,N_8305,N_8463);
and U9522 (N_9522,N_8031,N_7864);
and U9523 (N_9523,N_8862,N_8194);
or U9524 (N_9524,N_8068,N_8102);
xnor U9525 (N_9525,N_8182,N_8175);
or U9526 (N_9526,N_7749,N_8816);
xnor U9527 (N_9527,N_7722,N_7779);
nor U9528 (N_9528,N_7770,N_8242);
nand U9529 (N_9529,N_7530,N_7822);
or U9530 (N_9530,N_8058,N_7536);
nor U9531 (N_9531,N_7862,N_8334);
and U9532 (N_9532,N_8061,N_7602);
and U9533 (N_9533,N_8531,N_8976);
nand U9534 (N_9534,N_8203,N_7616);
or U9535 (N_9535,N_8255,N_8329);
or U9536 (N_9536,N_8012,N_7664);
and U9537 (N_9537,N_8469,N_7517);
xnor U9538 (N_9538,N_8872,N_7636);
nor U9539 (N_9539,N_8270,N_8322);
xor U9540 (N_9540,N_8774,N_7902);
nand U9541 (N_9541,N_7819,N_8891);
or U9542 (N_9542,N_7824,N_8413);
nand U9543 (N_9543,N_7943,N_8264);
or U9544 (N_9544,N_7942,N_8378);
or U9545 (N_9545,N_8100,N_8367);
nand U9546 (N_9546,N_8651,N_8758);
nand U9547 (N_9547,N_8054,N_8010);
or U9548 (N_9548,N_8389,N_7820);
and U9549 (N_9549,N_7546,N_8252);
and U9550 (N_9550,N_8311,N_7947);
xnor U9551 (N_9551,N_7919,N_7974);
xnor U9552 (N_9552,N_8120,N_8793);
or U9553 (N_9553,N_8600,N_8559);
and U9554 (N_9554,N_7577,N_8433);
and U9555 (N_9555,N_8317,N_8328);
and U9556 (N_9556,N_8324,N_7710);
nand U9557 (N_9557,N_8911,N_8857);
nand U9558 (N_9558,N_7597,N_8938);
xnor U9559 (N_9559,N_8694,N_7719);
and U9560 (N_9560,N_8586,N_8675);
or U9561 (N_9561,N_8532,N_8128);
nor U9562 (N_9562,N_7667,N_8282);
or U9563 (N_9563,N_7969,N_7966);
nor U9564 (N_9564,N_8508,N_7812);
nor U9565 (N_9565,N_7505,N_8941);
or U9566 (N_9566,N_7878,N_8447);
xnor U9567 (N_9567,N_8920,N_7741);
or U9568 (N_9568,N_7817,N_8126);
nand U9569 (N_9569,N_8442,N_7762);
and U9570 (N_9570,N_8730,N_8840);
nor U9571 (N_9571,N_7744,N_8109);
nand U9572 (N_9572,N_8644,N_8056);
nor U9573 (N_9573,N_7721,N_8147);
nor U9574 (N_9574,N_8896,N_7670);
and U9575 (N_9575,N_8266,N_8314);
or U9576 (N_9576,N_8475,N_7587);
nand U9577 (N_9577,N_7810,N_8721);
or U9578 (N_9578,N_8737,N_8915);
nor U9579 (N_9579,N_8501,N_8023);
nor U9580 (N_9580,N_8344,N_7962);
nor U9581 (N_9581,N_8258,N_8443);
and U9582 (N_9582,N_8952,N_7654);
nor U9583 (N_9583,N_8117,N_8259);
or U9584 (N_9584,N_8215,N_8083);
xor U9585 (N_9585,N_8346,N_8184);
or U9586 (N_9586,N_8155,N_7763);
xor U9587 (N_9587,N_8526,N_8436);
xnor U9588 (N_9588,N_8474,N_8551);
xor U9589 (N_9589,N_8234,N_8059);
nor U9590 (N_9590,N_8188,N_8536);
and U9591 (N_9591,N_8418,N_8296);
and U9592 (N_9592,N_8048,N_8878);
and U9593 (N_9593,N_8719,N_8856);
nor U9594 (N_9594,N_7933,N_8489);
or U9595 (N_9595,N_8701,N_8827);
or U9596 (N_9596,N_8979,N_7520);
or U9597 (N_9597,N_7567,N_8925);
nand U9598 (N_9598,N_7854,N_8377);
or U9599 (N_9599,N_8086,N_7604);
nor U9600 (N_9600,N_8472,N_8980);
or U9601 (N_9601,N_8766,N_7875);
or U9602 (N_9602,N_7709,N_8387);
or U9603 (N_9603,N_8165,N_8553);
nor U9604 (N_9604,N_8963,N_8902);
and U9605 (N_9605,N_8177,N_7987);
and U9606 (N_9606,N_8975,N_8173);
xnor U9607 (N_9607,N_7708,N_8265);
xnor U9608 (N_9608,N_8403,N_8854);
and U9609 (N_9609,N_8055,N_8254);
nand U9610 (N_9610,N_8283,N_7656);
xor U9611 (N_9611,N_8009,N_8799);
xnor U9612 (N_9612,N_7531,N_8492);
and U9613 (N_9613,N_7832,N_8534);
nor U9614 (N_9614,N_8310,N_8589);
and U9615 (N_9615,N_7607,N_7831);
and U9616 (N_9616,N_8399,N_8794);
or U9617 (N_9617,N_8609,N_8099);
or U9618 (N_9618,N_8246,N_8927);
or U9619 (N_9619,N_7993,N_8720);
nand U9620 (N_9620,N_7575,N_8160);
nor U9621 (N_9621,N_7588,N_7863);
and U9622 (N_9622,N_7759,N_8770);
nor U9623 (N_9623,N_7715,N_8193);
or U9624 (N_9624,N_7995,N_8304);
nand U9625 (N_9625,N_8640,N_8829);
nor U9626 (N_9626,N_8929,N_8875);
or U9627 (N_9627,N_7728,N_8823);
nor U9628 (N_9628,N_8563,N_8350);
nor U9629 (N_9629,N_7669,N_8732);
nor U9630 (N_9630,N_8449,N_8157);
or U9631 (N_9631,N_8168,N_7518);
nor U9632 (N_9632,N_8859,N_7928);
or U9633 (N_9633,N_8722,N_8670);
xnor U9634 (N_9634,N_8990,N_7608);
xor U9635 (N_9635,N_8456,N_8028);
nor U9636 (N_9636,N_7873,N_8444);
xnor U9637 (N_9637,N_8626,N_8582);
or U9638 (N_9638,N_7976,N_8114);
and U9639 (N_9639,N_7515,N_7861);
nand U9640 (N_9640,N_7706,N_8678);
nand U9641 (N_9641,N_7512,N_8655);
nor U9642 (N_9642,N_7733,N_8788);
nand U9643 (N_9643,N_8178,N_8129);
xnor U9644 (N_9644,N_7690,N_7882);
nor U9645 (N_9645,N_7571,N_8705);
or U9646 (N_9646,N_8320,N_7883);
xor U9647 (N_9647,N_8256,N_8402);
xor U9648 (N_9648,N_8151,N_7800);
xor U9649 (N_9649,N_8604,N_8522);
and U9650 (N_9650,N_8985,N_8476);
or U9651 (N_9651,N_8172,N_7742);
nand U9652 (N_9652,N_8619,N_7872);
or U9653 (N_9653,N_7677,N_7500);
nand U9654 (N_9654,N_8749,N_8122);
and U9655 (N_9655,N_7856,N_8139);
nor U9656 (N_9656,N_8738,N_8276);
or U9657 (N_9657,N_8153,N_8213);
nor U9658 (N_9658,N_8792,N_7829);
nor U9659 (N_9659,N_7813,N_8894);
and U9660 (N_9660,N_8740,N_7647);
or U9661 (N_9661,N_8222,N_8950);
and U9662 (N_9662,N_8362,N_8481);
or U9663 (N_9663,N_8690,N_8943);
and U9664 (N_9664,N_7984,N_8496);
or U9665 (N_9665,N_8303,N_8208);
or U9666 (N_9666,N_8949,N_8272);
nor U9667 (N_9667,N_7650,N_7879);
and U9668 (N_9668,N_7523,N_8284);
or U9669 (N_9669,N_8529,N_7950);
nand U9670 (N_9670,N_8629,N_8511);
nor U9671 (N_9671,N_8597,N_8865);
and U9672 (N_9672,N_8852,N_8986);
nand U9673 (N_9673,N_8106,N_7707);
or U9674 (N_9674,N_8581,N_7685);
xor U9675 (N_9675,N_7791,N_8863);
xor U9676 (N_9676,N_8071,N_8791);
or U9677 (N_9677,N_7717,N_7581);
xor U9678 (N_9678,N_7899,N_7516);
or U9679 (N_9679,N_8490,N_8965);
xor U9680 (N_9680,N_8409,N_8459);
xnor U9681 (N_9681,N_8954,N_8731);
xnor U9682 (N_9682,N_7874,N_8450);
and U9683 (N_9683,N_7574,N_8824);
nor U9684 (N_9684,N_8916,N_8781);
or U9685 (N_9685,N_7845,N_8672);
nand U9686 (N_9686,N_8812,N_7998);
or U9687 (N_9687,N_7569,N_7596);
xnor U9688 (N_9688,N_7949,N_8620);
or U9689 (N_9689,N_8163,N_8621);
and U9690 (N_9690,N_7758,N_7910);
nand U9691 (N_9691,N_8939,N_8478);
xnor U9692 (N_9692,N_8176,N_7692);
nor U9693 (N_9693,N_7507,N_8631);
nor U9694 (N_9694,N_7796,N_8212);
xnor U9695 (N_9695,N_7954,N_8578);
nor U9696 (N_9696,N_8198,N_8795);
nor U9697 (N_9697,N_8135,N_8637);
and U9698 (N_9698,N_7615,N_8942);
nand U9699 (N_9699,N_8785,N_8074);
or U9700 (N_9700,N_8886,N_8641);
and U9701 (N_9701,N_8517,N_8716);
nor U9702 (N_9702,N_7807,N_8972);
and U9703 (N_9703,N_7659,N_7508);
nor U9704 (N_9704,N_8997,N_8808);
or U9705 (N_9705,N_8652,N_8088);
or U9706 (N_9706,N_8944,N_8611);
xor U9707 (N_9707,N_8685,N_8473);
nand U9708 (N_9708,N_8333,N_7641);
or U9709 (N_9709,N_8885,N_8181);
nor U9710 (N_9710,N_8767,N_8041);
and U9711 (N_9711,N_7991,N_8119);
xor U9712 (N_9712,N_8901,N_8613);
nor U9713 (N_9713,N_8707,N_7612);
nor U9714 (N_9714,N_8174,N_8879);
xor U9715 (N_9715,N_8493,N_8364);
nand U9716 (N_9716,N_8904,N_8206);
or U9717 (N_9717,N_8595,N_8390);
nor U9718 (N_9718,N_8158,N_8541);
and U9719 (N_9719,N_7973,N_7957);
nor U9720 (N_9720,N_8392,N_8610);
nor U9721 (N_9721,N_7850,N_8510);
or U9722 (N_9722,N_8438,N_8034);
or U9723 (N_9723,N_8649,N_7609);
nand U9724 (N_9724,N_8783,N_8523);
nor U9725 (N_9725,N_7542,N_8703);
nand U9726 (N_9726,N_8834,N_8495);
nor U9727 (N_9727,N_8428,N_8970);
nor U9728 (N_9728,N_8345,N_8769);
or U9729 (N_9729,N_8226,N_7946);
and U9730 (N_9730,N_8483,N_8691);
nand U9731 (N_9731,N_7776,N_7802);
xor U9732 (N_9732,N_8464,N_8742);
nor U9733 (N_9733,N_7745,N_8787);
or U9734 (N_9734,N_7869,N_8587);
or U9735 (N_9735,N_7617,N_8216);
xnor U9736 (N_9736,N_8285,N_7686);
xor U9737 (N_9737,N_7890,N_7713);
and U9738 (N_9738,N_7751,N_8561);
or U9739 (N_9739,N_8555,N_8648);
nor U9740 (N_9740,N_8214,N_7880);
nand U9741 (N_9741,N_8771,N_7586);
nor U9742 (N_9742,N_8025,N_7887);
or U9743 (N_9743,N_7638,N_8584);
and U9744 (N_9744,N_7999,N_8388);
or U9745 (N_9745,N_8679,N_8035);
nor U9746 (N_9746,N_7620,N_8209);
nor U9747 (N_9747,N_7551,N_8191);
nor U9748 (N_9748,N_8415,N_7778);
nor U9749 (N_9749,N_7753,N_7814);
or U9750 (N_9750,N_8503,N_7694);
or U9751 (N_9751,N_7505,N_8946);
nand U9752 (N_9752,N_8123,N_8574);
xnor U9753 (N_9753,N_8786,N_8398);
nor U9754 (N_9754,N_8726,N_8243);
or U9755 (N_9755,N_8388,N_8122);
or U9756 (N_9756,N_7989,N_8418);
nand U9757 (N_9757,N_8278,N_7827);
nand U9758 (N_9758,N_8893,N_7636);
or U9759 (N_9759,N_8624,N_8442);
and U9760 (N_9760,N_7944,N_8629);
and U9761 (N_9761,N_8707,N_7516);
nor U9762 (N_9762,N_8677,N_8423);
nor U9763 (N_9763,N_8868,N_7590);
nor U9764 (N_9764,N_8935,N_8249);
xor U9765 (N_9765,N_8522,N_8533);
nor U9766 (N_9766,N_8962,N_8879);
nor U9767 (N_9767,N_8989,N_8529);
nand U9768 (N_9768,N_8441,N_8757);
nand U9769 (N_9769,N_7823,N_8316);
xnor U9770 (N_9770,N_8679,N_7707);
nand U9771 (N_9771,N_7677,N_8306);
xnor U9772 (N_9772,N_8187,N_8253);
xnor U9773 (N_9773,N_8702,N_7811);
nor U9774 (N_9774,N_8582,N_7736);
nand U9775 (N_9775,N_8171,N_7760);
and U9776 (N_9776,N_7882,N_8720);
nor U9777 (N_9777,N_7812,N_8069);
or U9778 (N_9778,N_8824,N_8601);
nand U9779 (N_9779,N_8744,N_8731);
nor U9780 (N_9780,N_8248,N_7787);
and U9781 (N_9781,N_8249,N_7593);
nand U9782 (N_9782,N_7630,N_8037);
or U9783 (N_9783,N_7732,N_7952);
or U9784 (N_9784,N_7855,N_8497);
xor U9785 (N_9785,N_7795,N_8454);
and U9786 (N_9786,N_8256,N_8705);
xnor U9787 (N_9787,N_8693,N_8575);
and U9788 (N_9788,N_8509,N_7566);
xor U9789 (N_9789,N_8868,N_7935);
or U9790 (N_9790,N_8170,N_8779);
xnor U9791 (N_9791,N_8699,N_7647);
xnor U9792 (N_9792,N_7721,N_8998);
nand U9793 (N_9793,N_8627,N_7687);
and U9794 (N_9794,N_8185,N_7780);
nand U9795 (N_9795,N_8444,N_8842);
nand U9796 (N_9796,N_8947,N_8379);
xor U9797 (N_9797,N_7828,N_8748);
nor U9798 (N_9798,N_8066,N_8834);
or U9799 (N_9799,N_7596,N_8055);
or U9800 (N_9800,N_8808,N_7788);
and U9801 (N_9801,N_7504,N_8998);
nand U9802 (N_9802,N_7703,N_8603);
nor U9803 (N_9803,N_7586,N_7958);
xor U9804 (N_9804,N_8139,N_8820);
or U9805 (N_9805,N_8410,N_8526);
nor U9806 (N_9806,N_8624,N_8492);
nand U9807 (N_9807,N_8001,N_8948);
nor U9808 (N_9808,N_8410,N_8508);
nor U9809 (N_9809,N_7883,N_8247);
and U9810 (N_9810,N_8933,N_7646);
nand U9811 (N_9811,N_8502,N_8930);
or U9812 (N_9812,N_7865,N_8542);
xor U9813 (N_9813,N_8649,N_7608);
nor U9814 (N_9814,N_7759,N_8567);
and U9815 (N_9815,N_8914,N_7730);
nand U9816 (N_9816,N_8459,N_7603);
or U9817 (N_9817,N_8839,N_8382);
and U9818 (N_9818,N_8213,N_8467);
xor U9819 (N_9819,N_8163,N_8667);
and U9820 (N_9820,N_8982,N_8445);
xnor U9821 (N_9821,N_8210,N_7975);
xor U9822 (N_9822,N_8944,N_8104);
and U9823 (N_9823,N_8662,N_7803);
nor U9824 (N_9824,N_8999,N_8900);
xor U9825 (N_9825,N_8159,N_8170);
nor U9826 (N_9826,N_8126,N_8029);
and U9827 (N_9827,N_8857,N_8816);
nand U9828 (N_9828,N_8385,N_8413);
nor U9829 (N_9829,N_8610,N_7655);
or U9830 (N_9830,N_8093,N_8260);
or U9831 (N_9831,N_8782,N_8920);
nand U9832 (N_9832,N_7858,N_7507);
nor U9833 (N_9833,N_8370,N_7859);
nand U9834 (N_9834,N_7714,N_7773);
or U9835 (N_9835,N_7555,N_7575);
or U9836 (N_9836,N_7938,N_8835);
nand U9837 (N_9837,N_8541,N_8670);
xnor U9838 (N_9838,N_8252,N_8869);
and U9839 (N_9839,N_8133,N_8681);
nor U9840 (N_9840,N_8276,N_8549);
nand U9841 (N_9841,N_8927,N_7785);
nor U9842 (N_9842,N_8933,N_8734);
xnor U9843 (N_9843,N_7838,N_7733);
nand U9844 (N_9844,N_8268,N_8055);
nor U9845 (N_9845,N_8798,N_8396);
or U9846 (N_9846,N_7610,N_8563);
nand U9847 (N_9847,N_8634,N_8748);
nand U9848 (N_9848,N_7529,N_7828);
xnor U9849 (N_9849,N_8346,N_8920);
or U9850 (N_9850,N_7931,N_8017);
nand U9851 (N_9851,N_7831,N_7645);
nor U9852 (N_9852,N_7776,N_7679);
and U9853 (N_9853,N_7849,N_8695);
xor U9854 (N_9854,N_8592,N_7727);
and U9855 (N_9855,N_8176,N_8390);
xnor U9856 (N_9856,N_8341,N_8725);
and U9857 (N_9857,N_8126,N_8746);
and U9858 (N_9858,N_8727,N_8415);
or U9859 (N_9859,N_8742,N_7955);
xnor U9860 (N_9860,N_8303,N_8144);
and U9861 (N_9861,N_8323,N_8595);
and U9862 (N_9862,N_7741,N_8757);
nor U9863 (N_9863,N_8090,N_8235);
and U9864 (N_9864,N_8174,N_8559);
or U9865 (N_9865,N_8613,N_8701);
xor U9866 (N_9866,N_8711,N_8583);
and U9867 (N_9867,N_8900,N_7725);
nor U9868 (N_9868,N_7866,N_8572);
nor U9869 (N_9869,N_7738,N_8848);
xnor U9870 (N_9870,N_8598,N_7819);
and U9871 (N_9871,N_7656,N_8635);
and U9872 (N_9872,N_8783,N_8146);
nor U9873 (N_9873,N_7922,N_8847);
or U9874 (N_9874,N_7545,N_8932);
nand U9875 (N_9875,N_7631,N_8893);
xnor U9876 (N_9876,N_8424,N_8490);
and U9877 (N_9877,N_8546,N_8216);
and U9878 (N_9878,N_8431,N_8398);
nand U9879 (N_9879,N_8830,N_8451);
nor U9880 (N_9880,N_7850,N_8519);
nand U9881 (N_9881,N_8292,N_7792);
or U9882 (N_9882,N_8141,N_8492);
nand U9883 (N_9883,N_8353,N_8959);
xor U9884 (N_9884,N_8184,N_8964);
xnor U9885 (N_9885,N_8272,N_8521);
nor U9886 (N_9886,N_8182,N_8049);
xnor U9887 (N_9887,N_7966,N_8121);
nand U9888 (N_9888,N_7605,N_7786);
or U9889 (N_9889,N_8664,N_8982);
nand U9890 (N_9890,N_7880,N_8358);
and U9891 (N_9891,N_8669,N_8629);
nand U9892 (N_9892,N_8263,N_8737);
and U9893 (N_9893,N_8748,N_7829);
xnor U9894 (N_9894,N_8137,N_7870);
xnor U9895 (N_9895,N_8249,N_7646);
or U9896 (N_9896,N_8329,N_8021);
xor U9897 (N_9897,N_8785,N_7563);
xor U9898 (N_9898,N_7888,N_8575);
nor U9899 (N_9899,N_7722,N_8381);
xnor U9900 (N_9900,N_7952,N_7631);
xnor U9901 (N_9901,N_8670,N_8126);
or U9902 (N_9902,N_8266,N_8197);
or U9903 (N_9903,N_7787,N_7923);
and U9904 (N_9904,N_8882,N_7741);
or U9905 (N_9905,N_7656,N_8131);
nand U9906 (N_9906,N_8694,N_7771);
or U9907 (N_9907,N_7549,N_7671);
or U9908 (N_9908,N_8329,N_8145);
xor U9909 (N_9909,N_8854,N_8112);
xor U9910 (N_9910,N_7873,N_8651);
xnor U9911 (N_9911,N_8130,N_7677);
or U9912 (N_9912,N_7748,N_8724);
or U9913 (N_9913,N_8678,N_8232);
and U9914 (N_9914,N_8743,N_8784);
xor U9915 (N_9915,N_8369,N_7913);
nand U9916 (N_9916,N_8022,N_7779);
nand U9917 (N_9917,N_8679,N_8845);
xor U9918 (N_9918,N_8489,N_8092);
or U9919 (N_9919,N_8562,N_8504);
and U9920 (N_9920,N_7697,N_8163);
nor U9921 (N_9921,N_7570,N_7625);
and U9922 (N_9922,N_7538,N_7948);
nor U9923 (N_9923,N_8440,N_8584);
xor U9924 (N_9924,N_7904,N_8344);
and U9925 (N_9925,N_7687,N_8301);
xnor U9926 (N_9926,N_8383,N_7978);
nand U9927 (N_9927,N_7939,N_8626);
and U9928 (N_9928,N_7765,N_8624);
nand U9929 (N_9929,N_8228,N_8807);
and U9930 (N_9930,N_8638,N_7625);
or U9931 (N_9931,N_7967,N_8858);
nor U9932 (N_9932,N_7539,N_8648);
nand U9933 (N_9933,N_8443,N_8015);
nand U9934 (N_9934,N_8530,N_8972);
nor U9935 (N_9935,N_8793,N_7939);
xor U9936 (N_9936,N_8656,N_8600);
xnor U9937 (N_9937,N_8006,N_7836);
and U9938 (N_9938,N_8926,N_8780);
xnor U9939 (N_9939,N_7700,N_7814);
or U9940 (N_9940,N_8136,N_7803);
nand U9941 (N_9941,N_8841,N_7853);
xnor U9942 (N_9942,N_8963,N_7716);
nor U9943 (N_9943,N_8087,N_8889);
and U9944 (N_9944,N_8593,N_8910);
or U9945 (N_9945,N_7756,N_8638);
or U9946 (N_9946,N_7873,N_8643);
nor U9947 (N_9947,N_8697,N_7782);
or U9948 (N_9948,N_8457,N_8774);
xnor U9949 (N_9949,N_8820,N_8299);
xor U9950 (N_9950,N_7956,N_8102);
or U9951 (N_9951,N_7884,N_7598);
nand U9952 (N_9952,N_7957,N_7844);
and U9953 (N_9953,N_7577,N_7623);
and U9954 (N_9954,N_8654,N_8101);
and U9955 (N_9955,N_8245,N_8418);
or U9956 (N_9956,N_8295,N_7521);
xor U9957 (N_9957,N_7659,N_8033);
nand U9958 (N_9958,N_8343,N_8833);
or U9959 (N_9959,N_7911,N_8895);
nor U9960 (N_9960,N_7764,N_7915);
and U9961 (N_9961,N_8751,N_8872);
or U9962 (N_9962,N_8579,N_8666);
nand U9963 (N_9963,N_7966,N_8966);
nor U9964 (N_9964,N_7766,N_8061);
nand U9965 (N_9965,N_8528,N_8031);
nand U9966 (N_9966,N_7725,N_7773);
nand U9967 (N_9967,N_8947,N_7981);
or U9968 (N_9968,N_7957,N_8889);
xnor U9969 (N_9969,N_7648,N_7880);
nor U9970 (N_9970,N_8140,N_8632);
and U9971 (N_9971,N_8928,N_8772);
or U9972 (N_9972,N_8584,N_8182);
nor U9973 (N_9973,N_7743,N_8404);
nand U9974 (N_9974,N_8580,N_8372);
xnor U9975 (N_9975,N_8416,N_8406);
or U9976 (N_9976,N_8240,N_8014);
and U9977 (N_9977,N_8718,N_7813);
nor U9978 (N_9978,N_7786,N_8258);
nand U9979 (N_9979,N_7697,N_7918);
or U9980 (N_9980,N_8785,N_7683);
xnor U9981 (N_9981,N_7904,N_7928);
nor U9982 (N_9982,N_8054,N_7903);
xnor U9983 (N_9983,N_8479,N_7946);
xnor U9984 (N_9984,N_8529,N_8746);
nand U9985 (N_9985,N_8527,N_8300);
or U9986 (N_9986,N_7608,N_8843);
nand U9987 (N_9987,N_8149,N_8744);
nor U9988 (N_9988,N_8091,N_7729);
and U9989 (N_9989,N_8778,N_8414);
and U9990 (N_9990,N_7626,N_7848);
and U9991 (N_9991,N_8385,N_8355);
xnor U9992 (N_9992,N_8340,N_8994);
or U9993 (N_9993,N_7758,N_8217);
xor U9994 (N_9994,N_8336,N_7672);
xor U9995 (N_9995,N_8174,N_8830);
and U9996 (N_9996,N_8370,N_7652);
and U9997 (N_9997,N_8013,N_7939);
and U9998 (N_9998,N_8208,N_8137);
nand U9999 (N_9999,N_8816,N_8098);
or U10000 (N_10000,N_8971,N_8097);
and U10001 (N_10001,N_7923,N_8037);
nand U10002 (N_10002,N_7824,N_8340);
and U10003 (N_10003,N_7793,N_8797);
nand U10004 (N_10004,N_7854,N_8200);
and U10005 (N_10005,N_8503,N_8975);
or U10006 (N_10006,N_8470,N_7590);
or U10007 (N_10007,N_8179,N_7808);
nand U10008 (N_10008,N_8940,N_8297);
and U10009 (N_10009,N_8960,N_7983);
or U10010 (N_10010,N_8531,N_8565);
or U10011 (N_10011,N_7820,N_8234);
nand U10012 (N_10012,N_8360,N_7697);
and U10013 (N_10013,N_8772,N_8909);
or U10014 (N_10014,N_7596,N_7692);
or U10015 (N_10015,N_8913,N_8996);
and U10016 (N_10016,N_8438,N_8352);
nor U10017 (N_10017,N_7553,N_8120);
nand U10018 (N_10018,N_8312,N_8722);
xnor U10019 (N_10019,N_8403,N_7540);
nand U10020 (N_10020,N_8899,N_8456);
or U10021 (N_10021,N_7619,N_8437);
and U10022 (N_10022,N_8976,N_8396);
xnor U10023 (N_10023,N_8971,N_7752);
nand U10024 (N_10024,N_7930,N_8398);
nand U10025 (N_10025,N_8748,N_7996);
and U10026 (N_10026,N_7816,N_7576);
or U10027 (N_10027,N_7922,N_8671);
nand U10028 (N_10028,N_8245,N_8271);
nand U10029 (N_10029,N_8861,N_7635);
nor U10030 (N_10030,N_8427,N_8010);
xor U10031 (N_10031,N_8574,N_8104);
xor U10032 (N_10032,N_8395,N_7573);
nor U10033 (N_10033,N_8239,N_8725);
xor U10034 (N_10034,N_8252,N_8320);
and U10035 (N_10035,N_7954,N_8458);
and U10036 (N_10036,N_7722,N_8717);
or U10037 (N_10037,N_7641,N_8241);
nor U10038 (N_10038,N_7697,N_7704);
nand U10039 (N_10039,N_8617,N_8439);
xor U10040 (N_10040,N_8668,N_8318);
nand U10041 (N_10041,N_8107,N_8275);
and U10042 (N_10042,N_7621,N_7874);
or U10043 (N_10043,N_8859,N_8039);
or U10044 (N_10044,N_8646,N_8121);
nor U10045 (N_10045,N_7823,N_8209);
and U10046 (N_10046,N_7863,N_7906);
nor U10047 (N_10047,N_8260,N_7597);
or U10048 (N_10048,N_8880,N_8452);
and U10049 (N_10049,N_8632,N_8128);
nand U10050 (N_10050,N_7622,N_8354);
nor U10051 (N_10051,N_8055,N_7852);
xnor U10052 (N_10052,N_7656,N_8424);
or U10053 (N_10053,N_8617,N_8272);
xnor U10054 (N_10054,N_8556,N_8896);
and U10055 (N_10055,N_8897,N_8412);
or U10056 (N_10056,N_8049,N_7798);
xnor U10057 (N_10057,N_8164,N_8417);
xor U10058 (N_10058,N_8671,N_7938);
and U10059 (N_10059,N_7754,N_7809);
xor U10060 (N_10060,N_8060,N_8890);
nor U10061 (N_10061,N_8623,N_7646);
or U10062 (N_10062,N_7758,N_7568);
and U10063 (N_10063,N_8259,N_8683);
nor U10064 (N_10064,N_8812,N_8735);
and U10065 (N_10065,N_8301,N_8116);
nor U10066 (N_10066,N_8972,N_8396);
xnor U10067 (N_10067,N_8073,N_8475);
or U10068 (N_10068,N_7999,N_8732);
nand U10069 (N_10069,N_8706,N_7513);
nor U10070 (N_10070,N_8335,N_8305);
nor U10071 (N_10071,N_7571,N_8380);
nor U10072 (N_10072,N_7919,N_7503);
nor U10073 (N_10073,N_7827,N_7877);
nand U10074 (N_10074,N_7914,N_8227);
nor U10075 (N_10075,N_8087,N_8192);
or U10076 (N_10076,N_8922,N_7758);
and U10077 (N_10077,N_7572,N_8093);
and U10078 (N_10078,N_8662,N_8188);
nor U10079 (N_10079,N_8498,N_7970);
and U10080 (N_10080,N_8653,N_7534);
nand U10081 (N_10081,N_7818,N_8543);
nand U10082 (N_10082,N_8281,N_8294);
nand U10083 (N_10083,N_8376,N_7714);
nand U10084 (N_10084,N_8063,N_8502);
or U10085 (N_10085,N_8249,N_8322);
xor U10086 (N_10086,N_8617,N_8973);
nand U10087 (N_10087,N_8472,N_8002);
xnor U10088 (N_10088,N_8612,N_7686);
or U10089 (N_10089,N_7533,N_8197);
nor U10090 (N_10090,N_7770,N_7645);
nand U10091 (N_10091,N_8159,N_8979);
or U10092 (N_10092,N_7985,N_8767);
nand U10093 (N_10093,N_7934,N_8218);
and U10094 (N_10094,N_8901,N_8667);
nand U10095 (N_10095,N_8536,N_7906);
or U10096 (N_10096,N_8259,N_8164);
nor U10097 (N_10097,N_8248,N_8755);
or U10098 (N_10098,N_7698,N_8630);
and U10099 (N_10099,N_8295,N_8660);
nand U10100 (N_10100,N_8918,N_8263);
or U10101 (N_10101,N_8663,N_7751);
and U10102 (N_10102,N_8378,N_7811);
nor U10103 (N_10103,N_8572,N_7738);
and U10104 (N_10104,N_7554,N_7507);
and U10105 (N_10105,N_7756,N_8450);
xnor U10106 (N_10106,N_7860,N_8699);
nor U10107 (N_10107,N_8088,N_8898);
xnor U10108 (N_10108,N_8616,N_7704);
or U10109 (N_10109,N_7812,N_7854);
nor U10110 (N_10110,N_8893,N_8212);
and U10111 (N_10111,N_8387,N_8952);
nand U10112 (N_10112,N_8696,N_8157);
nor U10113 (N_10113,N_8442,N_8164);
nand U10114 (N_10114,N_8904,N_8824);
nor U10115 (N_10115,N_7969,N_8106);
nor U10116 (N_10116,N_8862,N_8596);
and U10117 (N_10117,N_8048,N_8576);
nand U10118 (N_10118,N_8048,N_8570);
or U10119 (N_10119,N_7737,N_8723);
or U10120 (N_10120,N_7672,N_8841);
nand U10121 (N_10121,N_8296,N_8591);
nor U10122 (N_10122,N_8830,N_7542);
xor U10123 (N_10123,N_8793,N_7852);
xnor U10124 (N_10124,N_7660,N_8717);
xor U10125 (N_10125,N_7888,N_8623);
nor U10126 (N_10126,N_8064,N_7623);
nand U10127 (N_10127,N_8240,N_8380);
xor U10128 (N_10128,N_8621,N_7809);
nand U10129 (N_10129,N_8956,N_8270);
or U10130 (N_10130,N_8116,N_8550);
and U10131 (N_10131,N_7966,N_8769);
nor U10132 (N_10132,N_8770,N_8469);
nor U10133 (N_10133,N_8053,N_8303);
nand U10134 (N_10134,N_8907,N_8598);
and U10135 (N_10135,N_8448,N_8806);
or U10136 (N_10136,N_7577,N_8754);
or U10137 (N_10137,N_8437,N_7774);
nand U10138 (N_10138,N_7507,N_8362);
nand U10139 (N_10139,N_8200,N_8360);
nand U10140 (N_10140,N_8440,N_7696);
nor U10141 (N_10141,N_8468,N_8107);
and U10142 (N_10142,N_7618,N_7842);
nor U10143 (N_10143,N_7526,N_8543);
xor U10144 (N_10144,N_8042,N_7818);
nand U10145 (N_10145,N_7895,N_7557);
or U10146 (N_10146,N_8841,N_8956);
xor U10147 (N_10147,N_8968,N_8814);
xor U10148 (N_10148,N_8648,N_8154);
xnor U10149 (N_10149,N_8614,N_7530);
xnor U10150 (N_10150,N_8972,N_8568);
or U10151 (N_10151,N_8029,N_8442);
and U10152 (N_10152,N_8449,N_8855);
nand U10153 (N_10153,N_8549,N_8924);
and U10154 (N_10154,N_7602,N_8373);
xnor U10155 (N_10155,N_8908,N_8774);
and U10156 (N_10156,N_7550,N_7570);
nand U10157 (N_10157,N_7579,N_8260);
and U10158 (N_10158,N_7692,N_8533);
or U10159 (N_10159,N_8863,N_8671);
nand U10160 (N_10160,N_8038,N_8160);
and U10161 (N_10161,N_8162,N_8997);
and U10162 (N_10162,N_7595,N_8232);
xnor U10163 (N_10163,N_8029,N_7578);
xnor U10164 (N_10164,N_8681,N_8242);
nor U10165 (N_10165,N_8315,N_8728);
and U10166 (N_10166,N_8888,N_7695);
xnor U10167 (N_10167,N_8761,N_8941);
xnor U10168 (N_10168,N_8377,N_8909);
xnor U10169 (N_10169,N_8330,N_8904);
nand U10170 (N_10170,N_8149,N_7527);
nor U10171 (N_10171,N_7932,N_7572);
and U10172 (N_10172,N_7621,N_8026);
or U10173 (N_10173,N_7740,N_8377);
xnor U10174 (N_10174,N_7690,N_8441);
nand U10175 (N_10175,N_8505,N_7911);
nand U10176 (N_10176,N_8039,N_7577);
xnor U10177 (N_10177,N_8286,N_7807);
and U10178 (N_10178,N_8443,N_8593);
nand U10179 (N_10179,N_8281,N_8632);
and U10180 (N_10180,N_8881,N_7595);
or U10181 (N_10181,N_8842,N_8607);
nor U10182 (N_10182,N_7508,N_8416);
and U10183 (N_10183,N_8019,N_8868);
or U10184 (N_10184,N_8271,N_7526);
nand U10185 (N_10185,N_7617,N_8046);
or U10186 (N_10186,N_8911,N_8157);
nand U10187 (N_10187,N_8191,N_7680);
and U10188 (N_10188,N_7509,N_8602);
or U10189 (N_10189,N_8939,N_8433);
and U10190 (N_10190,N_8996,N_7775);
nand U10191 (N_10191,N_8814,N_7946);
nand U10192 (N_10192,N_7726,N_8914);
xnor U10193 (N_10193,N_7922,N_8740);
and U10194 (N_10194,N_8530,N_8760);
xnor U10195 (N_10195,N_8740,N_8863);
nor U10196 (N_10196,N_8009,N_8683);
or U10197 (N_10197,N_7921,N_8650);
nor U10198 (N_10198,N_8352,N_8479);
nand U10199 (N_10199,N_8240,N_7690);
and U10200 (N_10200,N_8766,N_7614);
xor U10201 (N_10201,N_8045,N_8984);
nor U10202 (N_10202,N_7719,N_7647);
and U10203 (N_10203,N_8754,N_8623);
nor U10204 (N_10204,N_8630,N_8278);
or U10205 (N_10205,N_8264,N_8801);
and U10206 (N_10206,N_8520,N_7668);
nor U10207 (N_10207,N_7715,N_8549);
nand U10208 (N_10208,N_7550,N_8282);
and U10209 (N_10209,N_8069,N_7751);
nor U10210 (N_10210,N_8527,N_7579);
xor U10211 (N_10211,N_8263,N_7620);
nand U10212 (N_10212,N_7975,N_8850);
nand U10213 (N_10213,N_8589,N_8099);
nor U10214 (N_10214,N_7808,N_8384);
nor U10215 (N_10215,N_8631,N_8572);
or U10216 (N_10216,N_7964,N_8313);
or U10217 (N_10217,N_8733,N_8120);
nand U10218 (N_10218,N_7755,N_7835);
nand U10219 (N_10219,N_8760,N_7708);
nand U10220 (N_10220,N_8985,N_8425);
or U10221 (N_10221,N_8914,N_8427);
or U10222 (N_10222,N_8737,N_8923);
nor U10223 (N_10223,N_8238,N_8788);
xor U10224 (N_10224,N_7978,N_7765);
or U10225 (N_10225,N_8058,N_8613);
nand U10226 (N_10226,N_8058,N_8953);
nor U10227 (N_10227,N_8529,N_7503);
nor U10228 (N_10228,N_7723,N_8298);
or U10229 (N_10229,N_8838,N_7531);
nand U10230 (N_10230,N_8613,N_7500);
nand U10231 (N_10231,N_8468,N_7997);
xor U10232 (N_10232,N_8481,N_8597);
nand U10233 (N_10233,N_7537,N_8418);
and U10234 (N_10234,N_8065,N_8158);
xor U10235 (N_10235,N_8920,N_8889);
nand U10236 (N_10236,N_8010,N_7795);
xnor U10237 (N_10237,N_8842,N_8763);
and U10238 (N_10238,N_7589,N_8247);
and U10239 (N_10239,N_7501,N_8201);
nor U10240 (N_10240,N_7950,N_8914);
nand U10241 (N_10241,N_7644,N_8238);
nor U10242 (N_10242,N_7679,N_8892);
or U10243 (N_10243,N_8579,N_8617);
or U10244 (N_10244,N_8484,N_8264);
xnor U10245 (N_10245,N_7579,N_8951);
xnor U10246 (N_10246,N_8513,N_7993);
nor U10247 (N_10247,N_7563,N_7917);
or U10248 (N_10248,N_8881,N_7610);
or U10249 (N_10249,N_8310,N_8114);
or U10250 (N_10250,N_8983,N_8901);
or U10251 (N_10251,N_7861,N_7986);
and U10252 (N_10252,N_7953,N_7693);
nor U10253 (N_10253,N_8971,N_8747);
xnor U10254 (N_10254,N_8520,N_8884);
or U10255 (N_10255,N_8886,N_7587);
xnor U10256 (N_10256,N_7666,N_8843);
and U10257 (N_10257,N_8214,N_7566);
xnor U10258 (N_10258,N_8403,N_8879);
nand U10259 (N_10259,N_8335,N_8469);
or U10260 (N_10260,N_8380,N_7787);
nor U10261 (N_10261,N_8410,N_8603);
nor U10262 (N_10262,N_7919,N_8373);
nand U10263 (N_10263,N_7763,N_8312);
nand U10264 (N_10264,N_8917,N_7900);
nor U10265 (N_10265,N_8048,N_8069);
or U10266 (N_10266,N_8025,N_8833);
nor U10267 (N_10267,N_8739,N_8854);
nor U10268 (N_10268,N_8752,N_7650);
or U10269 (N_10269,N_7738,N_8818);
or U10270 (N_10270,N_8811,N_8550);
or U10271 (N_10271,N_7778,N_7781);
or U10272 (N_10272,N_8738,N_8656);
and U10273 (N_10273,N_8395,N_8191);
nor U10274 (N_10274,N_8960,N_8456);
or U10275 (N_10275,N_8895,N_8300);
or U10276 (N_10276,N_7614,N_7505);
nand U10277 (N_10277,N_8099,N_7866);
or U10278 (N_10278,N_8929,N_7861);
nand U10279 (N_10279,N_7982,N_8671);
nand U10280 (N_10280,N_8045,N_8712);
nor U10281 (N_10281,N_8878,N_8947);
nand U10282 (N_10282,N_8300,N_7718);
nand U10283 (N_10283,N_8093,N_8583);
xor U10284 (N_10284,N_8730,N_7682);
nand U10285 (N_10285,N_8641,N_7885);
nor U10286 (N_10286,N_7733,N_7960);
nand U10287 (N_10287,N_8114,N_8999);
nand U10288 (N_10288,N_8141,N_8104);
nor U10289 (N_10289,N_8543,N_7532);
or U10290 (N_10290,N_8153,N_8491);
nor U10291 (N_10291,N_7770,N_8535);
xor U10292 (N_10292,N_7976,N_8517);
xor U10293 (N_10293,N_7779,N_7799);
xor U10294 (N_10294,N_8409,N_7572);
nand U10295 (N_10295,N_7516,N_8619);
nor U10296 (N_10296,N_8349,N_7662);
xor U10297 (N_10297,N_7844,N_8135);
or U10298 (N_10298,N_7630,N_7964);
and U10299 (N_10299,N_8791,N_7547);
and U10300 (N_10300,N_8153,N_8707);
nor U10301 (N_10301,N_7881,N_7813);
or U10302 (N_10302,N_8317,N_8045);
or U10303 (N_10303,N_8705,N_8672);
nor U10304 (N_10304,N_8496,N_8486);
nand U10305 (N_10305,N_8243,N_8121);
or U10306 (N_10306,N_8432,N_8069);
nor U10307 (N_10307,N_8530,N_8546);
and U10308 (N_10308,N_8330,N_8789);
xor U10309 (N_10309,N_7646,N_7947);
or U10310 (N_10310,N_8737,N_8654);
nand U10311 (N_10311,N_8117,N_8658);
and U10312 (N_10312,N_7601,N_7580);
nand U10313 (N_10313,N_8779,N_7901);
nor U10314 (N_10314,N_8151,N_7996);
or U10315 (N_10315,N_7825,N_8909);
nand U10316 (N_10316,N_8664,N_7600);
and U10317 (N_10317,N_8131,N_8838);
nor U10318 (N_10318,N_7590,N_8902);
or U10319 (N_10319,N_8621,N_8486);
and U10320 (N_10320,N_7875,N_7721);
nand U10321 (N_10321,N_8749,N_8588);
and U10322 (N_10322,N_7772,N_7823);
xnor U10323 (N_10323,N_8764,N_8786);
or U10324 (N_10324,N_7901,N_8689);
nor U10325 (N_10325,N_8075,N_7694);
xnor U10326 (N_10326,N_8261,N_8271);
xnor U10327 (N_10327,N_7978,N_7785);
and U10328 (N_10328,N_8768,N_8230);
nand U10329 (N_10329,N_7891,N_7697);
xnor U10330 (N_10330,N_7643,N_8352);
and U10331 (N_10331,N_8411,N_7516);
or U10332 (N_10332,N_8272,N_8847);
and U10333 (N_10333,N_7874,N_8500);
and U10334 (N_10334,N_7789,N_7650);
or U10335 (N_10335,N_8443,N_8159);
xor U10336 (N_10336,N_7680,N_8450);
or U10337 (N_10337,N_8488,N_8655);
or U10338 (N_10338,N_8935,N_7863);
or U10339 (N_10339,N_8777,N_8080);
nand U10340 (N_10340,N_7830,N_8624);
nand U10341 (N_10341,N_8745,N_8978);
nand U10342 (N_10342,N_7536,N_7540);
or U10343 (N_10343,N_8145,N_8573);
nand U10344 (N_10344,N_8429,N_8922);
and U10345 (N_10345,N_7746,N_8160);
or U10346 (N_10346,N_7882,N_8593);
and U10347 (N_10347,N_7524,N_7541);
nand U10348 (N_10348,N_8905,N_7627);
xnor U10349 (N_10349,N_7857,N_8136);
nor U10350 (N_10350,N_7726,N_8304);
nand U10351 (N_10351,N_8770,N_8253);
or U10352 (N_10352,N_8364,N_8554);
nand U10353 (N_10353,N_8596,N_8543);
nand U10354 (N_10354,N_8878,N_7533);
and U10355 (N_10355,N_8124,N_7532);
or U10356 (N_10356,N_8550,N_8737);
or U10357 (N_10357,N_7615,N_8586);
nor U10358 (N_10358,N_7871,N_8847);
nand U10359 (N_10359,N_8810,N_8605);
and U10360 (N_10360,N_8142,N_8930);
or U10361 (N_10361,N_7831,N_7727);
nor U10362 (N_10362,N_7792,N_7772);
xnor U10363 (N_10363,N_8261,N_8275);
xnor U10364 (N_10364,N_8904,N_8635);
nand U10365 (N_10365,N_8735,N_7733);
or U10366 (N_10366,N_8291,N_8135);
nor U10367 (N_10367,N_7710,N_8673);
nor U10368 (N_10368,N_8815,N_7882);
or U10369 (N_10369,N_7752,N_7643);
and U10370 (N_10370,N_8230,N_7515);
nand U10371 (N_10371,N_8537,N_8692);
or U10372 (N_10372,N_8807,N_8027);
or U10373 (N_10373,N_8401,N_8026);
nor U10374 (N_10374,N_7503,N_8286);
xnor U10375 (N_10375,N_8549,N_8294);
xor U10376 (N_10376,N_8657,N_8530);
nor U10377 (N_10377,N_8486,N_7526);
and U10378 (N_10378,N_7840,N_8930);
nand U10379 (N_10379,N_8885,N_7911);
nor U10380 (N_10380,N_7760,N_8004);
nor U10381 (N_10381,N_8712,N_8459);
and U10382 (N_10382,N_8636,N_8052);
nand U10383 (N_10383,N_7661,N_8482);
and U10384 (N_10384,N_7883,N_7557);
xnor U10385 (N_10385,N_7662,N_7725);
xnor U10386 (N_10386,N_8370,N_8970);
and U10387 (N_10387,N_8109,N_7739);
nor U10388 (N_10388,N_8317,N_8184);
or U10389 (N_10389,N_8850,N_8647);
nor U10390 (N_10390,N_8599,N_8202);
or U10391 (N_10391,N_8954,N_8029);
and U10392 (N_10392,N_7792,N_7710);
nand U10393 (N_10393,N_8941,N_7918);
and U10394 (N_10394,N_7861,N_8830);
nand U10395 (N_10395,N_8576,N_8311);
or U10396 (N_10396,N_7595,N_8514);
and U10397 (N_10397,N_8066,N_7650);
nand U10398 (N_10398,N_8456,N_8194);
nor U10399 (N_10399,N_8802,N_8135);
and U10400 (N_10400,N_8137,N_7955);
xor U10401 (N_10401,N_8055,N_8999);
nor U10402 (N_10402,N_7737,N_8719);
or U10403 (N_10403,N_7772,N_8903);
nor U10404 (N_10404,N_7827,N_8048);
or U10405 (N_10405,N_8172,N_8603);
or U10406 (N_10406,N_8380,N_8271);
nand U10407 (N_10407,N_7899,N_7629);
and U10408 (N_10408,N_8587,N_8085);
or U10409 (N_10409,N_7988,N_8882);
nor U10410 (N_10410,N_8746,N_8409);
and U10411 (N_10411,N_8909,N_8090);
nor U10412 (N_10412,N_7854,N_8645);
nand U10413 (N_10413,N_8259,N_8285);
nand U10414 (N_10414,N_8777,N_7504);
nand U10415 (N_10415,N_8120,N_8014);
nand U10416 (N_10416,N_7831,N_7691);
nor U10417 (N_10417,N_7885,N_8374);
and U10418 (N_10418,N_8413,N_8623);
nor U10419 (N_10419,N_8928,N_8388);
nor U10420 (N_10420,N_8907,N_8472);
or U10421 (N_10421,N_7845,N_7504);
nor U10422 (N_10422,N_8756,N_8622);
nor U10423 (N_10423,N_8973,N_8994);
xnor U10424 (N_10424,N_8149,N_8070);
or U10425 (N_10425,N_8239,N_7736);
or U10426 (N_10426,N_8892,N_8135);
nor U10427 (N_10427,N_7645,N_8006);
nor U10428 (N_10428,N_8455,N_8412);
and U10429 (N_10429,N_7771,N_7518);
nor U10430 (N_10430,N_8149,N_8645);
xnor U10431 (N_10431,N_8563,N_8539);
xnor U10432 (N_10432,N_7844,N_7905);
nor U10433 (N_10433,N_8864,N_8702);
xnor U10434 (N_10434,N_7771,N_7833);
and U10435 (N_10435,N_8564,N_8394);
and U10436 (N_10436,N_8735,N_7851);
and U10437 (N_10437,N_8454,N_7759);
or U10438 (N_10438,N_7920,N_7560);
nand U10439 (N_10439,N_8625,N_8189);
and U10440 (N_10440,N_8501,N_7680);
nand U10441 (N_10441,N_8227,N_8377);
and U10442 (N_10442,N_8919,N_8283);
and U10443 (N_10443,N_7755,N_8820);
and U10444 (N_10444,N_8549,N_7532);
nand U10445 (N_10445,N_8680,N_8176);
and U10446 (N_10446,N_8332,N_7814);
nor U10447 (N_10447,N_8792,N_7812);
nor U10448 (N_10448,N_7880,N_8131);
nand U10449 (N_10449,N_8023,N_8654);
and U10450 (N_10450,N_8844,N_8522);
or U10451 (N_10451,N_8253,N_8912);
nand U10452 (N_10452,N_8252,N_7772);
nand U10453 (N_10453,N_8631,N_8528);
nor U10454 (N_10454,N_8803,N_7782);
or U10455 (N_10455,N_7928,N_7999);
xor U10456 (N_10456,N_8214,N_7847);
nand U10457 (N_10457,N_8315,N_8011);
nand U10458 (N_10458,N_7833,N_8054);
xor U10459 (N_10459,N_7694,N_8279);
nor U10460 (N_10460,N_8712,N_7507);
xor U10461 (N_10461,N_8043,N_7989);
nand U10462 (N_10462,N_8930,N_7986);
or U10463 (N_10463,N_7972,N_8307);
and U10464 (N_10464,N_8096,N_7549);
nor U10465 (N_10465,N_8320,N_8841);
nor U10466 (N_10466,N_8185,N_8280);
nand U10467 (N_10467,N_7663,N_8483);
nand U10468 (N_10468,N_8012,N_8016);
nor U10469 (N_10469,N_7806,N_8859);
nand U10470 (N_10470,N_8396,N_8006);
xor U10471 (N_10471,N_8848,N_8640);
xor U10472 (N_10472,N_8046,N_7528);
nand U10473 (N_10473,N_8659,N_8971);
xnor U10474 (N_10474,N_8085,N_8398);
nand U10475 (N_10475,N_8950,N_8163);
nor U10476 (N_10476,N_7526,N_8569);
xnor U10477 (N_10477,N_7582,N_7529);
nand U10478 (N_10478,N_7694,N_8807);
nor U10479 (N_10479,N_7646,N_8024);
xor U10480 (N_10480,N_7894,N_7659);
and U10481 (N_10481,N_8898,N_7736);
nand U10482 (N_10482,N_8615,N_8445);
nor U10483 (N_10483,N_7513,N_8931);
xor U10484 (N_10484,N_8876,N_8914);
or U10485 (N_10485,N_8572,N_8475);
nand U10486 (N_10486,N_8537,N_7524);
nand U10487 (N_10487,N_8525,N_8036);
or U10488 (N_10488,N_8929,N_8553);
nand U10489 (N_10489,N_8263,N_8759);
and U10490 (N_10490,N_7516,N_7513);
xnor U10491 (N_10491,N_8174,N_8945);
and U10492 (N_10492,N_7899,N_8231);
or U10493 (N_10493,N_7629,N_8077);
or U10494 (N_10494,N_8220,N_8387);
xnor U10495 (N_10495,N_8171,N_8432);
nand U10496 (N_10496,N_7878,N_8442);
or U10497 (N_10497,N_8316,N_8868);
nand U10498 (N_10498,N_8233,N_8227);
nor U10499 (N_10499,N_8211,N_8867);
xor U10500 (N_10500,N_9384,N_10286);
or U10501 (N_10501,N_9534,N_9179);
or U10502 (N_10502,N_9140,N_10400);
or U10503 (N_10503,N_9945,N_9035);
nor U10504 (N_10504,N_10133,N_9898);
and U10505 (N_10505,N_10335,N_10442);
and U10506 (N_10506,N_10237,N_10075);
nand U10507 (N_10507,N_10326,N_9561);
xor U10508 (N_10508,N_10433,N_9076);
and U10509 (N_10509,N_10385,N_9505);
and U10510 (N_10510,N_9475,N_9065);
nor U10511 (N_10511,N_10211,N_9351);
and U10512 (N_10512,N_10159,N_9258);
and U10513 (N_10513,N_10432,N_10425);
and U10514 (N_10514,N_10239,N_10370);
nand U10515 (N_10515,N_9191,N_9488);
nand U10516 (N_10516,N_9409,N_10386);
nand U10517 (N_10517,N_10248,N_9102);
or U10518 (N_10518,N_9448,N_9425);
or U10519 (N_10519,N_9984,N_9469);
nor U10520 (N_10520,N_10052,N_9611);
or U10521 (N_10521,N_9257,N_9695);
xor U10522 (N_10522,N_9563,N_9702);
and U10523 (N_10523,N_9373,N_10156);
nand U10524 (N_10524,N_10293,N_9397);
nand U10525 (N_10525,N_9062,N_9283);
xnor U10526 (N_10526,N_9017,N_9345);
nor U10527 (N_10527,N_9300,N_9232);
or U10528 (N_10528,N_10255,N_9894);
or U10529 (N_10529,N_9596,N_9150);
xor U10530 (N_10530,N_9570,N_9325);
nor U10531 (N_10531,N_9506,N_9356);
nand U10532 (N_10532,N_9878,N_9946);
and U10533 (N_10533,N_9463,N_10294);
and U10534 (N_10534,N_9668,N_10138);
and U10535 (N_10535,N_10175,N_10061);
nand U10536 (N_10536,N_9437,N_10204);
and U10537 (N_10537,N_10201,N_10187);
nand U10538 (N_10538,N_9994,N_9950);
nand U10539 (N_10539,N_9739,N_10308);
and U10540 (N_10540,N_10339,N_9252);
and U10541 (N_10541,N_9004,N_10072);
or U10542 (N_10542,N_9848,N_10328);
xor U10543 (N_10543,N_9597,N_9548);
xor U10544 (N_10544,N_9074,N_9771);
or U10545 (N_10545,N_9453,N_9577);
and U10546 (N_10546,N_10194,N_10283);
nor U10547 (N_10547,N_9880,N_9395);
and U10548 (N_10548,N_10131,N_9508);
nor U10549 (N_10549,N_10404,N_10143);
xor U10550 (N_10550,N_9464,N_9827);
xor U10551 (N_10551,N_10276,N_10078);
nand U10552 (N_10552,N_9105,N_9800);
xnor U10553 (N_10553,N_10261,N_9610);
nand U10554 (N_10554,N_9981,N_9976);
nor U10555 (N_10555,N_9213,N_9954);
and U10556 (N_10556,N_9580,N_10338);
nor U10557 (N_10557,N_9914,N_9200);
xor U10558 (N_10558,N_9088,N_10142);
xnor U10559 (N_10559,N_9036,N_9816);
xnor U10560 (N_10560,N_9817,N_9371);
nor U10561 (N_10561,N_9788,N_9911);
xnor U10562 (N_10562,N_9229,N_9533);
xnor U10563 (N_10563,N_9503,N_9614);
and U10564 (N_10564,N_10110,N_9713);
or U10565 (N_10565,N_10352,N_9221);
and U10566 (N_10566,N_9810,N_9091);
or U10567 (N_10567,N_9941,N_9559);
nand U10568 (N_10568,N_9164,N_9467);
or U10569 (N_10569,N_9640,N_9882);
xnor U10570 (N_10570,N_9832,N_9658);
xor U10571 (N_10571,N_10354,N_10090);
nor U10572 (N_10572,N_9720,N_9731);
nand U10573 (N_10573,N_9360,N_9362);
or U10574 (N_10574,N_10266,N_10483);
nand U10575 (N_10575,N_9592,N_9532);
and U10576 (N_10576,N_9418,N_9947);
or U10577 (N_10577,N_10259,N_9896);
nand U10578 (N_10578,N_9414,N_9970);
xnor U10579 (N_10579,N_9645,N_9108);
or U10580 (N_10580,N_9473,N_10379);
nor U10581 (N_10581,N_9915,N_10240);
nand U10582 (N_10582,N_10149,N_10249);
xor U10583 (N_10583,N_9600,N_10340);
xnor U10584 (N_10584,N_9313,N_9187);
xor U10585 (N_10585,N_10049,N_9174);
xnor U10586 (N_10586,N_9378,N_9446);
nand U10587 (N_10587,N_10162,N_10079);
or U10588 (N_10588,N_9697,N_10295);
xor U10589 (N_10589,N_9244,N_10083);
or U10590 (N_10590,N_9392,N_9040);
and U10591 (N_10591,N_10123,N_10289);
nor U10592 (N_10592,N_9000,N_9312);
nor U10593 (N_10593,N_10322,N_9644);
or U10594 (N_10594,N_10384,N_9005);
xor U10595 (N_10595,N_10431,N_9401);
xnor U10596 (N_10596,N_10388,N_9888);
nand U10597 (N_10597,N_9028,N_9196);
xnor U10598 (N_10598,N_10472,N_10437);
nand U10599 (N_10599,N_9622,N_9456);
or U10600 (N_10600,N_9654,N_9704);
and U10601 (N_10601,N_9780,N_10378);
or U10602 (N_10602,N_10191,N_10490);
xnor U10603 (N_10603,N_9924,N_9309);
or U10604 (N_10604,N_9080,N_10224);
xor U10605 (N_10605,N_10387,N_9083);
and U10606 (N_10606,N_9770,N_9333);
xor U10607 (N_10607,N_9209,N_9698);
and U10608 (N_10608,N_9995,N_9515);
nand U10609 (N_10609,N_9122,N_9389);
or U10610 (N_10610,N_9149,N_9372);
nand U10611 (N_10611,N_9251,N_9834);
xnor U10612 (N_10612,N_10024,N_9651);
nor U10613 (N_10613,N_9912,N_9795);
nand U10614 (N_10614,N_9485,N_9661);
or U10615 (N_10615,N_9572,N_10485);
nor U10616 (N_10616,N_10051,N_9072);
and U10617 (N_10617,N_9230,N_9940);
xor U10618 (N_10618,N_9023,N_9850);
and U10619 (N_10619,N_9175,N_10145);
nand U10620 (N_10620,N_9528,N_9433);
and U10621 (N_10621,N_10214,N_9276);
nand U10622 (N_10622,N_9847,N_10252);
and U10623 (N_10623,N_10087,N_9001);
and U10624 (N_10624,N_10268,N_10334);
xnor U10625 (N_10625,N_9732,N_10190);
and U10626 (N_10626,N_10319,N_9775);
or U10627 (N_10627,N_9566,N_10174);
nor U10628 (N_10628,N_9239,N_9518);
xnor U10629 (N_10629,N_9181,N_9823);
xnor U10630 (N_10630,N_10172,N_10324);
xor U10631 (N_10631,N_10455,N_9165);
nand U10632 (N_10632,N_10153,N_10044);
nor U10633 (N_10633,N_10084,N_9055);
or U10634 (N_10634,N_9337,N_10081);
nor U10635 (N_10635,N_10107,N_10004);
and U10636 (N_10636,N_9346,N_9598);
xor U10637 (N_10637,N_10016,N_9594);
nand U10638 (N_10638,N_10235,N_10376);
and U10639 (N_10639,N_9728,N_9906);
nor U10640 (N_10640,N_10230,N_10048);
and U10641 (N_10641,N_9185,N_9854);
nand U10642 (N_10642,N_9682,N_10341);
nor U10643 (N_10643,N_9556,N_9820);
and U10644 (N_10644,N_9609,N_10140);
nor U10645 (N_10645,N_9747,N_10192);
nor U10646 (N_10646,N_9536,N_10114);
nor U10647 (N_10647,N_9043,N_9326);
nand U10648 (N_10648,N_10436,N_9218);
xnor U10649 (N_10649,N_10426,N_9367);
nand U10650 (N_10650,N_9988,N_9826);
nor U10651 (N_10651,N_9949,N_9694);
and U10652 (N_10652,N_9303,N_10070);
and U10653 (N_10653,N_10014,N_10113);
and U10654 (N_10654,N_9342,N_9909);
nand U10655 (N_10655,N_9078,N_10029);
or U10656 (N_10656,N_9321,N_10257);
and U10657 (N_10657,N_10375,N_9650);
nand U10658 (N_10658,N_9095,N_10023);
or U10659 (N_10659,N_9126,N_9989);
nor U10660 (N_10660,N_10305,N_10085);
and U10661 (N_10661,N_9860,N_9159);
or U10662 (N_10662,N_10095,N_9869);
xor U10663 (N_10663,N_9412,N_10122);
or U10664 (N_10664,N_10499,N_9586);
xnor U10665 (N_10665,N_9049,N_10273);
xor U10666 (N_10666,N_9639,N_9240);
xnor U10667 (N_10667,N_9838,N_9932);
xor U10668 (N_10668,N_9608,N_9765);
nor U10669 (N_10669,N_9544,N_10034);
or U10670 (N_10670,N_9601,N_9830);
xor U10671 (N_10671,N_9757,N_10112);
or U10672 (N_10672,N_9223,N_9242);
nor U10673 (N_10673,N_10045,N_9047);
or U10674 (N_10674,N_9376,N_9408);
or U10675 (N_10675,N_9510,N_10226);
nor U10676 (N_10676,N_9107,N_9605);
nor U10677 (N_10677,N_10050,N_9135);
nand U10678 (N_10678,N_9013,N_9216);
xnor U10679 (N_10679,N_10451,N_9393);
nor U10680 (N_10680,N_9099,N_9273);
nor U10681 (N_10681,N_10101,N_9226);
nand U10682 (N_10682,N_9018,N_10482);
nand U10683 (N_10683,N_9824,N_9841);
nor U10684 (N_10684,N_9477,N_9910);
nand U10685 (N_10685,N_9071,N_10017);
or U10686 (N_10686,N_9134,N_9426);
nor U10687 (N_10687,N_9328,N_9936);
nor U10688 (N_10688,N_9428,N_10054);
nor U10689 (N_10689,N_10285,N_9812);
xor U10690 (N_10690,N_9655,N_10018);
or U10691 (N_10691,N_9738,N_9501);
and U10692 (N_10692,N_9039,N_9669);
xor U10693 (N_10693,N_9724,N_9297);
nand U10694 (N_10694,N_10111,N_9247);
and U10695 (N_10695,N_10146,N_9246);
and U10696 (N_10696,N_9840,N_10011);
or U10697 (N_10697,N_10414,N_10181);
or U10698 (N_10698,N_9806,N_9522);
or U10699 (N_10699,N_10222,N_10027);
nor U10700 (N_10700,N_10343,N_10418);
and U10701 (N_10701,N_9543,N_10231);
nor U10702 (N_10702,N_9993,N_9278);
nor U10703 (N_10703,N_9427,N_9461);
nand U10704 (N_10704,N_9447,N_9194);
nor U10705 (N_10705,N_9969,N_9712);
nor U10706 (N_10706,N_9865,N_10148);
xor U10707 (N_10707,N_10361,N_10165);
or U10708 (N_10708,N_9589,N_9862);
nand U10709 (N_10709,N_10046,N_9861);
nor U10710 (N_10710,N_9130,N_9098);
and U10711 (N_10711,N_9541,N_9207);
nor U10712 (N_10712,N_10321,N_9803);
xor U10713 (N_10713,N_10368,N_10434);
nand U10714 (N_10714,N_9144,N_10058);
xor U10715 (N_10715,N_9934,N_9562);
and U10716 (N_10716,N_10307,N_9270);
nand U10717 (N_10717,N_10185,N_9998);
nor U10718 (N_10718,N_10401,N_9417);
and U10719 (N_10719,N_10106,N_9253);
xnor U10720 (N_10720,N_10118,N_9727);
nor U10721 (N_10721,N_10074,N_9415);
nor U10722 (N_10722,N_10120,N_9602);
xor U10723 (N_10723,N_9919,N_9929);
nand U10724 (N_10724,N_10177,N_9769);
nand U10725 (N_10725,N_9081,N_9920);
and U10726 (N_10726,N_10329,N_9009);
or U10727 (N_10727,N_10160,N_9784);
and U10728 (N_10728,N_9466,N_9131);
nor U10729 (N_10729,N_9203,N_9762);
or U10730 (N_10730,N_10117,N_10151);
nand U10731 (N_10731,N_9740,N_9670);
xnor U10732 (N_10732,N_9129,N_9112);
nor U10733 (N_10733,N_9643,N_9406);
nand U10734 (N_10734,N_9547,N_9517);
nand U10735 (N_10735,N_9452,N_10232);
nand U10736 (N_10736,N_9141,N_10141);
nor U10737 (N_10737,N_9354,N_10447);
xnor U10738 (N_10738,N_9899,N_10032);
nand U10739 (N_10739,N_9250,N_10492);
and U10740 (N_10740,N_9304,N_9237);
xnor U10741 (N_10741,N_10128,N_10465);
or U10742 (N_10742,N_9109,N_9343);
nand U10743 (N_10743,N_9523,N_9774);
and U10744 (N_10744,N_10258,N_10277);
nand U10745 (N_10745,N_9557,N_9335);
or U10746 (N_10746,N_10331,N_9167);
or U10747 (N_10747,N_9382,N_10167);
xnor U10748 (N_10748,N_10207,N_9590);
nand U10749 (N_10749,N_9012,N_10150);
or U10750 (N_10750,N_10275,N_9494);
and U10751 (N_10751,N_9269,N_9451);
or U10752 (N_10752,N_9220,N_10461);
and U10753 (N_10753,N_9821,N_10419);
and U10754 (N_10754,N_9917,N_9705);
xor U10755 (N_10755,N_10064,N_9444);
and U10756 (N_10756,N_9858,N_10394);
nand U10757 (N_10757,N_10456,N_9918);
nand U10758 (N_10758,N_9805,N_9472);
or U10759 (N_10759,N_10154,N_9199);
or U10760 (N_10760,N_10066,N_9400);
nand U10761 (N_10761,N_9569,N_9723);
or U10762 (N_10762,N_9222,N_9678);
nand U10763 (N_10763,N_10299,N_9845);
and U10764 (N_10764,N_9429,N_9646);
xnor U10765 (N_10765,N_9520,N_9966);
nand U10766 (N_10766,N_9010,N_9143);
and U10767 (N_10767,N_9708,N_10246);
nand U10768 (N_10768,N_9020,N_10126);
xnor U10769 (N_10769,N_9125,N_9127);
nor U10770 (N_10770,N_10247,N_9015);
nor U10771 (N_10771,N_9254,N_9474);
and U10772 (N_10772,N_9366,N_9613);
and U10773 (N_10773,N_9624,N_10309);
or U10774 (N_10774,N_9267,N_9975);
xor U10775 (N_10775,N_10065,N_9524);
xor U10776 (N_10776,N_10313,N_9011);
or U10777 (N_10777,N_9772,N_10033);
and U10778 (N_10778,N_9292,N_9443);
nor U10779 (N_10779,N_10330,N_10410);
nand U10780 (N_10780,N_10096,N_9776);
or U10781 (N_10781,N_9877,N_9266);
or U10782 (N_10782,N_10020,N_10038);
nand U10783 (N_10783,N_10274,N_9907);
or U10784 (N_10784,N_10306,N_9963);
nor U10785 (N_10785,N_9671,N_9576);
or U10786 (N_10786,N_9407,N_9208);
nand U10787 (N_10787,N_9859,N_10478);
and U10788 (N_10788,N_9552,N_10301);
nor U10789 (N_10789,N_9582,N_10069);
xor U10790 (N_10790,N_9275,N_9147);
nand U10791 (N_10791,N_9318,N_9837);
nor U10792 (N_10792,N_9980,N_10026);
nor U10793 (N_10793,N_9476,N_10443);
nor U10794 (N_10794,N_10345,N_10012);
and U10795 (N_10795,N_9166,N_9420);
nand U10796 (N_10796,N_10179,N_9883);
xnor U10797 (N_10797,N_10062,N_9169);
nand U10798 (N_10798,N_9014,N_9077);
and U10799 (N_10799,N_10407,N_10287);
xnor U10800 (N_10800,N_9692,N_9120);
nand U10801 (N_10801,N_10473,N_9884);
nor U10802 (N_10802,N_9939,N_10374);
nand U10803 (N_10803,N_9926,N_9627);
and U10804 (N_10804,N_9311,N_9060);
nor U10805 (N_10805,N_10008,N_10203);
and U10806 (N_10806,N_9227,N_10316);
nor U10807 (N_10807,N_10183,N_9491);
xnor U10808 (N_10808,N_9758,N_9736);
nor U10809 (N_10809,N_10007,N_9686);
xnor U10810 (N_10810,N_9688,N_9277);
and U10811 (N_10811,N_10489,N_9288);
nor U10812 (N_10812,N_9486,N_9113);
nand U10813 (N_10813,N_10362,N_9256);
or U10814 (N_10814,N_9804,N_9274);
nor U10815 (N_10815,N_9801,N_9449);
and U10816 (N_10816,N_9468,N_9104);
xnor U10817 (N_10817,N_9497,N_9396);
xnor U10818 (N_10818,N_10399,N_9419);
nand U10819 (N_10819,N_9892,N_9152);
nor U10820 (N_10820,N_9402,N_10464);
nor U10821 (N_10821,N_9195,N_9499);
xor U10822 (N_10822,N_9157,N_9905);
and U10823 (N_10823,N_9025,N_9148);
nor U10824 (N_10824,N_9302,N_9942);
nor U10825 (N_10825,N_9903,N_10363);
or U10826 (N_10826,N_10170,N_10225);
or U10827 (N_10827,N_10219,N_9819);
nor U10828 (N_10828,N_9068,N_9733);
nand U10829 (N_10829,N_9484,N_9279);
or U10830 (N_10830,N_9158,N_9089);
xnor U10831 (N_10831,N_9928,N_9349);
nor U10832 (N_10832,N_9070,N_9146);
and U10833 (N_10833,N_10221,N_9836);
nand U10834 (N_10834,N_9359,N_10344);
or U10835 (N_10835,N_9383,N_9599);
nor U10836 (N_10836,N_9923,N_9843);
or U10837 (N_10837,N_9663,N_9675);
xnor U10838 (N_10838,N_9405,N_10039);
nor U10839 (N_10839,N_9323,N_9991);
and U10840 (N_10840,N_9990,N_10280);
and U10841 (N_10841,N_9375,N_9096);
or U10842 (N_10842,N_9549,N_9377);
or U10843 (N_10843,N_9790,N_9137);
nand U10844 (N_10844,N_9162,N_9992);
xnor U10845 (N_10845,N_10152,N_9768);
nand U10846 (N_10846,N_9635,N_9709);
and U10847 (N_10847,N_9938,N_9489);
xor U10848 (N_10848,N_9585,N_9571);
nor U10849 (N_10849,N_9701,N_10139);
nor U10850 (N_10850,N_10291,N_9595);
nor U10851 (N_10851,N_9197,N_9783);
and U10852 (N_10852,N_9887,N_9974);
nand U10853 (N_10853,N_10184,N_10272);
xor U10854 (N_10854,N_10271,N_9616);
xor U10855 (N_10855,N_9295,N_9690);
and U10856 (N_10856,N_9703,N_9173);
nand U10857 (N_10857,N_9538,N_10071);
nor U10858 (N_10858,N_10041,N_10367);
nand U10859 (N_10859,N_10342,N_9050);
xnor U10860 (N_10860,N_10168,N_9742);
and U10861 (N_10861,N_10424,N_9511);
or U10862 (N_10862,N_9202,N_9927);
nand U10863 (N_10863,N_10470,N_9344);
nor U10864 (N_10864,N_9868,N_9657);
and U10865 (N_10865,N_9734,N_9455);
nand U10866 (N_10866,N_10360,N_9054);
nor U10867 (N_10867,N_10031,N_10390);
and U10868 (N_10868,N_10365,N_9641);
nor U10869 (N_10869,N_9492,N_9410);
nand U10870 (N_10870,N_10364,N_9893);
nor U10871 (N_10871,N_10264,N_9458);
xor U10872 (N_10872,N_9038,N_10245);
and U10873 (N_10873,N_9007,N_9959);
and U10874 (N_10874,N_9459,N_10318);
xnor U10875 (N_10875,N_9829,N_9554);
or U10876 (N_10876,N_9656,N_9867);
and U10877 (N_10877,N_9027,N_9440);
nand U10878 (N_10878,N_9773,N_9086);
or U10879 (N_10879,N_9358,N_10463);
nand U10880 (N_10880,N_9073,N_9537);
or U10881 (N_10881,N_9890,N_9735);
nand U10882 (N_10882,N_9003,N_9962);
or U10883 (N_10883,N_10242,N_9314);
nor U10884 (N_10884,N_9961,N_10163);
and U10885 (N_10885,N_9057,N_9673);
nor U10886 (N_10886,N_9215,N_9807);
nand U10887 (N_10887,N_9886,N_9211);
and U10888 (N_10888,N_10218,N_9293);
nand U10889 (N_10889,N_9363,N_10005);
xnor U10890 (N_10890,N_10125,N_9574);
nor U10891 (N_10891,N_9818,N_10395);
and U10892 (N_10892,N_10025,N_10169);
nor U10893 (N_10893,N_10358,N_9483);
and U10894 (N_10894,N_9863,N_9432);
nor U10895 (N_10895,N_9618,N_9638);
xor U10896 (N_10896,N_10406,N_9411);
nand U10897 (N_10897,N_9567,N_9982);
and U10898 (N_10898,N_10488,N_9802);
nand U10899 (N_10899,N_9857,N_9977);
and U10900 (N_10900,N_9891,N_9814);
xnor U10901 (N_10901,N_9353,N_10157);
nand U10902 (N_10902,N_10332,N_10474);
nand U10903 (N_10903,N_9948,N_10098);
nand U10904 (N_10904,N_9987,N_9636);
nor U10905 (N_10905,N_9403,N_9063);
xor U10906 (N_10906,N_9413,N_10173);
xor U10907 (N_10907,N_9759,N_10459);
nand U10908 (N_10908,N_9777,N_10348);
nor U10909 (N_10909,N_9394,N_9555);
and U10910 (N_10910,N_9214,N_9956);
xor U10911 (N_10911,N_10320,N_10333);
nor U10912 (N_10912,N_10284,N_9301);
nand U10913 (N_10913,N_9438,N_9512);
nor U10914 (N_10914,N_9271,N_10176);
nor U10915 (N_10915,N_9481,N_9404);
xor U10916 (N_10916,N_9016,N_9235);
nor U10917 (N_10917,N_9665,N_10228);
nand U10918 (N_10918,N_9593,N_9116);
nor U10919 (N_10919,N_9059,N_9714);
or U10920 (N_10920,N_9796,N_9324);
and U10921 (N_10921,N_9672,N_9763);
or U10922 (N_10922,N_9317,N_10270);
nand U10923 (N_10923,N_9051,N_9336);
xnor U10924 (N_10924,N_10389,N_9037);
and U10925 (N_10925,N_9677,N_10467);
nor U10926 (N_10926,N_10234,N_10415);
nand U10927 (N_10927,N_9550,N_10357);
nor U10928 (N_10928,N_9542,N_9008);
xor U10929 (N_10929,N_9730,N_9809);
xnor U10930 (N_10930,N_9531,N_9971);
and U10931 (N_10931,N_10346,N_9287);
and U10932 (N_10932,N_10337,N_9741);
xor U10933 (N_10933,N_9516,N_10212);
and U10934 (N_10934,N_9441,N_10380);
or U10935 (N_10935,N_9154,N_9846);
nor U10936 (N_10936,N_9509,N_9588);
and U10937 (N_10937,N_10208,N_9307);
and U10938 (N_10938,N_9424,N_9368);
nor U10939 (N_10939,N_10460,N_9815);
nor U10940 (N_10940,N_10077,N_9176);
or U10941 (N_10941,N_10427,N_9519);
and U10942 (N_10942,N_9500,N_9075);
xnor U10943 (N_10943,N_9831,N_9445);
nand U10944 (N_10944,N_9649,N_9299);
or U10945 (N_10945,N_9546,N_9183);
nand U10946 (N_10946,N_9067,N_9607);
nand U10947 (N_10947,N_10392,N_9679);
nand U10948 (N_10948,N_10093,N_9034);
nand U10949 (N_10949,N_9957,N_9902);
and U10950 (N_10950,N_9625,N_10178);
or U10951 (N_10951,N_9856,N_9729);
xnor U10952 (N_10952,N_10458,N_9755);
nand U10953 (N_10953,N_9718,N_10495);
or U10954 (N_10954,N_9338,N_9699);
nor U10955 (N_10955,N_9922,N_9983);
nand U10956 (N_10956,N_9289,N_9330);
xnor U10957 (N_10957,N_9390,N_10028);
or U10958 (N_10958,N_9296,N_10042);
and U10959 (N_10959,N_10466,N_10055);
or U10960 (N_10960,N_9716,N_9745);
nand U10961 (N_10961,N_9558,N_9069);
nor U10962 (N_10962,N_9233,N_9872);
and U10963 (N_10963,N_9357,N_9243);
nor U10964 (N_10964,N_9659,N_10241);
or U10965 (N_10965,N_10398,N_9327);
and U10966 (N_10966,N_9182,N_9308);
xnor U10967 (N_10967,N_10315,N_9931);
nor U10968 (N_10968,N_10198,N_10353);
and U10969 (N_10969,N_9913,N_9155);
nand U10970 (N_10970,N_10091,N_10010);
or U10971 (N_10971,N_10130,N_9794);
and U10972 (N_10972,N_10209,N_9999);
and U10973 (N_10973,N_9587,N_10484);
nor U10974 (N_10974,N_9092,N_9706);
or U10975 (N_10975,N_9921,N_9265);
and U10976 (N_10976,N_10336,N_9084);
nand U10977 (N_10977,N_9683,N_9791);
nand U10978 (N_10978,N_9666,N_9190);
nor U10979 (N_10979,N_9128,N_9689);
nor U10980 (N_10980,N_9482,N_9041);
and U10981 (N_10981,N_10200,N_10199);
xnor U10982 (N_10982,N_9870,N_9284);
or U10983 (N_10983,N_9851,N_9114);
and U10984 (N_10984,N_9132,N_9753);
nand U10985 (N_10985,N_10030,N_9535);
nor U10986 (N_10986,N_9767,N_9044);
xor U10987 (N_10987,N_9852,N_9591);
nand U10988 (N_10988,N_9103,N_9935);
and U10989 (N_10989,N_9052,N_9897);
xor U10990 (N_10990,N_9664,N_9217);
or U10991 (N_10991,N_9198,N_9434);
nor U10992 (N_10992,N_9876,N_9163);
xnor U10993 (N_10993,N_9853,N_9234);
or U10994 (N_10994,N_10469,N_9766);
xor U10995 (N_10995,N_9828,N_9178);
xor U10996 (N_10996,N_9145,N_9462);
and U10997 (N_10997,N_9093,N_9225);
xor U10998 (N_10998,N_10256,N_9136);
nor U10999 (N_10999,N_9539,N_10409);
nand U11000 (N_11000,N_9340,N_9514);
and U11001 (N_11001,N_10440,N_9204);
xor U11002 (N_11002,N_9507,N_10129);
nand U11003 (N_11003,N_9513,N_10099);
or U11004 (N_11004,N_9953,N_9952);
nor U11005 (N_11005,N_9889,N_10417);
nor U11006 (N_11006,N_9560,N_10086);
and U11007 (N_11007,N_10450,N_10223);
xor U11008 (N_11008,N_9281,N_10119);
nor U11009 (N_11009,N_9056,N_9298);
nand U11010 (N_11010,N_10251,N_9118);
nand U11011 (N_11011,N_10438,N_9231);
nand U11012 (N_11012,N_9684,N_9498);
or U11013 (N_11013,N_9652,N_10480);
or U11014 (N_11014,N_9026,N_9272);
or U11015 (N_11015,N_9031,N_9238);
and U11016 (N_11016,N_9808,N_10003);
nand U11017 (N_11017,N_9637,N_9294);
nor U11018 (N_11018,N_9626,N_9792);
nand U11019 (N_11019,N_10366,N_9110);
nor U11020 (N_11020,N_10359,N_9348);
xnor U11021 (N_11021,N_9264,N_10135);
xnor U11022 (N_11022,N_10314,N_9925);
and U11023 (N_11023,N_10381,N_10449);
and U11024 (N_11024,N_10193,N_10002);
or U11025 (N_11025,N_9454,N_9710);
xor U11026 (N_11026,N_9750,N_10080);
nand U11027 (N_11027,N_9642,N_9450);
xor U11028 (N_11028,N_10227,N_10448);
nor U11029 (N_11029,N_9979,N_9320);
or U11030 (N_11030,N_9748,N_10303);
nor U11031 (N_11031,N_10195,N_9119);
or U11032 (N_11032,N_10265,N_10116);
nor U11033 (N_11033,N_9781,N_10396);
or U11034 (N_11034,N_10403,N_10282);
nand U11035 (N_11035,N_9908,N_9530);
and U11036 (N_11036,N_9789,N_10053);
or U11037 (N_11037,N_9361,N_9575);
and U11038 (N_11038,N_9100,N_10136);
nor U11039 (N_11039,N_9881,N_9285);
and U11040 (N_11040,N_9142,N_9874);
nor U11041 (N_11041,N_10134,N_9681);
and U11042 (N_11042,N_9864,N_9612);
and U11043 (N_11043,N_9811,N_9839);
nor U11044 (N_11044,N_9540,N_10304);
nand U11045 (N_11045,N_9667,N_9717);
xnor U11046 (N_11046,N_10108,N_9579);
xnor U11047 (N_11047,N_9442,N_10009);
nor U11048 (N_11048,N_9944,N_9315);
nand U11049 (N_11049,N_10089,N_9900);
nor U11050 (N_11050,N_10263,N_9743);
xnor U11051 (N_11051,N_10144,N_9374);
nor U11052 (N_11052,N_9955,N_10260);
xnor U11053 (N_11053,N_9904,N_10323);
nand U11054 (N_11054,N_9787,N_9123);
xor U11055 (N_11055,N_9604,N_10453);
xor U11056 (N_11056,N_10121,N_10220);
or U11057 (N_11057,N_9722,N_9082);
nand U11058 (N_11058,N_10103,N_9436);
nand U11059 (N_11059,N_10059,N_9568);
nor U11060 (N_11060,N_9495,N_10372);
nor U11061 (N_11061,N_9496,N_9385);
and U11062 (N_11062,N_9282,N_9879);
nand U11063 (N_11063,N_9721,N_9306);
xnor U11064 (N_11064,N_10067,N_9212);
nor U11065 (N_11065,N_10006,N_9061);
nand U11066 (N_11066,N_9006,N_9521);
or U11067 (N_11067,N_10278,N_10104);
and U11068 (N_11068,N_9583,N_10371);
nand U11069 (N_11069,N_9172,N_10082);
nand U11070 (N_11070,N_9551,N_10296);
or U11071 (N_11071,N_9628,N_9490);
or U11072 (N_11072,N_10267,N_10088);
nor U11073 (N_11073,N_9855,N_10056);
xor U11074 (N_11074,N_10391,N_9779);
or U11075 (N_11075,N_10105,N_9364);
nor U11076 (N_11076,N_9117,N_9291);
or U11077 (N_11077,N_9460,N_9268);
and U11078 (N_11078,N_9606,N_9019);
xor U11079 (N_11079,N_9248,N_9584);
and U11080 (N_11080,N_9631,N_9310);
xnor U11081 (N_11081,N_9021,N_9901);
and U11082 (N_11082,N_10127,N_9316);
nand U11083 (N_11083,N_9978,N_9849);
nor U11084 (N_11084,N_9380,N_10182);
or U11085 (N_11085,N_9825,N_10327);
nor U11086 (N_11086,N_9687,N_10215);
or U11087 (N_11087,N_9798,N_10202);
xor U11088 (N_11088,N_10137,N_10197);
nand U11089 (N_11089,N_9219,N_9756);
xnor U11090 (N_11090,N_10040,N_10420);
or U11091 (N_11091,N_10413,N_9066);
xnor U11092 (N_11092,N_9097,N_9391);
or U11093 (N_11093,N_9032,N_9184);
nand U11094 (N_11094,N_10412,N_9228);
nand U11095 (N_11095,N_10422,N_9630);
and U11096 (N_11096,N_9746,N_9024);
and U11097 (N_11097,N_10408,N_10405);
nand U11098 (N_11098,N_9553,N_9261);
and U11099 (N_11099,N_9725,N_9972);
xnor U11100 (N_11100,N_9171,N_9002);
nand U11101 (N_11101,N_9087,N_9170);
xor U11102 (N_11102,N_9958,N_9526);
or U11103 (N_11103,N_9564,N_9799);
xnor U11104 (N_11104,N_9205,N_9262);
xor U11105 (N_11105,N_9465,N_9470);
nor U11106 (N_11106,N_9430,N_9662);
nor U11107 (N_11107,N_9933,N_9951);
or U11108 (N_11108,N_9964,N_9754);
nand U11109 (N_11109,N_10302,N_9193);
xnor U11110 (N_11110,N_9930,N_9201);
nor U11111 (N_11111,N_9480,N_9711);
nor U11112 (N_11112,N_10402,N_9633);
xor U11113 (N_11113,N_10430,N_9674);
xnor U11114 (N_11114,N_10188,N_10423);
xnor U11115 (N_11115,N_9332,N_10281);
or U11116 (N_11116,N_9439,N_10216);
and U11117 (N_11117,N_9022,N_10317);
and U11118 (N_11118,N_10076,N_9138);
or U11119 (N_11119,N_9350,N_10421);
or U11120 (N_11120,N_10429,N_9844);
nand U11121 (N_11121,N_9707,N_10253);
nand U11122 (N_11122,N_9545,N_10043);
and U11123 (N_11123,N_9079,N_9085);
or U11124 (N_11124,N_9186,N_10236);
nand U11125 (N_11125,N_9334,N_9786);
nor U11126 (N_11126,N_9967,N_10454);
or U11127 (N_11127,N_9280,N_9094);
xor U11128 (N_11128,N_10416,N_9115);
nor U11129 (N_11129,N_10397,N_10147);
and U11130 (N_11130,N_9968,N_9236);
or U11131 (N_11131,N_10494,N_10155);
xor U11132 (N_11132,N_10462,N_10097);
xor U11133 (N_11133,N_9479,N_9764);
nor U11134 (N_11134,N_9737,N_9504);
or U11135 (N_11135,N_10196,N_10164);
xnor U11136 (N_11136,N_9875,N_9156);
or U11137 (N_11137,N_10269,N_9685);
xnor U11138 (N_11138,N_9719,N_9153);
xor U11139 (N_11139,N_10060,N_10475);
nand U11140 (N_11140,N_10444,N_10471);
nor U11141 (N_11141,N_10325,N_9124);
and U11142 (N_11142,N_10254,N_9617);
xnor U11143 (N_11143,N_9744,N_9322);
nor U11144 (N_11144,N_9478,N_10486);
nand U11145 (N_11145,N_9048,N_9033);
xnor U11146 (N_11146,N_9160,N_9457);
xor U11147 (N_11147,N_9399,N_9660);
or U11148 (N_11148,N_10171,N_9778);
and U11149 (N_11149,N_9895,N_10382);
and U11150 (N_11150,N_9369,N_10102);
nand U11151 (N_11151,N_9139,N_9691);
xnor U11152 (N_11152,N_10001,N_9493);
and U11153 (N_11153,N_9259,N_9168);
nor U11154 (N_11154,N_9263,N_10349);
xor U11155 (N_11155,N_9177,N_9965);
and U11156 (N_11156,N_9916,N_9873);
nor U11157 (N_11157,N_9696,N_10393);
or U11158 (N_11158,N_9615,N_9603);
or U11159 (N_11159,N_9680,N_9997);
or U11160 (N_11160,N_9676,N_9749);
and U11161 (N_11161,N_10279,N_9943);
and U11162 (N_11162,N_9339,N_9106);
nor U11163 (N_11163,N_10292,N_10310);
xnor U11164 (N_11164,N_9937,N_9133);
or U11165 (N_11165,N_10022,N_9319);
xnor U11166 (N_11166,N_9621,N_9620);
nand U11167 (N_11167,N_10373,N_10238);
nor U11168 (N_11168,N_10037,N_10369);
and U11169 (N_11169,N_10481,N_10013);
and U11170 (N_11170,N_10262,N_9046);
and U11171 (N_11171,N_10019,N_9249);
and U11172 (N_11172,N_10498,N_9693);
nor U11173 (N_11173,N_10439,N_10468);
nor U11174 (N_11174,N_9782,N_10213);
and U11175 (N_11175,N_9151,N_10180);
xor U11176 (N_11176,N_10356,N_9797);
and U11177 (N_11177,N_10035,N_9305);
and U11178 (N_11178,N_9387,N_9341);
xnor U11179 (N_11179,N_10300,N_9111);
or U11180 (N_11180,N_9029,N_10476);
nand U11181 (N_11181,N_9822,N_9813);
xor U11182 (N_11182,N_10109,N_10411);
nor U11183 (N_11183,N_9206,N_10166);
xnor U11184 (N_11184,N_9578,N_10186);
and U11185 (N_11185,N_9527,N_9210);
or U11186 (N_11186,N_9290,N_10092);
nand U11187 (N_11187,N_9726,N_10205);
nor U11188 (N_11188,N_9189,N_9996);
nor U11189 (N_11189,N_9653,N_10250);
xnor U11190 (N_11190,N_10298,N_10161);
and U11191 (N_11191,N_9286,N_9416);
nand U11192 (N_11192,N_9623,N_9502);
xor U11193 (N_11193,N_9529,N_10446);
nor U11194 (N_11194,N_9370,N_10497);
and U11195 (N_11195,N_10347,N_10217);
nor U11196 (N_11196,N_10073,N_9647);
nor U11197 (N_11197,N_9121,N_9785);
or U11198 (N_11198,N_9715,N_9634);
or U11199 (N_11199,N_9700,N_10288);
nand U11200 (N_11200,N_9422,N_10063);
or U11201 (N_11201,N_10452,N_9423);
nand U11202 (N_11202,N_10015,N_9180);
nor U11203 (N_11203,N_9101,N_10115);
and U11204 (N_11204,N_9471,N_10000);
nor U11205 (N_11205,N_9381,N_10021);
nor U11206 (N_11206,N_10036,N_9632);
xnor U11207 (N_11207,N_10229,N_9986);
nand U11208 (N_11208,N_10158,N_9752);
or U11209 (N_11209,N_10311,N_9365);
and U11210 (N_11210,N_9090,N_10441);
nor U11211 (N_11211,N_9581,N_10297);
xor U11212 (N_11212,N_9355,N_9161);
nor U11213 (N_11213,N_9398,N_9042);
nand U11214 (N_11214,N_9487,N_9347);
xnor U11215 (N_11215,N_10244,N_10350);
and U11216 (N_11216,N_10210,N_10057);
nor U11217 (N_11217,N_10491,N_9629);
nand U11218 (N_11218,N_9379,N_10094);
xor U11219 (N_11219,N_10068,N_9565);
nor U11220 (N_11220,N_9619,N_9058);
nor U11221 (N_11221,N_10445,N_9260);
and U11222 (N_11222,N_10312,N_10100);
nand U11223 (N_11223,N_9573,N_10047);
nand U11224 (N_11224,N_10487,N_9331);
xor U11225 (N_11225,N_9431,N_9866);
nor U11226 (N_11226,N_9885,N_9835);
nand U11227 (N_11227,N_10124,N_9421);
nand U11228 (N_11228,N_9760,N_9030);
and U11229 (N_11229,N_9842,N_10189);
nor U11230 (N_11230,N_9224,N_10132);
nand U11231 (N_11231,N_10383,N_9188);
and U11232 (N_11232,N_10435,N_10355);
nand U11233 (N_11233,N_9329,N_9761);
and U11234 (N_11234,N_9793,N_9388);
nand U11235 (N_11235,N_9833,N_9648);
nand U11236 (N_11236,N_10290,N_10233);
or U11237 (N_11237,N_10479,N_9245);
nor U11238 (N_11238,N_10428,N_9960);
or U11239 (N_11239,N_9435,N_9255);
nand U11240 (N_11240,N_9525,N_9386);
nand U11241 (N_11241,N_9064,N_9973);
nand U11242 (N_11242,N_10496,N_9985);
and U11243 (N_11243,N_9241,N_9045);
and U11244 (N_11244,N_10457,N_10477);
nand U11245 (N_11245,N_9053,N_10493);
or U11246 (N_11246,N_10351,N_10243);
nor U11247 (N_11247,N_9352,N_9751);
or U11248 (N_11248,N_10377,N_9192);
and U11249 (N_11249,N_9871,N_10206);
nand U11250 (N_11250,N_9659,N_9403);
nor U11251 (N_11251,N_9962,N_10096);
xor U11252 (N_11252,N_9888,N_9943);
and U11253 (N_11253,N_9435,N_10061);
or U11254 (N_11254,N_9749,N_9359);
or U11255 (N_11255,N_10316,N_9559);
xnor U11256 (N_11256,N_9730,N_9817);
or U11257 (N_11257,N_10035,N_10122);
and U11258 (N_11258,N_10483,N_9856);
or U11259 (N_11259,N_10397,N_9837);
nor U11260 (N_11260,N_9101,N_9416);
nor U11261 (N_11261,N_9873,N_10129);
xor U11262 (N_11262,N_10206,N_10347);
nand U11263 (N_11263,N_9393,N_10476);
nand U11264 (N_11264,N_9140,N_10030);
xnor U11265 (N_11265,N_10311,N_9295);
or U11266 (N_11266,N_9251,N_9770);
or U11267 (N_11267,N_10450,N_10113);
xor U11268 (N_11268,N_9107,N_9600);
nor U11269 (N_11269,N_10238,N_9703);
xor U11270 (N_11270,N_10145,N_9033);
and U11271 (N_11271,N_10034,N_10308);
and U11272 (N_11272,N_9377,N_9764);
xor U11273 (N_11273,N_9589,N_10221);
and U11274 (N_11274,N_10173,N_10255);
and U11275 (N_11275,N_10347,N_10218);
xor U11276 (N_11276,N_9308,N_10141);
and U11277 (N_11277,N_9661,N_9066);
and U11278 (N_11278,N_9295,N_10275);
or U11279 (N_11279,N_9915,N_10297);
nand U11280 (N_11280,N_9393,N_9779);
xor U11281 (N_11281,N_10168,N_10055);
xnor U11282 (N_11282,N_9643,N_10260);
nand U11283 (N_11283,N_9011,N_9007);
or U11284 (N_11284,N_10297,N_10112);
or U11285 (N_11285,N_9391,N_9927);
and U11286 (N_11286,N_10459,N_9581);
or U11287 (N_11287,N_9558,N_9267);
nand U11288 (N_11288,N_9929,N_9490);
nand U11289 (N_11289,N_10036,N_9485);
xnor U11290 (N_11290,N_9918,N_9075);
and U11291 (N_11291,N_9401,N_10381);
nor U11292 (N_11292,N_9758,N_10467);
xnor U11293 (N_11293,N_9592,N_9046);
or U11294 (N_11294,N_9752,N_9834);
xor U11295 (N_11295,N_9855,N_9498);
and U11296 (N_11296,N_9078,N_9054);
and U11297 (N_11297,N_9289,N_10113);
nand U11298 (N_11298,N_10339,N_10135);
or U11299 (N_11299,N_9472,N_9822);
xnor U11300 (N_11300,N_9693,N_9965);
xnor U11301 (N_11301,N_10173,N_10428);
nor U11302 (N_11302,N_9370,N_9535);
xnor U11303 (N_11303,N_9538,N_9094);
and U11304 (N_11304,N_9847,N_9495);
nand U11305 (N_11305,N_9974,N_10099);
and U11306 (N_11306,N_10081,N_9552);
xor U11307 (N_11307,N_9479,N_10063);
nor U11308 (N_11308,N_9382,N_10091);
xor U11309 (N_11309,N_9040,N_9814);
and U11310 (N_11310,N_9143,N_10047);
nor U11311 (N_11311,N_9742,N_10262);
or U11312 (N_11312,N_10329,N_9621);
or U11313 (N_11313,N_9725,N_9163);
xnor U11314 (N_11314,N_9113,N_10181);
xor U11315 (N_11315,N_10137,N_9623);
nor U11316 (N_11316,N_10450,N_9351);
and U11317 (N_11317,N_10045,N_10067);
nor U11318 (N_11318,N_10395,N_10065);
nor U11319 (N_11319,N_9991,N_10261);
nor U11320 (N_11320,N_10375,N_10024);
and U11321 (N_11321,N_9330,N_9980);
nor U11322 (N_11322,N_9601,N_9320);
xor U11323 (N_11323,N_10135,N_9271);
nor U11324 (N_11324,N_9565,N_9164);
and U11325 (N_11325,N_9502,N_10281);
or U11326 (N_11326,N_9096,N_10423);
and U11327 (N_11327,N_9213,N_10107);
and U11328 (N_11328,N_10043,N_10282);
nand U11329 (N_11329,N_10404,N_9302);
xnor U11330 (N_11330,N_9542,N_9873);
nand U11331 (N_11331,N_10215,N_9544);
and U11332 (N_11332,N_9207,N_9407);
or U11333 (N_11333,N_9645,N_9460);
nand U11334 (N_11334,N_9777,N_10177);
nor U11335 (N_11335,N_9811,N_10360);
or U11336 (N_11336,N_9016,N_9316);
or U11337 (N_11337,N_9695,N_9622);
or U11338 (N_11338,N_10453,N_9460);
nor U11339 (N_11339,N_9189,N_9333);
or U11340 (N_11340,N_10356,N_9156);
xor U11341 (N_11341,N_9310,N_10028);
nor U11342 (N_11342,N_10201,N_9185);
or U11343 (N_11343,N_9148,N_9892);
and U11344 (N_11344,N_9973,N_10381);
nand U11345 (N_11345,N_9319,N_10328);
nand U11346 (N_11346,N_10170,N_9327);
or U11347 (N_11347,N_9335,N_9787);
nand U11348 (N_11348,N_9645,N_9271);
and U11349 (N_11349,N_9361,N_10077);
and U11350 (N_11350,N_10315,N_9502);
and U11351 (N_11351,N_10476,N_9780);
xor U11352 (N_11352,N_10005,N_9659);
and U11353 (N_11353,N_9516,N_9358);
nor U11354 (N_11354,N_9119,N_9923);
xnor U11355 (N_11355,N_9883,N_9343);
and U11356 (N_11356,N_10457,N_9822);
xnor U11357 (N_11357,N_10014,N_9759);
nor U11358 (N_11358,N_9375,N_9613);
and U11359 (N_11359,N_9388,N_9012);
xnor U11360 (N_11360,N_9402,N_10158);
nand U11361 (N_11361,N_9617,N_9080);
xnor U11362 (N_11362,N_9513,N_9145);
nand U11363 (N_11363,N_10494,N_9705);
or U11364 (N_11364,N_10408,N_10044);
nand U11365 (N_11365,N_10108,N_10348);
nand U11366 (N_11366,N_9625,N_10048);
nand U11367 (N_11367,N_10145,N_9659);
xor U11368 (N_11368,N_10265,N_10492);
xnor U11369 (N_11369,N_9716,N_9248);
or U11370 (N_11370,N_9779,N_9050);
and U11371 (N_11371,N_10268,N_10133);
nor U11372 (N_11372,N_9734,N_10204);
and U11373 (N_11373,N_9448,N_9836);
xnor U11374 (N_11374,N_10276,N_10063);
nor U11375 (N_11375,N_9882,N_10457);
nand U11376 (N_11376,N_10063,N_9248);
and U11377 (N_11377,N_9203,N_9838);
nor U11378 (N_11378,N_10170,N_9828);
and U11379 (N_11379,N_10207,N_9310);
xor U11380 (N_11380,N_10289,N_9112);
nand U11381 (N_11381,N_10238,N_10094);
nand U11382 (N_11382,N_9663,N_10368);
nand U11383 (N_11383,N_9723,N_9444);
nand U11384 (N_11384,N_9660,N_10176);
or U11385 (N_11385,N_10013,N_9119);
nand U11386 (N_11386,N_10467,N_9014);
nand U11387 (N_11387,N_9002,N_10446);
or U11388 (N_11388,N_9012,N_9078);
nor U11389 (N_11389,N_9569,N_9511);
xnor U11390 (N_11390,N_10044,N_9661);
nand U11391 (N_11391,N_9326,N_9154);
or U11392 (N_11392,N_9532,N_9788);
or U11393 (N_11393,N_9454,N_9786);
or U11394 (N_11394,N_9472,N_9160);
or U11395 (N_11395,N_9659,N_10348);
and U11396 (N_11396,N_10468,N_10336);
nor U11397 (N_11397,N_9347,N_10413);
nor U11398 (N_11398,N_9477,N_10310);
and U11399 (N_11399,N_10133,N_9909);
or U11400 (N_11400,N_9719,N_9898);
and U11401 (N_11401,N_9346,N_10225);
and U11402 (N_11402,N_9744,N_9894);
or U11403 (N_11403,N_10046,N_10390);
and U11404 (N_11404,N_10119,N_9324);
and U11405 (N_11405,N_9455,N_9806);
nor U11406 (N_11406,N_9799,N_10311);
and U11407 (N_11407,N_10195,N_9560);
nand U11408 (N_11408,N_10387,N_9635);
and U11409 (N_11409,N_9649,N_10147);
or U11410 (N_11410,N_9711,N_10386);
or U11411 (N_11411,N_9713,N_9424);
nand U11412 (N_11412,N_9181,N_9247);
or U11413 (N_11413,N_10266,N_9708);
nand U11414 (N_11414,N_9514,N_10467);
or U11415 (N_11415,N_9592,N_10086);
nand U11416 (N_11416,N_9469,N_10194);
and U11417 (N_11417,N_10474,N_9535);
nand U11418 (N_11418,N_9644,N_9526);
and U11419 (N_11419,N_10186,N_10097);
xor U11420 (N_11420,N_9448,N_9778);
nand U11421 (N_11421,N_10038,N_10478);
nor U11422 (N_11422,N_9160,N_9697);
nor U11423 (N_11423,N_9344,N_9618);
nand U11424 (N_11424,N_10011,N_10450);
or U11425 (N_11425,N_9068,N_9723);
and U11426 (N_11426,N_9118,N_10198);
or U11427 (N_11427,N_9658,N_9581);
and U11428 (N_11428,N_9724,N_9451);
or U11429 (N_11429,N_9897,N_9460);
or U11430 (N_11430,N_9505,N_10169);
and U11431 (N_11431,N_9608,N_10352);
xnor U11432 (N_11432,N_10029,N_9768);
nand U11433 (N_11433,N_9610,N_9794);
nor U11434 (N_11434,N_9091,N_9723);
and U11435 (N_11435,N_9867,N_9174);
nor U11436 (N_11436,N_9168,N_9210);
nand U11437 (N_11437,N_9152,N_9725);
nor U11438 (N_11438,N_9221,N_9209);
or U11439 (N_11439,N_10464,N_9006);
or U11440 (N_11440,N_9172,N_9603);
xor U11441 (N_11441,N_9719,N_9769);
nor U11442 (N_11442,N_9897,N_10471);
nand U11443 (N_11443,N_9515,N_10093);
nand U11444 (N_11444,N_9109,N_10106);
and U11445 (N_11445,N_9236,N_10334);
nand U11446 (N_11446,N_9998,N_9603);
nor U11447 (N_11447,N_10075,N_10163);
nor U11448 (N_11448,N_10328,N_9767);
and U11449 (N_11449,N_9752,N_9335);
or U11450 (N_11450,N_9367,N_9718);
nand U11451 (N_11451,N_10289,N_9288);
xor U11452 (N_11452,N_9487,N_10371);
nand U11453 (N_11453,N_9186,N_9083);
or U11454 (N_11454,N_9830,N_9017);
nand U11455 (N_11455,N_9856,N_9438);
or U11456 (N_11456,N_9864,N_9823);
and U11457 (N_11457,N_10459,N_10315);
or U11458 (N_11458,N_10123,N_9368);
nand U11459 (N_11459,N_10287,N_10213);
xnor U11460 (N_11460,N_9636,N_9444);
nand U11461 (N_11461,N_9973,N_9347);
nor U11462 (N_11462,N_10280,N_9503);
or U11463 (N_11463,N_10188,N_9267);
xor U11464 (N_11464,N_9774,N_9649);
xnor U11465 (N_11465,N_9975,N_9628);
nand U11466 (N_11466,N_10435,N_10344);
xor U11467 (N_11467,N_9035,N_9905);
nand U11468 (N_11468,N_9490,N_10449);
nand U11469 (N_11469,N_10411,N_9211);
nor U11470 (N_11470,N_10465,N_10010);
nor U11471 (N_11471,N_9673,N_9670);
nor U11472 (N_11472,N_9386,N_9337);
xnor U11473 (N_11473,N_10304,N_9083);
or U11474 (N_11474,N_10209,N_9360);
xor U11475 (N_11475,N_10390,N_9842);
xor U11476 (N_11476,N_9214,N_9626);
or U11477 (N_11477,N_9755,N_9248);
and U11478 (N_11478,N_9531,N_9299);
nor U11479 (N_11479,N_10237,N_9297);
or U11480 (N_11480,N_9683,N_9373);
nand U11481 (N_11481,N_9497,N_10387);
nor U11482 (N_11482,N_10037,N_9049);
or U11483 (N_11483,N_9102,N_9205);
nand U11484 (N_11484,N_10443,N_9756);
and U11485 (N_11485,N_9106,N_9924);
nand U11486 (N_11486,N_9151,N_9414);
and U11487 (N_11487,N_9971,N_9498);
nor U11488 (N_11488,N_9147,N_10301);
or U11489 (N_11489,N_9599,N_10497);
xnor U11490 (N_11490,N_9387,N_9690);
and U11491 (N_11491,N_9461,N_9294);
or U11492 (N_11492,N_9670,N_10129);
xor U11493 (N_11493,N_9702,N_9006);
or U11494 (N_11494,N_9716,N_9942);
and U11495 (N_11495,N_9417,N_9304);
or U11496 (N_11496,N_9342,N_9285);
and U11497 (N_11497,N_10484,N_9626);
nor U11498 (N_11498,N_9845,N_9673);
or U11499 (N_11499,N_10448,N_9908);
nor U11500 (N_11500,N_9390,N_10138);
nor U11501 (N_11501,N_10336,N_10170);
or U11502 (N_11502,N_9781,N_9965);
nand U11503 (N_11503,N_9892,N_10178);
xnor U11504 (N_11504,N_10081,N_10423);
xnor U11505 (N_11505,N_9665,N_9192);
nor U11506 (N_11506,N_10477,N_9514);
nand U11507 (N_11507,N_9844,N_9628);
xnor U11508 (N_11508,N_9243,N_9822);
nand U11509 (N_11509,N_9856,N_9370);
xnor U11510 (N_11510,N_10259,N_10399);
nand U11511 (N_11511,N_9803,N_10115);
xnor U11512 (N_11512,N_10453,N_9660);
xnor U11513 (N_11513,N_10122,N_9301);
xor U11514 (N_11514,N_9320,N_9452);
nor U11515 (N_11515,N_9385,N_9123);
and U11516 (N_11516,N_9145,N_9463);
nor U11517 (N_11517,N_9314,N_10195);
nor U11518 (N_11518,N_10269,N_9449);
nor U11519 (N_11519,N_10019,N_10499);
or U11520 (N_11520,N_10136,N_10055);
nand U11521 (N_11521,N_9135,N_9312);
and U11522 (N_11522,N_10075,N_9602);
or U11523 (N_11523,N_9067,N_10314);
xor U11524 (N_11524,N_10386,N_9177);
nand U11525 (N_11525,N_9817,N_9582);
nand U11526 (N_11526,N_9083,N_10083);
xnor U11527 (N_11527,N_9836,N_9368);
nand U11528 (N_11528,N_9455,N_9837);
or U11529 (N_11529,N_9348,N_9808);
or U11530 (N_11530,N_10165,N_9118);
nor U11531 (N_11531,N_9810,N_9813);
and U11532 (N_11532,N_9062,N_10053);
and U11533 (N_11533,N_10286,N_10400);
and U11534 (N_11534,N_9170,N_10440);
nand U11535 (N_11535,N_10266,N_9353);
nand U11536 (N_11536,N_9906,N_10341);
xnor U11537 (N_11537,N_10323,N_10443);
nor U11538 (N_11538,N_9721,N_9207);
nand U11539 (N_11539,N_9919,N_9581);
nand U11540 (N_11540,N_10249,N_9528);
nor U11541 (N_11541,N_9414,N_9977);
and U11542 (N_11542,N_10331,N_10091);
or U11543 (N_11543,N_9843,N_9699);
nor U11544 (N_11544,N_9061,N_9499);
nor U11545 (N_11545,N_10442,N_9752);
and U11546 (N_11546,N_10354,N_9153);
or U11547 (N_11547,N_9378,N_9319);
nor U11548 (N_11548,N_9632,N_9781);
or U11549 (N_11549,N_9199,N_10457);
nand U11550 (N_11550,N_9727,N_9927);
nand U11551 (N_11551,N_9035,N_9431);
nor U11552 (N_11552,N_10479,N_10196);
and U11553 (N_11553,N_9642,N_9204);
or U11554 (N_11554,N_9317,N_9414);
nor U11555 (N_11555,N_10142,N_10323);
xor U11556 (N_11556,N_10090,N_9503);
xnor U11557 (N_11557,N_10379,N_9030);
nand U11558 (N_11558,N_9478,N_9885);
nand U11559 (N_11559,N_10457,N_9109);
nand U11560 (N_11560,N_10155,N_10096);
nand U11561 (N_11561,N_9944,N_9038);
nor U11562 (N_11562,N_9761,N_9158);
nor U11563 (N_11563,N_9866,N_10437);
nand U11564 (N_11564,N_9152,N_9418);
nand U11565 (N_11565,N_10268,N_9111);
and U11566 (N_11566,N_9922,N_9389);
xor U11567 (N_11567,N_9716,N_10450);
or U11568 (N_11568,N_9395,N_9334);
nor U11569 (N_11569,N_9237,N_9103);
nand U11570 (N_11570,N_9603,N_10420);
nor U11571 (N_11571,N_10152,N_9178);
nand U11572 (N_11572,N_9553,N_10069);
nor U11573 (N_11573,N_9596,N_10346);
nor U11574 (N_11574,N_10014,N_9232);
and U11575 (N_11575,N_9898,N_10336);
nand U11576 (N_11576,N_9915,N_10411);
xnor U11577 (N_11577,N_10291,N_10334);
or U11578 (N_11578,N_9922,N_10322);
nand U11579 (N_11579,N_10286,N_9239);
nand U11580 (N_11580,N_9593,N_9882);
nand U11581 (N_11581,N_10482,N_9762);
nand U11582 (N_11582,N_9122,N_10134);
nor U11583 (N_11583,N_10472,N_9165);
xnor U11584 (N_11584,N_9874,N_9113);
nor U11585 (N_11585,N_10350,N_10053);
or U11586 (N_11586,N_10069,N_9942);
xor U11587 (N_11587,N_9591,N_9981);
nand U11588 (N_11588,N_9133,N_9895);
nand U11589 (N_11589,N_9682,N_10445);
xor U11590 (N_11590,N_10291,N_10337);
or U11591 (N_11591,N_9795,N_9826);
nor U11592 (N_11592,N_10446,N_9236);
nor U11593 (N_11593,N_9093,N_10264);
xor U11594 (N_11594,N_9576,N_10019);
nor U11595 (N_11595,N_10201,N_9807);
or U11596 (N_11596,N_9559,N_9434);
or U11597 (N_11597,N_9803,N_9155);
nand U11598 (N_11598,N_9201,N_9834);
nor U11599 (N_11599,N_9180,N_9475);
xnor U11600 (N_11600,N_9082,N_10071);
nor U11601 (N_11601,N_9131,N_10187);
nand U11602 (N_11602,N_10182,N_10076);
or U11603 (N_11603,N_9996,N_9989);
or U11604 (N_11604,N_9324,N_9905);
nor U11605 (N_11605,N_10251,N_10472);
nor U11606 (N_11606,N_9190,N_10089);
xnor U11607 (N_11607,N_9937,N_9732);
and U11608 (N_11608,N_10247,N_9865);
xnor U11609 (N_11609,N_9059,N_10059);
xor U11610 (N_11610,N_9944,N_9663);
nand U11611 (N_11611,N_9361,N_9587);
or U11612 (N_11612,N_9383,N_9647);
nor U11613 (N_11613,N_9781,N_10469);
and U11614 (N_11614,N_9343,N_10251);
or U11615 (N_11615,N_9930,N_9534);
nor U11616 (N_11616,N_9756,N_9168);
nor U11617 (N_11617,N_9404,N_9801);
or U11618 (N_11618,N_10099,N_10181);
xor U11619 (N_11619,N_9397,N_10380);
or U11620 (N_11620,N_10020,N_9499);
xnor U11621 (N_11621,N_9385,N_9382);
or U11622 (N_11622,N_9739,N_9161);
xor U11623 (N_11623,N_10063,N_9813);
and U11624 (N_11624,N_9172,N_9928);
xor U11625 (N_11625,N_10409,N_9866);
or U11626 (N_11626,N_9841,N_9637);
xnor U11627 (N_11627,N_10435,N_9783);
and U11628 (N_11628,N_9784,N_9725);
xor U11629 (N_11629,N_9533,N_9172);
nand U11630 (N_11630,N_9444,N_9465);
xor U11631 (N_11631,N_9841,N_10412);
and U11632 (N_11632,N_10495,N_9263);
nand U11633 (N_11633,N_9413,N_10438);
and U11634 (N_11634,N_9439,N_9154);
and U11635 (N_11635,N_10113,N_9588);
and U11636 (N_11636,N_9429,N_10202);
xor U11637 (N_11637,N_9970,N_9484);
nor U11638 (N_11638,N_9443,N_9944);
nor U11639 (N_11639,N_9519,N_9603);
and U11640 (N_11640,N_10417,N_9688);
and U11641 (N_11641,N_10088,N_9639);
xnor U11642 (N_11642,N_9680,N_10281);
nand U11643 (N_11643,N_10090,N_9545);
nand U11644 (N_11644,N_9543,N_9630);
or U11645 (N_11645,N_10221,N_9848);
nand U11646 (N_11646,N_10459,N_10461);
and U11647 (N_11647,N_9165,N_9608);
and U11648 (N_11648,N_10344,N_9584);
and U11649 (N_11649,N_9998,N_9697);
nor U11650 (N_11650,N_10323,N_10019);
or U11651 (N_11651,N_9232,N_9597);
nand U11652 (N_11652,N_9029,N_10495);
or U11653 (N_11653,N_9783,N_9740);
and U11654 (N_11654,N_10130,N_9539);
nor U11655 (N_11655,N_10079,N_9358);
nand U11656 (N_11656,N_9763,N_9442);
and U11657 (N_11657,N_10193,N_10015);
nand U11658 (N_11658,N_9786,N_9207);
nor U11659 (N_11659,N_10386,N_9437);
xor U11660 (N_11660,N_9209,N_10394);
and U11661 (N_11661,N_9538,N_9208);
nand U11662 (N_11662,N_10029,N_10302);
nand U11663 (N_11663,N_9757,N_9474);
nand U11664 (N_11664,N_9696,N_9873);
nor U11665 (N_11665,N_10461,N_10016);
or U11666 (N_11666,N_9902,N_9027);
xnor U11667 (N_11667,N_9693,N_9156);
or U11668 (N_11668,N_9825,N_9493);
nor U11669 (N_11669,N_10413,N_9885);
xor U11670 (N_11670,N_9084,N_9883);
nand U11671 (N_11671,N_9859,N_10267);
xor U11672 (N_11672,N_9134,N_9698);
and U11673 (N_11673,N_9936,N_10012);
nor U11674 (N_11674,N_9243,N_9077);
nand U11675 (N_11675,N_10142,N_10265);
or U11676 (N_11676,N_9049,N_10208);
or U11677 (N_11677,N_10016,N_9113);
and U11678 (N_11678,N_9873,N_9902);
nand U11679 (N_11679,N_10109,N_10162);
xnor U11680 (N_11680,N_10168,N_10405);
nand U11681 (N_11681,N_9540,N_9854);
and U11682 (N_11682,N_10401,N_10460);
nor U11683 (N_11683,N_9545,N_9427);
nand U11684 (N_11684,N_10020,N_9892);
and U11685 (N_11685,N_9216,N_9894);
and U11686 (N_11686,N_10211,N_10147);
nor U11687 (N_11687,N_10120,N_10107);
nor U11688 (N_11688,N_9681,N_10407);
xor U11689 (N_11689,N_9002,N_10451);
and U11690 (N_11690,N_9686,N_10121);
xor U11691 (N_11691,N_9907,N_9013);
nor U11692 (N_11692,N_9361,N_10001);
and U11693 (N_11693,N_9048,N_10462);
or U11694 (N_11694,N_9269,N_10138);
and U11695 (N_11695,N_9582,N_10145);
or U11696 (N_11696,N_9168,N_9776);
and U11697 (N_11697,N_9074,N_9722);
or U11698 (N_11698,N_10392,N_9831);
nor U11699 (N_11699,N_9080,N_9339);
or U11700 (N_11700,N_9707,N_9037);
and U11701 (N_11701,N_9636,N_9741);
and U11702 (N_11702,N_10147,N_10112);
xnor U11703 (N_11703,N_10193,N_9684);
and U11704 (N_11704,N_9785,N_9484);
nor U11705 (N_11705,N_9651,N_9214);
xnor U11706 (N_11706,N_9302,N_10136);
nand U11707 (N_11707,N_9602,N_10108);
or U11708 (N_11708,N_9770,N_9051);
nor U11709 (N_11709,N_10005,N_9442);
or U11710 (N_11710,N_9884,N_9889);
nand U11711 (N_11711,N_10146,N_10029);
nand U11712 (N_11712,N_9410,N_10156);
and U11713 (N_11713,N_9860,N_10042);
xor U11714 (N_11714,N_10297,N_10486);
xnor U11715 (N_11715,N_9201,N_9997);
xnor U11716 (N_11716,N_10378,N_9287);
or U11717 (N_11717,N_10294,N_9896);
xor U11718 (N_11718,N_9229,N_9214);
nand U11719 (N_11719,N_9075,N_9432);
xnor U11720 (N_11720,N_10283,N_9476);
and U11721 (N_11721,N_10284,N_10292);
xor U11722 (N_11722,N_9965,N_10087);
nor U11723 (N_11723,N_9184,N_9989);
xnor U11724 (N_11724,N_9350,N_10100);
nor U11725 (N_11725,N_9328,N_10310);
and U11726 (N_11726,N_10379,N_9297);
xnor U11727 (N_11727,N_9918,N_9603);
or U11728 (N_11728,N_9464,N_9801);
or U11729 (N_11729,N_10138,N_9083);
and U11730 (N_11730,N_9719,N_9700);
nand U11731 (N_11731,N_9310,N_9908);
nand U11732 (N_11732,N_9069,N_10047);
xnor U11733 (N_11733,N_10106,N_10112);
or U11734 (N_11734,N_9746,N_9499);
and U11735 (N_11735,N_10004,N_9316);
and U11736 (N_11736,N_9083,N_9868);
nand U11737 (N_11737,N_9876,N_9408);
and U11738 (N_11738,N_9347,N_10098);
or U11739 (N_11739,N_9396,N_9708);
nand U11740 (N_11740,N_10313,N_9066);
nand U11741 (N_11741,N_10412,N_9536);
nor U11742 (N_11742,N_9784,N_10283);
xnor U11743 (N_11743,N_9550,N_9129);
nand U11744 (N_11744,N_10338,N_9920);
and U11745 (N_11745,N_9786,N_9269);
and U11746 (N_11746,N_9147,N_10202);
and U11747 (N_11747,N_9893,N_10327);
and U11748 (N_11748,N_9345,N_9869);
and U11749 (N_11749,N_9559,N_10086);
or U11750 (N_11750,N_9044,N_10121);
xnor U11751 (N_11751,N_10236,N_9090);
nand U11752 (N_11752,N_9080,N_9558);
xnor U11753 (N_11753,N_9664,N_10242);
xor U11754 (N_11754,N_9733,N_9322);
xnor U11755 (N_11755,N_10148,N_9635);
nor U11756 (N_11756,N_10405,N_9598);
xor U11757 (N_11757,N_9235,N_9625);
nand U11758 (N_11758,N_10028,N_9053);
or U11759 (N_11759,N_9440,N_9719);
nand U11760 (N_11760,N_9357,N_10386);
and U11761 (N_11761,N_9831,N_10087);
or U11762 (N_11762,N_9084,N_9909);
or U11763 (N_11763,N_9203,N_9911);
xnor U11764 (N_11764,N_9115,N_9866);
xnor U11765 (N_11765,N_10151,N_10124);
nand U11766 (N_11766,N_10027,N_9477);
nor U11767 (N_11767,N_10475,N_10104);
or U11768 (N_11768,N_9591,N_9434);
and U11769 (N_11769,N_10409,N_9138);
or U11770 (N_11770,N_9272,N_9776);
nor U11771 (N_11771,N_10491,N_10479);
nor U11772 (N_11772,N_10350,N_10078);
xor U11773 (N_11773,N_9252,N_9875);
nand U11774 (N_11774,N_9621,N_9216);
or U11775 (N_11775,N_9420,N_10082);
or U11776 (N_11776,N_9111,N_9374);
nand U11777 (N_11777,N_9372,N_9316);
or U11778 (N_11778,N_9423,N_9623);
nand U11779 (N_11779,N_9927,N_9584);
nor U11780 (N_11780,N_9394,N_9443);
or U11781 (N_11781,N_10222,N_9433);
or U11782 (N_11782,N_10154,N_9675);
nand U11783 (N_11783,N_9359,N_9319);
nand U11784 (N_11784,N_9831,N_9629);
nor U11785 (N_11785,N_9383,N_9337);
or U11786 (N_11786,N_10391,N_9375);
xnor U11787 (N_11787,N_9100,N_9076);
nand U11788 (N_11788,N_10392,N_9264);
nand U11789 (N_11789,N_9923,N_10186);
xor U11790 (N_11790,N_9099,N_9071);
nor U11791 (N_11791,N_9874,N_9441);
nor U11792 (N_11792,N_9360,N_9482);
or U11793 (N_11793,N_9094,N_10048);
nor U11794 (N_11794,N_9320,N_10045);
and U11795 (N_11795,N_10194,N_9781);
and U11796 (N_11796,N_10121,N_9235);
xor U11797 (N_11797,N_9828,N_9092);
xnor U11798 (N_11798,N_10040,N_9480);
nor U11799 (N_11799,N_9783,N_9801);
nor U11800 (N_11800,N_9880,N_9605);
xor U11801 (N_11801,N_10047,N_9876);
nor U11802 (N_11802,N_9684,N_9550);
nor U11803 (N_11803,N_9790,N_9038);
nand U11804 (N_11804,N_9187,N_10132);
or U11805 (N_11805,N_9982,N_9445);
nor U11806 (N_11806,N_9524,N_9642);
nor U11807 (N_11807,N_10490,N_10272);
and U11808 (N_11808,N_10262,N_9727);
nor U11809 (N_11809,N_9076,N_9291);
and U11810 (N_11810,N_9408,N_9441);
xnor U11811 (N_11811,N_9742,N_10038);
nand U11812 (N_11812,N_9891,N_9268);
nor U11813 (N_11813,N_9967,N_9445);
nand U11814 (N_11814,N_10491,N_9722);
nor U11815 (N_11815,N_9459,N_9916);
nand U11816 (N_11816,N_10363,N_9567);
xor U11817 (N_11817,N_9949,N_9758);
and U11818 (N_11818,N_10403,N_9525);
nor U11819 (N_11819,N_9303,N_10199);
or U11820 (N_11820,N_9830,N_9583);
and U11821 (N_11821,N_9274,N_10038);
and U11822 (N_11822,N_9386,N_9184);
nand U11823 (N_11823,N_9093,N_9123);
nand U11824 (N_11824,N_9956,N_10199);
xor U11825 (N_11825,N_9184,N_10258);
or U11826 (N_11826,N_10260,N_9058);
xor U11827 (N_11827,N_9745,N_10202);
or U11828 (N_11828,N_10088,N_9109);
nor U11829 (N_11829,N_9732,N_9963);
nor U11830 (N_11830,N_9353,N_9466);
and U11831 (N_11831,N_10469,N_10250);
nand U11832 (N_11832,N_10213,N_10348);
nand U11833 (N_11833,N_9395,N_9107);
xnor U11834 (N_11834,N_10188,N_9950);
and U11835 (N_11835,N_10491,N_9021);
nor U11836 (N_11836,N_10055,N_9738);
and U11837 (N_11837,N_9191,N_9263);
and U11838 (N_11838,N_10412,N_10457);
nor U11839 (N_11839,N_10114,N_10390);
xnor U11840 (N_11840,N_9484,N_9575);
nor U11841 (N_11841,N_9871,N_9907);
or U11842 (N_11842,N_9418,N_9365);
nor U11843 (N_11843,N_9475,N_9787);
or U11844 (N_11844,N_9142,N_9699);
and U11845 (N_11845,N_9625,N_9671);
nor U11846 (N_11846,N_9777,N_9016);
nor U11847 (N_11847,N_9740,N_9765);
and U11848 (N_11848,N_9500,N_9763);
and U11849 (N_11849,N_9975,N_9418);
or U11850 (N_11850,N_9330,N_9414);
and U11851 (N_11851,N_9218,N_10235);
nand U11852 (N_11852,N_9763,N_10356);
and U11853 (N_11853,N_9766,N_9893);
and U11854 (N_11854,N_9249,N_9035);
nor U11855 (N_11855,N_9424,N_9321);
xor U11856 (N_11856,N_9314,N_9676);
xor U11857 (N_11857,N_9353,N_9523);
and U11858 (N_11858,N_9256,N_10375);
nand U11859 (N_11859,N_10017,N_9305);
and U11860 (N_11860,N_9166,N_10427);
nand U11861 (N_11861,N_9541,N_9268);
xnor U11862 (N_11862,N_10024,N_9446);
or U11863 (N_11863,N_9452,N_9678);
nand U11864 (N_11864,N_9758,N_10335);
or U11865 (N_11865,N_10417,N_9574);
nor U11866 (N_11866,N_10389,N_9733);
xor U11867 (N_11867,N_10311,N_9152);
nand U11868 (N_11868,N_9333,N_9001);
and U11869 (N_11869,N_9075,N_9312);
and U11870 (N_11870,N_10008,N_10464);
xor U11871 (N_11871,N_9407,N_10327);
xor U11872 (N_11872,N_10313,N_9955);
xnor U11873 (N_11873,N_9393,N_10358);
nand U11874 (N_11874,N_9786,N_9650);
xor U11875 (N_11875,N_9680,N_9425);
and U11876 (N_11876,N_9245,N_10238);
nor U11877 (N_11877,N_9221,N_10298);
nor U11878 (N_11878,N_9780,N_9139);
xnor U11879 (N_11879,N_9639,N_9481);
nand U11880 (N_11880,N_9573,N_10429);
xor U11881 (N_11881,N_9006,N_10435);
or U11882 (N_11882,N_10190,N_9927);
xor U11883 (N_11883,N_9488,N_10228);
nand U11884 (N_11884,N_9525,N_9845);
or U11885 (N_11885,N_10087,N_9148);
and U11886 (N_11886,N_10497,N_9447);
nor U11887 (N_11887,N_9974,N_10284);
and U11888 (N_11888,N_9776,N_9845);
and U11889 (N_11889,N_9211,N_9918);
or U11890 (N_11890,N_9454,N_9753);
or U11891 (N_11891,N_10170,N_9552);
and U11892 (N_11892,N_9558,N_9117);
or U11893 (N_11893,N_9416,N_10183);
and U11894 (N_11894,N_9439,N_10461);
or U11895 (N_11895,N_10373,N_10055);
xnor U11896 (N_11896,N_9725,N_9999);
xnor U11897 (N_11897,N_9114,N_9497);
nor U11898 (N_11898,N_10337,N_9045);
and U11899 (N_11899,N_9288,N_9917);
nand U11900 (N_11900,N_9349,N_9458);
xnor U11901 (N_11901,N_9830,N_10426);
xnor U11902 (N_11902,N_9082,N_9037);
xnor U11903 (N_11903,N_9891,N_10180);
nand U11904 (N_11904,N_10087,N_9054);
and U11905 (N_11905,N_9505,N_9258);
nor U11906 (N_11906,N_10165,N_9966);
and U11907 (N_11907,N_9628,N_9766);
nand U11908 (N_11908,N_9569,N_9393);
or U11909 (N_11909,N_9148,N_9569);
or U11910 (N_11910,N_10411,N_10107);
nor U11911 (N_11911,N_9121,N_9048);
or U11912 (N_11912,N_9363,N_9729);
or U11913 (N_11913,N_9755,N_10162);
or U11914 (N_11914,N_9177,N_9724);
xor U11915 (N_11915,N_9394,N_9572);
or U11916 (N_11916,N_10373,N_10376);
and U11917 (N_11917,N_10423,N_9919);
xor U11918 (N_11918,N_9816,N_9173);
xor U11919 (N_11919,N_10052,N_9549);
and U11920 (N_11920,N_10055,N_9086);
nor U11921 (N_11921,N_10311,N_10304);
or U11922 (N_11922,N_9365,N_9475);
nand U11923 (N_11923,N_9204,N_9641);
nand U11924 (N_11924,N_10336,N_9885);
xor U11925 (N_11925,N_9775,N_9168);
xor U11926 (N_11926,N_9390,N_9687);
nand U11927 (N_11927,N_10016,N_9201);
nand U11928 (N_11928,N_9142,N_9406);
and U11929 (N_11929,N_9684,N_9006);
nand U11930 (N_11930,N_10292,N_9181);
nor U11931 (N_11931,N_9767,N_10477);
xor U11932 (N_11932,N_10203,N_9605);
nand U11933 (N_11933,N_9976,N_9998);
and U11934 (N_11934,N_9635,N_9555);
and U11935 (N_11935,N_9050,N_9902);
xor U11936 (N_11936,N_9021,N_9998);
nor U11937 (N_11937,N_10145,N_10029);
xor U11938 (N_11938,N_9622,N_9289);
or U11939 (N_11939,N_9083,N_10314);
nand U11940 (N_11940,N_10211,N_9547);
and U11941 (N_11941,N_10046,N_9416);
and U11942 (N_11942,N_10124,N_9922);
nor U11943 (N_11943,N_10053,N_9987);
or U11944 (N_11944,N_10036,N_10496);
nand U11945 (N_11945,N_9868,N_9525);
or U11946 (N_11946,N_10378,N_10388);
xor U11947 (N_11947,N_9668,N_9355);
xor U11948 (N_11948,N_9295,N_9177);
xnor U11949 (N_11949,N_10039,N_10136);
nor U11950 (N_11950,N_9505,N_10258);
or U11951 (N_11951,N_9605,N_9327);
xor U11952 (N_11952,N_9246,N_9212);
or U11953 (N_11953,N_10436,N_9223);
or U11954 (N_11954,N_10308,N_9728);
or U11955 (N_11955,N_10295,N_10166);
xor U11956 (N_11956,N_9489,N_10259);
xnor U11957 (N_11957,N_9068,N_9106);
and U11958 (N_11958,N_10473,N_9639);
nor U11959 (N_11959,N_10107,N_9379);
and U11960 (N_11960,N_10289,N_10224);
xor U11961 (N_11961,N_9012,N_9062);
nand U11962 (N_11962,N_10197,N_9587);
nor U11963 (N_11963,N_10215,N_9001);
nor U11964 (N_11964,N_9443,N_10254);
nor U11965 (N_11965,N_9174,N_9729);
nor U11966 (N_11966,N_9071,N_9685);
xor U11967 (N_11967,N_9167,N_9402);
and U11968 (N_11968,N_9906,N_10323);
nor U11969 (N_11969,N_10334,N_9315);
nor U11970 (N_11970,N_10058,N_9852);
and U11971 (N_11971,N_10072,N_9756);
or U11972 (N_11972,N_9745,N_9965);
nand U11973 (N_11973,N_10032,N_9726);
nand U11974 (N_11974,N_9967,N_10093);
nor U11975 (N_11975,N_10048,N_10401);
and U11976 (N_11976,N_9715,N_9859);
or U11977 (N_11977,N_9734,N_10142);
nor U11978 (N_11978,N_10399,N_9395);
nand U11979 (N_11979,N_9080,N_10177);
and U11980 (N_11980,N_9205,N_10252);
nor U11981 (N_11981,N_9348,N_10063);
xnor U11982 (N_11982,N_9983,N_9677);
xnor U11983 (N_11983,N_9839,N_9822);
nor U11984 (N_11984,N_9168,N_9256);
and U11985 (N_11985,N_9346,N_9748);
and U11986 (N_11986,N_9528,N_10460);
nand U11987 (N_11987,N_9710,N_10218);
nand U11988 (N_11988,N_10198,N_9887);
xor U11989 (N_11989,N_10076,N_10487);
and U11990 (N_11990,N_9515,N_10259);
or U11991 (N_11991,N_10447,N_10190);
nand U11992 (N_11992,N_10139,N_9269);
xnor U11993 (N_11993,N_10300,N_10346);
and U11994 (N_11994,N_9595,N_9176);
xor U11995 (N_11995,N_9799,N_10220);
nand U11996 (N_11996,N_9310,N_10405);
nand U11997 (N_11997,N_9993,N_9510);
and U11998 (N_11998,N_10021,N_10283);
xor U11999 (N_11999,N_9506,N_10149);
nor U12000 (N_12000,N_11258,N_11436);
nand U12001 (N_12001,N_11508,N_11214);
or U12002 (N_12002,N_10521,N_10835);
or U12003 (N_12003,N_11804,N_11105);
nand U12004 (N_12004,N_11148,N_10815);
and U12005 (N_12005,N_10853,N_11832);
and U12006 (N_12006,N_11530,N_11601);
xnor U12007 (N_12007,N_10593,N_11376);
nand U12008 (N_12008,N_10543,N_10505);
nor U12009 (N_12009,N_11224,N_10712);
nand U12010 (N_12010,N_11235,N_11317);
xor U12011 (N_12011,N_11864,N_11116);
or U12012 (N_12012,N_11468,N_11411);
xor U12013 (N_12013,N_11130,N_11218);
nand U12014 (N_12014,N_11519,N_11527);
or U12015 (N_12015,N_10807,N_11842);
or U12016 (N_12016,N_11573,N_11078);
and U12017 (N_12017,N_10889,N_11338);
and U12018 (N_12018,N_10918,N_11264);
and U12019 (N_12019,N_11337,N_10939);
and U12020 (N_12020,N_10869,N_11967);
xnor U12021 (N_12021,N_11268,N_11921);
xnor U12022 (N_12022,N_11675,N_11686);
or U12023 (N_12023,N_11551,N_11388);
nand U12024 (N_12024,N_11061,N_11090);
or U12025 (N_12025,N_11257,N_11498);
xor U12026 (N_12026,N_11941,N_11109);
xor U12027 (N_12027,N_10854,N_11205);
nor U12028 (N_12028,N_10502,N_11533);
and U12029 (N_12029,N_11641,N_11795);
nand U12030 (N_12030,N_11774,N_11415);
nor U12031 (N_12031,N_11696,N_11473);
nor U12032 (N_12032,N_11964,N_11299);
or U12033 (N_12033,N_11836,N_11475);
and U12034 (N_12034,N_11825,N_11757);
or U12035 (N_12035,N_11611,N_11986);
and U12036 (N_12036,N_11897,N_10604);
nand U12037 (N_12037,N_11555,N_10759);
xor U12038 (N_12038,N_11994,N_10898);
nand U12039 (N_12039,N_11894,N_11007);
nand U12040 (N_12040,N_10744,N_11561);
xnor U12041 (N_12041,N_10689,N_11820);
or U12042 (N_12042,N_10594,N_11386);
xor U12043 (N_12043,N_11673,N_11700);
or U12044 (N_12044,N_11588,N_11636);
and U12045 (N_12045,N_10784,N_10617);
and U12046 (N_12046,N_11187,N_10722);
nand U12047 (N_12047,N_10925,N_10978);
and U12048 (N_12048,N_10522,N_11068);
and U12049 (N_12049,N_11741,N_11311);
and U12050 (N_12050,N_10568,N_10945);
or U12051 (N_12051,N_10861,N_10799);
or U12052 (N_12052,N_10651,N_11401);
nand U12053 (N_12053,N_10739,N_11371);
nor U12054 (N_12054,N_10950,N_11694);
nor U12055 (N_12055,N_11069,N_10813);
or U12056 (N_12056,N_10782,N_11233);
nor U12057 (N_12057,N_11521,N_10652);
nor U12058 (N_12058,N_10922,N_11703);
and U12059 (N_12059,N_11926,N_11946);
nand U12060 (N_12060,N_11378,N_11279);
or U12061 (N_12061,N_11719,N_11310);
and U12062 (N_12062,N_11333,N_11639);
or U12063 (N_12063,N_11977,N_11975);
and U12064 (N_12064,N_11810,N_11502);
nand U12065 (N_12065,N_10921,N_11140);
nor U12066 (N_12066,N_10805,N_11306);
xnor U12067 (N_12067,N_10866,N_11443);
or U12068 (N_12068,N_10672,N_10542);
or U12069 (N_12069,N_10536,N_10724);
nor U12070 (N_12070,N_11709,N_10673);
nor U12071 (N_12071,N_10947,N_11195);
nand U12072 (N_12072,N_11623,N_11176);
xnor U12073 (N_12073,N_11330,N_11652);
xnor U12074 (N_12074,N_10880,N_10964);
and U12075 (N_12075,N_11746,N_10633);
and U12076 (N_12076,N_11331,N_11617);
xor U12077 (N_12077,N_11322,N_11245);
or U12078 (N_12078,N_10909,N_11228);
xor U12079 (N_12079,N_11984,N_11917);
xnor U12080 (N_12080,N_11285,N_11682);
or U12081 (N_12081,N_11458,N_11942);
nand U12082 (N_12082,N_11039,N_11165);
nor U12083 (N_12083,N_11324,N_11379);
nand U12084 (N_12084,N_11489,N_11188);
and U12085 (N_12085,N_11840,N_10506);
xnor U12086 (N_12086,N_10707,N_11113);
or U12087 (N_12087,N_11053,N_11363);
or U12088 (N_12088,N_11035,N_11036);
or U12089 (N_12089,N_10680,N_10579);
nand U12090 (N_12090,N_10641,N_10924);
nor U12091 (N_12091,N_11303,N_11427);
xor U12092 (N_12092,N_11341,N_11689);
nor U12093 (N_12093,N_10589,N_11824);
and U12094 (N_12094,N_11631,N_11387);
xor U12095 (N_12095,N_10840,N_11500);
and U12096 (N_12096,N_11275,N_11396);
nor U12097 (N_12097,N_11990,N_11978);
and U12098 (N_12098,N_10768,N_11438);
and U12099 (N_12099,N_11868,N_11626);
xnor U12100 (N_12100,N_11852,N_10914);
nand U12101 (N_12101,N_10546,N_11841);
xnor U12102 (N_12102,N_11229,N_11687);
nor U12103 (N_12103,N_10802,N_11449);
xnor U12104 (N_12104,N_10678,N_10573);
or U12105 (N_12105,N_11750,N_11143);
xnor U12106 (N_12106,N_11759,N_11645);
or U12107 (N_12107,N_11567,N_11129);
or U12108 (N_12108,N_11353,N_11848);
and U12109 (N_12109,N_10990,N_10740);
nor U12110 (N_12110,N_11422,N_11726);
or U12111 (N_12111,N_11585,N_11779);
xor U12112 (N_12112,N_11787,N_11723);
xnor U12113 (N_12113,N_10870,N_11507);
or U12114 (N_12114,N_11718,N_10826);
nor U12115 (N_12115,N_10586,N_10620);
and U12116 (N_12116,N_10953,N_11535);
nor U12117 (N_12117,N_10640,N_10555);
or U12118 (N_12118,N_11908,N_11592);
xor U12119 (N_12119,N_10609,N_11497);
nor U12120 (N_12120,N_11118,N_11531);
xor U12121 (N_12121,N_11951,N_11125);
nor U12122 (N_12122,N_10837,N_11866);
xor U12123 (N_12123,N_11448,N_11248);
xnor U12124 (N_12124,N_11861,N_11334);
nor U12125 (N_12125,N_11360,N_11123);
xor U12126 (N_12126,N_11442,N_10954);
or U12127 (N_12127,N_11809,N_11751);
nand U12128 (N_12128,N_10537,N_11604);
or U12129 (N_12129,N_11667,N_11242);
and U12130 (N_12130,N_11054,N_10725);
xor U12131 (N_12131,N_11083,N_11421);
and U12132 (N_12132,N_10734,N_11781);
or U12133 (N_12133,N_11895,N_10756);
nor U12134 (N_12134,N_11262,N_11393);
or U12135 (N_12135,N_11857,N_10694);
or U12136 (N_12136,N_11838,N_10550);
xor U12137 (N_12137,N_11528,N_11877);
xor U12138 (N_12138,N_10762,N_11407);
or U12139 (N_12139,N_11150,N_11738);
nand U12140 (N_12140,N_11156,N_11405);
and U12141 (N_12141,N_11451,N_11162);
xor U12142 (N_12142,N_11288,N_11822);
or U12143 (N_12143,N_11354,N_11426);
xnor U12144 (N_12144,N_11052,N_10871);
xnor U12145 (N_12145,N_11104,N_11831);
nand U12146 (N_12146,N_11370,N_11134);
and U12147 (N_12147,N_11615,N_11047);
nor U12148 (N_12148,N_10686,N_10966);
or U12149 (N_12149,N_11818,N_10750);
or U12150 (N_12150,N_11349,N_11979);
and U12151 (N_12151,N_11313,N_11119);
or U12152 (N_12152,N_10822,N_11766);
or U12153 (N_12153,N_11812,N_11901);
or U12154 (N_12154,N_11582,N_11352);
or U12155 (N_12155,N_11128,N_11513);
and U12156 (N_12156,N_10504,N_11999);
nor U12157 (N_12157,N_10597,N_11972);
xnor U12158 (N_12158,N_11111,N_10612);
nand U12159 (N_12159,N_11465,N_11762);
nor U12160 (N_12160,N_10570,N_10723);
nor U12161 (N_12161,N_11849,N_11587);
nor U12162 (N_12162,N_11676,N_11256);
xor U12163 (N_12163,N_11931,N_11291);
nor U12164 (N_12164,N_11860,N_11121);
nand U12165 (N_12165,N_10908,N_11169);
and U12166 (N_12166,N_11575,N_10749);
nand U12167 (N_12167,N_11705,N_11200);
nand U12168 (N_12168,N_11085,N_11879);
or U12169 (N_12169,N_10708,N_11525);
nor U12170 (N_12170,N_10703,N_11270);
and U12171 (N_12171,N_10995,N_11219);
nand U12172 (N_12172,N_11938,N_11568);
xor U12173 (N_12173,N_11115,N_10501);
or U12174 (N_12174,N_11876,N_11891);
xnor U12175 (N_12175,N_10821,N_11295);
or U12176 (N_12176,N_11058,N_11539);
nor U12177 (N_12177,N_11817,N_10600);
xnor U12178 (N_12178,N_11204,N_10529);
nand U12179 (N_12179,N_11996,N_11212);
xor U12180 (N_12180,N_10661,N_11347);
or U12181 (N_12181,N_10698,N_11292);
nor U12182 (N_12182,N_10659,N_11230);
nor U12183 (N_12183,N_10516,N_11127);
nand U12184 (N_12184,N_11412,N_10900);
xor U12185 (N_12185,N_10862,N_11905);
and U12186 (N_12186,N_11546,N_10713);
and U12187 (N_12187,N_11960,N_11179);
xnor U12188 (N_12188,N_11699,N_11114);
nor U12189 (N_12189,N_10763,N_11710);
nor U12190 (N_12190,N_10654,N_11314);
nand U12191 (N_12191,N_11494,N_11046);
or U12192 (N_12192,N_10719,N_11428);
nor U12193 (N_12193,N_11461,N_10704);
or U12194 (N_12194,N_11173,N_10977);
nor U12195 (N_12195,N_11470,N_11171);
nand U12196 (N_12196,N_11010,N_11981);
nand U12197 (N_12197,N_11610,N_11020);
nand U12198 (N_12198,N_11798,N_11492);
or U12199 (N_12199,N_10812,N_10872);
or U12200 (N_12200,N_11948,N_11348);
or U12201 (N_12201,N_10811,N_11080);
or U12202 (N_12202,N_10518,N_10688);
and U12203 (N_12203,N_11862,N_11903);
or U12204 (N_12204,N_11537,N_11563);
nor U12205 (N_12205,N_11032,N_11161);
and U12206 (N_12206,N_11987,N_11009);
xor U12207 (N_12207,N_11190,N_11736);
and U12208 (N_12208,N_10970,N_10904);
xnor U12209 (N_12209,N_11441,N_11289);
xnor U12210 (N_12210,N_10888,N_10669);
nand U12211 (N_12211,N_11957,N_11067);
nor U12212 (N_12212,N_10843,N_11029);
nand U12213 (N_12213,N_11778,N_11803);
nand U12214 (N_12214,N_11936,N_11909);
nor U12215 (N_12215,N_11425,N_11655);
nor U12216 (N_12216,N_10645,N_10991);
nand U12217 (N_12217,N_11924,N_11199);
or U12218 (N_12218,N_11012,N_10591);
xor U12219 (N_12219,N_11406,N_11579);
nor U12220 (N_12220,N_11139,N_11340);
nand U12221 (N_12221,N_11151,N_10779);
xor U12222 (N_12222,N_11087,N_11560);
xnor U12223 (N_12223,N_10683,N_10517);
nand U12224 (N_12224,N_10539,N_11439);
nor U12225 (N_12225,N_11079,N_10531);
xnor U12226 (N_12226,N_11328,N_10758);
and U12227 (N_12227,N_11577,N_11532);
or U12228 (N_12228,N_10877,N_11210);
nand U12229 (N_12229,N_10817,N_11088);
or U12230 (N_12230,N_10751,N_10974);
nor U12231 (N_12231,N_11512,N_10608);
and U12232 (N_12232,N_11496,N_10797);
and U12233 (N_12233,N_11761,N_11431);
xor U12234 (N_12234,N_10632,N_11594);
or U12235 (N_12235,N_11843,N_11095);
and U12236 (N_12236,N_11714,N_11770);
nor U12237 (N_12237,N_11707,N_11284);
nor U12238 (N_12238,N_11409,N_11932);
and U12239 (N_12239,N_11720,N_11410);
nor U12240 (N_12240,N_10735,N_11157);
or U12241 (N_12241,N_11074,N_11472);
and U12242 (N_12242,N_11137,N_11886);
xor U12243 (N_12243,N_11811,N_10775);
or U12244 (N_12244,N_11064,N_11293);
nand U12245 (N_12245,N_11627,N_11983);
xor U12246 (N_12246,N_11158,N_10728);
xor U12247 (N_12247,N_10733,N_11679);
or U12248 (N_12248,N_11316,N_10601);
and U12249 (N_12249,N_10985,N_11455);
nor U12250 (N_12250,N_10520,N_10796);
nand U12251 (N_12251,N_10684,N_11066);
xor U12252 (N_12252,N_11906,N_10527);
or U12253 (N_12253,N_11858,N_11395);
and U12254 (N_12254,N_11685,N_11380);
nor U12255 (N_12255,N_11101,N_11584);
nand U12256 (N_12256,N_10702,N_11359);
nor U12257 (N_12257,N_10780,N_11193);
nor U12258 (N_12258,N_11596,N_11106);
nor U12259 (N_12259,N_10687,N_10844);
or U12260 (N_12260,N_11706,N_10538);
nor U12261 (N_12261,N_10878,N_10653);
nand U12262 (N_12262,N_10814,N_10833);
or U12263 (N_12263,N_11375,N_11605);
or U12264 (N_12264,N_11806,N_10618);
xnor U12265 (N_12265,N_11944,N_11658);
nor U12266 (N_12266,N_11142,N_11730);
and U12267 (N_12267,N_10623,N_11612);
nand U12268 (N_12268,N_10923,N_11098);
nor U12269 (N_12269,N_11377,N_10544);
nor U12270 (N_12270,N_11267,N_11578);
or U12271 (N_12271,N_10852,N_11780);
xnor U12272 (N_12272,N_10530,N_11050);
nor U12273 (N_12273,N_10647,N_11929);
or U12274 (N_12274,N_11883,N_10806);
nor U12275 (N_12275,N_11246,N_10549);
nor U12276 (N_12276,N_11572,N_11011);
or U12277 (N_12277,N_11429,N_11044);
or U12278 (N_12278,N_11965,N_11756);
nand U12279 (N_12279,N_10690,N_11765);
or U12280 (N_12280,N_11261,N_11466);
xnor U12281 (N_12281,N_11342,N_11608);
xor U12282 (N_12282,N_11355,N_11834);
nand U12283 (N_12283,N_10790,N_10886);
nand U12284 (N_12284,N_10519,N_11164);
or U12285 (N_12285,N_10524,N_11005);
or U12286 (N_12286,N_11775,N_11453);
xor U12287 (N_12287,N_11589,N_10509);
or U12288 (N_12288,N_10746,N_11754);
xor U12289 (N_12289,N_10860,N_11786);
nand U12290 (N_12290,N_11599,N_10511);
and U12291 (N_12291,N_11097,N_10767);
nand U12292 (N_12292,N_10610,N_11110);
or U12293 (N_12293,N_11629,N_11251);
and U12294 (N_12294,N_11661,N_11571);
xor U12295 (N_12295,N_11628,N_11403);
nand U12296 (N_12296,N_11919,N_11159);
or U12297 (N_12297,N_10983,N_11417);
xor U12298 (N_12298,N_11548,N_11487);
and U12299 (N_12299,N_10629,N_11241);
nor U12300 (N_12300,N_10679,N_10658);
nand U12301 (N_12301,N_10582,N_11345);
nand U12302 (N_12302,N_11656,N_10644);
and U12303 (N_12303,N_10564,N_10829);
nor U12304 (N_12304,N_11928,N_10863);
xnor U12305 (N_12305,N_11748,N_11872);
xnor U12306 (N_12306,N_11554,N_10613);
nand U12307 (N_12307,N_11659,N_11025);
or U12308 (N_12308,N_10500,N_10783);
or U12309 (N_12309,N_11138,N_11691);
and U12310 (N_12310,N_11454,N_10956);
nor U12311 (N_12311,N_11911,N_10596);
nor U12312 (N_12312,N_11100,N_10699);
xor U12313 (N_12313,N_10742,N_11174);
nand U12314 (N_12314,N_11620,N_11398);
or U12315 (N_12315,N_10875,N_11201);
and U12316 (N_12316,N_11900,N_11447);
xor U12317 (N_12317,N_11501,N_11968);
and U12318 (N_12318,N_10607,N_11526);
and U12319 (N_12319,N_11935,N_10948);
xnor U12320 (N_12320,N_11096,N_11021);
xor U12321 (N_12321,N_11988,N_11553);
and U12322 (N_12322,N_10599,N_11969);
nor U12323 (N_12323,N_11499,N_11185);
nor U12324 (N_12324,N_11055,N_11493);
or U12325 (N_12325,N_11189,N_11690);
nand U12326 (N_12326,N_11504,N_11002);
nand U12327 (N_12327,N_11239,N_10532);
or U12328 (N_12328,N_11073,N_10588);
and U12329 (N_12329,N_11456,N_11305);
or U12330 (N_12330,N_10515,N_11638);
or U12331 (N_12331,N_11072,N_11597);
nor U12332 (N_12332,N_11662,N_10507);
and U12333 (N_12333,N_11024,N_11800);
or U12334 (N_12334,N_10973,N_11789);
nand U12335 (N_12335,N_11059,N_10913);
xnor U12336 (N_12336,N_11813,N_11191);
xnor U12337 (N_12337,N_11226,N_11013);
or U12338 (N_12338,N_11146,N_11767);
and U12339 (N_12339,N_10828,N_11595);
nand U12340 (N_12340,N_10598,N_10634);
nor U12341 (N_12341,N_10905,N_11819);
or U12342 (N_12342,N_11327,N_10576);
nor U12343 (N_12343,N_11048,N_11484);
xor U12344 (N_12344,N_10938,N_10748);
xnor U12345 (N_12345,N_11215,N_11445);
and U12346 (N_12346,N_11735,N_11529);
xnor U12347 (N_12347,N_11265,N_11593);
xor U12348 (N_12348,N_10585,N_11792);
and U12349 (N_12349,N_10789,N_11520);
xor U12350 (N_12350,N_10621,N_11287);
nor U12351 (N_12351,N_11920,N_10868);
xnor U12352 (N_12352,N_10741,N_11339);
and U12353 (N_12353,N_11263,N_11785);
nand U12354 (N_12354,N_10571,N_11853);
and U12355 (N_12355,N_11566,N_11829);
or U12356 (N_12356,N_11252,N_10794);
and U12357 (N_12357,N_10839,N_11701);
nor U12358 (N_12358,N_10916,N_11565);
xor U12359 (N_12359,N_11890,N_11351);
or U12360 (N_12360,N_11916,N_11372);
xnor U12361 (N_12361,N_11135,N_11414);
nor U12362 (N_12362,N_11168,N_11478);
nor U12363 (N_12363,N_11434,N_11037);
and U12364 (N_12364,N_11896,N_10876);
nor U12365 (N_12365,N_11049,N_11077);
nand U12366 (N_12366,N_10931,N_11297);
xor U12367 (N_12367,N_10615,N_11962);
nand U12368 (N_12368,N_11361,N_11556);
xnor U12369 (N_12369,N_11003,N_11249);
nand U12370 (N_12370,N_11060,N_11826);
or U12371 (N_12371,N_11618,N_11616);
nand U12372 (N_12372,N_10772,N_11231);
or U12373 (N_12373,N_11963,N_11885);
nor U12374 (N_12374,N_10584,N_10693);
nor U12375 (N_12375,N_10747,N_11488);
nor U12376 (N_12376,N_11286,N_11283);
nand U12377 (N_12377,N_10567,N_11126);
xor U12378 (N_12378,N_11300,N_10663);
xnor U12379 (N_12379,N_10562,N_10533);
nor U12380 (N_12380,N_11315,N_11713);
nor U12381 (N_12381,N_10930,N_10649);
and U12382 (N_12382,N_11621,N_11402);
xor U12383 (N_12383,N_10552,N_10765);
and U12384 (N_12384,N_11536,N_11390);
or U12385 (N_12385,N_10920,N_10874);
or U12386 (N_12386,N_11892,N_11301);
nand U12387 (N_12387,N_11332,N_10668);
nor U12388 (N_12388,N_11093,N_11178);
and U12389 (N_12389,N_11518,N_11132);
or U12390 (N_12390,N_11040,N_10984);
and U12391 (N_12391,N_11665,N_11477);
xor U12392 (N_12392,N_10910,N_11708);
or U12393 (N_12393,N_10626,N_11057);
and U12394 (N_12394,N_11144,N_11904);
xor U12395 (N_12395,N_10657,N_11859);
nand U12396 (N_12396,N_11271,N_10674);
nor U12397 (N_12397,N_11801,N_11590);
or U12398 (N_12398,N_10893,N_10541);
xnor U12399 (N_12399,N_11574,N_10513);
or U12400 (N_12400,N_10896,N_10580);
nor U12401 (N_12401,N_11383,N_11654);
or U12402 (N_12402,N_11084,N_11793);
or U12403 (N_12403,N_11506,N_10906);
nand U12404 (N_12404,N_10770,N_11211);
nor U12405 (N_12405,N_10718,N_11523);
or U12406 (N_12406,N_10720,N_11391);
and U12407 (N_12407,N_11298,N_11545);
nor U12408 (N_12408,N_11103,N_11490);
or U12409 (N_12409,N_11277,N_11019);
nor U12410 (N_12410,N_10932,N_10992);
and U12411 (N_12411,N_11273,N_10903);
and U12412 (N_12412,N_11145,N_11635);
nor U12413 (N_12413,N_10709,N_11408);
nor U12414 (N_12414,N_11304,N_11294);
xnor U12415 (N_12415,N_10838,N_10830);
and U12416 (N_12416,N_11915,N_11711);
xor U12417 (N_12417,N_10535,N_11399);
nand U12418 (N_12418,N_11515,N_10755);
xor U12419 (N_12419,N_11630,N_11882);
or U12420 (N_12420,N_11991,N_11668);
xnor U12421 (N_12421,N_11296,N_11516);
nor U12422 (N_12422,N_10897,N_11006);
or U12423 (N_12423,N_10561,N_11389);
or U12424 (N_12424,N_11244,N_11698);
xnor U12425 (N_12425,N_11870,N_10969);
or U12426 (N_12426,N_11091,N_10666);
or U12427 (N_12427,N_11544,N_11216);
nor U12428 (N_12428,N_11480,N_11954);
xnor U12429 (N_12429,N_11569,N_11839);
nand U12430 (N_12430,N_11649,N_10771);
nand U12431 (N_12431,N_11881,N_10655);
or U12432 (N_12432,N_10614,N_11949);
nand U12433 (N_12433,N_11336,N_11460);
nor U12434 (N_12434,N_11666,N_10660);
nand U12435 (N_12435,N_11182,N_11956);
or U12436 (N_12436,N_11647,N_10941);
nor U12437 (N_12437,N_11462,N_10986);
and U12438 (N_12438,N_10936,N_10656);
xnor U12439 (N_12439,N_11483,N_10882);
nor U12440 (N_12440,N_10793,N_10711);
or U12441 (N_12441,N_11683,N_10961);
nor U12442 (N_12442,N_11154,N_10899);
and U12443 (N_12443,N_11416,N_10671);
and U12444 (N_12444,N_11722,N_10757);
or U12445 (N_12445,N_11763,N_10976);
and U12446 (N_12446,N_10548,N_10534);
and U12447 (N_12447,N_11082,N_10846);
or U12448 (N_12448,N_11790,N_11744);
xnor U12449 (N_12449,N_11603,N_11481);
or U12450 (N_12450,N_11889,N_11815);
xor U12451 (N_12451,N_10760,N_11671);
nand U12452 (N_12452,N_10583,N_11446);
xor U12453 (N_12453,N_11833,N_10943);
nor U12454 (N_12454,N_11541,N_10551);
and U12455 (N_12455,N_11910,N_10745);
nand U12456 (N_12456,N_11232,N_11640);
nand U12457 (N_12457,N_11240,N_10818);
nand U12458 (N_12458,N_11643,N_11613);
xnor U12459 (N_12459,N_11381,N_10892);
and U12460 (N_12460,N_11657,N_11995);
and U12461 (N_12461,N_10628,N_11511);
nor U12462 (N_12462,N_11018,N_11642);
xor U12463 (N_12463,N_10957,N_11878);
xnor U12464 (N_12464,N_10692,N_10761);
xnor U12465 (N_12465,N_11221,N_11937);
nor U12466 (N_12466,N_10940,N_11576);
xnor U12467 (N_12467,N_10710,N_11733);
nand U12468 (N_12468,N_11914,N_11384);
xor U12469 (N_12469,N_10503,N_10752);
nor U12470 (N_12470,N_11695,N_11973);
nor U12471 (N_12471,N_10849,N_10685);
xnor U12472 (N_12472,N_11343,N_10949);
or U12473 (N_12473,N_11782,N_10885);
and U12474 (N_12474,N_10553,N_11653);
and U12475 (N_12475,N_11491,N_11867);
xnor U12476 (N_12476,N_11562,N_11607);
or U12477 (N_12477,N_11888,N_11681);
nand U12478 (N_12478,N_11042,N_11847);
nand U12479 (N_12479,N_11464,N_11747);
or U12480 (N_12480,N_10935,N_11828);
nand U12481 (N_12481,N_11043,N_10512);
nor U12482 (N_12482,N_10842,N_11259);
nand U12483 (N_12483,N_11606,N_11729);
and U12484 (N_12484,N_11209,N_11753);
and U12485 (N_12485,N_10791,N_11776);
xnor U12486 (N_12486,N_11958,N_11855);
and U12487 (N_12487,N_11837,N_11227);
and U12488 (N_12488,N_11547,N_10879);
and U12489 (N_12489,N_10616,N_11312);
or U12490 (N_12490,N_11930,N_11993);
and U12491 (N_12491,N_10737,N_11543);
nand U12492 (N_12492,N_11898,N_10894);
xnor U12493 (N_12493,N_10795,N_10631);
or U12494 (N_12494,N_11250,N_10556);
and U12495 (N_12495,N_10662,N_10982);
or U12496 (N_12496,N_10891,N_10559);
xor U12497 (N_12497,N_11236,N_10639);
or U12498 (N_12498,N_11773,N_11266);
nand U12499 (N_12499,N_10526,N_11764);
and U12500 (N_12500,N_11184,N_11133);
and U12501 (N_12501,N_11382,N_11457);
xnor U12502 (N_12502,N_10540,N_11581);
and U12503 (N_12503,N_11940,N_11194);
nand U12504 (N_12504,N_10731,N_10510);
nand U12505 (N_12505,N_11459,N_10971);
xnor U12506 (N_12506,N_11816,N_10836);
nand U12507 (N_12507,N_11147,N_11344);
and U12508 (N_12508,N_11945,N_11413);
and U12509 (N_12509,N_10774,N_10624);
nor U12510 (N_12510,N_10994,N_11622);
xnor U12511 (N_12511,N_11664,N_10851);
and U12512 (N_12512,N_11646,N_10525);
nand U12513 (N_12513,N_10958,N_11777);
xor U12514 (N_12514,N_11791,N_10798);
xnor U12515 (N_12515,N_11163,N_11369);
or U12516 (N_12516,N_11023,N_10727);
or U12517 (N_12517,N_11486,N_11208);
nor U12518 (N_12518,N_11749,N_11180);
or U12519 (N_12519,N_11452,N_11805);
and U12520 (N_12520,N_10873,N_10820);
xor U12521 (N_12521,N_10965,N_10809);
nor U12522 (N_12522,N_11835,N_11927);
or U12523 (N_12523,N_11959,N_11220);
and U12524 (N_12524,N_10827,N_11350);
xnor U12525 (N_12525,N_11444,N_11274);
or U12526 (N_12526,N_11902,N_11688);
nor U12527 (N_12527,N_10960,N_10787);
nand U12528 (N_12528,N_10706,N_11014);
xor U12529 (N_12529,N_10587,N_10831);
or U12530 (N_12530,N_11160,N_11075);
nor U12531 (N_12531,N_11318,N_10590);
nor U12532 (N_12532,N_10732,N_11329);
and U12533 (N_12533,N_11364,N_11794);
and U12534 (N_12534,N_11614,N_10676);
or U12535 (N_12535,N_10636,N_11557);
nand U12536 (N_12536,N_11953,N_10895);
nor U12537 (N_12537,N_11712,N_11015);
and U12538 (N_12538,N_10804,N_11223);
nor U12539 (N_12539,N_11056,N_11362);
xnor U12540 (N_12540,N_10638,N_11112);
or U12541 (N_12541,N_10946,N_11739);
and U12542 (N_12542,N_10738,N_11392);
and U12543 (N_12543,N_11419,N_10781);
xor U12544 (N_12544,N_11998,N_10721);
or U12545 (N_12545,N_11827,N_10574);
and U12546 (N_12546,N_11365,N_11648);
or U12547 (N_12547,N_10776,N_11206);
or U12548 (N_12548,N_11394,N_10753);
nand U12549 (N_12549,N_11192,N_11884);
or U12550 (N_12550,N_11071,N_11684);
nand U12551 (N_12551,N_11923,N_11674);
nor U12552 (N_12552,N_11326,N_11846);
nor U12553 (N_12553,N_11213,N_11971);
xnor U12554 (N_12554,N_10834,N_11717);
nor U12555 (N_12555,N_11081,N_11070);
and U12556 (N_12556,N_10917,N_11469);
nand U12557 (N_12557,N_10605,N_10792);
nor U12558 (N_12558,N_10808,N_11089);
and U12559 (N_12559,N_10927,N_10801);
nor U12560 (N_12560,N_11913,N_11821);
nor U12561 (N_12561,N_11814,N_10715);
and U12562 (N_12562,N_11505,N_10595);
or U12563 (N_12563,N_10998,N_10902);
and U12564 (N_12564,N_10602,N_11918);
and U12565 (N_12565,N_11474,N_11400);
xor U12566 (N_12566,N_10508,N_11122);
xor U12567 (N_12567,N_10566,N_10968);
or U12568 (N_12568,N_10635,N_11323);
xor U12569 (N_12569,N_11772,N_10942);
or U12570 (N_12570,N_11702,N_11272);
or U12571 (N_12571,N_11358,N_11933);
xor U12572 (N_12572,N_11385,N_10558);
nand U12573 (N_12573,N_11437,N_11045);
nand U12574 (N_12574,N_11022,N_11247);
xor U12575 (N_12575,N_10858,N_11278);
and U12576 (N_12576,N_10743,N_11253);
xnor U12577 (N_12577,N_11760,N_10824);
nor U12578 (N_12578,N_10816,N_11207);
nor U12579 (N_12579,N_10883,N_10667);
or U12580 (N_12580,N_10554,N_11865);
nand U12581 (N_12581,N_10850,N_11307);
xnor U12582 (N_12582,N_10944,N_11788);
nand U12583 (N_12583,N_10845,N_11619);
nand U12584 (N_12584,N_11716,N_11424);
nor U12585 (N_12585,N_10865,N_11514);
and U12586 (N_12586,N_10592,N_11309);
xor U12587 (N_12587,N_11583,N_10810);
nand U12588 (N_12588,N_11797,N_10773);
and U12589 (N_12589,N_10786,N_11509);
and U12590 (N_12590,N_11644,N_10980);
or U12591 (N_12591,N_10847,N_11107);
or U12592 (N_12592,N_10857,N_11041);
or U12593 (N_12593,N_11875,N_11238);
and U12594 (N_12594,N_10643,N_11534);
or U12595 (N_12595,N_11752,N_11680);
nor U12596 (N_12596,N_11731,N_10929);
or U12597 (N_12597,N_11542,N_11989);
nor U12598 (N_12598,N_11034,N_10681);
xor U12599 (N_12599,N_10545,N_10864);
or U12600 (N_12600,N_11108,N_11260);
nor U12601 (N_12601,N_11471,N_11368);
and U12602 (N_12602,N_10975,N_10716);
xor U12603 (N_12603,N_11784,N_11724);
or U12604 (N_12604,N_10993,N_11255);
xor U12605 (N_12605,N_11570,N_11136);
nand U12606 (N_12606,N_11734,N_10578);
and U12607 (N_12607,N_11692,N_11149);
nor U12608 (N_12608,N_11198,N_11925);
xnor U12609 (N_12609,N_10979,N_10856);
xnor U12610 (N_12610,N_11863,N_10557);
and U12611 (N_12611,N_11650,N_11177);
xnor U12612 (N_12612,N_11704,N_11482);
nand U12613 (N_12613,N_10611,N_11290);
nand U12614 (N_12614,N_10928,N_11065);
nand U12615 (N_12615,N_11552,N_11030);
and U12616 (N_12616,N_11463,N_11167);
and U12617 (N_12617,N_10766,N_11302);
and U12618 (N_12618,N_11558,N_11076);
nor U12619 (N_12619,N_11001,N_11099);
xnor U12620 (N_12620,N_10581,N_10547);
or U12621 (N_12621,N_10823,N_11966);
nor U12622 (N_12622,N_11016,N_10696);
or U12623 (N_12623,N_11715,N_11856);
nor U12624 (N_12624,N_11524,N_11893);
nand U12625 (N_12625,N_11970,N_11120);
nand U12626 (N_12626,N_11321,N_11672);
xnor U12627 (N_12627,N_11141,N_11181);
and U12628 (N_12628,N_11743,N_11063);
or U12629 (N_12629,N_11155,N_11669);
or U12630 (N_12630,N_11559,N_10700);
xnor U12631 (N_12631,N_11017,N_11243);
and U12632 (N_12632,N_10569,N_10560);
nand U12633 (N_12633,N_11008,N_11907);
nor U12634 (N_12634,N_11950,N_11922);
or U12635 (N_12635,N_11550,N_10987);
and U12636 (N_12636,N_10695,N_11591);
nand U12637 (N_12637,N_10890,N_11325);
nor U12638 (N_12638,N_11732,N_11033);
nand U12639 (N_12639,N_11728,N_10981);
xnor U12640 (N_12640,N_11026,N_10952);
nor U12641 (N_12641,N_11830,N_10937);
xnor U12642 (N_12642,N_10627,N_10729);
nand U12643 (N_12643,N_11912,N_11000);
nand U12644 (N_12644,N_11467,N_11980);
and U12645 (N_12645,N_11280,N_10800);
nand U12646 (N_12646,N_11538,N_11237);
or U12647 (N_12647,N_10717,N_10785);
and U12648 (N_12648,N_11598,N_10951);
or U12649 (N_12649,N_11225,N_11976);
or U12650 (N_12650,N_10972,N_10884);
nand U12651 (N_12651,N_11004,N_10705);
and U12652 (N_12652,N_11783,N_10650);
and U12653 (N_12653,N_11432,N_11540);
nor U12654 (N_12654,N_10777,N_11586);
or U12655 (N_12655,N_11366,N_10901);
or U12656 (N_12656,N_11102,N_10514);
nor U12657 (N_12657,N_10934,N_10637);
or U12658 (N_12658,N_10887,N_11503);
xnor U12659 (N_12659,N_10625,N_11397);
and U12660 (N_12660,N_11479,N_10603);
nor U12661 (N_12661,N_11028,N_11485);
and U12662 (N_12662,N_10963,N_10682);
and U12663 (N_12663,N_10577,N_11153);
nand U12664 (N_12664,N_10726,N_11880);
or U12665 (N_12665,N_10962,N_11276);
xor U12666 (N_12666,N_11697,N_10565);
xnor U12667 (N_12667,N_10642,N_11367);
and U12668 (N_12668,N_10881,N_11771);
nand U12669 (N_12669,N_11660,N_11952);
or U12670 (N_12670,N_10630,N_11196);
or U12671 (N_12671,N_11282,N_11740);
and U12672 (N_12672,N_11721,N_11742);
nor U12673 (N_12673,N_10572,N_11845);
and U12674 (N_12674,N_11038,N_11281);
nor U12675 (N_12675,N_11420,N_10575);
or U12676 (N_12676,N_11166,N_11869);
nand U12677 (N_12677,N_11637,N_11476);
or U12678 (N_12678,N_10867,N_11678);
nor U12679 (N_12679,N_11899,N_11939);
nor U12680 (N_12680,N_10911,N_10907);
nor U12681 (N_12681,N_11887,N_11651);
xnor U12682 (N_12682,N_10677,N_11423);
and U12683 (N_12683,N_10848,N_11131);
and U12684 (N_12684,N_11632,N_11495);
or U12685 (N_12685,N_10528,N_11997);
and U12686 (N_12686,N_10730,N_11677);
or U12687 (N_12687,N_11985,N_11624);
or U12688 (N_12688,N_10989,N_11440);
nand U12689 (N_12689,N_11955,N_11269);
xor U12690 (N_12690,N_10997,N_11357);
nand U12691 (N_12691,N_10714,N_11152);
xor U12692 (N_12692,N_11943,N_11609);
or U12693 (N_12693,N_11086,N_10855);
or U12694 (N_12694,N_10803,N_11808);
nand U12695 (N_12695,N_11725,N_11693);
and U12696 (N_12696,N_10926,N_11117);
nor U12697 (N_12697,N_11796,N_11799);
and U12698 (N_12698,N_11124,N_11450);
xnor U12699 (N_12699,N_11758,N_11418);
or U12700 (N_12700,N_10736,N_11373);
xor U12701 (N_12701,N_11850,N_11768);
or U12702 (N_12702,N_11092,N_10664);
xnor U12703 (N_12703,N_11308,N_10915);
xor U12704 (N_12704,N_10919,N_11961);
nand U12705 (N_12705,N_10648,N_10691);
and U12706 (N_12706,N_11745,N_11335);
xnor U12707 (N_12707,N_11346,N_11992);
or U12708 (N_12708,N_10933,N_10646);
nand U12709 (N_12709,N_11974,N_11737);
nor U12710 (N_12710,N_10754,N_11802);
nand U12711 (N_12711,N_11320,N_11769);
xor U12712 (N_12712,N_11510,N_10955);
and U12713 (N_12713,N_10670,N_10778);
nor U12714 (N_12714,N_11430,N_10622);
nand U12715 (N_12715,N_11854,N_11186);
nand U12716 (N_12716,N_11874,N_11602);
nor U12717 (N_12717,N_10832,N_10769);
nand U12718 (N_12718,N_10859,N_11823);
or U12719 (N_12719,N_11947,N_10959);
nor U12720 (N_12720,N_11175,N_11183);
or U12721 (N_12721,N_11634,N_11051);
and U12722 (N_12722,N_10665,N_11217);
and U12723 (N_12723,N_11433,N_11670);
and U12724 (N_12724,N_11934,N_11522);
or U12725 (N_12725,N_10606,N_11356);
nor U12726 (N_12726,N_10841,N_11549);
nand U12727 (N_12727,N_10563,N_11873);
nor U12728 (N_12728,N_10523,N_11172);
or U12729 (N_12729,N_11625,N_11663);
or U12730 (N_12730,N_10967,N_10988);
nor U12731 (N_12731,N_10675,N_11564);
and U12732 (N_12732,N_11027,N_10912);
nor U12733 (N_12733,N_11435,N_10764);
nand U12734 (N_12734,N_11374,N_11727);
nand U12735 (N_12735,N_11202,N_10788);
xor U12736 (N_12736,N_11600,N_11319);
nand U12737 (N_12737,N_11851,N_11197);
nand U12738 (N_12738,N_11982,N_11254);
or U12739 (N_12739,N_11517,N_11844);
nand U12740 (N_12740,N_10819,N_11203);
and U12741 (N_12741,N_11580,N_11170);
and U12742 (N_12742,N_10619,N_11633);
and U12743 (N_12743,N_11062,N_11234);
and U12744 (N_12744,N_11755,N_11404);
nor U12745 (N_12745,N_11031,N_10996);
and U12746 (N_12746,N_10999,N_11094);
nor U12747 (N_12747,N_10697,N_10701);
nand U12748 (N_12748,N_10825,N_11871);
nand U12749 (N_12749,N_11222,N_11807);
or U12750 (N_12750,N_11639,N_11393);
or U12751 (N_12751,N_10875,N_11286);
and U12752 (N_12752,N_11958,N_10620);
nor U12753 (N_12753,N_11672,N_11056);
nor U12754 (N_12754,N_11369,N_11142);
nor U12755 (N_12755,N_11912,N_10875);
xnor U12756 (N_12756,N_11172,N_11946);
and U12757 (N_12757,N_11465,N_10541);
nand U12758 (N_12758,N_11289,N_10566);
or U12759 (N_12759,N_10817,N_11968);
nor U12760 (N_12760,N_10992,N_10848);
or U12761 (N_12761,N_11718,N_10747);
and U12762 (N_12762,N_11804,N_11689);
nand U12763 (N_12763,N_11190,N_10584);
nor U12764 (N_12764,N_10794,N_10798);
nor U12765 (N_12765,N_11632,N_11128);
and U12766 (N_12766,N_11816,N_11218);
nand U12767 (N_12767,N_11453,N_10778);
and U12768 (N_12768,N_11937,N_11511);
or U12769 (N_12769,N_11580,N_11376);
or U12770 (N_12770,N_11130,N_11469);
xnor U12771 (N_12771,N_11006,N_11856);
nand U12772 (N_12772,N_11314,N_11455);
xor U12773 (N_12773,N_11215,N_11129);
or U12774 (N_12774,N_11732,N_11114);
xnor U12775 (N_12775,N_11222,N_11977);
nor U12776 (N_12776,N_11928,N_10886);
nor U12777 (N_12777,N_11661,N_11021);
and U12778 (N_12778,N_11028,N_11834);
or U12779 (N_12779,N_11496,N_11079);
or U12780 (N_12780,N_11261,N_10549);
and U12781 (N_12781,N_11768,N_11740);
or U12782 (N_12782,N_11549,N_11632);
and U12783 (N_12783,N_10627,N_11108);
or U12784 (N_12784,N_10770,N_11917);
nand U12785 (N_12785,N_11807,N_11378);
nor U12786 (N_12786,N_11962,N_11935);
and U12787 (N_12787,N_10923,N_11878);
nand U12788 (N_12788,N_10963,N_10946);
xnor U12789 (N_12789,N_11417,N_10868);
xnor U12790 (N_12790,N_10754,N_11266);
and U12791 (N_12791,N_11634,N_11419);
and U12792 (N_12792,N_11481,N_11687);
or U12793 (N_12793,N_11676,N_11033);
and U12794 (N_12794,N_11579,N_11107);
xor U12795 (N_12795,N_11461,N_11773);
nand U12796 (N_12796,N_10706,N_10592);
nor U12797 (N_12797,N_10902,N_11791);
nand U12798 (N_12798,N_10771,N_11892);
nor U12799 (N_12799,N_11315,N_10860);
and U12800 (N_12800,N_10790,N_11796);
and U12801 (N_12801,N_11472,N_11248);
nor U12802 (N_12802,N_11478,N_11050);
xnor U12803 (N_12803,N_10883,N_11417);
nor U12804 (N_12804,N_11417,N_11032);
and U12805 (N_12805,N_10795,N_10793);
or U12806 (N_12806,N_11513,N_10735);
nor U12807 (N_12807,N_10641,N_11720);
and U12808 (N_12808,N_11501,N_11434);
or U12809 (N_12809,N_10661,N_10914);
or U12810 (N_12810,N_10675,N_10945);
and U12811 (N_12811,N_11340,N_11722);
nor U12812 (N_12812,N_11352,N_11884);
and U12813 (N_12813,N_11741,N_11681);
nor U12814 (N_12814,N_11408,N_11068);
nand U12815 (N_12815,N_10675,N_11372);
xnor U12816 (N_12816,N_11074,N_11217);
and U12817 (N_12817,N_10870,N_11262);
or U12818 (N_12818,N_11110,N_11189);
nor U12819 (N_12819,N_11331,N_10593);
nor U12820 (N_12820,N_10716,N_11882);
and U12821 (N_12821,N_11749,N_11341);
or U12822 (N_12822,N_11482,N_10834);
and U12823 (N_12823,N_11364,N_11957);
or U12824 (N_12824,N_11999,N_11313);
xnor U12825 (N_12825,N_11256,N_10539);
xnor U12826 (N_12826,N_10837,N_11727);
nand U12827 (N_12827,N_11865,N_10711);
and U12828 (N_12828,N_11011,N_11911);
nor U12829 (N_12829,N_11163,N_11145);
and U12830 (N_12830,N_11311,N_11415);
nand U12831 (N_12831,N_10599,N_10820);
nor U12832 (N_12832,N_11204,N_10734);
nand U12833 (N_12833,N_10845,N_11950);
nand U12834 (N_12834,N_10907,N_11356);
xnor U12835 (N_12835,N_11324,N_11655);
nand U12836 (N_12836,N_11082,N_10703);
and U12837 (N_12837,N_11261,N_10764);
xnor U12838 (N_12838,N_10682,N_10701);
xor U12839 (N_12839,N_10554,N_10708);
nand U12840 (N_12840,N_10612,N_11478);
and U12841 (N_12841,N_11725,N_11579);
nand U12842 (N_12842,N_10571,N_11864);
nor U12843 (N_12843,N_11078,N_11622);
nor U12844 (N_12844,N_10820,N_11566);
xnor U12845 (N_12845,N_11034,N_10571);
nand U12846 (N_12846,N_10515,N_10592);
and U12847 (N_12847,N_11946,N_10635);
nand U12848 (N_12848,N_11667,N_10690);
and U12849 (N_12849,N_11252,N_10982);
and U12850 (N_12850,N_11355,N_10925);
xor U12851 (N_12851,N_10537,N_11912);
nand U12852 (N_12852,N_11170,N_11136);
xor U12853 (N_12853,N_11918,N_10557);
nand U12854 (N_12854,N_10840,N_11190);
nand U12855 (N_12855,N_10521,N_10708);
or U12856 (N_12856,N_10825,N_11003);
and U12857 (N_12857,N_11822,N_11496);
or U12858 (N_12858,N_11001,N_11451);
and U12859 (N_12859,N_10757,N_11121);
or U12860 (N_12860,N_11771,N_10599);
nor U12861 (N_12861,N_10720,N_10723);
xor U12862 (N_12862,N_11036,N_10580);
xnor U12863 (N_12863,N_11414,N_11138);
nor U12864 (N_12864,N_11747,N_11900);
nand U12865 (N_12865,N_11010,N_11409);
or U12866 (N_12866,N_10503,N_10794);
nand U12867 (N_12867,N_11691,N_10581);
nor U12868 (N_12868,N_11865,N_10567);
or U12869 (N_12869,N_10621,N_10601);
or U12870 (N_12870,N_11888,N_11484);
nor U12871 (N_12871,N_10889,N_11587);
xnor U12872 (N_12872,N_11788,N_11265);
nor U12873 (N_12873,N_10921,N_10508);
nand U12874 (N_12874,N_10617,N_11698);
or U12875 (N_12875,N_10713,N_11190);
nand U12876 (N_12876,N_11947,N_10894);
nand U12877 (N_12877,N_11701,N_11585);
or U12878 (N_12878,N_11542,N_11537);
xnor U12879 (N_12879,N_11482,N_11125);
and U12880 (N_12880,N_11618,N_10597);
and U12881 (N_12881,N_11324,N_11873);
xor U12882 (N_12882,N_11347,N_11374);
nand U12883 (N_12883,N_11181,N_11688);
xor U12884 (N_12884,N_11957,N_10831);
xor U12885 (N_12885,N_11199,N_11940);
nor U12886 (N_12886,N_11369,N_11677);
and U12887 (N_12887,N_10922,N_11349);
xor U12888 (N_12888,N_10596,N_11018);
xnor U12889 (N_12889,N_11114,N_11186);
or U12890 (N_12890,N_11708,N_11907);
nor U12891 (N_12891,N_10653,N_11922);
or U12892 (N_12892,N_11436,N_11483);
or U12893 (N_12893,N_11538,N_11568);
or U12894 (N_12894,N_11185,N_11250);
xor U12895 (N_12895,N_11072,N_11722);
nor U12896 (N_12896,N_11310,N_10510);
or U12897 (N_12897,N_11132,N_10573);
or U12898 (N_12898,N_11211,N_10926);
nand U12899 (N_12899,N_11435,N_11860);
xor U12900 (N_12900,N_11234,N_10847);
and U12901 (N_12901,N_11271,N_11296);
and U12902 (N_12902,N_11299,N_10643);
or U12903 (N_12903,N_11773,N_11514);
xnor U12904 (N_12904,N_11170,N_11956);
nor U12905 (N_12905,N_11022,N_11543);
or U12906 (N_12906,N_11176,N_10593);
or U12907 (N_12907,N_10973,N_11337);
and U12908 (N_12908,N_11229,N_11110);
and U12909 (N_12909,N_10785,N_11982);
nand U12910 (N_12910,N_11011,N_11744);
xor U12911 (N_12911,N_11037,N_11052);
and U12912 (N_12912,N_11409,N_11865);
xor U12913 (N_12913,N_10723,N_11896);
nor U12914 (N_12914,N_11907,N_10734);
nand U12915 (N_12915,N_10641,N_10779);
nor U12916 (N_12916,N_11357,N_11819);
or U12917 (N_12917,N_11091,N_10601);
nand U12918 (N_12918,N_11839,N_11083);
nand U12919 (N_12919,N_11492,N_11834);
nor U12920 (N_12920,N_10848,N_10644);
and U12921 (N_12921,N_11696,N_10842);
nor U12922 (N_12922,N_11663,N_10881);
xor U12923 (N_12923,N_10645,N_11205);
and U12924 (N_12924,N_11956,N_11437);
nor U12925 (N_12925,N_10893,N_11980);
nor U12926 (N_12926,N_10926,N_11493);
nor U12927 (N_12927,N_10862,N_11136);
nand U12928 (N_12928,N_11052,N_11148);
nor U12929 (N_12929,N_11086,N_11204);
and U12930 (N_12930,N_10997,N_10572);
nor U12931 (N_12931,N_10708,N_11021);
and U12932 (N_12932,N_11108,N_11729);
and U12933 (N_12933,N_11866,N_11460);
and U12934 (N_12934,N_10661,N_11695);
or U12935 (N_12935,N_11653,N_11586);
or U12936 (N_12936,N_11543,N_11657);
nand U12937 (N_12937,N_11535,N_10616);
and U12938 (N_12938,N_11628,N_11574);
and U12939 (N_12939,N_11495,N_11656);
and U12940 (N_12940,N_10916,N_10897);
or U12941 (N_12941,N_11849,N_10992);
nor U12942 (N_12942,N_11366,N_11597);
and U12943 (N_12943,N_10925,N_11813);
or U12944 (N_12944,N_11586,N_11035);
xor U12945 (N_12945,N_11441,N_10780);
xnor U12946 (N_12946,N_11593,N_11868);
nand U12947 (N_12947,N_11850,N_11668);
and U12948 (N_12948,N_10638,N_10831);
and U12949 (N_12949,N_11184,N_11736);
nand U12950 (N_12950,N_11157,N_11386);
or U12951 (N_12951,N_11300,N_11182);
and U12952 (N_12952,N_11051,N_11832);
nand U12953 (N_12953,N_10720,N_11938);
or U12954 (N_12954,N_11996,N_11008);
xor U12955 (N_12955,N_11368,N_11389);
or U12956 (N_12956,N_11389,N_10888);
and U12957 (N_12957,N_11234,N_11510);
nor U12958 (N_12958,N_11926,N_11475);
nor U12959 (N_12959,N_10995,N_11690);
or U12960 (N_12960,N_10773,N_11173);
nand U12961 (N_12961,N_11756,N_11290);
and U12962 (N_12962,N_10891,N_10715);
nand U12963 (N_12963,N_11329,N_10845);
or U12964 (N_12964,N_10683,N_10946);
or U12965 (N_12965,N_11694,N_11535);
and U12966 (N_12966,N_10553,N_11405);
nand U12967 (N_12967,N_11406,N_10747);
or U12968 (N_12968,N_11753,N_11860);
nor U12969 (N_12969,N_10667,N_11184);
xnor U12970 (N_12970,N_10897,N_11572);
nand U12971 (N_12971,N_11370,N_11556);
nor U12972 (N_12972,N_11215,N_11994);
xnor U12973 (N_12973,N_11598,N_11638);
xnor U12974 (N_12974,N_11966,N_11033);
and U12975 (N_12975,N_11567,N_11640);
xnor U12976 (N_12976,N_11576,N_11088);
xor U12977 (N_12977,N_11258,N_11983);
or U12978 (N_12978,N_11218,N_11453);
nand U12979 (N_12979,N_10926,N_11990);
and U12980 (N_12980,N_11882,N_10596);
and U12981 (N_12981,N_11180,N_11096);
or U12982 (N_12982,N_11987,N_11407);
or U12983 (N_12983,N_10645,N_10723);
nand U12984 (N_12984,N_11793,N_11910);
xnor U12985 (N_12985,N_11885,N_10818);
and U12986 (N_12986,N_11088,N_11715);
or U12987 (N_12987,N_11632,N_11451);
and U12988 (N_12988,N_10943,N_11717);
nand U12989 (N_12989,N_10831,N_11847);
or U12990 (N_12990,N_10602,N_11169);
nand U12991 (N_12991,N_10719,N_10863);
nor U12992 (N_12992,N_11115,N_11398);
or U12993 (N_12993,N_10872,N_11271);
nand U12994 (N_12994,N_11637,N_10974);
nor U12995 (N_12995,N_10825,N_10944);
nand U12996 (N_12996,N_10692,N_11558);
xor U12997 (N_12997,N_10958,N_11535);
nor U12998 (N_12998,N_11831,N_11187);
nor U12999 (N_12999,N_10584,N_10757);
and U13000 (N_13000,N_10548,N_11616);
nor U13001 (N_13001,N_11955,N_10858);
xnor U13002 (N_13002,N_11335,N_10969);
and U13003 (N_13003,N_11832,N_11843);
nand U13004 (N_13004,N_11311,N_11889);
nand U13005 (N_13005,N_11143,N_11014);
or U13006 (N_13006,N_10669,N_11612);
and U13007 (N_13007,N_11642,N_11824);
nand U13008 (N_13008,N_11558,N_10703);
and U13009 (N_13009,N_10503,N_11367);
nor U13010 (N_13010,N_11850,N_10938);
and U13011 (N_13011,N_11615,N_11451);
nor U13012 (N_13012,N_11812,N_11434);
xor U13013 (N_13013,N_11592,N_11206);
nor U13014 (N_13014,N_11750,N_11621);
and U13015 (N_13015,N_11921,N_11428);
xor U13016 (N_13016,N_11925,N_10890);
nand U13017 (N_13017,N_11300,N_10696);
or U13018 (N_13018,N_11132,N_11525);
xor U13019 (N_13019,N_11891,N_11837);
or U13020 (N_13020,N_11934,N_11764);
nor U13021 (N_13021,N_10957,N_11332);
nor U13022 (N_13022,N_10696,N_11412);
or U13023 (N_13023,N_10659,N_10638);
or U13024 (N_13024,N_11795,N_10582);
nand U13025 (N_13025,N_11725,N_11190);
nand U13026 (N_13026,N_11897,N_10577);
nand U13027 (N_13027,N_11707,N_11736);
nand U13028 (N_13028,N_11476,N_11499);
or U13029 (N_13029,N_11970,N_11105);
nand U13030 (N_13030,N_11721,N_10649);
or U13031 (N_13031,N_10765,N_11867);
xnor U13032 (N_13032,N_10660,N_11087);
or U13033 (N_13033,N_10636,N_11727);
or U13034 (N_13034,N_10935,N_11367);
nand U13035 (N_13035,N_11964,N_10620);
or U13036 (N_13036,N_10663,N_11843);
nand U13037 (N_13037,N_11522,N_11062);
or U13038 (N_13038,N_11349,N_10587);
or U13039 (N_13039,N_10606,N_11223);
nor U13040 (N_13040,N_11276,N_11839);
xor U13041 (N_13041,N_11023,N_10801);
and U13042 (N_13042,N_10737,N_11068);
nand U13043 (N_13043,N_11792,N_11745);
nor U13044 (N_13044,N_10903,N_10793);
or U13045 (N_13045,N_10591,N_11408);
xnor U13046 (N_13046,N_10989,N_10634);
or U13047 (N_13047,N_10842,N_11179);
and U13048 (N_13048,N_11407,N_10825);
nand U13049 (N_13049,N_11670,N_11210);
xnor U13050 (N_13050,N_11340,N_11839);
and U13051 (N_13051,N_10850,N_11156);
xor U13052 (N_13052,N_11502,N_10905);
xnor U13053 (N_13053,N_10558,N_11446);
nor U13054 (N_13054,N_11598,N_10847);
and U13055 (N_13055,N_11857,N_11098);
or U13056 (N_13056,N_11066,N_11902);
nand U13057 (N_13057,N_11747,N_10586);
nor U13058 (N_13058,N_11272,N_11383);
or U13059 (N_13059,N_11547,N_10987);
xor U13060 (N_13060,N_10989,N_11391);
nand U13061 (N_13061,N_10666,N_11963);
nor U13062 (N_13062,N_10865,N_11364);
xor U13063 (N_13063,N_10761,N_11025);
nor U13064 (N_13064,N_11484,N_10509);
and U13065 (N_13065,N_10928,N_11610);
nand U13066 (N_13066,N_11971,N_11618);
nand U13067 (N_13067,N_10772,N_11668);
nor U13068 (N_13068,N_11528,N_11290);
nor U13069 (N_13069,N_11455,N_10890);
xnor U13070 (N_13070,N_11515,N_11982);
and U13071 (N_13071,N_11263,N_11064);
xnor U13072 (N_13072,N_11888,N_11183);
xnor U13073 (N_13073,N_11440,N_10877);
and U13074 (N_13074,N_11730,N_11602);
nand U13075 (N_13075,N_11453,N_10593);
xnor U13076 (N_13076,N_11957,N_10640);
and U13077 (N_13077,N_10520,N_11641);
and U13078 (N_13078,N_10784,N_11639);
xnor U13079 (N_13079,N_10885,N_11332);
nor U13080 (N_13080,N_10792,N_10535);
or U13081 (N_13081,N_10531,N_11433);
xor U13082 (N_13082,N_11292,N_10696);
xnor U13083 (N_13083,N_11096,N_10580);
nand U13084 (N_13084,N_11502,N_11867);
nand U13085 (N_13085,N_11626,N_11998);
xor U13086 (N_13086,N_10892,N_11108);
nand U13087 (N_13087,N_11797,N_11845);
xor U13088 (N_13088,N_11625,N_11021);
and U13089 (N_13089,N_11267,N_10702);
nand U13090 (N_13090,N_10903,N_11199);
or U13091 (N_13091,N_11704,N_10936);
nor U13092 (N_13092,N_11907,N_11307);
and U13093 (N_13093,N_11741,N_11772);
and U13094 (N_13094,N_10902,N_10838);
nor U13095 (N_13095,N_11095,N_11860);
nand U13096 (N_13096,N_11896,N_10964);
or U13097 (N_13097,N_10517,N_11723);
nand U13098 (N_13098,N_11139,N_11380);
nor U13099 (N_13099,N_10527,N_10697);
xor U13100 (N_13100,N_10855,N_10873);
nor U13101 (N_13101,N_11517,N_11657);
nor U13102 (N_13102,N_10550,N_11654);
xor U13103 (N_13103,N_11296,N_11675);
nand U13104 (N_13104,N_11828,N_11222);
or U13105 (N_13105,N_11056,N_11801);
nand U13106 (N_13106,N_10867,N_11895);
or U13107 (N_13107,N_11938,N_11453);
xnor U13108 (N_13108,N_11281,N_11086);
xor U13109 (N_13109,N_11254,N_10871);
xor U13110 (N_13110,N_11519,N_10599);
xor U13111 (N_13111,N_11366,N_10671);
and U13112 (N_13112,N_10627,N_11330);
or U13113 (N_13113,N_11535,N_11089);
or U13114 (N_13114,N_11255,N_11975);
and U13115 (N_13115,N_10893,N_11067);
xnor U13116 (N_13116,N_11698,N_10765);
nor U13117 (N_13117,N_11706,N_10747);
nor U13118 (N_13118,N_10528,N_10988);
nor U13119 (N_13119,N_10912,N_11526);
and U13120 (N_13120,N_11945,N_11214);
and U13121 (N_13121,N_10621,N_11697);
nor U13122 (N_13122,N_10850,N_11139);
nand U13123 (N_13123,N_11705,N_11762);
or U13124 (N_13124,N_10633,N_11802);
or U13125 (N_13125,N_10783,N_11885);
nor U13126 (N_13126,N_11564,N_11347);
or U13127 (N_13127,N_10832,N_10625);
nor U13128 (N_13128,N_11594,N_10708);
nor U13129 (N_13129,N_10632,N_11842);
nand U13130 (N_13130,N_11211,N_10685);
nand U13131 (N_13131,N_11381,N_11838);
nor U13132 (N_13132,N_10725,N_11520);
nand U13133 (N_13133,N_10737,N_11911);
xor U13134 (N_13134,N_10692,N_11488);
and U13135 (N_13135,N_10676,N_10546);
or U13136 (N_13136,N_11457,N_10675);
nand U13137 (N_13137,N_11376,N_11714);
nand U13138 (N_13138,N_11626,N_11208);
nand U13139 (N_13139,N_11602,N_11269);
nor U13140 (N_13140,N_10843,N_11925);
and U13141 (N_13141,N_11991,N_11437);
nand U13142 (N_13142,N_11702,N_11765);
nor U13143 (N_13143,N_11798,N_11639);
nand U13144 (N_13144,N_11972,N_10636);
nand U13145 (N_13145,N_10670,N_10578);
or U13146 (N_13146,N_10537,N_11193);
nor U13147 (N_13147,N_10629,N_11110);
or U13148 (N_13148,N_11501,N_11296);
and U13149 (N_13149,N_11576,N_11176);
and U13150 (N_13150,N_11472,N_11891);
xnor U13151 (N_13151,N_11302,N_10751);
and U13152 (N_13152,N_11135,N_11997);
or U13153 (N_13153,N_11562,N_10792);
nor U13154 (N_13154,N_10796,N_10627);
xnor U13155 (N_13155,N_10915,N_11175);
nand U13156 (N_13156,N_10889,N_10539);
nor U13157 (N_13157,N_11716,N_11006);
or U13158 (N_13158,N_11918,N_10905);
nand U13159 (N_13159,N_11923,N_10955);
nand U13160 (N_13160,N_11078,N_11926);
and U13161 (N_13161,N_11957,N_10586);
xnor U13162 (N_13162,N_11755,N_11545);
nor U13163 (N_13163,N_11795,N_10853);
nand U13164 (N_13164,N_10805,N_10984);
and U13165 (N_13165,N_10535,N_10806);
nand U13166 (N_13166,N_11661,N_11989);
xnor U13167 (N_13167,N_10980,N_11777);
xnor U13168 (N_13168,N_11795,N_11726);
or U13169 (N_13169,N_11706,N_10938);
nand U13170 (N_13170,N_11807,N_10972);
xor U13171 (N_13171,N_11576,N_11267);
and U13172 (N_13172,N_10793,N_11027);
xnor U13173 (N_13173,N_11358,N_10886);
nand U13174 (N_13174,N_11092,N_11976);
and U13175 (N_13175,N_11484,N_11935);
xnor U13176 (N_13176,N_11785,N_11720);
nor U13177 (N_13177,N_10672,N_10971);
nor U13178 (N_13178,N_10848,N_11269);
nand U13179 (N_13179,N_11409,N_11417);
xor U13180 (N_13180,N_11125,N_11174);
and U13181 (N_13181,N_11701,N_11794);
or U13182 (N_13182,N_10522,N_11217);
xor U13183 (N_13183,N_11111,N_10893);
or U13184 (N_13184,N_10657,N_10575);
nor U13185 (N_13185,N_10637,N_11375);
and U13186 (N_13186,N_11610,N_11937);
nor U13187 (N_13187,N_11274,N_10977);
nor U13188 (N_13188,N_11175,N_11630);
nor U13189 (N_13189,N_10774,N_11405);
nor U13190 (N_13190,N_10707,N_10864);
nand U13191 (N_13191,N_11973,N_11295);
and U13192 (N_13192,N_11851,N_11080);
and U13193 (N_13193,N_11602,N_10535);
nand U13194 (N_13194,N_11914,N_11810);
nand U13195 (N_13195,N_10875,N_11503);
xor U13196 (N_13196,N_10705,N_10711);
nor U13197 (N_13197,N_11705,N_11757);
nor U13198 (N_13198,N_11363,N_11043);
nor U13199 (N_13199,N_11148,N_11590);
and U13200 (N_13200,N_11566,N_11704);
nor U13201 (N_13201,N_11498,N_10912);
nor U13202 (N_13202,N_11315,N_11843);
xnor U13203 (N_13203,N_11771,N_11255);
xnor U13204 (N_13204,N_11228,N_10725);
nand U13205 (N_13205,N_10881,N_10853);
nor U13206 (N_13206,N_10729,N_11327);
nor U13207 (N_13207,N_11982,N_11584);
xor U13208 (N_13208,N_10801,N_11386);
nand U13209 (N_13209,N_11744,N_11694);
or U13210 (N_13210,N_11724,N_11916);
nand U13211 (N_13211,N_11359,N_10757);
xnor U13212 (N_13212,N_11650,N_11515);
or U13213 (N_13213,N_11795,N_10952);
or U13214 (N_13214,N_11337,N_11651);
and U13215 (N_13215,N_11634,N_10816);
and U13216 (N_13216,N_11260,N_11598);
and U13217 (N_13217,N_11076,N_11535);
or U13218 (N_13218,N_11324,N_11573);
xnor U13219 (N_13219,N_11191,N_11332);
xnor U13220 (N_13220,N_11800,N_11365);
nand U13221 (N_13221,N_11706,N_11206);
nor U13222 (N_13222,N_10537,N_11094);
nor U13223 (N_13223,N_11717,N_11127);
xor U13224 (N_13224,N_11770,N_10582);
nand U13225 (N_13225,N_11585,N_11139);
and U13226 (N_13226,N_11473,N_11684);
nor U13227 (N_13227,N_11951,N_11212);
xnor U13228 (N_13228,N_11843,N_11373);
xnor U13229 (N_13229,N_11891,N_11932);
nor U13230 (N_13230,N_11505,N_11680);
and U13231 (N_13231,N_11468,N_11499);
xnor U13232 (N_13232,N_11075,N_10565);
nand U13233 (N_13233,N_11601,N_11313);
nand U13234 (N_13234,N_10724,N_11038);
xor U13235 (N_13235,N_10829,N_11381);
or U13236 (N_13236,N_11676,N_11092);
nor U13237 (N_13237,N_11081,N_11532);
or U13238 (N_13238,N_11725,N_10543);
or U13239 (N_13239,N_11204,N_11359);
nor U13240 (N_13240,N_11924,N_10941);
or U13241 (N_13241,N_11191,N_10916);
or U13242 (N_13242,N_11133,N_10879);
and U13243 (N_13243,N_11545,N_10501);
nand U13244 (N_13244,N_10998,N_10973);
nor U13245 (N_13245,N_10586,N_10938);
nor U13246 (N_13246,N_10901,N_10561);
nand U13247 (N_13247,N_10840,N_10869);
nor U13248 (N_13248,N_11134,N_11034);
xor U13249 (N_13249,N_11045,N_10883);
nand U13250 (N_13250,N_11471,N_11931);
or U13251 (N_13251,N_10613,N_10789);
nor U13252 (N_13252,N_10736,N_10572);
or U13253 (N_13253,N_11692,N_11844);
nor U13254 (N_13254,N_10983,N_11925);
nor U13255 (N_13255,N_11241,N_11313);
nand U13256 (N_13256,N_10695,N_11775);
nor U13257 (N_13257,N_10904,N_11775);
nand U13258 (N_13258,N_11767,N_11253);
nand U13259 (N_13259,N_11106,N_11528);
nand U13260 (N_13260,N_11739,N_11288);
or U13261 (N_13261,N_11124,N_11216);
or U13262 (N_13262,N_11308,N_11245);
nand U13263 (N_13263,N_11753,N_11222);
nor U13264 (N_13264,N_11502,N_10795);
or U13265 (N_13265,N_10872,N_11887);
and U13266 (N_13266,N_11633,N_11397);
nor U13267 (N_13267,N_10806,N_11209);
nand U13268 (N_13268,N_11425,N_10690);
and U13269 (N_13269,N_11200,N_11438);
xnor U13270 (N_13270,N_11373,N_11045);
xor U13271 (N_13271,N_11553,N_10742);
nor U13272 (N_13272,N_10980,N_11256);
nand U13273 (N_13273,N_11997,N_10938);
nand U13274 (N_13274,N_10872,N_11059);
nor U13275 (N_13275,N_11917,N_11685);
and U13276 (N_13276,N_11373,N_11992);
xor U13277 (N_13277,N_11834,N_11822);
nor U13278 (N_13278,N_11767,N_10745);
and U13279 (N_13279,N_11583,N_10530);
xor U13280 (N_13280,N_11147,N_10563);
nor U13281 (N_13281,N_10639,N_11102);
nand U13282 (N_13282,N_11660,N_11559);
nand U13283 (N_13283,N_11790,N_10818);
nor U13284 (N_13284,N_11869,N_11058);
nor U13285 (N_13285,N_11820,N_11129);
nor U13286 (N_13286,N_11773,N_10546);
nand U13287 (N_13287,N_11548,N_10848);
nand U13288 (N_13288,N_10818,N_11600);
and U13289 (N_13289,N_11930,N_10983);
nor U13290 (N_13290,N_10552,N_11219);
and U13291 (N_13291,N_10766,N_11875);
and U13292 (N_13292,N_11860,N_11311);
nand U13293 (N_13293,N_10597,N_11928);
nand U13294 (N_13294,N_11438,N_11407);
nor U13295 (N_13295,N_10616,N_11954);
or U13296 (N_13296,N_10549,N_10681);
or U13297 (N_13297,N_11094,N_10937);
xor U13298 (N_13298,N_11843,N_10578);
and U13299 (N_13299,N_11709,N_10953);
nand U13300 (N_13300,N_11550,N_11553);
nor U13301 (N_13301,N_11005,N_11635);
or U13302 (N_13302,N_11654,N_11117);
and U13303 (N_13303,N_10826,N_11004);
and U13304 (N_13304,N_11337,N_11161);
xnor U13305 (N_13305,N_11833,N_11551);
or U13306 (N_13306,N_11756,N_11980);
xnor U13307 (N_13307,N_11248,N_11256);
xnor U13308 (N_13308,N_11449,N_11237);
and U13309 (N_13309,N_11983,N_10667);
and U13310 (N_13310,N_11325,N_10857);
nor U13311 (N_13311,N_11003,N_11912);
or U13312 (N_13312,N_11602,N_11748);
and U13313 (N_13313,N_11913,N_10674);
and U13314 (N_13314,N_11478,N_11031);
or U13315 (N_13315,N_11204,N_11706);
nand U13316 (N_13316,N_11343,N_11801);
xor U13317 (N_13317,N_10704,N_10705);
xor U13318 (N_13318,N_11323,N_11767);
xnor U13319 (N_13319,N_10725,N_11766);
xor U13320 (N_13320,N_11782,N_10659);
or U13321 (N_13321,N_11443,N_10820);
and U13322 (N_13322,N_11083,N_11616);
xor U13323 (N_13323,N_10668,N_10658);
nand U13324 (N_13324,N_11918,N_10703);
nor U13325 (N_13325,N_11813,N_10903);
nor U13326 (N_13326,N_11903,N_11187);
or U13327 (N_13327,N_10558,N_10915);
or U13328 (N_13328,N_11188,N_11573);
nor U13329 (N_13329,N_11291,N_11987);
xor U13330 (N_13330,N_10743,N_11193);
and U13331 (N_13331,N_11462,N_11485);
or U13332 (N_13332,N_10513,N_11655);
and U13333 (N_13333,N_10673,N_11150);
nor U13334 (N_13334,N_11976,N_10875);
or U13335 (N_13335,N_11283,N_10760);
nor U13336 (N_13336,N_10646,N_11129);
nand U13337 (N_13337,N_10740,N_11214);
xor U13338 (N_13338,N_10891,N_11061);
xor U13339 (N_13339,N_11640,N_10527);
or U13340 (N_13340,N_11316,N_11781);
or U13341 (N_13341,N_11207,N_11204);
nand U13342 (N_13342,N_10885,N_11169);
or U13343 (N_13343,N_10816,N_11043);
nor U13344 (N_13344,N_11369,N_10977);
and U13345 (N_13345,N_11053,N_11350);
or U13346 (N_13346,N_10680,N_10710);
or U13347 (N_13347,N_11190,N_11617);
xnor U13348 (N_13348,N_11688,N_11915);
and U13349 (N_13349,N_11807,N_11979);
or U13350 (N_13350,N_11478,N_11849);
and U13351 (N_13351,N_11415,N_11146);
or U13352 (N_13352,N_11332,N_10558);
nand U13353 (N_13353,N_11821,N_11628);
nand U13354 (N_13354,N_10629,N_11657);
nand U13355 (N_13355,N_11504,N_11196);
and U13356 (N_13356,N_10546,N_11225);
or U13357 (N_13357,N_11227,N_11881);
nor U13358 (N_13358,N_10519,N_10802);
nand U13359 (N_13359,N_11449,N_11821);
xor U13360 (N_13360,N_11668,N_11981);
xor U13361 (N_13361,N_11923,N_11813);
nand U13362 (N_13362,N_10877,N_11844);
and U13363 (N_13363,N_10969,N_10977);
nor U13364 (N_13364,N_10902,N_10636);
or U13365 (N_13365,N_10750,N_11442);
and U13366 (N_13366,N_10586,N_10503);
or U13367 (N_13367,N_11045,N_11040);
nand U13368 (N_13368,N_10662,N_11600);
and U13369 (N_13369,N_11218,N_11134);
or U13370 (N_13370,N_11173,N_11591);
and U13371 (N_13371,N_11794,N_11987);
nand U13372 (N_13372,N_11878,N_11959);
nor U13373 (N_13373,N_11944,N_11251);
and U13374 (N_13374,N_10874,N_11472);
xor U13375 (N_13375,N_11030,N_10693);
or U13376 (N_13376,N_10693,N_10766);
nand U13377 (N_13377,N_11333,N_11200);
xor U13378 (N_13378,N_11894,N_11706);
nor U13379 (N_13379,N_11303,N_11349);
nand U13380 (N_13380,N_11470,N_11761);
nand U13381 (N_13381,N_10809,N_10758);
nand U13382 (N_13382,N_11190,N_11766);
or U13383 (N_13383,N_11675,N_10625);
or U13384 (N_13384,N_11567,N_10683);
and U13385 (N_13385,N_11037,N_11297);
nand U13386 (N_13386,N_11929,N_11962);
nand U13387 (N_13387,N_11728,N_11267);
and U13388 (N_13388,N_10524,N_10901);
or U13389 (N_13389,N_10778,N_10603);
xor U13390 (N_13390,N_10549,N_11739);
nand U13391 (N_13391,N_11707,N_10703);
or U13392 (N_13392,N_11315,N_10605);
and U13393 (N_13393,N_11548,N_11650);
xnor U13394 (N_13394,N_10664,N_11037);
xor U13395 (N_13395,N_10762,N_11637);
or U13396 (N_13396,N_10870,N_10653);
xor U13397 (N_13397,N_11049,N_11700);
or U13398 (N_13398,N_11560,N_11444);
nand U13399 (N_13399,N_11988,N_11449);
nor U13400 (N_13400,N_11267,N_11943);
and U13401 (N_13401,N_11338,N_11279);
or U13402 (N_13402,N_11990,N_11731);
nand U13403 (N_13403,N_10922,N_11542);
or U13404 (N_13404,N_11892,N_11845);
nand U13405 (N_13405,N_11934,N_11863);
xor U13406 (N_13406,N_11546,N_11116);
and U13407 (N_13407,N_11961,N_10777);
and U13408 (N_13408,N_10858,N_10711);
nand U13409 (N_13409,N_11451,N_11459);
nand U13410 (N_13410,N_11707,N_11482);
and U13411 (N_13411,N_11785,N_11450);
and U13412 (N_13412,N_11154,N_10713);
nor U13413 (N_13413,N_10783,N_11734);
nor U13414 (N_13414,N_11433,N_10972);
nor U13415 (N_13415,N_10746,N_10697);
xor U13416 (N_13416,N_10619,N_11216);
nand U13417 (N_13417,N_11250,N_10987);
or U13418 (N_13418,N_10905,N_11203);
and U13419 (N_13419,N_10681,N_11548);
or U13420 (N_13420,N_11811,N_11407);
nor U13421 (N_13421,N_11955,N_11611);
or U13422 (N_13422,N_11784,N_11360);
xor U13423 (N_13423,N_11339,N_10512);
nand U13424 (N_13424,N_10803,N_11412);
nor U13425 (N_13425,N_11314,N_10899);
nand U13426 (N_13426,N_11602,N_11876);
or U13427 (N_13427,N_11703,N_10557);
nand U13428 (N_13428,N_10989,N_11769);
or U13429 (N_13429,N_11367,N_10794);
xnor U13430 (N_13430,N_11554,N_10657);
nand U13431 (N_13431,N_10574,N_11050);
or U13432 (N_13432,N_11449,N_11673);
or U13433 (N_13433,N_11594,N_11588);
and U13434 (N_13434,N_10637,N_10904);
and U13435 (N_13435,N_11134,N_11889);
or U13436 (N_13436,N_11277,N_11059);
or U13437 (N_13437,N_11864,N_10890);
xnor U13438 (N_13438,N_11236,N_10977);
or U13439 (N_13439,N_11464,N_11806);
or U13440 (N_13440,N_11538,N_11424);
nor U13441 (N_13441,N_10874,N_11208);
and U13442 (N_13442,N_11392,N_11671);
nor U13443 (N_13443,N_11869,N_10544);
or U13444 (N_13444,N_11263,N_10871);
nand U13445 (N_13445,N_11648,N_10834);
or U13446 (N_13446,N_11071,N_11679);
and U13447 (N_13447,N_11309,N_10864);
xor U13448 (N_13448,N_11397,N_11501);
nand U13449 (N_13449,N_10590,N_11925);
nand U13450 (N_13450,N_11344,N_11974);
nand U13451 (N_13451,N_11988,N_11432);
and U13452 (N_13452,N_10628,N_11548);
or U13453 (N_13453,N_11319,N_11837);
xnor U13454 (N_13454,N_10825,N_11834);
or U13455 (N_13455,N_11150,N_11745);
or U13456 (N_13456,N_11875,N_11756);
xor U13457 (N_13457,N_11601,N_10860);
xnor U13458 (N_13458,N_11486,N_11370);
and U13459 (N_13459,N_11180,N_10548);
xor U13460 (N_13460,N_11375,N_11041);
and U13461 (N_13461,N_11552,N_11515);
or U13462 (N_13462,N_11528,N_10600);
and U13463 (N_13463,N_10515,N_11203);
and U13464 (N_13464,N_10549,N_11752);
nor U13465 (N_13465,N_11140,N_11075);
xnor U13466 (N_13466,N_11990,N_10560);
xor U13467 (N_13467,N_11070,N_11488);
and U13468 (N_13468,N_10735,N_11452);
nor U13469 (N_13469,N_10554,N_11171);
and U13470 (N_13470,N_11560,N_11745);
xnor U13471 (N_13471,N_10568,N_10598);
nor U13472 (N_13472,N_11246,N_10757);
nand U13473 (N_13473,N_11477,N_11155);
nor U13474 (N_13474,N_11489,N_11924);
nand U13475 (N_13475,N_10686,N_11412);
nand U13476 (N_13476,N_11518,N_11816);
nor U13477 (N_13477,N_11823,N_11301);
and U13478 (N_13478,N_11956,N_11545);
and U13479 (N_13479,N_11298,N_10672);
or U13480 (N_13480,N_11637,N_11053);
nand U13481 (N_13481,N_11514,N_11561);
xnor U13482 (N_13482,N_10952,N_11308);
nor U13483 (N_13483,N_11089,N_11970);
or U13484 (N_13484,N_10763,N_11835);
nor U13485 (N_13485,N_11716,N_11479);
and U13486 (N_13486,N_11715,N_11022);
xnor U13487 (N_13487,N_11483,N_10702);
and U13488 (N_13488,N_11818,N_11136);
nand U13489 (N_13489,N_10745,N_10657);
and U13490 (N_13490,N_11713,N_11855);
or U13491 (N_13491,N_11638,N_11965);
and U13492 (N_13492,N_11402,N_10525);
and U13493 (N_13493,N_11236,N_11161);
xor U13494 (N_13494,N_10629,N_10873);
xor U13495 (N_13495,N_10659,N_11819);
and U13496 (N_13496,N_10503,N_11038);
nor U13497 (N_13497,N_11440,N_10506);
nor U13498 (N_13498,N_11770,N_11948);
or U13499 (N_13499,N_11482,N_11611);
xnor U13500 (N_13500,N_13003,N_13384);
and U13501 (N_13501,N_13364,N_12665);
and U13502 (N_13502,N_12717,N_12377);
and U13503 (N_13503,N_12913,N_12146);
nor U13504 (N_13504,N_12293,N_13398);
nand U13505 (N_13505,N_12882,N_12877);
nor U13506 (N_13506,N_12100,N_12962);
nor U13507 (N_13507,N_12308,N_13028);
nor U13508 (N_13508,N_12197,N_13413);
nand U13509 (N_13509,N_13172,N_12501);
xor U13510 (N_13510,N_12283,N_13060);
and U13511 (N_13511,N_12020,N_12787);
nand U13512 (N_13512,N_12195,N_12997);
nor U13513 (N_13513,N_13263,N_12686);
nand U13514 (N_13514,N_12772,N_12475);
or U13515 (N_13515,N_12738,N_12822);
xnor U13516 (N_13516,N_12433,N_13156);
nor U13517 (N_13517,N_12984,N_12104);
or U13518 (N_13518,N_12545,N_12906);
nor U13519 (N_13519,N_13297,N_12780);
and U13520 (N_13520,N_12758,N_13025);
xnor U13521 (N_13521,N_13498,N_12769);
nand U13522 (N_13522,N_12472,N_12103);
and U13523 (N_13523,N_12762,N_13442);
or U13524 (N_13524,N_12929,N_12641);
nor U13525 (N_13525,N_12234,N_12672);
and U13526 (N_13526,N_13270,N_13248);
or U13527 (N_13527,N_13479,N_13457);
xor U13528 (N_13528,N_12843,N_13010);
xnor U13529 (N_13529,N_12830,N_13326);
nor U13530 (N_13530,N_13088,N_12141);
or U13531 (N_13531,N_12371,N_13021);
or U13532 (N_13532,N_12278,N_12809);
xor U13533 (N_13533,N_12098,N_12801);
nand U13534 (N_13534,N_12645,N_13085);
xor U13535 (N_13535,N_12420,N_12647);
xor U13536 (N_13536,N_13487,N_12824);
or U13537 (N_13537,N_12189,N_13080);
nor U13538 (N_13538,N_13011,N_13052);
xnor U13539 (N_13539,N_12477,N_13046);
nand U13540 (N_13540,N_12664,N_13233);
xnor U13541 (N_13541,N_13460,N_12749);
xor U13542 (N_13542,N_12237,N_12701);
nand U13543 (N_13543,N_13024,N_12423);
or U13544 (N_13544,N_13219,N_13311);
nor U13545 (N_13545,N_12200,N_13063);
xor U13546 (N_13546,N_12855,N_12192);
nand U13547 (N_13547,N_13295,N_12960);
nor U13548 (N_13548,N_12188,N_12368);
nand U13549 (N_13549,N_12306,N_13342);
or U13550 (N_13550,N_12562,N_13375);
and U13551 (N_13551,N_12771,N_12430);
nand U13552 (N_13552,N_12727,N_13058);
or U13553 (N_13553,N_13212,N_12886);
nand U13554 (N_13554,N_13417,N_12417);
and U13555 (N_13555,N_12298,N_12059);
or U13556 (N_13556,N_13471,N_13069);
or U13557 (N_13557,N_12112,N_12601);
and U13558 (N_13558,N_13045,N_12279);
nor U13559 (N_13559,N_12421,N_13374);
or U13560 (N_13560,N_12041,N_12054);
nand U13561 (N_13561,N_12217,N_12144);
or U13562 (N_13562,N_12643,N_12186);
or U13563 (N_13563,N_12201,N_12770);
or U13564 (N_13564,N_13369,N_13341);
or U13565 (N_13565,N_13053,N_12367);
nor U13566 (N_13566,N_12205,N_12966);
xor U13567 (N_13567,N_13307,N_12702);
or U13568 (N_13568,N_12479,N_12937);
nand U13569 (N_13569,N_12779,N_13397);
nor U13570 (N_13570,N_13102,N_13113);
xor U13571 (N_13571,N_12334,N_12943);
nand U13572 (N_13572,N_12783,N_12190);
or U13573 (N_13573,N_12220,N_13409);
or U13574 (N_13574,N_12628,N_12925);
or U13575 (N_13575,N_13392,N_12303);
or U13576 (N_13576,N_12097,N_13218);
and U13577 (N_13577,N_12276,N_12044);
nor U13578 (N_13578,N_12030,N_12229);
xor U13579 (N_13579,N_12038,N_12720);
nor U13580 (N_13580,N_12951,N_12765);
xor U13581 (N_13581,N_12734,N_12244);
nor U13582 (N_13582,N_12979,N_13288);
xor U13583 (N_13583,N_12255,N_12135);
or U13584 (N_13584,N_13244,N_13198);
and U13585 (N_13585,N_13148,N_13388);
or U13586 (N_13586,N_12795,N_13267);
xor U13587 (N_13587,N_12386,N_12311);
or U13588 (N_13588,N_12267,N_13072);
and U13589 (N_13589,N_12662,N_13387);
or U13590 (N_13590,N_12378,N_12581);
or U13591 (N_13591,N_12870,N_13395);
or U13592 (N_13592,N_12360,N_13211);
nor U13593 (N_13593,N_13182,N_13140);
or U13594 (N_13594,N_12549,N_12998);
nand U13595 (N_13595,N_12976,N_12441);
or U13596 (N_13596,N_12968,N_12494);
nand U13597 (N_13597,N_12031,N_13178);
and U13598 (N_13598,N_12039,N_12499);
and U13599 (N_13599,N_12495,N_12698);
nand U13600 (N_13600,N_13147,N_13343);
xor U13601 (N_13601,N_12596,N_12766);
xnor U13602 (N_13602,N_12397,N_12573);
nor U13603 (N_13603,N_12070,N_12989);
or U13604 (N_13604,N_12275,N_12470);
and U13605 (N_13605,N_12793,N_12113);
or U13606 (N_13606,N_13418,N_12558);
and U13607 (N_13607,N_12816,N_13097);
and U13608 (N_13608,N_13016,N_12362);
or U13609 (N_13609,N_13189,N_12695);
xor U13610 (N_13610,N_12151,N_13377);
xor U13611 (N_13611,N_12357,N_12295);
xor U13612 (N_13612,N_12159,N_12706);
nand U13613 (N_13613,N_12277,N_12489);
nand U13614 (N_13614,N_12388,N_12831);
nor U13615 (N_13615,N_12256,N_12033);
nor U13616 (N_13616,N_13253,N_13474);
xor U13617 (N_13617,N_12332,N_12867);
xor U13618 (N_13618,N_12061,N_12453);
xor U13619 (N_13619,N_12956,N_12704);
nand U13620 (N_13620,N_12076,N_13443);
or U13621 (N_13621,N_12443,N_12316);
nor U13622 (N_13622,N_13290,N_12953);
xor U13623 (N_13623,N_12000,N_13365);
nor U13624 (N_13624,N_13208,N_12243);
or U13625 (N_13625,N_12526,N_12163);
nand U13626 (N_13626,N_12811,N_12437);
nand U13627 (N_13627,N_12454,N_13345);
and U13628 (N_13628,N_13152,N_12651);
xnor U13629 (N_13629,N_12580,N_12162);
nor U13630 (N_13630,N_13252,N_13020);
and U13631 (N_13631,N_12525,N_12292);
xnor U13632 (N_13632,N_13214,N_13420);
or U13633 (N_13633,N_12637,N_13389);
nand U13634 (N_13634,N_12546,N_13122);
xor U13635 (N_13635,N_13023,N_12006);
and U13636 (N_13636,N_13470,N_13157);
nand U13637 (N_13637,N_13273,N_12012);
and U13638 (N_13638,N_12358,N_12516);
or U13639 (N_13639,N_12755,N_12253);
or U13640 (N_13640,N_12920,N_12908);
or U13641 (N_13641,N_12524,N_12819);
and U13642 (N_13642,N_13476,N_12015);
and U13643 (N_13643,N_13117,N_13034);
xnor U13644 (N_13644,N_12222,N_12642);
nand U13645 (N_13645,N_12861,N_12062);
or U13646 (N_13646,N_12575,N_12345);
nand U13647 (N_13647,N_12291,N_12782);
nand U13648 (N_13648,N_12744,N_12668);
xnor U13649 (N_13649,N_13256,N_12846);
nor U13650 (N_13650,N_13031,N_12406);
or U13651 (N_13651,N_13475,N_12338);
and U13652 (N_13652,N_12586,N_12235);
xor U13653 (N_13653,N_12482,N_12434);
or U13654 (N_13654,N_13049,N_12412);
xor U13655 (N_13655,N_12804,N_12119);
and U13656 (N_13656,N_12851,N_12810);
xor U13657 (N_13657,N_13142,N_12569);
nand U13658 (N_13658,N_12607,N_12604);
xor U13659 (N_13659,N_12543,N_12284);
or U13660 (N_13660,N_12595,N_12307);
and U13661 (N_13661,N_12792,N_12413);
nor U13662 (N_13662,N_13136,N_13126);
and U13663 (N_13663,N_12093,N_13357);
nand U13664 (N_13664,N_13184,N_13416);
nand U13665 (N_13665,N_12722,N_12899);
nand U13666 (N_13666,N_12796,N_12981);
nand U13667 (N_13667,N_12785,N_12414);
xnor U13668 (N_13668,N_12258,N_13149);
nand U13669 (N_13669,N_13170,N_12947);
xor U13670 (N_13670,N_12603,N_12468);
nand U13671 (N_13671,N_12590,N_12829);
and U13672 (N_13672,N_13481,N_12600);
nand U13673 (N_13673,N_13463,N_13455);
xnor U13674 (N_13674,N_13105,N_13332);
nand U13675 (N_13675,N_12820,N_12964);
nand U13676 (N_13676,N_13322,N_12376);
and U13677 (N_13677,N_12393,N_13019);
nor U13678 (N_13678,N_12732,N_13177);
and U13679 (N_13679,N_12660,N_12449);
or U13680 (N_13680,N_13445,N_12252);
nand U13681 (N_13681,N_13245,N_12321);
nand U13682 (N_13682,N_12339,N_12124);
and U13683 (N_13683,N_13161,N_12812);
xnor U13684 (N_13684,N_12418,N_12958);
nand U13685 (N_13685,N_12954,N_12272);
xor U13686 (N_13686,N_13108,N_13123);
or U13687 (N_13687,N_12176,N_12024);
xor U13688 (N_13688,N_12193,N_12398);
nor U13689 (N_13689,N_12950,N_13289);
nand U13690 (N_13690,N_12260,N_13279);
xor U13691 (N_13691,N_12289,N_13319);
nand U13692 (N_13692,N_12326,N_12138);
xor U13693 (N_13693,N_12930,N_12225);
xnor U13694 (N_13694,N_13220,N_12152);
or U13695 (N_13695,N_12860,N_12745);
and U13696 (N_13696,N_12659,N_12207);
or U13697 (N_13697,N_12158,N_13489);
nand U13698 (N_13698,N_12040,N_12356);
or U13699 (N_13699,N_12347,N_12876);
nand U13700 (N_13700,N_13465,N_12832);
nand U13701 (N_13701,N_13380,N_13201);
and U13702 (N_13702,N_12444,N_13124);
nor U13703 (N_13703,N_12194,N_12187);
nand U13704 (N_13704,N_12791,N_13217);
or U13705 (N_13705,N_12409,N_13317);
and U13706 (N_13706,N_13160,N_13026);
nand U13707 (N_13707,N_12707,N_13158);
nor U13708 (N_13708,N_13431,N_12459);
and U13709 (N_13709,N_13154,N_12667);
and U13710 (N_13710,N_13368,N_13180);
and U13711 (N_13711,N_12153,N_13404);
or U13712 (N_13712,N_12521,N_13411);
or U13713 (N_13713,N_12233,N_12463);
nand U13714 (N_13714,N_12730,N_12605);
nor U13715 (N_13715,N_12161,N_12602);
and U13716 (N_13716,N_12327,N_12130);
or U13717 (N_13717,N_12508,N_12952);
or U13718 (N_13718,N_12369,N_12895);
nor U13719 (N_13719,N_12705,N_12648);
and U13720 (N_13720,N_13286,N_12328);
xnor U13721 (N_13721,N_13354,N_13268);
nor U13722 (N_13722,N_12089,N_12673);
and U13723 (N_13723,N_12560,N_12210);
nand U13724 (N_13724,N_12513,N_12268);
or U13725 (N_13725,N_12676,N_12317);
xnor U13726 (N_13726,N_13153,N_12211);
nand U13727 (N_13727,N_12383,N_12561);
nand U13728 (N_13728,N_12416,N_12985);
and U13729 (N_13729,N_13310,N_13283);
nand U13730 (N_13730,N_12788,N_12827);
or U13731 (N_13731,N_12106,N_13190);
nor U13732 (N_13732,N_12552,N_13036);
xnor U13733 (N_13733,N_12864,N_12419);
xor U13734 (N_13734,N_12689,N_13287);
or U13735 (N_13735,N_12498,N_13433);
or U13736 (N_13736,N_12946,N_12068);
or U13737 (N_13737,N_12131,N_13439);
or U13738 (N_13738,N_12885,N_12528);
or U13739 (N_13739,N_13008,N_12105);
or U13740 (N_13740,N_12122,N_12630);
and U13741 (N_13741,N_12900,N_12938);
nand U13742 (N_13742,N_13095,N_12715);
nand U13743 (N_13743,N_13356,N_12879);
nand U13744 (N_13744,N_12294,N_13089);
and U13745 (N_13745,N_12052,N_13456);
nor U13746 (N_13746,N_12612,N_13394);
and U13747 (N_13747,N_12426,N_12786);
nand U13748 (N_13748,N_12752,N_13259);
xor U13749 (N_13749,N_12476,N_12904);
or U13750 (N_13750,N_13472,N_13367);
xnor U13751 (N_13751,N_12107,N_13043);
nand U13752 (N_13752,N_12571,N_12018);
and U13753 (N_13753,N_12535,N_12842);
xor U13754 (N_13754,N_12522,N_12675);
and U13755 (N_13755,N_12799,N_12335);
nor U13756 (N_13756,N_12891,N_12688);
xnor U13757 (N_13757,N_12593,N_12523);
nand U13758 (N_13758,N_12139,N_12736);
and U13759 (N_13759,N_13320,N_13340);
or U13760 (N_13760,N_12324,N_13206);
nand U13761 (N_13761,N_12578,N_12036);
xnor U13762 (N_13762,N_12491,N_12646);
xnor U13763 (N_13763,N_12723,N_12432);
xnor U13764 (N_13764,N_13249,N_13141);
nor U13765 (N_13765,N_12540,N_12965);
or U13766 (N_13766,N_12719,N_12505);
nand U13767 (N_13767,N_12023,N_13005);
nor U13768 (N_13768,N_12574,N_13174);
nand U13769 (N_13769,N_13099,N_12315);
nand U13770 (N_13770,N_13318,N_12261);
or U13771 (N_13771,N_12503,N_12692);
xor U13772 (N_13772,N_13001,N_12032);
nor U13773 (N_13773,N_13315,N_13084);
and U13774 (N_13774,N_13347,N_12741);
nor U13775 (N_13775,N_12905,N_12974);
and U13776 (N_13776,N_12007,N_12082);
xnor U13777 (N_13777,N_12086,N_12019);
nand U13778 (N_13778,N_12889,N_12557);
nand U13779 (N_13779,N_12435,N_13469);
nor U13780 (N_13780,N_12663,N_12504);
xor U13781 (N_13781,N_13071,N_13261);
or U13782 (N_13782,N_12721,N_12208);
and U13783 (N_13783,N_12175,N_12057);
xnor U13784 (N_13784,N_13302,N_13027);
nor U13785 (N_13785,N_12839,N_12797);
or U13786 (N_13786,N_13401,N_12457);
nand U13787 (N_13787,N_13371,N_13109);
or U13788 (N_13788,N_13379,N_12478);
or U13789 (N_13789,N_12712,N_12892);
nor U13790 (N_13790,N_12325,N_12680);
xor U13791 (N_13791,N_13304,N_13223);
and U13792 (N_13792,N_13065,N_12548);
or U13793 (N_13793,N_12168,N_12365);
nand U13794 (N_13794,N_12221,N_12507);
or U13795 (N_13795,N_12613,N_13306);
or U13796 (N_13796,N_12322,N_12568);
and U13797 (N_13797,N_13130,N_12149);
nand U13798 (N_13798,N_12655,N_12066);
xor U13799 (N_13799,N_13265,N_12399);
and U13800 (N_13800,N_13493,N_13004);
or U13801 (N_13801,N_13482,N_13251);
nand U13802 (N_13802,N_13055,N_13144);
or U13803 (N_13803,N_13056,N_13477);
nand U13804 (N_13804,N_12699,N_12865);
and U13805 (N_13805,N_12037,N_12579);
xnor U13806 (N_13806,N_12681,N_12658);
and U13807 (N_13807,N_13258,N_12703);
xor U13808 (N_13808,N_12653,N_13281);
nor U13809 (N_13809,N_12051,N_13224);
or U13810 (N_13810,N_13014,N_13271);
nand U13811 (N_13811,N_12509,N_13323);
xor U13812 (N_13812,N_12354,N_13274);
xor U13813 (N_13813,N_12074,N_12431);
nor U13814 (N_13814,N_12775,N_12942);
nor U13815 (N_13815,N_13061,N_13074);
nor U13816 (N_13816,N_13007,N_12085);
and U13817 (N_13817,N_12405,N_12374);
xnor U13818 (N_13818,N_13429,N_12777);
nand U13819 (N_13819,N_12693,N_13419);
and U13820 (N_13820,N_12169,N_13305);
nor U13821 (N_13821,N_12348,N_12577);
nor U13822 (N_13822,N_12994,N_12746);
nor U13823 (N_13823,N_12228,N_13185);
xor U13824 (N_13824,N_12259,N_13484);
xor U13825 (N_13825,N_13137,N_13264);
nor U13826 (N_13826,N_12333,N_13353);
nand U13827 (N_13827,N_12296,N_13490);
and U13828 (N_13828,N_12921,N_12778);
and U13829 (N_13829,N_13066,N_12003);
and U13830 (N_13830,N_12697,N_12618);
nand U13831 (N_13831,N_13446,N_12133);
or U13832 (N_13832,N_12203,N_12683);
nand U13833 (N_13833,N_12456,N_13448);
and U13834 (N_13834,N_13114,N_13164);
xor U13835 (N_13835,N_12366,N_13018);
xor U13836 (N_13836,N_12922,N_12747);
xnor U13837 (N_13837,N_12875,N_12972);
xor U13838 (N_13838,N_13090,N_12271);
nand U13839 (N_13839,N_12868,N_13216);
nor U13840 (N_13840,N_12013,N_13068);
or U13841 (N_13841,N_12874,N_12530);
nand U13842 (N_13842,N_12671,N_13346);
or U13843 (N_13843,N_12171,N_13497);
xor U13844 (N_13844,N_12670,N_12733);
nand U13845 (N_13845,N_12091,N_13193);
or U13846 (N_13846,N_12533,N_13146);
nor U13847 (N_13847,N_12464,N_12485);
nand U13848 (N_13848,N_13403,N_12323);
xnor U13849 (N_13849,N_12532,N_13405);
and U13850 (N_13850,N_13111,N_12969);
or U13851 (N_13851,N_13150,N_12599);
or U13852 (N_13852,N_12402,N_13225);
and U13853 (N_13853,N_12845,N_12781);
nor U13854 (N_13854,N_12666,N_13250);
xnor U13855 (N_13855,N_13076,N_12735);
nand U13856 (N_13856,N_12725,N_13232);
and U13857 (N_13857,N_12807,N_12551);
xor U13858 (N_13858,N_13255,N_13228);
and U13859 (N_13859,N_13143,N_13187);
and U13860 (N_13860,N_13030,N_13352);
or U13861 (N_13861,N_13293,N_12948);
nand U13862 (N_13862,N_13086,N_13183);
and U13863 (N_13863,N_12240,N_13314);
nand U13864 (N_13864,N_13370,N_13176);
nand U13865 (N_13865,N_12336,N_13402);
and U13866 (N_13866,N_12320,N_12045);
or U13867 (N_13867,N_12390,N_12587);
nand U13868 (N_13868,N_12455,N_12896);
nand U13869 (N_13869,N_12841,N_12739);
or U13870 (N_13870,N_12635,N_13213);
nand U13871 (N_13871,N_12588,N_12751);
xnor U13872 (N_13872,N_12955,N_12639);
nor U13873 (N_13873,N_12330,N_13412);
and U13874 (N_13874,N_13033,N_13070);
nand U13875 (N_13875,N_13309,N_13231);
or U13876 (N_13876,N_13427,N_12917);
or U13877 (N_13877,N_12273,N_13096);
or U13878 (N_13878,N_12346,N_12465);
xor U13879 (N_13879,N_12134,N_13362);
or U13880 (N_13880,N_12123,N_12626);
nor U13881 (N_13881,N_13091,N_12199);
nand U13882 (N_13882,N_12800,N_12887);
or U13883 (N_13883,N_13390,N_12392);
xor U13884 (N_13884,N_13236,N_13499);
xnor U13885 (N_13885,N_12999,N_12056);
xnor U13886 (N_13886,N_13344,N_12314);
nor U13887 (N_13887,N_12511,N_13151);
nand U13888 (N_13888,N_12411,N_12679);
nand U13889 (N_13889,N_13054,N_12591);
xor U13890 (N_13890,N_12669,N_12083);
xor U13891 (N_13891,N_12170,N_12617);
and U13892 (N_13892,N_13348,N_13135);
or U13893 (N_13893,N_12844,N_12894);
xnor U13894 (N_13894,N_13366,N_13494);
nand U13895 (N_13895,N_13194,N_13222);
and U13896 (N_13896,N_12983,N_13040);
or U13897 (N_13897,N_12026,N_12309);
and U13898 (N_13898,N_12961,N_13107);
or U13899 (N_13899,N_13278,N_12394);
nor U13900 (N_13900,N_13022,N_12803);
nor U13901 (N_13901,N_13234,N_13204);
nor U13902 (N_13902,N_12154,N_12143);
nand U13903 (N_13903,N_12118,N_12035);
nor U13904 (N_13904,N_13078,N_13128);
or U13905 (N_13905,N_12515,N_13284);
or U13906 (N_13906,N_12991,N_12784);
or U13907 (N_13907,N_12262,N_12183);
nor U13908 (N_13908,N_13257,N_13408);
nand U13909 (N_13909,N_13262,N_12564);
and U13910 (N_13910,N_13386,N_12767);
nor U13911 (N_13911,N_12427,N_12075);
nand U13912 (N_13912,N_12461,N_13254);
nand U13913 (N_13913,N_13075,N_12077);
nor U13914 (N_13914,N_12901,N_13452);
and U13915 (N_13915,N_13199,N_12125);
xnor U13916 (N_13916,N_12517,N_12849);
or U13917 (N_13917,N_12471,N_12836);
and U13918 (N_13918,N_12400,N_13067);
or U13919 (N_13919,N_12854,N_13424);
nor U13920 (N_13920,N_12108,N_12047);
or U13921 (N_13921,N_12179,N_12084);
nand U13922 (N_13922,N_13202,N_13064);
nand U13923 (N_13923,N_12565,N_12361);
and U13924 (N_13924,N_12167,N_12387);
nor U13925 (N_13925,N_12483,N_12970);
or U13926 (N_13926,N_12069,N_12542);
or U13927 (N_13927,N_12389,N_13167);
or U13928 (N_13928,N_13324,N_12848);
xnor U13929 (N_13929,N_12490,N_13426);
nor U13930 (N_13930,N_12835,N_13294);
nand U13931 (N_13931,N_12288,N_12608);
xor U13932 (N_13932,N_13101,N_12282);
or U13933 (N_13933,N_12251,N_13327);
or U13934 (N_13934,N_12754,N_13467);
nand U13935 (N_13935,N_12949,N_13132);
xor U13936 (N_13936,N_12518,N_13051);
nor U13937 (N_13937,N_13393,N_12213);
xnor U13938 (N_13938,N_12709,N_12934);
and U13939 (N_13939,N_12928,N_12563);
nor U13940 (N_13940,N_13119,N_13079);
xor U13941 (N_13941,N_12761,N_13331);
or U13942 (N_13942,N_12813,N_12614);
and U13943 (N_13943,N_13459,N_12227);
xor U13944 (N_13944,N_12241,N_12724);
nand U13945 (N_13945,N_13300,N_12806);
xor U13946 (N_13946,N_12014,N_12164);
and U13947 (N_13947,N_12174,N_12768);
xor U13948 (N_13948,N_12594,N_12980);
and U13949 (N_13949,N_12497,N_12931);
or U13950 (N_13950,N_12945,N_12440);
xor U13951 (N_13951,N_13350,N_12001);
nand U13952 (N_13952,N_12910,N_13104);
nand U13953 (N_13953,N_12756,N_12514);
or U13954 (N_13954,N_12691,N_12678);
nand U13955 (N_13955,N_12919,N_12500);
nand U13956 (N_13956,N_13308,N_12340);
nor U13957 (N_13957,N_12857,N_12297);
xnor U13958 (N_13958,N_13441,N_12396);
xor U13959 (N_13959,N_13243,N_12988);
nand U13960 (N_13960,N_13133,N_12407);
and U13961 (N_13961,N_12450,N_12902);
nand U13962 (N_13962,N_12353,N_12238);
nor U13963 (N_13963,N_12342,N_12993);
or U13964 (N_13964,N_13428,N_12852);
nand U13965 (N_13965,N_13292,N_12088);
nor U13966 (N_13966,N_13335,N_12971);
xor U13967 (N_13967,N_13449,N_12274);
or U13968 (N_13968,N_12246,N_12058);
nor U13969 (N_13969,N_12621,N_13351);
or U13970 (N_13970,N_12833,N_12422);
nand U13971 (N_13971,N_12247,N_12519);
nand U13972 (N_13972,N_13235,N_12764);
nor U13973 (N_13973,N_13103,N_12429);
nand U13974 (N_13974,N_12110,N_13165);
or U13975 (N_13975,N_12257,N_13480);
nand U13976 (N_13976,N_12537,N_13129);
nor U13977 (N_13977,N_13435,N_12156);
nor U13978 (N_13978,N_12230,N_12381);
nor U13979 (N_13979,N_13047,N_13399);
and U13980 (N_13980,N_12496,N_12239);
nand U13981 (N_13981,N_12684,N_12428);
or U13982 (N_13982,N_12281,N_12616);
nand U13983 (N_13983,N_12567,N_13376);
and U13984 (N_13984,N_12566,N_12099);
nor U13985 (N_13985,N_13296,N_12534);
nor U13986 (N_13986,N_12863,N_12140);
nor U13987 (N_13987,N_12584,N_12615);
nor U13988 (N_13988,N_12620,N_12790);
xnor U13989 (N_13989,N_13423,N_12926);
nor U13990 (N_13990,N_13196,N_12555);
nand U13991 (N_13991,N_12656,N_12029);
or U13992 (N_13992,N_13159,N_12351);
and U13993 (N_13993,N_12576,N_13203);
nor U13994 (N_13994,N_13112,N_13221);
xor U13995 (N_13995,N_13358,N_12448);
nor U13996 (N_13996,N_12128,N_13451);
nand U13997 (N_13997,N_12978,N_12990);
nor U13998 (N_13998,N_12763,N_12250);
or U13999 (N_13999,N_12529,N_13163);
and U14000 (N_14000,N_13266,N_13175);
or U14001 (N_14001,N_12939,N_13215);
nand U14002 (N_14002,N_13121,N_12583);
or U14003 (N_14003,N_12034,N_12606);
xnor U14004 (N_14004,N_12331,N_12280);
nand U14005 (N_14005,N_13138,N_12743);
and U14006 (N_14006,N_12017,N_12789);
nor U14007 (N_14007,N_12714,N_12137);
nor U14008 (N_14008,N_12060,N_13385);
or U14009 (N_14009,N_12359,N_12710);
nand U14010 (N_14010,N_13316,N_12927);
nor U14011 (N_14011,N_12285,N_13237);
nand U14012 (N_14012,N_12467,N_12126);
nor U14013 (N_14013,N_12963,N_12313);
xor U14014 (N_14014,N_13000,N_12299);
or U14015 (N_14015,N_12090,N_12087);
nand U14016 (N_14016,N_12157,N_12236);
xor U14017 (N_14017,N_12264,N_12729);
xnor U14018 (N_14018,N_12166,N_13087);
or U14019 (N_14019,N_13230,N_12975);
nand U14020 (N_14020,N_13372,N_12198);
and U14021 (N_14021,N_12403,N_13125);
nor U14022 (N_14022,N_12700,N_12242);
nand U14023 (N_14023,N_12941,N_13410);
xnor U14024 (N_14024,N_13328,N_13062);
and U14025 (N_14025,N_12484,N_12650);
xor U14026 (N_14026,N_12932,N_12716);
or U14027 (N_14027,N_13081,N_12341);
and U14028 (N_14028,N_12410,N_12881);
xor U14029 (N_14029,N_12798,N_12597);
and U14030 (N_14030,N_12794,N_12363);
xor U14031 (N_14031,N_13313,N_13325);
xor U14032 (N_14032,N_12249,N_12506);
nand U14033 (N_14033,N_13241,N_12310);
nand U14034 (N_14034,N_12973,N_12638);
or U14035 (N_14035,N_12872,N_12748);
nor U14036 (N_14036,N_12592,N_12224);
nor U14037 (N_14037,N_12654,N_13162);
nand U14038 (N_14038,N_12266,N_13029);
nor U14039 (N_14039,N_13171,N_12996);
nor U14040 (N_14040,N_12726,N_13363);
or U14041 (N_14041,N_13422,N_12028);
and U14042 (N_14042,N_13032,N_12212);
or U14043 (N_14043,N_13116,N_12053);
and U14044 (N_14044,N_12344,N_13077);
xnor U14045 (N_14045,N_12048,N_12185);
xor U14046 (N_14046,N_12269,N_13276);
nor U14047 (N_14047,N_12102,N_12907);
or U14048 (N_14048,N_12916,N_12817);
or U14049 (N_14049,N_13436,N_12384);
or U14050 (N_14050,N_12550,N_12880);
or U14051 (N_14051,N_13042,N_12218);
and U14052 (N_14052,N_13118,N_13006);
or U14053 (N_14053,N_12094,N_13382);
or U14054 (N_14054,N_12395,N_12531);
and U14055 (N_14055,N_13491,N_12116);
or U14056 (N_14056,N_13106,N_13181);
nor U14057 (N_14057,N_12987,N_12536);
nor U14058 (N_14058,N_13450,N_12226);
xor U14059 (N_14059,N_12553,N_12178);
or U14060 (N_14060,N_12632,N_13333);
xnor U14061 (N_14061,N_12967,N_12375);
and U14062 (N_14062,N_12101,N_13039);
nor U14063 (N_14063,N_13083,N_12847);
or U14064 (N_14064,N_12914,N_12424);
and U14065 (N_14065,N_12888,N_13186);
and U14066 (N_14066,N_12859,N_12918);
nand U14067 (N_14067,N_12011,N_13155);
nor U14068 (N_14068,N_12862,N_12370);
nand U14069 (N_14069,N_12502,N_12512);
nand U14070 (N_14070,N_12206,N_12776);
and U14071 (N_14071,N_12823,N_12120);
nand U14072 (N_14072,N_12300,N_12570);
and U14073 (N_14073,N_12674,N_13173);
nand U14074 (N_14074,N_12290,N_12415);
nand U14075 (N_14075,N_12995,N_13462);
xnor U14076 (N_14076,N_12538,N_12598);
xnor U14077 (N_14077,N_12147,N_12286);
xor U14078 (N_14078,N_13437,N_13396);
or U14079 (N_14079,N_12223,N_13229);
nand U14080 (N_14080,N_12073,N_12840);
nor U14081 (N_14081,N_13330,N_12451);
or U14082 (N_14082,N_12191,N_12898);
xor U14083 (N_14083,N_13478,N_13337);
and U14084 (N_14084,N_12959,N_12231);
nor U14085 (N_14085,N_12355,N_13192);
nand U14086 (N_14086,N_13495,N_12046);
xor U14087 (N_14087,N_13269,N_12682);
xor U14088 (N_14088,N_12111,N_12148);
and U14089 (N_14089,N_13383,N_12095);
nor U14090 (N_14090,N_13239,N_13207);
nand U14091 (N_14091,N_12760,N_12629);
nand U14092 (N_14092,N_12890,N_12155);
and U14093 (N_14093,N_12677,N_12263);
xor U14094 (N_14094,N_12821,N_12380);
and U14095 (N_14095,N_13406,N_12458);
xnor U14096 (N_14096,N_12856,N_12711);
nor U14097 (N_14097,N_13098,N_12544);
nand U14098 (N_14098,N_12740,N_12866);
nor U14099 (N_14099,N_12957,N_12633);
nand U14100 (N_14100,N_12172,N_13421);
nor U14101 (N_14101,N_12923,N_12869);
or U14102 (N_14102,N_12287,N_12109);
or U14103 (N_14103,N_12759,N_13355);
nand U14104 (N_14104,N_12127,N_12850);
nand U14105 (N_14105,N_12644,N_13009);
and U14106 (N_14106,N_12488,N_12805);
and U14107 (N_14107,N_13359,N_13169);
or U14108 (N_14108,N_13247,N_12343);
nand U14109 (N_14109,N_12142,N_13440);
nor U14110 (N_14110,N_12265,N_12622);
nor U14111 (N_14111,N_12634,N_12072);
and U14112 (N_14112,N_12025,N_12559);
nor U14113 (N_14113,N_13246,N_13301);
and U14114 (N_14114,N_12005,N_12652);
and U14115 (N_14115,N_12903,N_13110);
and U14116 (N_14116,N_12232,N_13361);
or U14117 (N_14117,N_13461,N_13483);
and U14118 (N_14118,N_12802,N_12893);
nand U14119 (N_14119,N_13059,N_12373);
xnor U14120 (N_14120,N_13464,N_12619);
nand U14121 (N_14121,N_13226,N_12572);
or U14122 (N_14122,N_13092,N_12818);
nor U14123 (N_14123,N_12318,N_12911);
xor U14124 (N_14124,N_13329,N_12474);
nor U14125 (N_14125,N_12442,N_13093);
and U14126 (N_14126,N_12742,N_12204);
and U14127 (N_14127,N_12897,N_13468);
or U14128 (N_14128,N_12067,N_12556);
nand U14129 (N_14129,N_13280,N_12636);
and U14130 (N_14130,N_12912,N_13127);
nand U14131 (N_14131,N_13205,N_12096);
xnor U14132 (N_14132,N_13275,N_12021);
xor U14133 (N_14133,N_12944,N_12352);
xnor U14134 (N_14134,N_12049,N_13299);
and U14135 (N_14135,N_12080,N_12115);
nand U14136 (N_14136,N_12462,N_12436);
nand U14137 (N_14137,N_13488,N_12337);
nor U14138 (N_14138,N_12270,N_12022);
xor U14139 (N_14139,N_12828,N_12129);
xnor U14140 (N_14140,N_13458,N_13002);
and U14141 (N_14141,N_12438,N_12349);
nand U14142 (N_14142,N_12002,N_13038);
nand U14143 (N_14143,N_12486,N_13139);
or U14144 (N_14144,N_12182,N_13486);
xnor U14145 (N_14145,N_12042,N_12473);
and U14146 (N_14146,N_13338,N_12214);
and U14147 (N_14147,N_12871,N_12982);
xnor U14148 (N_14148,N_12624,N_13188);
nand U14149 (N_14149,N_12731,N_12016);
xor U14150 (N_14150,N_13179,N_12582);
nor U14151 (N_14151,N_12547,N_13227);
or U14152 (N_14152,N_13291,N_12184);
or U14153 (N_14153,N_12181,N_12245);
nand U14154 (N_14154,N_12145,N_12657);
nor U14155 (N_14155,N_12936,N_13240);
nand U14156 (N_14156,N_13438,N_12884);
xor U14157 (N_14157,N_13013,N_12004);
nand U14158 (N_14158,N_13191,N_12510);
nor U14159 (N_14159,N_12858,N_12649);
nand U14160 (N_14160,N_12132,N_13378);
or U14161 (N_14161,N_12302,N_12425);
and U14162 (N_14162,N_12625,N_12728);
xor U14163 (N_14163,N_12718,N_13131);
xor U14164 (N_14164,N_13432,N_12696);
nand U14165 (N_14165,N_13037,N_12690);
nand U14166 (N_14166,N_12064,N_12364);
or U14167 (N_14167,N_13360,N_12554);
or U14168 (N_14168,N_13415,N_12750);
nor U14169 (N_14169,N_12623,N_12254);
nand U14170 (N_14170,N_12439,N_12445);
xnor U14171 (N_14171,N_13017,N_12446);
nor U14172 (N_14172,N_12611,N_13082);
or U14173 (N_14173,N_13492,N_13434);
nand U14174 (N_14174,N_13303,N_12010);
xnor U14175 (N_14175,N_13485,N_12055);
xnor U14176 (N_14176,N_12924,N_13200);
or U14177 (N_14177,N_13447,N_12493);
or U14178 (N_14178,N_12304,N_12935);
nor U14179 (N_14179,N_12492,N_13115);
nor U14180 (N_14180,N_12992,N_13195);
or U14181 (N_14181,N_12382,N_12117);
or U14182 (N_14182,N_12050,N_13400);
nor U14183 (N_14183,N_13145,N_12737);
nor U14184 (N_14184,N_12460,N_12873);
nor U14185 (N_14185,N_12079,N_12121);
and U14186 (N_14186,N_13166,N_12814);
or U14187 (N_14187,N_13050,N_12977);
nor U14188 (N_14188,N_12520,N_12305);
and U14189 (N_14189,N_13430,N_13298);
nor U14190 (N_14190,N_12640,N_12940);
nand U14191 (N_14191,N_12808,N_13414);
and U14192 (N_14192,N_13312,N_12092);
and U14193 (N_14193,N_12114,N_12986);
nor U14194 (N_14194,N_12216,N_12661);
and U14195 (N_14195,N_12329,N_13349);
or U14196 (N_14196,N_12408,N_12379);
nand U14197 (N_14197,N_12466,N_12773);
nor U14198 (N_14198,N_12527,N_12173);
or U14199 (N_14199,N_13334,N_13073);
nand U14200 (N_14200,N_12196,N_12627);
nand U14201 (N_14201,N_12215,N_12312);
or U14202 (N_14202,N_12915,N_12469);
nor U14203 (N_14203,N_12909,N_13453);
nand U14204 (N_14204,N_12071,N_12165);
and U14205 (N_14205,N_13321,N_13391);
and U14206 (N_14206,N_12319,N_12883);
and U14207 (N_14207,N_13238,N_12404);
nor U14208 (N_14208,N_12853,N_13407);
xnor U14209 (N_14209,N_13425,N_12826);
nand U14210 (N_14210,N_12825,N_12150);
xor U14211 (N_14211,N_12480,N_12708);
and U14212 (N_14212,N_12008,N_12609);
nand U14213 (N_14213,N_13168,N_12878);
nand U14214 (N_14214,N_13100,N_12401);
nand U14215 (N_14215,N_12063,N_13260);
nand U14216 (N_14216,N_13044,N_13242);
or U14217 (N_14217,N_13041,N_13057);
nand U14218 (N_14218,N_12043,N_13381);
nor U14219 (N_14219,N_13035,N_13339);
nor U14220 (N_14220,N_12372,N_12065);
xor U14221 (N_14221,N_12539,N_12487);
xnor U14222 (N_14222,N_12180,N_12585);
and U14223 (N_14223,N_13197,N_13373);
nor U14224 (N_14224,N_13444,N_12589);
xor U14225 (N_14225,N_12209,N_12301);
nand U14226 (N_14226,N_13473,N_12027);
and U14227 (N_14227,N_12248,N_12447);
or U14228 (N_14228,N_12838,N_13272);
nand U14229 (N_14229,N_12452,N_12757);
nand U14230 (N_14230,N_12009,N_12631);
or U14231 (N_14231,N_12713,N_13210);
and U14232 (N_14232,N_12541,N_13277);
xnor U14233 (N_14233,N_13336,N_12774);
xor U14234 (N_14234,N_12160,N_13015);
and U14235 (N_14235,N_12078,N_13120);
nor U14236 (N_14236,N_12391,N_12081);
and U14237 (N_14237,N_13094,N_12753);
nor U14238 (N_14238,N_13209,N_12687);
nand U14239 (N_14239,N_13454,N_12219);
nand U14240 (N_14240,N_12202,N_13282);
nand U14241 (N_14241,N_13285,N_12837);
xnor U14242 (N_14242,N_13134,N_12610);
nor U14243 (N_14243,N_12350,N_12177);
and U14244 (N_14244,N_12694,N_12685);
or U14245 (N_14245,N_13012,N_12481);
and U14246 (N_14246,N_13496,N_12136);
xor U14247 (N_14247,N_12385,N_12834);
xor U14248 (N_14248,N_12933,N_12815);
xnor U14249 (N_14249,N_13466,N_13048);
or U14250 (N_14250,N_12861,N_12079);
or U14251 (N_14251,N_12690,N_12241);
xnor U14252 (N_14252,N_12464,N_12251);
and U14253 (N_14253,N_13354,N_12494);
nand U14254 (N_14254,N_12705,N_13404);
and U14255 (N_14255,N_13152,N_12514);
or U14256 (N_14256,N_12915,N_12625);
nor U14257 (N_14257,N_12006,N_13088);
and U14258 (N_14258,N_13131,N_13206);
and U14259 (N_14259,N_12328,N_12806);
nor U14260 (N_14260,N_12668,N_12387);
or U14261 (N_14261,N_12463,N_13044);
and U14262 (N_14262,N_13437,N_12171);
xnor U14263 (N_14263,N_12248,N_12769);
or U14264 (N_14264,N_12016,N_12288);
nand U14265 (N_14265,N_12917,N_13075);
or U14266 (N_14266,N_12873,N_13366);
xor U14267 (N_14267,N_13419,N_12219);
and U14268 (N_14268,N_12706,N_12092);
or U14269 (N_14269,N_12810,N_12773);
xnor U14270 (N_14270,N_13480,N_13379);
nand U14271 (N_14271,N_13415,N_12811);
or U14272 (N_14272,N_13079,N_12911);
nor U14273 (N_14273,N_12008,N_12747);
or U14274 (N_14274,N_12996,N_12680);
nand U14275 (N_14275,N_13427,N_12285);
xor U14276 (N_14276,N_13108,N_13449);
or U14277 (N_14277,N_12976,N_12245);
nor U14278 (N_14278,N_12413,N_13178);
nand U14279 (N_14279,N_13095,N_12121);
xor U14280 (N_14280,N_12384,N_12070);
and U14281 (N_14281,N_12387,N_12879);
nor U14282 (N_14282,N_12735,N_12460);
nor U14283 (N_14283,N_12770,N_13224);
nand U14284 (N_14284,N_12869,N_12863);
or U14285 (N_14285,N_12294,N_13259);
xnor U14286 (N_14286,N_12139,N_13314);
and U14287 (N_14287,N_12302,N_12318);
xnor U14288 (N_14288,N_13460,N_12384);
and U14289 (N_14289,N_12995,N_12363);
or U14290 (N_14290,N_13294,N_12469);
xnor U14291 (N_14291,N_13046,N_12102);
xor U14292 (N_14292,N_12303,N_12089);
nand U14293 (N_14293,N_13225,N_13103);
nor U14294 (N_14294,N_12935,N_12529);
or U14295 (N_14295,N_13357,N_12698);
nand U14296 (N_14296,N_12764,N_12321);
xnor U14297 (N_14297,N_12285,N_12570);
and U14298 (N_14298,N_12395,N_12434);
nor U14299 (N_14299,N_12003,N_12991);
nand U14300 (N_14300,N_12728,N_12198);
nor U14301 (N_14301,N_13022,N_13194);
and U14302 (N_14302,N_13137,N_12934);
nand U14303 (N_14303,N_12879,N_13220);
and U14304 (N_14304,N_12802,N_13185);
nand U14305 (N_14305,N_12400,N_13033);
nor U14306 (N_14306,N_13108,N_12956);
or U14307 (N_14307,N_13305,N_12797);
nor U14308 (N_14308,N_13081,N_12725);
and U14309 (N_14309,N_12443,N_13144);
or U14310 (N_14310,N_12225,N_12585);
and U14311 (N_14311,N_12760,N_12147);
nor U14312 (N_14312,N_12186,N_12411);
xor U14313 (N_14313,N_12758,N_13423);
nor U14314 (N_14314,N_13365,N_13122);
nor U14315 (N_14315,N_13159,N_13079);
nand U14316 (N_14316,N_12295,N_12234);
nand U14317 (N_14317,N_12215,N_12868);
and U14318 (N_14318,N_12571,N_12917);
xor U14319 (N_14319,N_13346,N_13074);
nor U14320 (N_14320,N_13488,N_13243);
nand U14321 (N_14321,N_12354,N_12370);
nor U14322 (N_14322,N_12933,N_13352);
or U14323 (N_14323,N_12789,N_13304);
or U14324 (N_14324,N_13368,N_12358);
nor U14325 (N_14325,N_12402,N_12750);
or U14326 (N_14326,N_12521,N_13327);
and U14327 (N_14327,N_12576,N_13152);
nor U14328 (N_14328,N_12044,N_12185);
nor U14329 (N_14329,N_13390,N_13294);
xnor U14330 (N_14330,N_12478,N_12787);
or U14331 (N_14331,N_12164,N_13043);
nand U14332 (N_14332,N_12001,N_13028);
or U14333 (N_14333,N_12644,N_13269);
nor U14334 (N_14334,N_12406,N_13004);
nand U14335 (N_14335,N_13449,N_12929);
and U14336 (N_14336,N_12672,N_12830);
nand U14337 (N_14337,N_12522,N_12972);
nor U14338 (N_14338,N_12774,N_12552);
nor U14339 (N_14339,N_13445,N_12671);
xnor U14340 (N_14340,N_13312,N_12031);
or U14341 (N_14341,N_13440,N_12203);
and U14342 (N_14342,N_13057,N_12687);
xnor U14343 (N_14343,N_12868,N_12306);
nor U14344 (N_14344,N_13373,N_12751);
nand U14345 (N_14345,N_12902,N_13150);
and U14346 (N_14346,N_12896,N_13026);
or U14347 (N_14347,N_13303,N_12942);
nor U14348 (N_14348,N_12247,N_12517);
xnor U14349 (N_14349,N_12649,N_13037);
xor U14350 (N_14350,N_13160,N_12866);
or U14351 (N_14351,N_13290,N_13070);
xnor U14352 (N_14352,N_12563,N_13020);
or U14353 (N_14353,N_13104,N_12744);
nand U14354 (N_14354,N_12972,N_12057);
xor U14355 (N_14355,N_12101,N_12582);
nor U14356 (N_14356,N_13265,N_12057);
nand U14357 (N_14357,N_12638,N_13284);
nand U14358 (N_14358,N_13132,N_12138);
nor U14359 (N_14359,N_12974,N_12470);
and U14360 (N_14360,N_12797,N_13495);
or U14361 (N_14361,N_12487,N_12622);
nor U14362 (N_14362,N_12378,N_13150);
xnor U14363 (N_14363,N_12785,N_12194);
and U14364 (N_14364,N_13361,N_12443);
and U14365 (N_14365,N_12099,N_13456);
nand U14366 (N_14366,N_13272,N_12468);
nor U14367 (N_14367,N_12717,N_13230);
or U14368 (N_14368,N_12523,N_13053);
nor U14369 (N_14369,N_12135,N_12151);
nand U14370 (N_14370,N_13018,N_12382);
nand U14371 (N_14371,N_12155,N_13493);
nor U14372 (N_14372,N_13123,N_12027);
or U14373 (N_14373,N_12554,N_12224);
xnor U14374 (N_14374,N_12910,N_13317);
xnor U14375 (N_14375,N_12939,N_13271);
nor U14376 (N_14376,N_12339,N_12668);
xor U14377 (N_14377,N_13282,N_12768);
xnor U14378 (N_14378,N_12028,N_12495);
and U14379 (N_14379,N_13242,N_13301);
nor U14380 (N_14380,N_12049,N_13276);
or U14381 (N_14381,N_12855,N_12148);
nor U14382 (N_14382,N_13057,N_12198);
or U14383 (N_14383,N_12986,N_13207);
or U14384 (N_14384,N_12096,N_12257);
xnor U14385 (N_14385,N_13386,N_12007);
nand U14386 (N_14386,N_13178,N_13023);
nand U14387 (N_14387,N_12701,N_12620);
nor U14388 (N_14388,N_13457,N_12360);
and U14389 (N_14389,N_12593,N_12323);
xnor U14390 (N_14390,N_12744,N_12934);
xor U14391 (N_14391,N_12524,N_12715);
and U14392 (N_14392,N_12734,N_12831);
or U14393 (N_14393,N_13461,N_12903);
nor U14394 (N_14394,N_12398,N_12184);
or U14395 (N_14395,N_13347,N_12824);
nor U14396 (N_14396,N_12529,N_12951);
xnor U14397 (N_14397,N_12495,N_12441);
nand U14398 (N_14398,N_13148,N_13391);
nor U14399 (N_14399,N_12748,N_12488);
xor U14400 (N_14400,N_12773,N_12868);
and U14401 (N_14401,N_12463,N_13030);
or U14402 (N_14402,N_12963,N_12735);
or U14403 (N_14403,N_12661,N_12434);
and U14404 (N_14404,N_12911,N_12929);
nor U14405 (N_14405,N_12900,N_13362);
or U14406 (N_14406,N_12679,N_13365);
nor U14407 (N_14407,N_12952,N_13101);
nand U14408 (N_14408,N_12841,N_12429);
nor U14409 (N_14409,N_12892,N_13148);
nor U14410 (N_14410,N_12037,N_12929);
nor U14411 (N_14411,N_12415,N_13266);
xnor U14412 (N_14412,N_12072,N_12186);
or U14413 (N_14413,N_13476,N_12713);
or U14414 (N_14414,N_12902,N_13380);
or U14415 (N_14415,N_12380,N_12236);
or U14416 (N_14416,N_12012,N_12035);
xnor U14417 (N_14417,N_13495,N_12828);
or U14418 (N_14418,N_13197,N_13250);
and U14419 (N_14419,N_12479,N_12368);
xor U14420 (N_14420,N_12013,N_13270);
xor U14421 (N_14421,N_12633,N_12339);
nor U14422 (N_14422,N_13150,N_12205);
or U14423 (N_14423,N_12377,N_13479);
nor U14424 (N_14424,N_13042,N_13255);
xor U14425 (N_14425,N_12193,N_13363);
xor U14426 (N_14426,N_13462,N_13072);
nor U14427 (N_14427,N_12397,N_12063);
or U14428 (N_14428,N_13019,N_13086);
or U14429 (N_14429,N_13230,N_12982);
nand U14430 (N_14430,N_12769,N_12637);
and U14431 (N_14431,N_12654,N_12594);
nand U14432 (N_14432,N_12967,N_13275);
and U14433 (N_14433,N_12589,N_13002);
or U14434 (N_14434,N_12376,N_12621);
xor U14435 (N_14435,N_12579,N_12474);
and U14436 (N_14436,N_12242,N_13136);
and U14437 (N_14437,N_13254,N_12760);
nand U14438 (N_14438,N_12902,N_12716);
xor U14439 (N_14439,N_12791,N_12093);
and U14440 (N_14440,N_13255,N_13286);
or U14441 (N_14441,N_12536,N_12881);
xor U14442 (N_14442,N_12086,N_12575);
nand U14443 (N_14443,N_12505,N_12345);
and U14444 (N_14444,N_13062,N_12442);
or U14445 (N_14445,N_13404,N_12617);
nor U14446 (N_14446,N_12241,N_12337);
nor U14447 (N_14447,N_13497,N_13007);
nor U14448 (N_14448,N_12981,N_13098);
and U14449 (N_14449,N_12045,N_13282);
and U14450 (N_14450,N_13134,N_12951);
or U14451 (N_14451,N_12023,N_12880);
nand U14452 (N_14452,N_13420,N_12995);
nand U14453 (N_14453,N_13430,N_12731);
xnor U14454 (N_14454,N_13491,N_13268);
or U14455 (N_14455,N_12285,N_12772);
xnor U14456 (N_14456,N_12034,N_12018);
and U14457 (N_14457,N_12489,N_12127);
xnor U14458 (N_14458,N_12184,N_13151);
nand U14459 (N_14459,N_12972,N_13128);
nand U14460 (N_14460,N_13353,N_13275);
and U14461 (N_14461,N_12543,N_12125);
nand U14462 (N_14462,N_12022,N_12420);
or U14463 (N_14463,N_12876,N_12636);
nor U14464 (N_14464,N_13245,N_12875);
nand U14465 (N_14465,N_12117,N_13197);
or U14466 (N_14466,N_12083,N_12950);
and U14467 (N_14467,N_12618,N_13029);
xnor U14468 (N_14468,N_12930,N_13083);
nand U14469 (N_14469,N_13128,N_13392);
nand U14470 (N_14470,N_12404,N_12374);
or U14471 (N_14471,N_12829,N_13090);
nor U14472 (N_14472,N_12684,N_13400);
and U14473 (N_14473,N_12255,N_12941);
or U14474 (N_14474,N_13421,N_12157);
xor U14475 (N_14475,N_12615,N_12175);
nand U14476 (N_14476,N_13461,N_13311);
nand U14477 (N_14477,N_12292,N_12965);
xnor U14478 (N_14478,N_13423,N_12978);
and U14479 (N_14479,N_13408,N_13279);
or U14480 (N_14480,N_13159,N_12824);
nor U14481 (N_14481,N_12121,N_13344);
nand U14482 (N_14482,N_13261,N_13119);
xor U14483 (N_14483,N_12877,N_12536);
nor U14484 (N_14484,N_13163,N_12134);
or U14485 (N_14485,N_12630,N_12556);
nor U14486 (N_14486,N_12639,N_12398);
xnor U14487 (N_14487,N_13082,N_12759);
or U14488 (N_14488,N_13000,N_12637);
nor U14489 (N_14489,N_12890,N_13044);
and U14490 (N_14490,N_12716,N_12646);
nand U14491 (N_14491,N_12723,N_12155);
xnor U14492 (N_14492,N_12300,N_13058);
nand U14493 (N_14493,N_12649,N_13021);
or U14494 (N_14494,N_12131,N_12178);
and U14495 (N_14495,N_13381,N_13055);
nor U14496 (N_14496,N_12861,N_12424);
xor U14497 (N_14497,N_13270,N_12709);
xnor U14498 (N_14498,N_12530,N_12124);
nor U14499 (N_14499,N_12462,N_12364);
nor U14500 (N_14500,N_12134,N_13333);
nor U14501 (N_14501,N_13373,N_12590);
or U14502 (N_14502,N_13378,N_12205);
nor U14503 (N_14503,N_12036,N_12236);
xor U14504 (N_14504,N_12782,N_12059);
xnor U14505 (N_14505,N_13058,N_12317);
xnor U14506 (N_14506,N_12657,N_12577);
and U14507 (N_14507,N_12892,N_13462);
xor U14508 (N_14508,N_12948,N_12324);
nor U14509 (N_14509,N_13456,N_13141);
nand U14510 (N_14510,N_12600,N_12876);
nor U14511 (N_14511,N_12130,N_12552);
nor U14512 (N_14512,N_12346,N_12072);
or U14513 (N_14513,N_12498,N_12296);
nand U14514 (N_14514,N_12068,N_13275);
and U14515 (N_14515,N_13188,N_12010);
or U14516 (N_14516,N_13283,N_12206);
xnor U14517 (N_14517,N_12381,N_13495);
or U14518 (N_14518,N_12251,N_13257);
xor U14519 (N_14519,N_12310,N_13206);
and U14520 (N_14520,N_13495,N_12457);
nor U14521 (N_14521,N_12046,N_13221);
nand U14522 (N_14522,N_13352,N_12668);
and U14523 (N_14523,N_13339,N_12220);
xor U14524 (N_14524,N_12321,N_12582);
xor U14525 (N_14525,N_13088,N_12092);
xnor U14526 (N_14526,N_13052,N_13004);
nand U14527 (N_14527,N_12874,N_12000);
and U14528 (N_14528,N_13139,N_12604);
and U14529 (N_14529,N_12379,N_12336);
xor U14530 (N_14530,N_12834,N_13066);
and U14531 (N_14531,N_12767,N_13109);
nor U14532 (N_14532,N_12944,N_12671);
nand U14533 (N_14533,N_12024,N_12234);
xor U14534 (N_14534,N_13336,N_12824);
and U14535 (N_14535,N_12106,N_12303);
or U14536 (N_14536,N_12340,N_12937);
nor U14537 (N_14537,N_12496,N_12771);
xor U14538 (N_14538,N_13293,N_12851);
xor U14539 (N_14539,N_12992,N_12879);
nand U14540 (N_14540,N_13202,N_12319);
nand U14541 (N_14541,N_12515,N_12669);
or U14542 (N_14542,N_12307,N_13069);
or U14543 (N_14543,N_13363,N_12691);
or U14544 (N_14544,N_12839,N_12200);
and U14545 (N_14545,N_12400,N_12160);
nand U14546 (N_14546,N_13268,N_12069);
nor U14547 (N_14547,N_12087,N_12306);
nand U14548 (N_14548,N_12632,N_12173);
xnor U14549 (N_14549,N_12000,N_12545);
xor U14550 (N_14550,N_13496,N_12385);
xor U14551 (N_14551,N_12466,N_12949);
xnor U14552 (N_14552,N_12004,N_12264);
and U14553 (N_14553,N_12644,N_13270);
and U14554 (N_14554,N_12809,N_12922);
or U14555 (N_14555,N_12709,N_12453);
nand U14556 (N_14556,N_13345,N_12594);
xnor U14557 (N_14557,N_12509,N_12041);
and U14558 (N_14558,N_12675,N_13334);
and U14559 (N_14559,N_13165,N_13414);
and U14560 (N_14560,N_12490,N_12102);
nand U14561 (N_14561,N_12498,N_12754);
and U14562 (N_14562,N_12747,N_12723);
nor U14563 (N_14563,N_12077,N_12308);
nor U14564 (N_14564,N_13442,N_13252);
nand U14565 (N_14565,N_12564,N_12466);
nor U14566 (N_14566,N_13161,N_12784);
and U14567 (N_14567,N_12129,N_12190);
and U14568 (N_14568,N_12545,N_13128);
nor U14569 (N_14569,N_13365,N_13190);
xor U14570 (N_14570,N_12550,N_12618);
xor U14571 (N_14571,N_12653,N_13115);
nand U14572 (N_14572,N_12372,N_12379);
and U14573 (N_14573,N_12169,N_13161);
nand U14574 (N_14574,N_13214,N_13080);
nor U14575 (N_14575,N_12223,N_12463);
and U14576 (N_14576,N_13072,N_12107);
xnor U14577 (N_14577,N_12198,N_12236);
nand U14578 (N_14578,N_13189,N_13219);
xnor U14579 (N_14579,N_13210,N_13451);
nor U14580 (N_14580,N_12807,N_12247);
and U14581 (N_14581,N_13184,N_12769);
or U14582 (N_14582,N_13095,N_13410);
xor U14583 (N_14583,N_12297,N_13371);
and U14584 (N_14584,N_13196,N_12245);
xnor U14585 (N_14585,N_12029,N_12333);
and U14586 (N_14586,N_12153,N_12070);
and U14587 (N_14587,N_12487,N_13423);
xnor U14588 (N_14588,N_12735,N_12693);
nand U14589 (N_14589,N_12199,N_13423);
nor U14590 (N_14590,N_12894,N_13480);
and U14591 (N_14591,N_13232,N_12586);
nor U14592 (N_14592,N_12473,N_13339);
nor U14593 (N_14593,N_12006,N_12993);
and U14594 (N_14594,N_13372,N_12349);
and U14595 (N_14595,N_12054,N_12447);
nand U14596 (N_14596,N_12098,N_12797);
nor U14597 (N_14597,N_13168,N_12603);
nor U14598 (N_14598,N_13044,N_13016);
or U14599 (N_14599,N_12236,N_12113);
nand U14600 (N_14600,N_12608,N_12006);
and U14601 (N_14601,N_12462,N_13384);
nand U14602 (N_14602,N_13143,N_12749);
or U14603 (N_14603,N_13278,N_12781);
and U14604 (N_14604,N_13180,N_12661);
nor U14605 (N_14605,N_12114,N_13330);
and U14606 (N_14606,N_13111,N_13473);
nor U14607 (N_14607,N_13128,N_12563);
nor U14608 (N_14608,N_12865,N_12210);
or U14609 (N_14609,N_12695,N_13181);
nand U14610 (N_14610,N_12594,N_13221);
or U14611 (N_14611,N_12900,N_12090);
nand U14612 (N_14612,N_13237,N_12961);
or U14613 (N_14613,N_12452,N_12513);
and U14614 (N_14614,N_13434,N_12356);
or U14615 (N_14615,N_12721,N_12671);
nor U14616 (N_14616,N_12753,N_13029);
xor U14617 (N_14617,N_12446,N_12590);
nand U14618 (N_14618,N_12174,N_12230);
nand U14619 (N_14619,N_13253,N_13075);
or U14620 (N_14620,N_12941,N_12171);
nor U14621 (N_14621,N_12923,N_13110);
xor U14622 (N_14622,N_13156,N_12081);
nor U14623 (N_14623,N_12267,N_12794);
xnor U14624 (N_14624,N_12215,N_12645);
and U14625 (N_14625,N_12009,N_12564);
xnor U14626 (N_14626,N_12814,N_13250);
nand U14627 (N_14627,N_12044,N_12704);
and U14628 (N_14628,N_12708,N_12461);
xnor U14629 (N_14629,N_12138,N_13211);
nor U14630 (N_14630,N_12962,N_13498);
nand U14631 (N_14631,N_13066,N_12429);
and U14632 (N_14632,N_12206,N_12688);
nand U14633 (N_14633,N_12550,N_12483);
or U14634 (N_14634,N_13090,N_13386);
and U14635 (N_14635,N_13121,N_12759);
nor U14636 (N_14636,N_13426,N_13433);
xnor U14637 (N_14637,N_12679,N_12350);
nand U14638 (N_14638,N_12866,N_12704);
nor U14639 (N_14639,N_13196,N_12742);
xnor U14640 (N_14640,N_12795,N_12986);
or U14641 (N_14641,N_12783,N_12605);
or U14642 (N_14642,N_13167,N_12681);
nor U14643 (N_14643,N_12358,N_13374);
nor U14644 (N_14644,N_13354,N_13386);
xnor U14645 (N_14645,N_12400,N_13208);
nand U14646 (N_14646,N_13053,N_12070);
or U14647 (N_14647,N_12741,N_12308);
nand U14648 (N_14648,N_12407,N_12446);
or U14649 (N_14649,N_12249,N_12240);
nor U14650 (N_14650,N_12161,N_12259);
nand U14651 (N_14651,N_12674,N_12894);
and U14652 (N_14652,N_13093,N_12593);
and U14653 (N_14653,N_12315,N_13403);
nand U14654 (N_14654,N_12967,N_13034);
xor U14655 (N_14655,N_12676,N_12354);
nor U14656 (N_14656,N_12597,N_13498);
xor U14657 (N_14657,N_12918,N_12008);
xnor U14658 (N_14658,N_12612,N_13396);
nand U14659 (N_14659,N_13459,N_12479);
nand U14660 (N_14660,N_12869,N_12499);
nor U14661 (N_14661,N_12766,N_12247);
and U14662 (N_14662,N_12542,N_13116);
nand U14663 (N_14663,N_13450,N_12861);
and U14664 (N_14664,N_12391,N_12933);
and U14665 (N_14665,N_12221,N_12364);
nand U14666 (N_14666,N_12702,N_12210);
nor U14667 (N_14667,N_13071,N_12616);
xor U14668 (N_14668,N_12727,N_12397);
and U14669 (N_14669,N_12330,N_13365);
or U14670 (N_14670,N_13466,N_13404);
nand U14671 (N_14671,N_12269,N_12240);
nand U14672 (N_14672,N_12729,N_12781);
and U14673 (N_14673,N_12913,N_12771);
and U14674 (N_14674,N_12977,N_12116);
xor U14675 (N_14675,N_13371,N_13167);
nor U14676 (N_14676,N_12683,N_12925);
or U14677 (N_14677,N_13290,N_13334);
xnor U14678 (N_14678,N_13006,N_12124);
nand U14679 (N_14679,N_13453,N_13401);
or U14680 (N_14680,N_12288,N_13068);
nor U14681 (N_14681,N_13305,N_13459);
xnor U14682 (N_14682,N_13346,N_12480);
nand U14683 (N_14683,N_12197,N_12937);
or U14684 (N_14684,N_12329,N_12250);
and U14685 (N_14685,N_12343,N_12262);
nand U14686 (N_14686,N_12345,N_12008);
xnor U14687 (N_14687,N_13350,N_12144);
nor U14688 (N_14688,N_12512,N_12373);
and U14689 (N_14689,N_12856,N_12332);
xor U14690 (N_14690,N_12015,N_13238);
and U14691 (N_14691,N_12762,N_12484);
or U14692 (N_14692,N_13145,N_12809);
nor U14693 (N_14693,N_12805,N_13458);
and U14694 (N_14694,N_12740,N_13172);
or U14695 (N_14695,N_12805,N_12260);
or U14696 (N_14696,N_13372,N_12674);
nand U14697 (N_14697,N_12510,N_13003);
and U14698 (N_14698,N_12908,N_12446);
and U14699 (N_14699,N_12675,N_13370);
nand U14700 (N_14700,N_13159,N_13146);
nor U14701 (N_14701,N_12956,N_12648);
nor U14702 (N_14702,N_12684,N_13057);
nand U14703 (N_14703,N_13448,N_12591);
or U14704 (N_14704,N_12864,N_13076);
xnor U14705 (N_14705,N_13026,N_12121);
xnor U14706 (N_14706,N_12007,N_12870);
nand U14707 (N_14707,N_12333,N_12354);
xor U14708 (N_14708,N_12549,N_13270);
nor U14709 (N_14709,N_12595,N_12964);
nand U14710 (N_14710,N_13331,N_12819);
or U14711 (N_14711,N_12922,N_12537);
or U14712 (N_14712,N_12545,N_12731);
nor U14713 (N_14713,N_12363,N_12369);
nand U14714 (N_14714,N_13097,N_12369);
nand U14715 (N_14715,N_13058,N_12278);
or U14716 (N_14716,N_12847,N_12113);
nand U14717 (N_14717,N_12660,N_12730);
or U14718 (N_14718,N_12835,N_12232);
xnor U14719 (N_14719,N_12803,N_13090);
and U14720 (N_14720,N_12765,N_12940);
nand U14721 (N_14721,N_12010,N_12856);
nor U14722 (N_14722,N_12754,N_12341);
and U14723 (N_14723,N_13382,N_13283);
nand U14724 (N_14724,N_13265,N_12805);
nand U14725 (N_14725,N_13008,N_13372);
nor U14726 (N_14726,N_13154,N_13313);
nor U14727 (N_14727,N_13285,N_12748);
and U14728 (N_14728,N_12937,N_12306);
xor U14729 (N_14729,N_13161,N_13018);
nand U14730 (N_14730,N_13431,N_12429);
xnor U14731 (N_14731,N_12791,N_13041);
nand U14732 (N_14732,N_12943,N_12011);
xnor U14733 (N_14733,N_12177,N_12656);
nor U14734 (N_14734,N_12972,N_12161);
nand U14735 (N_14735,N_12476,N_12098);
xnor U14736 (N_14736,N_13166,N_12279);
xor U14737 (N_14737,N_12744,N_13118);
or U14738 (N_14738,N_12452,N_12765);
or U14739 (N_14739,N_12113,N_12257);
and U14740 (N_14740,N_13314,N_12729);
xnor U14741 (N_14741,N_12054,N_12634);
nor U14742 (N_14742,N_13193,N_12624);
nor U14743 (N_14743,N_12239,N_12997);
and U14744 (N_14744,N_12285,N_12112);
xor U14745 (N_14745,N_13405,N_13145);
nand U14746 (N_14746,N_13413,N_13420);
nand U14747 (N_14747,N_12806,N_13265);
or U14748 (N_14748,N_12886,N_12151);
nor U14749 (N_14749,N_12293,N_12010);
nor U14750 (N_14750,N_12677,N_12306);
nor U14751 (N_14751,N_12366,N_12548);
and U14752 (N_14752,N_12872,N_13338);
and U14753 (N_14753,N_12358,N_12590);
or U14754 (N_14754,N_12365,N_12588);
nand U14755 (N_14755,N_12246,N_12565);
or U14756 (N_14756,N_12944,N_13223);
nand U14757 (N_14757,N_13377,N_13072);
or U14758 (N_14758,N_12861,N_13309);
and U14759 (N_14759,N_13224,N_12254);
nand U14760 (N_14760,N_12059,N_12058);
nand U14761 (N_14761,N_13283,N_12160);
or U14762 (N_14762,N_13155,N_13225);
nor U14763 (N_14763,N_12271,N_12175);
nand U14764 (N_14764,N_13474,N_12531);
and U14765 (N_14765,N_12852,N_13191);
and U14766 (N_14766,N_12230,N_12001);
and U14767 (N_14767,N_12645,N_12377);
nor U14768 (N_14768,N_13434,N_12839);
nor U14769 (N_14769,N_12503,N_13496);
nand U14770 (N_14770,N_13321,N_12137);
nor U14771 (N_14771,N_12481,N_12906);
xor U14772 (N_14772,N_12268,N_12969);
nor U14773 (N_14773,N_13286,N_12253);
nor U14774 (N_14774,N_12236,N_13358);
nand U14775 (N_14775,N_12243,N_12159);
or U14776 (N_14776,N_12406,N_12780);
nor U14777 (N_14777,N_12902,N_12094);
nand U14778 (N_14778,N_12860,N_12829);
nor U14779 (N_14779,N_13146,N_13463);
xor U14780 (N_14780,N_12681,N_13261);
xnor U14781 (N_14781,N_13131,N_12564);
xnor U14782 (N_14782,N_13113,N_12638);
nor U14783 (N_14783,N_13002,N_12692);
or U14784 (N_14784,N_13123,N_12382);
nor U14785 (N_14785,N_12999,N_12444);
and U14786 (N_14786,N_12173,N_12578);
nand U14787 (N_14787,N_13202,N_12165);
xor U14788 (N_14788,N_12610,N_12515);
and U14789 (N_14789,N_12878,N_13474);
nor U14790 (N_14790,N_13155,N_12839);
or U14791 (N_14791,N_13207,N_12201);
xor U14792 (N_14792,N_12313,N_13180);
nor U14793 (N_14793,N_12878,N_13289);
or U14794 (N_14794,N_12566,N_12030);
xnor U14795 (N_14795,N_13314,N_12021);
or U14796 (N_14796,N_12174,N_12390);
xnor U14797 (N_14797,N_13348,N_13178);
nand U14798 (N_14798,N_12866,N_12215);
xnor U14799 (N_14799,N_12320,N_12954);
or U14800 (N_14800,N_13051,N_13493);
nand U14801 (N_14801,N_12786,N_13161);
nand U14802 (N_14802,N_13401,N_12663);
and U14803 (N_14803,N_12958,N_13385);
or U14804 (N_14804,N_13249,N_13174);
nor U14805 (N_14805,N_12487,N_12977);
xor U14806 (N_14806,N_12178,N_13314);
and U14807 (N_14807,N_12137,N_12590);
and U14808 (N_14808,N_12975,N_13152);
nor U14809 (N_14809,N_12358,N_13262);
or U14810 (N_14810,N_13126,N_12553);
nand U14811 (N_14811,N_12336,N_12687);
nand U14812 (N_14812,N_12030,N_12961);
or U14813 (N_14813,N_13054,N_13311);
or U14814 (N_14814,N_12159,N_12918);
and U14815 (N_14815,N_12059,N_12717);
nand U14816 (N_14816,N_13431,N_12406);
nor U14817 (N_14817,N_13033,N_12705);
nor U14818 (N_14818,N_13071,N_13060);
xor U14819 (N_14819,N_12463,N_13084);
nand U14820 (N_14820,N_12903,N_12562);
nor U14821 (N_14821,N_12415,N_13067);
and U14822 (N_14822,N_13175,N_12299);
nand U14823 (N_14823,N_12219,N_12238);
or U14824 (N_14824,N_12369,N_13288);
xor U14825 (N_14825,N_13241,N_12452);
or U14826 (N_14826,N_12938,N_12866);
and U14827 (N_14827,N_12764,N_12490);
nor U14828 (N_14828,N_12525,N_12231);
xor U14829 (N_14829,N_12773,N_12483);
nor U14830 (N_14830,N_13436,N_12995);
or U14831 (N_14831,N_12111,N_12957);
nor U14832 (N_14832,N_12996,N_13124);
and U14833 (N_14833,N_12012,N_12897);
or U14834 (N_14834,N_12984,N_12811);
or U14835 (N_14835,N_12182,N_13033);
nand U14836 (N_14836,N_12332,N_12544);
or U14837 (N_14837,N_12667,N_12203);
nor U14838 (N_14838,N_12830,N_12351);
and U14839 (N_14839,N_12601,N_13256);
nand U14840 (N_14840,N_13361,N_12878);
nor U14841 (N_14841,N_12630,N_12365);
xor U14842 (N_14842,N_12604,N_12382);
and U14843 (N_14843,N_12159,N_12246);
nand U14844 (N_14844,N_13110,N_13325);
nand U14845 (N_14845,N_12673,N_12922);
or U14846 (N_14846,N_13498,N_13119);
xor U14847 (N_14847,N_12516,N_12923);
nand U14848 (N_14848,N_12961,N_12989);
xor U14849 (N_14849,N_12620,N_12634);
xnor U14850 (N_14850,N_12859,N_12251);
nand U14851 (N_14851,N_12675,N_12509);
or U14852 (N_14852,N_12068,N_13199);
or U14853 (N_14853,N_13348,N_12003);
and U14854 (N_14854,N_12320,N_12021);
or U14855 (N_14855,N_13009,N_13012);
nand U14856 (N_14856,N_13391,N_12581);
or U14857 (N_14857,N_13020,N_13091);
nor U14858 (N_14858,N_12386,N_12074);
or U14859 (N_14859,N_12948,N_12481);
and U14860 (N_14860,N_13108,N_12177);
nand U14861 (N_14861,N_12134,N_12551);
nand U14862 (N_14862,N_12148,N_12217);
nor U14863 (N_14863,N_12239,N_12856);
or U14864 (N_14864,N_13125,N_12727);
nand U14865 (N_14865,N_12264,N_13452);
or U14866 (N_14866,N_13483,N_12823);
and U14867 (N_14867,N_12598,N_12362);
and U14868 (N_14868,N_12485,N_12691);
or U14869 (N_14869,N_12653,N_12621);
or U14870 (N_14870,N_12562,N_12143);
xor U14871 (N_14871,N_12181,N_12997);
nand U14872 (N_14872,N_13056,N_12294);
and U14873 (N_14873,N_12340,N_12099);
or U14874 (N_14874,N_13082,N_13373);
xnor U14875 (N_14875,N_13155,N_12438);
and U14876 (N_14876,N_12380,N_13166);
or U14877 (N_14877,N_13218,N_13401);
or U14878 (N_14878,N_12197,N_13416);
xnor U14879 (N_14879,N_13293,N_13181);
xnor U14880 (N_14880,N_13154,N_12897);
xnor U14881 (N_14881,N_12028,N_12715);
nand U14882 (N_14882,N_12561,N_12966);
nor U14883 (N_14883,N_12484,N_13169);
nand U14884 (N_14884,N_13218,N_12868);
or U14885 (N_14885,N_12560,N_12104);
or U14886 (N_14886,N_13214,N_12715);
nand U14887 (N_14887,N_12096,N_13391);
and U14888 (N_14888,N_12134,N_12294);
nor U14889 (N_14889,N_12222,N_12014);
or U14890 (N_14890,N_13488,N_12885);
nor U14891 (N_14891,N_12327,N_13483);
xor U14892 (N_14892,N_12653,N_12945);
and U14893 (N_14893,N_12668,N_12426);
or U14894 (N_14894,N_13470,N_13302);
xnor U14895 (N_14895,N_13177,N_12984);
nand U14896 (N_14896,N_12228,N_12148);
xor U14897 (N_14897,N_12972,N_12213);
nand U14898 (N_14898,N_13374,N_13042);
or U14899 (N_14899,N_12730,N_12878);
xor U14900 (N_14900,N_12082,N_12420);
or U14901 (N_14901,N_12177,N_12822);
nand U14902 (N_14902,N_13388,N_12313);
and U14903 (N_14903,N_13462,N_12514);
xnor U14904 (N_14904,N_13044,N_12299);
or U14905 (N_14905,N_13189,N_12754);
xnor U14906 (N_14906,N_12238,N_12754);
and U14907 (N_14907,N_12066,N_12611);
nor U14908 (N_14908,N_13284,N_12662);
xor U14909 (N_14909,N_13353,N_12424);
nand U14910 (N_14910,N_13396,N_12646);
and U14911 (N_14911,N_12708,N_12483);
nand U14912 (N_14912,N_13084,N_12973);
xor U14913 (N_14913,N_12386,N_12242);
xnor U14914 (N_14914,N_12593,N_12809);
or U14915 (N_14915,N_12837,N_12880);
nand U14916 (N_14916,N_12475,N_12756);
nor U14917 (N_14917,N_13434,N_13097);
xnor U14918 (N_14918,N_13143,N_12986);
and U14919 (N_14919,N_12799,N_12222);
nor U14920 (N_14920,N_12985,N_13026);
nor U14921 (N_14921,N_13161,N_13001);
and U14922 (N_14922,N_12736,N_12398);
and U14923 (N_14923,N_12108,N_13060);
nand U14924 (N_14924,N_13274,N_12628);
nor U14925 (N_14925,N_13211,N_12403);
nand U14926 (N_14926,N_13117,N_13131);
and U14927 (N_14927,N_12635,N_12304);
nor U14928 (N_14928,N_12152,N_13213);
nand U14929 (N_14929,N_12021,N_13309);
xnor U14930 (N_14930,N_12216,N_12562);
nand U14931 (N_14931,N_12068,N_12596);
or U14932 (N_14932,N_12008,N_13306);
nor U14933 (N_14933,N_13231,N_12900);
xor U14934 (N_14934,N_12265,N_12067);
xnor U14935 (N_14935,N_13168,N_13338);
nand U14936 (N_14936,N_13245,N_12390);
and U14937 (N_14937,N_12674,N_13417);
xor U14938 (N_14938,N_13017,N_13213);
and U14939 (N_14939,N_12036,N_12144);
nand U14940 (N_14940,N_13325,N_13149);
xnor U14941 (N_14941,N_12121,N_12478);
or U14942 (N_14942,N_13215,N_12803);
xor U14943 (N_14943,N_13385,N_13013);
xor U14944 (N_14944,N_12559,N_12767);
nand U14945 (N_14945,N_12805,N_12621);
nor U14946 (N_14946,N_13442,N_13268);
nand U14947 (N_14947,N_13230,N_13362);
and U14948 (N_14948,N_12216,N_12560);
nor U14949 (N_14949,N_13232,N_12736);
xnor U14950 (N_14950,N_13184,N_12215);
xor U14951 (N_14951,N_12140,N_12289);
nor U14952 (N_14952,N_13274,N_13398);
nor U14953 (N_14953,N_12712,N_12988);
nand U14954 (N_14954,N_13081,N_12116);
or U14955 (N_14955,N_12974,N_12781);
nand U14956 (N_14956,N_12520,N_12779);
and U14957 (N_14957,N_12836,N_12004);
and U14958 (N_14958,N_12359,N_12080);
or U14959 (N_14959,N_12694,N_12797);
and U14960 (N_14960,N_12730,N_13318);
nor U14961 (N_14961,N_13370,N_12945);
nor U14962 (N_14962,N_12184,N_12426);
nand U14963 (N_14963,N_12208,N_13495);
or U14964 (N_14964,N_12570,N_12171);
and U14965 (N_14965,N_13191,N_12679);
nand U14966 (N_14966,N_12662,N_13119);
and U14967 (N_14967,N_12192,N_13317);
xor U14968 (N_14968,N_12711,N_12415);
and U14969 (N_14969,N_13162,N_13123);
nor U14970 (N_14970,N_12962,N_12885);
or U14971 (N_14971,N_12962,N_12383);
nand U14972 (N_14972,N_12706,N_12687);
xor U14973 (N_14973,N_12838,N_13186);
nor U14974 (N_14974,N_13273,N_13413);
nor U14975 (N_14975,N_12773,N_13263);
nor U14976 (N_14976,N_12271,N_12263);
xor U14977 (N_14977,N_13063,N_12825);
nand U14978 (N_14978,N_12016,N_12067);
and U14979 (N_14979,N_12812,N_12026);
xor U14980 (N_14980,N_13161,N_12201);
or U14981 (N_14981,N_13136,N_12322);
nand U14982 (N_14982,N_13400,N_12868);
nor U14983 (N_14983,N_13043,N_13340);
nor U14984 (N_14984,N_12350,N_12308);
nor U14985 (N_14985,N_12221,N_12385);
xor U14986 (N_14986,N_13270,N_12374);
nor U14987 (N_14987,N_12817,N_13321);
or U14988 (N_14988,N_12139,N_13263);
nand U14989 (N_14989,N_13416,N_13465);
and U14990 (N_14990,N_13439,N_12158);
nand U14991 (N_14991,N_13015,N_12262);
xnor U14992 (N_14992,N_12109,N_12421);
and U14993 (N_14993,N_12009,N_12615);
nor U14994 (N_14994,N_12428,N_12374);
nor U14995 (N_14995,N_12019,N_12089);
nand U14996 (N_14996,N_13283,N_13495);
xnor U14997 (N_14997,N_12733,N_12247);
and U14998 (N_14998,N_13385,N_12720);
xnor U14999 (N_14999,N_12759,N_12021);
and U15000 (N_15000,N_13729,N_13634);
nor U15001 (N_15001,N_14477,N_14917);
and U15002 (N_15002,N_14869,N_13614);
xnor U15003 (N_15003,N_13793,N_14146);
xor U15004 (N_15004,N_14778,N_14200);
xnor U15005 (N_15005,N_13609,N_13982);
and U15006 (N_15006,N_14002,N_13551);
xor U15007 (N_15007,N_14198,N_14615);
and U15008 (N_15008,N_13763,N_14057);
or U15009 (N_15009,N_13834,N_13718);
nor U15010 (N_15010,N_14991,N_13595);
or U15011 (N_15011,N_13738,N_14124);
and U15012 (N_15012,N_13954,N_13528);
or U15013 (N_15013,N_13856,N_14399);
and U15014 (N_15014,N_14192,N_14912);
and U15015 (N_15015,N_14532,N_14302);
or U15016 (N_15016,N_14375,N_14468);
xor U15017 (N_15017,N_14382,N_14098);
nand U15018 (N_15018,N_14653,N_14469);
or U15019 (N_15019,N_14233,N_14748);
or U15020 (N_15020,N_14423,N_14079);
xnor U15021 (N_15021,N_13711,N_13734);
and U15022 (N_15022,N_14516,N_14414);
or U15023 (N_15023,N_14854,N_14319);
and U15024 (N_15024,N_14901,N_14930);
xor U15025 (N_15025,N_14228,N_14520);
nand U15026 (N_15026,N_14792,N_14288);
nand U15027 (N_15027,N_14088,N_14260);
xor U15028 (N_15028,N_13893,N_13612);
nand U15029 (N_15029,N_13717,N_13749);
xor U15030 (N_15030,N_14505,N_14310);
xnor U15031 (N_15031,N_13599,N_13555);
and U15032 (N_15032,N_13603,N_14637);
nand U15033 (N_15033,N_13929,N_14305);
xor U15034 (N_15034,N_13988,N_13987);
xor U15035 (N_15035,N_13968,N_13716);
nand U15036 (N_15036,N_13650,N_14307);
xnor U15037 (N_15037,N_14551,N_13668);
and U15038 (N_15038,N_14764,N_14159);
xnor U15039 (N_15039,N_13955,N_13723);
nand U15040 (N_15040,N_14900,N_13784);
nand U15041 (N_15041,N_14841,N_13583);
nor U15042 (N_15042,N_14301,N_14056);
xor U15043 (N_15043,N_13715,N_13516);
nand U15044 (N_15044,N_14862,N_13775);
nand U15045 (N_15045,N_14938,N_13890);
and U15046 (N_15046,N_13867,N_14657);
or U15047 (N_15047,N_14689,N_14191);
nand U15048 (N_15048,N_14309,N_13624);
and U15049 (N_15049,N_13864,N_14654);
nor U15050 (N_15050,N_14485,N_14276);
xnor U15051 (N_15051,N_14958,N_14173);
or U15052 (N_15052,N_13931,N_14776);
and U15053 (N_15053,N_13602,N_14867);
nor U15054 (N_15054,N_14224,N_13917);
xor U15055 (N_15055,N_13670,N_14840);
nor U15056 (N_15056,N_13985,N_14091);
nor U15057 (N_15057,N_14422,N_14230);
and U15058 (N_15058,N_14899,N_13637);
xnor U15059 (N_15059,N_14864,N_14095);
or U15060 (N_15060,N_13753,N_14565);
xnor U15061 (N_15061,N_13582,N_14506);
or U15062 (N_15062,N_14832,N_13888);
xor U15063 (N_15063,N_14717,N_14069);
or U15064 (N_15064,N_13903,N_13740);
or U15065 (N_15065,N_13674,N_14743);
and U15066 (N_15066,N_14096,N_13689);
xor U15067 (N_15067,N_14438,N_13607);
xnor U15068 (N_15068,N_14784,N_14659);
nor U15069 (N_15069,N_14861,N_14045);
nor U15070 (N_15070,N_14221,N_14700);
and U15071 (N_15071,N_14461,N_14491);
and U15072 (N_15072,N_13735,N_13896);
nor U15073 (N_15073,N_14694,N_13511);
nor U15074 (N_15074,N_14142,N_13664);
or U15075 (N_15075,N_14464,N_14061);
xor U15076 (N_15076,N_13643,N_13894);
xor U15077 (N_15077,N_13709,N_13900);
xnor U15078 (N_15078,N_14392,N_13855);
nand U15079 (N_15079,N_13550,N_13764);
xor U15080 (N_15080,N_13733,N_14679);
and U15081 (N_15081,N_14342,N_13916);
xor U15082 (N_15082,N_13933,N_14430);
or U15083 (N_15083,N_14165,N_14686);
xnor U15084 (N_15084,N_13810,N_13536);
and U15085 (N_15085,N_13826,N_13750);
nor U15086 (N_15086,N_13564,N_14327);
or U15087 (N_15087,N_14182,N_14108);
and U15088 (N_15088,N_14160,N_14356);
nor U15089 (N_15089,N_14785,N_14406);
and U15090 (N_15090,N_13649,N_14676);
nor U15091 (N_15091,N_13849,N_13539);
or U15092 (N_15092,N_14289,N_14730);
nand U15093 (N_15093,N_14795,N_14097);
nand U15094 (N_15094,N_13660,N_14023);
and U15095 (N_15095,N_13781,N_14136);
or U15096 (N_15096,N_14408,N_13795);
and U15097 (N_15097,N_14512,N_13932);
and U15098 (N_15098,N_13658,N_13532);
nor U15099 (N_15099,N_14950,N_14021);
and U15100 (N_15100,N_14932,N_14070);
and U15101 (N_15101,N_14398,N_14454);
nor U15102 (N_15102,N_14456,N_14556);
or U15103 (N_15103,N_14740,N_14597);
xnor U15104 (N_15104,N_14533,N_14897);
or U15105 (N_15105,N_13760,N_13548);
and U15106 (N_15106,N_14129,N_14251);
and U15107 (N_15107,N_14404,N_13818);
xor U15108 (N_15108,N_14199,N_14627);
nand U15109 (N_15109,N_14280,N_13676);
xor U15110 (N_15110,N_14662,N_14985);
and U15111 (N_15111,N_14890,N_14559);
xnor U15112 (N_15112,N_14265,N_13882);
nor U15113 (N_15113,N_14871,N_13611);
and U15114 (N_15114,N_14889,N_13927);
or U15115 (N_15115,N_14314,N_14360);
or U15116 (N_15116,N_13728,N_14286);
nand U15117 (N_15117,N_14735,N_14243);
and U15118 (N_15118,N_14519,N_14384);
and U15119 (N_15119,N_14587,N_14352);
xnor U15120 (N_15120,N_13571,N_14872);
and U15121 (N_15121,N_14183,N_14621);
and U15122 (N_15122,N_14388,N_13820);
nand U15123 (N_15123,N_13765,N_14037);
xnor U15124 (N_15124,N_14853,N_14705);
nand U15125 (N_15125,N_13759,N_13581);
nand U15126 (N_15126,N_13525,N_13566);
nand U15127 (N_15127,N_14883,N_13947);
xnor U15128 (N_15128,N_13799,N_13556);
xnor U15129 (N_15129,N_14568,N_14445);
or U15130 (N_15130,N_14990,N_13881);
or U15131 (N_15131,N_13731,N_13825);
nor U15132 (N_15132,N_14790,N_14306);
xnor U15133 (N_15133,N_14172,N_14936);
nand U15134 (N_15134,N_14452,N_14364);
and U15135 (N_15135,N_14649,N_14857);
nor U15136 (N_15136,N_14378,N_14698);
xnor U15137 (N_15137,N_14143,N_14361);
nor U15138 (N_15138,N_14053,N_14294);
nand U15139 (N_15139,N_14651,N_14094);
nor U15140 (N_15140,N_13833,N_13842);
nor U15141 (N_15141,N_14726,N_14973);
nor U15142 (N_15142,N_14328,N_14955);
or U15143 (N_15143,N_13863,N_14300);
nor U15144 (N_15144,N_14333,N_14193);
or U15145 (N_15145,N_13552,N_13696);
or U15146 (N_15146,N_14610,N_13938);
or U15147 (N_15147,N_14994,N_14161);
xor U15148 (N_15148,N_13596,N_14522);
nor U15149 (N_15149,N_13802,N_14514);
nand U15150 (N_15150,N_14970,N_14104);
nor U15151 (N_15151,N_14761,N_14571);
nand U15152 (N_15152,N_13990,N_14063);
nor U15153 (N_15153,N_13590,N_14196);
or U15154 (N_15154,N_14755,N_14606);
xor U15155 (N_15155,N_14805,N_14148);
xor U15156 (N_15156,N_14455,N_14308);
nand U15157 (N_15157,N_14575,N_13514);
nor U15158 (N_15158,N_13610,N_13621);
nand U15159 (N_15159,N_14424,N_14678);
or U15160 (N_15160,N_14989,N_14670);
and U15161 (N_15161,N_13994,N_13857);
nand U15162 (N_15162,N_14020,N_13714);
xnor U15163 (N_15163,N_14187,N_14004);
and U15164 (N_15164,N_14526,N_13789);
xor U15165 (N_15165,N_14561,N_14586);
nand U15166 (N_15166,N_14368,N_13526);
nand U15167 (N_15167,N_14879,N_14636);
nand U15168 (N_15168,N_14113,N_14137);
nand U15169 (N_15169,N_14799,N_14134);
nand U15170 (N_15170,N_14335,N_13577);
nand U15171 (N_15171,N_14017,N_14708);
nor U15172 (N_15172,N_13706,N_14599);
nor U15173 (N_15173,N_14975,N_14554);
or U15174 (N_15174,N_13667,N_13541);
nor U15175 (N_15175,N_14577,N_14403);
or U15176 (N_15176,N_13817,N_14614);
xnor U15177 (N_15177,N_14434,N_13791);
or U15178 (N_15178,N_14866,N_14236);
or U15179 (N_15179,N_14838,N_13622);
xor U15180 (N_15180,N_14706,N_13724);
xnor U15181 (N_15181,N_14470,N_14696);
and U15182 (N_15182,N_13743,N_14734);
or U15183 (N_15183,N_14081,N_13854);
and U15184 (N_15184,N_14536,N_14644);
xnor U15185 (N_15185,N_14481,N_14446);
nor U15186 (N_15186,N_14849,N_13995);
xnor U15187 (N_15187,N_14812,N_14978);
nand U15188 (N_15188,N_14660,N_14727);
or U15189 (N_15189,N_14055,N_13771);
nor U15190 (N_15190,N_13895,N_14279);
and U15191 (N_15191,N_13687,N_14138);
nand U15192 (N_15192,N_14295,N_14895);
nand U15193 (N_15193,N_14839,N_14631);
nor U15194 (N_15194,N_13754,N_13673);
nor U15195 (N_15195,N_13682,N_13510);
or U15196 (N_15196,N_13695,N_14515);
xnor U15197 (N_15197,N_14436,N_13902);
nor U15198 (N_15198,N_14254,N_14664);
or U15199 (N_15199,N_14147,N_14802);
nand U15200 (N_15200,N_13892,N_14035);
or U15201 (N_15201,N_13959,N_14478);
xnor U15202 (N_15202,N_13936,N_14121);
xor U15203 (N_15203,N_14546,N_13592);
or U15204 (N_15204,N_14873,N_13549);
or U15205 (N_15205,N_13584,N_14892);
nor U15206 (N_15206,N_13942,N_14847);
nor U15207 (N_15207,N_14845,N_14639);
xor U15208 (N_15208,N_14471,N_14721);
xor U15209 (N_15209,N_13821,N_14151);
xnor U15210 (N_15210,N_14980,N_14894);
and U15211 (N_15211,N_14934,N_14229);
xor U15212 (N_15212,N_13605,N_14407);
nor U15213 (N_15213,N_14632,N_13944);
xnor U15214 (N_15214,N_13779,N_14163);
xnor U15215 (N_15215,N_13559,N_13964);
xor U15216 (N_15216,N_14579,N_14701);
or U15217 (N_15217,N_14150,N_14099);
and U15218 (N_15218,N_13647,N_14219);
or U15219 (N_15219,N_14258,N_14339);
and U15220 (N_15220,N_13688,N_14774);
or U15221 (N_15221,N_14829,N_14492);
xor U15222 (N_15222,N_13578,N_14363);
xnor U15223 (N_15223,N_14842,N_13924);
nor U15224 (N_15224,N_14034,N_14607);
nand U15225 (N_15225,N_14154,N_14806);
nand U15226 (N_15226,N_14036,N_14572);
nand U15227 (N_15227,N_14024,N_14549);
or U15228 (N_15228,N_14501,N_13980);
xor U15229 (N_15229,N_14177,N_14405);
and U15230 (N_15230,N_14139,N_14181);
nand U15231 (N_15231,N_14011,N_14888);
or U15232 (N_15232,N_13970,N_13651);
and U15233 (N_15233,N_14126,N_13846);
nor U15234 (N_15234,N_13998,N_14449);
or U15235 (N_15235,N_13946,N_14529);
or U15236 (N_15236,N_14935,N_14715);
nand U15237 (N_15237,N_13827,N_14178);
or U15238 (N_15238,N_14112,N_14072);
or U15239 (N_15239,N_13748,N_14902);
xnor U15240 (N_15240,N_14441,N_13692);
and U15241 (N_15241,N_14703,N_14331);
and U15242 (N_15242,N_13758,N_14106);
nand U15243 (N_15243,N_13652,N_14603);
nor U15244 (N_15244,N_13679,N_14860);
or U15245 (N_15245,N_13572,N_14823);
nand U15246 (N_15246,N_14028,N_14346);
xor U15247 (N_15247,N_14118,N_14428);
nand U15248 (N_15248,N_13515,N_13693);
nor U15249 (N_15249,N_13619,N_14981);
and U15250 (N_15250,N_14995,N_14006);
and U15251 (N_15251,N_14074,N_13905);
nor U15252 (N_15252,N_13604,N_13782);
nor U15253 (N_15253,N_14322,N_14227);
xor U15254 (N_15254,N_14604,N_14525);
and U15255 (N_15255,N_13989,N_13783);
nand U15256 (N_15256,N_14493,N_14809);
or U15257 (N_15257,N_14218,N_13567);
xnor U15258 (N_15258,N_13589,N_13992);
xor U15259 (N_15259,N_13770,N_13505);
nand U15260 (N_15260,N_14252,N_14366);
xor U15261 (N_15261,N_14521,N_13823);
and U15262 (N_15262,N_14680,N_14313);
xor U15263 (N_15263,N_14576,N_14672);
and U15264 (N_15264,N_14026,N_14600);
or U15265 (N_15265,N_13645,N_13865);
and U15266 (N_15266,N_14401,N_14467);
nor U15267 (N_15267,N_14073,N_14082);
nor U15268 (N_15268,N_13587,N_14462);
nand U15269 (N_15269,N_14215,N_14728);
nand U15270 (N_15270,N_14951,N_14831);
nand U15271 (N_15271,N_13869,N_14284);
nor U15272 (N_15272,N_13840,N_14810);
or U15273 (N_15273,N_14570,N_13851);
or U15274 (N_15274,N_14966,N_14263);
xnor U15275 (N_15275,N_14661,N_14292);
xor U15276 (N_15276,N_14065,N_14420);
and U15277 (N_15277,N_13755,N_14647);
nor U15278 (N_15278,N_14591,N_14330);
or U15279 (N_15279,N_13616,N_14646);
nor U15280 (N_15280,N_14350,N_13730);
nand U15281 (N_15281,N_14722,N_14933);
xnor U15282 (N_15282,N_14757,N_13701);
nor U15283 (N_15283,N_14153,N_14402);
and U15284 (N_15284,N_14231,N_14830);
nor U15285 (N_15285,N_14920,N_14624);
nor U15286 (N_15286,N_14808,N_14453);
or U15287 (N_15287,N_13935,N_13613);
nor U15288 (N_15288,N_14185,N_14396);
xnor U15289 (N_15289,N_13641,N_13597);
nor U15290 (N_15290,N_14787,N_14584);
nand U15291 (N_15291,N_13626,N_13986);
nor U15292 (N_15292,N_14737,N_14358);
nand U15293 (N_15293,N_14983,N_14690);
and U15294 (N_15294,N_14553,N_13503);
xor U15295 (N_15295,N_14960,N_14253);
xor U15296 (N_15296,N_13797,N_14495);
or U15297 (N_15297,N_14658,N_14334);
xor U15298 (N_15298,N_14448,N_14870);
xor U15299 (N_15299,N_13639,N_14859);
or U15300 (N_15300,N_14176,N_14798);
nor U15301 (N_15301,N_14131,N_14329);
or U15302 (N_15302,N_14201,N_14685);
or U15303 (N_15303,N_14896,N_14645);
nor U15304 (N_15304,N_14472,N_14796);
xnor U15305 (N_15305,N_14673,N_13521);
nor U15306 (N_15306,N_14628,N_14816);
and U15307 (N_15307,N_14391,N_14232);
or U15308 (N_15308,N_13952,N_13950);
and U15309 (N_15309,N_14166,N_14344);
xor U15310 (N_15310,N_14648,N_14054);
or U15311 (N_15311,N_13777,N_14484);
and U15312 (N_15312,N_13500,N_14527);
xor U15313 (N_15313,N_13625,N_14775);
and U15314 (N_15314,N_14238,N_14372);
nor U15315 (N_15315,N_13686,N_14101);
nand U15316 (N_15316,N_14188,N_14692);
or U15317 (N_15317,N_13966,N_14874);
or U15318 (N_15318,N_14272,N_13608);
nor U15319 (N_15319,N_13662,N_14655);
xnor U15320 (N_15320,N_14145,N_14789);
or U15321 (N_15321,N_14959,N_13948);
nor U15322 (N_15322,N_14969,N_14267);
nand U15323 (N_15323,N_14542,N_14270);
xnor U15324 (N_15324,N_14791,N_14915);
and U15325 (N_15325,N_13756,N_14601);
xor U15326 (N_15326,N_14751,N_14777);
nand U15327 (N_15327,N_14713,N_14943);
xnor U15328 (N_15328,N_14049,N_14788);
and U15329 (N_15329,N_14547,N_13772);
nor U15330 (N_15330,N_13681,N_13690);
nor U15331 (N_15331,N_14819,N_14758);
nand U15332 (N_15332,N_14204,N_14050);
nor U15333 (N_15333,N_14007,N_14793);
and U15334 (N_15334,N_14911,N_14080);
or U15335 (N_15335,N_14630,N_13832);
and U15336 (N_15336,N_14089,N_14588);
nor U15337 (N_15337,N_13553,N_14910);
or U15338 (N_15338,N_14103,N_13787);
or U15339 (N_15339,N_13803,N_13830);
and U15340 (N_15340,N_14189,N_14589);
nor U15341 (N_15341,N_14596,N_13722);
xor U15342 (N_15342,N_13909,N_14602);
xnor U15343 (N_15343,N_14765,N_14773);
xnor U15344 (N_15344,N_14325,N_14693);
xnor U15345 (N_15345,N_14827,N_14675);
and U15346 (N_15346,N_14535,N_14040);
nand U15347 (N_15347,N_14687,N_14707);
or U15348 (N_15348,N_14937,N_13545);
xnor U15349 (N_15349,N_14038,N_13628);
nand U15350 (N_15350,N_13940,N_14821);
and U15351 (N_15351,N_14197,N_13638);
nor U15352 (N_15352,N_14848,N_14837);
nand U15353 (N_15353,N_14507,N_14371);
or U15354 (N_15354,N_13860,N_13742);
or U15355 (N_15355,N_14993,N_13691);
nor U15356 (N_15356,N_14179,N_13801);
nand U15357 (N_15357,N_14413,N_13920);
nor U15358 (N_15358,N_13725,N_13642);
or U15359 (N_15359,N_13565,N_14987);
and U15360 (N_15360,N_13848,N_14580);
nand U15361 (N_15361,N_14184,N_13809);
nor U15362 (N_15362,N_13540,N_14212);
and U15363 (N_15363,N_14931,N_14421);
or U15364 (N_15364,N_14504,N_13757);
and U15365 (N_15365,N_14092,N_14563);
nor U15366 (N_15366,N_13977,N_14926);
nand U15367 (N_15367,N_14068,N_13873);
nand U15368 (N_15368,N_13862,N_13804);
or U15369 (N_15369,N_13533,N_14362);
nor U15370 (N_15370,N_14583,N_14030);
and U15371 (N_15371,N_14043,N_13618);
nand U15372 (N_15372,N_13535,N_14724);
nand U15373 (N_15373,N_14474,N_14473);
xor U15374 (N_15374,N_14451,N_14817);
xnor U15375 (N_15375,N_14419,N_14475);
or U15376 (N_15376,N_14303,N_14248);
nand U15377 (N_15377,N_13623,N_13847);
or U15378 (N_15378,N_13767,N_14127);
and U15379 (N_15379,N_14115,N_14585);
xnor U15380 (N_15380,N_14875,N_14427);
or U15381 (N_15381,N_13704,N_14534);
nor U15382 (N_15382,N_14105,N_14711);
or U15383 (N_15383,N_14818,N_14483);
xnor U15384 (N_15384,N_14369,N_14290);
nor U15385 (N_15385,N_13575,N_13560);
and U15386 (N_15386,N_13635,N_14415);
and U15387 (N_15387,N_14768,N_14738);
nand U15388 (N_15388,N_14626,N_13737);
and U15389 (N_15389,N_13684,N_13877);
xor U15390 (N_15390,N_14465,N_14394);
nand U15391 (N_15391,N_14444,N_13680);
and U15392 (N_15392,N_14545,N_14919);
xor U15393 (N_15393,N_14435,N_14064);
or U15394 (N_15394,N_14235,N_14928);
nand U15395 (N_15395,N_13844,N_13726);
and U15396 (N_15396,N_14623,N_13698);
nor U15397 (N_15397,N_14479,N_14552);
xnor U15398 (N_15398,N_13627,N_14843);
or U15399 (N_15399,N_13752,N_14638);
nand U15400 (N_15400,N_14425,N_14059);
and U15401 (N_15401,N_13914,N_14117);
nand U15402 (N_15402,N_13963,N_14353);
and U15403 (N_15403,N_14225,N_13972);
nor U15404 (N_15404,N_14858,N_14929);
nand U15405 (N_15405,N_14923,N_14813);
nor U15406 (N_15406,N_13591,N_13800);
and U15407 (N_15407,N_14149,N_14834);
nand U15408 (N_15408,N_14365,N_14865);
nor U15409 (N_15409,N_13538,N_13746);
and U15410 (N_15410,N_14760,N_14119);
xnor U15411 (N_15411,N_13710,N_14367);
nand U15412 (N_15412,N_14801,N_14027);
and U15413 (N_15413,N_14523,N_13594);
or U15414 (N_15414,N_14195,N_13871);
or U15415 (N_15415,N_14605,N_13805);
or U15416 (N_15416,N_14291,N_14123);
nand U15417 (N_15417,N_14982,N_14262);
xnor U15418 (N_15418,N_14110,N_14544);
xor U15419 (N_15419,N_14264,N_14732);
or U15420 (N_15420,N_13557,N_14835);
nand U15421 (N_15421,N_13798,N_13580);
nand U15422 (N_15422,N_13501,N_13837);
nand U15423 (N_15423,N_13786,N_14752);
or U15424 (N_15424,N_14964,N_14348);
nand U15425 (N_15425,N_14921,N_14271);
nand U15426 (N_15426,N_14261,N_13831);
xor U15427 (N_15427,N_13901,N_14749);
nor U15428 (N_15428,N_14487,N_14001);
or U15429 (N_15429,N_14744,N_14736);
or U15430 (N_15430,N_13700,N_14885);
or U15431 (N_15431,N_14868,N_14574);
and U15432 (N_15432,N_14620,N_14642);
xnor U15433 (N_15433,N_14725,N_14255);
or U15434 (N_15434,N_14343,N_14754);
nor U15435 (N_15435,N_14640,N_14712);
nor U15436 (N_15436,N_14132,N_13960);
nor U15437 (N_15437,N_13945,N_13744);
or U15438 (N_15438,N_14663,N_13984);
or U15439 (N_15439,N_14100,N_14380);
nor U15440 (N_15440,N_13579,N_14560);
xnor U15441 (N_15441,N_14731,N_14439);
or U15442 (N_15442,N_13979,N_14742);
nor U15443 (N_15443,N_14668,N_13928);
nor U15444 (N_15444,N_14312,N_14087);
nand U15445 (N_15445,N_14741,N_14220);
and U15446 (N_15446,N_14245,N_14440);
nor U15447 (N_15447,N_13675,N_13762);
or U15448 (N_15448,N_13876,N_14476);
nor U15449 (N_15449,N_14277,N_14315);
nand U15450 (N_15450,N_14332,N_14498);
xnor U15451 (N_15451,N_14511,N_13769);
and U15452 (N_15452,N_14852,N_14695);
nor U15453 (N_15453,N_14275,N_14846);
and U15454 (N_15454,N_14450,N_14223);
nand U15455 (N_15455,N_14746,N_14499);
nand U15456 (N_15456,N_13586,N_13712);
nand U15457 (N_15457,N_14674,N_13570);
nor U15458 (N_15458,N_13736,N_14268);
and U15459 (N_15459,N_14433,N_13519);
and U15460 (N_15460,N_14359,N_14769);
xnor U15461 (N_15461,N_14633,N_14617);
nand U15462 (N_15462,N_13739,N_14397);
xor U15463 (N_15463,N_14939,N_14076);
xnor U15464 (N_15464,N_14878,N_14999);
nor U15465 (N_15465,N_13546,N_14759);
nand U15466 (N_15466,N_14581,N_13671);
xnor U15467 (N_15467,N_13513,N_13918);
nor U15468 (N_15468,N_14242,N_14257);
xor U15469 (N_15469,N_14297,N_14052);
and U15470 (N_15470,N_13962,N_13907);
and U15471 (N_15471,N_14259,N_14984);
nor U15472 (N_15472,N_13665,N_14656);
nand U15473 (N_15473,N_14084,N_13631);
nand U15474 (N_15474,N_14977,N_13646);
or U15475 (N_15475,N_14318,N_13983);
nor U15476 (N_15476,N_14000,N_14357);
or U15477 (N_15477,N_14800,N_14085);
nor U15478 (N_15478,N_14032,N_13796);
xor U15479 (N_15479,N_14285,N_13785);
xor U15480 (N_15480,N_14273,N_13657);
nand U15481 (N_15481,N_14202,N_14164);
nor U15482 (N_15482,N_14767,N_14347);
nor U15483 (N_15483,N_13926,N_14460);
nor U15484 (N_15484,N_14590,N_14437);
or U15485 (N_15485,N_14756,N_14083);
xnor U15486 (N_15486,N_14611,N_13841);
nor U15487 (N_15487,N_13884,N_14609);
and U15488 (N_15488,N_14381,N_14836);
xor U15489 (N_15489,N_14207,N_13845);
or U15490 (N_15490,N_13792,N_14906);
nand U15491 (N_15491,N_14412,N_14458);
and U15492 (N_15492,N_14893,N_14826);
nand U15493 (N_15493,N_14152,N_14377);
nand U15494 (N_15494,N_14947,N_14781);
nand U15495 (N_15495,N_14005,N_13562);
nor U15496 (N_15496,N_14033,N_14247);
xnor U15497 (N_15497,N_13527,N_13694);
or U15498 (N_15498,N_14316,N_13858);
or U15499 (N_15499,N_14107,N_13617);
xor U15500 (N_15500,N_14772,N_14718);
nand U15501 (N_15501,N_13741,N_13886);
nand U15502 (N_15502,N_13534,N_13835);
and U15503 (N_15503,N_14688,N_14321);
nand U15504 (N_15504,N_14822,N_14903);
and U15505 (N_15505,N_13653,N_14913);
and U15506 (N_15506,N_14887,N_14691);
xnor U15507 (N_15507,N_13520,N_13941);
and U15508 (N_15508,N_14595,N_14907);
nand U15509 (N_15509,N_13878,N_13910);
or U15510 (N_15510,N_13975,N_14952);
and U15511 (N_15511,N_14962,N_13922);
and U15512 (N_15512,N_14447,N_14416);
nor U15513 (N_15513,N_14763,N_13707);
and U15514 (N_15514,N_13951,N_14237);
nor U15515 (N_15515,N_13518,N_14042);
and U15516 (N_15516,N_14109,N_13504);
and U15517 (N_15517,N_14953,N_13713);
nor U15518 (N_15518,N_14783,N_14022);
and U15519 (N_15519,N_13554,N_14592);
xor U15520 (N_15520,N_14634,N_13685);
xnor U15521 (N_15521,N_14945,N_14528);
nor U15522 (N_15522,N_14048,N_14373);
nor U15523 (N_15523,N_14029,N_13719);
and U15524 (N_15524,N_13766,N_14569);
nor U15525 (N_15525,N_14010,N_13879);
nand U15526 (N_15526,N_14374,N_13531);
nor U15527 (N_15527,N_13891,N_13828);
nor U15528 (N_15528,N_13861,N_14567);
and U15529 (N_15529,N_14666,N_13666);
xnor U15530 (N_15530,N_14782,N_13981);
nand U15531 (N_15531,N_14619,N_14881);
or U15532 (N_15532,N_14217,N_14954);
nor U15533 (N_15533,N_13507,N_14283);
xnor U15534 (N_15534,N_14250,N_14431);
and U15535 (N_15535,N_14530,N_13997);
nor U15536 (N_15536,N_14208,N_13522);
or U15537 (N_15537,N_13558,N_13898);
nand U15538 (N_15538,N_13508,N_14779);
and U15539 (N_15539,N_14612,N_13561);
or U15540 (N_15540,N_14747,N_14786);
or U15541 (N_15541,N_14824,N_14988);
and U15542 (N_15542,N_14909,N_13773);
nor U15543 (N_15543,N_14976,N_13829);
nand U15544 (N_15544,N_14086,N_14961);
or U15545 (N_15545,N_14019,N_14209);
nor U15546 (N_15546,N_13868,N_14650);
nor U15547 (N_15547,N_13976,N_13655);
nand U15548 (N_15548,N_14269,N_14974);
xnor U15549 (N_15549,N_14256,N_14041);
xor U15550 (N_15550,N_14298,N_14968);
nor U15551 (N_15551,N_13836,N_14524);
nor U15552 (N_15552,N_13925,N_13957);
nand U15553 (N_15553,N_14697,N_13768);
xnor U15554 (N_15554,N_14635,N_13529);
xnor U15555 (N_15555,N_14426,N_13958);
nor U15556 (N_15556,N_13678,N_14457);
nor U15557 (N_15557,N_14877,N_13672);
or U15558 (N_15558,N_13996,N_14213);
xnor U15559 (N_15559,N_14510,N_13794);
nand U15560 (N_15560,N_13661,N_14488);
xnor U15561 (N_15561,N_14598,N_13588);
xnor U15562 (N_15562,N_14067,N_14039);
or U15563 (N_15563,N_13654,N_13934);
or U15564 (N_15564,N_14157,N_13636);
nand U15565 (N_15565,N_14677,N_14558);
nand U15566 (N_15566,N_14665,N_13509);
nand U15567 (N_15567,N_14946,N_13852);
or U15568 (N_15568,N_14417,N_13887);
xor U15569 (N_15569,N_14031,N_14682);
nor U15570 (N_15570,N_14003,N_14803);
and U15571 (N_15571,N_13912,N_14180);
nand U15572 (N_15572,N_14739,N_13923);
nand U15573 (N_15573,N_13648,N_14905);
nand U15574 (N_15574,N_14513,N_14497);
nor U15575 (N_15575,N_13573,N_14863);
nor U15576 (N_15576,N_14214,N_13967);
xnor U15577 (N_15577,N_13523,N_14616);
xor U15578 (N_15578,N_14443,N_14766);
and U15579 (N_15579,N_13727,N_14750);
xnor U15580 (N_15580,N_14745,N_14564);
nor U15581 (N_15581,N_13904,N_13745);
or U15582 (N_15582,N_13524,N_14156);
nand U15583 (N_15583,N_14720,N_14876);
or U15584 (N_15584,N_14855,N_14386);
and U15585 (N_15585,N_14566,N_14170);
nor U15586 (N_15586,N_13897,N_14194);
or U15587 (N_15587,N_13872,N_14578);
xnor U15588 (N_15588,N_13574,N_13517);
xnor U15589 (N_15589,N_14016,N_14916);
nor U15590 (N_15590,N_14770,N_13838);
nor U15591 (N_15591,N_14379,N_14389);
or U15592 (N_15592,N_14797,N_13542);
xnor U15593 (N_15593,N_14130,N_13512);
xor U15594 (N_15594,N_13973,N_13859);
xor U15595 (N_15595,N_14013,N_14942);
and U15596 (N_15596,N_14502,N_14794);
nor U15597 (N_15597,N_13790,N_13993);
nor U15598 (N_15598,N_13953,N_13883);
or U15599 (N_15599,N_14376,N_13811);
xnor U15600 (N_15600,N_13816,N_14851);
nand U15601 (N_15601,N_14608,N_14486);
nand U15602 (N_15602,N_14992,N_14186);
nand U15603 (N_15603,N_13915,N_14856);
nor U15604 (N_15604,N_14667,N_14941);
nor U15605 (N_15605,N_14008,N_14044);
xnor U15606 (N_15606,N_14466,N_13999);
or U15607 (N_15607,N_14296,N_14540);
and U15608 (N_15608,N_14886,N_14282);
xor U15609 (N_15609,N_13969,N_14062);
xnor U15610 (N_15610,N_13620,N_14222);
nor U15611 (N_15611,N_14326,N_13808);
xnor U15612 (N_15612,N_13850,N_14494);
and U15613 (N_15613,N_14811,N_13813);
xor U15614 (N_15614,N_14249,N_14411);
or U15615 (N_15615,N_14979,N_14908);
nand U15616 (N_15616,N_14239,N_13815);
or U15617 (N_15617,N_14128,N_14996);
or U15618 (N_15618,N_13822,N_14924);
or U15619 (N_15619,N_14395,N_13606);
nand U15620 (N_15620,N_13615,N_14241);
xnor U15621 (N_15621,N_14240,N_14090);
or U15622 (N_15622,N_14354,N_14683);
nand U15623 (N_15623,N_13839,N_14557);
or U15624 (N_15624,N_14771,N_13965);
xor U15625 (N_15625,N_13544,N_14463);
xor U15626 (N_15626,N_14226,N_14216);
xor U15627 (N_15627,N_14393,N_14336);
nand U15628 (N_15628,N_13576,N_13978);
nand U15629 (N_15629,N_14370,N_14046);
or U15630 (N_15630,N_14681,N_14009);
and U15631 (N_15631,N_13563,N_13502);
or U15632 (N_15632,N_14957,N_13761);
or U15633 (N_15633,N_14060,N_14555);
xnor U15634 (N_15634,N_14317,N_14211);
nand U15635 (N_15635,N_14135,N_13683);
or U15636 (N_15636,N_14387,N_13908);
or U15637 (N_15637,N_14815,N_14629);
and U15638 (N_15638,N_13547,N_14490);
nor U15639 (N_15639,N_14704,N_14116);
and U15640 (N_15640,N_14078,N_14714);
or U15641 (N_15641,N_14918,N_13956);
xnor U15642 (N_15642,N_13824,N_14710);
and U15643 (N_15643,N_14355,N_14496);
or U15644 (N_15644,N_13598,N_14833);
nand U15645 (N_15645,N_14169,N_13780);
or U15646 (N_15646,N_14550,N_14168);
nor U15647 (N_15647,N_14593,N_13921);
nand U15648 (N_15648,N_14158,N_13677);
nor U15649 (N_15649,N_14120,N_14543);
or U15650 (N_15650,N_13778,N_14442);
nor U15651 (N_15651,N_13885,N_14927);
nand U15652 (N_15652,N_14641,N_14963);
and U15653 (N_15653,N_13656,N_14155);
or U15654 (N_15654,N_14716,N_13663);
and U15655 (N_15655,N_14102,N_14025);
or U15656 (N_15656,N_14986,N_14274);
xnor U15657 (N_15657,N_13939,N_14266);
xor U15658 (N_15658,N_13600,N_14538);
nand U15659 (N_15659,N_14015,N_14093);
nand U15660 (N_15660,N_13880,N_14014);
and U15661 (N_15661,N_14531,N_14828);
or U15662 (N_15662,N_14548,N_13991);
nand U15663 (N_15663,N_14998,N_14537);
nor U15664 (N_15664,N_14884,N_14825);
nand U15665 (N_15665,N_13974,N_14904);
or U15666 (N_15666,N_13788,N_14669);
nand U15667 (N_15667,N_14345,N_14971);
or U15668 (N_15668,N_14012,N_14234);
xor U15669 (N_15669,N_13543,N_14482);
xnor U15670 (N_15670,N_14489,N_14429);
nor U15671 (N_15671,N_13568,N_13630);
or U15672 (N_15672,N_14807,N_14071);
and U15673 (N_15673,N_14293,N_14432);
nand U15674 (N_15674,N_14949,N_13506);
xor U15675 (N_15675,N_13774,N_14622);
nand U15676 (N_15676,N_14400,N_14652);
or U15677 (N_15677,N_13569,N_14337);
or U15678 (N_15678,N_14925,N_13593);
and U15679 (N_15679,N_14162,N_14144);
or U15680 (N_15680,N_14594,N_14018);
xor U15681 (N_15681,N_14205,N_14965);
nand U15682 (N_15682,N_13530,N_14287);
nand U15683 (N_15683,N_13632,N_13919);
xnor U15684 (N_15684,N_14844,N_14340);
xnor U15685 (N_15685,N_14804,N_13721);
nor U15686 (N_15686,N_14780,N_13697);
nand U15687 (N_15687,N_14410,N_13819);
nand U15688 (N_15688,N_14509,N_14114);
and U15689 (N_15689,N_14244,N_13870);
and U15690 (N_15690,N_13708,N_14891);
xnor U15691 (N_15691,N_13937,N_14541);
or U15692 (N_15692,N_14324,N_14210);
or U15693 (N_15693,N_14281,N_13812);
nand U15694 (N_15694,N_14967,N_14304);
nor U15695 (N_15695,N_14753,N_13702);
or U15696 (N_15696,N_13659,N_13889);
and U15697 (N_15697,N_13906,N_14699);
and U15698 (N_15698,N_14539,N_14880);
nor U15699 (N_15699,N_13629,N_14206);
nand U15700 (N_15700,N_14122,N_13776);
nand U15701 (N_15701,N_14850,N_14517);
and U15702 (N_15702,N_13911,N_13806);
xor U15703 (N_15703,N_14323,N_13913);
and U15704 (N_15704,N_13537,N_13703);
nor U15705 (N_15705,N_14643,N_14503);
or U15706 (N_15706,N_14625,N_13961);
or U15707 (N_15707,N_14141,N_14882);
xor U15708 (N_15708,N_14723,N_14203);
or U15709 (N_15709,N_14500,N_14278);
nor U15710 (N_15710,N_14047,N_14684);
or U15711 (N_15711,N_14671,N_14898);
and U15712 (N_15712,N_14075,N_14762);
xor U15713 (N_15713,N_14733,N_14058);
and U15714 (N_15714,N_14190,N_14175);
nor U15715 (N_15715,N_14922,N_14338);
xnor U15716 (N_15716,N_13640,N_13949);
or U15717 (N_15717,N_14729,N_14351);
nor U15718 (N_15718,N_14167,N_14562);
or U15719 (N_15719,N_14480,N_14944);
nor U15720 (N_15720,N_14618,N_14997);
and U15721 (N_15721,N_14582,N_14418);
nand U15722 (N_15722,N_13585,N_14940);
and U15723 (N_15723,N_14914,N_14066);
or U15724 (N_15724,N_14349,N_13601);
nand U15725 (N_15725,N_13866,N_13875);
and U15726 (N_15726,N_14133,N_14383);
and U15727 (N_15727,N_14508,N_13843);
nor U15728 (N_15728,N_14171,N_13732);
nor U15729 (N_15729,N_14409,N_14299);
xor U15730 (N_15730,N_13720,N_14174);
and U15731 (N_15731,N_13930,N_13751);
and U15732 (N_15732,N_14311,N_14459);
or U15733 (N_15733,N_13699,N_13669);
and U15734 (N_15734,N_13899,N_14709);
xor U15735 (N_15735,N_14246,N_14814);
xor U15736 (N_15736,N_14613,N_14390);
nor U15737 (N_15737,N_14125,N_13943);
and U15738 (N_15738,N_14956,N_14820);
and U15739 (N_15739,N_14341,N_14719);
xnor U15740 (N_15740,N_14518,N_13747);
or U15741 (N_15741,N_14111,N_13705);
nor U15742 (N_15742,N_13971,N_13807);
nand U15743 (N_15743,N_14385,N_14702);
or U15744 (N_15744,N_13644,N_13814);
xor U15745 (N_15745,N_14573,N_13874);
xnor U15746 (N_15746,N_14948,N_14051);
nand U15747 (N_15747,N_14140,N_13853);
nand U15748 (N_15748,N_14077,N_14320);
or U15749 (N_15749,N_14972,N_13633);
nor U15750 (N_15750,N_14528,N_13953);
and U15751 (N_15751,N_14427,N_13928);
nor U15752 (N_15752,N_14651,N_14322);
nor U15753 (N_15753,N_14546,N_14402);
nand U15754 (N_15754,N_14179,N_13510);
nand U15755 (N_15755,N_14303,N_14280);
xnor U15756 (N_15756,N_14214,N_14342);
and U15757 (N_15757,N_14694,N_13838);
or U15758 (N_15758,N_14026,N_14704);
or U15759 (N_15759,N_14967,N_14002);
nor U15760 (N_15760,N_13740,N_14963);
xnor U15761 (N_15761,N_14635,N_14242);
and U15762 (N_15762,N_14752,N_14291);
and U15763 (N_15763,N_14628,N_14663);
xor U15764 (N_15764,N_13626,N_13848);
or U15765 (N_15765,N_14832,N_14988);
and U15766 (N_15766,N_14185,N_13949);
nor U15767 (N_15767,N_14178,N_14080);
nand U15768 (N_15768,N_14478,N_14409);
xor U15769 (N_15769,N_14231,N_13966);
xnor U15770 (N_15770,N_13855,N_13884);
and U15771 (N_15771,N_14141,N_14633);
nand U15772 (N_15772,N_14664,N_14353);
xnor U15773 (N_15773,N_13844,N_13608);
or U15774 (N_15774,N_14375,N_13556);
or U15775 (N_15775,N_13561,N_14232);
and U15776 (N_15776,N_14467,N_13974);
and U15777 (N_15777,N_13843,N_14273);
and U15778 (N_15778,N_13654,N_13748);
xor U15779 (N_15779,N_14120,N_14080);
xor U15780 (N_15780,N_14664,N_14156);
or U15781 (N_15781,N_14677,N_14369);
and U15782 (N_15782,N_14703,N_14983);
xor U15783 (N_15783,N_14251,N_13509);
nand U15784 (N_15784,N_14748,N_14421);
and U15785 (N_15785,N_14193,N_13778);
nor U15786 (N_15786,N_14107,N_14768);
nand U15787 (N_15787,N_14935,N_14824);
nand U15788 (N_15788,N_14031,N_14034);
nand U15789 (N_15789,N_14115,N_13945);
nor U15790 (N_15790,N_13709,N_13633);
or U15791 (N_15791,N_14464,N_14102);
or U15792 (N_15792,N_14209,N_14905);
nor U15793 (N_15793,N_13925,N_14670);
or U15794 (N_15794,N_13893,N_13716);
nor U15795 (N_15795,N_14270,N_14242);
nor U15796 (N_15796,N_14353,N_13918);
nand U15797 (N_15797,N_14271,N_13971);
nor U15798 (N_15798,N_14920,N_13543);
xor U15799 (N_15799,N_14977,N_14606);
nand U15800 (N_15800,N_14529,N_14156);
nand U15801 (N_15801,N_13824,N_14575);
nor U15802 (N_15802,N_13706,N_14284);
or U15803 (N_15803,N_13538,N_13939);
or U15804 (N_15804,N_14575,N_14715);
nor U15805 (N_15805,N_14153,N_13504);
nand U15806 (N_15806,N_14064,N_13880);
and U15807 (N_15807,N_13601,N_14022);
nor U15808 (N_15808,N_14230,N_13825);
xor U15809 (N_15809,N_14275,N_14714);
or U15810 (N_15810,N_14334,N_14849);
nand U15811 (N_15811,N_14571,N_14073);
or U15812 (N_15812,N_14414,N_14439);
xor U15813 (N_15813,N_14728,N_14853);
nand U15814 (N_15814,N_14940,N_13614);
nand U15815 (N_15815,N_13714,N_13746);
nand U15816 (N_15816,N_14332,N_14279);
or U15817 (N_15817,N_14217,N_14517);
xor U15818 (N_15818,N_13709,N_13534);
and U15819 (N_15819,N_13943,N_14301);
or U15820 (N_15820,N_14696,N_13923);
and U15821 (N_15821,N_13554,N_13957);
nand U15822 (N_15822,N_13785,N_13922);
xnor U15823 (N_15823,N_14532,N_14085);
xor U15824 (N_15824,N_14159,N_14222);
and U15825 (N_15825,N_14121,N_14778);
xor U15826 (N_15826,N_13882,N_14294);
xor U15827 (N_15827,N_13870,N_14216);
xor U15828 (N_15828,N_14180,N_14057);
nand U15829 (N_15829,N_13652,N_14756);
and U15830 (N_15830,N_14487,N_14579);
and U15831 (N_15831,N_14667,N_14799);
nor U15832 (N_15832,N_13718,N_13758);
xor U15833 (N_15833,N_14092,N_13793);
or U15834 (N_15834,N_14144,N_14709);
nand U15835 (N_15835,N_14166,N_14940);
or U15836 (N_15836,N_14800,N_14896);
and U15837 (N_15837,N_13757,N_14640);
nand U15838 (N_15838,N_14296,N_14736);
xnor U15839 (N_15839,N_13785,N_13792);
or U15840 (N_15840,N_13603,N_13683);
nand U15841 (N_15841,N_14048,N_13855);
or U15842 (N_15842,N_14069,N_14203);
nor U15843 (N_15843,N_14181,N_14596);
nor U15844 (N_15844,N_14576,N_14887);
nor U15845 (N_15845,N_14533,N_14890);
nor U15846 (N_15846,N_14484,N_14183);
xnor U15847 (N_15847,N_14923,N_13795);
or U15848 (N_15848,N_14410,N_13588);
xnor U15849 (N_15849,N_13696,N_14816);
xor U15850 (N_15850,N_13745,N_13900);
or U15851 (N_15851,N_14267,N_14466);
xnor U15852 (N_15852,N_14702,N_14236);
or U15853 (N_15853,N_14578,N_13602);
xor U15854 (N_15854,N_14771,N_14702);
nor U15855 (N_15855,N_14948,N_14311);
nand U15856 (N_15856,N_14004,N_13683);
xor U15857 (N_15857,N_14406,N_13819);
or U15858 (N_15858,N_14730,N_14885);
and U15859 (N_15859,N_14994,N_13962);
and U15860 (N_15860,N_13843,N_14694);
xnor U15861 (N_15861,N_14358,N_13521);
or U15862 (N_15862,N_13889,N_13767);
or U15863 (N_15863,N_13805,N_14465);
and U15864 (N_15864,N_13800,N_14263);
nor U15865 (N_15865,N_13882,N_13838);
and U15866 (N_15866,N_13762,N_14500);
or U15867 (N_15867,N_13637,N_14325);
or U15868 (N_15868,N_14382,N_14533);
nor U15869 (N_15869,N_13935,N_13595);
and U15870 (N_15870,N_14952,N_14825);
and U15871 (N_15871,N_14848,N_14249);
or U15872 (N_15872,N_13593,N_14993);
or U15873 (N_15873,N_14138,N_14855);
nand U15874 (N_15874,N_13967,N_14020);
nor U15875 (N_15875,N_13776,N_14520);
and U15876 (N_15876,N_14583,N_13968);
nand U15877 (N_15877,N_13650,N_14406);
nor U15878 (N_15878,N_14206,N_13881);
or U15879 (N_15879,N_14325,N_13539);
and U15880 (N_15880,N_14536,N_14917);
or U15881 (N_15881,N_14586,N_13955);
nand U15882 (N_15882,N_13945,N_14701);
or U15883 (N_15883,N_14751,N_13976);
xnor U15884 (N_15884,N_14760,N_14073);
nor U15885 (N_15885,N_13941,N_14665);
xor U15886 (N_15886,N_14807,N_14635);
nand U15887 (N_15887,N_14979,N_14889);
xor U15888 (N_15888,N_14782,N_13984);
and U15889 (N_15889,N_14581,N_14574);
or U15890 (N_15890,N_13558,N_14989);
or U15891 (N_15891,N_13554,N_14470);
xnor U15892 (N_15892,N_13864,N_14270);
and U15893 (N_15893,N_13881,N_14874);
nor U15894 (N_15894,N_13961,N_14247);
nor U15895 (N_15895,N_14726,N_14051);
and U15896 (N_15896,N_14633,N_13745);
nor U15897 (N_15897,N_13746,N_13718);
or U15898 (N_15898,N_14139,N_14122);
xnor U15899 (N_15899,N_14666,N_14635);
or U15900 (N_15900,N_14990,N_14045);
nor U15901 (N_15901,N_14336,N_14734);
or U15902 (N_15902,N_14917,N_13844);
nand U15903 (N_15903,N_13748,N_14141);
nand U15904 (N_15904,N_14715,N_13974);
or U15905 (N_15905,N_14787,N_14487);
nand U15906 (N_15906,N_14346,N_13690);
nor U15907 (N_15907,N_14428,N_13681);
or U15908 (N_15908,N_13576,N_13844);
nand U15909 (N_15909,N_13683,N_14339);
or U15910 (N_15910,N_13821,N_14131);
xor U15911 (N_15911,N_14689,N_14658);
or U15912 (N_15912,N_13727,N_14582);
xor U15913 (N_15913,N_14757,N_14373);
xnor U15914 (N_15914,N_14671,N_14769);
nor U15915 (N_15915,N_14587,N_13928);
or U15916 (N_15916,N_14292,N_13937);
nor U15917 (N_15917,N_13979,N_13903);
or U15918 (N_15918,N_13569,N_14843);
and U15919 (N_15919,N_13814,N_14982);
xor U15920 (N_15920,N_14391,N_13955);
nand U15921 (N_15921,N_14029,N_14376);
or U15922 (N_15922,N_13810,N_14701);
or U15923 (N_15923,N_13583,N_14077);
nor U15924 (N_15924,N_14700,N_14845);
xnor U15925 (N_15925,N_14868,N_13989);
nand U15926 (N_15926,N_13743,N_14756);
nand U15927 (N_15927,N_14985,N_14497);
nand U15928 (N_15928,N_14928,N_14312);
xor U15929 (N_15929,N_13679,N_14748);
nor U15930 (N_15930,N_13631,N_14882);
xor U15931 (N_15931,N_14113,N_13704);
nand U15932 (N_15932,N_13820,N_13688);
and U15933 (N_15933,N_13916,N_13886);
nand U15934 (N_15934,N_13865,N_14189);
xor U15935 (N_15935,N_14465,N_14212);
nand U15936 (N_15936,N_14275,N_13849);
xor U15937 (N_15937,N_13585,N_14395);
nand U15938 (N_15938,N_13883,N_13631);
nor U15939 (N_15939,N_14902,N_13839);
or U15940 (N_15940,N_13834,N_14009);
nor U15941 (N_15941,N_14701,N_14867);
nand U15942 (N_15942,N_13867,N_14691);
and U15943 (N_15943,N_14250,N_14050);
or U15944 (N_15944,N_14128,N_14716);
xor U15945 (N_15945,N_14627,N_13991);
nand U15946 (N_15946,N_14968,N_14922);
or U15947 (N_15947,N_14586,N_14628);
and U15948 (N_15948,N_14879,N_14720);
and U15949 (N_15949,N_13640,N_13521);
nand U15950 (N_15950,N_14903,N_13538);
and U15951 (N_15951,N_14792,N_14305);
or U15952 (N_15952,N_14758,N_14672);
nor U15953 (N_15953,N_14888,N_13676);
xnor U15954 (N_15954,N_13532,N_14307);
or U15955 (N_15955,N_13539,N_13946);
and U15956 (N_15956,N_14508,N_14070);
and U15957 (N_15957,N_14424,N_14326);
and U15958 (N_15958,N_14773,N_14757);
nor U15959 (N_15959,N_14868,N_13991);
and U15960 (N_15960,N_14311,N_14355);
nor U15961 (N_15961,N_14261,N_13601);
xor U15962 (N_15962,N_13683,N_13698);
nand U15963 (N_15963,N_14483,N_14303);
nor U15964 (N_15964,N_14918,N_13713);
and U15965 (N_15965,N_14913,N_13782);
or U15966 (N_15966,N_14305,N_13643);
nand U15967 (N_15967,N_13694,N_14326);
nand U15968 (N_15968,N_14966,N_14643);
and U15969 (N_15969,N_14654,N_14159);
and U15970 (N_15970,N_14478,N_14252);
nor U15971 (N_15971,N_14999,N_14957);
nand U15972 (N_15972,N_14103,N_14142);
nor U15973 (N_15973,N_14712,N_14503);
xor U15974 (N_15974,N_13746,N_14816);
nor U15975 (N_15975,N_13771,N_13742);
and U15976 (N_15976,N_13697,N_14716);
nand U15977 (N_15977,N_14845,N_13920);
xor U15978 (N_15978,N_14388,N_14343);
and U15979 (N_15979,N_14295,N_13958);
nor U15980 (N_15980,N_14848,N_14445);
or U15981 (N_15981,N_14641,N_13717);
nor U15982 (N_15982,N_14858,N_13913);
and U15983 (N_15983,N_13715,N_13955);
nand U15984 (N_15984,N_14524,N_14689);
and U15985 (N_15985,N_14436,N_13885);
nand U15986 (N_15986,N_13805,N_14003);
nand U15987 (N_15987,N_13995,N_13817);
nor U15988 (N_15988,N_14442,N_14053);
xnor U15989 (N_15989,N_14908,N_14584);
or U15990 (N_15990,N_14207,N_13744);
or U15991 (N_15991,N_13603,N_13921);
xnor U15992 (N_15992,N_14339,N_14696);
and U15993 (N_15993,N_14520,N_14080);
nor U15994 (N_15994,N_14262,N_13593);
nor U15995 (N_15995,N_13656,N_14918);
xnor U15996 (N_15996,N_14411,N_13683);
and U15997 (N_15997,N_14447,N_13887);
nor U15998 (N_15998,N_13881,N_14706);
or U15999 (N_15999,N_13787,N_14430);
xor U16000 (N_16000,N_13922,N_14019);
xnor U16001 (N_16001,N_14052,N_13531);
nand U16002 (N_16002,N_13975,N_14472);
nor U16003 (N_16003,N_14185,N_14646);
nand U16004 (N_16004,N_14334,N_14923);
nand U16005 (N_16005,N_13561,N_14203);
nor U16006 (N_16006,N_13604,N_13620);
or U16007 (N_16007,N_14347,N_14181);
xnor U16008 (N_16008,N_13642,N_14699);
nand U16009 (N_16009,N_14870,N_13705);
nor U16010 (N_16010,N_13607,N_14752);
nand U16011 (N_16011,N_14436,N_14626);
and U16012 (N_16012,N_13736,N_13713);
nand U16013 (N_16013,N_14647,N_14984);
xor U16014 (N_16014,N_13867,N_13987);
xor U16015 (N_16015,N_14385,N_13889);
xnor U16016 (N_16016,N_13994,N_14022);
or U16017 (N_16017,N_14496,N_14500);
and U16018 (N_16018,N_14183,N_13542);
and U16019 (N_16019,N_14636,N_14298);
or U16020 (N_16020,N_14969,N_14997);
xnor U16021 (N_16021,N_14873,N_14281);
xnor U16022 (N_16022,N_14944,N_14727);
or U16023 (N_16023,N_14952,N_13667);
xor U16024 (N_16024,N_14883,N_14615);
or U16025 (N_16025,N_14466,N_14403);
xor U16026 (N_16026,N_14775,N_13603);
xor U16027 (N_16027,N_13957,N_13598);
and U16028 (N_16028,N_13799,N_14681);
nor U16029 (N_16029,N_13812,N_14294);
nor U16030 (N_16030,N_14994,N_14677);
xor U16031 (N_16031,N_13576,N_13765);
xor U16032 (N_16032,N_14746,N_14095);
nand U16033 (N_16033,N_14437,N_14854);
xnor U16034 (N_16034,N_14598,N_13853);
nor U16035 (N_16035,N_14076,N_14684);
or U16036 (N_16036,N_13687,N_14822);
and U16037 (N_16037,N_14584,N_13905);
nor U16038 (N_16038,N_14680,N_14160);
or U16039 (N_16039,N_14650,N_13556);
xor U16040 (N_16040,N_13858,N_14172);
xor U16041 (N_16041,N_13991,N_14989);
or U16042 (N_16042,N_14803,N_14263);
xnor U16043 (N_16043,N_14972,N_13625);
or U16044 (N_16044,N_14086,N_13605);
and U16045 (N_16045,N_14040,N_14728);
xor U16046 (N_16046,N_14430,N_14979);
nor U16047 (N_16047,N_14855,N_14058);
xnor U16048 (N_16048,N_14021,N_14266);
and U16049 (N_16049,N_13657,N_14236);
or U16050 (N_16050,N_14419,N_14298);
or U16051 (N_16051,N_13695,N_13855);
or U16052 (N_16052,N_13759,N_14843);
xor U16053 (N_16053,N_14087,N_14298);
nor U16054 (N_16054,N_14031,N_14290);
xor U16055 (N_16055,N_14341,N_13796);
xor U16056 (N_16056,N_13832,N_13940);
nand U16057 (N_16057,N_14640,N_13920);
xor U16058 (N_16058,N_14098,N_14454);
nor U16059 (N_16059,N_13744,N_14009);
nor U16060 (N_16060,N_14540,N_14139);
nor U16061 (N_16061,N_13703,N_14681);
xnor U16062 (N_16062,N_13834,N_14814);
nor U16063 (N_16063,N_14605,N_13548);
nand U16064 (N_16064,N_14669,N_14489);
or U16065 (N_16065,N_14881,N_13724);
or U16066 (N_16066,N_14529,N_14743);
or U16067 (N_16067,N_13563,N_13812);
xor U16068 (N_16068,N_14030,N_14711);
nand U16069 (N_16069,N_14539,N_13633);
or U16070 (N_16070,N_14471,N_14246);
or U16071 (N_16071,N_14563,N_13633);
nand U16072 (N_16072,N_14430,N_14683);
nand U16073 (N_16073,N_14646,N_13684);
nand U16074 (N_16074,N_14603,N_14927);
nor U16075 (N_16075,N_13823,N_13615);
and U16076 (N_16076,N_14522,N_14232);
nor U16077 (N_16077,N_14240,N_14826);
and U16078 (N_16078,N_14914,N_13695);
and U16079 (N_16079,N_13728,N_13715);
nand U16080 (N_16080,N_14299,N_13789);
nand U16081 (N_16081,N_14432,N_14194);
xnor U16082 (N_16082,N_14659,N_14024);
nand U16083 (N_16083,N_14652,N_14923);
xor U16084 (N_16084,N_14175,N_14045);
or U16085 (N_16085,N_14193,N_13748);
nand U16086 (N_16086,N_14088,N_13576);
and U16087 (N_16087,N_13901,N_14724);
or U16088 (N_16088,N_14574,N_14788);
and U16089 (N_16089,N_14550,N_13891);
or U16090 (N_16090,N_14603,N_13599);
nor U16091 (N_16091,N_14349,N_14367);
xnor U16092 (N_16092,N_14701,N_14802);
xor U16093 (N_16093,N_13938,N_13513);
or U16094 (N_16094,N_14848,N_14370);
nand U16095 (N_16095,N_14422,N_14490);
nor U16096 (N_16096,N_14544,N_14151);
and U16097 (N_16097,N_13719,N_14786);
xor U16098 (N_16098,N_13992,N_14472);
nor U16099 (N_16099,N_14235,N_14909);
xnor U16100 (N_16100,N_14529,N_14417);
xor U16101 (N_16101,N_14183,N_13664);
or U16102 (N_16102,N_14552,N_14795);
and U16103 (N_16103,N_13831,N_14413);
nor U16104 (N_16104,N_14061,N_14796);
nor U16105 (N_16105,N_13924,N_13749);
or U16106 (N_16106,N_14135,N_14536);
or U16107 (N_16107,N_13582,N_13618);
nor U16108 (N_16108,N_14238,N_13659);
nor U16109 (N_16109,N_13622,N_13905);
nand U16110 (N_16110,N_14308,N_14299);
xnor U16111 (N_16111,N_13722,N_13771);
and U16112 (N_16112,N_14799,N_14704);
nor U16113 (N_16113,N_13708,N_14344);
xnor U16114 (N_16114,N_14319,N_13753);
or U16115 (N_16115,N_14860,N_14704);
nand U16116 (N_16116,N_14204,N_13803);
nor U16117 (N_16117,N_14856,N_14800);
nand U16118 (N_16118,N_14236,N_14923);
xor U16119 (N_16119,N_13770,N_13982);
xor U16120 (N_16120,N_14495,N_14718);
and U16121 (N_16121,N_14413,N_13777);
or U16122 (N_16122,N_14365,N_14788);
or U16123 (N_16123,N_13502,N_14531);
nand U16124 (N_16124,N_14261,N_14236);
xor U16125 (N_16125,N_14620,N_14413);
nand U16126 (N_16126,N_14258,N_14950);
and U16127 (N_16127,N_13615,N_14455);
xor U16128 (N_16128,N_14541,N_13924);
and U16129 (N_16129,N_14704,N_14853);
nor U16130 (N_16130,N_14845,N_14437);
nand U16131 (N_16131,N_14185,N_14765);
xor U16132 (N_16132,N_14218,N_13650);
nand U16133 (N_16133,N_13623,N_14206);
nor U16134 (N_16134,N_14363,N_14993);
nand U16135 (N_16135,N_14606,N_13912);
xor U16136 (N_16136,N_14340,N_14085);
nand U16137 (N_16137,N_14815,N_13735);
xor U16138 (N_16138,N_14737,N_14322);
xnor U16139 (N_16139,N_14057,N_14700);
nor U16140 (N_16140,N_13784,N_14544);
nor U16141 (N_16141,N_13578,N_13790);
nor U16142 (N_16142,N_13545,N_13798);
or U16143 (N_16143,N_14423,N_14894);
or U16144 (N_16144,N_13612,N_13682);
nand U16145 (N_16145,N_14873,N_14534);
or U16146 (N_16146,N_14520,N_13901);
nand U16147 (N_16147,N_14738,N_13668);
or U16148 (N_16148,N_13873,N_14261);
nor U16149 (N_16149,N_13692,N_14659);
xor U16150 (N_16150,N_13632,N_14963);
or U16151 (N_16151,N_14864,N_13863);
nor U16152 (N_16152,N_13807,N_14680);
nor U16153 (N_16153,N_13744,N_13959);
xor U16154 (N_16154,N_13622,N_14422);
and U16155 (N_16155,N_14093,N_14153);
nor U16156 (N_16156,N_13883,N_14541);
xor U16157 (N_16157,N_14244,N_14232);
nor U16158 (N_16158,N_14474,N_13558);
and U16159 (N_16159,N_14711,N_13979);
and U16160 (N_16160,N_14491,N_13806);
and U16161 (N_16161,N_14683,N_14425);
nor U16162 (N_16162,N_13876,N_14116);
nand U16163 (N_16163,N_13683,N_14747);
and U16164 (N_16164,N_14222,N_14529);
and U16165 (N_16165,N_14703,N_14875);
or U16166 (N_16166,N_14071,N_14416);
or U16167 (N_16167,N_13650,N_14087);
nor U16168 (N_16168,N_14133,N_14085);
nand U16169 (N_16169,N_14515,N_14836);
or U16170 (N_16170,N_13920,N_14433);
nor U16171 (N_16171,N_13532,N_14082);
nand U16172 (N_16172,N_14884,N_14024);
nand U16173 (N_16173,N_14808,N_13508);
nor U16174 (N_16174,N_13750,N_14542);
and U16175 (N_16175,N_14220,N_14164);
nand U16176 (N_16176,N_14989,N_14595);
xor U16177 (N_16177,N_14037,N_14181);
and U16178 (N_16178,N_14702,N_13708);
xnor U16179 (N_16179,N_14281,N_14606);
nor U16180 (N_16180,N_14699,N_14610);
xnor U16181 (N_16181,N_14291,N_13890);
nand U16182 (N_16182,N_14629,N_14717);
nor U16183 (N_16183,N_14191,N_14235);
xnor U16184 (N_16184,N_14661,N_13586);
nor U16185 (N_16185,N_14883,N_13899);
or U16186 (N_16186,N_14483,N_14717);
and U16187 (N_16187,N_14447,N_13663);
nor U16188 (N_16188,N_14590,N_14324);
nor U16189 (N_16189,N_14165,N_14327);
or U16190 (N_16190,N_13760,N_14967);
xnor U16191 (N_16191,N_13696,N_14235);
nand U16192 (N_16192,N_14195,N_13542);
or U16193 (N_16193,N_14822,N_14021);
or U16194 (N_16194,N_14180,N_14566);
nand U16195 (N_16195,N_14098,N_13774);
nor U16196 (N_16196,N_14980,N_14631);
nand U16197 (N_16197,N_13529,N_14296);
or U16198 (N_16198,N_14227,N_14290);
or U16199 (N_16199,N_13771,N_14037);
xor U16200 (N_16200,N_14297,N_14368);
and U16201 (N_16201,N_14031,N_13700);
or U16202 (N_16202,N_14534,N_13723);
or U16203 (N_16203,N_13723,N_13833);
nand U16204 (N_16204,N_14172,N_13824);
and U16205 (N_16205,N_14664,N_14988);
nor U16206 (N_16206,N_14881,N_14094);
or U16207 (N_16207,N_14643,N_14443);
and U16208 (N_16208,N_14344,N_14920);
nand U16209 (N_16209,N_14667,N_13951);
and U16210 (N_16210,N_14455,N_13974);
nor U16211 (N_16211,N_14572,N_14146);
nor U16212 (N_16212,N_13836,N_14240);
nor U16213 (N_16213,N_13705,N_14788);
xnor U16214 (N_16214,N_14160,N_14527);
and U16215 (N_16215,N_13773,N_13767);
and U16216 (N_16216,N_14851,N_14475);
nor U16217 (N_16217,N_13926,N_14205);
nand U16218 (N_16218,N_14697,N_14967);
nand U16219 (N_16219,N_14144,N_14578);
nor U16220 (N_16220,N_13847,N_14933);
nand U16221 (N_16221,N_13811,N_14747);
xnor U16222 (N_16222,N_14327,N_14692);
nor U16223 (N_16223,N_14961,N_14699);
and U16224 (N_16224,N_14953,N_14893);
and U16225 (N_16225,N_14758,N_14430);
nand U16226 (N_16226,N_14808,N_13525);
xnor U16227 (N_16227,N_14255,N_14296);
nand U16228 (N_16228,N_14666,N_14164);
nand U16229 (N_16229,N_14454,N_13915);
xor U16230 (N_16230,N_14546,N_13876);
nand U16231 (N_16231,N_13809,N_14387);
xnor U16232 (N_16232,N_14688,N_13854);
or U16233 (N_16233,N_13589,N_14254);
and U16234 (N_16234,N_14283,N_14018);
and U16235 (N_16235,N_14885,N_14466);
or U16236 (N_16236,N_14100,N_14120);
nor U16237 (N_16237,N_14922,N_13807);
or U16238 (N_16238,N_13759,N_14279);
nand U16239 (N_16239,N_13824,N_13662);
and U16240 (N_16240,N_14670,N_14897);
nor U16241 (N_16241,N_14452,N_14700);
and U16242 (N_16242,N_14677,N_14967);
and U16243 (N_16243,N_14597,N_13790);
nor U16244 (N_16244,N_13880,N_14076);
nand U16245 (N_16245,N_14042,N_13828);
nor U16246 (N_16246,N_13897,N_13645);
nand U16247 (N_16247,N_14860,N_14394);
nor U16248 (N_16248,N_14364,N_13538);
and U16249 (N_16249,N_13745,N_13654);
and U16250 (N_16250,N_13663,N_14042);
and U16251 (N_16251,N_14904,N_14141);
xor U16252 (N_16252,N_14073,N_13627);
xor U16253 (N_16253,N_13655,N_14283);
and U16254 (N_16254,N_14998,N_13638);
or U16255 (N_16255,N_14468,N_14733);
and U16256 (N_16256,N_13517,N_14509);
or U16257 (N_16257,N_14453,N_14540);
xor U16258 (N_16258,N_14565,N_13626);
and U16259 (N_16259,N_13979,N_13656);
nand U16260 (N_16260,N_13838,N_14697);
or U16261 (N_16261,N_14778,N_14298);
or U16262 (N_16262,N_14334,N_14696);
xor U16263 (N_16263,N_13909,N_14293);
xnor U16264 (N_16264,N_13698,N_14492);
and U16265 (N_16265,N_14150,N_13832);
or U16266 (N_16266,N_14450,N_13667);
or U16267 (N_16267,N_14740,N_14938);
or U16268 (N_16268,N_13519,N_13980);
nand U16269 (N_16269,N_14171,N_14701);
or U16270 (N_16270,N_13600,N_14575);
and U16271 (N_16271,N_14366,N_14215);
nand U16272 (N_16272,N_14506,N_14308);
or U16273 (N_16273,N_14674,N_13865);
or U16274 (N_16274,N_14461,N_14247);
nand U16275 (N_16275,N_13937,N_14471);
nand U16276 (N_16276,N_13601,N_13827);
or U16277 (N_16277,N_14014,N_13686);
nand U16278 (N_16278,N_13895,N_13883);
or U16279 (N_16279,N_13634,N_14868);
xor U16280 (N_16280,N_14108,N_13953);
nor U16281 (N_16281,N_14683,N_14378);
nand U16282 (N_16282,N_14550,N_14383);
nor U16283 (N_16283,N_14771,N_13658);
nand U16284 (N_16284,N_13813,N_14651);
xnor U16285 (N_16285,N_14738,N_13899);
nor U16286 (N_16286,N_13786,N_14091);
and U16287 (N_16287,N_14255,N_14413);
or U16288 (N_16288,N_14878,N_14602);
and U16289 (N_16289,N_14709,N_14153);
xnor U16290 (N_16290,N_14694,N_14307);
nand U16291 (N_16291,N_13744,N_14965);
nand U16292 (N_16292,N_13816,N_14785);
nand U16293 (N_16293,N_14454,N_13543);
xor U16294 (N_16294,N_14039,N_13740);
nand U16295 (N_16295,N_14114,N_14807);
nor U16296 (N_16296,N_14506,N_14509);
or U16297 (N_16297,N_13560,N_13912);
or U16298 (N_16298,N_14173,N_14983);
or U16299 (N_16299,N_14781,N_14764);
or U16300 (N_16300,N_14373,N_14471);
xor U16301 (N_16301,N_14941,N_13703);
and U16302 (N_16302,N_13532,N_14831);
and U16303 (N_16303,N_14744,N_13918);
xnor U16304 (N_16304,N_14290,N_14810);
nor U16305 (N_16305,N_14377,N_14272);
or U16306 (N_16306,N_13820,N_14995);
or U16307 (N_16307,N_14430,N_14665);
and U16308 (N_16308,N_14570,N_14679);
nor U16309 (N_16309,N_14928,N_13674);
xor U16310 (N_16310,N_14328,N_13528);
or U16311 (N_16311,N_14048,N_14890);
xor U16312 (N_16312,N_14207,N_14785);
and U16313 (N_16313,N_14107,N_13847);
and U16314 (N_16314,N_14781,N_13897);
nand U16315 (N_16315,N_13575,N_14006);
and U16316 (N_16316,N_14941,N_13680);
xnor U16317 (N_16317,N_13610,N_14309);
xor U16318 (N_16318,N_14170,N_13752);
nand U16319 (N_16319,N_13646,N_13681);
nor U16320 (N_16320,N_13678,N_14466);
nand U16321 (N_16321,N_13969,N_14746);
nor U16322 (N_16322,N_14286,N_14818);
or U16323 (N_16323,N_14833,N_14838);
nor U16324 (N_16324,N_14200,N_14494);
and U16325 (N_16325,N_14333,N_14242);
or U16326 (N_16326,N_14923,N_13858);
xnor U16327 (N_16327,N_14810,N_14458);
and U16328 (N_16328,N_14306,N_13568);
nor U16329 (N_16329,N_14234,N_13678);
and U16330 (N_16330,N_14201,N_14055);
or U16331 (N_16331,N_14605,N_13582);
or U16332 (N_16332,N_14264,N_13858);
xor U16333 (N_16333,N_14397,N_14750);
nand U16334 (N_16334,N_13726,N_13918);
xnor U16335 (N_16335,N_13793,N_14232);
nand U16336 (N_16336,N_13626,N_14286);
or U16337 (N_16337,N_14124,N_14166);
xnor U16338 (N_16338,N_14700,N_14545);
or U16339 (N_16339,N_14722,N_13534);
nor U16340 (N_16340,N_13547,N_14657);
xnor U16341 (N_16341,N_13804,N_13999);
nor U16342 (N_16342,N_13678,N_13512);
nor U16343 (N_16343,N_13660,N_14157);
nor U16344 (N_16344,N_14907,N_14490);
or U16345 (N_16345,N_13677,N_14799);
nand U16346 (N_16346,N_14567,N_14737);
or U16347 (N_16347,N_13977,N_14424);
nor U16348 (N_16348,N_14267,N_14773);
nand U16349 (N_16349,N_14548,N_13717);
nor U16350 (N_16350,N_13659,N_14195);
nor U16351 (N_16351,N_14391,N_13979);
nor U16352 (N_16352,N_13531,N_13548);
nor U16353 (N_16353,N_14862,N_14415);
or U16354 (N_16354,N_14480,N_13714);
nor U16355 (N_16355,N_14783,N_13570);
nand U16356 (N_16356,N_13509,N_14007);
nand U16357 (N_16357,N_14162,N_14628);
nor U16358 (N_16358,N_13696,N_13633);
or U16359 (N_16359,N_14301,N_14323);
nor U16360 (N_16360,N_13610,N_13716);
xor U16361 (N_16361,N_14521,N_14329);
xnor U16362 (N_16362,N_14060,N_14484);
xnor U16363 (N_16363,N_14494,N_13668);
or U16364 (N_16364,N_14015,N_13824);
xnor U16365 (N_16365,N_13933,N_14891);
or U16366 (N_16366,N_14113,N_14188);
xor U16367 (N_16367,N_14243,N_14277);
and U16368 (N_16368,N_14846,N_14422);
xnor U16369 (N_16369,N_14977,N_14745);
and U16370 (N_16370,N_13545,N_14085);
xor U16371 (N_16371,N_14891,N_14296);
xor U16372 (N_16372,N_13629,N_14552);
nand U16373 (N_16373,N_13848,N_13750);
nor U16374 (N_16374,N_13635,N_14212);
xor U16375 (N_16375,N_13814,N_14090);
or U16376 (N_16376,N_13673,N_14741);
and U16377 (N_16377,N_14057,N_13706);
nor U16378 (N_16378,N_13751,N_14272);
nor U16379 (N_16379,N_13960,N_14998);
nand U16380 (N_16380,N_14133,N_13523);
or U16381 (N_16381,N_14735,N_14928);
or U16382 (N_16382,N_13547,N_14973);
and U16383 (N_16383,N_14616,N_14270);
or U16384 (N_16384,N_13917,N_14732);
or U16385 (N_16385,N_13725,N_14043);
or U16386 (N_16386,N_14215,N_14095);
and U16387 (N_16387,N_13580,N_13766);
xnor U16388 (N_16388,N_14351,N_13682);
nor U16389 (N_16389,N_13553,N_14619);
or U16390 (N_16390,N_13532,N_14876);
nand U16391 (N_16391,N_13702,N_14228);
nand U16392 (N_16392,N_14596,N_14071);
xor U16393 (N_16393,N_14676,N_13892);
or U16394 (N_16394,N_14210,N_14779);
or U16395 (N_16395,N_14587,N_14684);
nor U16396 (N_16396,N_14580,N_13667);
nor U16397 (N_16397,N_14686,N_14385);
or U16398 (N_16398,N_14195,N_13999);
or U16399 (N_16399,N_14635,N_14131);
xor U16400 (N_16400,N_14191,N_14485);
xnor U16401 (N_16401,N_14577,N_14817);
nand U16402 (N_16402,N_14328,N_14830);
and U16403 (N_16403,N_14330,N_14187);
and U16404 (N_16404,N_14617,N_13964);
nor U16405 (N_16405,N_14956,N_14525);
nor U16406 (N_16406,N_14858,N_14096);
or U16407 (N_16407,N_14965,N_14315);
and U16408 (N_16408,N_14148,N_13997);
and U16409 (N_16409,N_14264,N_14525);
nor U16410 (N_16410,N_13733,N_14645);
nand U16411 (N_16411,N_14771,N_13905);
nor U16412 (N_16412,N_14014,N_14009);
xnor U16413 (N_16413,N_14644,N_14296);
or U16414 (N_16414,N_14591,N_13773);
nand U16415 (N_16415,N_14287,N_13532);
xor U16416 (N_16416,N_14041,N_14292);
and U16417 (N_16417,N_14453,N_13850);
nor U16418 (N_16418,N_14558,N_14632);
nand U16419 (N_16419,N_14133,N_13688);
nand U16420 (N_16420,N_13691,N_14029);
and U16421 (N_16421,N_14606,N_14200);
xnor U16422 (N_16422,N_13995,N_13583);
xor U16423 (N_16423,N_14634,N_13566);
nand U16424 (N_16424,N_14324,N_14853);
xnor U16425 (N_16425,N_13745,N_14971);
nand U16426 (N_16426,N_14842,N_14480);
and U16427 (N_16427,N_14410,N_14676);
xnor U16428 (N_16428,N_14133,N_14647);
or U16429 (N_16429,N_13857,N_13930);
or U16430 (N_16430,N_13891,N_13830);
and U16431 (N_16431,N_14110,N_14849);
nand U16432 (N_16432,N_14676,N_14782);
nand U16433 (N_16433,N_14949,N_14844);
xor U16434 (N_16434,N_13692,N_14268);
xor U16435 (N_16435,N_14595,N_14670);
or U16436 (N_16436,N_14797,N_13692);
and U16437 (N_16437,N_14487,N_13696);
nor U16438 (N_16438,N_13825,N_14455);
xnor U16439 (N_16439,N_14945,N_13802);
nand U16440 (N_16440,N_13711,N_14587);
nand U16441 (N_16441,N_14462,N_14640);
xor U16442 (N_16442,N_14240,N_14594);
or U16443 (N_16443,N_13501,N_13518);
nand U16444 (N_16444,N_14346,N_14247);
nor U16445 (N_16445,N_13555,N_14558);
nand U16446 (N_16446,N_13949,N_14990);
xor U16447 (N_16447,N_14607,N_14606);
and U16448 (N_16448,N_14644,N_13953);
nand U16449 (N_16449,N_14168,N_14216);
or U16450 (N_16450,N_14696,N_14275);
nand U16451 (N_16451,N_13678,N_14711);
nand U16452 (N_16452,N_14812,N_13506);
nand U16453 (N_16453,N_13543,N_14480);
xnor U16454 (N_16454,N_14715,N_13579);
or U16455 (N_16455,N_14212,N_14147);
xnor U16456 (N_16456,N_14382,N_14195);
nor U16457 (N_16457,N_14725,N_14050);
nor U16458 (N_16458,N_13840,N_14336);
nand U16459 (N_16459,N_13696,N_13867);
xor U16460 (N_16460,N_14890,N_13796);
nor U16461 (N_16461,N_13752,N_13726);
xor U16462 (N_16462,N_14471,N_14908);
and U16463 (N_16463,N_14605,N_13718);
nor U16464 (N_16464,N_13625,N_14508);
nand U16465 (N_16465,N_14935,N_13880);
xor U16466 (N_16466,N_14819,N_14344);
or U16467 (N_16467,N_14405,N_14640);
and U16468 (N_16468,N_13796,N_13716);
or U16469 (N_16469,N_14616,N_14280);
nand U16470 (N_16470,N_14089,N_14077);
and U16471 (N_16471,N_14039,N_13683);
nor U16472 (N_16472,N_13532,N_14750);
and U16473 (N_16473,N_13875,N_13503);
or U16474 (N_16474,N_13771,N_14085);
and U16475 (N_16475,N_14825,N_14523);
xnor U16476 (N_16476,N_14649,N_14426);
and U16477 (N_16477,N_13767,N_14146);
or U16478 (N_16478,N_14772,N_13856);
nor U16479 (N_16479,N_14310,N_14573);
xnor U16480 (N_16480,N_14203,N_14029);
nand U16481 (N_16481,N_14435,N_13934);
and U16482 (N_16482,N_13918,N_14095);
nor U16483 (N_16483,N_14634,N_14660);
nand U16484 (N_16484,N_14226,N_14657);
xnor U16485 (N_16485,N_13608,N_13574);
and U16486 (N_16486,N_14697,N_13921);
or U16487 (N_16487,N_13873,N_14853);
and U16488 (N_16488,N_14829,N_14213);
and U16489 (N_16489,N_13631,N_13915);
or U16490 (N_16490,N_14113,N_14568);
nand U16491 (N_16491,N_13503,N_14819);
xor U16492 (N_16492,N_14703,N_13668);
nand U16493 (N_16493,N_14464,N_13834);
xnor U16494 (N_16494,N_13964,N_14838);
nor U16495 (N_16495,N_13940,N_14842);
and U16496 (N_16496,N_14412,N_13868);
or U16497 (N_16497,N_14499,N_14634);
and U16498 (N_16498,N_14518,N_13752);
nand U16499 (N_16499,N_13832,N_13612);
nor U16500 (N_16500,N_15674,N_15506);
nand U16501 (N_16501,N_16308,N_15536);
nor U16502 (N_16502,N_15466,N_15941);
and U16503 (N_16503,N_15170,N_15479);
and U16504 (N_16504,N_15884,N_16250);
nor U16505 (N_16505,N_15269,N_15007);
nand U16506 (N_16506,N_15091,N_15526);
nor U16507 (N_16507,N_15923,N_16443);
nor U16508 (N_16508,N_16026,N_15796);
and U16509 (N_16509,N_15021,N_16191);
xnor U16510 (N_16510,N_15003,N_15816);
nor U16511 (N_16511,N_15186,N_15885);
xor U16512 (N_16512,N_15891,N_15621);
or U16513 (N_16513,N_15283,N_15915);
and U16514 (N_16514,N_15857,N_15864);
or U16515 (N_16515,N_15082,N_15998);
or U16516 (N_16516,N_16396,N_16243);
and U16517 (N_16517,N_15121,N_16272);
xor U16518 (N_16518,N_15057,N_16051);
nand U16519 (N_16519,N_15415,N_15012);
and U16520 (N_16520,N_16167,N_15435);
nor U16521 (N_16521,N_16166,N_16011);
and U16522 (N_16522,N_15390,N_15689);
nand U16523 (N_16523,N_16284,N_16365);
xor U16524 (N_16524,N_15959,N_15574);
xor U16525 (N_16525,N_16182,N_15434);
and U16526 (N_16526,N_15395,N_16100);
or U16527 (N_16527,N_16296,N_15510);
or U16528 (N_16528,N_15639,N_15317);
nand U16529 (N_16529,N_15344,N_15203);
or U16530 (N_16530,N_16499,N_15356);
and U16531 (N_16531,N_16490,N_16138);
and U16532 (N_16532,N_15773,N_15538);
xor U16533 (N_16533,N_15267,N_15131);
nor U16534 (N_16534,N_16417,N_15784);
nand U16535 (N_16535,N_15762,N_15543);
xor U16536 (N_16536,N_15032,N_15111);
and U16537 (N_16537,N_15625,N_16486);
xor U16538 (N_16538,N_16299,N_16291);
nor U16539 (N_16539,N_16127,N_16162);
xnor U16540 (N_16540,N_16257,N_15198);
or U16541 (N_16541,N_15914,N_15527);
or U16542 (N_16542,N_16027,N_15491);
nand U16543 (N_16543,N_15164,N_16203);
and U16544 (N_16544,N_16117,N_15367);
and U16545 (N_16545,N_15238,N_15893);
nand U16546 (N_16546,N_16367,N_15063);
nand U16547 (N_16547,N_15712,N_15160);
or U16548 (N_16548,N_15078,N_15787);
xnor U16549 (N_16549,N_16454,N_15004);
and U16550 (N_16550,N_15558,N_16295);
and U16551 (N_16551,N_15006,N_15951);
and U16552 (N_16552,N_15060,N_16074);
nor U16553 (N_16553,N_15874,N_15447);
nand U16554 (N_16554,N_15464,N_15691);
nand U16555 (N_16555,N_16334,N_16481);
and U16556 (N_16556,N_16458,N_16316);
or U16557 (N_16557,N_16252,N_15336);
nor U16558 (N_16558,N_15204,N_16081);
nand U16559 (N_16559,N_15022,N_16022);
nand U16560 (N_16560,N_16105,N_16495);
nor U16561 (N_16561,N_16063,N_15109);
nand U16562 (N_16562,N_15715,N_16285);
nor U16563 (N_16563,N_15886,N_15542);
and U16564 (N_16564,N_15263,N_16419);
nor U16565 (N_16565,N_16180,N_15023);
xnor U16566 (N_16566,N_15226,N_16216);
nand U16567 (N_16567,N_15183,N_15671);
nor U16568 (N_16568,N_15988,N_15056);
and U16569 (N_16569,N_15562,N_16336);
and U16570 (N_16570,N_15942,N_15989);
nand U16571 (N_16571,N_15709,N_15075);
nor U16572 (N_16572,N_15058,N_16092);
nand U16573 (N_16573,N_15155,N_15190);
nor U16574 (N_16574,N_15159,N_15619);
or U16575 (N_16575,N_16229,N_15142);
nand U16576 (N_16576,N_15047,N_15644);
nand U16577 (N_16577,N_16386,N_15167);
and U16578 (N_16578,N_15286,N_15632);
and U16579 (N_16579,N_15778,N_16469);
and U16580 (N_16580,N_15532,N_15423);
and U16581 (N_16581,N_15281,N_16075);
xnor U16582 (N_16582,N_15152,N_15410);
nor U16583 (N_16583,N_15900,N_15494);
nor U16584 (N_16584,N_15848,N_15605);
nand U16585 (N_16585,N_15929,N_15404);
or U16586 (N_16586,N_15401,N_15596);
and U16587 (N_16587,N_15337,N_16032);
and U16588 (N_16588,N_15749,N_15855);
nor U16589 (N_16589,N_16165,N_15595);
xnor U16590 (N_16590,N_16418,N_15364);
and U16591 (N_16591,N_16094,N_16258);
and U16592 (N_16592,N_15661,N_16220);
or U16593 (N_16593,N_15085,N_15747);
and U16594 (N_16594,N_15055,N_15355);
xor U16595 (N_16595,N_16466,N_16485);
xor U16596 (N_16596,N_15833,N_16259);
nor U16597 (N_16597,N_15346,N_15373);
xor U16598 (N_16598,N_15692,N_15242);
or U16599 (N_16599,N_15617,N_16201);
or U16600 (N_16600,N_15975,N_16263);
and U16601 (N_16601,N_15991,N_15489);
and U16602 (N_16602,N_16325,N_15655);
nand U16603 (N_16603,N_15609,N_15456);
nor U16604 (N_16604,N_15546,N_16280);
and U16605 (N_16605,N_15037,N_16215);
or U16606 (N_16606,N_15629,N_15973);
or U16607 (N_16607,N_15398,N_15407);
and U16608 (N_16608,N_15842,N_15110);
xor U16609 (N_16609,N_15278,N_16471);
or U16610 (N_16610,N_15256,N_16474);
nor U16611 (N_16611,N_15241,N_15432);
or U16612 (N_16612,N_16430,N_16268);
nor U16613 (N_16613,N_15473,N_15174);
nor U16614 (N_16614,N_15406,N_16479);
nor U16615 (N_16615,N_16369,N_15879);
xnor U16616 (N_16616,N_15245,N_15880);
nand U16617 (N_16617,N_15881,N_15062);
nand U16618 (N_16618,N_16449,N_15871);
or U16619 (N_16619,N_16040,N_15824);
nor U16620 (N_16620,N_16424,N_15729);
xnor U16621 (N_16621,N_16394,N_15262);
and U16622 (N_16622,N_15995,N_16298);
nand U16623 (N_16623,N_16275,N_16120);
or U16624 (N_16624,N_15394,N_15053);
xor U16625 (N_16625,N_15901,N_15803);
nor U16626 (N_16626,N_16076,N_16340);
xor U16627 (N_16627,N_15334,N_15916);
and U16628 (N_16628,N_16233,N_16303);
or U16629 (N_16629,N_16234,N_16118);
or U16630 (N_16630,N_15505,N_16457);
xnor U16631 (N_16631,N_15522,N_15184);
xor U16632 (N_16632,N_15614,N_15737);
xnor U16633 (N_16633,N_15259,N_15011);
nor U16634 (N_16634,N_15601,N_16393);
nand U16635 (N_16635,N_15633,N_15268);
xnor U16636 (N_16636,N_16402,N_16213);
and U16637 (N_16637,N_15939,N_16097);
nor U16638 (N_16638,N_15731,N_16139);
nor U16639 (N_16639,N_15829,N_16315);
xor U16640 (N_16640,N_16082,N_15877);
nand U16641 (N_16641,N_15583,N_15497);
nand U16642 (N_16642,N_16174,N_15149);
nor U16643 (N_16643,N_15271,N_15636);
xnor U16644 (N_16644,N_15044,N_15104);
or U16645 (N_16645,N_16416,N_15986);
xnor U16646 (N_16646,N_15191,N_15845);
and U16647 (N_16647,N_15687,N_15124);
nand U16648 (N_16648,N_16008,N_16484);
xnor U16649 (N_16649,N_16169,N_16373);
xnor U16650 (N_16650,N_16281,N_15429);
or U16651 (N_16651,N_16143,N_15635);
and U16652 (N_16652,N_15148,N_15284);
nor U16653 (N_16653,N_15958,N_16384);
nand U16654 (N_16654,N_15428,N_16231);
or U16655 (N_16655,N_15113,N_16378);
or U16656 (N_16656,N_15924,N_16133);
nor U16657 (N_16657,N_15163,N_16435);
or U16658 (N_16658,N_15875,N_16072);
nand U16659 (N_16659,N_15618,N_15675);
nor U16660 (N_16660,N_15345,N_16034);
or U16661 (N_16661,N_15348,N_15150);
nor U16662 (N_16662,N_15000,N_15586);
nor U16663 (N_16663,N_15561,N_15457);
or U16664 (N_16664,N_16159,N_15422);
or U16665 (N_16665,N_15120,N_15265);
nand U16666 (N_16666,N_16442,N_15570);
and U16667 (N_16667,N_15782,N_16193);
nand U16668 (N_16668,N_15903,N_15417);
and U16669 (N_16669,N_16327,N_15067);
or U16670 (N_16670,N_15579,N_15726);
xor U16671 (N_16671,N_15734,N_15649);
nand U16672 (N_16672,N_15297,N_15952);
nor U16673 (N_16673,N_15819,N_15869);
or U16674 (N_16674,N_16031,N_15978);
and U16675 (N_16675,N_16428,N_16119);
and U16676 (N_16676,N_16462,N_16246);
and U16677 (N_16677,N_15324,N_15468);
xor U16678 (N_16678,N_15828,N_15225);
xnor U16679 (N_16679,N_15507,N_16056);
nand U16680 (N_16680,N_15197,N_16225);
nor U16681 (N_16681,N_15380,N_15928);
nand U16682 (N_16682,N_15698,N_15100);
nand U16683 (N_16683,N_16226,N_15512);
nor U16684 (N_16684,N_16144,N_15530);
xnor U16685 (N_16685,N_16247,N_15910);
nor U16686 (N_16686,N_15332,N_15308);
and U16687 (N_16687,N_16307,N_15779);
nand U16688 (N_16688,N_16088,N_15246);
or U16689 (N_16689,N_16354,N_15703);
and U16690 (N_16690,N_15654,N_15972);
xnor U16691 (N_16691,N_15450,N_16021);
nor U16692 (N_16692,N_15774,N_16161);
and U16693 (N_16693,N_15837,N_16408);
nand U16694 (N_16694,N_15823,N_15894);
nor U16695 (N_16695,N_15384,N_15327);
xnor U16696 (N_16696,N_15331,N_15354);
xnor U16697 (N_16697,N_16173,N_15573);
or U16698 (N_16698,N_15385,N_15790);
nand U16699 (N_16699,N_15777,N_15187);
and U16700 (N_16700,N_15863,N_15818);
nor U16701 (N_16701,N_16440,N_15430);
and U16702 (N_16702,N_16194,N_15335);
xor U16703 (N_16703,N_15213,N_16218);
nand U16704 (N_16704,N_15666,N_15568);
nor U16705 (N_16705,N_16413,N_15069);
nand U16706 (N_16706,N_16253,N_15396);
xor U16707 (N_16707,N_15288,N_16172);
xnor U16708 (N_16708,N_16184,N_15850);
or U16709 (N_16709,N_16489,N_15841);
nor U16710 (N_16710,N_15189,N_16439);
and U16711 (N_16711,N_15377,N_16477);
nor U16712 (N_16712,N_15471,N_15014);
nand U16713 (N_16713,N_15305,N_16112);
and U16714 (N_16714,N_15851,N_16451);
or U16715 (N_16715,N_15071,N_15125);
nand U16716 (N_16716,N_16244,N_15813);
nor U16717 (N_16717,N_16330,N_15755);
nor U16718 (N_16718,N_16175,N_16374);
xnor U16719 (N_16719,N_15146,N_15815);
and U16720 (N_16720,N_15221,N_15553);
and U16721 (N_16721,N_16324,N_15376);
xor U16722 (N_16722,N_16322,N_15209);
and U16723 (N_16723,N_15472,N_15514);
and U16724 (N_16724,N_15165,N_16211);
xnor U16725 (N_16725,N_15275,N_16065);
nand U16726 (N_16726,N_16420,N_15386);
xnor U16727 (N_16727,N_15157,N_15810);
xnor U16728 (N_16728,N_15913,N_16106);
or U16729 (N_16729,N_15746,N_15511);
or U16730 (N_16730,N_15442,N_15220);
nand U16731 (N_16731,N_16238,N_15858);
or U16732 (N_16732,N_15902,N_16096);
or U16733 (N_16733,N_16041,N_15904);
nor U16734 (N_16734,N_15086,N_15660);
or U16735 (N_16735,N_15919,N_16493);
nand U16736 (N_16736,N_15252,N_16292);
and U16737 (N_16737,N_16107,N_15413);
xnor U16738 (N_16738,N_15525,N_16068);
or U16739 (N_16739,N_16048,N_15482);
nand U16740 (N_16740,N_15716,N_15343);
xor U16741 (N_16741,N_16332,N_15061);
nand U16742 (N_16742,N_15616,N_15683);
nand U16743 (N_16743,N_15748,N_15678);
nand U16744 (N_16744,N_15054,N_16249);
nor U16745 (N_16745,N_15711,N_15483);
xnor U16746 (N_16746,N_15719,N_15201);
nand U16747 (N_16747,N_16488,N_15688);
or U16748 (N_16748,N_15300,N_15768);
nand U16749 (N_16749,N_15892,N_15177);
nor U16750 (N_16750,N_15772,N_16000);
nand U16751 (N_16751,N_16223,N_15452);
or U16752 (N_16752,N_16104,N_16015);
and U16753 (N_16753,N_15378,N_15066);
and U16754 (N_16754,N_15969,N_15135);
xnor U16755 (N_16755,N_16411,N_15436);
xnor U16756 (N_16756,N_15200,N_16344);
nor U16757 (N_16757,N_15025,N_15362);
nand U16758 (N_16758,N_15865,N_16261);
or U16759 (N_16759,N_16183,N_15215);
nor U16760 (N_16760,N_16073,N_15883);
nand U16761 (N_16761,N_15714,N_15295);
and U16762 (N_16762,N_16084,N_15079);
nor U16763 (N_16763,N_16412,N_15218);
or U16764 (N_16764,N_15908,N_16338);
and U16765 (N_16765,N_15577,N_15622);
or U16766 (N_16766,N_15230,N_16140);
and U16767 (N_16767,N_16160,N_16079);
or U16768 (N_16768,N_16029,N_16236);
and U16769 (N_16769,N_15722,N_15946);
or U16770 (N_16770,N_15580,N_16239);
nand U16771 (N_16771,N_15383,N_16460);
and U16772 (N_16772,N_15103,N_15002);
and U16773 (N_16773,N_15582,N_15181);
nand U16774 (N_16774,N_15860,N_16347);
and U16775 (N_16775,N_15329,N_15807);
xnor U16776 (N_16776,N_15279,N_15500);
nand U16777 (N_16777,N_15227,N_15013);
nor U16778 (N_16778,N_15584,N_15647);
nor U16779 (N_16779,N_15788,N_15909);
or U16780 (N_16780,N_16364,N_16152);
and U16781 (N_16781,N_16366,N_15094);
or U16782 (N_16782,N_16099,N_15208);
nand U16783 (N_16783,N_15294,N_16108);
and U16784 (N_16784,N_15027,N_15859);
xnor U16785 (N_16785,N_16059,N_16320);
xor U16786 (N_16786,N_15597,N_16156);
nand U16787 (N_16787,N_16482,N_16046);
and U16788 (N_16788,N_16290,N_16300);
nand U16789 (N_16789,N_15598,N_15721);
and U16790 (N_16790,N_15475,N_15708);
or U16791 (N_16791,N_15825,N_16012);
and U16792 (N_16792,N_15992,N_16102);
xor U16793 (N_16793,N_15224,N_15485);
or U16794 (N_16794,N_15264,N_16389);
xor U16795 (N_16795,N_15431,N_15634);
nor U16796 (N_16796,N_15166,N_15347);
xor U16797 (N_16797,N_16128,N_16494);
nand U16798 (N_16798,N_15667,N_15775);
xor U16799 (N_16799,N_15339,N_16078);
and U16800 (N_16800,N_16197,N_15766);
nor U16801 (N_16801,N_15814,N_15196);
and U16802 (N_16802,N_15374,N_15802);
or U16803 (N_16803,N_16400,N_15890);
nor U16804 (N_16804,N_16368,N_16464);
and U16805 (N_16805,N_15141,N_15742);
or U16806 (N_16806,N_16328,N_16235);
xor U16807 (N_16807,N_15576,N_15707);
nor U16808 (N_16808,N_15136,N_16309);
and U16809 (N_16809,N_15296,N_16002);
and U16810 (N_16810,N_15981,N_16221);
and U16811 (N_16811,N_15730,N_15897);
xor U16812 (N_16812,N_15693,N_16438);
xnor U16813 (N_16813,N_15838,N_16276);
or U16814 (N_16814,N_16146,N_15682);
or U16815 (N_16815,N_15304,N_16245);
nand U16816 (N_16816,N_15441,N_15963);
nor U16817 (N_16817,N_16318,N_15448);
nor U16818 (N_16818,N_15817,N_15761);
nand U16819 (N_16819,N_15470,N_15361);
nor U16820 (N_16820,N_16080,N_15794);
nor U16821 (N_16821,N_15797,N_16129);
nor U16822 (N_16822,N_15178,N_16122);
nor U16823 (N_16823,N_15199,N_16007);
nor U16824 (N_16824,N_15455,N_15499);
and U16825 (N_16825,N_15798,N_15076);
and U16826 (N_16826,N_15535,N_16093);
nand U16827 (N_16827,N_16004,N_15031);
or U16828 (N_16828,N_15509,N_15623);
xnor U16829 (N_16829,N_16432,N_15559);
nand U16830 (N_16830,N_15397,N_15926);
or U16831 (N_16831,N_15849,N_16423);
xnor U16832 (N_16832,N_15552,N_15938);
or U16833 (N_16833,N_15306,N_15095);
and U16834 (N_16834,N_15982,N_15905);
and U16835 (N_16835,N_16351,N_16209);
nor U16836 (N_16836,N_15566,N_16358);
xor U16837 (N_16837,N_15481,N_15631);
nand U16838 (N_16838,N_15314,N_15805);
nand U16839 (N_16839,N_15759,N_16025);
and U16840 (N_16840,N_16042,N_15811);
or U16841 (N_16841,N_15302,N_15469);
nor U16842 (N_16842,N_16446,N_15289);
xor U16843 (N_16843,N_16331,N_15366);
nand U16844 (N_16844,N_15180,N_16110);
and U16845 (N_16845,N_15912,N_15705);
and U16846 (N_16846,N_15443,N_15740);
nand U16847 (N_16847,N_16049,N_16288);
xor U16848 (N_16848,N_15960,N_15188);
nand U16849 (N_16849,N_15993,N_15602);
and U16850 (N_16850,N_16476,N_15114);
and U16851 (N_16851,N_15389,N_16103);
xnor U16852 (N_16852,N_16382,N_15222);
and U16853 (N_16853,N_16465,N_16343);
and U16854 (N_16854,N_15676,N_16111);
nand U16855 (N_16855,N_15801,N_16035);
xor U16856 (N_16856,N_15462,N_16434);
xor U16857 (N_16857,N_15641,N_16200);
or U16858 (N_16858,N_16459,N_16228);
xor U16859 (N_16859,N_15359,N_15502);
or U16860 (N_16860,N_16188,N_15418);
nor U16861 (N_16861,N_15301,N_15783);
nand U16862 (N_16862,N_16426,N_16240);
nand U16863 (N_16863,N_15706,N_15353);
nand U16864 (N_16864,N_15550,N_15133);
and U16865 (N_16865,N_15997,N_15700);
or U16866 (N_16866,N_16461,N_16095);
nor U16867 (N_16867,N_16199,N_16154);
nor U16868 (N_16868,N_16405,N_16131);
nand U16869 (N_16869,N_15876,N_15433);
nand U16870 (N_16870,N_16468,N_15255);
nand U16871 (N_16871,N_15216,N_15854);
nor U16872 (N_16872,N_16187,N_15690);
nor U16873 (N_16873,N_16085,N_15681);
nor U16874 (N_16874,N_15987,N_16248);
or U16875 (N_16875,N_16254,N_16134);
xor U16876 (N_16876,N_16319,N_16089);
xor U16877 (N_16877,N_15097,N_16415);
and U16878 (N_16878,N_15424,N_15889);
or U16879 (N_16879,N_15717,N_15239);
xor U16880 (N_16880,N_15931,N_15513);
xnor U16881 (N_16881,N_15474,N_15024);
xnor U16882 (N_16882,N_16407,N_16487);
xnor U16883 (N_16883,N_16064,N_15843);
xnor U16884 (N_16884,N_16398,N_15699);
nand U16885 (N_16885,N_16157,N_15323);
or U16886 (N_16886,N_15786,N_15036);
nand U16887 (N_16887,N_16053,N_16342);
nand U16888 (N_16888,N_16219,N_15615);
and U16889 (N_16889,N_15957,N_15650);
and U16890 (N_16890,N_15657,N_16353);
nand U16891 (N_16891,N_16345,N_15882);
xnor U16892 (N_16892,N_15272,N_16142);
xnor U16893 (N_16893,N_15836,N_15990);
nand U16894 (N_16894,N_15454,N_15234);
xnor U16895 (N_16895,N_15028,N_15545);
xnor U16896 (N_16896,N_15669,N_15080);
or U16897 (N_16897,N_15211,N_16313);
or U16898 (N_16898,N_15585,N_15974);
nand U16899 (N_16899,N_16116,N_16274);
nor U16900 (N_16900,N_15064,N_15034);
and U16901 (N_16901,N_15092,N_16020);
xor U16902 (N_16902,N_15822,N_15808);
or U16903 (N_16903,N_15358,N_16033);
xnor U16904 (N_16904,N_15273,N_16388);
xnor U16905 (N_16905,N_15467,N_16312);
xor U16906 (N_16906,N_16043,N_15516);
nor U16907 (N_16907,N_16086,N_15756);
xor U16908 (N_16908,N_15073,N_16463);
nor U16909 (N_16909,N_15735,N_16297);
nor U16910 (N_16910,N_15106,N_15587);
xor U16911 (N_16911,N_15593,N_15459);
xnor U16912 (N_16912,N_16287,N_16314);
nand U16913 (N_16913,N_15194,N_15920);
or U16914 (N_16914,N_15059,N_15307);
xnor U16915 (N_16915,N_16385,N_16409);
xnor U16916 (N_16916,N_15446,N_16017);
or U16917 (N_16917,N_15704,N_15572);
xnor U16918 (N_16918,N_15090,N_16179);
nand U16919 (N_16919,N_15371,N_15476);
xor U16920 (N_16920,N_16425,N_15870);
and U16921 (N_16921,N_16422,N_15101);
nor U16922 (N_16922,N_15463,N_16185);
xor U16923 (N_16923,N_15340,N_15927);
nand U16924 (N_16924,N_15640,N_16371);
nand U16925 (N_16925,N_16052,N_15233);
or U16926 (N_16926,N_15804,N_15438);
or U16927 (N_16927,N_15795,N_15846);
xnor U16928 (N_16928,N_15967,N_16195);
xor U16929 (N_16929,N_15381,N_15770);
and U16930 (N_16930,N_16153,N_15503);
nand U16931 (N_16931,N_15590,N_16189);
nor U16932 (N_16932,N_16497,N_15139);
nand U16933 (N_16933,N_16141,N_15531);
xnor U16934 (N_16934,N_15961,N_16136);
nor U16935 (N_16935,N_16237,N_15065);
and U16936 (N_16936,N_15309,N_16436);
or U16937 (N_16937,N_15117,N_15820);
and U16938 (N_16938,N_16202,N_15979);
and U16939 (N_16939,N_15932,N_16121);
nor U16940 (N_16940,N_15628,N_15895);
xnor U16941 (N_16941,N_16427,N_15405);
nand U16942 (N_16942,N_15030,N_15498);
and U16943 (N_16943,N_15293,N_15051);
nor U16944 (N_16944,N_15556,N_15486);
and U16945 (N_16945,N_15607,N_15564);
and U16946 (N_16946,N_15099,N_16145);
nor U16947 (N_16947,N_15392,N_15781);
nand U16948 (N_16948,N_15368,N_15533);
or U16949 (N_16949,N_16289,N_15320);
and U16950 (N_16950,N_15282,N_15352);
nor U16951 (N_16951,N_16387,N_15548);
or U16952 (N_16952,N_15231,N_15557);
nand U16953 (N_16953,N_15236,N_15119);
and U16954 (N_16954,N_16380,N_15411);
nor U16955 (N_16955,N_16491,N_15757);
or U16956 (N_16956,N_16270,N_15753);
xnor U16957 (N_16957,N_15020,N_15672);
or U16958 (N_16958,N_15444,N_16058);
xnor U16959 (N_16959,N_16083,N_15754);
nor U16960 (N_16960,N_15313,N_15738);
and U16961 (N_16961,N_15330,N_15555);
nor U16962 (N_16962,N_15484,N_15287);
and U16963 (N_16963,N_16264,N_16186);
nand U16964 (N_16964,N_15154,N_15250);
and U16965 (N_16965,N_15780,N_16473);
nor U16966 (N_16966,N_16356,N_15326);
nand U16967 (N_16967,N_15243,N_16294);
or U16968 (N_16968,N_15249,N_15713);
nor U16969 (N_16969,N_15899,N_15769);
or U16970 (N_16970,N_15604,N_15945);
xor U16971 (N_16971,N_15541,N_16355);
xor U16972 (N_16972,N_15303,N_15720);
or U16973 (N_16973,N_15663,N_16359);
nor U16974 (N_16974,N_15126,N_15840);
or U16975 (N_16975,N_15276,N_15581);
or U16976 (N_16976,N_16109,N_16467);
nand U16977 (N_16977,N_15478,N_16406);
nand U16978 (N_16978,N_16403,N_16341);
nand U16979 (N_16979,N_15789,N_16024);
and U16980 (N_16980,N_16410,N_15785);
or U16981 (N_16981,N_15019,N_15270);
or U16982 (N_16982,N_16256,N_15116);
and U16983 (N_16983,N_15985,N_15685);
nand U16984 (N_16984,N_16311,N_15937);
xnor U16985 (N_16985,N_16452,N_15936);
or U16986 (N_16986,N_15962,N_15944);
xnor U16987 (N_16987,N_15156,N_15943);
or U16988 (N_16988,N_15567,N_15068);
or U16989 (N_16989,N_15257,N_15399);
nor U16990 (N_16990,N_15247,N_15529);
and U16991 (N_16991,N_15112,N_15161);
and U16992 (N_16992,N_16126,N_15763);
nand U16993 (N_16993,N_15862,N_15016);
or U16994 (N_16994,N_16321,N_16090);
and U16995 (N_16995,N_16448,N_16401);
xnor U16996 (N_16996,N_16492,N_16196);
or U16997 (N_16997,N_15603,N_16204);
nand U16998 (N_16998,N_15048,N_16114);
and U16999 (N_16999,N_16445,N_15369);
nand U17000 (N_17000,N_15659,N_15606);
xor U17001 (N_17001,N_15643,N_15311);
or U17002 (N_17002,N_15005,N_15906);
nand U17003 (N_17003,N_15665,N_15084);
and U17004 (N_17004,N_16306,N_16010);
nand U17005 (N_17005,N_15624,N_15206);
and U17006 (N_17006,N_16352,N_15724);
or U17007 (N_17007,N_15743,N_16333);
and U17008 (N_17008,N_15844,N_15158);
xnor U17009 (N_17009,N_15662,N_15108);
nor U17010 (N_17010,N_16171,N_15725);
nand U17011 (N_17011,N_16301,N_16164);
nand U17012 (N_17012,N_15192,N_16363);
xnor U17013 (N_17013,N_15129,N_16055);
nor U17014 (N_17014,N_15096,N_15280);
or U17015 (N_17015,N_15228,N_15664);
or U17016 (N_17016,N_16148,N_15964);
or U17017 (N_17017,N_15925,N_15151);
xor U17018 (N_17018,N_15977,N_15569);
nand U17019 (N_17019,N_15518,N_15420);
or U17020 (N_17020,N_16057,N_16441);
xnor U17021 (N_17021,N_16496,N_15695);
and U17022 (N_17022,N_15809,N_15852);
or U17023 (N_17023,N_16421,N_15767);
and U17024 (N_17024,N_16036,N_15451);
or U17025 (N_17025,N_15984,N_15918);
nand U17026 (N_17026,N_16016,N_16271);
xor U17027 (N_17027,N_15656,N_15949);
and U17028 (N_17028,N_15517,N_16050);
nor U17029 (N_17029,N_15077,N_15922);
or U17030 (N_17030,N_15029,N_16071);
and U17031 (N_17031,N_15940,N_15427);
xor U17032 (N_17032,N_15350,N_15515);
or U17033 (N_17033,N_15393,N_16431);
xor U17034 (N_17034,N_15147,N_15537);
and U17035 (N_17035,N_15832,N_15646);
nor U17036 (N_17036,N_16390,N_16286);
or U17037 (N_17037,N_16267,N_15701);
or U17038 (N_17038,N_15207,N_16391);
nand U17039 (N_17039,N_16155,N_15038);
nor U17040 (N_17040,N_16087,N_15608);
nand U17041 (N_17041,N_15684,N_16232);
nand U17042 (N_17042,N_15403,N_15169);
or U17043 (N_17043,N_16381,N_16113);
or U17044 (N_17044,N_15519,N_15130);
nand U17045 (N_17045,N_15254,N_16001);
xnor U17046 (N_17046,N_15727,N_15145);
nor U17047 (N_17047,N_15360,N_15834);
or U17048 (N_17048,N_15520,N_15477);
or U17049 (N_17049,N_15523,N_15179);
nor U17050 (N_17050,N_15449,N_15122);
nor U17051 (N_17051,N_15847,N_16061);
nand U17052 (N_17052,N_16210,N_16009);
xnor U17053 (N_17053,N_15524,N_15043);
or U17054 (N_17054,N_16135,N_16003);
and U17055 (N_17055,N_15261,N_15081);
and U17056 (N_17056,N_15668,N_15202);
xnor U17057 (N_17057,N_16149,N_16060);
and U17058 (N_17058,N_15439,N_16323);
or U17059 (N_17059,N_16310,N_15793);
xnor U17060 (N_17060,N_15052,N_15137);
nand U17061 (N_17061,N_15102,N_15492);
and U17062 (N_17062,N_15504,N_15322);
nand U17063 (N_17063,N_16392,N_15887);
nand U17064 (N_17064,N_15930,N_16326);
nand U17065 (N_17065,N_15547,N_15501);
nand U17066 (N_17066,N_15277,N_15496);
nand U17067 (N_17067,N_15440,N_15408);
and U17068 (N_17068,N_16349,N_15610);
xnor U17069 (N_17069,N_16335,N_15637);
or U17070 (N_17070,N_15045,N_15312);
or U17071 (N_17071,N_15266,N_15839);
xor U17072 (N_17072,N_15934,N_15175);
or U17073 (N_17073,N_15445,N_16013);
nor U17074 (N_17074,N_15379,N_15115);
and U17075 (N_17075,N_15049,N_16177);
or U17076 (N_17076,N_15588,N_16251);
nor U17077 (N_17077,N_15365,N_15765);
nor U17078 (N_17078,N_16455,N_16337);
and U17079 (N_17079,N_15351,N_15853);
xor U17080 (N_17080,N_15866,N_15193);
nor U17081 (N_17081,N_15315,N_16444);
or U17082 (N_17082,N_15465,N_16070);
xnor U17083 (N_17083,N_16038,N_15258);
nor U17084 (N_17084,N_15911,N_15458);
or U17085 (N_17085,N_16293,N_15341);
nand U17086 (N_17086,N_16147,N_15764);
nor U17087 (N_17087,N_15143,N_15260);
nand U17088 (N_17088,N_15645,N_15253);
and U17089 (N_17089,N_16151,N_15409);
or U17090 (N_17090,N_16091,N_16304);
and U17091 (N_17091,N_15642,N_16170);
nand U17092 (N_17092,N_15093,N_15888);
xor U17093 (N_17093,N_15954,N_15419);
xnor U17094 (N_17094,N_15968,N_15387);
or U17095 (N_17095,N_15402,N_15589);
xnor U17096 (N_17096,N_15375,N_15074);
xor U17097 (N_17097,N_15776,N_15627);
nand U17098 (N_17098,N_16005,N_16150);
and U17099 (N_17099,N_16348,N_15026);
or U17100 (N_17100,N_15907,N_15771);
and U17101 (N_17101,N_15040,N_15630);
nor U17102 (N_17102,N_15976,N_15460);
nor U17103 (N_17103,N_15599,N_15338);
nor U17104 (N_17104,N_16475,N_15235);
nand U17105 (N_17105,N_15240,N_15551);
nor U17106 (N_17106,N_15425,N_15349);
xor U17107 (N_17107,N_15575,N_15274);
nor U17108 (N_17108,N_16023,N_15563);
and U17109 (N_17109,N_16230,N_15921);
and U17110 (N_17110,N_15996,N_15412);
nor U17111 (N_17111,N_15758,N_15947);
nor U17112 (N_17112,N_15736,N_16453);
or U17113 (N_17113,N_16192,N_15299);
xor U17114 (N_17114,N_16450,N_16039);
nand U17115 (N_17115,N_16357,N_15290);
or U17116 (N_17116,N_15744,N_16255);
nor U17117 (N_17117,N_15799,N_16047);
and U17118 (N_17118,N_15008,N_15089);
nor U17119 (N_17119,N_16397,N_15237);
nand U17120 (N_17120,N_16329,N_15426);
nand U17121 (N_17121,N_16376,N_15176);
xor U17122 (N_17122,N_15072,N_16273);
or U17123 (N_17123,N_16483,N_16456);
nand U17124 (N_17124,N_15565,N_15826);
nand U17125 (N_17125,N_15751,N_16217);
or U17126 (N_17126,N_15001,N_16437);
or U17127 (N_17127,N_15856,N_15953);
nand U17128 (N_17128,N_15105,N_16429);
nor U17129 (N_17129,N_15251,N_15153);
nand U17130 (N_17130,N_16176,N_15041);
and U17131 (N_17131,N_15528,N_15223);
or U17132 (N_17132,N_15521,N_15493);
nor U17133 (N_17133,N_15752,N_16018);
xnor U17134 (N_17134,N_15098,N_15050);
xnor U17135 (N_17135,N_15718,N_15232);
xnor U17136 (N_17136,N_16350,N_16472);
xnor U17137 (N_17137,N_15611,N_15333);
nor U17138 (N_17138,N_15612,N_15214);
and U17139 (N_17139,N_16379,N_16361);
and U17140 (N_17140,N_15980,N_16006);
xor U17141 (N_17141,N_15830,N_15453);
nor U17142 (N_17142,N_15391,N_16399);
or U17143 (N_17143,N_15806,N_16066);
xnor U17144 (N_17144,N_15873,N_15310);
or U17145 (N_17145,N_15679,N_15594);
or U17146 (N_17146,N_15620,N_16178);
or U17147 (N_17147,N_16190,N_15745);
and U17148 (N_17148,N_15549,N_15070);
nand U17149 (N_17149,N_16124,N_15971);
or U17150 (N_17150,N_15400,N_16480);
nand U17151 (N_17151,N_16214,N_15298);
or U17152 (N_17152,N_15950,N_15741);
xor U17153 (N_17153,N_16241,N_16123);
nor U17154 (N_17154,N_16222,N_16282);
nor U17155 (N_17155,N_15896,N_16054);
or U17156 (N_17156,N_15321,N_15219);
nor U17157 (N_17157,N_15087,N_16278);
xor U17158 (N_17158,N_15686,N_15461);
xor U17159 (N_17159,N_16375,N_15680);
and U17160 (N_17160,N_15898,N_16265);
xnor U17161 (N_17161,N_15983,N_15750);
xor U17162 (N_17162,N_15651,N_15325);
xor U17163 (N_17163,N_16205,N_15123);
nand U17164 (N_17164,N_16395,N_16069);
and U17165 (N_17165,N_15677,N_16206);
xor U17166 (N_17166,N_15694,N_16125);
or U17167 (N_17167,N_15172,N_15917);
nand U17168 (N_17168,N_15128,N_15015);
and U17169 (N_17169,N_15970,N_15118);
xnor U17170 (N_17170,N_16370,N_16478);
and U17171 (N_17171,N_16158,N_15878);
nor U17172 (N_17172,N_15956,N_16062);
xnor U17173 (N_17173,N_16163,N_15046);
nor U17174 (N_17174,N_15812,N_15591);
and U17175 (N_17175,N_15723,N_15653);
nand U17176 (N_17176,N_16101,N_15861);
nand U17177 (N_17177,N_15370,N_15144);
nor U17178 (N_17178,N_16433,N_15539);
xnor U17179 (N_17179,N_15955,N_16212);
or U17180 (N_17180,N_15648,N_16181);
nor U17181 (N_17181,N_16019,N_15658);
nor U17182 (N_17182,N_15792,N_16470);
and U17183 (N_17183,N_16132,N_15437);
and U17184 (N_17184,N_15292,N_15107);
or U17185 (N_17185,N_15244,N_15592);
xor U17186 (N_17186,N_15010,N_15088);
and U17187 (N_17187,N_16414,N_16317);
nor U17188 (N_17188,N_16067,N_15217);
and U17189 (N_17189,N_15132,N_15821);
nand U17190 (N_17190,N_15488,N_15033);
and U17191 (N_17191,N_15933,N_16044);
xor U17192 (N_17192,N_15127,N_15480);
or U17193 (N_17193,N_15372,N_15318);
or U17194 (N_17194,N_16227,N_15554);
xor U17195 (N_17195,N_15171,N_16262);
or U17196 (N_17196,N_15739,N_15138);
or U17197 (N_17197,N_15017,N_16269);
nand U17198 (N_17198,N_16198,N_16045);
xnor U17199 (N_17199,N_15652,N_16305);
nor U17200 (N_17200,N_15319,N_15702);
nand U17201 (N_17201,N_15508,N_15134);
nand U17202 (N_17202,N_16098,N_15328);
nor U17203 (N_17203,N_15414,N_15416);
xor U17204 (N_17204,N_15835,N_15600);
xor U17205 (N_17205,N_15534,N_15999);
and U17206 (N_17206,N_15827,N_16266);
xnor U17207 (N_17207,N_15966,N_16037);
nor U17208 (N_17208,N_15935,N_16302);
or U17209 (N_17209,N_15800,N_16242);
nand U17210 (N_17210,N_15018,N_16168);
nor U17211 (N_17211,N_16028,N_15673);
xnor U17212 (N_17212,N_15831,N_15560);
or U17213 (N_17213,N_15039,N_15638);
nand U17214 (N_17214,N_15626,N_15421);
nand U17215 (N_17215,N_15490,N_15316);
nor U17216 (N_17216,N_15162,N_16498);
and U17217 (N_17217,N_15697,N_15382);
nor U17218 (N_17218,N_16115,N_16207);
or U17219 (N_17219,N_15195,N_15760);
nand U17220 (N_17220,N_15363,N_15868);
and U17221 (N_17221,N_16447,N_15791);
xnor U17222 (N_17222,N_16224,N_15544);
and U17223 (N_17223,N_15285,N_15291);
or U17224 (N_17224,N_16360,N_15495);
xnor U17225 (N_17225,N_16377,N_15571);
nor U17226 (N_17226,N_15948,N_15696);
and U17227 (N_17227,N_15388,N_15670);
or U17228 (N_17228,N_15083,N_16279);
and U17229 (N_17229,N_15613,N_15168);
nor U17230 (N_17230,N_15185,N_16283);
or U17231 (N_17231,N_15867,N_16014);
or U17232 (N_17232,N_15173,N_15540);
and U17233 (N_17233,N_15035,N_15872);
nand U17234 (N_17234,N_16030,N_15229);
nand U17235 (N_17235,N_16137,N_16130);
or U17236 (N_17236,N_15342,N_15487);
and U17237 (N_17237,N_15009,N_15733);
xnor U17238 (N_17238,N_15140,N_16339);
nand U17239 (N_17239,N_15578,N_15182);
xor U17240 (N_17240,N_16277,N_16362);
xnor U17241 (N_17241,N_16372,N_16260);
nor U17242 (N_17242,N_15248,N_15965);
xnor U17243 (N_17243,N_15994,N_16404);
xor U17244 (N_17244,N_16346,N_15210);
nor U17245 (N_17245,N_15732,N_15728);
or U17246 (N_17246,N_15205,N_15042);
xor U17247 (N_17247,N_16383,N_15212);
or U17248 (N_17248,N_15357,N_16208);
or U17249 (N_17249,N_15710,N_16077);
or U17250 (N_17250,N_15507,N_15401);
nand U17251 (N_17251,N_15790,N_15362);
or U17252 (N_17252,N_15782,N_15688);
nand U17253 (N_17253,N_16081,N_16330);
and U17254 (N_17254,N_16344,N_15542);
xnor U17255 (N_17255,N_15190,N_15123);
xor U17256 (N_17256,N_15414,N_16438);
or U17257 (N_17257,N_16380,N_16361);
or U17258 (N_17258,N_15882,N_15042);
or U17259 (N_17259,N_15572,N_15745);
xnor U17260 (N_17260,N_15970,N_15993);
nor U17261 (N_17261,N_16061,N_15063);
or U17262 (N_17262,N_15970,N_15247);
or U17263 (N_17263,N_16155,N_16164);
xor U17264 (N_17264,N_15113,N_15953);
nand U17265 (N_17265,N_15361,N_16242);
and U17266 (N_17266,N_15512,N_16079);
and U17267 (N_17267,N_15063,N_15869);
and U17268 (N_17268,N_16060,N_15082);
xor U17269 (N_17269,N_15097,N_15207);
nor U17270 (N_17270,N_15830,N_16339);
nor U17271 (N_17271,N_15147,N_15067);
nand U17272 (N_17272,N_16420,N_15492);
or U17273 (N_17273,N_16351,N_16146);
nand U17274 (N_17274,N_15089,N_16057);
nand U17275 (N_17275,N_16361,N_15126);
xnor U17276 (N_17276,N_15207,N_15197);
or U17277 (N_17277,N_16144,N_16065);
xor U17278 (N_17278,N_15414,N_15053);
nor U17279 (N_17279,N_15716,N_15968);
and U17280 (N_17280,N_15234,N_15910);
or U17281 (N_17281,N_15635,N_16135);
and U17282 (N_17282,N_15263,N_16211);
nor U17283 (N_17283,N_15168,N_16378);
xor U17284 (N_17284,N_15191,N_15957);
xor U17285 (N_17285,N_15561,N_15135);
xor U17286 (N_17286,N_15560,N_16181);
and U17287 (N_17287,N_16412,N_15405);
or U17288 (N_17288,N_15655,N_15756);
or U17289 (N_17289,N_15412,N_16470);
and U17290 (N_17290,N_16473,N_15348);
or U17291 (N_17291,N_15055,N_16379);
or U17292 (N_17292,N_15956,N_15306);
nand U17293 (N_17293,N_15942,N_15890);
nand U17294 (N_17294,N_16380,N_15793);
nor U17295 (N_17295,N_15191,N_16110);
nand U17296 (N_17296,N_15546,N_16189);
nor U17297 (N_17297,N_16166,N_15994);
nor U17298 (N_17298,N_16002,N_15909);
or U17299 (N_17299,N_16475,N_15302);
nor U17300 (N_17300,N_15394,N_15093);
nor U17301 (N_17301,N_16109,N_15906);
xnor U17302 (N_17302,N_16217,N_15611);
xor U17303 (N_17303,N_15121,N_15729);
and U17304 (N_17304,N_15334,N_15575);
xor U17305 (N_17305,N_15953,N_15007);
nor U17306 (N_17306,N_16357,N_15268);
or U17307 (N_17307,N_16400,N_16386);
nor U17308 (N_17308,N_15346,N_16466);
nor U17309 (N_17309,N_15172,N_15502);
nand U17310 (N_17310,N_16314,N_15861);
or U17311 (N_17311,N_15994,N_15125);
and U17312 (N_17312,N_16258,N_15794);
nor U17313 (N_17313,N_15195,N_15197);
or U17314 (N_17314,N_15949,N_16447);
or U17315 (N_17315,N_15102,N_15260);
xnor U17316 (N_17316,N_16494,N_15037);
and U17317 (N_17317,N_16144,N_15076);
and U17318 (N_17318,N_16216,N_16069);
nand U17319 (N_17319,N_16155,N_15673);
or U17320 (N_17320,N_15007,N_16143);
nand U17321 (N_17321,N_15411,N_16497);
and U17322 (N_17322,N_16389,N_16084);
nand U17323 (N_17323,N_16026,N_15783);
nor U17324 (N_17324,N_15063,N_15062);
xnor U17325 (N_17325,N_15481,N_15388);
or U17326 (N_17326,N_15936,N_15956);
or U17327 (N_17327,N_16185,N_15475);
and U17328 (N_17328,N_16099,N_16156);
xnor U17329 (N_17329,N_16499,N_15947);
nand U17330 (N_17330,N_15219,N_15717);
and U17331 (N_17331,N_15924,N_15043);
nor U17332 (N_17332,N_16209,N_16409);
or U17333 (N_17333,N_15377,N_16305);
nor U17334 (N_17334,N_15523,N_16204);
nor U17335 (N_17335,N_15058,N_15850);
xor U17336 (N_17336,N_15850,N_15665);
or U17337 (N_17337,N_15681,N_15109);
nand U17338 (N_17338,N_16318,N_15072);
nor U17339 (N_17339,N_15507,N_15484);
nand U17340 (N_17340,N_16433,N_16190);
or U17341 (N_17341,N_15251,N_15714);
nor U17342 (N_17342,N_16029,N_16496);
or U17343 (N_17343,N_15416,N_16242);
and U17344 (N_17344,N_16248,N_16341);
xnor U17345 (N_17345,N_16003,N_15420);
or U17346 (N_17346,N_15205,N_15953);
nand U17347 (N_17347,N_16131,N_15731);
and U17348 (N_17348,N_16060,N_16193);
nor U17349 (N_17349,N_15133,N_15779);
xor U17350 (N_17350,N_15177,N_16401);
nand U17351 (N_17351,N_16241,N_15931);
nor U17352 (N_17352,N_15160,N_15937);
or U17353 (N_17353,N_15412,N_15975);
nand U17354 (N_17354,N_15329,N_15745);
nand U17355 (N_17355,N_15302,N_15752);
and U17356 (N_17356,N_15113,N_16337);
nor U17357 (N_17357,N_15435,N_15809);
xnor U17358 (N_17358,N_16178,N_16477);
nand U17359 (N_17359,N_16344,N_16366);
or U17360 (N_17360,N_15512,N_16032);
nand U17361 (N_17361,N_15870,N_15172);
nor U17362 (N_17362,N_16250,N_15505);
or U17363 (N_17363,N_16459,N_15223);
or U17364 (N_17364,N_16449,N_16276);
nor U17365 (N_17365,N_16404,N_16427);
xor U17366 (N_17366,N_16132,N_15653);
nor U17367 (N_17367,N_15963,N_15242);
nand U17368 (N_17368,N_15693,N_16379);
nand U17369 (N_17369,N_15908,N_15323);
xor U17370 (N_17370,N_15624,N_16449);
nand U17371 (N_17371,N_16487,N_15791);
or U17372 (N_17372,N_15913,N_16498);
or U17373 (N_17373,N_15564,N_16359);
xor U17374 (N_17374,N_16337,N_16253);
or U17375 (N_17375,N_16205,N_15292);
xor U17376 (N_17376,N_16041,N_16027);
nand U17377 (N_17377,N_16319,N_15383);
nor U17378 (N_17378,N_15322,N_16208);
and U17379 (N_17379,N_15376,N_16140);
nand U17380 (N_17380,N_15685,N_15642);
or U17381 (N_17381,N_15938,N_15446);
xnor U17382 (N_17382,N_15001,N_15692);
xor U17383 (N_17383,N_15326,N_16472);
and U17384 (N_17384,N_15615,N_16376);
nand U17385 (N_17385,N_16179,N_15596);
nor U17386 (N_17386,N_15666,N_15680);
and U17387 (N_17387,N_16312,N_15573);
xor U17388 (N_17388,N_15352,N_15690);
and U17389 (N_17389,N_15338,N_16090);
xnor U17390 (N_17390,N_16483,N_15080);
nand U17391 (N_17391,N_15920,N_16482);
nor U17392 (N_17392,N_16402,N_16170);
nor U17393 (N_17393,N_16397,N_15030);
xnor U17394 (N_17394,N_15697,N_15128);
nor U17395 (N_17395,N_15042,N_15314);
xor U17396 (N_17396,N_16160,N_15092);
or U17397 (N_17397,N_16440,N_15856);
nand U17398 (N_17398,N_15400,N_15201);
nor U17399 (N_17399,N_15274,N_15458);
and U17400 (N_17400,N_15581,N_15823);
nor U17401 (N_17401,N_15450,N_15602);
and U17402 (N_17402,N_16467,N_15421);
nand U17403 (N_17403,N_16393,N_16251);
or U17404 (N_17404,N_15451,N_16122);
xnor U17405 (N_17405,N_16170,N_15726);
xor U17406 (N_17406,N_16491,N_15523);
xnor U17407 (N_17407,N_16163,N_15003);
and U17408 (N_17408,N_15727,N_15360);
nor U17409 (N_17409,N_15123,N_15741);
or U17410 (N_17410,N_15969,N_16478);
or U17411 (N_17411,N_15341,N_15432);
xor U17412 (N_17412,N_16233,N_15878);
nand U17413 (N_17413,N_15803,N_15054);
nor U17414 (N_17414,N_15558,N_16462);
and U17415 (N_17415,N_15350,N_15338);
nor U17416 (N_17416,N_15821,N_16264);
nand U17417 (N_17417,N_15239,N_15881);
or U17418 (N_17418,N_16397,N_16036);
xor U17419 (N_17419,N_16202,N_15615);
nand U17420 (N_17420,N_15344,N_16123);
nor U17421 (N_17421,N_16425,N_15016);
xor U17422 (N_17422,N_15849,N_16137);
xnor U17423 (N_17423,N_16182,N_15739);
or U17424 (N_17424,N_15548,N_15115);
nor U17425 (N_17425,N_15425,N_15506);
xor U17426 (N_17426,N_15706,N_15776);
nand U17427 (N_17427,N_16387,N_15007);
or U17428 (N_17428,N_15688,N_16422);
nor U17429 (N_17429,N_15932,N_15814);
and U17430 (N_17430,N_15225,N_15544);
xor U17431 (N_17431,N_15050,N_15901);
nor U17432 (N_17432,N_16117,N_16059);
nand U17433 (N_17433,N_16397,N_16215);
and U17434 (N_17434,N_15813,N_15093);
nand U17435 (N_17435,N_15792,N_16463);
nand U17436 (N_17436,N_15673,N_15553);
xnor U17437 (N_17437,N_16324,N_15290);
nand U17438 (N_17438,N_15115,N_16409);
nor U17439 (N_17439,N_15231,N_15510);
and U17440 (N_17440,N_15645,N_15130);
nand U17441 (N_17441,N_15049,N_15669);
nand U17442 (N_17442,N_15218,N_15506);
or U17443 (N_17443,N_15555,N_15518);
xnor U17444 (N_17444,N_16230,N_15102);
or U17445 (N_17445,N_15152,N_15500);
nor U17446 (N_17446,N_15164,N_15939);
and U17447 (N_17447,N_16241,N_16099);
nand U17448 (N_17448,N_15117,N_15514);
nand U17449 (N_17449,N_15261,N_15365);
nor U17450 (N_17450,N_16421,N_15753);
nor U17451 (N_17451,N_15648,N_15772);
or U17452 (N_17452,N_15003,N_15349);
and U17453 (N_17453,N_15496,N_16413);
or U17454 (N_17454,N_16259,N_15765);
nand U17455 (N_17455,N_15988,N_16146);
nand U17456 (N_17456,N_15370,N_15722);
nand U17457 (N_17457,N_15960,N_16130);
or U17458 (N_17458,N_15028,N_15075);
nor U17459 (N_17459,N_16424,N_16415);
nor U17460 (N_17460,N_15790,N_16314);
and U17461 (N_17461,N_16406,N_15580);
or U17462 (N_17462,N_16232,N_15561);
or U17463 (N_17463,N_15081,N_15324);
or U17464 (N_17464,N_15408,N_15698);
or U17465 (N_17465,N_15528,N_15369);
nor U17466 (N_17466,N_16342,N_15518);
and U17467 (N_17467,N_16198,N_16168);
nand U17468 (N_17468,N_16176,N_15389);
nor U17469 (N_17469,N_15913,N_16064);
xor U17470 (N_17470,N_16130,N_15834);
xnor U17471 (N_17471,N_15450,N_15662);
and U17472 (N_17472,N_15368,N_15507);
or U17473 (N_17473,N_15045,N_15653);
nand U17474 (N_17474,N_15213,N_16402);
xor U17475 (N_17475,N_15730,N_16498);
and U17476 (N_17476,N_15973,N_16264);
xnor U17477 (N_17477,N_15542,N_16385);
nand U17478 (N_17478,N_16192,N_16166);
or U17479 (N_17479,N_15323,N_15171);
or U17480 (N_17480,N_16252,N_15563);
or U17481 (N_17481,N_15355,N_16159);
nor U17482 (N_17482,N_15882,N_15249);
nor U17483 (N_17483,N_15497,N_15001);
nor U17484 (N_17484,N_15124,N_16471);
and U17485 (N_17485,N_15576,N_15353);
xor U17486 (N_17486,N_15052,N_15856);
nand U17487 (N_17487,N_15276,N_15900);
and U17488 (N_17488,N_15030,N_15830);
nor U17489 (N_17489,N_15104,N_15611);
and U17490 (N_17490,N_15017,N_16443);
or U17491 (N_17491,N_15936,N_15202);
or U17492 (N_17492,N_15051,N_15507);
nand U17493 (N_17493,N_16200,N_15675);
nor U17494 (N_17494,N_16089,N_15155);
and U17495 (N_17495,N_15806,N_15084);
and U17496 (N_17496,N_16141,N_15762);
and U17497 (N_17497,N_16076,N_16327);
and U17498 (N_17498,N_16211,N_15281);
and U17499 (N_17499,N_15535,N_16399);
and U17500 (N_17500,N_16245,N_15143);
nor U17501 (N_17501,N_15402,N_16387);
and U17502 (N_17502,N_15012,N_15555);
and U17503 (N_17503,N_16499,N_15627);
nor U17504 (N_17504,N_15056,N_16185);
xor U17505 (N_17505,N_15123,N_15507);
and U17506 (N_17506,N_15945,N_15560);
or U17507 (N_17507,N_15208,N_15663);
xor U17508 (N_17508,N_16199,N_15402);
xor U17509 (N_17509,N_15071,N_16262);
nand U17510 (N_17510,N_15679,N_15654);
and U17511 (N_17511,N_15637,N_15616);
and U17512 (N_17512,N_16246,N_15705);
or U17513 (N_17513,N_15013,N_15137);
and U17514 (N_17514,N_15145,N_15118);
nor U17515 (N_17515,N_16389,N_16062);
nor U17516 (N_17516,N_16319,N_15721);
xnor U17517 (N_17517,N_16449,N_16091);
and U17518 (N_17518,N_16379,N_15586);
nand U17519 (N_17519,N_15385,N_15895);
nand U17520 (N_17520,N_15914,N_15056);
nand U17521 (N_17521,N_15237,N_15721);
or U17522 (N_17522,N_16194,N_16060);
nor U17523 (N_17523,N_15588,N_15582);
nor U17524 (N_17524,N_15883,N_15810);
nand U17525 (N_17525,N_15910,N_15261);
nor U17526 (N_17526,N_15047,N_16052);
nor U17527 (N_17527,N_16291,N_16436);
or U17528 (N_17528,N_15243,N_16145);
and U17529 (N_17529,N_16225,N_15697);
nor U17530 (N_17530,N_15545,N_15185);
xor U17531 (N_17531,N_16330,N_15673);
nand U17532 (N_17532,N_15275,N_16164);
nor U17533 (N_17533,N_15808,N_16414);
and U17534 (N_17534,N_15756,N_15707);
nand U17535 (N_17535,N_16265,N_15121);
nand U17536 (N_17536,N_16218,N_15985);
nor U17537 (N_17537,N_15137,N_15831);
nor U17538 (N_17538,N_15164,N_15395);
xor U17539 (N_17539,N_15238,N_16474);
nand U17540 (N_17540,N_15737,N_15251);
nand U17541 (N_17541,N_15805,N_15382);
and U17542 (N_17542,N_16264,N_15015);
xnor U17543 (N_17543,N_16263,N_16257);
nor U17544 (N_17544,N_15403,N_15575);
and U17545 (N_17545,N_16470,N_15699);
and U17546 (N_17546,N_15885,N_16177);
and U17547 (N_17547,N_15490,N_15296);
nand U17548 (N_17548,N_16209,N_15238);
or U17549 (N_17549,N_15179,N_15706);
nor U17550 (N_17550,N_15682,N_15478);
nor U17551 (N_17551,N_16377,N_15831);
or U17552 (N_17552,N_15019,N_15871);
nand U17553 (N_17553,N_15057,N_15095);
or U17554 (N_17554,N_15210,N_15506);
nand U17555 (N_17555,N_15198,N_15022);
and U17556 (N_17556,N_16150,N_15297);
and U17557 (N_17557,N_15053,N_16395);
and U17558 (N_17558,N_15465,N_16168);
nand U17559 (N_17559,N_15543,N_16234);
or U17560 (N_17560,N_15876,N_15850);
and U17561 (N_17561,N_15225,N_15618);
and U17562 (N_17562,N_15567,N_15066);
nor U17563 (N_17563,N_16080,N_15353);
nand U17564 (N_17564,N_15147,N_15298);
nor U17565 (N_17565,N_15901,N_15805);
or U17566 (N_17566,N_15764,N_16046);
nand U17567 (N_17567,N_15087,N_15026);
nor U17568 (N_17568,N_16082,N_15799);
or U17569 (N_17569,N_15659,N_15575);
or U17570 (N_17570,N_16338,N_15747);
and U17571 (N_17571,N_15788,N_16380);
or U17572 (N_17572,N_15832,N_15691);
xor U17573 (N_17573,N_15445,N_16173);
nor U17574 (N_17574,N_15947,N_16123);
and U17575 (N_17575,N_16121,N_15783);
and U17576 (N_17576,N_15774,N_16244);
nor U17577 (N_17577,N_15060,N_16325);
or U17578 (N_17578,N_16395,N_15331);
xor U17579 (N_17579,N_16441,N_15760);
nor U17580 (N_17580,N_15095,N_15637);
or U17581 (N_17581,N_16037,N_15592);
nor U17582 (N_17582,N_15702,N_15264);
nor U17583 (N_17583,N_16490,N_15456);
and U17584 (N_17584,N_15201,N_15094);
and U17585 (N_17585,N_15080,N_15682);
nor U17586 (N_17586,N_16193,N_15058);
xnor U17587 (N_17587,N_15071,N_16259);
and U17588 (N_17588,N_16159,N_15911);
and U17589 (N_17589,N_15764,N_16140);
nand U17590 (N_17590,N_16149,N_15601);
or U17591 (N_17591,N_15918,N_15068);
and U17592 (N_17592,N_15969,N_15877);
or U17593 (N_17593,N_15599,N_15407);
or U17594 (N_17594,N_15102,N_16486);
or U17595 (N_17595,N_16455,N_15693);
nor U17596 (N_17596,N_16062,N_15939);
and U17597 (N_17597,N_15667,N_15085);
nor U17598 (N_17598,N_15476,N_15638);
or U17599 (N_17599,N_15693,N_15664);
or U17600 (N_17600,N_15322,N_16044);
nand U17601 (N_17601,N_16219,N_15966);
xnor U17602 (N_17602,N_15498,N_15852);
xnor U17603 (N_17603,N_15070,N_16063);
or U17604 (N_17604,N_16282,N_16001);
nand U17605 (N_17605,N_15432,N_15575);
xor U17606 (N_17606,N_16170,N_15070);
or U17607 (N_17607,N_15254,N_15923);
and U17608 (N_17608,N_15507,N_15057);
nand U17609 (N_17609,N_15285,N_16252);
and U17610 (N_17610,N_15296,N_15784);
and U17611 (N_17611,N_15967,N_15149);
nor U17612 (N_17612,N_15477,N_15534);
or U17613 (N_17613,N_16281,N_16224);
nor U17614 (N_17614,N_15944,N_15891);
nor U17615 (N_17615,N_16295,N_15637);
xor U17616 (N_17616,N_16347,N_16052);
nand U17617 (N_17617,N_15101,N_15717);
xor U17618 (N_17618,N_16188,N_16001);
and U17619 (N_17619,N_15282,N_15369);
nor U17620 (N_17620,N_16067,N_15232);
or U17621 (N_17621,N_16227,N_16020);
nor U17622 (N_17622,N_16043,N_15656);
or U17623 (N_17623,N_15927,N_15929);
nor U17624 (N_17624,N_15511,N_15647);
and U17625 (N_17625,N_16495,N_16365);
or U17626 (N_17626,N_16126,N_15598);
nand U17627 (N_17627,N_15781,N_15248);
and U17628 (N_17628,N_15935,N_15117);
xnor U17629 (N_17629,N_15768,N_15829);
and U17630 (N_17630,N_15734,N_16366);
and U17631 (N_17631,N_15974,N_15091);
or U17632 (N_17632,N_15886,N_15238);
nor U17633 (N_17633,N_16039,N_16318);
and U17634 (N_17634,N_16232,N_16051);
xor U17635 (N_17635,N_15772,N_16456);
nor U17636 (N_17636,N_15650,N_16228);
or U17637 (N_17637,N_16403,N_16255);
and U17638 (N_17638,N_15715,N_16228);
nor U17639 (N_17639,N_15119,N_16307);
xnor U17640 (N_17640,N_16235,N_15111);
nor U17641 (N_17641,N_15987,N_15799);
nand U17642 (N_17642,N_15225,N_15688);
and U17643 (N_17643,N_16361,N_16112);
nor U17644 (N_17644,N_15825,N_16122);
nor U17645 (N_17645,N_15343,N_15757);
and U17646 (N_17646,N_15166,N_15946);
nor U17647 (N_17647,N_16190,N_15155);
nand U17648 (N_17648,N_15499,N_15091);
nand U17649 (N_17649,N_16002,N_15587);
nor U17650 (N_17650,N_16305,N_15481);
xor U17651 (N_17651,N_16099,N_15428);
or U17652 (N_17652,N_15461,N_15540);
xor U17653 (N_17653,N_15071,N_16420);
xnor U17654 (N_17654,N_15306,N_16374);
and U17655 (N_17655,N_15563,N_16249);
and U17656 (N_17656,N_15146,N_16383);
nor U17657 (N_17657,N_15659,N_15681);
nor U17658 (N_17658,N_15507,N_15300);
nor U17659 (N_17659,N_15393,N_15733);
nand U17660 (N_17660,N_15800,N_15653);
nand U17661 (N_17661,N_15695,N_15963);
and U17662 (N_17662,N_16288,N_15626);
or U17663 (N_17663,N_15706,N_15251);
or U17664 (N_17664,N_15485,N_16347);
or U17665 (N_17665,N_15351,N_15659);
nand U17666 (N_17666,N_16233,N_15024);
and U17667 (N_17667,N_15805,N_15848);
nand U17668 (N_17668,N_15857,N_15089);
or U17669 (N_17669,N_15047,N_15717);
nand U17670 (N_17670,N_15775,N_15982);
xnor U17671 (N_17671,N_15553,N_15741);
and U17672 (N_17672,N_16444,N_16114);
xnor U17673 (N_17673,N_15553,N_15762);
or U17674 (N_17674,N_15371,N_16429);
nor U17675 (N_17675,N_15942,N_15377);
or U17676 (N_17676,N_15500,N_15966);
and U17677 (N_17677,N_15921,N_15924);
or U17678 (N_17678,N_15501,N_15025);
and U17679 (N_17679,N_15600,N_15156);
nor U17680 (N_17680,N_15547,N_15114);
nor U17681 (N_17681,N_15350,N_15862);
or U17682 (N_17682,N_16409,N_15553);
nand U17683 (N_17683,N_15244,N_15860);
and U17684 (N_17684,N_15855,N_15600);
or U17685 (N_17685,N_15924,N_15530);
or U17686 (N_17686,N_16474,N_15587);
nand U17687 (N_17687,N_15545,N_15183);
or U17688 (N_17688,N_15426,N_15154);
xor U17689 (N_17689,N_15265,N_16494);
nand U17690 (N_17690,N_15866,N_16450);
xnor U17691 (N_17691,N_16383,N_16205);
nand U17692 (N_17692,N_16006,N_16359);
nand U17693 (N_17693,N_16167,N_15940);
xnor U17694 (N_17694,N_15640,N_15360);
xnor U17695 (N_17695,N_15045,N_15774);
or U17696 (N_17696,N_15944,N_16234);
and U17697 (N_17697,N_15202,N_15277);
and U17698 (N_17698,N_15810,N_15422);
and U17699 (N_17699,N_16365,N_16453);
xor U17700 (N_17700,N_15783,N_15805);
or U17701 (N_17701,N_15176,N_15319);
and U17702 (N_17702,N_16244,N_16411);
and U17703 (N_17703,N_15101,N_15467);
xnor U17704 (N_17704,N_15612,N_15080);
or U17705 (N_17705,N_15199,N_15899);
and U17706 (N_17706,N_15307,N_15969);
and U17707 (N_17707,N_15422,N_16142);
xnor U17708 (N_17708,N_16184,N_15909);
nand U17709 (N_17709,N_16012,N_15651);
and U17710 (N_17710,N_15901,N_15668);
and U17711 (N_17711,N_15379,N_15554);
nand U17712 (N_17712,N_16093,N_15776);
nor U17713 (N_17713,N_15216,N_15014);
xnor U17714 (N_17714,N_16211,N_16321);
and U17715 (N_17715,N_15376,N_16337);
nand U17716 (N_17716,N_15933,N_15673);
xnor U17717 (N_17717,N_15906,N_15883);
xnor U17718 (N_17718,N_15308,N_16399);
and U17719 (N_17719,N_15108,N_15420);
or U17720 (N_17720,N_16122,N_15494);
nor U17721 (N_17721,N_15366,N_15917);
xnor U17722 (N_17722,N_15549,N_15644);
and U17723 (N_17723,N_15020,N_15253);
or U17724 (N_17724,N_15065,N_16440);
nor U17725 (N_17725,N_15632,N_16359);
xnor U17726 (N_17726,N_16175,N_15360);
xnor U17727 (N_17727,N_16272,N_15181);
or U17728 (N_17728,N_15038,N_15406);
nor U17729 (N_17729,N_15355,N_15096);
nor U17730 (N_17730,N_15624,N_15198);
nor U17731 (N_17731,N_15079,N_16080);
nand U17732 (N_17732,N_15244,N_16209);
and U17733 (N_17733,N_15054,N_15141);
xor U17734 (N_17734,N_15978,N_15904);
xnor U17735 (N_17735,N_15014,N_16096);
nand U17736 (N_17736,N_15958,N_15327);
xor U17737 (N_17737,N_16138,N_15337);
and U17738 (N_17738,N_15767,N_15487);
nand U17739 (N_17739,N_15804,N_16290);
nor U17740 (N_17740,N_15179,N_15366);
or U17741 (N_17741,N_15698,N_15159);
xnor U17742 (N_17742,N_16434,N_15095);
nand U17743 (N_17743,N_16377,N_15363);
nand U17744 (N_17744,N_16316,N_16287);
or U17745 (N_17745,N_15535,N_15512);
nor U17746 (N_17746,N_15513,N_16137);
and U17747 (N_17747,N_16131,N_16087);
and U17748 (N_17748,N_15341,N_15009);
and U17749 (N_17749,N_15064,N_16057);
nand U17750 (N_17750,N_15525,N_16342);
nor U17751 (N_17751,N_16164,N_16458);
xnor U17752 (N_17752,N_15737,N_15369);
nand U17753 (N_17753,N_16440,N_15708);
and U17754 (N_17754,N_15760,N_15315);
or U17755 (N_17755,N_15069,N_15009);
nor U17756 (N_17756,N_15792,N_16004);
xor U17757 (N_17757,N_15867,N_15706);
nand U17758 (N_17758,N_15699,N_15902);
xnor U17759 (N_17759,N_15520,N_16036);
and U17760 (N_17760,N_15207,N_16485);
and U17761 (N_17761,N_15961,N_16175);
and U17762 (N_17762,N_15756,N_15847);
nand U17763 (N_17763,N_15381,N_15242);
xnor U17764 (N_17764,N_15390,N_15839);
and U17765 (N_17765,N_15874,N_16320);
xor U17766 (N_17766,N_15534,N_16334);
xnor U17767 (N_17767,N_15665,N_15160);
nand U17768 (N_17768,N_15959,N_16448);
nor U17769 (N_17769,N_15001,N_15391);
xnor U17770 (N_17770,N_15959,N_15089);
nand U17771 (N_17771,N_15774,N_15746);
nand U17772 (N_17772,N_15410,N_16428);
nor U17773 (N_17773,N_15175,N_15837);
xnor U17774 (N_17774,N_16071,N_15757);
and U17775 (N_17775,N_16284,N_15702);
nand U17776 (N_17776,N_15429,N_16032);
nand U17777 (N_17777,N_15967,N_15134);
nand U17778 (N_17778,N_15954,N_15113);
or U17779 (N_17779,N_15993,N_15522);
nand U17780 (N_17780,N_15042,N_15377);
and U17781 (N_17781,N_15181,N_15365);
or U17782 (N_17782,N_15398,N_15842);
nor U17783 (N_17783,N_16477,N_16092);
nor U17784 (N_17784,N_16404,N_15703);
and U17785 (N_17785,N_15181,N_15820);
or U17786 (N_17786,N_15391,N_15075);
or U17787 (N_17787,N_16417,N_15613);
nand U17788 (N_17788,N_16266,N_15939);
nand U17789 (N_17789,N_16198,N_15988);
xnor U17790 (N_17790,N_16478,N_15572);
nor U17791 (N_17791,N_16111,N_16186);
xor U17792 (N_17792,N_15565,N_16396);
xnor U17793 (N_17793,N_15179,N_15018);
or U17794 (N_17794,N_16208,N_16342);
or U17795 (N_17795,N_15837,N_16418);
nand U17796 (N_17796,N_16203,N_16460);
and U17797 (N_17797,N_15804,N_15491);
xnor U17798 (N_17798,N_15766,N_15123);
xor U17799 (N_17799,N_16224,N_15916);
xnor U17800 (N_17800,N_16393,N_15438);
or U17801 (N_17801,N_15805,N_15732);
or U17802 (N_17802,N_16388,N_15144);
or U17803 (N_17803,N_16433,N_15745);
or U17804 (N_17804,N_16314,N_16076);
xnor U17805 (N_17805,N_15486,N_15959);
nor U17806 (N_17806,N_15995,N_16119);
and U17807 (N_17807,N_15969,N_16485);
nand U17808 (N_17808,N_16075,N_15729);
and U17809 (N_17809,N_15139,N_16416);
nand U17810 (N_17810,N_15082,N_16367);
nand U17811 (N_17811,N_15137,N_15640);
nor U17812 (N_17812,N_15102,N_15842);
and U17813 (N_17813,N_16108,N_16332);
xnor U17814 (N_17814,N_15799,N_16451);
and U17815 (N_17815,N_16116,N_16026);
or U17816 (N_17816,N_16486,N_16489);
nor U17817 (N_17817,N_15832,N_15095);
and U17818 (N_17818,N_16465,N_15653);
or U17819 (N_17819,N_15466,N_15682);
and U17820 (N_17820,N_15292,N_15706);
nor U17821 (N_17821,N_15554,N_16459);
and U17822 (N_17822,N_15797,N_15456);
or U17823 (N_17823,N_16320,N_16453);
or U17824 (N_17824,N_16120,N_15610);
or U17825 (N_17825,N_15357,N_16131);
or U17826 (N_17826,N_16248,N_15891);
nor U17827 (N_17827,N_16124,N_15641);
nand U17828 (N_17828,N_15366,N_15922);
and U17829 (N_17829,N_15705,N_16211);
or U17830 (N_17830,N_16066,N_16490);
nor U17831 (N_17831,N_15833,N_16001);
and U17832 (N_17832,N_15346,N_16338);
xor U17833 (N_17833,N_16160,N_16304);
or U17834 (N_17834,N_16188,N_15244);
or U17835 (N_17835,N_15195,N_15674);
nor U17836 (N_17836,N_16242,N_15807);
nor U17837 (N_17837,N_16440,N_16387);
xnor U17838 (N_17838,N_16318,N_15147);
nand U17839 (N_17839,N_15738,N_16024);
xnor U17840 (N_17840,N_16285,N_16250);
and U17841 (N_17841,N_15294,N_16269);
nor U17842 (N_17842,N_16354,N_16369);
xor U17843 (N_17843,N_16288,N_16385);
or U17844 (N_17844,N_15868,N_15497);
and U17845 (N_17845,N_16149,N_15719);
nand U17846 (N_17846,N_15849,N_16325);
xnor U17847 (N_17847,N_16380,N_15926);
and U17848 (N_17848,N_15115,N_15008);
xnor U17849 (N_17849,N_16233,N_15349);
nand U17850 (N_17850,N_15757,N_15133);
or U17851 (N_17851,N_15413,N_15132);
and U17852 (N_17852,N_16396,N_16350);
nor U17853 (N_17853,N_16426,N_15388);
nand U17854 (N_17854,N_16462,N_15238);
xor U17855 (N_17855,N_15907,N_15306);
and U17856 (N_17856,N_16208,N_15915);
and U17857 (N_17857,N_15287,N_15005);
nand U17858 (N_17858,N_15573,N_15366);
nand U17859 (N_17859,N_15558,N_15465);
nand U17860 (N_17860,N_16474,N_15716);
nor U17861 (N_17861,N_15432,N_16204);
nor U17862 (N_17862,N_16364,N_15073);
and U17863 (N_17863,N_15741,N_15844);
or U17864 (N_17864,N_15452,N_15537);
and U17865 (N_17865,N_15479,N_16471);
and U17866 (N_17866,N_15722,N_15153);
nand U17867 (N_17867,N_15839,N_16204);
or U17868 (N_17868,N_15348,N_16209);
and U17869 (N_17869,N_16451,N_15070);
nor U17870 (N_17870,N_15426,N_15885);
or U17871 (N_17871,N_16184,N_15698);
and U17872 (N_17872,N_15218,N_16365);
and U17873 (N_17873,N_16122,N_16029);
nand U17874 (N_17874,N_15302,N_15275);
nor U17875 (N_17875,N_16393,N_15950);
or U17876 (N_17876,N_15939,N_15163);
nor U17877 (N_17877,N_15625,N_15158);
and U17878 (N_17878,N_16262,N_16271);
xnor U17879 (N_17879,N_15926,N_16282);
and U17880 (N_17880,N_15080,N_16011);
xnor U17881 (N_17881,N_15344,N_16186);
xnor U17882 (N_17882,N_15455,N_16293);
and U17883 (N_17883,N_15853,N_16413);
nand U17884 (N_17884,N_15562,N_15507);
nand U17885 (N_17885,N_16006,N_15386);
and U17886 (N_17886,N_15883,N_15715);
or U17887 (N_17887,N_16120,N_15358);
nand U17888 (N_17888,N_15680,N_15290);
nand U17889 (N_17889,N_16204,N_15284);
xor U17890 (N_17890,N_15915,N_15373);
nand U17891 (N_17891,N_16074,N_15901);
or U17892 (N_17892,N_15621,N_15250);
or U17893 (N_17893,N_16042,N_16172);
and U17894 (N_17894,N_15804,N_15445);
and U17895 (N_17895,N_15245,N_15428);
and U17896 (N_17896,N_15002,N_16002);
nor U17897 (N_17897,N_15790,N_15504);
nand U17898 (N_17898,N_15506,N_16391);
nor U17899 (N_17899,N_16051,N_15299);
xnor U17900 (N_17900,N_15720,N_15565);
nand U17901 (N_17901,N_16474,N_16082);
nand U17902 (N_17902,N_15532,N_15151);
xnor U17903 (N_17903,N_15434,N_15355);
nor U17904 (N_17904,N_16238,N_15539);
or U17905 (N_17905,N_16347,N_15567);
nor U17906 (N_17906,N_15591,N_16057);
nor U17907 (N_17907,N_15764,N_16440);
xnor U17908 (N_17908,N_16315,N_16097);
nand U17909 (N_17909,N_16129,N_15734);
nand U17910 (N_17910,N_15991,N_16089);
nor U17911 (N_17911,N_16339,N_16007);
or U17912 (N_17912,N_15921,N_15975);
or U17913 (N_17913,N_15760,N_15291);
nor U17914 (N_17914,N_16000,N_15582);
xnor U17915 (N_17915,N_15656,N_16291);
xor U17916 (N_17916,N_16030,N_15110);
and U17917 (N_17917,N_15910,N_16287);
or U17918 (N_17918,N_15757,N_15767);
nand U17919 (N_17919,N_16115,N_15724);
or U17920 (N_17920,N_16141,N_15264);
nor U17921 (N_17921,N_15574,N_16049);
nand U17922 (N_17922,N_15861,N_15304);
or U17923 (N_17923,N_16021,N_15110);
or U17924 (N_17924,N_16022,N_16416);
nor U17925 (N_17925,N_15380,N_15263);
or U17926 (N_17926,N_15917,N_15836);
or U17927 (N_17927,N_16092,N_16451);
xnor U17928 (N_17928,N_15553,N_15693);
nor U17929 (N_17929,N_15503,N_15208);
and U17930 (N_17930,N_16402,N_16278);
and U17931 (N_17931,N_16454,N_16301);
or U17932 (N_17932,N_15376,N_15201);
xor U17933 (N_17933,N_16215,N_16161);
xnor U17934 (N_17934,N_15875,N_16355);
nand U17935 (N_17935,N_15654,N_15830);
and U17936 (N_17936,N_15821,N_15562);
nand U17937 (N_17937,N_16186,N_15508);
and U17938 (N_17938,N_15152,N_15192);
nand U17939 (N_17939,N_15195,N_16011);
or U17940 (N_17940,N_15256,N_15780);
xor U17941 (N_17941,N_15544,N_16085);
nor U17942 (N_17942,N_16271,N_16100);
nand U17943 (N_17943,N_15686,N_16272);
or U17944 (N_17944,N_15414,N_15104);
nand U17945 (N_17945,N_15507,N_15514);
nor U17946 (N_17946,N_16151,N_16312);
nand U17947 (N_17947,N_16268,N_15540);
nand U17948 (N_17948,N_15466,N_15910);
xor U17949 (N_17949,N_15860,N_15427);
and U17950 (N_17950,N_15704,N_15880);
nand U17951 (N_17951,N_16215,N_15440);
and U17952 (N_17952,N_16396,N_16235);
nand U17953 (N_17953,N_16089,N_16031);
and U17954 (N_17954,N_15061,N_15958);
xor U17955 (N_17955,N_15642,N_16100);
or U17956 (N_17956,N_16208,N_15957);
nor U17957 (N_17957,N_16327,N_16268);
and U17958 (N_17958,N_15869,N_15149);
or U17959 (N_17959,N_15454,N_15917);
nor U17960 (N_17960,N_15032,N_16130);
nor U17961 (N_17961,N_15567,N_15706);
or U17962 (N_17962,N_15855,N_16426);
xnor U17963 (N_17963,N_15669,N_15528);
nand U17964 (N_17964,N_15602,N_16454);
and U17965 (N_17965,N_15762,N_16015);
and U17966 (N_17966,N_15835,N_15872);
or U17967 (N_17967,N_15854,N_15142);
nor U17968 (N_17968,N_15014,N_15712);
nor U17969 (N_17969,N_15903,N_15777);
nand U17970 (N_17970,N_15646,N_15813);
nor U17971 (N_17971,N_16327,N_16435);
and U17972 (N_17972,N_15158,N_15413);
nand U17973 (N_17973,N_16352,N_16305);
xnor U17974 (N_17974,N_15469,N_15715);
xnor U17975 (N_17975,N_15749,N_15013);
nand U17976 (N_17976,N_16471,N_15659);
nor U17977 (N_17977,N_16341,N_15371);
nand U17978 (N_17978,N_16034,N_16457);
or U17979 (N_17979,N_15605,N_15691);
nand U17980 (N_17980,N_16344,N_15958);
nor U17981 (N_17981,N_16114,N_15536);
xor U17982 (N_17982,N_15485,N_15652);
nand U17983 (N_17983,N_15598,N_16363);
and U17984 (N_17984,N_16071,N_15572);
nand U17985 (N_17985,N_15193,N_16411);
nand U17986 (N_17986,N_15277,N_15640);
or U17987 (N_17987,N_15445,N_16181);
xor U17988 (N_17988,N_16041,N_15496);
xnor U17989 (N_17989,N_15591,N_15993);
xor U17990 (N_17990,N_15976,N_15767);
xnor U17991 (N_17991,N_15947,N_15390);
or U17992 (N_17992,N_15750,N_16053);
nand U17993 (N_17993,N_15210,N_16315);
and U17994 (N_17994,N_15172,N_15540);
xor U17995 (N_17995,N_16397,N_15228);
or U17996 (N_17996,N_16204,N_15913);
or U17997 (N_17997,N_15043,N_15280);
and U17998 (N_17998,N_15275,N_15068);
or U17999 (N_17999,N_15961,N_15455);
xor U18000 (N_18000,N_16589,N_16770);
xor U18001 (N_18001,N_16914,N_17770);
and U18002 (N_18002,N_17390,N_17794);
and U18003 (N_18003,N_17829,N_17881);
and U18004 (N_18004,N_16663,N_17949);
nor U18005 (N_18005,N_17907,N_17352);
xnor U18006 (N_18006,N_16524,N_17162);
and U18007 (N_18007,N_17408,N_17825);
nor U18008 (N_18008,N_16968,N_16884);
xnor U18009 (N_18009,N_16941,N_17261);
or U18010 (N_18010,N_17207,N_17773);
or U18011 (N_18011,N_17266,N_17220);
nand U18012 (N_18012,N_16995,N_17014);
nand U18013 (N_18013,N_17425,N_17602);
nor U18014 (N_18014,N_16961,N_17945);
nand U18015 (N_18015,N_17336,N_17995);
nor U18016 (N_18016,N_16763,N_17037);
nand U18017 (N_18017,N_16579,N_16774);
and U18018 (N_18018,N_16544,N_17484);
nor U18019 (N_18019,N_17099,N_16803);
and U18020 (N_18020,N_16867,N_16890);
nor U18021 (N_18021,N_16925,N_17096);
xnor U18022 (N_18022,N_16768,N_17471);
or U18023 (N_18023,N_17447,N_17004);
or U18024 (N_18024,N_16590,N_17255);
nand U18025 (N_18025,N_16719,N_17275);
xnor U18026 (N_18026,N_17653,N_17195);
nor U18027 (N_18027,N_17637,N_17520);
and U18028 (N_18028,N_17790,N_16892);
and U18029 (N_18029,N_17048,N_17380);
or U18030 (N_18030,N_17963,N_16906);
and U18031 (N_18031,N_17397,N_16611);
and U18032 (N_18032,N_17572,N_17280);
nor U18033 (N_18033,N_16536,N_16607);
nor U18034 (N_18034,N_17036,N_17596);
xor U18035 (N_18035,N_17574,N_16622);
and U18036 (N_18036,N_17118,N_17171);
nand U18037 (N_18037,N_17712,N_17548);
and U18038 (N_18038,N_17553,N_17312);
nor U18039 (N_18039,N_17922,N_16564);
and U18040 (N_18040,N_17507,N_17353);
or U18041 (N_18041,N_17231,N_16862);
nand U18042 (N_18042,N_16554,N_16736);
nand U18043 (N_18043,N_17369,N_17143);
nor U18044 (N_18044,N_16828,N_17796);
nor U18045 (N_18045,N_17102,N_17466);
and U18046 (N_18046,N_17684,N_16682);
nor U18047 (N_18047,N_16819,N_17402);
nor U18048 (N_18048,N_17492,N_17209);
or U18049 (N_18049,N_16658,N_16636);
or U18050 (N_18050,N_17550,N_17139);
nor U18051 (N_18051,N_16548,N_17713);
and U18052 (N_18052,N_17021,N_17599);
nand U18053 (N_18053,N_17687,N_17430);
xnor U18054 (N_18054,N_17244,N_17023);
nor U18055 (N_18055,N_17594,N_17513);
or U18056 (N_18056,N_17233,N_17362);
xnor U18057 (N_18057,N_17477,N_16566);
and U18058 (N_18058,N_17678,N_17670);
or U18059 (N_18059,N_17677,N_17854);
xor U18060 (N_18060,N_17952,N_17866);
and U18061 (N_18061,N_17075,N_16982);
nor U18062 (N_18062,N_17785,N_16532);
and U18063 (N_18063,N_16660,N_16778);
and U18064 (N_18064,N_17958,N_17029);
or U18065 (N_18065,N_16650,N_16716);
or U18066 (N_18066,N_17315,N_16729);
or U18067 (N_18067,N_17210,N_17725);
xnor U18068 (N_18068,N_17201,N_17235);
xnor U18069 (N_18069,N_17338,N_16707);
nor U18070 (N_18070,N_17337,N_17531);
and U18071 (N_18071,N_17535,N_17869);
nor U18072 (N_18072,N_17126,N_16528);
or U18073 (N_18073,N_16508,N_17192);
and U18074 (N_18074,N_17019,N_17011);
nor U18075 (N_18075,N_17765,N_17614);
and U18076 (N_18076,N_16573,N_17135);
and U18077 (N_18077,N_17278,N_16933);
nor U18078 (N_18078,N_17122,N_17121);
nor U18079 (N_18079,N_16558,N_16702);
and U18080 (N_18080,N_17087,N_17200);
xnor U18081 (N_18081,N_17310,N_16989);
and U18082 (N_18082,N_16733,N_17746);
xor U18083 (N_18083,N_17705,N_17003);
nor U18084 (N_18084,N_17153,N_16671);
nor U18085 (N_18085,N_17988,N_17845);
and U18086 (N_18086,N_17470,N_16980);
or U18087 (N_18087,N_17015,N_17459);
xnor U18088 (N_18088,N_17095,N_17600);
nand U18089 (N_18089,N_16743,N_16724);
nor U18090 (N_18090,N_16758,N_17354);
and U18091 (N_18091,N_17818,N_16851);
nor U18092 (N_18092,N_16720,N_16593);
and U18093 (N_18093,N_16891,N_16744);
or U18094 (N_18094,N_16969,N_16553);
nand U18095 (N_18095,N_17168,N_17814);
and U18096 (N_18096,N_17647,N_17069);
xnor U18097 (N_18097,N_17419,N_17867);
nor U18098 (N_18098,N_16538,N_17581);
nor U18099 (N_18099,N_16986,N_16509);
or U18100 (N_18100,N_17117,N_17643);
or U18101 (N_18101,N_17788,N_17538);
xor U18102 (N_18102,N_16617,N_17875);
nand U18103 (N_18103,N_17455,N_17721);
or U18104 (N_18104,N_17717,N_16813);
nor U18105 (N_18105,N_16975,N_17180);
xnor U18106 (N_18106,N_17667,N_17883);
nor U18107 (N_18107,N_17410,N_17100);
and U18108 (N_18108,N_17161,N_17253);
and U18109 (N_18109,N_17114,N_17435);
xnor U18110 (N_18110,N_17987,N_17157);
nor U18111 (N_18111,N_17227,N_17248);
and U18112 (N_18112,N_16978,N_17944);
nand U18113 (N_18113,N_17979,N_17294);
xnor U18114 (N_18114,N_17049,N_17732);
or U18115 (N_18115,N_17859,N_17286);
or U18116 (N_18116,N_17758,N_16821);
or U18117 (N_18117,N_17541,N_16935);
nor U18118 (N_18118,N_16754,N_17324);
and U18119 (N_18119,N_16565,N_17912);
xor U18120 (N_18120,N_16859,N_16854);
nand U18121 (N_18121,N_17730,N_17413);
nand U18122 (N_18122,N_17570,N_17909);
and U18123 (N_18123,N_17656,N_16529);
or U18124 (N_18124,N_17849,N_16793);
xnor U18125 (N_18125,N_17177,N_16789);
nor U18126 (N_18126,N_17360,N_17368);
or U18127 (N_18127,N_17272,N_17482);
or U18128 (N_18128,N_16574,N_16567);
xor U18129 (N_18129,N_17199,N_17065);
nand U18130 (N_18130,N_16857,N_17468);
xor U18131 (N_18131,N_17813,N_17018);
nor U18132 (N_18132,N_17504,N_17137);
and U18133 (N_18133,N_17031,N_17777);
and U18134 (N_18134,N_17565,N_17042);
xnor U18135 (N_18135,N_17150,N_17152);
and U18136 (N_18136,N_17924,N_17532);
and U18137 (N_18137,N_17142,N_16928);
xor U18138 (N_18138,N_17851,N_17499);
or U18139 (N_18139,N_17288,N_17107);
nor U18140 (N_18140,N_16637,N_17819);
xor U18141 (N_18141,N_17415,N_17968);
nand U18142 (N_18142,N_16505,N_16570);
nand U18143 (N_18143,N_16753,N_16837);
nand U18144 (N_18144,N_17835,N_17622);
or U18145 (N_18145,N_17495,N_17269);
xor U18146 (N_18146,N_16632,N_17283);
xnor U18147 (N_18147,N_17690,N_17146);
xor U18148 (N_18148,N_17865,N_17632);
and U18149 (N_18149,N_17915,N_17775);
xor U18150 (N_18150,N_16742,N_16706);
or U18151 (N_18151,N_17542,N_17399);
and U18152 (N_18152,N_17159,N_17009);
nand U18153 (N_18153,N_16901,N_16945);
and U18154 (N_18154,N_17557,N_17301);
or U18155 (N_18155,N_16893,N_16705);
xor U18156 (N_18156,N_17054,N_17704);
nor U18157 (N_18157,N_17084,N_17970);
nor U18158 (N_18158,N_17229,N_17772);
nand U18159 (N_18159,N_16873,N_16820);
nand U18160 (N_18160,N_17809,N_17497);
nor U18161 (N_18161,N_17722,N_17676);
and U18162 (N_18162,N_16985,N_16839);
nand U18163 (N_18163,N_16501,N_17262);
nand U18164 (N_18164,N_16780,N_17365);
nor U18165 (N_18165,N_16988,N_16846);
nand U18166 (N_18166,N_17234,N_16701);
nor U18167 (N_18167,N_17940,N_16895);
xnor U18168 (N_18168,N_17181,N_16542);
xnor U18169 (N_18169,N_17252,N_17428);
nor U18170 (N_18170,N_17088,N_17708);
or U18171 (N_18171,N_17744,N_17645);
nor U18172 (N_18172,N_17680,N_16588);
xnor U18173 (N_18173,N_17997,N_16539);
nor U18174 (N_18174,N_17321,N_17190);
and U18175 (N_18175,N_17887,N_17382);
nor U18176 (N_18176,N_17032,N_17464);
nor U18177 (N_18177,N_16664,N_16878);
and U18178 (N_18178,N_17188,N_17742);
and U18179 (N_18179,N_17584,N_17747);
xor U18180 (N_18180,N_17033,N_16904);
and U18181 (N_18181,N_17378,N_16722);
and U18182 (N_18182,N_17879,N_16540);
nand U18183 (N_18183,N_17836,N_16619);
or U18184 (N_18184,N_17026,N_17085);
xor U18185 (N_18185,N_17441,N_17595);
xnor U18186 (N_18186,N_17969,N_17892);
xor U18187 (N_18187,N_17649,N_17285);
nand U18188 (N_18188,N_17268,N_16673);
and U18189 (N_18189,N_17582,N_17832);
nor U18190 (N_18190,N_17764,N_16812);
nor U18191 (N_18191,N_16731,N_16970);
or U18192 (N_18192,N_17433,N_17757);
xnor U18193 (N_18193,N_17446,N_16992);
and U18194 (N_18194,N_16861,N_16534);
or U18195 (N_18195,N_17536,N_17573);
xor U18196 (N_18196,N_17238,N_17342);
or U18197 (N_18197,N_17502,N_16687);
xor U18198 (N_18198,N_17058,N_16718);
xor U18199 (N_18199,N_16858,N_17218);
nor U18200 (N_18200,N_16603,N_16960);
nand U18201 (N_18201,N_16657,N_16515);
and U18202 (N_18202,N_17906,N_17039);
nor U18203 (N_18203,N_16734,N_16535);
or U18204 (N_18204,N_16947,N_17568);
xnor U18205 (N_18205,N_17804,N_17379);
nor U18206 (N_18206,N_17245,N_17184);
xnor U18207 (N_18207,N_17440,N_17938);
or U18208 (N_18208,N_16677,N_17861);
nand U18209 (N_18209,N_16596,N_17366);
and U18210 (N_18210,N_16900,N_16816);
and U18211 (N_18211,N_16546,N_17005);
nand U18212 (N_18212,N_16836,N_17127);
xnor U18213 (N_18213,N_17800,N_17799);
and U18214 (N_18214,N_17696,N_16759);
or U18215 (N_18215,N_17025,N_16949);
nor U18216 (N_18216,N_16678,N_17490);
nor U18217 (N_18217,N_16685,N_17897);
xor U18218 (N_18218,N_17350,N_17916);
xnor U18219 (N_18219,N_16956,N_17606);
or U18220 (N_18220,N_17871,N_16880);
and U18221 (N_18221,N_17453,N_16633);
nor U18222 (N_18222,N_17682,N_17700);
nand U18223 (N_18223,N_17839,N_16962);
or U18224 (N_18224,N_16958,N_16620);
nand U18225 (N_18225,N_17899,N_17050);
nand U18226 (N_18226,N_17279,N_17450);
nand U18227 (N_18227,N_17345,N_17489);
or U18228 (N_18228,N_17351,N_17304);
and U18229 (N_18229,N_17903,N_17109);
nor U18230 (N_18230,N_17780,N_17609);
and U18231 (N_18231,N_16679,N_16690);
nand U18232 (N_18232,N_17567,N_16994);
or U18233 (N_18233,N_17635,N_17044);
xor U18234 (N_18234,N_17067,N_17098);
nor U18235 (N_18235,N_17518,N_17588);
and U18236 (N_18236,N_16543,N_16751);
or U18237 (N_18237,N_16915,N_17931);
nor U18238 (N_18238,N_17858,N_16898);
nor U18239 (N_18239,N_17840,N_16955);
or U18240 (N_18240,N_17982,N_17000);
nor U18241 (N_18241,N_17904,N_17344);
nor U18242 (N_18242,N_17683,N_17741);
nand U18243 (N_18243,N_17295,N_17715);
nor U18244 (N_18244,N_17271,N_17474);
and U18245 (N_18245,N_16797,N_17193);
xnor U18246 (N_18246,N_17723,N_17424);
nor U18247 (N_18247,N_17309,N_16764);
nor U18248 (N_18248,N_17779,N_17418);
and U18249 (N_18249,N_17605,N_17138);
xnor U18250 (N_18250,N_16921,N_17080);
and U18251 (N_18251,N_17259,N_17112);
nand U18252 (N_18252,N_17144,N_16923);
and U18253 (N_18253,N_17506,N_17731);
and U18254 (N_18254,N_17828,N_17287);
nor U18255 (N_18255,N_17738,N_16834);
xor U18256 (N_18256,N_16569,N_16772);
nand U18257 (N_18257,N_17737,N_17028);
nand U18258 (N_18258,N_17562,N_17620);
nor U18259 (N_18259,N_17421,N_16644);
and U18260 (N_18260,N_17985,N_17675);
nor U18261 (N_18261,N_17590,N_17954);
and U18262 (N_18262,N_16516,N_17894);
nand U18263 (N_18263,N_17079,N_17078);
or U18264 (N_18264,N_17370,N_16831);
nor U18265 (N_18265,N_17243,N_17946);
nor U18266 (N_18266,N_17320,N_17327);
and U18267 (N_18267,N_17561,N_16531);
and U18268 (N_18268,N_16625,N_16571);
xor U18269 (N_18269,N_17060,N_16957);
and U18270 (N_18270,N_16779,N_17325);
and U18271 (N_18271,N_17575,N_16506);
nor U18272 (N_18272,N_17061,N_16922);
nand U18273 (N_18273,N_17801,N_16630);
and U18274 (N_18274,N_16612,N_17577);
and U18275 (N_18275,N_17727,N_16563);
and U18276 (N_18276,N_17108,N_16905);
nor U18277 (N_18277,N_17333,N_16510);
nor U18278 (N_18278,N_17367,N_17558);
nand U18279 (N_18279,N_17444,N_17148);
nand U18280 (N_18280,N_17795,N_16885);
xor U18281 (N_18281,N_17579,N_16715);
or U18282 (N_18282,N_17630,N_17202);
nand U18283 (N_18283,N_16902,N_17305);
xor U18284 (N_18284,N_17487,N_16776);
xor U18285 (N_18285,N_17791,N_17443);
or U18286 (N_18286,N_16940,N_16568);
nor U18287 (N_18287,N_16502,N_17330);
and U18288 (N_18288,N_17983,N_17260);
or U18289 (N_18289,N_17874,N_17921);
nand U18290 (N_18290,N_17179,N_16965);
nand U18291 (N_18291,N_17256,N_17047);
nand U18292 (N_18292,N_16886,N_17569);
xor U18293 (N_18293,N_17759,N_17053);
or U18294 (N_18294,N_17823,N_16887);
and U18295 (N_18295,N_17090,N_17356);
or U18296 (N_18296,N_17638,N_17774);
nand U18297 (N_18297,N_16786,N_17523);
nand U18298 (N_18298,N_17401,N_16547);
nor U18299 (N_18299,N_16848,N_17101);
and U18300 (N_18300,N_17007,N_17756);
or U18301 (N_18301,N_17884,N_17170);
nand U18302 (N_18302,N_16911,N_16913);
and U18303 (N_18303,N_16642,N_17480);
nand U18304 (N_18304,N_16907,N_17514);
or U18305 (N_18305,N_17965,N_17830);
nand U18306 (N_18306,N_16586,N_17412);
or U18307 (N_18307,N_17010,N_17918);
or U18308 (N_18308,N_17461,N_17300);
nor U18309 (N_18309,N_17237,N_17826);
nor U18310 (N_18310,N_16598,N_16578);
or U18311 (N_18311,N_17664,N_17314);
xnor U18312 (N_18312,N_16576,N_16967);
nand U18313 (N_18313,N_17926,N_17786);
and U18314 (N_18314,N_17002,N_16641);
nor U18315 (N_18315,N_17782,N_17546);
nand U18316 (N_18316,N_17593,N_17598);
and U18317 (N_18317,N_17893,N_17284);
and U18318 (N_18318,N_17824,N_16708);
and U18319 (N_18319,N_17355,N_17068);
nand U18320 (N_18320,N_16806,N_16616);
and U18321 (N_18321,N_17665,N_17257);
or U18322 (N_18322,N_16748,N_17749);
xnor U18323 (N_18323,N_17613,N_16977);
nor U18324 (N_18324,N_17890,N_16815);
or U18325 (N_18325,N_17844,N_17947);
or U18326 (N_18326,N_17317,N_16870);
nor U18327 (N_18327,N_16608,N_16920);
nor U18328 (N_18328,N_16561,N_16910);
xnor U18329 (N_18329,N_17640,N_16691);
and U18330 (N_18330,N_16631,N_16807);
nor U18331 (N_18331,N_16931,N_17174);
xor U18332 (N_18332,N_17977,N_17163);
or U18333 (N_18333,N_17674,N_16953);
nor U18334 (N_18334,N_17547,N_17156);
and U18335 (N_18335,N_17386,N_17703);
and U18336 (N_18336,N_16613,N_17205);
xor U18337 (N_18337,N_16794,N_17197);
nand U18338 (N_18338,N_16583,N_17335);
or U18339 (N_18339,N_17962,N_17071);
or U18340 (N_18340,N_16939,N_17755);
nand U18341 (N_18341,N_17392,N_17426);
and U18342 (N_18342,N_17629,N_17974);
nor U18343 (N_18343,N_17034,N_17996);
and U18344 (N_18344,N_17374,N_16645);
or U18345 (N_18345,N_16897,N_17463);
nand U18346 (N_18346,N_16952,N_16799);
and U18347 (N_18347,N_16626,N_17914);
nor U18348 (N_18348,N_17213,N_17967);
xnor U18349 (N_18349,N_17339,N_17394);
and U18350 (N_18350,N_17376,N_17847);
or U18351 (N_18351,N_17817,N_17763);
or U18352 (N_18352,N_17022,N_16627);
or U18353 (N_18353,N_16654,N_16700);
nor U18354 (N_18354,N_17024,N_17057);
xnor U18355 (N_18355,N_16926,N_17383);
xnor U18356 (N_18356,N_17306,N_17978);
nand U18357 (N_18357,N_16943,N_17950);
and U18358 (N_18358,N_17064,N_17494);
nor U18359 (N_18359,N_16903,N_17539);
nand U18360 (N_18360,N_17270,N_16863);
nand U18361 (N_18361,N_17743,N_16647);
and U18362 (N_18362,N_17885,N_16849);
and U18363 (N_18363,N_16643,N_17693);
xor U18364 (N_18364,N_17132,N_16711);
and U18365 (N_18365,N_17939,N_17694);
or U18366 (N_18366,N_17391,N_16600);
or U18367 (N_18367,N_16545,N_17343);
nand U18368 (N_18368,N_17739,N_17106);
or U18369 (N_18369,N_17241,N_17820);
nand U18370 (N_18370,N_17580,N_16788);
and U18371 (N_18371,N_16996,N_16971);
nand U18372 (N_18372,N_17120,N_16818);
nand U18373 (N_18373,N_16549,N_17527);
and U18374 (N_18374,N_17214,N_17224);
nand U18375 (N_18375,N_17349,N_17886);
xnor U18376 (N_18376,N_17510,N_16514);
nor U18377 (N_18377,N_16888,N_17056);
xnor U18378 (N_18378,N_17642,N_17429);
nand U18379 (N_18379,N_17512,N_16765);
nand U18380 (N_18380,N_16979,N_17230);
nor U18381 (N_18381,N_16973,N_16683);
and U18382 (N_18382,N_17329,N_17027);
and U18383 (N_18383,N_17559,N_17864);
or U18384 (N_18384,N_17290,N_17431);
and U18385 (N_18385,N_17853,N_17151);
nor U18386 (N_18386,N_16692,N_16746);
xnor U18387 (N_18387,N_17930,N_17388);
xnor U18388 (N_18388,N_16530,N_17655);
or U18389 (N_18389,N_16963,N_16597);
or U18390 (N_18390,N_16595,N_17628);
nand U18391 (N_18391,N_17937,N_17631);
nand U18392 (N_18392,N_16503,N_17020);
nand U18393 (N_18393,N_16784,N_16875);
or U18394 (N_18394,N_17895,N_17129);
or U18395 (N_18395,N_17902,N_17189);
xor U18396 (N_18396,N_17863,N_17277);
and U18397 (N_18397,N_16823,N_17439);
or U18398 (N_18398,N_16688,N_17891);
nand U18399 (N_18399,N_16850,N_16752);
nor U18400 (N_18400,N_17718,N_17971);
nand U18401 (N_18401,N_17724,N_17533);
and U18402 (N_18402,N_16518,N_17528);
and U18403 (N_18403,N_17017,N_17695);
nor U18404 (N_18404,N_17934,N_17852);
nor U18405 (N_18405,N_17292,N_17610);
and U18406 (N_18406,N_17882,N_17409);
and U18407 (N_18407,N_16695,N_16762);
nand U18408 (N_18408,N_16916,N_16826);
nand U18409 (N_18409,N_17267,N_17781);
nand U18410 (N_18410,N_16811,N_16845);
or U18411 (N_18411,N_16699,N_17991);
or U18412 (N_18412,N_16801,N_17877);
and U18413 (N_18413,N_17077,N_17748);
nor U18414 (N_18414,N_16712,N_16517);
nand U18415 (N_18415,N_17929,N_17908);
and U18416 (N_18416,N_16852,N_17707);
nor U18417 (N_18417,N_16822,N_16577);
and U18418 (N_18418,N_17543,N_16721);
or U18419 (N_18419,N_17933,N_16966);
or U18420 (N_18420,N_17264,N_17445);
nor U18421 (N_18421,N_16594,N_16838);
nand U18422 (N_18422,N_16787,N_17932);
and U18423 (N_18423,N_17046,N_16500);
xnor U18424 (N_18424,N_16855,N_16937);
nor U18425 (N_18425,N_17697,N_16810);
xnor U18426 (N_18426,N_17611,N_16656);
nor U18427 (N_18427,N_16552,N_17927);
and U18428 (N_18428,N_17709,N_17663);
nand U18429 (N_18429,N_17167,N_17016);
xnor U18430 (N_18430,N_17407,N_17955);
nor U18431 (N_18431,N_16841,N_16761);
or U18432 (N_18432,N_17298,N_17837);
and U18433 (N_18433,N_16615,N_17767);
or U18434 (N_18434,N_17639,N_16640);
nand U18435 (N_18435,N_16842,N_17462);
and U18436 (N_18436,N_17282,N_17432);
and U18437 (N_18437,N_16714,N_16868);
or U18438 (N_18438,N_17936,N_17784);
and U18439 (N_18439,N_16580,N_17797);
nor U18440 (N_18440,N_17816,N_17500);
or U18441 (N_18441,N_16649,N_17975);
and U18442 (N_18442,N_17448,N_17364);
nand U18443 (N_18443,N_17460,N_17951);
xnor U18444 (N_18444,N_17242,N_16782);
or U18445 (N_18445,N_17805,N_16676);
or U18446 (N_18446,N_17681,N_16581);
or U18447 (N_18447,N_17634,N_16882);
nand U18448 (N_18448,N_16843,N_17993);
xnor U18449 (N_18449,N_17396,N_17627);
nand U18450 (N_18450,N_16525,N_17615);
xor U18451 (N_18451,N_16974,N_16766);
nor U18452 (N_18452,N_17263,N_16934);
nor U18453 (N_18453,N_17030,N_17651);
nor U18454 (N_18454,N_17302,N_17650);
xor U18455 (N_18455,N_16541,N_16638);
xor U18456 (N_18456,N_17953,N_16659);
and U18457 (N_18457,N_17092,N_16662);
xnor U18458 (N_18458,N_17052,N_16520);
xor U18459 (N_18459,N_17081,N_17398);
and U18460 (N_18460,N_17423,N_17941);
and U18461 (N_18461,N_16653,N_16521);
or U18462 (N_18462,N_17469,N_17232);
or U18463 (N_18463,N_17815,N_17076);
nor U18464 (N_18464,N_17070,N_17994);
or U18465 (N_18465,N_17652,N_17761);
xnor U18466 (N_18466,N_16769,N_17160);
xor U18467 (N_18467,N_16800,N_17481);
and U18468 (N_18468,N_17551,N_17155);
or U18469 (N_18469,N_16930,N_17740);
nand U18470 (N_18470,N_17359,N_17679);
nor U18471 (N_18471,N_17373,N_17072);
nor U18472 (N_18472,N_17515,N_17789);
or U18473 (N_18473,N_17013,N_17555);
xnor U18474 (N_18474,N_16555,N_17608);
and U18475 (N_18475,N_17778,N_17729);
nor U18476 (N_18476,N_17458,N_17750);
nor U18477 (N_18477,N_17714,N_17091);
nor U18478 (N_18478,N_16628,N_16767);
xor U18479 (N_18479,N_17841,N_17073);
and U18480 (N_18480,N_17659,N_16672);
nor U18481 (N_18481,N_17066,N_17623);
xnor U18482 (N_18482,N_17124,N_16757);
nand U18483 (N_18483,N_16665,N_16550);
nand U18484 (N_18484,N_17178,N_16728);
or U18485 (N_18485,N_17654,N_17411);
nand U18486 (N_18486,N_16735,N_17089);
and U18487 (N_18487,N_16591,N_17191);
nor U18488 (N_18488,N_16526,N_16924);
and U18489 (N_18489,N_16829,N_16918);
and U18490 (N_18490,N_16959,N_17525);
nor U18491 (N_18491,N_17254,N_16732);
nand U18492 (N_18492,N_17530,N_16512);
and U18493 (N_18493,N_17503,N_17491);
or U18494 (N_18494,N_16796,N_17662);
nand U18495 (N_18495,N_17603,N_16981);
and U18496 (N_18496,N_17827,N_17299);
nor U18497 (N_18497,N_17597,N_16755);
or U18498 (N_18498,N_17483,N_17303);
or U18499 (N_18499,N_17094,N_17736);
and U18500 (N_18500,N_17668,N_17769);
xnor U18501 (N_18501,N_17706,N_16670);
xor U18502 (N_18502,N_16572,N_16646);
xnor U18503 (N_18503,N_16869,N_17571);
nand U18504 (N_18504,N_16750,N_17719);
and U18505 (N_18505,N_17900,N_16781);
or U18506 (N_18506,N_17416,N_17692);
and U18507 (N_18507,N_17296,N_17641);
xnor U18508 (N_18508,N_17710,N_16775);
xor U18509 (N_18509,N_17176,N_17318);
nand U18510 (N_18510,N_16871,N_17658);
or U18511 (N_18511,N_17164,N_17855);
nand U18512 (N_18512,N_17751,N_17529);
or U18513 (N_18513,N_16738,N_17626);
xnor U18514 (N_18514,N_16533,N_17843);
nand U18515 (N_18515,N_17592,N_16777);
nand U18516 (N_18516,N_17116,N_16609);
nand U18517 (N_18517,N_16999,N_16639);
nand U18518 (N_18518,N_16704,N_17905);
or U18519 (N_18519,N_17083,N_17226);
nand U18520 (N_18520,N_17964,N_17880);
nor U18521 (N_18521,N_17957,N_17361);
or U18522 (N_18522,N_17848,N_17012);
xnor U18523 (N_18523,N_16946,N_16693);
nand U18524 (N_18524,N_16511,N_16606);
xnor U18525 (N_18525,N_17265,N_17646);
xnor U18526 (N_18526,N_16749,N_17768);
nor U18527 (N_18527,N_17434,N_16876);
nor U18528 (N_18528,N_17702,N_17842);
or U18529 (N_18529,N_17297,N_17385);
nor U18530 (N_18530,N_17616,N_17806);
and U18531 (N_18531,N_17347,N_17896);
and U18532 (N_18532,N_17564,N_17086);
xor U18533 (N_18533,N_17872,N_17006);
nor U18534 (N_18534,N_17976,N_16584);
or U18535 (N_18535,N_16889,N_17943);
and U18536 (N_18536,N_17621,N_17901);
nand U18537 (N_18537,N_17633,N_17522);
nand U18538 (N_18538,N_17607,N_17456);
nand U18539 (N_18539,N_16537,N_16623);
nor U18540 (N_18540,N_16987,N_16948);
nor U18541 (N_18541,N_17959,N_16527);
or U18542 (N_18542,N_17688,N_17850);
nand U18543 (N_18543,N_16804,N_16675);
or U18544 (N_18544,N_17473,N_17147);
and U18545 (N_18545,N_17215,N_17661);
nand U18546 (N_18546,N_16835,N_17175);
nand U18547 (N_18547,N_17545,N_16710);
nor U18548 (N_18548,N_17485,N_16856);
xor U18549 (N_18549,N_16652,N_17111);
and U18550 (N_18550,N_17313,N_16909);
or U18551 (N_18551,N_17043,N_17403);
xnor U18552 (N_18552,N_17984,N_16703);
and U18553 (N_18553,N_17348,N_17776);
nand U18554 (N_18554,N_17141,N_16551);
xnor U18555 (N_18555,N_17136,N_17406);
and U18556 (N_18556,N_17517,N_16944);
and U18557 (N_18557,N_16814,N_16562);
xnor U18558 (N_18558,N_17666,N_17720);
xor U18559 (N_18559,N_17618,N_17149);
nor U18560 (N_18560,N_17115,N_17182);
nand U18561 (N_18561,N_17082,N_17534);
and U18562 (N_18562,N_17158,N_17436);
or U18563 (N_18563,N_17113,N_17041);
xnor U18564 (N_18564,N_17563,N_17986);
and U18565 (N_18565,N_17123,N_16864);
nand U18566 (N_18566,N_17960,N_17363);
xor U18567 (N_18567,N_17173,N_17183);
xor U18568 (N_18568,N_17258,N_17334);
or U18569 (N_18569,N_17357,N_17508);
nor U18570 (N_18570,N_17326,N_16932);
and U18571 (N_18571,N_17249,N_16817);
or U18572 (N_18572,N_17236,N_17711);
xor U18573 (N_18573,N_17217,N_17478);
or U18574 (N_18574,N_16592,N_17625);
and U18575 (N_18575,N_16651,N_16942);
or U18576 (N_18576,N_17870,N_17998);
xnor U18577 (N_18577,N_17689,N_17228);
and U18578 (N_18578,N_17308,N_16783);
nand U18579 (N_18579,N_16618,N_16634);
and U18580 (N_18580,N_17657,N_17372);
nor U18581 (N_18581,N_17587,N_17917);
or U18582 (N_18582,N_16785,N_16602);
or U18583 (N_18583,N_16976,N_17898);
nand U18584 (N_18584,N_17311,N_17001);
nor U18585 (N_18585,N_16833,N_17221);
xor U18586 (N_18586,N_16927,N_16559);
or U18587 (N_18587,N_17810,N_17920);
or U18588 (N_18588,N_16773,N_17194);
nand U18589 (N_18589,N_17185,N_17556);
nor U18590 (N_18590,N_16661,N_16727);
nor U18591 (N_18591,N_17222,N_17822);
or U18592 (N_18592,N_17624,N_17038);
xor U18593 (N_18593,N_17204,N_17422);
or U18594 (N_18594,N_17648,N_16587);
or U18595 (N_18595,N_16899,N_17636);
or U18596 (N_18596,N_17289,N_16840);
xor U18597 (N_18597,N_16938,N_17673);
nor U18598 (N_18598,N_16635,N_17701);
or U18599 (N_18599,N_17726,N_17671);
xnor U18600 (N_18600,N_17619,N_17035);
and U18601 (N_18601,N_16853,N_17857);
xnor U18602 (N_18602,N_17812,N_17427);
nand U18603 (N_18603,N_16929,N_16791);
or U18604 (N_18604,N_17753,N_17125);
and U18605 (N_18605,N_17913,N_16740);
nor U18606 (N_18606,N_17246,N_17454);
nor U18607 (N_18607,N_17479,N_17208);
nor U18608 (N_18608,N_17437,N_17923);
nand U18609 (N_18609,N_17856,N_16624);
or U18610 (N_18610,N_17511,N_16582);
nand U18611 (N_18611,N_17381,N_17465);
xor U18612 (N_18612,N_17496,N_16998);
nor U18613 (N_18613,N_17811,N_17273);
nand U18614 (N_18614,N_17216,N_16771);
nor U18615 (N_18615,N_17762,N_17405);
or U18616 (N_18616,N_17400,N_17910);
xor U18617 (N_18617,N_17519,N_16655);
nand U18618 (N_18618,N_17389,N_16792);
nor U18619 (N_18619,N_17544,N_17860);
or U18620 (N_18620,N_17583,N_17752);
nand U18621 (N_18621,N_17206,N_17862);
or U18622 (N_18622,N_17808,N_17990);
or U18623 (N_18623,N_17239,N_17888);
nand U18624 (N_18624,N_17322,N_17644);
nand U18625 (N_18625,N_16824,N_16832);
nand U18626 (N_18626,N_16954,N_16557);
and U18627 (N_18627,N_16725,N_16798);
nand U18628 (N_18628,N_17585,N_17062);
and U18629 (N_18629,N_16827,N_17251);
nand U18630 (N_18630,N_16737,N_17733);
and U18631 (N_18631,N_17104,N_17420);
and U18632 (N_18632,N_17307,N_17766);
nand U18633 (N_18633,N_16601,N_17505);
nor U18634 (N_18634,N_17074,N_16713);
and U18635 (N_18635,N_16681,N_17591);
nor U18636 (N_18636,N_16604,N_17404);
nand U18637 (N_18637,N_17291,N_17669);
and U18638 (N_18638,N_16760,N_17375);
and U18639 (N_18639,N_16717,N_17807);
or U18640 (N_18640,N_17219,N_17754);
xnor U18641 (N_18641,N_17956,N_16684);
nor U18642 (N_18642,N_17735,N_17240);
and U18643 (N_18643,N_17604,N_17250);
and U18644 (N_18644,N_17873,N_17745);
or U18645 (N_18645,N_17728,N_16830);
or U18646 (N_18646,N_17973,N_17942);
and U18647 (N_18647,N_16860,N_17516);
xor U18648 (N_18648,N_16556,N_17783);
nand U18649 (N_18649,N_17760,N_17451);
nand U18650 (N_18650,N_17716,N_16865);
or U18651 (N_18651,N_16805,N_17103);
nand U18652 (N_18652,N_17699,N_17792);
or U18653 (N_18653,N_16666,N_16648);
and U18654 (N_18654,N_17878,N_17377);
or U18655 (N_18655,N_16698,N_16726);
nor U18656 (N_18656,N_16809,N_17803);
and U18657 (N_18657,N_17560,N_17475);
nor U18658 (N_18658,N_17549,N_17387);
or U18659 (N_18659,N_17110,N_16519);
xnor U18660 (N_18660,N_16872,N_16993);
nand U18661 (N_18661,N_17328,N_17055);
xor U18662 (N_18662,N_16605,N_17274);
xor U18663 (N_18663,N_16723,N_17128);
nand U18664 (N_18664,N_17578,N_17332);
and U18665 (N_18665,N_17169,N_17948);
nor U18666 (N_18666,N_17384,N_17966);
nand U18667 (N_18667,N_16741,N_17196);
or U18668 (N_18668,N_17846,N_17051);
xnor U18669 (N_18669,N_16739,N_16694);
xnor U18670 (N_18670,N_17276,N_17488);
nand U18671 (N_18671,N_16983,N_17576);
and U18672 (N_18672,N_16790,N_16560);
nand U18673 (N_18673,N_17524,N_17552);
nand U18674 (N_18674,N_17371,N_17172);
xnor U18675 (N_18675,N_17911,N_16745);
and U18676 (N_18676,N_17008,N_17838);
nor U18677 (N_18677,N_17414,N_16686);
xor U18678 (N_18678,N_16866,N_16629);
xor U18679 (N_18679,N_17417,N_17198);
or U18680 (N_18680,N_17145,N_16879);
nor U18681 (N_18681,N_17889,N_16919);
or U18682 (N_18682,N_17589,N_17247);
nor U18683 (N_18683,N_16680,N_17586);
xnor U18684 (N_18684,N_16883,N_16847);
and U18685 (N_18685,N_16674,N_17316);
or U18686 (N_18686,N_16756,N_17438);
or U18687 (N_18687,N_17685,N_16844);
nor U18688 (N_18688,N_16513,N_17919);
xnor U18689 (N_18689,N_17612,N_17045);
nor U18690 (N_18690,N_17063,N_17134);
and U18691 (N_18691,N_17566,N_16991);
and U18692 (N_18692,N_17734,N_17698);
nor U18693 (N_18693,N_17493,N_17961);
or U18694 (N_18694,N_16621,N_17980);
nor U18695 (N_18695,N_17130,N_16747);
nand U18696 (N_18696,N_17452,N_17457);
or U18697 (N_18697,N_16877,N_16668);
xor U18698 (N_18698,N_17340,N_16802);
nand U18699 (N_18699,N_16917,N_16984);
or U18700 (N_18700,N_17358,N_16522);
nor U18701 (N_18701,N_16507,N_17105);
and U18702 (N_18702,N_17554,N_16950);
nor U18703 (N_18703,N_17449,N_17617);
and U18704 (N_18704,N_17833,N_17119);
xor U18705 (N_18705,N_16874,N_17672);
xor U18706 (N_18706,N_17876,N_17187);
xnor U18707 (N_18707,N_17526,N_16709);
nor U18708 (N_18708,N_17989,N_17140);
and U18709 (N_18709,N_16585,N_17097);
or U18710 (N_18710,N_17133,N_17154);
nor U18711 (N_18711,N_17834,N_16912);
nand U18712 (N_18712,N_16689,N_17999);
and U18713 (N_18713,N_17793,N_17686);
and U18714 (N_18714,N_17691,N_16599);
xor U18715 (N_18715,N_16669,N_17281);
nand U18716 (N_18716,N_17831,N_17211);
and U18717 (N_18717,N_16896,N_17802);
and U18718 (N_18718,N_17319,N_17992);
or U18719 (N_18719,N_17165,N_17498);
and U18720 (N_18720,N_17203,N_17928);
xor U18721 (N_18721,N_16808,N_16951);
nor U18722 (N_18722,N_17501,N_17467);
nor U18723 (N_18723,N_16894,N_16504);
or U18724 (N_18724,N_16697,N_17787);
nor U18725 (N_18725,N_17476,N_17771);
or U18726 (N_18726,N_17393,N_16575);
and U18727 (N_18727,N_17059,N_17223);
or U18728 (N_18728,N_17166,N_17186);
nor U18729 (N_18729,N_16667,N_16972);
nand U18730 (N_18730,N_17395,N_17935);
and U18731 (N_18731,N_17225,N_16964);
nand U18732 (N_18732,N_17521,N_17472);
or U18733 (N_18733,N_17486,N_17868);
nand U18734 (N_18734,N_16795,N_16610);
and U18735 (N_18735,N_17972,N_16936);
nand U18736 (N_18736,N_16997,N_17821);
nor U18737 (N_18737,N_16825,N_17341);
nor U18738 (N_18738,N_17040,N_16990);
xor U18739 (N_18739,N_16881,N_17131);
or U18740 (N_18740,N_17925,N_16523);
nand U18741 (N_18741,N_17346,N_16614);
xor U18742 (N_18742,N_17093,N_17212);
nand U18743 (N_18743,N_17537,N_17442);
xnor U18744 (N_18744,N_16730,N_17798);
or U18745 (N_18745,N_17540,N_17660);
nand U18746 (N_18746,N_17331,N_16696);
or U18747 (N_18747,N_17981,N_16908);
xnor U18748 (N_18748,N_17509,N_17323);
or U18749 (N_18749,N_17293,N_17601);
and U18750 (N_18750,N_17375,N_16660);
nand U18751 (N_18751,N_16758,N_17010);
nand U18752 (N_18752,N_17272,N_16817);
nand U18753 (N_18753,N_16984,N_17832);
or U18754 (N_18754,N_17414,N_16871);
nand U18755 (N_18755,N_17097,N_17783);
nand U18756 (N_18756,N_17062,N_17887);
nand U18757 (N_18757,N_17524,N_17359);
xor U18758 (N_18758,N_17396,N_16777);
nor U18759 (N_18759,N_17731,N_17272);
and U18760 (N_18760,N_16668,N_16569);
and U18761 (N_18761,N_17501,N_17240);
or U18762 (N_18762,N_17618,N_16639);
nand U18763 (N_18763,N_17928,N_16919);
nand U18764 (N_18764,N_16526,N_16939);
nor U18765 (N_18765,N_16662,N_17657);
or U18766 (N_18766,N_17927,N_17686);
nor U18767 (N_18767,N_16559,N_16666);
and U18768 (N_18768,N_17933,N_17791);
and U18769 (N_18769,N_17147,N_16655);
nor U18770 (N_18770,N_17328,N_17837);
or U18771 (N_18771,N_16702,N_16565);
nand U18772 (N_18772,N_17091,N_17711);
and U18773 (N_18773,N_16553,N_17622);
and U18774 (N_18774,N_17518,N_17278);
and U18775 (N_18775,N_16865,N_17875);
nand U18776 (N_18776,N_16554,N_17901);
nor U18777 (N_18777,N_16556,N_17094);
nand U18778 (N_18778,N_16713,N_16964);
nand U18779 (N_18779,N_17105,N_16749);
and U18780 (N_18780,N_17383,N_17317);
or U18781 (N_18781,N_17771,N_16948);
nor U18782 (N_18782,N_16767,N_17952);
nand U18783 (N_18783,N_16596,N_17678);
xor U18784 (N_18784,N_16577,N_17332);
nand U18785 (N_18785,N_17838,N_16532);
nor U18786 (N_18786,N_16789,N_17004);
xor U18787 (N_18787,N_17985,N_17624);
nand U18788 (N_18788,N_17475,N_16686);
and U18789 (N_18789,N_17424,N_17029);
and U18790 (N_18790,N_17308,N_16631);
xnor U18791 (N_18791,N_17599,N_16542);
xnor U18792 (N_18792,N_17373,N_17036);
nand U18793 (N_18793,N_17915,N_17669);
nor U18794 (N_18794,N_17234,N_17682);
xor U18795 (N_18795,N_17760,N_16816);
nor U18796 (N_18796,N_17557,N_16912);
or U18797 (N_18797,N_16549,N_16682);
nor U18798 (N_18798,N_16781,N_17418);
and U18799 (N_18799,N_16805,N_17797);
nand U18800 (N_18800,N_17607,N_17202);
and U18801 (N_18801,N_17767,N_16794);
or U18802 (N_18802,N_17886,N_16501);
nand U18803 (N_18803,N_16549,N_17528);
and U18804 (N_18804,N_17656,N_17800);
nand U18805 (N_18805,N_16662,N_17142);
nand U18806 (N_18806,N_16734,N_17221);
nand U18807 (N_18807,N_16802,N_17849);
nor U18808 (N_18808,N_17735,N_16822);
xnor U18809 (N_18809,N_17854,N_17654);
xnor U18810 (N_18810,N_17777,N_17299);
xnor U18811 (N_18811,N_17924,N_17734);
nor U18812 (N_18812,N_17562,N_17225);
xor U18813 (N_18813,N_17160,N_17495);
or U18814 (N_18814,N_17732,N_17529);
or U18815 (N_18815,N_17399,N_16672);
nor U18816 (N_18816,N_16933,N_16738);
nor U18817 (N_18817,N_17930,N_17936);
or U18818 (N_18818,N_17606,N_17660);
and U18819 (N_18819,N_17965,N_17861);
nor U18820 (N_18820,N_17467,N_16564);
xnor U18821 (N_18821,N_17273,N_17024);
and U18822 (N_18822,N_17992,N_17805);
or U18823 (N_18823,N_17326,N_17944);
xor U18824 (N_18824,N_16948,N_17349);
xnor U18825 (N_18825,N_17393,N_17795);
nand U18826 (N_18826,N_16735,N_16619);
or U18827 (N_18827,N_16938,N_17127);
or U18828 (N_18828,N_17722,N_17232);
and U18829 (N_18829,N_16993,N_17282);
xnor U18830 (N_18830,N_17738,N_16792);
nand U18831 (N_18831,N_16950,N_17937);
and U18832 (N_18832,N_17245,N_17147);
or U18833 (N_18833,N_17593,N_16909);
nand U18834 (N_18834,N_16769,N_16832);
nand U18835 (N_18835,N_16712,N_17199);
xnor U18836 (N_18836,N_16777,N_17092);
xnor U18837 (N_18837,N_17679,N_17999);
or U18838 (N_18838,N_17718,N_16973);
xnor U18839 (N_18839,N_17541,N_17489);
and U18840 (N_18840,N_17931,N_16573);
xnor U18841 (N_18841,N_16887,N_17643);
nand U18842 (N_18842,N_17449,N_16876);
or U18843 (N_18843,N_17334,N_17830);
nor U18844 (N_18844,N_17925,N_16585);
or U18845 (N_18845,N_17976,N_17575);
or U18846 (N_18846,N_17940,N_17102);
nand U18847 (N_18847,N_17771,N_16709);
or U18848 (N_18848,N_17108,N_17686);
nor U18849 (N_18849,N_17294,N_16852);
xnor U18850 (N_18850,N_17447,N_16769);
nor U18851 (N_18851,N_16820,N_17360);
or U18852 (N_18852,N_17465,N_16841);
nand U18853 (N_18853,N_16631,N_17601);
nand U18854 (N_18854,N_17779,N_17099);
nand U18855 (N_18855,N_17031,N_16959);
nand U18856 (N_18856,N_17230,N_17552);
nor U18857 (N_18857,N_17065,N_16882);
xor U18858 (N_18858,N_17647,N_17725);
or U18859 (N_18859,N_17523,N_17794);
nand U18860 (N_18860,N_17870,N_17957);
and U18861 (N_18861,N_17338,N_16726);
nor U18862 (N_18862,N_17114,N_16959);
or U18863 (N_18863,N_17444,N_16783);
nor U18864 (N_18864,N_17747,N_17526);
nand U18865 (N_18865,N_17573,N_17022);
or U18866 (N_18866,N_17606,N_16833);
or U18867 (N_18867,N_16570,N_17039);
and U18868 (N_18868,N_17131,N_16638);
xnor U18869 (N_18869,N_16587,N_17881);
nor U18870 (N_18870,N_17021,N_17886);
or U18871 (N_18871,N_16716,N_16800);
and U18872 (N_18872,N_17674,N_16732);
nand U18873 (N_18873,N_16646,N_17658);
nand U18874 (N_18874,N_17079,N_17736);
or U18875 (N_18875,N_17850,N_17671);
or U18876 (N_18876,N_17023,N_17242);
nor U18877 (N_18877,N_16854,N_17332);
nand U18878 (N_18878,N_16993,N_16641);
and U18879 (N_18879,N_17920,N_17345);
nor U18880 (N_18880,N_17383,N_17217);
nor U18881 (N_18881,N_17790,N_16877);
nand U18882 (N_18882,N_16903,N_17777);
or U18883 (N_18883,N_16965,N_16993);
and U18884 (N_18884,N_17214,N_17396);
and U18885 (N_18885,N_17284,N_17364);
xnor U18886 (N_18886,N_16546,N_16776);
nand U18887 (N_18887,N_17118,N_17330);
nand U18888 (N_18888,N_17436,N_17616);
and U18889 (N_18889,N_16927,N_17215);
or U18890 (N_18890,N_17532,N_17613);
and U18891 (N_18891,N_17966,N_17844);
nor U18892 (N_18892,N_17775,N_17810);
nand U18893 (N_18893,N_17479,N_17688);
xnor U18894 (N_18894,N_16655,N_16677);
or U18895 (N_18895,N_17212,N_17545);
xor U18896 (N_18896,N_17322,N_17093);
and U18897 (N_18897,N_17892,N_16815);
nand U18898 (N_18898,N_17556,N_16581);
nor U18899 (N_18899,N_16674,N_16915);
and U18900 (N_18900,N_16784,N_16714);
nor U18901 (N_18901,N_17962,N_17637);
nor U18902 (N_18902,N_17953,N_17325);
or U18903 (N_18903,N_17953,N_17068);
nor U18904 (N_18904,N_16763,N_17728);
xnor U18905 (N_18905,N_16506,N_16951);
nor U18906 (N_18906,N_17986,N_16749);
nor U18907 (N_18907,N_17480,N_16906);
and U18908 (N_18908,N_17371,N_17017);
nand U18909 (N_18909,N_17103,N_17611);
xnor U18910 (N_18910,N_16722,N_17757);
xnor U18911 (N_18911,N_17588,N_17708);
nor U18912 (N_18912,N_17016,N_17666);
and U18913 (N_18913,N_17132,N_17918);
nor U18914 (N_18914,N_17395,N_17984);
and U18915 (N_18915,N_17265,N_17266);
and U18916 (N_18916,N_17387,N_17800);
nand U18917 (N_18917,N_16980,N_16736);
nand U18918 (N_18918,N_17083,N_16549);
or U18919 (N_18919,N_16687,N_17864);
nand U18920 (N_18920,N_17837,N_17712);
and U18921 (N_18921,N_17472,N_17646);
nand U18922 (N_18922,N_17453,N_17629);
and U18923 (N_18923,N_16697,N_17421);
xor U18924 (N_18924,N_17877,N_16594);
or U18925 (N_18925,N_16696,N_16516);
nor U18926 (N_18926,N_17376,N_17921);
nand U18927 (N_18927,N_17594,N_16503);
xnor U18928 (N_18928,N_17117,N_17554);
or U18929 (N_18929,N_16592,N_17924);
xnor U18930 (N_18930,N_17133,N_16634);
or U18931 (N_18931,N_17669,N_16806);
and U18932 (N_18932,N_17516,N_16874);
and U18933 (N_18933,N_16999,N_16908);
nand U18934 (N_18934,N_17555,N_17215);
or U18935 (N_18935,N_17686,N_17305);
nor U18936 (N_18936,N_16519,N_17760);
and U18937 (N_18937,N_17454,N_17184);
and U18938 (N_18938,N_17739,N_17031);
and U18939 (N_18939,N_17914,N_17995);
xor U18940 (N_18940,N_17307,N_17160);
and U18941 (N_18941,N_17409,N_16777);
xnor U18942 (N_18942,N_16748,N_16938);
xnor U18943 (N_18943,N_17211,N_17016);
xor U18944 (N_18944,N_17072,N_17238);
or U18945 (N_18945,N_17096,N_17482);
nor U18946 (N_18946,N_17004,N_16883);
and U18947 (N_18947,N_17090,N_17399);
xnor U18948 (N_18948,N_16994,N_17095);
nand U18949 (N_18949,N_17069,N_17491);
or U18950 (N_18950,N_16623,N_16602);
nor U18951 (N_18951,N_16510,N_16875);
xor U18952 (N_18952,N_17728,N_17424);
nand U18953 (N_18953,N_16912,N_16836);
nand U18954 (N_18954,N_16754,N_16929);
xor U18955 (N_18955,N_17742,N_17289);
nand U18956 (N_18956,N_17733,N_17806);
nor U18957 (N_18957,N_17551,N_17523);
xor U18958 (N_18958,N_17133,N_16648);
and U18959 (N_18959,N_17826,N_17944);
nor U18960 (N_18960,N_17981,N_17820);
xnor U18961 (N_18961,N_17003,N_16698);
nand U18962 (N_18962,N_17599,N_17667);
nand U18963 (N_18963,N_17511,N_16520);
and U18964 (N_18964,N_16947,N_16798);
nor U18965 (N_18965,N_17600,N_17821);
or U18966 (N_18966,N_17146,N_16987);
and U18967 (N_18967,N_17316,N_17791);
xnor U18968 (N_18968,N_17588,N_17392);
xnor U18969 (N_18969,N_16606,N_17797);
xor U18970 (N_18970,N_17312,N_17762);
nand U18971 (N_18971,N_17760,N_16622);
or U18972 (N_18972,N_17851,N_17681);
nor U18973 (N_18973,N_16996,N_17876);
nor U18974 (N_18974,N_17355,N_16722);
or U18975 (N_18975,N_17220,N_16608);
and U18976 (N_18976,N_17162,N_16541);
xor U18977 (N_18977,N_16657,N_17210);
nor U18978 (N_18978,N_17146,N_16984);
nor U18979 (N_18979,N_17732,N_17145);
xnor U18980 (N_18980,N_17025,N_17274);
nand U18981 (N_18981,N_17585,N_17355);
and U18982 (N_18982,N_17153,N_16575);
or U18983 (N_18983,N_17851,N_17280);
and U18984 (N_18984,N_17584,N_17752);
nand U18985 (N_18985,N_16712,N_17357);
nor U18986 (N_18986,N_17817,N_17656);
and U18987 (N_18987,N_16923,N_16768);
or U18988 (N_18988,N_17649,N_16527);
and U18989 (N_18989,N_17705,N_17323);
or U18990 (N_18990,N_17155,N_16854);
xor U18991 (N_18991,N_17289,N_17951);
nand U18992 (N_18992,N_17143,N_16581);
or U18993 (N_18993,N_16612,N_16967);
nand U18994 (N_18994,N_17302,N_16927);
xor U18995 (N_18995,N_17283,N_16756);
xnor U18996 (N_18996,N_17979,N_17714);
xnor U18997 (N_18997,N_17233,N_17654);
nor U18998 (N_18998,N_17345,N_17218);
xnor U18999 (N_18999,N_16785,N_16754);
or U19000 (N_19000,N_16905,N_17178);
and U19001 (N_19001,N_17469,N_17987);
nand U19002 (N_19002,N_17693,N_17033);
nor U19003 (N_19003,N_17208,N_16538);
xnor U19004 (N_19004,N_17236,N_17952);
or U19005 (N_19005,N_17106,N_17192);
nand U19006 (N_19006,N_16904,N_17368);
and U19007 (N_19007,N_17753,N_17967);
nand U19008 (N_19008,N_17527,N_17317);
xnor U19009 (N_19009,N_17557,N_16761);
nand U19010 (N_19010,N_17680,N_16559);
nand U19011 (N_19011,N_17384,N_17297);
nand U19012 (N_19012,N_16937,N_17993);
or U19013 (N_19013,N_17797,N_17546);
nand U19014 (N_19014,N_17283,N_17269);
nor U19015 (N_19015,N_17786,N_17315);
nand U19016 (N_19016,N_17533,N_17212);
nand U19017 (N_19017,N_16908,N_17949);
nand U19018 (N_19018,N_17360,N_16705);
nand U19019 (N_19019,N_17025,N_17368);
xnor U19020 (N_19020,N_17666,N_17964);
xor U19021 (N_19021,N_16501,N_17795);
or U19022 (N_19022,N_17496,N_17211);
and U19023 (N_19023,N_16818,N_16926);
and U19024 (N_19024,N_17564,N_16765);
and U19025 (N_19025,N_16981,N_16533);
or U19026 (N_19026,N_17809,N_17302);
or U19027 (N_19027,N_16841,N_17709);
xnor U19028 (N_19028,N_17573,N_16501);
xnor U19029 (N_19029,N_17168,N_16599);
xor U19030 (N_19030,N_16658,N_17341);
nor U19031 (N_19031,N_17271,N_17804);
or U19032 (N_19032,N_17646,N_17244);
nor U19033 (N_19033,N_16667,N_17085);
nor U19034 (N_19034,N_17418,N_16897);
or U19035 (N_19035,N_17592,N_16767);
nand U19036 (N_19036,N_16991,N_17661);
and U19037 (N_19037,N_17772,N_17266);
nor U19038 (N_19038,N_16836,N_17915);
nor U19039 (N_19039,N_16876,N_16598);
nand U19040 (N_19040,N_17219,N_17321);
nand U19041 (N_19041,N_17072,N_16834);
or U19042 (N_19042,N_17897,N_17069);
and U19043 (N_19043,N_17367,N_17109);
nand U19044 (N_19044,N_17299,N_17617);
nor U19045 (N_19045,N_16859,N_17776);
nand U19046 (N_19046,N_16672,N_17357);
xnor U19047 (N_19047,N_16796,N_16713);
nand U19048 (N_19048,N_17130,N_16619);
xor U19049 (N_19049,N_17531,N_17046);
or U19050 (N_19050,N_16765,N_17046);
nand U19051 (N_19051,N_16800,N_17206);
nand U19052 (N_19052,N_17550,N_16986);
xnor U19053 (N_19053,N_17074,N_17506);
and U19054 (N_19054,N_16961,N_17181);
or U19055 (N_19055,N_17756,N_17647);
xor U19056 (N_19056,N_17522,N_16855);
and U19057 (N_19057,N_17371,N_16508);
or U19058 (N_19058,N_16762,N_17228);
nor U19059 (N_19059,N_16760,N_16742);
and U19060 (N_19060,N_17124,N_17742);
nor U19061 (N_19061,N_16593,N_17130);
and U19062 (N_19062,N_16742,N_16692);
nand U19063 (N_19063,N_17014,N_17288);
or U19064 (N_19064,N_16866,N_17377);
and U19065 (N_19065,N_17078,N_17623);
nor U19066 (N_19066,N_16839,N_17775);
nand U19067 (N_19067,N_16954,N_16957);
nor U19068 (N_19068,N_16614,N_16775);
xor U19069 (N_19069,N_16664,N_16917);
nor U19070 (N_19070,N_17644,N_16815);
nand U19071 (N_19071,N_17601,N_16932);
xor U19072 (N_19072,N_17654,N_17565);
and U19073 (N_19073,N_17678,N_17901);
nand U19074 (N_19074,N_17184,N_17448);
xnor U19075 (N_19075,N_17638,N_16754);
nor U19076 (N_19076,N_17719,N_16875);
nor U19077 (N_19077,N_16614,N_17730);
and U19078 (N_19078,N_16991,N_16912);
nor U19079 (N_19079,N_16769,N_16633);
nand U19080 (N_19080,N_17897,N_16544);
or U19081 (N_19081,N_17749,N_16751);
or U19082 (N_19082,N_17470,N_17398);
or U19083 (N_19083,N_17002,N_17837);
or U19084 (N_19084,N_16571,N_17274);
xnor U19085 (N_19085,N_16811,N_16624);
or U19086 (N_19086,N_16963,N_17702);
or U19087 (N_19087,N_16652,N_17014);
xor U19088 (N_19088,N_17346,N_16627);
xnor U19089 (N_19089,N_17335,N_17909);
or U19090 (N_19090,N_16917,N_17427);
nand U19091 (N_19091,N_16862,N_17415);
or U19092 (N_19092,N_16681,N_17500);
nand U19093 (N_19093,N_16601,N_16637);
or U19094 (N_19094,N_17979,N_17734);
xnor U19095 (N_19095,N_17448,N_16759);
or U19096 (N_19096,N_16699,N_17226);
nand U19097 (N_19097,N_16502,N_16571);
xor U19098 (N_19098,N_17016,N_17896);
xnor U19099 (N_19099,N_17407,N_16574);
nand U19100 (N_19100,N_17476,N_17366);
xnor U19101 (N_19101,N_17054,N_17213);
nand U19102 (N_19102,N_17706,N_17200);
xor U19103 (N_19103,N_17562,N_17548);
or U19104 (N_19104,N_17662,N_16715);
and U19105 (N_19105,N_17153,N_16530);
and U19106 (N_19106,N_16903,N_16692);
and U19107 (N_19107,N_17175,N_16773);
and U19108 (N_19108,N_16520,N_17485);
xnor U19109 (N_19109,N_17650,N_17894);
nor U19110 (N_19110,N_17335,N_17360);
nor U19111 (N_19111,N_17953,N_17268);
or U19112 (N_19112,N_17334,N_16945);
nand U19113 (N_19113,N_16719,N_16673);
nand U19114 (N_19114,N_16523,N_17734);
and U19115 (N_19115,N_17700,N_17764);
or U19116 (N_19116,N_17793,N_17796);
and U19117 (N_19117,N_16765,N_16518);
nor U19118 (N_19118,N_17660,N_17238);
nor U19119 (N_19119,N_17015,N_16742);
nand U19120 (N_19120,N_16518,N_17565);
nor U19121 (N_19121,N_17016,N_17097);
xor U19122 (N_19122,N_17007,N_17284);
and U19123 (N_19123,N_17309,N_17751);
xor U19124 (N_19124,N_16526,N_16538);
nand U19125 (N_19125,N_17373,N_17661);
nand U19126 (N_19126,N_16628,N_17303);
nor U19127 (N_19127,N_17444,N_16673);
or U19128 (N_19128,N_16648,N_16862);
nor U19129 (N_19129,N_17580,N_17178);
xnor U19130 (N_19130,N_16592,N_17784);
nand U19131 (N_19131,N_16583,N_16577);
or U19132 (N_19132,N_17054,N_16712);
or U19133 (N_19133,N_16571,N_17064);
nand U19134 (N_19134,N_16740,N_16638);
or U19135 (N_19135,N_17349,N_17831);
nand U19136 (N_19136,N_16863,N_17402);
and U19137 (N_19137,N_17330,N_17974);
and U19138 (N_19138,N_16655,N_16943);
nand U19139 (N_19139,N_16787,N_17545);
and U19140 (N_19140,N_16808,N_17824);
nand U19141 (N_19141,N_17187,N_16810);
nand U19142 (N_19142,N_17832,N_16716);
nand U19143 (N_19143,N_17224,N_17051);
nor U19144 (N_19144,N_17147,N_16539);
nand U19145 (N_19145,N_17453,N_17152);
nor U19146 (N_19146,N_16630,N_16502);
and U19147 (N_19147,N_17148,N_17709);
or U19148 (N_19148,N_17186,N_17405);
nand U19149 (N_19149,N_16512,N_16880);
nand U19150 (N_19150,N_17266,N_17286);
and U19151 (N_19151,N_16679,N_17602);
nor U19152 (N_19152,N_16872,N_17466);
xnor U19153 (N_19153,N_16673,N_16979);
xor U19154 (N_19154,N_17251,N_17510);
xnor U19155 (N_19155,N_17645,N_16963);
and U19156 (N_19156,N_17522,N_17638);
nor U19157 (N_19157,N_16751,N_17573);
or U19158 (N_19158,N_16800,N_17064);
and U19159 (N_19159,N_17866,N_17968);
nor U19160 (N_19160,N_17006,N_16717);
nand U19161 (N_19161,N_17416,N_17516);
xnor U19162 (N_19162,N_17357,N_17106);
nand U19163 (N_19163,N_17972,N_16501);
xnor U19164 (N_19164,N_17744,N_17093);
nor U19165 (N_19165,N_17511,N_17425);
nand U19166 (N_19166,N_17550,N_17542);
nand U19167 (N_19167,N_16701,N_16766);
xnor U19168 (N_19168,N_16857,N_17303);
nand U19169 (N_19169,N_17722,N_16782);
and U19170 (N_19170,N_17363,N_16799);
nand U19171 (N_19171,N_17024,N_17010);
and U19172 (N_19172,N_17631,N_17186);
nor U19173 (N_19173,N_17626,N_16779);
nor U19174 (N_19174,N_16537,N_16939);
and U19175 (N_19175,N_17426,N_17273);
xor U19176 (N_19176,N_16562,N_17488);
and U19177 (N_19177,N_17573,N_16665);
nand U19178 (N_19178,N_17840,N_17977);
and U19179 (N_19179,N_17994,N_16741);
or U19180 (N_19180,N_17859,N_17066);
and U19181 (N_19181,N_16664,N_16723);
and U19182 (N_19182,N_17089,N_16868);
and U19183 (N_19183,N_17960,N_17492);
and U19184 (N_19184,N_17916,N_17954);
nand U19185 (N_19185,N_17118,N_17570);
nor U19186 (N_19186,N_16740,N_17220);
and U19187 (N_19187,N_17405,N_17151);
nor U19188 (N_19188,N_17104,N_17946);
nor U19189 (N_19189,N_17984,N_16612);
or U19190 (N_19190,N_16595,N_17926);
nand U19191 (N_19191,N_16516,N_17541);
xor U19192 (N_19192,N_17968,N_17362);
nand U19193 (N_19193,N_17311,N_17421);
xor U19194 (N_19194,N_16646,N_17578);
and U19195 (N_19195,N_16596,N_16535);
xor U19196 (N_19196,N_16882,N_17894);
xor U19197 (N_19197,N_17733,N_17359);
xor U19198 (N_19198,N_16820,N_16668);
nand U19199 (N_19199,N_17653,N_17013);
xor U19200 (N_19200,N_17521,N_17176);
or U19201 (N_19201,N_17171,N_16882);
nor U19202 (N_19202,N_16678,N_17725);
or U19203 (N_19203,N_17550,N_17574);
and U19204 (N_19204,N_16753,N_17882);
or U19205 (N_19205,N_17626,N_16902);
or U19206 (N_19206,N_17725,N_17095);
nand U19207 (N_19207,N_17454,N_17572);
and U19208 (N_19208,N_16962,N_17249);
or U19209 (N_19209,N_17521,N_17778);
xnor U19210 (N_19210,N_17483,N_17289);
nand U19211 (N_19211,N_16675,N_17406);
and U19212 (N_19212,N_17711,N_17996);
or U19213 (N_19213,N_17618,N_17723);
or U19214 (N_19214,N_17011,N_16800);
or U19215 (N_19215,N_17271,N_17288);
or U19216 (N_19216,N_16605,N_16933);
xnor U19217 (N_19217,N_17220,N_17466);
or U19218 (N_19218,N_17283,N_17900);
and U19219 (N_19219,N_17617,N_17665);
and U19220 (N_19220,N_17287,N_16979);
nand U19221 (N_19221,N_16954,N_17244);
and U19222 (N_19222,N_17621,N_17458);
nor U19223 (N_19223,N_16582,N_17739);
xor U19224 (N_19224,N_17186,N_16832);
nand U19225 (N_19225,N_17602,N_16823);
nor U19226 (N_19226,N_17277,N_17508);
xor U19227 (N_19227,N_17705,N_16794);
or U19228 (N_19228,N_17024,N_16893);
or U19229 (N_19229,N_17794,N_17080);
nand U19230 (N_19230,N_16618,N_17588);
or U19231 (N_19231,N_16904,N_16694);
xor U19232 (N_19232,N_16934,N_16796);
nor U19233 (N_19233,N_17569,N_16538);
and U19234 (N_19234,N_17669,N_17665);
xnor U19235 (N_19235,N_16563,N_16999);
xor U19236 (N_19236,N_17996,N_17337);
nand U19237 (N_19237,N_17923,N_16915);
and U19238 (N_19238,N_16716,N_17635);
xnor U19239 (N_19239,N_17697,N_17141);
nor U19240 (N_19240,N_17396,N_17165);
nor U19241 (N_19241,N_17414,N_17784);
and U19242 (N_19242,N_16747,N_17623);
or U19243 (N_19243,N_16826,N_17001);
xnor U19244 (N_19244,N_17838,N_16930);
and U19245 (N_19245,N_17995,N_17270);
and U19246 (N_19246,N_17002,N_17621);
nor U19247 (N_19247,N_17830,N_17885);
nand U19248 (N_19248,N_17378,N_17178);
nand U19249 (N_19249,N_17479,N_16875);
xnor U19250 (N_19250,N_17188,N_17722);
nand U19251 (N_19251,N_16993,N_17057);
and U19252 (N_19252,N_17207,N_17423);
nand U19253 (N_19253,N_16924,N_17388);
nand U19254 (N_19254,N_17545,N_17054);
and U19255 (N_19255,N_17240,N_17478);
nor U19256 (N_19256,N_16654,N_17784);
nand U19257 (N_19257,N_17845,N_17044);
nand U19258 (N_19258,N_17865,N_17020);
nor U19259 (N_19259,N_16872,N_17269);
nand U19260 (N_19260,N_17263,N_16800);
or U19261 (N_19261,N_16624,N_17381);
nor U19262 (N_19262,N_16793,N_16933);
nor U19263 (N_19263,N_17599,N_16707);
xor U19264 (N_19264,N_17142,N_17259);
nor U19265 (N_19265,N_17889,N_17879);
nand U19266 (N_19266,N_17116,N_17442);
nand U19267 (N_19267,N_16921,N_16860);
and U19268 (N_19268,N_17330,N_17476);
or U19269 (N_19269,N_17437,N_17064);
xnor U19270 (N_19270,N_17518,N_16780);
or U19271 (N_19271,N_17895,N_17861);
or U19272 (N_19272,N_17455,N_17242);
or U19273 (N_19273,N_17033,N_17177);
nor U19274 (N_19274,N_17648,N_17429);
or U19275 (N_19275,N_17069,N_16589);
or U19276 (N_19276,N_17619,N_17363);
xnor U19277 (N_19277,N_17775,N_16710);
or U19278 (N_19278,N_17914,N_16511);
nand U19279 (N_19279,N_17754,N_17361);
and U19280 (N_19280,N_17518,N_16607);
xor U19281 (N_19281,N_17188,N_17155);
nor U19282 (N_19282,N_17991,N_17738);
or U19283 (N_19283,N_16936,N_17836);
or U19284 (N_19284,N_16563,N_16617);
and U19285 (N_19285,N_17025,N_16589);
nor U19286 (N_19286,N_17758,N_17408);
nor U19287 (N_19287,N_16799,N_16629);
nor U19288 (N_19288,N_17493,N_16509);
and U19289 (N_19289,N_17449,N_17980);
nor U19290 (N_19290,N_17847,N_17339);
and U19291 (N_19291,N_17402,N_17822);
and U19292 (N_19292,N_17902,N_17906);
and U19293 (N_19293,N_17042,N_17081);
xor U19294 (N_19294,N_17211,N_17981);
nor U19295 (N_19295,N_17519,N_17201);
nand U19296 (N_19296,N_17538,N_16816);
nor U19297 (N_19297,N_17421,N_16972);
or U19298 (N_19298,N_17501,N_17440);
or U19299 (N_19299,N_17024,N_17238);
and U19300 (N_19300,N_17625,N_16673);
and U19301 (N_19301,N_16916,N_16603);
or U19302 (N_19302,N_16793,N_16547);
and U19303 (N_19303,N_17694,N_17605);
xor U19304 (N_19304,N_16698,N_17949);
and U19305 (N_19305,N_16905,N_17367);
xnor U19306 (N_19306,N_16627,N_17370);
or U19307 (N_19307,N_17798,N_17181);
xnor U19308 (N_19308,N_16845,N_17722);
xor U19309 (N_19309,N_16649,N_16981);
or U19310 (N_19310,N_16566,N_17863);
nand U19311 (N_19311,N_16722,N_16844);
and U19312 (N_19312,N_16970,N_17126);
nor U19313 (N_19313,N_17842,N_16870);
or U19314 (N_19314,N_17751,N_17083);
and U19315 (N_19315,N_17605,N_17362);
or U19316 (N_19316,N_17312,N_16851);
xor U19317 (N_19317,N_17425,N_17240);
xnor U19318 (N_19318,N_17084,N_17327);
nor U19319 (N_19319,N_17836,N_17388);
xor U19320 (N_19320,N_17236,N_17341);
xnor U19321 (N_19321,N_17996,N_17459);
and U19322 (N_19322,N_16626,N_17042);
nand U19323 (N_19323,N_17692,N_16526);
and U19324 (N_19324,N_17705,N_17801);
xnor U19325 (N_19325,N_16902,N_17224);
nor U19326 (N_19326,N_17745,N_17645);
xnor U19327 (N_19327,N_17774,N_17738);
or U19328 (N_19328,N_17375,N_17458);
xnor U19329 (N_19329,N_17551,N_17166);
nand U19330 (N_19330,N_17413,N_16981);
and U19331 (N_19331,N_17126,N_17594);
or U19332 (N_19332,N_17985,N_16587);
xnor U19333 (N_19333,N_17133,N_16598);
nor U19334 (N_19334,N_17172,N_17167);
or U19335 (N_19335,N_16514,N_17346);
and U19336 (N_19336,N_17156,N_17539);
or U19337 (N_19337,N_17631,N_17654);
and U19338 (N_19338,N_17123,N_16942);
nand U19339 (N_19339,N_16649,N_17112);
xnor U19340 (N_19340,N_17179,N_17092);
xor U19341 (N_19341,N_17395,N_17943);
and U19342 (N_19342,N_17216,N_17134);
nand U19343 (N_19343,N_17513,N_17567);
xnor U19344 (N_19344,N_17867,N_16762);
nor U19345 (N_19345,N_17221,N_17471);
and U19346 (N_19346,N_17178,N_16941);
or U19347 (N_19347,N_17110,N_17231);
or U19348 (N_19348,N_16847,N_16932);
and U19349 (N_19349,N_17215,N_17839);
xor U19350 (N_19350,N_17372,N_17660);
nor U19351 (N_19351,N_17426,N_17009);
or U19352 (N_19352,N_17576,N_17078);
nand U19353 (N_19353,N_17819,N_17766);
and U19354 (N_19354,N_17058,N_17623);
and U19355 (N_19355,N_17055,N_17439);
nor U19356 (N_19356,N_17968,N_17496);
or U19357 (N_19357,N_17533,N_17391);
xnor U19358 (N_19358,N_17118,N_17104);
nor U19359 (N_19359,N_17459,N_17946);
nand U19360 (N_19360,N_16969,N_17935);
nor U19361 (N_19361,N_16649,N_17696);
and U19362 (N_19362,N_16908,N_17770);
xnor U19363 (N_19363,N_17550,N_17215);
nand U19364 (N_19364,N_17041,N_17849);
nand U19365 (N_19365,N_16660,N_17793);
and U19366 (N_19366,N_16926,N_16517);
or U19367 (N_19367,N_16780,N_16935);
nor U19368 (N_19368,N_17553,N_17865);
or U19369 (N_19369,N_16894,N_16599);
and U19370 (N_19370,N_17909,N_17674);
and U19371 (N_19371,N_17947,N_17720);
or U19372 (N_19372,N_17928,N_17934);
and U19373 (N_19373,N_17791,N_17307);
xor U19374 (N_19374,N_16758,N_16646);
nor U19375 (N_19375,N_16618,N_17894);
or U19376 (N_19376,N_17452,N_17729);
xnor U19377 (N_19377,N_17246,N_17561);
nand U19378 (N_19378,N_17691,N_17323);
nor U19379 (N_19379,N_16712,N_16602);
nand U19380 (N_19380,N_17006,N_17501);
nand U19381 (N_19381,N_16965,N_16547);
xor U19382 (N_19382,N_16977,N_16858);
nand U19383 (N_19383,N_17047,N_17595);
nor U19384 (N_19384,N_17387,N_17467);
and U19385 (N_19385,N_17944,N_17620);
or U19386 (N_19386,N_16928,N_16780);
nor U19387 (N_19387,N_17790,N_17401);
and U19388 (N_19388,N_17777,N_17587);
xnor U19389 (N_19389,N_17134,N_17517);
nor U19390 (N_19390,N_17305,N_16957);
nor U19391 (N_19391,N_17686,N_17723);
nand U19392 (N_19392,N_17423,N_17755);
nor U19393 (N_19393,N_16967,N_16541);
nor U19394 (N_19394,N_16537,N_17034);
xor U19395 (N_19395,N_17145,N_17993);
nand U19396 (N_19396,N_17146,N_17996);
and U19397 (N_19397,N_17836,N_16637);
xnor U19398 (N_19398,N_17501,N_17267);
nor U19399 (N_19399,N_17552,N_17759);
or U19400 (N_19400,N_17198,N_16506);
nor U19401 (N_19401,N_17806,N_16985);
xnor U19402 (N_19402,N_16772,N_17793);
or U19403 (N_19403,N_17825,N_16911);
and U19404 (N_19404,N_16563,N_16897);
nor U19405 (N_19405,N_17061,N_17995);
nand U19406 (N_19406,N_16863,N_17948);
or U19407 (N_19407,N_17197,N_17252);
nor U19408 (N_19408,N_17762,N_17308);
nor U19409 (N_19409,N_17880,N_17302);
and U19410 (N_19410,N_17396,N_17333);
or U19411 (N_19411,N_16624,N_17262);
and U19412 (N_19412,N_17838,N_16782);
nand U19413 (N_19413,N_17525,N_17357);
nor U19414 (N_19414,N_16990,N_17507);
nor U19415 (N_19415,N_17047,N_16898);
xnor U19416 (N_19416,N_17135,N_17965);
xnor U19417 (N_19417,N_17497,N_16737);
nor U19418 (N_19418,N_17902,N_17325);
or U19419 (N_19419,N_17888,N_17204);
nand U19420 (N_19420,N_16643,N_16888);
or U19421 (N_19421,N_17326,N_17383);
nor U19422 (N_19422,N_17987,N_17370);
or U19423 (N_19423,N_16813,N_17903);
and U19424 (N_19424,N_17381,N_16550);
nor U19425 (N_19425,N_17601,N_17873);
nand U19426 (N_19426,N_17250,N_17566);
nor U19427 (N_19427,N_16938,N_16647);
or U19428 (N_19428,N_17089,N_17571);
nor U19429 (N_19429,N_17257,N_17854);
or U19430 (N_19430,N_16974,N_17925);
or U19431 (N_19431,N_17885,N_17284);
and U19432 (N_19432,N_17329,N_17823);
and U19433 (N_19433,N_16980,N_16988);
xnor U19434 (N_19434,N_16936,N_17541);
nand U19435 (N_19435,N_17254,N_17999);
nand U19436 (N_19436,N_17915,N_17616);
nand U19437 (N_19437,N_16778,N_16727);
nand U19438 (N_19438,N_17508,N_17522);
and U19439 (N_19439,N_17285,N_17358);
and U19440 (N_19440,N_17969,N_17395);
nor U19441 (N_19441,N_17349,N_16539);
xor U19442 (N_19442,N_17317,N_16588);
and U19443 (N_19443,N_16731,N_17144);
or U19444 (N_19444,N_17497,N_16612);
nand U19445 (N_19445,N_17735,N_17886);
xor U19446 (N_19446,N_16642,N_17145);
nor U19447 (N_19447,N_17686,N_16755);
nand U19448 (N_19448,N_17830,N_16974);
nor U19449 (N_19449,N_17861,N_16833);
xnor U19450 (N_19450,N_17654,N_16835);
or U19451 (N_19451,N_17349,N_16993);
nor U19452 (N_19452,N_16958,N_16540);
nand U19453 (N_19453,N_17993,N_17090);
xnor U19454 (N_19454,N_16658,N_17496);
nand U19455 (N_19455,N_17002,N_17883);
or U19456 (N_19456,N_17895,N_17297);
or U19457 (N_19457,N_17095,N_17668);
nand U19458 (N_19458,N_17847,N_17348);
xor U19459 (N_19459,N_16746,N_17096);
xor U19460 (N_19460,N_16971,N_17091);
nor U19461 (N_19461,N_16730,N_17578);
and U19462 (N_19462,N_17127,N_17128);
xnor U19463 (N_19463,N_17804,N_17436);
or U19464 (N_19464,N_17591,N_16816);
nand U19465 (N_19465,N_17139,N_17333);
nor U19466 (N_19466,N_17901,N_17313);
or U19467 (N_19467,N_17365,N_16823);
nor U19468 (N_19468,N_17349,N_17523);
nand U19469 (N_19469,N_17729,N_17039);
or U19470 (N_19470,N_16593,N_16523);
or U19471 (N_19471,N_17066,N_17610);
xor U19472 (N_19472,N_17208,N_17304);
nand U19473 (N_19473,N_17203,N_16684);
and U19474 (N_19474,N_17062,N_17146);
and U19475 (N_19475,N_17766,N_17639);
nand U19476 (N_19476,N_17253,N_17339);
xor U19477 (N_19477,N_17025,N_17914);
nor U19478 (N_19478,N_16965,N_17226);
nand U19479 (N_19479,N_16882,N_17705);
and U19480 (N_19480,N_16532,N_17433);
nor U19481 (N_19481,N_17918,N_16778);
nor U19482 (N_19482,N_16580,N_16958);
nor U19483 (N_19483,N_16729,N_17624);
xnor U19484 (N_19484,N_16531,N_17512);
nor U19485 (N_19485,N_16535,N_16768);
nor U19486 (N_19486,N_17818,N_16984);
xnor U19487 (N_19487,N_16761,N_17072);
nand U19488 (N_19488,N_17510,N_16864);
xnor U19489 (N_19489,N_16630,N_17275);
nand U19490 (N_19490,N_17827,N_16748);
xnor U19491 (N_19491,N_17232,N_16844);
nand U19492 (N_19492,N_17526,N_17406);
nor U19493 (N_19493,N_16725,N_17496);
and U19494 (N_19494,N_17568,N_16598);
xnor U19495 (N_19495,N_17448,N_17028);
nor U19496 (N_19496,N_16573,N_17454);
and U19497 (N_19497,N_17361,N_17760);
xnor U19498 (N_19498,N_17409,N_17742);
nor U19499 (N_19499,N_17494,N_16993);
nor U19500 (N_19500,N_18669,N_18055);
or U19501 (N_19501,N_18438,N_18005);
nor U19502 (N_19502,N_19406,N_19364);
nand U19503 (N_19503,N_19113,N_18768);
nor U19504 (N_19504,N_18785,N_19156);
nand U19505 (N_19505,N_19437,N_19476);
nor U19506 (N_19506,N_18367,N_18011);
or U19507 (N_19507,N_18806,N_18665);
xor U19508 (N_19508,N_18819,N_18988);
nand U19509 (N_19509,N_19439,N_18387);
and U19510 (N_19510,N_19092,N_18719);
and U19511 (N_19511,N_18182,N_19365);
and U19512 (N_19512,N_18181,N_18897);
and U19513 (N_19513,N_18158,N_18923);
nand U19514 (N_19514,N_18696,N_18906);
nor U19515 (N_19515,N_18036,N_18341);
or U19516 (N_19516,N_18389,N_18363);
xor U19517 (N_19517,N_18787,N_18645);
nand U19518 (N_19518,N_19350,N_18807);
nand U19519 (N_19519,N_18965,N_18809);
nand U19520 (N_19520,N_18144,N_18022);
or U19521 (N_19521,N_18938,N_18945);
nand U19522 (N_19522,N_18166,N_18304);
and U19523 (N_19523,N_18732,N_18789);
or U19524 (N_19524,N_19182,N_18340);
xor U19525 (N_19525,N_18921,N_18691);
nand U19526 (N_19526,N_19420,N_18744);
xor U19527 (N_19527,N_18268,N_19486);
or U19528 (N_19528,N_18640,N_18274);
and U19529 (N_19529,N_18335,N_18790);
nand U19530 (N_19530,N_18277,N_19009);
and U19531 (N_19531,N_18107,N_18431);
and U19532 (N_19532,N_18541,N_18685);
nand U19533 (N_19533,N_18175,N_18489);
nand U19534 (N_19534,N_18153,N_19396);
nand U19535 (N_19535,N_18936,N_18991);
or U19536 (N_19536,N_18009,N_18003);
nor U19537 (N_19537,N_18602,N_19292);
nor U19538 (N_19538,N_18636,N_18714);
nor U19539 (N_19539,N_18984,N_18034);
nor U19540 (N_19540,N_18128,N_18373);
nor U19541 (N_19541,N_18400,N_18237);
and U19542 (N_19542,N_18279,N_18875);
and U19543 (N_19543,N_18288,N_19033);
or U19544 (N_19544,N_18186,N_18197);
xor U19545 (N_19545,N_19171,N_18347);
and U19546 (N_19546,N_18683,N_19190);
or U19547 (N_19547,N_19006,N_18354);
nand U19548 (N_19548,N_18667,N_18899);
nand U19549 (N_19549,N_19431,N_19013);
and U19550 (N_19550,N_18550,N_19327);
nor U19551 (N_19551,N_18090,N_19127);
xnor U19552 (N_19552,N_18693,N_19151);
or U19553 (N_19553,N_18738,N_18520);
and U19554 (N_19554,N_19496,N_18468);
xnor U19555 (N_19555,N_19294,N_18466);
or U19556 (N_19556,N_18053,N_19371);
and U19557 (N_19557,N_19441,N_18653);
nand U19558 (N_19558,N_18699,N_18599);
xor U19559 (N_19559,N_18631,N_18731);
nor U19560 (N_19560,N_18678,N_19107);
nor U19561 (N_19561,N_18384,N_19287);
nand U19562 (N_19562,N_18303,N_19362);
nand U19563 (N_19563,N_18914,N_18476);
nand U19564 (N_19564,N_18014,N_18568);
nand U19565 (N_19565,N_18278,N_18089);
xnor U19566 (N_19566,N_19453,N_19491);
nand U19567 (N_19567,N_19068,N_18574);
nand U19568 (N_19568,N_18276,N_18345);
nor U19569 (N_19569,N_19048,N_18001);
or U19570 (N_19570,N_18503,N_19197);
or U19571 (N_19571,N_19320,N_19025);
xnor U19572 (N_19572,N_18954,N_18536);
nor U19573 (N_19573,N_18007,N_19326);
and U19574 (N_19574,N_18200,N_18717);
nor U19575 (N_19575,N_19429,N_18123);
and U19576 (N_19576,N_19099,N_19374);
nor U19577 (N_19577,N_18156,N_19458);
xor U19578 (N_19578,N_18904,N_18490);
xor U19579 (N_19579,N_18828,N_19049);
and U19580 (N_19580,N_18085,N_18800);
xnor U19581 (N_19581,N_18511,N_19062);
nand U19582 (N_19582,N_19153,N_18901);
xor U19583 (N_19583,N_18894,N_18791);
and U19584 (N_19584,N_19051,N_19154);
nand U19585 (N_19585,N_18759,N_19200);
nor U19586 (N_19586,N_18600,N_18168);
or U19587 (N_19587,N_18404,N_18213);
and U19588 (N_19588,N_19319,N_19030);
nand U19589 (N_19589,N_19040,N_18573);
xnor U19590 (N_19590,N_18896,N_19100);
or U19591 (N_19591,N_19264,N_19426);
nand U19592 (N_19592,N_18539,N_18078);
nor U19593 (N_19593,N_18134,N_18098);
and U19594 (N_19594,N_18544,N_19240);
nand U19595 (N_19595,N_18730,N_18967);
nand U19596 (N_19596,N_18149,N_19367);
nand U19597 (N_19597,N_18758,N_19119);
nand U19598 (N_19598,N_18285,N_18233);
xor U19599 (N_19599,N_18530,N_19355);
xnor U19600 (N_19600,N_18068,N_18677);
nor U19601 (N_19601,N_19370,N_19072);
and U19602 (N_19602,N_18690,N_18486);
nand U19603 (N_19603,N_18666,N_18358);
xor U19604 (N_19604,N_18747,N_19340);
or U19605 (N_19605,N_18646,N_18911);
and U19606 (N_19606,N_18483,N_19415);
and U19607 (N_19607,N_19216,N_18112);
and U19608 (N_19608,N_18760,N_18119);
and U19609 (N_19609,N_19424,N_18905);
xor U19610 (N_19610,N_18810,N_18224);
nand U19611 (N_19611,N_19202,N_19306);
and U19612 (N_19612,N_19465,N_18617);
nand U19613 (N_19613,N_19477,N_18299);
nor U19614 (N_19614,N_18701,N_18004);
xnor U19615 (N_19615,N_18023,N_19313);
and U19616 (N_19616,N_18604,N_19311);
or U19617 (N_19617,N_18019,N_18969);
nor U19618 (N_19618,N_18915,N_19086);
xnor U19619 (N_19619,N_18368,N_18577);
nor U19620 (N_19620,N_18942,N_18359);
and U19621 (N_19621,N_19198,N_19463);
and U19622 (N_19622,N_18079,N_18879);
nor U19623 (N_19623,N_18727,N_19170);
nand U19624 (N_19624,N_19008,N_19121);
and U19625 (N_19625,N_18515,N_19281);
or U19626 (N_19626,N_19417,N_19318);
or U19627 (N_19627,N_18674,N_18458);
xor U19628 (N_19628,N_19215,N_18523);
or U19629 (N_19629,N_18201,N_18205);
nand U19630 (N_19630,N_18083,N_18661);
or U19631 (N_19631,N_18649,N_18910);
nand U19632 (N_19632,N_19032,N_19308);
or U19633 (N_19633,N_18793,N_18049);
or U19634 (N_19634,N_18664,N_19179);
nand U19635 (N_19635,N_18320,N_18086);
xnor U19636 (N_19636,N_19332,N_19066);
or U19637 (N_19637,N_18099,N_18397);
and U19638 (N_19638,N_18075,N_18115);
nor U19639 (N_19639,N_18337,N_18560);
nand U19640 (N_19640,N_18021,N_18094);
xnor U19641 (N_19641,N_18888,N_19225);
nor U19642 (N_19642,N_18297,N_18704);
or U19643 (N_19643,N_19296,N_18977);
or U19644 (N_19644,N_19079,N_19189);
nand U19645 (N_19645,N_19139,N_19118);
nor U19646 (N_19646,N_18111,N_18870);
and U19647 (N_19647,N_18774,N_18162);
and U19648 (N_19648,N_18949,N_19137);
or U19649 (N_19649,N_18006,N_18582);
nor U19650 (N_19650,N_19065,N_18203);
nor U19651 (N_19651,N_19193,N_19247);
and U19652 (N_19652,N_18627,N_19445);
or U19653 (N_19653,N_18456,N_18709);
nor U19654 (N_19654,N_18041,N_18048);
nand U19655 (N_19655,N_18628,N_19352);
and U19656 (N_19656,N_18644,N_18650);
xor U19657 (N_19657,N_18686,N_18794);
nor U19658 (N_19658,N_19255,N_18545);
and U19659 (N_19659,N_19490,N_18390);
nor U19660 (N_19660,N_18054,N_18620);
nand U19661 (N_19661,N_18495,N_18918);
or U19662 (N_19662,N_18808,N_18972);
nand U19663 (N_19663,N_18947,N_18286);
xor U19664 (N_19664,N_19253,N_18343);
and U19665 (N_19665,N_19495,N_18242);
nand U19666 (N_19666,N_18223,N_19372);
xnor U19667 (N_19667,N_19229,N_18147);
and U19668 (N_19668,N_18331,N_18926);
or U19669 (N_19669,N_19147,N_19257);
and U19670 (N_19670,N_18766,N_18246);
nor U19671 (N_19671,N_18916,N_19163);
nor U19672 (N_19672,N_18210,N_18258);
nor U19673 (N_19673,N_19405,N_18776);
nand U19674 (N_19674,N_18694,N_18513);
xor U19675 (N_19675,N_19011,N_19322);
nor U19676 (N_19676,N_18035,N_19010);
xor U19677 (N_19677,N_19203,N_19389);
nand U19678 (N_19678,N_19132,N_18333);
and U19679 (N_19679,N_18026,N_18624);
and U19680 (N_19680,N_19452,N_19358);
nand U19681 (N_19681,N_19135,N_18430);
nor U19682 (N_19682,N_18263,N_19440);
xor U19683 (N_19683,N_19271,N_18161);
nand U19684 (N_19684,N_19462,N_18931);
or U19685 (N_19685,N_19239,N_18994);
xor U19686 (N_19686,N_18204,N_18253);
xor U19687 (N_19687,N_19401,N_18629);
or U19688 (N_19688,N_18831,N_18950);
and U19689 (N_19689,N_19446,N_19469);
nand U19690 (N_19690,N_19096,N_19078);
or U19691 (N_19691,N_18270,N_19076);
or U19692 (N_19692,N_19386,N_18913);
nor U19693 (N_19693,N_19000,N_18217);
xnor U19694 (N_19694,N_18289,N_19456);
nand U19695 (N_19695,N_18872,N_19464);
nand U19696 (N_19696,N_18908,N_19003);
nor U19697 (N_19697,N_18618,N_19468);
xor U19698 (N_19698,N_18956,N_18136);
or U19699 (N_19699,N_19316,N_19375);
xor U19700 (N_19700,N_18883,N_18642);
nor U19701 (N_19701,N_18777,N_18236);
nand U19702 (N_19702,N_19212,N_18648);
and U19703 (N_19703,N_18855,N_18378);
xnor U19704 (N_19704,N_18064,N_18142);
and U19705 (N_19705,N_18403,N_18124);
and U19706 (N_19706,N_18255,N_18429);
and U19707 (N_19707,N_18589,N_18386);
nand U19708 (N_19708,N_18316,N_18804);
nand U19709 (N_19709,N_18816,N_18414);
and U19710 (N_19710,N_18542,N_19023);
and U19711 (N_19711,N_18532,N_19043);
and U19712 (N_19712,N_18585,N_19174);
or U19713 (N_19713,N_18273,N_18101);
nand U19714 (N_19714,N_18056,N_19273);
xnor U19715 (N_19715,N_18247,N_18010);
xnor U19716 (N_19716,N_18865,N_19054);
and U19717 (N_19717,N_19303,N_18659);
and U19718 (N_19718,N_18463,N_19339);
nor U19719 (N_19719,N_18952,N_18257);
and U19720 (N_19720,N_18427,N_18575);
nor U19721 (N_19721,N_18238,N_18951);
nor U19722 (N_19722,N_19394,N_18141);
or U19723 (N_19723,N_19489,N_18769);
and U19724 (N_19724,N_18753,N_19480);
nand U19725 (N_19725,N_18548,N_18394);
xor U19726 (N_19726,N_18016,N_18770);
nor U19727 (N_19727,N_18300,N_18578);
xor U19728 (N_19728,N_19085,N_19252);
and U19729 (N_19729,N_18746,N_18622);
or U19730 (N_19730,N_19412,N_19473);
xor U19731 (N_19731,N_18105,N_19335);
nand U19732 (N_19732,N_19492,N_19034);
xnor U19733 (N_19733,N_18993,N_18597);
or U19734 (N_19734,N_18876,N_19334);
or U19735 (N_19735,N_18195,N_19046);
or U19736 (N_19736,N_19019,N_19083);
and U19737 (N_19737,N_18507,N_18177);
or U19738 (N_19738,N_18346,N_18061);
nor U19739 (N_19739,N_18570,N_18528);
or U19740 (N_19740,N_18164,N_18139);
and U19741 (N_19741,N_18292,N_19047);
or U19742 (N_19742,N_18469,N_18324);
nor U19743 (N_19743,N_18351,N_19413);
nor U19744 (N_19744,N_18820,N_19106);
nor U19745 (N_19745,N_19346,N_19377);
and U19746 (N_19746,N_18836,N_19014);
or U19747 (N_19747,N_18409,N_19162);
xor U19748 (N_19748,N_18423,N_19237);
xor U19749 (N_19749,N_18565,N_18997);
xor U19750 (N_19750,N_18877,N_19390);
xor U19751 (N_19751,N_19290,N_18579);
nor U19752 (N_19752,N_18580,N_19075);
nand U19753 (N_19753,N_18125,N_18380);
xor U19754 (N_19754,N_18256,N_18318);
nand U19755 (N_19755,N_18937,N_18264);
nand U19756 (N_19756,N_18670,N_18927);
xnor U19757 (N_19757,N_18971,N_18799);
xor U19758 (N_19758,N_18681,N_18554);
nor U19759 (N_19759,N_19353,N_19382);
or U19760 (N_19760,N_19180,N_18027);
and U19761 (N_19761,N_18750,N_18127);
nand U19762 (N_19762,N_19055,N_19282);
nand U19763 (N_19763,N_18756,N_18823);
xor U19764 (N_19764,N_18344,N_18473);
nand U19765 (N_19765,N_18606,N_18571);
or U19766 (N_19766,N_18232,N_18191);
or U19767 (N_19767,N_18953,N_18812);
xor U19768 (N_19768,N_18765,N_19475);
or U19769 (N_19769,N_19288,N_18451);
or U19770 (N_19770,N_18454,N_18013);
or U19771 (N_19771,N_18307,N_18843);
xnor U19772 (N_19772,N_19089,N_18516);
nand U19773 (N_19773,N_18562,N_19020);
nand U19774 (N_19774,N_19368,N_18095);
or U19775 (N_19775,N_19410,N_18266);
or U19776 (N_19776,N_19001,N_18296);
nor U19777 (N_19777,N_19487,N_18033);
nor U19778 (N_19778,N_19238,N_18801);
nand U19779 (N_19779,N_18803,N_18859);
or U19780 (N_19780,N_19122,N_18445);
nand U19781 (N_19781,N_18712,N_18830);
or U19782 (N_19782,N_19451,N_19117);
nor U19783 (N_19783,N_18948,N_18214);
and U19784 (N_19784,N_19423,N_19038);
or U19785 (N_19785,N_18609,N_18382);
and U19786 (N_19786,N_19095,N_18538);
nor U19787 (N_19787,N_18902,N_18240);
and U19788 (N_19788,N_18424,N_18421);
and U19789 (N_19789,N_18850,N_18272);
xor U19790 (N_19790,N_19012,N_18484);
or U19791 (N_19791,N_18728,N_18504);
nor U19792 (N_19792,N_18754,N_18371);
and U19793 (N_19793,N_18248,N_18946);
and U19794 (N_19794,N_18074,N_19044);
or U19795 (N_19795,N_18715,N_18975);
nand U19796 (N_19796,N_19158,N_19267);
xnor U19797 (N_19797,N_19289,N_18356);
or U19798 (N_19798,N_18833,N_18482);
nor U19799 (N_19799,N_19347,N_19067);
nand U19800 (N_19800,N_19063,N_18692);
nor U19801 (N_19801,N_18928,N_18861);
nor U19802 (N_19802,N_18925,N_18442);
and U19803 (N_19803,N_19447,N_18187);
xor U19804 (N_19804,N_18325,N_18720);
and U19805 (N_19805,N_18109,N_19443);
and U19806 (N_19806,N_18673,N_18172);
and U19807 (N_19807,N_18372,N_19005);
and U19808 (N_19808,N_19138,N_18935);
xnor U19809 (N_19809,N_18349,N_19256);
nand U19810 (N_19810,N_18283,N_18710);
and U19811 (N_19811,N_19201,N_19110);
or U19812 (N_19812,N_19333,N_19425);
xor U19813 (N_19813,N_18867,N_19091);
nand U19814 (N_19814,N_18917,N_18436);
nor U19815 (N_19815,N_18996,N_18837);
nand U19816 (N_19816,N_19157,N_18183);
xor U19817 (N_19817,N_19233,N_19042);
nand U19818 (N_19818,N_18676,N_18329);
nand U19819 (N_19819,N_18675,N_19130);
nand U19820 (N_19820,N_18813,N_18543);
nor U19821 (N_19821,N_18634,N_19213);
xnor U19822 (N_19822,N_18966,N_18057);
nor U19823 (N_19823,N_19112,N_19472);
nand U19824 (N_19824,N_18594,N_19188);
and U19825 (N_19825,N_19265,N_18239);
or U19826 (N_19826,N_18145,N_18208);
and U19827 (N_19827,N_18494,N_18851);
and U19828 (N_19828,N_18798,N_18982);
and U19829 (N_19829,N_19435,N_18868);
and U19830 (N_19830,N_18360,N_18215);
nand U19831 (N_19831,N_18392,N_18651);
xnor U19832 (N_19832,N_18121,N_18632);
and U19833 (N_19833,N_18206,N_18566);
and U19834 (N_19834,N_18062,N_19403);
xor U19835 (N_19835,N_18418,N_19183);
and U19836 (N_19836,N_18417,N_19027);
xnor U19837 (N_19837,N_19259,N_19204);
and U19838 (N_19838,N_18961,N_18118);
nand U19839 (N_19839,N_18024,N_19285);
or U19840 (N_19840,N_18797,N_19116);
nor U19841 (N_19841,N_18225,N_18352);
and U19842 (N_19842,N_18050,N_19341);
nor U19843 (N_19843,N_19309,N_19422);
or U19844 (N_19844,N_18262,N_18437);
and U19845 (N_19845,N_19167,N_18012);
and U19846 (N_19846,N_19416,N_18940);
xnor U19847 (N_19847,N_18102,N_19330);
and U19848 (N_19848,N_18254,N_18018);
nand U19849 (N_19849,N_18500,N_18401);
xor U19850 (N_19850,N_18148,N_18002);
xnor U19851 (N_19851,N_18508,N_18137);
nand U19852 (N_19852,N_18827,N_18824);
nor U19853 (N_19853,N_18932,N_18663);
or U19854 (N_19854,N_19058,N_18796);
or U19855 (N_19855,N_18885,N_18561);
or U19856 (N_19856,N_18025,N_19369);
and U19857 (N_19857,N_19053,N_19208);
xnor U19858 (N_19858,N_18764,N_18601);
or U19859 (N_19859,N_19457,N_18457);
nor U19860 (N_19860,N_19421,N_19077);
or U19861 (N_19861,N_18964,N_19442);
xnor U19862 (N_19862,N_18871,N_18419);
xnor U19863 (N_19863,N_18779,N_18432);
nor U19864 (N_19864,N_18396,N_18983);
or U19865 (N_19865,N_18505,N_18775);
and U19866 (N_19866,N_18697,N_18093);
nor U19867 (N_19867,N_18815,N_19307);
xor U19868 (N_19868,N_19186,N_18610);
xnor U19869 (N_19869,N_18608,N_19094);
nand U19870 (N_19870,N_19232,N_18480);
nor U19871 (N_19871,N_19050,N_18771);
and U19872 (N_19872,N_19101,N_19280);
and U19873 (N_19873,N_19254,N_18350);
or U19874 (N_19874,N_19278,N_18847);
and U19875 (N_19875,N_18630,N_18596);
xor U19876 (N_19876,N_18448,N_19249);
and U19877 (N_19877,N_18999,N_18310);
nor U19878 (N_19878,N_18903,N_18422);
or U19879 (N_19879,N_18829,N_19070);
nand U19880 (N_19880,N_18465,N_18555);
nor U19881 (N_19881,N_19268,N_18740);
nand U19882 (N_19882,N_19366,N_19428);
nor U19883 (N_19883,N_18471,N_18188);
nand U19884 (N_19884,N_18146,N_18178);
or U19885 (N_19885,N_18377,N_19344);
xnor U19886 (N_19886,N_19105,N_19342);
nor U19887 (N_19887,N_18958,N_19337);
xnor U19888 (N_19888,N_19177,N_18595);
and U19889 (N_19889,N_18082,N_19402);
and U19890 (N_19890,N_18176,N_18512);
or U19891 (N_19891,N_18159,N_18261);
and U19892 (N_19892,N_18718,N_18687);
nor U19893 (N_19893,N_18348,N_19430);
nor U19894 (N_19894,N_18839,N_18639);
xnor U19895 (N_19895,N_19497,N_18455);
nand U19896 (N_19896,N_18235,N_19397);
and U19897 (N_19897,N_18518,N_18660);
nor U19898 (N_19898,N_19470,N_18415);
or U19899 (N_19899,N_19178,N_19297);
or U19900 (N_19900,N_19084,N_18581);
nand U19901 (N_19901,N_18493,N_18474);
xor U19902 (N_19902,N_19387,N_18569);
and U19903 (N_19903,N_18822,N_18679);
xnor U19904 (N_19904,N_18864,N_19228);
nor U19905 (N_19905,N_18780,N_18374);
xor U19906 (N_19906,N_18492,N_18623);
nand U19907 (N_19907,N_19449,N_18962);
nor U19908 (N_19908,N_19260,N_18980);
nand U19909 (N_19909,N_18267,N_18821);
nand U19910 (N_19910,N_18282,N_18192);
and U19911 (N_19911,N_19392,N_18547);
xor U19912 (N_19912,N_18751,N_18987);
or U19913 (N_19913,N_19018,N_19209);
or U19914 (N_19914,N_18381,N_18860);
or U19915 (N_19915,N_18849,N_18234);
xor U19916 (N_19916,N_18295,N_19155);
nor U19917 (N_19917,N_19459,N_19279);
or U19918 (N_19918,N_18856,N_18305);
or U19919 (N_19919,N_18652,N_18680);
or U19920 (N_19920,N_19136,N_18963);
or U19921 (N_19921,N_19324,N_18853);
nor U19922 (N_19922,N_18130,N_19131);
and U19923 (N_19923,N_18499,N_18100);
nand U19924 (N_19924,N_18167,N_19007);
and U19925 (N_19925,N_18889,N_19109);
or U19926 (N_19926,N_19373,N_18106);
nand U19927 (N_19927,N_18173,N_18353);
or U19928 (N_19928,N_18986,N_18138);
nor U19929 (N_19929,N_19120,N_18472);
and U19930 (N_19930,N_18995,N_19248);
nand U19931 (N_19931,N_18723,N_18895);
or U19932 (N_19932,N_19483,N_18781);
or U19933 (N_19933,N_18668,N_18301);
xnor U19934 (N_19934,N_18244,N_18981);
and U19935 (N_19935,N_18231,N_19080);
and U19936 (N_19936,N_19409,N_19404);
xor U19937 (N_19937,N_19388,N_19059);
nor U19938 (N_19938,N_18375,N_18185);
nand U19939 (N_19939,N_18230,N_19045);
xnor U19940 (N_19940,N_18334,N_18160);
xnor U19941 (N_19941,N_19196,N_19286);
xor U19942 (N_19942,N_18912,N_18391);
nand U19943 (N_19943,N_19126,N_18332);
nor U19944 (N_19944,N_19272,N_18655);
xor U19945 (N_19945,N_18294,N_18312);
nor U19946 (N_19946,N_18893,N_18924);
nor U19947 (N_19947,N_19321,N_19102);
nand U19948 (N_19948,N_19315,N_19444);
and U19949 (N_19949,N_18713,N_19169);
and U19950 (N_19950,N_18603,N_18703);
xor U19951 (N_19951,N_18184,N_18941);
nand U19952 (N_19952,N_18092,N_18757);
nor U19953 (N_19953,N_19220,N_19134);
nand U19954 (N_19954,N_19395,N_19357);
nand U19955 (N_19955,N_19354,N_19300);
xor U19956 (N_19956,N_18260,N_18748);
and U19957 (N_19957,N_18408,N_18411);
xor U19958 (N_19958,N_18046,N_18008);
or U19959 (N_19959,N_19205,N_18251);
nand U19960 (N_19960,N_19244,N_19363);
xor U19961 (N_19961,N_18302,N_19037);
and U19962 (N_19962,N_18654,N_18383);
and U19963 (N_19963,N_19312,N_19277);
or U19964 (N_19964,N_18042,N_19262);
nand U19965 (N_19965,N_18647,N_18453);
and U19966 (N_19966,N_18920,N_18281);
and U19967 (N_19967,N_19436,N_19211);
nor U19968 (N_19968,N_18132,N_18506);
or U19969 (N_19969,N_19251,N_19242);
nor U19970 (N_19970,N_18459,N_18362);
or U19971 (N_19971,N_19378,N_18762);
or U19972 (N_19972,N_18722,N_19207);
and U19973 (N_19973,N_18845,N_19041);
nor U19974 (N_19974,N_18939,N_18501);
and U19975 (N_19975,N_18514,N_18517);
nand U19976 (N_19976,N_18306,N_19418);
or U19977 (N_19977,N_19199,N_19103);
or U19978 (N_19978,N_18416,N_18040);
xnor U19979 (N_19979,N_18792,N_18052);
and U19980 (N_19980,N_19093,N_18892);
nor U19981 (N_19981,N_18854,N_19400);
nor U19982 (N_19982,N_18122,N_19223);
or U19983 (N_19983,N_18084,N_19407);
or U19984 (N_19984,N_18342,N_18739);
nor U19985 (N_19985,N_18587,N_19221);
nor U19986 (N_19986,N_19226,N_19356);
or U19987 (N_19987,N_18733,N_18711);
xnor U19988 (N_19988,N_19039,N_18406);
nand U19989 (N_19989,N_18841,N_19304);
xor U19990 (N_19990,N_18015,N_19329);
xnor U19991 (N_19991,N_18104,N_18564);
and U19992 (N_19992,N_19293,N_18060);
nand U19993 (N_19993,N_18811,N_18328);
and U19994 (N_19994,N_18180,N_18549);
and U19995 (N_19995,N_19438,N_18081);
nor U19996 (N_19996,N_18510,N_18366);
or U19997 (N_19997,N_18327,N_19236);
xnor U19998 (N_19998,N_18783,N_18126);
and U19999 (N_19999,N_18702,N_18832);
nor U20000 (N_20000,N_18546,N_18103);
nor U20001 (N_20001,N_19150,N_19029);
nor U20002 (N_20002,N_19361,N_19159);
and U20003 (N_20003,N_18955,N_18452);
nor U20004 (N_20004,N_19071,N_18443);
nand U20005 (N_20005,N_18221,N_18491);
nor U20006 (N_20006,N_19467,N_19275);
nand U20007 (N_20007,N_19082,N_19219);
xor U20008 (N_20008,N_18643,N_18179);
and U20009 (N_20009,N_18464,N_19172);
xor U20010 (N_20010,N_19291,N_18527);
or U20011 (N_20011,N_19064,N_19482);
nor U20012 (N_20012,N_18633,N_18818);
and U20013 (N_20013,N_18243,N_18529);
nor U20014 (N_20014,N_19379,N_19028);
and U20015 (N_20015,N_18428,N_18943);
nor U20016 (N_20016,N_18393,N_18250);
nor U20017 (N_20017,N_19176,N_18802);
and U20018 (N_20018,N_18891,N_18973);
xor U20019 (N_20019,N_18045,N_19185);
or U20020 (N_20020,N_18716,N_18735);
or U20021 (N_20021,N_18450,N_19230);
nand U20022 (N_20022,N_18157,N_18583);
nor U20023 (N_20023,N_18605,N_18135);
xor U20024 (N_20024,N_18576,N_18992);
nand U20025 (N_20025,N_18866,N_18155);
nand U20026 (N_20026,N_18858,N_18881);
nand U20027 (N_20027,N_18795,N_18189);
nand U20028 (N_20028,N_18198,N_18117);
and U20029 (N_20029,N_18884,N_19061);
nand U20030 (N_20030,N_19385,N_19128);
nor U20031 (N_20031,N_18029,N_18657);
xnor U20032 (N_20032,N_18322,N_19274);
or U20033 (N_20033,N_18559,N_18638);
and U20034 (N_20034,N_18567,N_18619);
nor U20035 (N_20035,N_18398,N_19414);
nand U20036 (N_20036,N_18689,N_18190);
or U20037 (N_20037,N_18497,N_19325);
xor U20038 (N_20038,N_18944,N_19144);
nor U20039 (N_20039,N_18591,N_18120);
xnor U20040 (N_20040,N_18193,N_18410);
nor U20041 (N_20041,N_18425,N_18778);
nand U20042 (N_20042,N_18535,N_18309);
nor U20043 (N_20043,N_18534,N_19434);
or U20044 (N_20044,N_18129,N_18152);
and U20045 (N_20045,N_18626,N_19234);
and U20046 (N_20046,N_18817,N_18226);
nand U20047 (N_20047,N_18848,N_19036);
and U20048 (N_20048,N_19493,N_19148);
or U20049 (N_20049,N_19129,N_18399);
nand U20050 (N_20050,N_18761,N_19466);
and U20051 (N_20051,N_19022,N_18043);
nand U20052 (N_20052,N_19191,N_18069);
nor U20053 (N_20053,N_18874,N_18929);
xor U20054 (N_20054,N_18611,N_18695);
or U20055 (N_20055,N_19460,N_18336);
nand U20056 (N_20056,N_19181,N_18752);
xor U20057 (N_20057,N_19192,N_18708);
or U20058 (N_20058,N_18140,N_18194);
xor U20059 (N_20059,N_18065,N_19302);
or U20060 (N_20060,N_18835,N_18502);
nand U20061 (N_20061,N_18900,N_19419);
nand U20062 (N_20062,N_18321,N_18073);
nand U20063 (N_20063,N_18444,N_19266);
xnor U20064 (N_20064,N_18290,N_18852);
nor U20065 (N_20065,N_18773,N_18586);
or U20066 (N_20066,N_18096,N_18734);
or U20067 (N_20067,N_19301,N_18435);
nand U20068 (N_20068,N_18970,N_18772);
nor U20069 (N_20069,N_19145,N_19031);
nand U20070 (N_20070,N_19152,N_18524);
nand U20071 (N_20071,N_19125,N_18265);
nor U20072 (N_20072,N_18447,N_19142);
and U20073 (N_20073,N_18998,N_18227);
nand U20074 (N_20074,N_18684,N_18960);
nor U20075 (N_20075,N_18979,N_18658);
and U20076 (N_20076,N_18976,N_18616);
xor U20077 (N_20077,N_18402,N_18315);
xor U20078 (N_20078,N_18475,N_19195);
and U20079 (N_20079,N_18533,N_18553);
and U20080 (N_20080,N_18478,N_19164);
or U20081 (N_20081,N_18047,N_18834);
xor U20082 (N_20082,N_18044,N_19427);
xnor U20083 (N_20083,N_18072,N_18165);
nor U20084 (N_20084,N_18485,N_18249);
and U20085 (N_20085,N_18280,N_18641);
nand U20086 (N_20086,N_18786,N_19269);
and U20087 (N_20087,N_18275,N_19359);
and U20088 (N_20088,N_18174,N_19398);
or U20089 (N_20089,N_18873,N_19168);
xnor U20090 (N_20090,N_19243,N_19245);
xnor U20091 (N_20091,N_18886,N_19017);
and U20092 (N_20092,N_18537,N_19218);
nor U20093 (N_20093,N_18840,N_18028);
nand U20094 (N_20094,N_18558,N_19052);
nor U20095 (N_20095,N_19448,N_18440);
nand U20096 (N_20096,N_18339,N_19149);
or U20097 (N_20097,N_19433,N_18934);
nor U20098 (N_20098,N_19283,N_18196);
xor U20099 (N_20099,N_18039,N_18308);
or U20100 (N_20100,N_18228,N_19250);
and U20101 (N_20101,N_18017,N_18370);
or U20102 (N_20102,N_18826,N_19222);
nor U20103 (N_20103,N_18671,N_19073);
xnor U20104 (N_20104,N_18287,N_19270);
nor U20105 (N_20105,N_18059,N_18488);
and U20106 (N_20106,N_19026,N_19305);
nand U20107 (N_20107,N_18625,N_19175);
and U20108 (N_20108,N_18097,N_19024);
or U20109 (N_20109,N_19471,N_18171);
xor U20110 (N_20110,N_19081,N_18269);
and U20111 (N_20111,N_18707,N_19349);
or U20112 (N_20112,N_18271,N_18705);
nand U20113 (N_20113,N_19360,N_19166);
xnor U20114 (N_20114,N_19002,N_18978);
or U20115 (N_20115,N_18729,N_18087);
or U20116 (N_20116,N_18919,N_19124);
and U20117 (N_20117,N_18369,N_18637);
nor U20118 (N_20118,N_18323,N_18038);
or U20119 (N_20119,N_19114,N_18110);
or U20120 (N_20120,N_18070,N_18379);
or U20121 (N_20121,N_19224,N_18498);
and U20122 (N_20122,N_18907,N_19016);
nor U20123 (N_20123,N_19381,N_18202);
xnor U20124 (N_20124,N_18842,N_19348);
xor U20125 (N_20125,N_18863,N_18199);
nor U20126 (N_20126,N_19484,N_19056);
nor U20127 (N_20127,N_19108,N_19133);
or U20128 (N_20128,N_18433,N_18749);
or U20129 (N_20129,N_18607,N_19376);
nand U20130 (N_20130,N_19345,N_18688);
xor U20131 (N_20131,N_18030,N_19104);
or U20132 (N_20132,N_18319,N_19097);
or U20133 (N_20133,N_18487,N_18846);
and U20134 (N_20134,N_18588,N_18838);
and U20135 (N_20135,N_18020,N_18496);
or U20136 (N_20136,N_19485,N_18439);
nor U20137 (N_20137,N_18721,N_18788);
nand U20138 (N_20138,N_18170,N_18593);
nand U20139 (N_20139,N_18216,N_18080);
nand U20140 (N_20140,N_18755,N_19123);
xnor U20141 (N_20141,N_18388,N_18890);
xnor U20142 (N_20142,N_19488,N_19478);
and U20143 (N_20143,N_18742,N_19184);
or U20144 (N_20144,N_19317,N_18526);
and U20145 (N_20145,N_18259,N_19261);
nor U20146 (N_20146,N_18477,N_19450);
xor U20147 (N_20147,N_18311,N_18481);
and U20148 (N_20148,N_19194,N_19074);
nand U20149 (N_20149,N_18462,N_19217);
nor U20150 (N_20150,N_18051,N_19391);
nor U20151 (N_20151,N_19454,N_18169);
xnor U20152 (N_20152,N_19035,N_18154);
and U20153 (N_20153,N_19399,N_18000);
nand U20154 (N_20154,N_18441,N_18521);
nor U20155 (N_20155,N_18869,N_18698);
and U20156 (N_20156,N_19231,N_19090);
nand U20157 (N_20157,N_18212,N_18385);
xnor U20158 (N_20158,N_19069,N_18116);
or U20159 (N_20159,N_19380,N_19111);
xor U20160 (N_20160,N_18814,N_18114);
or U20161 (N_20161,N_19455,N_18887);
nor U20162 (N_20162,N_18959,N_18844);
xor U20163 (N_20163,N_18218,N_18420);
nand U20164 (N_20164,N_18784,N_19258);
and U20165 (N_20165,N_19299,N_18460);
and U20166 (N_20166,N_18922,N_19165);
xor U20167 (N_20167,N_18229,N_18479);
nor U20168 (N_20168,N_18706,N_18291);
xor U20169 (N_20169,N_18133,N_18071);
nor U20170 (N_20170,N_18615,N_18077);
or U20171 (N_20171,N_19057,N_18898);
nand U20172 (N_20172,N_19015,N_18314);
xnor U20173 (N_20173,N_18211,N_18509);
nand U20174 (N_20174,N_18878,N_18930);
and U20175 (N_20175,N_18741,N_18556);
and U20176 (N_20176,N_18066,N_19310);
xnor U20177 (N_20177,N_18405,N_18222);
xnor U20178 (N_20178,N_18143,N_19408);
or U20179 (N_20179,N_19336,N_19088);
and U20180 (N_20180,N_18880,N_19474);
nand U20181 (N_20181,N_18067,N_19004);
nor U20182 (N_20182,N_18909,N_18682);
and U20183 (N_20183,N_18635,N_18862);
nor U20184 (N_20184,N_18598,N_18163);
and U20185 (N_20185,N_18434,N_19461);
nand U20186 (N_20186,N_18317,N_19338);
nand U20187 (N_20187,N_18551,N_19498);
and U20188 (N_20188,N_18426,N_18736);
nor U20189 (N_20189,N_19206,N_18209);
nor U20190 (N_20190,N_19393,N_18407);
and U20191 (N_20191,N_18449,N_18395);
nor U20192 (N_20192,N_19323,N_18252);
and U20193 (N_20193,N_19331,N_19060);
and U20194 (N_20194,N_18743,N_18245);
or U20195 (N_20195,N_18376,N_18525);
nand U20196 (N_20196,N_18522,N_18326);
nand U20197 (N_20197,N_18412,N_18063);
nor U20198 (N_20198,N_18365,N_18150);
or U20199 (N_20199,N_18284,N_19481);
nand U20200 (N_20200,N_18357,N_18298);
nand U20201 (N_20201,N_18572,N_19173);
nand U20202 (N_20202,N_18058,N_19140);
nand U20203 (N_20203,N_19227,N_19351);
nand U20204 (N_20204,N_18662,N_18767);
or U20205 (N_20205,N_19295,N_18700);
nor U20206 (N_20206,N_19087,N_18990);
nor U20207 (N_20207,N_18737,N_18364);
or U20208 (N_20208,N_19214,N_18293);
xor U20209 (N_20209,N_19432,N_19314);
and U20210 (N_20210,N_18857,N_19210);
or U20211 (N_20211,N_18540,N_18933);
xnor U20212 (N_20212,N_18220,N_19494);
or U20213 (N_20213,N_18088,N_18151);
and U20214 (N_20214,N_19263,N_18131);
or U20215 (N_20215,N_18355,N_18985);
nor U20216 (N_20216,N_18656,N_18338);
xnor U20217 (N_20217,N_19187,N_18968);
and U20218 (N_20218,N_18207,N_18563);
and U20219 (N_20219,N_19384,N_18590);
nor U20220 (N_20220,N_19383,N_18091);
or U20221 (N_20221,N_18612,N_18584);
or U20222 (N_20222,N_18825,N_18076);
nand U20223 (N_20223,N_18467,N_18519);
or U20224 (N_20224,N_19143,N_19343);
nand U20225 (N_20225,N_18805,N_18725);
or U20226 (N_20226,N_18241,N_18413);
and U20227 (N_20227,N_19499,N_18672);
nand U20228 (N_20228,N_18724,N_18592);
and U20229 (N_20229,N_19021,N_19235);
or U20230 (N_20230,N_19115,N_18957);
or U20231 (N_20231,N_19141,N_18614);
xnor U20232 (N_20232,N_18113,N_18989);
nor U20233 (N_20233,N_19284,N_19098);
xor U20234 (N_20234,N_19328,N_18782);
nand U20235 (N_20235,N_18531,N_19161);
or U20236 (N_20236,N_18461,N_18745);
nor U20237 (N_20237,N_18032,N_18470);
xnor U20238 (N_20238,N_18313,N_18361);
xor U20239 (N_20239,N_19246,N_18037);
xor U20240 (N_20240,N_19160,N_19298);
nor U20241 (N_20241,N_19479,N_18613);
xor U20242 (N_20242,N_18552,N_18031);
nand U20243 (N_20243,N_18726,N_19241);
xnor U20244 (N_20244,N_18219,N_18557);
xor U20245 (N_20245,N_18621,N_18330);
or U20246 (N_20246,N_19146,N_18974);
or U20247 (N_20247,N_18446,N_18882);
or U20248 (N_20248,N_18108,N_19411);
xor U20249 (N_20249,N_18763,N_19276);
nor U20250 (N_20250,N_18053,N_18664);
and U20251 (N_20251,N_19393,N_18207);
nand U20252 (N_20252,N_18884,N_18518);
and U20253 (N_20253,N_19322,N_19122);
nor U20254 (N_20254,N_19175,N_18219);
xnor U20255 (N_20255,N_19135,N_19430);
nand U20256 (N_20256,N_18832,N_18274);
and U20257 (N_20257,N_18888,N_19128);
nor U20258 (N_20258,N_18839,N_19326);
or U20259 (N_20259,N_19167,N_18941);
nor U20260 (N_20260,N_18068,N_18611);
or U20261 (N_20261,N_18019,N_18098);
nor U20262 (N_20262,N_18416,N_18803);
or U20263 (N_20263,N_18991,N_18770);
or U20264 (N_20264,N_18276,N_18450);
nand U20265 (N_20265,N_19099,N_18112);
xor U20266 (N_20266,N_18230,N_19343);
nor U20267 (N_20267,N_19329,N_18542);
nand U20268 (N_20268,N_18326,N_18682);
and U20269 (N_20269,N_18636,N_18596);
nand U20270 (N_20270,N_18721,N_18612);
nand U20271 (N_20271,N_18723,N_18611);
or U20272 (N_20272,N_19247,N_18036);
and U20273 (N_20273,N_18886,N_18819);
and U20274 (N_20274,N_18739,N_19459);
or U20275 (N_20275,N_18901,N_18829);
nand U20276 (N_20276,N_19223,N_18910);
or U20277 (N_20277,N_18589,N_19048);
nor U20278 (N_20278,N_18472,N_18273);
nor U20279 (N_20279,N_18278,N_19280);
nand U20280 (N_20280,N_18796,N_19012);
and U20281 (N_20281,N_18602,N_18587);
nand U20282 (N_20282,N_18130,N_18749);
xnor U20283 (N_20283,N_18844,N_18046);
nor U20284 (N_20284,N_18879,N_19442);
nor U20285 (N_20285,N_18138,N_18913);
or U20286 (N_20286,N_18666,N_18644);
or U20287 (N_20287,N_18236,N_18304);
and U20288 (N_20288,N_18961,N_18800);
nor U20289 (N_20289,N_18700,N_19303);
and U20290 (N_20290,N_19014,N_19372);
nand U20291 (N_20291,N_19143,N_18650);
nand U20292 (N_20292,N_19086,N_18408);
xor U20293 (N_20293,N_19062,N_18913);
nor U20294 (N_20294,N_19011,N_19387);
nor U20295 (N_20295,N_18916,N_18970);
or U20296 (N_20296,N_19442,N_18056);
nand U20297 (N_20297,N_18422,N_18442);
or U20298 (N_20298,N_19013,N_18653);
or U20299 (N_20299,N_18718,N_18797);
nor U20300 (N_20300,N_18604,N_19206);
xor U20301 (N_20301,N_18134,N_19322);
nor U20302 (N_20302,N_18773,N_19427);
or U20303 (N_20303,N_18497,N_18817);
and U20304 (N_20304,N_18910,N_18973);
nor U20305 (N_20305,N_18443,N_18849);
nand U20306 (N_20306,N_18058,N_18797);
xnor U20307 (N_20307,N_19069,N_19402);
and U20308 (N_20308,N_18641,N_18213);
and U20309 (N_20309,N_18676,N_19144);
xor U20310 (N_20310,N_18021,N_18541);
nor U20311 (N_20311,N_18289,N_18143);
xor U20312 (N_20312,N_18322,N_18170);
and U20313 (N_20313,N_18977,N_18703);
nor U20314 (N_20314,N_19052,N_18684);
xor U20315 (N_20315,N_18731,N_18826);
nand U20316 (N_20316,N_19212,N_18460);
or U20317 (N_20317,N_18079,N_18988);
or U20318 (N_20318,N_19108,N_18719);
or U20319 (N_20319,N_19035,N_19130);
nor U20320 (N_20320,N_19008,N_18831);
nand U20321 (N_20321,N_19354,N_19346);
xnor U20322 (N_20322,N_19074,N_18165);
nand U20323 (N_20323,N_19440,N_19292);
nor U20324 (N_20324,N_18236,N_19035);
xnor U20325 (N_20325,N_19303,N_18315);
nand U20326 (N_20326,N_18101,N_18268);
and U20327 (N_20327,N_18754,N_18331);
nand U20328 (N_20328,N_18924,N_18474);
nor U20329 (N_20329,N_18062,N_19168);
or U20330 (N_20330,N_18377,N_19033);
or U20331 (N_20331,N_19452,N_18058);
and U20332 (N_20332,N_18861,N_18067);
nand U20333 (N_20333,N_18458,N_19212);
xor U20334 (N_20334,N_18736,N_18043);
xnor U20335 (N_20335,N_18793,N_19265);
or U20336 (N_20336,N_18031,N_18938);
or U20337 (N_20337,N_18314,N_18994);
and U20338 (N_20338,N_18902,N_19131);
nand U20339 (N_20339,N_18730,N_18263);
nand U20340 (N_20340,N_18863,N_18330);
nand U20341 (N_20341,N_18927,N_18065);
nand U20342 (N_20342,N_18384,N_18027);
or U20343 (N_20343,N_18478,N_19461);
or U20344 (N_20344,N_18030,N_18344);
nand U20345 (N_20345,N_18949,N_18440);
nor U20346 (N_20346,N_19371,N_19165);
or U20347 (N_20347,N_19180,N_18403);
nand U20348 (N_20348,N_19461,N_19203);
nor U20349 (N_20349,N_18102,N_19350);
and U20350 (N_20350,N_18695,N_18451);
or U20351 (N_20351,N_19425,N_19466);
nand U20352 (N_20352,N_18162,N_19155);
and U20353 (N_20353,N_18167,N_18927);
nor U20354 (N_20354,N_18121,N_18838);
nand U20355 (N_20355,N_18671,N_18748);
nand U20356 (N_20356,N_18505,N_18754);
or U20357 (N_20357,N_18445,N_18775);
xnor U20358 (N_20358,N_18036,N_18697);
and U20359 (N_20359,N_19059,N_18987);
nand U20360 (N_20360,N_18061,N_19269);
and U20361 (N_20361,N_19168,N_18050);
nor U20362 (N_20362,N_18009,N_18831);
nand U20363 (N_20363,N_18329,N_19499);
and U20364 (N_20364,N_18040,N_18472);
or U20365 (N_20365,N_19120,N_18563);
nor U20366 (N_20366,N_19400,N_18479);
and U20367 (N_20367,N_18652,N_18191);
xor U20368 (N_20368,N_18071,N_19465);
xor U20369 (N_20369,N_18429,N_19010);
and U20370 (N_20370,N_18173,N_18707);
nor U20371 (N_20371,N_18987,N_19094);
xor U20372 (N_20372,N_18899,N_19353);
xor U20373 (N_20373,N_18372,N_18048);
and U20374 (N_20374,N_19166,N_18181);
xnor U20375 (N_20375,N_18295,N_19444);
xor U20376 (N_20376,N_18277,N_18263);
and U20377 (N_20377,N_18606,N_18662);
or U20378 (N_20378,N_18721,N_18075);
and U20379 (N_20379,N_18792,N_19406);
nor U20380 (N_20380,N_19242,N_19155);
nor U20381 (N_20381,N_19082,N_18446);
xnor U20382 (N_20382,N_18589,N_19442);
xor U20383 (N_20383,N_19390,N_18269);
xor U20384 (N_20384,N_18650,N_19420);
or U20385 (N_20385,N_19112,N_18371);
and U20386 (N_20386,N_19462,N_19377);
or U20387 (N_20387,N_19031,N_18476);
or U20388 (N_20388,N_18025,N_18821);
xor U20389 (N_20389,N_19318,N_19048);
or U20390 (N_20390,N_18399,N_18250);
or U20391 (N_20391,N_18666,N_18764);
and U20392 (N_20392,N_19160,N_19135);
nand U20393 (N_20393,N_18589,N_19253);
xnor U20394 (N_20394,N_18029,N_18110);
or U20395 (N_20395,N_19309,N_18186);
xor U20396 (N_20396,N_18089,N_18212);
nand U20397 (N_20397,N_19476,N_18520);
nor U20398 (N_20398,N_19085,N_19166);
nor U20399 (N_20399,N_19457,N_18869);
nand U20400 (N_20400,N_19156,N_18860);
nor U20401 (N_20401,N_18243,N_19365);
and U20402 (N_20402,N_19253,N_19208);
and U20403 (N_20403,N_18195,N_19482);
or U20404 (N_20404,N_18171,N_19029);
or U20405 (N_20405,N_19438,N_19188);
and U20406 (N_20406,N_18993,N_18498);
or U20407 (N_20407,N_18426,N_18153);
xor U20408 (N_20408,N_18732,N_18687);
xor U20409 (N_20409,N_19352,N_19421);
nand U20410 (N_20410,N_19120,N_18690);
xor U20411 (N_20411,N_18266,N_19026);
nor U20412 (N_20412,N_18977,N_19197);
and U20413 (N_20413,N_18026,N_18072);
or U20414 (N_20414,N_18577,N_18763);
xnor U20415 (N_20415,N_19367,N_18485);
or U20416 (N_20416,N_19083,N_18091);
xnor U20417 (N_20417,N_18581,N_18906);
or U20418 (N_20418,N_19486,N_18583);
nand U20419 (N_20419,N_19146,N_18252);
or U20420 (N_20420,N_18792,N_18069);
and U20421 (N_20421,N_18139,N_18118);
or U20422 (N_20422,N_18442,N_19031);
nand U20423 (N_20423,N_18190,N_18879);
nor U20424 (N_20424,N_18083,N_19015);
nor U20425 (N_20425,N_18276,N_18501);
or U20426 (N_20426,N_18103,N_18501);
nand U20427 (N_20427,N_19217,N_18154);
or U20428 (N_20428,N_18832,N_18950);
and U20429 (N_20429,N_18626,N_18457);
or U20430 (N_20430,N_18424,N_18103);
and U20431 (N_20431,N_18477,N_18835);
or U20432 (N_20432,N_18054,N_18882);
nand U20433 (N_20433,N_19401,N_18312);
nand U20434 (N_20434,N_19136,N_18760);
nand U20435 (N_20435,N_19330,N_19085);
or U20436 (N_20436,N_18037,N_19188);
or U20437 (N_20437,N_19070,N_18229);
or U20438 (N_20438,N_18185,N_18361);
or U20439 (N_20439,N_18034,N_19410);
xor U20440 (N_20440,N_18553,N_19001);
and U20441 (N_20441,N_18468,N_19344);
xnor U20442 (N_20442,N_19070,N_18505);
or U20443 (N_20443,N_18597,N_19497);
nand U20444 (N_20444,N_18775,N_19167);
nand U20445 (N_20445,N_18327,N_18928);
nor U20446 (N_20446,N_19418,N_18446);
and U20447 (N_20447,N_18028,N_18365);
xnor U20448 (N_20448,N_18005,N_19260);
xnor U20449 (N_20449,N_19112,N_18725);
and U20450 (N_20450,N_18882,N_19378);
nor U20451 (N_20451,N_18251,N_18216);
or U20452 (N_20452,N_18375,N_18296);
xnor U20453 (N_20453,N_19480,N_18245);
nand U20454 (N_20454,N_18724,N_18491);
nand U20455 (N_20455,N_19065,N_18153);
or U20456 (N_20456,N_18153,N_18290);
nor U20457 (N_20457,N_18276,N_18546);
xor U20458 (N_20458,N_18820,N_18952);
and U20459 (N_20459,N_18838,N_18073);
nand U20460 (N_20460,N_18308,N_18910);
and U20461 (N_20461,N_18505,N_19499);
or U20462 (N_20462,N_18048,N_18149);
nand U20463 (N_20463,N_19411,N_18480);
nand U20464 (N_20464,N_18733,N_18155);
nor U20465 (N_20465,N_18049,N_18026);
and U20466 (N_20466,N_18714,N_19399);
or U20467 (N_20467,N_18310,N_19387);
nor U20468 (N_20468,N_18299,N_18454);
and U20469 (N_20469,N_19397,N_18301);
or U20470 (N_20470,N_18225,N_19434);
and U20471 (N_20471,N_19432,N_19403);
nor U20472 (N_20472,N_18042,N_18466);
xor U20473 (N_20473,N_18955,N_18169);
nand U20474 (N_20474,N_18045,N_18496);
nand U20475 (N_20475,N_18701,N_18142);
nand U20476 (N_20476,N_18392,N_18558);
nand U20477 (N_20477,N_18464,N_18244);
nor U20478 (N_20478,N_19427,N_19460);
nor U20479 (N_20479,N_18975,N_18520);
or U20480 (N_20480,N_19425,N_18635);
nand U20481 (N_20481,N_18135,N_18911);
or U20482 (N_20482,N_18457,N_18693);
nor U20483 (N_20483,N_18171,N_18995);
or U20484 (N_20484,N_18274,N_18483);
xor U20485 (N_20485,N_18247,N_18206);
nor U20486 (N_20486,N_18252,N_18266);
and U20487 (N_20487,N_18101,N_18823);
or U20488 (N_20488,N_18985,N_18807);
xor U20489 (N_20489,N_19331,N_18999);
and U20490 (N_20490,N_18918,N_18892);
or U20491 (N_20491,N_18919,N_18060);
or U20492 (N_20492,N_19011,N_19450);
and U20493 (N_20493,N_18949,N_18643);
xnor U20494 (N_20494,N_18576,N_19013);
or U20495 (N_20495,N_19360,N_19347);
nor U20496 (N_20496,N_18388,N_18149);
nor U20497 (N_20497,N_18487,N_18731);
and U20498 (N_20498,N_18334,N_19397);
nor U20499 (N_20499,N_19473,N_19449);
or U20500 (N_20500,N_19461,N_18372);
xnor U20501 (N_20501,N_18559,N_18869);
and U20502 (N_20502,N_18061,N_18820);
nand U20503 (N_20503,N_18308,N_18846);
nor U20504 (N_20504,N_18843,N_18372);
nor U20505 (N_20505,N_18124,N_19495);
and U20506 (N_20506,N_18619,N_18404);
and U20507 (N_20507,N_18156,N_19446);
or U20508 (N_20508,N_18820,N_18576);
nand U20509 (N_20509,N_18329,N_19301);
nand U20510 (N_20510,N_19227,N_19311);
nand U20511 (N_20511,N_18137,N_18337);
or U20512 (N_20512,N_18294,N_19440);
or U20513 (N_20513,N_18497,N_18122);
or U20514 (N_20514,N_19475,N_18576);
nor U20515 (N_20515,N_18683,N_19229);
and U20516 (N_20516,N_18566,N_18737);
nand U20517 (N_20517,N_19359,N_18702);
or U20518 (N_20518,N_19464,N_18841);
or U20519 (N_20519,N_18550,N_18269);
nor U20520 (N_20520,N_18111,N_18649);
xnor U20521 (N_20521,N_18815,N_18910);
nand U20522 (N_20522,N_19340,N_19223);
nand U20523 (N_20523,N_18226,N_18695);
xnor U20524 (N_20524,N_18258,N_19465);
nor U20525 (N_20525,N_19173,N_18457);
or U20526 (N_20526,N_19431,N_18531);
nand U20527 (N_20527,N_18808,N_18801);
and U20528 (N_20528,N_19109,N_19322);
nand U20529 (N_20529,N_18022,N_19089);
and U20530 (N_20530,N_18558,N_18635);
nor U20531 (N_20531,N_18732,N_19011);
nor U20532 (N_20532,N_18516,N_18570);
nand U20533 (N_20533,N_19487,N_18955);
nand U20534 (N_20534,N_18419,N_18288);
and U20535 (N_20535,N_19007,N_18746);
and U20536 (N_20536,N_19421,N_18648);
or U20537 (N_20537,N_18759,N_18295);
nand U20538 (N_20538,N_19210,N_18971);
and U20539 (N_20539,N_18874,N_18562);
xor U20540 (N_20540,N_19361,N_18901);
xor U20541 (N_20541,N_18309,N_18363);
xnor U20542 (N_20542,N_18860,N_18742);
or U20543 (N_20543,N_18958,N_18303);
nand U20544 (N_20544,N_18316,N_18828);
nand U20545 (N_20545,N_19179,N_18692);
nor U20546 (N_20546,N_18858,N_18049);
nand U20547 (N_20547,N_18996,N_19052);
or U20548 (N_20548,N_18778,N_19460);
or U20549 (N_20549,N_18120,N_18135);
and U20550 (N_20550,N_18924,N_18046);
or U20551 (N_20551,N_18326,N_18016);
or U20552 (N_20552,N_18498,N_18410);
or U20553 (N_20553,N_18588,N_18223);
or U20554 (N_20554,N_19258,N_18044);
and U20555 (N_20555,N_19202,N_19075);
nor U20556 (N_20556,N_18852,N_18546);
nand U20557 (N_20557,N_18033,N_19088);
nor U20558 (N_20558,N_19160,N_19334);
xnor U20559 (N_20559,N_18072,N_18687);
nand U20560 (N_20560,N_18196,N_19182);
nand U20561 (N_20561,N_18225,N_19328);
nand U20562 (N_20562,N_18017,N_18898);
or U20563 (N_20563,N_19064,N_19133);
or U20564 (N_20564,N_18578,N_18508);
and U20565 (N_20565,N_18017,N_18773);
or U20566 (N_20566,N_19204,N_18252);
or U20567 (N_20567,N_18728,N_18560);
or U20568 (N_20568,N_19318,N_19039);
nor U20569 (N_20569,N_18539,N_19179);
and U20570 (N_20570,N_18307,N_18656);
and U20571 (N_20571,N_19047,N_19207);
nand U20572 (N_20572,N_18347,N_18907);
or U20573 (N_20573,N_18303,N_18246);
xor U20574 (N_20574,N_18357,N_19020);
nor U20575 (N_20575,N_19332,N_18528);
nor U20576 (N_20576,N_19084,N_19146);
nor U20577 (N_20577,N_18377,N_19412);
xnor U20578 (N_20578,N_18423,N_18398);
or U20579 (N_20579,N_19062,N_18533);
xnor U20580 (N_20580,N_18214,N_19047);
and U20581 (N_20581,N_19234,N_19317);
xor U20582 (N_20582,N_19444,N_19013);
or U20583 (N_20583,N_18231,N_18687);
and U20584 (N_20584,N_18759,N_18521);
nor U20585 (N_20585,N_19132,N_18363);
nor U20586 (N_20586,N_19196,N_19452);
and U20587 (N_20587,N_19317,N_18415);
nor U20588 (N_20588,N_19442,N_18711);
nand U20589 (N_20589,N_18443,N_19494);
nand U20590 (N_20590,N_19419,N_18834);
and U20591 (N_20591,N_18694,N_18682);
and U20592 (N_20592,N_19415,N_18551);
and U20593 (N_20593,N_18814,N_18696);
nor U20594 (N_20594,N_18634,N_18970);
xnor U20595 (N_20595,N_18272,N_19166);
xor U20596 (N_20596,N_18628,N_18126);
nor U20597 (N_20597,N_18377,N_18439);
xor U20598 (N_20598,N_18474,N_18100);
nor U20599 (N_20599,N_18332,N_18576);
xnor U20600 (N_20600,N_18236,N_18900);
xor U20601 (N_20601,N_19379,N_18536);
and U20602 (N_20602,N_18807,N_18724);
and U20603 (N_20603,N_19002,N_19404);
nand U20604 (N_20604,N_18915,N_18994);
nor U20605 (N_20605,N_19156,N_18685);
or U20606 (N_20606,N_19073,N_18703);
xnor U20607 (N_20607,N_18358,N_18470);
and U20608 (N_20608,N_19129,N_19415);
or U20609 (N_20609,N_18077,N_19241);
nor U20610 (N_20610,N_18651,N_19158);
nand U20611 (N_20611,N_18831,N_19365);
and U20612 (N_20612,N_18178,N_18179);
nand U20613 (N_20613,N_18751,N_19227);
xnor U20614 (N_20614,N_19015,N_19330);
nor U20615 (N_20615,N_18471,N_19376);
nor U20616 (N_20616,N_19390,N_18603);
or U20617 (N_20617,N_18031,N_19282);
nand U20618 (N_20618,N_19274,N_18833);
xnor U20619 (N_20619,N_18496,N_19268);
or U20620 (N_20620,N_18010,N_19306);
nor U20621 (N_20621,N_19387,N_19333);
nand U20622 (N_20622,N_19079,N_18699);
nor U20623 (N_20623,N_18770,N_18381);
nor U20624 (N_20624,N_19120,N_19156);
or U20625 (N_20625,N_18224,N_18144);
nand U20626 (N_20626,N_18262,N_19193);
xor U20627 (N_20627,N_19272,N_19465);
and U20628 (N_20628,N_18545,N_19439);
or U20629 (N_20629,N_18134,N_18303);
nor U20630 (N_20630,N_19021,N_18452);
and U20631 (N_20631,N_18234,N_18742);
or U20632 (N_20632,N_19172,N_18568);
and U20633 (N_20633,N_18340,N_19185);
xor U20634 (N_20634,N_19113,N_19302);
nand U20635 (N_20635,N_18620,N_18736);
xor U20636 (N_20636,N_19095,N_18452);
or U20637 (N_20637,N_18951,N_19249);
and U20638 (N_20638,N_18522,N_19001);
or U20639 (N_20639,N_19094,N_18884);
nand U20640 (N_20640,N_18713,N_19449);
nor U20641 (N_20641,N_18021,N_18126);
nand U20642 (N_20642,N_19021,N_19495);
nor U20643 (N_20643,N_18208,N_19003);
and U20644 (N_20644,N_19339,N_18539);
nand U20645 (N_20645,N_19176,N_19202);
xnor U20646 (N_20646,N_19189,N_18988);
nand U20647 (N_20647,N_18011,N_18850);
xnor U20648 (N_20648,N_19252,N_19143);
or U20649 (N_20649,N_18743,N_19474);
xnor U20650 (N_20650,N_18563,N_19017);
and U20651 (N_20651,N_19076,N_18047);
nand U20652 (N_20652,N_19097,N_19210);
nand U20653 (N_20653,N_19051,N_18141);
and U20654 (N_20654,N_18008,N_19204);
xnor U20655 (N_20655,N_19029,N_18298);
xor U20656 (N_20656,N_18281,N_19104);
and U20657 (N_20657,N_19065,N_18099);
nor U20658 (N_20658,N_18005,N_18256);
nor U20659 (N_20659,N_19057,N_19027);
nor U20660 (N_20660,N_18856,N_18558);
and U20661 (N_20661,N_18207,N_19033);
nand U20662 (N_20662,N_18907,N_18229);
or U20663 (N_20663,N_19151,N_18029);
or U20664 (N_20664,N_19414,N_18731);
nor U20665 (N_20665,N_18293,N_18493);
nand U20666 (N_20666,N_18769,N_19377);
and U20667 (N_20667,N_19230,N_18319);
and U20668 (N_20668,N_19397,N_18653);
nor U20669 (N_20669,N_19375,N_18295);
xnor U20670 (N_20670,N_18183,N_19189);
nand U20671 (N_20671,N_18464,N_18570);
nor U20672 (N_20672,N_18787,N_18471);
and U20673 (N_20673,N_19125,N_18760);
or U20674 (N_20674,N_19485,N_19342);
xnor U20675 (N_20675,N_18559,N_19009);
or U20676 (N_20676,N_18039,N_18239);
and U20677 (N_20677,N_19453,N_18228);
or U20678 (N_20678,N_18132,N_18802);
nand U20679 (N_20679,N_19401,N_18061);
nand U20680 (N_20680,N_19025,N_18130);
xor U20681 (N_20681,N_18654,N_18407);
nand U20682 (N_20682,N_19019,N_18174);
or U20683 (N_20683,N_19478,N_18157);
and U20684 (N_20684,N_18144,N_18267);
or U20685 (N_20685,N_19010,N_18493);
nor U20686 (N_20686,N_18224,N_18867);
or U20687 (N_20687,N_19448,N_19022);
and U20688 (N_20688,N_18986,N_18122);
or U20689 (N_20689,N_19277,N_19349);
or U20690 (N_20690,N_18652,N_19257);
or U20691 (N_20691,N_18901,N_19466);
nand U20692 (N_20692,N_18021,N_18303);
nor U20693 (N_20693,N_18671,N_18005);
xnor U20694 (N_20694,N_19130,N_19359);
nand U20695 (N_20695,N_18106,N_19220);
or U20696 (N_20696,N_19442,N_18482);
and U20697 (N_20697,N_19249,N_19398);
or U20698 (N_20698,N_18237,N_18815);
nor U20699 (N_20699,N_18308,N_19225);
nor U20700 (N_20700,N_19132,N_18228);
nor U20701 (N_20701,N_19300,N_18877);
nand U20702 (N_20702,N_18952,N_18667);
nor U20703 (N_20703,N_19186,N_18487);
and U20704 (N_20704,N_18769,N_18605);
xnor U20705 (N_20705,N_18186,N_19073);
nor U20706 (N_20706,N_19268,N_19179);
nor U20707 (N_20707,N_19386,N_19070);
nor U20708 (N_20708,N_18808,N_18101);
xnor U20709 (N_20709,N_19156,N_18466);
nand U20710 (N_20710,N_18816,N_19377);
nand U20711 (N_20711,N_18989,N_18056);
or U20712 (N_20712,N_18153,N_19230);
nand U20713 (N_20713,N_18003,N_18475);
xor U20714 (N_20714,N_18173,N_18885);
and U20715 (N_20715,N_19004,N_18730);
nor U20716 (N_20716,N_18346,N_18263);
xor U20717 (N_20717,N_18333,N_19068);
or U20718 (N_20718,N_19296,N_18602);
nor U20719 (N_20719,N_19198,N_18641);
xor U20720 (N_20720,N_18364,N_18221);
nor U20721 (N_20721,N_18796,N_19021);
nor U20722 (N_20722,N_19140,N_19152);
nand U20723 (N_20723,N_18282,N_18342);
xnor U20724 (N_20724,N_18034,N_18795);
xor U20725 (N_20725,N_18634,N_18826);
nor U20726 (N_20726,N_18133,N_18420);
xor U20727 (N_20727,N_18274,N_18767);
or U20728 (N_20728,N_18408,N_18453);
and U20729 (N_20729,N_18263,N_19489);
nand U20730 (N_20730,N_18808,N_19411);
nand U20731 (N_20731,N_18262,N_18653);
and U20732 (N_20732,N_18213,N_19449);
nor U20733 (N_20733,N_18824,N_18825);
nor U20734 (N_20734,N_19107,N_19373);
or U20735 (N_20735,N_19126,N_19377);
nor U20736 (N_20736,N_18794,N_19475);
xnor U20737 (N_20737,N_19036,N_19143);
or U20738 (N_20738,N_18966,N_18097);
nor U20739 (N_20739,N_18721,N_18704);
nor U20740 (N_20740,N_19409,N_19302);
or U20741 (N_20741,N_18389,N_18902);
nand U20742 (N_20742,N_18365,N_18808);
or U20743 (N_20743,N_18593,N_18136);
nor U20744 (N_20744,N_18119,N_18671);
xnor U20745 (N_20745,N_18070,N_19073);
xnor U20746 (N_20746,N_18569,N_18210);
or U20747 (N_20747,N_19381,N_18851);
or U20748 (N_20748,N_19146,N_18759);
nand U20749 (N_20749,N_19439,N_18311);
and U20750 (N_20750,N_19350,N_18107);
nand U20751 (N_20751,N_18330,N_18670);
and U20752 (N_20752,N_19300,N_18568);
nor U20753 (N_20753,N_18169,N_19129);
nand U20754 (N_20754,N_19117,N_18292);
xnor U20755 (N_20755,N_18606,N_18435);
xnor U20756 (N_20756,N_18097,N_19092);
xnor U20757 (N_20757,N_18186,N_18055);
and U20758 (N_20758,N_19157,N_19213);
nor U20759 (N_20759,N_18589,N_19462);
nand U20760 (N_20760,N_19084,N_18757);
nand U20761 (N_20761,N_18028,N_19101);
or U20762 (N_20762,N_19075,N_18965);
nand U20763 (N_20763,N_19066,N_19100);
nand U20764 (N_20764,N_18273,N_18383);
nand U20765 (N_20765,N_18064,N_19440);
and U20766 (N_20766,N_19397,N_19106);
nor U20767 (N_20767,N_18725,N_18357);
nand U20768 (N_20768,N_18999,N_18785);
xnor U20769 (N_20769,N_19496,N_18425);
nand U20770 (N_20770,N_18310,N_18707);
nand U20771 (N_20771,N_18993,N_18906);
xor U20772 (N_20772,N_18992,N_18594);
and U20773 (N_20773,N_18803,N_19442);
and U20774 (N_20774,N_18220,N_19333);
nor U20775 (N_20775,N_18423,N_18460);
nand U20776 (N_20776,N_19118,N_18360);
and U20777 (N_20777,N_19293,N_19345);
nor U20778 (N_20778,N_18882,N_19449);
or U20779 (N_20779,N_18743,N_19293);
nor U20780 (N_20780,N_18992,N_18507);
or U20781 (N_20781,N_18005,N_18061);
and U20782 (N_20782,N_18568,N_19011);
nor U20783 (N_20783,N_18464,N_18537);
xor U20784 (N_20784,N_18804,N_19295);
or U20785 (N_20785,N_19152,N_19284);
nand U20786 (N_20786,N_19491,N_19052);
and U20787 (N_20787,N_19324,N_18443);
xor U20788 (N_20788,N_18330,N_19488);
xor U20789 (N_20789,N_19366,N_18078);
nor U20790 (N_20790,N_18781,N_18632);
or U20791 (N_20791,N_18187,N_19395);
xnor U20792 (N_20792,N_19270,N_18908);
or U20793 (N_20793,N_18761,N_19210);
or U20794 (N_20794,N_18550,N_19259);
nand U20795 (N_20795,N_18066,N_18784);
nand U20796 (N_20796,N_18357,N_18576);
nand U20797 (N_20797,N_19372,N_18414);
and U20798 (N_20798,N_19361,N_19105);
and U20799 (N_20799,N_18161,N_18002);
nor U20800 (N_20800,N_18268,N_18354);
and U20801 (N_20801,N_18690,N_18865);
and U20802 (N_20802,N_18374,N_19343);
nand U20803 (N_20803,N_19215,N_18258);
nand U20804 (N_20804,N_18884,N_19092);
nand U20805 (N_20805,N_18049,N_19085);
and U20806 (N_20806,N_18635,N_19234);
or U20807 (N_20807,N_19034,N_18576);
nand U20808 (N_20808,N_18758,N_18840);
nor U20809 (N_20809,N_18265,N_19285);
xor U20810 (N_20810,N_19398,N_18874);
nor U20811 (N_20811,N_19344,N_18440);
nor U20812 (N_20812,N_19412,N_18283);
nand U20813 (N_20813,N_19176,N_18152);
nor U20814 (N_20814,N_18226,N_19412);
nor U20815 (N_20815,N_19111,N_19183);
nand U20816 (N_20816,N_18445,N_18006);
and U20817 (N_20817,N_18461,N_19126);
nand U20818 (N_20818,N_18932,N_19152);
nand U20819 (N_20819,N_18891,N_18442);
and U20820 (N_20820,N_18352,N_18596);
nor U20821 (N_20821,N_18352,N_18623);
and U20822 (N_20822,N_19070,N_18556);
nor U20823 (N_20823,N_18416,N_19280);
xnor U20824 (N_20824,N_18759,N_19038);
nand U20825 (N_20825,N_18945,N_19159);
xor U20826 (N_20826,N_19377,N_18694);
nand U20827 (N_20827,N_18096,N_18746);
xor U20828 (N_20828,N_19210,N_18303);
and U20829 (N_20829,N_18498,N_18727);
nor U20830 (N_20830,N_18468,N_18719);
nor U20831 (N_20831,N_19012,N_18578);
nand U20832 (N_20832,N_19174,N_19185);
xor U20833 (N_20833,N_19065,N_18085);
nand U20834 (N_20834,N_18362,N_18518);
nor U20835 (N_20835,N_19061,N_18605);
nor U20836 (N_20836,N_19198,N_19017);
or U20837 (N_20837,N_18965,N_18949);
xor U20838 (N_20838,N_19037,N_18066);
and U20839 (N_20839,N_18484,N_19277);
or U20840 (N_20840,N_18519,N_19065);
nand U20841 (N_20841,N_18188,N_18538);
or U20842 (N_20842,N_18524,N_18249);
nor U20843 (N_20843,N_18582,N_19281);
nor U20844 (N_20844,N_18001,N_19378);
xor U20845 (N_20845,N_18932,N_19384);
nor U20846 (N_20846,N_18673,N_18056);
nand U20847 (N_20847,N_19491,N_19288);
nor U20848 (N_20848,N_18684,N_18440);
nor U20849 (N_20849,N_19016,N_19233);
nor U20850 (N_20850,N_18998,N_18357);
nor U20851 (N_20851,N_18795,N_18599);
xnor U20852 (N_20852,N_18027,N_19186);
nand U20853 (N_20853,N_18236,N_18482);
nor U20854 (N_20854,N_18808,N_19450);
nand U20855 (N_20855,N_18608,N_18309);
xor U20856 (N_20856,N_18954,N_18496);
or U20857 (N_20857,N_18005,N_18156);
nor U20858 (N_20858,N_18633,N_18327);
nand U20859 (N_20859,N_18029,N_18312);
and U20860 (N_20860,N_19429,N_18745);
xor U20861 (N_20861,N_19058,N_18750);
nand U20862 (N_20862,N_18315,N_18612);
nand U20863 (N_20863,N_18904,N_19256);
xor U20864 (N_20864,N_19285,N_18509);
nor U20865 (N_20865,N_18408,N_18040);
and U20866 (N_20866,N_18060,N_18651);
xor U20867 (N_20867,N_18364,N_18291);
or U20868 (N_20868,N_18779,N_19263);
or U20869 (N_20869,N_19357,N_19204);
and U20870 (N_20870,N_18258,N_18795);
xor U20871 (N_20871,N_18472,N_18801);
nor U20872 (N_20872,N_19325,N_19058);
or U20873 (N_20873,N_18969,N_19138);
and U20874 (N_20874,N_18103,N_18472);
and U20875 (N_20875,N_18264,N_19236);
xor U20876 (N_20876,N_19401,N_19243);
and U20877 (N_20877,N_18360,N_18103);
nor U20878 (N_20878,N_19172,N_18370);
nand U20879 (N_20879,N_18818,N_18651);
nor U20880 (N_20880,N_19258,N_19027);
or U20881 (N_20881,N_18036,N_18817);
xor U20882 (N_20882,N_18565,N_18553);
nand U20883 (N_20883,N_19476,N_19012);
xor U20884 (N_20884,N_18425,N_18772);
nand U20885 (N_20885,N_18373,N_18193);
xor U20886 (N_20886,N_18950,N_18214);
or U20887 (N_20887,N_18762,N_19423);
nor U20888 (N_20888,N_18672,N_18805);
nor U20889 (N_20889,N_19058,N_18911);
or U20890 (N_20890,N_19041,N_18855);
nor U20891 (N_20891,N_18840,N_19408);
or U20892 (N_20892,N_18661,N_18866);
nand U20893 (N_20893,N_19020,N_19447);
and U20894 (N_20894,N_19479,N_18308);
nor U20895 (N_20895,N_18839,N_19351);
nor U20896 (N_20896,N_18013,N_19155);
xnor U20897 (N_20897,N_18529,N_19439);
nor U20898 (N_20898,N_18073,N_18390);
nor U20899 (N_20899,N_18623,N_18727);
and U20900 (N_20900,N_18504,N_19300);
nor U20901 (N_20901,N_19046,N_19466);
nor U20902 (N_20902,N_18050,N_19250);
nand U20903 (N_20903,N_18829,N_18381);
nor U20904 (N_20904,N_18652,N_19125);
nand U20905 (N_20905,N_19440,N_19009);
nand U20906 (N_20906,N_18782,N_18266);
xor U20907 (N_20907,N_18855,N_18084);
nand U20908 (N_20908,N_18874,N_18237);
xor U20909 (N_20909,N_19020,N_18959);
or U20910 (N_20910,N_18408,N_18272);
xnor U20911 (N_20911,N_18312,N_18402);
nand U20912 (N_20912,N_18662,N_18968);
or U20913 (N_20913,N_18644,N_18691);
nor U20914 (N_20914,N_18437,N_18734);
xnor U20915 (N_20915,N_18624,N_18539);
nand U20916 (N_20916,N_18900,N_18051);
xnor U20917 (N_20917,N_18473,N_19122);
nand U20918 (N_20918,N_18949,N_19427);
or U20919 (N_20919,N_18168,N_18422);
nor U20920 (N_20920,N_19398,N_18211);
xor U20921 (N_20921,N_18602,N_18870);
xor U20922 (N_20922,N_19488,N_18427);
xor U20923 (N_20923,N_19334,N_19359);
and U20924 (N_20924,N_18543,N_18897);
nor U20925 (N_20925,N_19278,N_18632);
nand U20926 (N_20926,N_19211,N_18306);
nor U20927 (N_20927,N_19405,N_18981);
xor U20928 (N_20928,N_18773,N_18194);
xor U20929 (N_20929,N_19368,N_19447);
or U20930 (N_20930,N_18115,N_18941);
or U20931 (N_20931,N_19480,N_18531);
nor U20932 (N_20932,N_18581,N_18944);
nand U20933 (N_20933,N_18372,N_19000);
xnor U20934 (N_20934,N_18804,N_18221);
xnor U20935 (N_20935,N_18498,N_19347);
and U20936 (N_20936,N_18205,N_18482);
xor U20937 (N_20937,N_18973,N_18210);
nand U20938 (N_20938,N_18161,N_18303);
xnor U20939 (N_20939,N_19283,N_19197);
nor U20940 (N_20940,N_18997,N_19147);
or U20941 (N_20941,N_18843,N_18834);
or U20942 (N_20942,N_18887,N_19050);
xnor U20943 (N_20943,N_18605,N_19352);
and U20944 (N_20944,N_19316,N_18999);
and U20945 (N_20945,N_18599,N_19383);
nand U20946 (N_20946,N_18391,N_18473);
or U20947 (N_20947,N_18489,N_18363);
or U20948 (N_20948,N_18272,N_18458);
and U20949 (N_20949,N_18063,N_19407);
xnor U20950 (N_20950,N_19406,N_18542);
nand U20951 (N_20951,N_18928,N_18503);
nor U20952 (N_20952,N_18035,N_19426);
xnor U20953 (N_20953,N_19051,N_18167);
nor U20954 (N_20954,N_19345,N_19186);
nand U20955 (N_20955,N_18471,N_18850);
nand U20956 (N_20956,N_19257,N_19094);
nor U20957 (N_20957,N_19206,N_18463);
or U20958 (N_20958,N_19078,N_19330);
xnor U20959 (N_20959,N_19201,N_19358);
nand U20960 (N_20960,N_19051,N_18173);
xor U20961 (N_20961,N_18217,N_19325);
nand U20962 (N_20962,N_18038,N_18770);
or U20963 (N_20963,N_18344,N_18849);
or U20964 (N_20964,N_18259,N_19325);
nor U20965 (N_20965,N_18966,N_18615);
nor U20966 (N_20966,N_18165,N_18193);
xor U20967 (N_20967,N_18138,N_18930);
or U20968 (N_20968,N_18077,N_18087);
and U20969 (N_20969,N_18022,N_19068);
nor U20970 (N_20970,N_19197,N_19469);
and U20971 (N_20971,N_18470,N_18943);
and U20972 (N_20972,N_18600,N_18701);
and U20973 (N_20973,N_19260,N_18454);
nand U20974 (N_20974,N_18998,N_18619);
and U20975 (N_20975,N_19326,N_18677);
and U20976 (N_20976,N_18743,N_18891);
or U20977 (N_20977,N_19233,N_19364);
nand U20978 (N_20978,N_18065,N_18604);
and U20979 (N_20979,N_18170,N_18606);
nand U20980 (N_20980,N_19210,N_19465);
or U20981 (N_20981,N_18605,N_19166);
or U20982 (N_20982,N_19238,N_19201);
xor U20983 (N_20983,N_18408,N_18686);
nand U20984 (N_20984,N_18441,N_18212);
nand U20985 (N_20985,N_18756,N_18999);
or U20986 (N_20986,N_19395,N_18737);
nor U20987 (N_20987,N_18451,N_18621);
nor U20988 (N_20988,N_18311,N_18527);
nor U20989 (N_20989,N_19003,N_18912);
xor U20990 (N_20990,N_18726,N_18183);
and U20991 (N_20991,N_19345,N_18140);
and U20992 (N_20992,N_18999,N_19371);
and U20993 (N_20993,N_18573,N_19479);
and U20994 (N_20994,N_18986,N_18644);
nor U20995 (N_20995,N_18015,N_18564);
or U20996 (N_20996,N_18990,N_19253);
nand U20997 (N_20997,N_18576,N_19062);
nand U20998 (N_20998,N_19106,N_19214);
nand U20999 (N_20999,N_19438,N_19180);
and U21000 (N_21000,N_20049,N_19721);
or U21001 (N_21001,N_19698,N_20168);
nor U21002 (N_21002,N_20899,N_19792);
nor U21003 (N_21003,N_19837,N_20266);
and U21004 (N_21004,N_19677,N_20896);
xor U21005 (N_21005,N_19811,N_20632);
xor U21006 (N_21006,N_19529,N_20914);
xnor U21007 (N_21007,N_20047,N_20620);
nor U21008 (N_21008,N_19901,N_20677);
and U21009 (N_21009,N_20234,N_19625);
xnor U21010 (N_21010,N_20495,N_20935);
or U21011 (N_21011,N_20441,N_19937);
or U21012 (N_21012,N_20415,N_20088);
nand U21013 (N_21013,N_19528,N_19858);
and U21014 (N_21014,N_20449,N_20253);
or U21015 (N_21015,N_20068,N_20530);
nor U21016 (N_21016,N_20925,N_20455);
or U21017 (N_21017,N_19820,N_20547);
nand U21018 (N_21018,N_20522,N_20348);
and U21019 (N_21019,N_20431,N_20172);
nor U21020 (N_21020,N_19533,N_19801);
or U21021 (N_21021,N_20447,N_19601);
nor U21022 (N_21022,N_19657,N_19594);
nor U21023 (N_21023,N_19644,N_20135);
nor U21024 (N_21024,N_20341,N_19946);
xnor U21025 (N_21025,N_20216,N_19587);
nand U21026 (N_21026,N_20351,N_20148);
nand U21027 (N_21027,N_20195,N_20802);
xnor U21028 (N_21028,N_20332,N_19852);
or U21029 (N_21029,N_19932,N_20854);
and U21030 (N_21030,N_20395,N_20772);
or U21031 (N_21031,N_20983,N_20911);
or U21032 (N_21032,N_19616,N_20523);
nand U21033 (N_21033,N_20967,N_20895);
nand U21034 (N_21034,N_20577,N_20394);
nor U21035 (N_21035,N_20964,N_20612);
xor U21036 (N_21036,N_19526,N_19910);
nor U21037 (N_21037,N_19595,N_20885);
nand U21038 (N_21038,N_19544,N_20053);
and U21039 (N_21039,N_20735,N_19695);
nor U21040 (N_21040,N_20477,N_19621);
or U21041 (N_21041,N_20786,N_19753);
or U21042 (N_21042,N_19553,N_20258);
or U21043 (N_21043,N_20104,N_20132);
xnor U21044 (N_21044,N_20506,N_20963);
and U21045 (N_21045,N_20862,N_19715);
or U21046 (N_21046,N_19936,N_19527);
nor U21047 (N_21047,N_20936,N_20666);
xnor U21048 (N_21048,N_19978,N_20569);
nor U21049 (N_21049,N_20947,N_20466);
and U21050 (N_21050,N_19797,N_20169);
nor U21051 (N_21051,N_20217,N_20407);
and U21052 (N_21052,N_20634,N_20099);
nand U21053 (N_21053,N_20614,N_19796);
and U21054 (N_21054,N_20278,N_19531);
and U21055 (N_21055,N_20091,N_20405);
nor U21056 (N_21056,N_20003,N_20417);
and U21057 (N_21057,N_19726,N_20762);
xor U21058 (N_21058,N_20568,N_20685);
and U21059 (N_21059,N_20669,N_20374);
nand U21060 (N_21060,N_19517,N_20815);
nand U21061 (N_21061,N_19502,N_20820);
or U21062 (N_21062,N_19506,N_20887);
nand U21063 (N_21063,N_20363,N_19536);
xor U21064 (N_21064,N_20814,N_19777);
nand U21065 (N_21065,N_19923,N_19520);
or U21066 (N_21066,N_20376,N_20458);
nor U21067 (N_21067,N_20763,N_20442);
nand U21068 (N_21068,N_20870,N_19821);
nand U21069 (N_21069,N_20048,N_20776);
and U21070 (N_21070,N_20838,N_19975);
and U21071 (N_21071,N_20354,N_20636);
and U21072 (N_21072,N_20052,N_20187);
xor U21073 (N_21073,N_19738,N_20412);
or U21074 (N_21074,N_19793,N_19831);
nand U21075 (N_21075,N_20603,N_19573);
or U21076 (N_21076,N_20328,N_20849);
nand U21077 (N_21077,N_20098,N_20750);
nor U21078 (N_21078,N_20753,N_19805);
nor U21079 (N_21079,N_20828,N_20630);
nor U21080 (N_21080,N_20290,N_20504);
and U21081 (N_21081,N_20615,N_20212);
xor U21082 (N_21082,N_20336,N_19762);
or U21083 (N_21083,N_19739,N_20327);
and U21084 (N_21084,N_20650,N_20136);
xor U21085 (N_21085,N_20832,N_20400);
or U21086 (N_21086,N_20661,N_20489);
xor U21087 (N_21087,N_20659,N_20611);
nand U21088 (N_21088,N_19586,N_20714);
nand U21089 (N_21089,N_20360,N_20557);
and U21090 (N_21090,N_20652,N_20060);
nand U21091 (N_21091,N_20399,N_19897);
nor U21092 (N_21092,N_20573,N_20528);
or U21093 (N_21093,N_20939,N_19948);
nand U21094 (N_21094,N_20289,N_19769);
and U21095 (N_21095,N_19909,N_20641);
nand U21096 (N_21096,N_20196,N_20825);
xor U21097 (N_21097,N_20841,N_19547);
nor U21098 (N_21098,N_20368,N_20457);
nand U21099 (N_21099,N_20170,N_19825);
and U21100 (N_21100,N_20715,N_20416);
nand U21101 (N_21101,N_20233,N_20987);
nand U21102 (N_21102,N_20688,N_20241);
nand U21103 (N_21103,N_20749,N_19955);
nor U21104 (N_21104,N_20892,N_19731);
or U21105 (N_21105,N_20302,N_20796);
and U21106 (N_21106,N_20260,N_20141);
or U21107 (N_21107,N_20338,N_20094);
or U21108 (N_21108,N_20004,N_19645);
xnor U21109 (N_21109,N_19578,N_20282);
xnor U21110 (N_21110,N_19708,N_19914);
and U21111 (N_21111,N_20497,N_20009);
nor U21112 (N_21112,N_19511,N_19600);
nand U21113 (N_21113,N_19917,N_20675);
xor U21114 (N_21114,N_20792,N_19944);
or U21115 (N_21115,N_19921,N_19829);
and U21116 (N_21116,N_20272,N_20460);
xnor U21117 (N_21117,N_20462,N_20519);
nand U21118 (N_21118,N_19765,N_20056);
nor U21119 (N_21119,N_20432,N_19760);
or U21120 (N_21120,N_20668,N_20888);
and U21121 (N_21121,N_20662,N_20345);
nand U21122 (N_21122,N_20469,N_20700);
or U21123 (N_21123,N_20909,N_20687);
nor U21124 (N_21124,N_20891,N_19892);
and U21125 (N_21125,N_20686,N_20508);
nand U21126 (N_21126,N_20798,N_20954);
or U21127 (N_21127,N_20836,N_20193);
nand U21128 (N_21128,N_19570,N_20534);
nand U21129 (N_21129,N_20034,N_20191);
or U21130 (N_21130,N_20719,N_20128);
or U21131 (N_21131,N_20230,N_20767);
and U21132 (N_21132,N_20186,N_20576);
nand U21133 (N_21133,N_19809,N_20218);
and U21134 (N_21134,N_19919,N_19579);
nor U21135 (N_21135,N_20766,N_20387);
xor U21136 (N_21136,N_20134,N_20257);
nand U21137 (N_21137,N_20222,N_19860);
xor U21138 (N_21138,N_19856,N_19729);
nand U21139 (N_21139,N_19803,N_20246);
nor U21140 (N_21140,N_20799,N_20592);
and U21141 (N_21141,N_19754,N_20959);
and U21142 (N_21142,N_19552,N_20574);
or U21143 (N_21143,N_19588,N_19840);
and U21144 (N_21144,N_19626,N_19709);
and U21145 (N_21145,N_20850,N_19795);
and U21146 (N_21146,N_19734,N_20153);
and U21147 (N_21147,N_20251,N_20130);
and U21148 (N_21148,N_20985,N_19942);
nor U21149 (N_21149,N_20424,N_20177);
or U21150 (N_21150,N_20001,N_20520);
or U21151 (N_21151,N_20627,N_20404);
or U21152 (N_21152,N_20924,N_20751);
and U21153 (N_21153,N_19717,N_19778);
and U21154 (N_21154,N_19664,N_20100);
nand U21155 (N_21155,N_20044,N_19999);
nor U21156 (N_21156,N_20894,N_20065);
or U21157 (N_21157,N_20537,N_20331);
or U21158 (N_21158,N_19624,N_20918);
nand U21159 (N_21159,N_19641,N_20024);
xnor U21160 (N_21160,N_20140,N_19655);
and U21161 (N_21161,N_20079,N_20090);
or U21162 (N_21162,N_20950,N_20554);
nor U21163 (N_21163,N_19742,N_20274);
nand U21164 (N_21164,N_19539,N_20518);
nand U21165 (N_21165,N_20043,N_20882);
nand U21166 (N_21166,N_20402,N_19808);
or U21167 (N_21167,N_20821,N_20538);
or U21168 (N_21168,N_20966,N_19913);
nor U21169 (N_21169,N_19679,N_19973);
nand U21170 (N_21170,N_19611,N_20998);
or U21171 (N_21171,N_20645,N_20463);
and U21172 (N_21172,N_20237,N_19776);
and U21173 (N_21173,N_19962,N_20549);
nand U21174 (N_21174,N_19918,N_20335);
or U21175 (N_21175,N_20635,N_20531);
xnor U21176 (N_21176,N_20294,N_20361);
nor U21177 (N_21177,N_20955,N_20639);
nand U21178 (N_21178,N_20107,N_20840);
or U21179 (N_21179,N_20931,N_20901);
and U21180 (N_21180,N_20865,N_20898);
xor U21181 (N_21181,N_19814,N_20689);
nor U21182 (N_21182,N_19927,N_20834);
nand U21183 (N_21183,N_20525,N_19972);
nand U21184 (N_21184,N_20667,N_20968);
or U21185 (N_21185,N_20926,N_20558);
or U21186 (N_21186,N_19564,N_20622);
nand U21187 (N_21187,N_20031,N_20581);
and U21188 (N_21188,N_20422,N_20378);
xor U21189 (N_21189,N_19929,N_20929);
xnor U21190 (N_21190,N_20900,N_19841);
nand U21191 (N_21191,N_19538,N_20372);
xor U21192 (N_21192,N_20874,N_20490);
and U21193 (N_21193,N_20481,N_19543);
or U21194 (N_21194,N_19646,N_19741);
or U21195 (N_21195,N_19806,N_19675);
and U21196 (N_21196,N_20309,N_19690);
or U21197 (N_21197,N_19710,N_20124);
xnor U21198 (N_21198,N_20949,N_20316);
nand U21199 (N_21199,N_20300,N_20026);
or U21200 (N_21200,N_20129,N_20224);
and U21201 (N_21201,N_20103,N_20919);
xnor U21202 (N_21202,N_19969,N_20190);
nor U21203 (N_21203,N_20265,N_20349);
or U21204 (N_21204,N_20702,N_19866);
xnor U21205 (N_21205,N_19749,N_19783);
or U21206 (N_21206,N_20252,N_19562);
nand U21207 (N_21207,N_20151,N_20268);
and U21208 (N_21208,N_20511,N_19876);
and U21209 (N_21209,N_20121,N_20994);
xor U21210 (N_21210,N_20369,N_20638);
nand U21211 (N_21211,N_20479,N_20228);
xnor U21212 (N_21212,N_19525,N_20464);
or U21213 (N_21213,N_19782,N_19571);
and U21214 (N_21214,N_20733,N_20775);
xor U21215 (N_21215,N_19583,N_20209);
nor U21216 (N_21216,N_20419,N_20500);
nand U21217 (N_21217,N_19702,N_19557);
or U21218 (N_21218,N_20958,N_20198);
nor U21219 (N_21219,N_20742,N_20683);
nor U21220 (N_21220,N_20414,N_20277);
or U21221 (N_21221,N_20080,N_19683);
xnor U21222 (N_21222,N_20055,N_20250);
nor U21223 (N_21223,N_20889,N_20308);
or U21224 (N_21224,N_20002,N_19712);
xnor U21225 (N_21225,N_19874,N_19643);
and U21226 (N_21226,N_20197,N_20629);
or U21227 (N_21227,N_19967,N_20072);
and U21228 (N_21228,N_20851,N_20516);
nor U21229 (N_21229,N_20058,N_20513);
or U21230 (N_21230,N_19505,N_19771);
and U21231 (N_21231,N_20752,N_20303);
nand U21232 (N_21232,N_19680,N_19569);
nand U21233 (N_21233,N_20108,N_20243);
nor U21234 (N_21234,N_20712,N_20708);
or U21235 (N_21235,N_20319,N_19745);
and U21236 (N_21236,N_19963,N_19576);
and U21237 (N_21237,N_19691,N_20773);
or U21238 (N_21238,N_19839,N_19891);
xor U21239 (N_21239,N_19639,N_19790);
xor U21240 (N_21240,N_19950,N_20541);
nor U21241 (N_21241,N_20498,N_20934);
xor U21242 (N_21242,N_20709,N_20176);
nand U21243 (N_21243,N_20096,N_20219);
xnor U21244 (N_21244,N_20470,N_20310);
and U21245 (N_21245,N_19697,N_20928);
xor U21246 (N_21246,N_19908,N_20305);
nand U21247 (N_21247,N_19609,N_20904);
xor U21248 (N_21248,N_19733,N_19668);
nor U21249 (N_21249,N_20232,N_20208);
nor U21250 (N_21250,N_19599,N_20721);
or U21251 (N_21251,N_20586,N_20609);
nor U21252 (N_21252,N_19747,N_20684);
xnor U21253 (N_21253,N_19836,N_19575);
or U21254 (N_21254,N_20467,N_19509);
nand U21255 (N_21255,N_20306,N_20077);
or U21256 (N_21256,N_19849,N_19758);
nor U21257 (N_21257,N_20724,N_19898);
nor U21258 (N_21258,N_20383,N_20656);
nand U21259 (N_21259,N_19642,N_19584);
nor U21260 (N_21260,N_20435,N_20548);
nor U21261 (N_21261,N_20138,N_19510);
xnor U21262 (N_21262,N_20855,N_20120);
xor U21263 (N_21263,N_20015,N_20720);
nor U21264 (N_21264,N_20736,N_19947);
nor U21265 (N_21265,N_19991,N_20203);
or U21266 (N_21266,N_20981,N_20366);
xor U21267 (N_21267,N_19530,N_19902);
xnor U21268 (N_21268,N_19682,N_20014);
and U21269 (N_21269,N_20391,N_20384);
and U21270 (N_21270,N_19514,N_20322);
xnor U21271 (N_21271,N_20800,N_20254);
xor U21272 (N_21272,N_19723,N_20403);
or U21273 (N_21273,N_20174,N_20550);
xnor U21274 (N_21274,N_20073,N_20754);
and U21275 (N_21275,N_20608,N_19925);
or U21276 (N_21276,N_19663,N_20990);
nand U21277 (N_21277,N_19537,N_19830);
nand U21278 (N_21278,N_19983,N_20494);
nor U21279 (N_21279,N_19623,N_20633);
nor U21280 (N_21280,N_20823,N_19686);
and U21281 (N_21281,N_20364,N_20941);
nand U21282 (N_21282,N_19722,N_19951);
and U21283 (N_21283,N_20595,N_20381);
nor U21284 (N_21284,N_20006,N_20373);
nor U21285 (N_21285,N_20621,N_20235);
nor U21286 (N_21286,N_20822,N_19501);
or U21287 (N_21287,N_20734,N_19546);
and U21288 (N_21288,N_20587,N_20081);
nor U21289 (N_21289,N_19627,N_20488);
and U21290 (N_21290,N_19684,N_20582);
or U21291 (N_21291,N_19842,N_19662);
or U21292 (N_21292,N_19992,N_20758);
and U21293 (N_21293,N_20710,N_19581);
and U21294 (N_21294,N_20816,N_19693);
nand U21295 (N_21295,N_19816,N_20651);
nand U21296 (N_21296,N_20122,N_20281);
nor U21297 (N_21297,N_19784,N_20672);
nand U21298 (N_21298,N_20510,N_19613);
and U21299 (N_21299,N_20562,N_20160);
nand U21300 (N_21300,N_20917,N_20594);
or U21301 (N_21301,N_19629,N_20897);
or U21302 (N_21302,N_20201,N_20439);
or U21303 (N_21303,N_19632,N_19622);
and U21304 (N_21304,N_19890,N_20564);
nand U21305 (N_21305,N_19545,N_19615);
nor U21306 (N_21306,N_20401,N_20676);
and U21307 (N_21307,N_19988,N_20681);
or U21308 (N_21308,N_20358,N_19807);
xor U21309 (N_21309,N_20061,N_20739);
nand U21310 (N_21310,N_20385,N_20357);
xnor U21311 (N_21311,N_20591,N_20748);
and U21312 (N_21312,N_19945,N_20083);
xor U21313 (N_21313,N_20829,N_19519);
xnor U21314 (N_21314,N_20480,N_20299);
nor U21315 (N_21315,N_19879,N_20790);
or U21316 (N_21316,N_20741,N_20386);
and U21317 (N_21317,N_19672,N_20301);
or U21318 (N_21318,N_20451,N_20330);
xor U21319 (N_21319,N_19798,N_19648);
nand U21320 (N_21320,N_20082,N_19713);
xor U21321 (N_21321,N_20040,N_20916);
and U21322 (N_21322,N_20379,N_19877);
nand U21323 (N_21323,N_20101,N_19563);
and U21324 (N_21324,N_20596,N_20264);
xnor U21325 (N_21325,N_19549,N_20054);
or U21326 (N_21326,N_20810,N_20943);
and U21327 (N_21327,N_20476,N_20215);
xor U21328 (N_21328,N_20315,N_20852);
nor U21329 (N_21329,N_19888,N_20037);
and U21330 (N_21330,N_20437,N_20291);
and U21331 (N_21331,N_19521,N_20788);
and U21332 (N_21332,N_20042,N_19503);
nor U21333 (N_21333,N_20370,N_20655);
nand U21334 (N_21334,N_19922,N_20613);
xor U21335 (N_21335,N_19755,N_20050);
nand U21336 (N_21336,N_20872,N_20071);
nor U21337 (N_21337,N_20161,N_20755);
nand U21338 (N_21338,N_19705,N_20743);
xnor U21339 (N_21339,N_20869,N_20746);
xor U21340 (N_21340,N_20567,N_19912);
or U21341 (N_21341,N_19787,N_20062);
nand U21342 (N_21342,N_19985,N_20344);
and U21343 (N_21343,N_19899,N_20848);
and U21344 (N_21344,N_20933,N_20337);
or U21345 (N_21345,N_19746,N_20324);
xor U21346 (N_21346,N_19968,N_20286);
xnor U21347 (N_21347,N_20013,N_20540);
xnor U21348 (N_21348,N_20678,N_20262);
nand U21349 (N_21349,N_20199,N_20304);
or U21350 (N_21350,N_19904,N_19822);
xor U21351 (N_21351,N_20493,N_20146);
nand U21352 (N_21352,N_20078,N_20539);
and U21353 (N_21353,N_19590,N_20382);
nor U21354 (N_21354,N_19631,N_20877);
nand U21355 (N_21355,N_19554,N_20318);
nand U21356 (N_21356,N_19979,N_20867);
nor U21357 (N_21357,N_20857,N_20915);
nand U21358 (N_21358,N_20843,N_20842);
or U21359 (N_21359,N_20142,N_20988);
and U21360 (N_21360,N_19670,N_20962);
nand U21361 (N_21361,N_19804,N_20975);
or U21362 (N_21362,N_20565,N_20809);
nand U21363 (N_21363,N_20007,N_20965);
nand U21364 (N_21364,N_19728,N_20737);
and U21365 (N_21365,N_20827,N_20626);
nand U21366 (N_21366,N_20946,N_20893);
nand U21367 (N_21367,N_20163,N_20923);
or U21368 (N_21368,N_20350,N_20273);
xnor U21369 (N_21369,N_20325,N_20542);
xnor U21370 (N_21370,N_20041,N_20692);
nor U21371 (N_21371,N_20427,N_20317);
nor U21372 (N_21372,N_19850,N_20646);
nand U21373 (N_21373,N_20993,N_19938);
nor U21374 (N_21374,N_20057,N_19522);
or U21375 (N_21375,N_19534,N_19886);
and U21376 (N_21376,N_19513,N_20856);
and U21377 (N_21377,N_19943,N_20440);
or U21378 (N_21378,N_20927,N_20205);
xor U21379 (N_21379,N_20601,N_19916);
or U21380 (N_21380,N_20572,N_20529);
nor U21381 (N_21381,N_19652,N_20147);
and U21382 (N_21382,N_20269,N_20509);
and U21383 (N_21383,N_20863,N_20438);
xnor U21384 (N_21384,N_20178,N_19714);
nor U21385 (N_21385,N_19561,N_20871);
nor U21386 (N_21386,N_20214,N_19884);
nand U21387 (N_21387,N_20207,N_20543);
or U21388 (N_21388,N_20181,N_19628);
xnor U21389 (N_21389,N_20499,N_20145);
nor U21390 (N_21390,N_20512,N_20027);
nor U21391 (N_21391,N_20211,N_20606);
or U21392 (N_21392,N_19794,N_19567);
xor U21393 (N_21393,N_20535,N_19920);
nor U21394 (N_21394,N_19960,N_19614);
nor U21395 (N_21395,N_19685,N_20271);
nor U21396 (N_21396,N_19558,N_20579);
or U21397 (N_21397,N_19833,N_20756);
and U21398 (N_21398,N_20296,N_20297);
nor U21399 (N_21399,N_20903,N_20960);
nor U21400 (N_21400,N_19752,N_20977);
nand U21401 (N_21401,N_20256,N_20673);
nor U21402 (N_21402,N_20314,N_19889);
xor U21403 (N_21403,N_20456,N_19961);
or U21404 (N_21404,N_20210,N_20410);
nor U21405 (N_21405,N_20443,N_20846);
or U21406 (N_21406,N_19924,N_19666);
nor U21407 (N_21407,N_20760,N_20768);
and U21408 (N_21408,N_20298,N_19870);
xor U21409 (N_21409,N_20182,N_20359);
nor U21410 (N_21410,N_20797,N_20227);
nor U21411 (N_21411,N_20165,N_19676);
nand U21412 (N_21412,N_20355,N_19812);
nand U21413 (N_21413,N_20409,N_20021);
nor U21414 (N_21414,N_20022,N_20032);
xnor U21415 (N_21415,N_19550,N_20571);
xor U21416 (N_21416,N_19989,N_20236);
xor U21417 (N_21417,N_19634,N_19949);
nand U21418 (N_21418,N_20194,N_20649);
xor U21419 (N_21419,N_19618,N_20831);
nand U21420 (N_21420,N_20745,N_20334);
or U21421 (N_21421,N_20783,N_19857);
nand U21422 (N_21422,N_19681,N_19802);
nand U21423 (N_21423,N_20905,N_19810);
nand U21424 (N_21424,N_20902,N_20551);
nand U21425 (N_21425,N_19848,N_19774);
and U21426 (N_21426,N_20570,N_19737);
nor U21427 (N_21427,N_20794,N_20206);
and U21428 (N_21428,N_20245,N_19518);
nand U21429 (N_21429,N_20853,N_20801);
or U21430 (N_21430,N_19987,N_20389);
nand U21431 (N_21431,N_20944,N_20890);
or U21432 (N_21432,N_20747,N_19751);
or U21433 (N_21433,N_20039,N_20883);
or U21434 (N_21434,N_20450,N_19523);
and U21435 (N_21435,N_19846,N_20703);
and U21436 (N_21436,N_19743,N_20942);
xnor U21437 (N_21437,N_20657,N_19720);
or U21438 (N_21438,N_20392,N_20818);
and U21439 (N_21439,N_20940,N_20175);
or U21440 (N_21440,N_20095,N_19535);
or U21441 (N_21441,N_19871,N_20010);
nor U21442 (N_21442,N_19881,N_20578);
nor U21443 (N_21443,N_19582,N_20459);
nor U21444 (N_21444,N_20362,N_20732);
or U21445 (N_21445,N_20804,N_19864);
xnor U21446 (N_21446,N_20276,N_20616);
nor U21447 (N_21447,N_20292,N_20461);
nand U21448 (N_21448,N_19838,N_20320);
nor U21449 (N_21449,N_20553,N_20604);
or U21450 (N_21450,N_20496,N_20283);
or U21451 (N_21451,N_20448,N_19926);
nand U21452 (N_21452,N_20782,N_20280);
xnor U21453 (N_21453,N_20559,N_19667);
or U21454 (N_21454,N_19637,N_19964);
nor U21455 (N_21455,N_19786,N_19761);
nor U21456 (N_21456,N_20220,N_19669);
or U21457 (N_21457,N_20602,N_19735);
and U21458 (N_21458,N_20131,N_20225);
nand U21459 (N_21459,N_20371,N_19993);
nor U21460 (N_21460,N_19748,N_20847);
nor U21461 (N_21461,N_20259,N_20473);
and U21462 (N_21462,N_20787,N_19568);
and U21463 (N_21463,N_20589,N_20653);
nor U21464 (N_21464,N_20434,N_20817);
or U21465 (N_21465,N_20482,N_20430);
or U21466 (N_21466,N_20221,N_19701);
nand U21467 (N_21467,N_20507,N_20670);
nand U21468 (N_21468,N_19865,N_20046);
nand U21469 (N_21469,N_20599,N_19930);
nor U21470 (N_21470,N_19872,N_19934);
nor U21471 (N_21471,N_20491,N_20696);
nand U21472 (N_21472,N_19704,N_19556);
and U21473 (N_21473,N_20664,N_20418);
and U21474 (N_21474,N_20029,N_20793);
nand U21475 (N_21475,N_19559,N_20390);
nor U21476 (N_21476,N_19608,N_19661);
nor U21477 (N_21477,N_20556,N_20575);
or U21478 (N_21478,N_19508,N_20426);
and U21479 (N_21479,N_20969,N_19855);
or U21480 (N_21480,N_20223,N_20726);
xor U21481 (N_21481,N_19727,N_19656);
and U21482 (N_21482,N_20485,N_20682);
nor U21483 (N_21483,N_20008,N_19935);
xor U21484 (N_21484,N_19647,N_19966);
nor U21485 (N_21485,N_19791,N_19998);
and U21486 (N_21486,N_20204,N_20167);
nor U21487 (N_21487,N_20560,N_19818);
nor U21488 (N_21488,N_19744,N_19566);
or U21489 (N_21489,N_20938,N_20546);
or U21490 (N_21490,N_20974,N_20654);
or U21491 (N_21491,N_19903,N_20270);
nor U21492 (N_21492,N_20979,N_20429);
nand U21493 (N_21493,N_20555,N_19980);
and U21494 (N_21494,N_20835,N_20515);
xor U21495 (N_21495,N_19853,N_20119);
or U21496 (N_21496,N_20116,N_20102);
nor U21497 (N_21497,N_19653,N_20527);
xnor U21498 (N_21498,N_20805,N_19635);
and U21499 (N_21499,N_20478,N_20671);
and U21500 (N_21500,N_20992,N_20033);
nor U21501 (N_21501,N_19994,N_19835);
or U21502 (N_21502,N_19823,N_19885);
and U21503 (N_21503,N_20113,N_20143);
nand U21504 (N_21504,N_20106,N_20020);
xnor U21505 (N_21505,N_20860,N_19931);
nand U21506 (N_21506,N_19580,N_20566);
and U21507 (N_21507,N_20665,N_19990);
nand U21508 (N_21508,N_19906,N_20833);
nor U21509 (N_21509,N_20859,N_20069);
and U21510 (N_21510,N_20038,N_19772);
xnor U21511 (N_21511,N_20097,N_20408);
and U21512 (N_21512,N_19766,N_20624);
xor U21513 (N_21513,N_20213,N_19828);
or U21514 (N_21514,N_19671,N_19939);
and U21515 (N_21515,N_20738,N_19716);
xnor U21516 (N_21516,N_19707,N_20789);
xnor U21517 (N_21517,N_19928,N_19799);
or U21518 (N_21518,N_20023,N_19813);
and U21519 (N_21519,N_20875,N_20761);
and U21520 (N_21520,N_20723,N_20533);
nor U21521 (N_21521,N_20806,N_20631);
and U21522 (N_21522,N_20740,N_20718);
or U21523 (N_21523,N_19541,N_19894);
or U21524 (N_21524,N_20779,N_20619);
xnor U21525 (N_21525,N_19834,N_20770);
or U21526 (N_21526,N_20179,N_20680);
and U21527 (N_21527,N_19785,N_19658);
nor U21528 (N_21528,N_20200,N_19996);
xnor U21529 (N_21529,N_20580,N_19605);
and U21530 (N_21530,N_20123,N_20706);
and U21531 (N_21531,N_19540,N_20144);
or U21532 (N_21532,N_20545,N_19706);
or U21533 (N_21533,N_20995,N_20293);
or U21534 (N_21534,N_19941,N_20873);
nor U21535 (N_21535,N_20625,N_20731);
nand U21536 (N_21536,N_19863,N_20413);
nand U21537 (N_21537,N_20980,N_20694);
nor U21538 (N_21538,N_19598,N_20238);
xnor U21539 (N_21539,N_20285,N_20725);
nor U21540 (N_21540,N_20468,N_19878);
nor U21541 (N_21541,N_20991,N_20000);
xnor U21542 (N_21542,N_20247,N_20628);
xor U21543 (N_21543,N_19574,N_20644);
or U21544 (N_21544,N_20311,N_20728);
nand U21545 (N_21545,N_20879,N_19606);
nand U21546 (N_21546,N_19775,N_20445);
xnor U21547 (N_21547,N_20713,N_20164);
xor U21548 (N_21548,N_20780,N_20192);
xnor U21549 (N_21549,N_20312,N_20089);
nand U21550 (N_21550,N_19532,N_19887);
nor U21551 (N_21551,N_19861,N_20830);
or U21552 (N_21552,N_20640,N_19515);
nand U21553 (N_21553,N_20858,N_19699);
nor U21554 (N_21554,N_20249,N_19593);
nand U21555 (N_21555,N_20396,N_20663);
nand U21556 (N_21556,N_20005,N_19824);
xor U21557 (N_21557,N_19957,N_20184);
nor U21558 (N_21558,N_20397,N_19620);
nand U21559 (N_21559,N_20398,N_20948);
xor U21560 (N_21560,N_20791,N_20876);
nor U21561 (N_21561,N_19832,N_20242);
nor U21562 (N_21562,N_20411,N_20826);
nor U21563 (N_21563,N_20552,N_20287);
and U21564 (N_21564,N_20110,N_20084);
xor U21565 (N_21565,N_20922,N_20261);
nand U21566 (N_21566,N_19696,N_20154);
or U21567 (N_21567,N_20333,N_20453);
nand U21568 (N_21568,N_19893,N_20126);
xor U21569 (N_21569,N_20326,N_20813);
xnor U21570 (N_21570,N_20016,N_20781);
xnor U21571 (N_21571,N_20824,N_19597);
nand U21572 (N_21572,N_20807,N_20536);
nor U21573 (N_21573,N_19585,N_20059);
nor U21574 (N_21574,N_20035,N_19859);
or U21575 (N_21575,N_19630,N_20393);
nor U21576 (N_21576,N_20839,N_20421);
or U21577 (N_21577,N_20526,N_20295);
xor U21578 (N_21578,N_20452,N_20971);
and U21579 (N_21579,N_20377,N_19572);
xor U21580 (N_21580,N_20118,N_20986);
nor U21581 (N_21581,N_20777,N_20025);
nor U21582 (N_21582,N_20617,N_20679);
nor U21583 (N_21583,N_20563,N_20699);
nand U21584 (N_21584,N_20584,N_20637);
or U21585 (N_21585,N_20505,N_20342);
and U21586 (N_21586,N_20610,N_20158);
xnor U21587 (N_21587,N_19907,N_19565);
nor U21588 (N_21588,N_20999,N_20972);
nor U21589 (N_21589,N_20045,N_20880);
xnor U21590 (N_21590,N_20070,N_19781);
and U21591 (N_21591,N_19952,N_20018);
nand U21592 (N_21592,N_19958,N_20705);
xor U21593 (N_21593,N_20866,N_20433);
xnor U21594 (N_21594,N_20544,N_19736);
or U21595 (N_21595,N_20861,N_20159);
and U21596 (N_21596,N_20593,N_20837);
or U21597 (N_21597,N_19757,N_20881);
and U21598 (N_21598,N_20913,N_20139);
nor U21599 (N_21599,N_20600,N_20884);
nand U21600 (N_21600,N_19965,N_19933);
and U21601 (N_21601,N_20690,N_20803);
nor U21602 (N_21602,N_20996,N_19504);
or U21603 (N_21603,N_20716,N_20133);
and U21604 (N_21604,N_19843,N_20471);
or U21605 (N_21605,N_20774,N_20722);
nand U21606 (N_21606,N_19640,N_19869);
and U21607 (N_21607,N_20329,N_20486);
or U21608 (N_21608,N_20180,N_19665);
and U21609 (N_21609,N_19724,N_20585);
and U21610 (N_21610,N_20087,N_19854);
and U21611 (N_21611,N_20465,N_20795);
and U21612 (N_21612,N_20906,N_20605);
xnor U21613 (N_21613,N_20502,N_20845);
and U21614 (N_21614,N_20693,N_19953);
xnor U21615 (N_21615,N_20156,N_20819);
or U21616 (N_21616,N_20727,N_20590);
nor U21617 (N_21617,N_19789,N_19763);
xor U21618 (N_21618,N_19700,N_20085);
xor U21619 (N_21619,N_20517,N_20989);
nand U21620 (N_21620,N_19500,N_20019);
nor U21621 (N_21621,N_19984,N_20910);
or U21622 (N_21622,N_20945,N_19788);
or U21623 (N_21623,N_19548,N_20263);
xor U21624 (N_21624,N_19905,N_20982);
or U21625 (N_21625,N_20248,N_19542);
nor U21626 (N_21626,N_19560,N_20340);
and U21627 (N_21627,N_20811,N_19896);
nor U21628 (N_21628,N_19880,N_20279);
and U21629 (N_21629,N_19694,N_20707);
and U21630 (N_21630,N_19940,N_20086);
nor U21631 (N_21631,N_20239,N_19844);
or U21632 (N_21632,N_20937,N_20583);
and U21633 (N_21633,N_19826,N_19800);
xnor U21634 (N_21634,N_19827,N_20514);
and U21635 (N_21635,N_20375,N_20997);
and U21636 (N_21636,N_20588,N_19911);
xnor U21637 (N_21637,N_19780,N_19768);
or U21638 (N_21638,N_20127,N_19633);
or U21639 (N_21639,N_20492,N_19971);
or U21640 (N_21640,N_20484,N_20367);
or U21641 (N_21641,N_20423,N_20808);
xor U21642 (N_21642,N_20764,N_20561);
xor U21643 (N_21643,N_20704,N_20030);
and U21644 (N_21644,N_20189,N_20356);
xnor U21645 (N_21645,N_19524,N_19956);
nor U21646 (N_21646,N_20487,N_20011);
xor U21647 (N_21647,N_20921,N_20597);
nand U21648 (N_21648,N_20912,N_20844);
xnor U21649 (N_21649,N_20643,N_19718);
xnor U21650 (N_21650,N_20436,N_20691);
or U21651 (N_21651,N_19650,N_20474);
nor U21652 (N_21652,N_19602,N_20729);
and U21653 (N_21653,N_19607,N_20307);
nor U21654 (N_21654,N_19970,N_20155);
or U21655 (N_21655,N_20313,N_19900);
and U21656 (N_21656,N_20076,N_20162);
nand U21657 (N_21657,N_19982,N_20137);
or U21658 (N_21658,N_20886,N_19847);
nor U21659 (N_21659,N_19959,N_19719);
and U21660 (N_21660,N_20166,N_20623);
and U21661 (N_21661,N_20864,N_20765);
or U21662 (N_21662,N_20951,N_20647);
and U21663 (N_21663,N_19591,N_20769);
nand U21664 (N_21664,N_20064,N_19740);
and U21665 (N_21665,N_20347,N_19895);
nor U21666 (N_21666,N_20778,N_19756);
and U21667 (N_21667,N_19678,N_20607);
nand U21668 (N_21668,N_20173,N_19977);
nand U21669 (N_21669,N_20051,N_19817);
and U21670 (N_21670,N_19725,N_20028);
and U21671 (N_21671,N_19551,N_19767);
nand U21672 (N_21672,N_20771,N_19868);
nor U21673 (N_21673,N_20017,N_20920);
nor U21674 (N_21674,N_19619,N_20117);
nand U21675 (N_21675,N_20229,N_20503);
or U21676 (N_21676,N_19692,N_19770);
nand U21677 (N_21677,N_19711,N_20475);
and U21678 (N_21678,N_20420,N_20483);
or U21679 (N_21679,N_19875,N_20878);
or U21680 (N_21680,N_20598,N_20642);
or U21681 (N_21681,N_19759,N_20012);
xnor U21682 (N_21682,N_20244,N_20532);
and U21683 (N_21683,N_20932,N_19882);
and U21684 (N_21684,N_19883,N_20472);
nand U21685 (N_21685,N_20150,N_20618);
xor U21686 (N_21686,N_20425,N_19660);
nand U21687 (N_21687,N_20152,N_20365);
nor U21688 (N_21688,N_19976,N_20701);
and U21689 (N_21689,N_20114,N_20388);
xor U21690 (N_21690,N_20125,N_20953);
and U21691 (N_21691,N_19819,N_20868);
and U21692 (N_21692,N_20105,N_20171);
xor U21693 (N_21693,N_19507,N_19995);
and U21694 (N_21694,N_20074,N_19636);
xnor U21695 (N_21695,N_19764,N_19815);
nand U21696 (N_21696,N_20744,N_20711);
xor U21697 (N_21697,N_20428,N_20255);
and U21698 (N_21698,N_20202,N_19688);
nor U21699 (N_21699,N_20063,N_20648);
and U21700 (N_21700,N_19589,N_20231);
and U21701 (N_21701,N_20343,N_20759);
or U21702 (N_21702,N_20674,N_19687);
nor U21703 (N_21703,N_20785,N_20406);
xor U21704 (N_21704,N_20267,N_20717);
and U21705 (N_21705,N_20157,N_20036);
nor U21706 (N_21706,N_20183,N_20757);
or U21707 (N_21707,N_20188,N_20976);
nand U21708 (N_21708,N_19596,N_20115);
xnor U21709 (N_21709,N_20521,N_20784);
nand U21710 (N_21710,N_20957,N_20730);
or U21711 (N_21711,N_20501,N_20984);
nand U21712 (N_21712,N_20284,N_20111);
and U21713 (N_21713,N_19516,N_20697);
xor U21714 (N_21714,N_20956,N_19703);
nand U21715 (N_21715,N_19997,N_19638);
or U21716 (N_21716,N_20093,N_19974);
or U21717 (N_21717,N_20444,N_19651);
or U21718 (N_21718,N_20973,N_19617);
or U21719 (N_21719,N_20353,N_19773);
and U21720 (N_21720,N_20112,N_20454);
nand U21721 (N_21721,N_20066,N_20698);
or U21722 (N_21722,N_20346,N_20185);
or U21723 (N_21723,N_19654,N_20961);
and U21724 (N_21724,N_19873,N_20952);
nand U21725 (N_21725,N_20524,N_19577);
nor U21726 (N_21726,N_20092,N_20930);
and U21727 (N_21727,N_20695,N_20908);
nand U21728 (N_21728,N_20812,N_20352);
nor U21729 (N_21729,N_19750,N_20275);
or U21730 (N_21730,N_19674,N_20075);
xnor U21731 (N_21731,N_20660,N_19512);
or U21732 (N_21732,N_19659,N_20226);
nor U21733 (N_21733,N_19730,N_19604);
xor U21734 (N_21734,N_20339,N_19689);
xor U21735 (N_21735,N_20109,N_19862);
nand U21736 (N_21736,N_20380,N_20978);
xor U21737 (N_21737,N_19592,N_19603);
nor U21738 (N_21738,N_19986,N_19954);
or U21739 (N_21739,N_20446,N_19981);
xnor U21740 (N_21740,N_20658,N_20321);
xor U21741 (N_21741,N_19673,N_19612);
and U21742 (N_21742,N_20323,N_19845);
nand U21743 (N_21743,N_19867,N_20970);
and U21744 (N_21744,N_19732,N_20240);
nand U21745 (N_21745,N_19610,N_20907);
and U21746 (N_21746,N_19649,N_20067);
or U21747 (N_21747,N_19915,N_20149);
nand U21748 (N_21748,N_19555,N_19851);
and U21749 (N_21749,N_19779,N_20288);
and U21750 (N_21750,N_20013,N_20872);
or U21751 (N_21751,N_20827,N_20964);
or U21752 (N_21752,N_20217,N_20652);
xnor U21753 (N_21753,N_19845,N_20785);
nand U21754 (N_21754,N_19647,N_20097);
xor U21755 (N_21755,N_19600,N_19617);
nor U21756 (N_21756,N_19738,N_20809);
or U21757 (N_21757,N_19908,N_20393);
nor U21758 (N_21758,N_20994,N_20397);
or U21759 (N_21759,N_20850,N_20727);
and U21760 (N_21760,N_20541,N_19833);
nor U21761 (N_21761,N_20718,N_20001);
or U21762 (N_21762,N_19719,N_20387);
or U21763 (N_21763,N_19844,N_20844);
xnor U21764 (N_21764,N_20915,N_20635);
and U21765 (N_21765,N_20573,N_20316);
nand U21766 (N_21766,N_20578,N_20600);
or U21767 (N_21767,N_20942,N_19887);
xnor U21768 (N_21768,N_19758,N_19763);
nand U21769 (N_21769,N_20088,N_19670);
and U21770 (N_21770,N_20183,N_20255);
nand U21771 (N_21771,N_20512,N_20175);
nand U21772 (N_21772,N_20050,N_20223);
and U21773 (N_21773,N_19526,N_20631);
xnor U21774 (N_21774,N_19733,N_19703);
xor U21775 (N_21775,N_19647,N_20693);
and U21776 (N_21776,N_20535,N_20857);
nand U21777 (N_21777,N_20111,N_20943);
and U21778 (N_21778,N_20355,N_20437);
nand U21779 (N_21779,N_20015,N_20861);
nand U21780 (N_21780,N_20439,N_19646);
nor U21781 (N_21781,N_20022,N_20450);
nand U21782 (N_21782,N_20385,N_20210);
or U21783 (N_21783,N_20655,N_20246);
or U21784 (N_21784,N_19549,N_20417);
or U21785 (N_21785,N_20798,N_20975);
xnor U21786 (N_21786,N_20273,N_19741);
nor U21787 (N_21787,N_19877,N_20139);
or U21788 (N_21788,N_20907,N_20757);
nor U21789 (N_21789,N_20931,N_19789);
or U21790 (N_21790,N_19928,N_20272);
nand U21791 (N_21791,N_20211,N_19521);
and U21792 (N_21792,N_20268,N_19632);
nor U21793 (N_21793,N_20306,N_19940);
xor U21794 (N_21794,N_20584,N_19560);
nor U21795 (N_21795,N_19525,N_20542);
and U21796 (N_21796,N_20897,N_20040);
and U21797 (N_21797,N_19746,N_19682);
xor U21798 (N_21798,N_19981,N_20481);
nor U21799 (N_21799,N_20315,N_20965);
nor U21800 (N_21800,N_20614,N_20131);
nor U21801 (N_21801,N_20805,N_19546);
nor U21802 (N_21802,N_19505,N_19531);
and U21803 (N_21803,N_20692,N_19557);
nor U21804 (N_21804,N_20314,N_20752);
or U21805 (N_21805,N_20976,N_19651);
nor U21806 (N_21806,N_20172,N_19987);
and U21807 (N_21807,N_20252,N_20812);
xor U21808 (N_21808,N_20087,N_20085);
nor U21809 (N_21809,N_20546,N_19702);
xnor U21810 (N_21810,N_20749,N_20705);
nand U21811 (N_21811,N_20884,N_19510);
xnor U21812 (N_21812,N_20105,N_20943);
nor U21813 (N_21813,N_19864,N_19666);
nand U21814 (N_21814,N_20134,N_20202);
nand U21815 (N_21815,N_19709,N_20602);
or U21816 (N_21816,N_20070,N_20290);
and U21817 (N_21817,N_19751,N_20785);
nand U21818 (N_21818,N_20315,N_20722);
or U21819 (N_21819,N_20182,N_20549);
xnor U21820 (N_21820,N_20110,N_20418);
nand U21821 (N_21821,N_20452,N_20309);
xnor U21822 (N_21822,N_20380,N_19632);
or U21823 (N_21823,N_19615,N_20485);
or U21824 (N_21824,N_20230,N_19561);
or U21825 (N_21825,N_19989,N_20660);
nor U21826 (N_21826,N_20344,N_20277);
and U21827 (N_21827,N_20886,N_20932);
or U21828 (N_21828,N_19887,N_20118);
xnor U21829 (N_21829,N_19547,N_20922);
nor U21830 (N_21830,N_20814,N_19967);
nand U21831 (N_21831,N_20564,N_20341);
xnor U21832 (N_21832,N_19716,N_20430);
and U21833 (N_21833,N_20887,N_20056);
and U21834 (N_21834,N_19783,N_20737);
and U21835 (N_21835,N_20163,N_20252);
xnor U21836 (N_21836,N_19592,N_20506);
and U21837 (N_21837,N_20306,N_20410);
and U21838 (N_21838,N_20068,N_19742);
nor U21839 (N_21839,N_19647,N_20823);
or U21840 (N_21840,N_20984,N_20129);
nand U21841 (N_21841,N_20044,N_19701);
xnor U21842 (N_21842,N_20826,N_19875);
and U21843 (N_21843,N_20062,N_20209);
or U21844 (N_21844,N_19640,N_20463);
nor U21845 (N_21845,N_19863,N_20288);
nand U21846 (N_21846,N_19863,N_20780);
and U21847 (N_21847,N_20734,N_19905);
nor U21848 (N_21848,N_20385,N_20605);
xor U21849 (N_21849,N_20941,N_20105);
xnor U21850 (N_21850,N_19724,N_20143);
and U21851 (N_21851,N_20969,N_20452);
or U21852 (N_21852,N_20543,N_19561);
nor U21853 (N_21853,N_19713,N_20881);
and U21854 (N_21854,N_20573,N_19867);
xor U21855 (N_21855,N_20468,N_20675);
and U21856 (N_21856,N_20309,N_20963);
nand U21857 (N_21857,N_20861,N_20101);
xor U21858 (N_21858,N_20577,N_20766);
and U21859 (N_21859,N_20192,N_19691);
and U21860 (N_21860,N_20338,N_20133);
xor U21861 (N_21861,N_20721,N_20890);
nand U21862 (N_21862,N_20978,N_20927);
nand U21863 (N_21863,N_20173,N_20713);
or U21864 (N_21864,N_20631,N_19530);
nor U21865 (N_21865,N_20860,N_19508);
and U21866 (N_21866,N_19997,N_20484);
nor U21867 (N_21867,N_19506,N_20959);
nand U21868 (N_21868,N_20687,N_19525);
nor U21869 (N_21869,N_19588,N_19510);
nor U21870 (N_21870,N_19755,N_19954);
nand U21871 (N_21871,N_19536,N_20585);
nand U21872 (N_21872,N_19955,N_20178);
or U21873 (N_21873,N_20688,N_20826);
xor U21874 (N_21874,N_20204,N_20259);
nand U21875 (N_21875,N_19916,N_20008);
nand U21876 (N_21876,N_20970,N_20946);
and U21877 (N_21877,N_19968,N_20344);
or U21878 (N_21878,N_20701,N_20735);
nand U21879 (N_21879,N_19874,N_20189);
and U21880 (N_21880,N_19540,N_20773);
and U21881 (N_21881,N_20710,N_19779);
and U21882 (N_21882,N_19554,N_19619);
or U21883 (N_21883,N_20494,N_20084);
nor U21884 (N_21884,N_20161,N_20789);
nand U21885 (N_21885,N_20416,N_20229);
nor U21886 (N_21886,N_20471,N_20068);
xor U21887 (N_21887,N_19505,N_20049);
nor U21888 (N_21888,N_20223,N_20705);
xor U21889 (N_21889,N_20437,N_20744);
nor U21890 (N_21890,N_20629,N_19979);
nand U21891 (N_21891,N_19586,N_20360);
xor U21892 (N_21892,N_20579,N_20058);
xnor U21893 (N_21893,N_19819,N_20530);
nor U21894 (N_21894,N_19785,N_19929);
nor U21895 (N_21895,N_20951,N_20928);
nor U21896 (N_21896,N_20310,N_19934);
and U21897 (N_21897,N_20945,N_20922);
nand U21898 (N_21898,N_20729,N_20022);
nor U21899 (N_21899,N_20973,N_19589);
nor U21900 (N_21900,N_19564,N_20301);
and U21901 (N_21901,N_20386,N_19866);
or U21902 (N_21902,N_20192,N_19885);
or U21903 (N_21903,N_20194,N_20292);
and U21904 (N_21904,N_20857,N_20974);
and U21905 (N_21905,N_20501,N_19934);
and U21906 (N_21906,N_20301,N_20823);
nor U21907 (N_21907,N_20599,N_19918);
and U21908 (N_21908,N_19803,N_19547);
nor U21909 (N_21909,N_19977,N_20694);
xor U21910 (N_21910,N_20738,N_20334);
nor U21911 (N_21911,N_19566,N_20702);
nand U21912 (N_21912,N_19591,N_20298);
or U21913 (N_21913,N_19790,N_20391);
nor U21914 (N_21914,N_20262,N_19750);
xnor U21915 (N_21915,N_19771,N_20666);
or U21916 (N_21916,N_20556,N_19870);
nor U21917 (N_21917,N_20450,N_19733);
or U21918 (N_21918,N_19806,N_19841);
or U21919 (N_21919,N_19851,N_20324);
xor U21920 (N_21920,N_20133,N_20268);
or U21921 (N_21921,N_20679,N_20066);
nand U21922 (N_21922,N_20000,N_20466);
and U21923 (N_21923,N_20829,N_19680);
and U21924 (N_21924,N_20273,N_20538);
xor U21925 (N_21925,N_19877,N_20820);
or U21926 (N_21926,N_20599,N_19774);
and U21927 (N_21927,N_20671,N_20829);
or U21928 (N_21928,N_19789,N_20047);
nor U21929 (N_21929,N_20575,N_20879);
nor U21930 (N_21930,N_20124,N_19686);
nor U21931 (N_21931,N_20218,N_20864);
or U21932 (N_21932,N_20307,N_20093);
nor U21933 (N_21933,N_20954,N_20816);
or U21934 (N_21934,N_20930,N_19673);
and U21935 (N_21935,N_20977,N_20496);
and U21936 (N_21936,N_20779,N_20679);
xnor U21937 (N_21937,N_20622,N_20978);
or U21938 (N_21938,N_19679,N_20958);
or U21939 (N_21939,N_20383,N_20591);
or U21940 (N_21940,N_20550,N_20125);
or U21941 (N_21941,N_19676,N_20881);
xnor U21942 (N_21942,N_20918,N_20062);
nand U21943 (N_21943,N_20101,N_19818);
nor U21944 (N_21944,N_20772,N_19572);
nand U21945 (N_21945,N_20946,N_20278);
xnor U21946 (N_21946,N_20488,N_19545);
and U21947 (N_21947,N_20550,N_20814);
nor U21948 (N_21948,N_20272,N_19547);
nor U21949 (N_21949,N_20768,N_20458);
nand U21950 (N_21950,N_20946,N_20938);
nand U21951 (N_21951,N_20317,N_19774);
nand U21952 (N_21952,N_20801,N_20008);
and U21953 (N_21953,N_19601,N_20060);
nand U21954 (N_21954,N_19658,N_20375);
nor U21955 (N_21955,N_19790,N_20661);
or U21956 (N_21956,N_20090,N_20547);
nor U21957 (N_21957,N_19597,N_20755);
and U21958 (N_21958,N_19522,N_20112);
or U21959 (N_21959,N_19845,N_19743);
nor U21960 (N_21960,N_19611,N_20748);
or U21961 (N_21961,N_20753,N_20709);
and U21962 (N_21962,N_19813,N_20536);
xor U21963 (N_21963,N_19910,N_19681);
nand U21964 (N_21964,N_19631,N_19540);
or U21965 (N_21965,N_20570,N_20974);
nand U21966 (N_21966,N_20775,N_19501);
xor U21967 (N_21967,N_19523,N_20934);
and U21968 (N_21968,N_20194,N_20570);
or U21969 (N_21969,N_20931,N_20778);
xnor U21970 (N_21970,N_19684,N_20950);
nand U21971 (N_21971,N_20672,N_19596);
and U21972 (N_21972,N_20268,N_20279);
or U21973 (N_21973,N_20014,N_19575);
or U21974 (N_21974,N_20812,N_19665);
nor U21975 (N_21975,N_19725,N_20696);
nor U21976 (N_21976,N_20430,N_19982);
xor U21977 (N_21977,N_20966,N_20060);
and U21978 (N_21978,N_19523,N_20483);
nand U21979 (N_21979,N_20579,N_20177);
and U21980 (N_21980,N_19950,N_20588);
nand U21981 (N_21981,N_20268,N_19605);
nor U21982 (N_21982,N_19862,N_19641);
and U21983 (N_21983,N_20876,N_20251);
nor U21984 (N_21984,N_20766,N_20093);
xnor U21985 (N_21985,N_19643,N_20759);
nand U21986 (N_21986,N_20770,N_20631);
and U21987 (N_21987,N_20825,N_19985);
xor U21988 (N_21988,N_19814,N_20334);
xor U21989 (N_21989,N_19731,N_19908);
nand U21990 (N_21990,N_19993,N_20846);
xnor U21991 (N_21991,N_20532,N_20719);
or U21992 (N_21992,N_19618,N_20024);
or U21993 (N_21993,N_20561,N_20650);
nand U21994 (N_21994,N_20717,N_19756);
and U21995 (N_21995,N_20799,N_20442);
xnor U21996 (N_21996,N_20674,N_19692);
nor U21997 (N_21997,N_20924,N_20364);
nor U21998 (N_21998,N_19696,N_20568);
or U21999 (N_21999,N_19664,N_20234);
or U22000 (N_22000,N_19531,N_20869);
or U22001 (N_22001,N_20618,N_19814);
and U22002 (N_22002,N_19769,N_20362);
nor U22003 (N_22003,N_19920,N_20034);
nor U22004 (N_22004,N_19827,N_20518);
nor U22005 (N_22005,N_19610,N_20499);
and U22006 (N_22006,N_20509,N_19975);
nor U22007 (N_22007,N_20880,N_20981);
and U22008 (N_22008,N_19995,N_19816);
nor U22009 (N_22009,N_20928,N_19911);
nor U22010 (N_22010,N_20161,N_20906);
nand U22011 (N_22011,N_19782,N_20491);
nor U22012 (N_22012,N_20851,N_19668);
nand U22013 (N_22013,N_20883,N_20556);
xnor U22014 (N_22014,N_19967,N_20411);
nand U22015 (N_22015,N_20075,N_19905);
and U22016 (N_22016,N_20884,N_20503);
nor U22017 (N_22017,N_19512,N_20775);
nand U22018 (N_22018,N_19643,N_19975);
or U22019 (N_22019,N_20812,N_20836);
or U22020 (N_22020,N_19945,N_19780);
nand U22021 (N_22021,N_20743,N_20473);
nand U22022 (N_22022,N_20974,N_19582);
or U22023 (N_22023,N_20779,N_19936);
nor U22024 (N_22024,N_19590,N_20126);
xnor U22025 (N_22025,N_20042,N_19931);
and U22026 (N_22026,N_20871,N_20772);
nor U22027 (N_22027,N_20971,N_19697);
nor U22028 (N_22028,N_19584,N_20770);
nand U22029 (N_22029,N_19621,N_20518);
or U22030 (N_22030,N_20450,N_19924);
and U22031 (N_22031,N_19813,N_19500);
nor U22032 (N_22032,N_20525,N_20583);
or U22033 (N_22033,N_20594,N_20410);
nor U22034 (N_22034,N_20028,N_19791);
nor U22035 (N_22035,N_20589,N_20624);
or U22036 (N_22036,N_19959,N_19658);
and U22037 (N_22037,N_20816,N_20767);
xor U22038 (N_22038,N_20188,N_20934);
xor U22039 (N_22039,N_20202,N_20471);
nor U22040 (N_22040,N_20859,N_19500);
and U22041 (N_22041,N_20237,N_19863);
nor U22042 (N_22042,N_20125,N_20973);
or U22043 (N_22043,N_20655,N_19993);
or U22044 (N_22044,N_20832,N_20396);
nor U22045 (N_22045,N_19531,N_20301);
or U22046 (N_22046,N_20649,N_20981);
xor U22047 (N_22047,N_19832,N_20421);
and U22048 (N_22048,N_20374,N_19679);
or U22049 (N_22049,N_20981,N_20622);
xnor U22050 (N_22050,N_20489,N_19959);
or U22051 (N_22051,N_20185,N_20041);
nor U22052 (N_22052,N_19732,N_19538);
or U22053 (N_22053,N_20240,N_19515);
nor U22054 (N_22054,N_20443,N_20835);
and U22055 (N_22055,N_19534,N_20930);
nand U22056 (N_22056,N_19950,N_20758);
xnor U22057 (N_22057,N_20973,N_20481);
nand U22058 (N_22058,N_20548,N_20164);
and U22059 (N_22059,N_20740,N_19547);
or U22060 (N_22060,N_20282,N_19680);
nor U22061 (N_22061,N_19676,N_20492);
xor U22062 (N_22062,N_20361,N_19942);
nor U22063 (N_22063,N_20770,N_19971);
and U22064 (N_22064,N_19931,N_19919);
or U22065 (N_22065,N_20873,N_20743);
nand U22066 (N_22066,N_19767,N_19856);
xnor U22067 (N_22067,N_20139,N_19912);
xnor U22068 (N_22068,N_20159,N_20712);
nand U22069 (N_22069,N_20405,N_20768);
nand U22070 (N_22070,N_20537,N_20275);
nand U22071 (N_22071,N_20322,N_20412);
and U22072 (N_22072,N_20679,N_20294);
and U22073 (N_22073,N_20174,N_19896);
xor U22074 (N_22074,N_20468,N_20609);
and U22075 (N_22075,N_19978,N_19714);
nor U22076 (N_22076,N_19878,N_20782);
or U22077 (N_22077,N_20885,N_20877);
nand U22078 (N_22078,N_19723,N_20740);
nor U22079 (N_22079,N_20890,N_19998);
nor U22080 (N_22080,N_19581,N_20253);
or U22081 (N_22081,N_19783,N_20094);
xnor U22082 (N_22082,N_19855,N_20593);
xor U22083 (N_22083,N_19884,N_20744);
nor U22084 (N_22084,N_19841,N_20767);
xnor U22085 (N_22085,N_19744,N_19550);
nor U22086 (N_22086,N_19988,N_19843);
nor U22087 (N_22087,N_20721,N_20410);
nand U22088 (N_22088,N_19918,N_19904);
nand U22089 (N_22089,N_19832,N_19577);
or U22090 (N_22090,N_19970,N_20045);
and U22091 (N_22091,N_20317,N_19873);
nor U22092 (N_22092,N_20703,N_20335);
or U22093 (N_22093,N_20457,N_20919);
xor U22094 (N_22094,N_19840,N_20190);
nand U22095 (N_22095,N_20806,N_19977);
or U22096 (N_22096,N_20714,N_19701);
xor U22097 (N_22097,N_19969,N_20318);
xnor U22098 (N_22098,N_19613,N_19781);
nand U22099 (N_22099,N_20125,N_20200);
and U22100 (N_22100,N_20410,N_19783);
and U22101 (N_22101,N_20938,N_20094);
xnor U22102 (N_22102,N_20933,N_20930);
or U22103 (N_22103,N_20472,N_19574);
or U22104 (N_22104,N_20017,N_19867);
xor U22105 (N_22105,N_19885,N_19785);
nand U22106 (N_22106,N_19858,N_20423);
and U22107 (N_22107,N_19978,N_19727);
nor U22108 (N_22108,N_20391,N_19680);
xor U22109 (N_22109,N_20328,N_19601);
xor U22110 (N_22110,N_20011,N_20785);
or U22111 (N_22111,N_20743,N_20226);
and U22112 (N_22112,N_20390,N_19545);
nor U22113 (N_22113,N_20786,N_20891);
nor U22114 (N_22114,N_19815,N_19513);
nand U22115 (N_22115,N_20521,N_19681);
nor U22116 (N_22116,N_20152,N_20564);
nor U22117 (N_22117,N_19858,N_19552);
nor U22118 (N_22118,N_20674,N_20528);
xnor U22119 (N_22119,N_20246,N_20592);
nand U22120 (N_22120,N_20269,N_20055);
nand U22121 (N_22121,N_20935,N_20297);
xor U22122 (N_22122,N_19575,N_20628);
nand U22123 (N_22123,N_20194,N_19596);
or U22124 (N_22124,N_19578,N_20174);
nor U22125 (N_22125,N_19550,N_20037);
or U22126 (N_22126,N_19523,N_19856);
xnor U22127 (N_22127,N_19798,N_20643);
nor U22128 (N_22128,N_20604,N_20194);
and U22129 (N_22129,N_20971,N_20281);
nand U22130 (N_22130,N_20291,N_20989);
nand U22131 (N_22131,N_19666,N_20369);
xnor U22132 (N_22132,N_20642,N_20797);
xnor U22133 (N_22133,N_20252,N_19721);
or U22134 (N_22134,N_19758,N_19508);
or U22135 (N_22135,N_20352,N_20833);
nor U22136 (N_22136,N_20052,N_20159);
nand U22137 (N_22137,N_19589,N_19540);
nand U22138 (N_22138,N_19703,N_20190);
nor U22139 (N_22139,N_19800,N_20570);
or U22140 (N_22140,N_19823,N_20927);
nor U22141 (N_22141,N_20806,N_20108);
nand U22142 (N_22142,N_20353,N_20086);
xor U22143 (N_22143,N_20852,N_19529);
nand U22144 (N_22144,N_19629,N_20715);
xor U22145 (N_22145,N_19661,N_20808);
or U22146 (N_22146,N_20979,N_20660);
nand U22147 (N_22147,N_20249,N_20499);
nand U22148 (N_22148,N_20405,N_20324);
xor U22149 (N_22149,N_19710,N_20121);
or U22150 (N_22150,N_20303,N_19545);
or U22151 (N_22151,N_20417,N_20349);
nor U22152 (N_22152,N_19739,N_20807);
xor U22153 (N_22153,N_20440,N_20545);
nor U22154 (N_22154,N_19840,N_20758);
and U22155 (N_22155,N_20318,N_20192);
or U22156 (N_22156,N_20945,N_19748);
and U22157 (N_22157,N_20447,N_20769);
xnor U22158 (N_22158,N_19526,N_19764);
and U22159 (N_22159,N_20747,N_20985);
and U22160 (N_22160,N_20479,N_20978);
nor U22161 (N_22161,N_20742,N_19718);
xnor U22162 (N_22162,N_20121,N_20086);
or U22163 (N_22163,N_20517,N_20017);
nor U22164 (N_22164,N_20328,N_20534);
xor U22165 (N_22165,N_20976,N_19891);
or U22166 (N_22166,N_19642,N_20105);
or U22167 (N_22167,N_20548,N_19653);
nor U22168 (N_22168,N_20881,N_20782);
and U22169 (N_22169,N_20788,N_19699);
nand U22170 (N_22170,N_20897,N_19537);
nand U22171 (N_22171,N_20985,N_20864);
xor U22172 (N_22172,N_20337,N_19889);
xor U22173 (N_22173,N_20124,N_20291);
nand U22174 (N_22174,N_20887,N_19798);
and U22175 (N_22175,N_19659,N_19857);
xor U22176 (N_22176,N_20569,N_20124);
nand U22177 (N_22177,N_20458,N_20446);
nand U22178 (N_22178,N_19555,N_19726);
and U22179 (N_22179,N_20661,N_20840);
nand U22180 (N_22180,N_19882,N_20169);
and U22181 (N_22181,N_20648,N_20457);
nor U22182 (N_22182,N_20417,N_20713);
or U22183 (N_22183,N_20786,N_20453);
or U22184 (N_22184,N_19863,N_19634);
nor U22185 (N_22185,N_19711,N_20703);
or U22186 (N_22186,N_20261,N_19730);
xor U22187 (N_22187,N_20215,N_20880);
nor U22188 (N_22188,N_19562,N_19820);
nand U22189 (N_22189,N_19785,N_19831);
and U22190 (N_22190,N_19597,N_19877);
and U22191 (N_22191,N_20546,N_20626);
xnor U22192 (N_22192,N_19610,N_19818);
nor U22193 (N_22193,N_20742,N_20555);
nor U22194 (N_22194,N_20200,N_20660);
xor U22195 (N_22195,N_20556,N_20512);
and U22196 (N_22196,N_19686,N_20511);
nor U22197 (N_22197,N_19501,N_20339);
nand U22198 (N_22198,N_19690,N_19662);
or U22199 (N_22199,N_20953,N_20203);
nand U22200 (N_22200,N_20235,N_19703);
nand U22201 (N_22201,N_20111,N_19778);
or U22202 (N_22202,N_20910,N_20981);
and U22203 (N_22203,N_20478,N_20870);
or U22204 (N_22204,N_20699,N_19897);
and U22205 (N_22205,N_19865,N_20439);
xnor U22206 (N_22206,N_20018,N_20174);
nor U22207 (N_22207,N_20995,N_19692);
xnor U22208 (N_22208,N_20214,N_20476);
or U22209 (N_22209,N_20139,N_20619);
xnor U22210 (N_22210,N_20848,N_20602);
nand U22211 (N_22211,N_19786,N_19626);
or U22212 (N_22212,N_20673,N_19959);
or U22213 (N_22213,N_19959,N_20875);
xnor U22214 (N_22214,N_19758,N_19547);
nand U22215 (N_22215,N_20433,N_19963);
xor U22216 (N_22216,N_19584,N_20308);
or U22217 (N_22217,N_19639,N_19574);
or U22218 (N_22218,N_20281,N_20501);
nor U22219 (N_22219,N_20121,N_19601);
or U22220 (N_22220,N_19844,N_20729);
nand U22221 (N_22221,N_19692,N_19666);
xnor U22222 (N_22222,N_19599,N_20826);
and U22223 (N_22223,N_20078,N_19629);
or U22224 (N_22224,N_20930,N_19979);
or U22225 (N_22225,N_20787,N_20472);
xnor U22226 (N_22226,N_20270,N_20134);
xor U22227 (N_22227,N_20391,N_20920);
or U22228 (N_22228,N_19576,N_19587);
and U22229 (N_22229,N_19536,N_20286);
nand U22230 (N_22230,N_20930,N_20245);
nor U22231 (N_22231,N_19917,N_19596);
nand U22232 (N_22232,N_19860,N_19512);
xnor U22233 (N_22233,N_19771,N_20703);
and U22234 (N_22234,N_20832,N_19997);
xnor U22235 (N_22235,N_19543,N_20096);
nor U22236 (N_22236,N_20831,N_19687);
nand U22237 (N_22237,N_19652,N_19568);
and U22238 (N_22238,N_20979,N_19912);
nor U22239 (N_22239,N_20807,N_19619);
xor U22240 (N_22240,N_20851,N_20679);
or U22241 (N_22241,N_20120,N_20175);
xor U22242 (N_22242,N_20269,N_20959);
nand U22243 (N_22243,N_19717,N_20104);
or U22244 (N_22244,N_20478,N_19821);
or U22245 (N_22245,N_20332,N_20542);
and U22246 (N_22246,N_20075,N_20202);
and U22247 (N_22247,N_19799,N_20920);
or U22248 (N_22248,N_20387,N_19869);
xor U22249 (N_22249,N_20022,N_19541);
xnor U22250 (N_22250,N_19948,N_19798);
nor U22251 (N_22251,N_20643,N_20553);
nand U22252 (N_22252,N_20774,N_20561);
and U22253 (N_22253,N_20302,N_20013);
nand U22254 (N_22254,N_19536,N_20584);
and U22255 (N_22255,N_19582,N_20240);
nand U22256 (N_22256,N_19966,N_19901);
and U22257 (N_22257,N_19625,N_20777);
nor U22258 (N_22258,N_20180,N_20281);
nor U22259 (N_22259,N_19697,N_20103);
or U22260 (N_22260,N_20651,N_20395);
xor U22261 (N_22261,N_20024,N_19588);
nand U22262 (N_22262,N_20357,N_20468);
xor U22263 (N_22263,N_20426,N_20247);
or U22264 (N_22264,N_20741,N_20888);
or U22265 (N_22265,N_20574,N_20893);
and U22266 (N_22266,N_19911,N_20010);
and U22267 (N_22267,N_19682,N_19724);
nor U22268 (N_22268,N_20862,N_19813);
nand U22269 (N_22269,N_20426,N_20145);
nor U22270 (N_22270,N_20522,N_19963);
nor U22271 (N_22271,N_19723,N_20739);
and U22272 (N_22272,N_20269,N_19826);
and U22273 (N_22273,N_19667,N_20756);
xor U22274 (N_22274,N_19836,N_20992);
xor U22275 (N_22275,N_20411,N_19634);
xor U22276 (N_22276,N_19551,N_19769);
xor U22277 (N_22277,N_20266,N_20998);
and U22278 (N_22278,N_20631,N_20471);
nor U22279 (N_22279,N_19663,N_20121);
nor U22280 (N_22280,N_19913,N_20713);
nand U22281 (N_22281,N_19577,N_20473);
nor U22282 (N_22282,N_19547,N_19822);
nand U22283 (N_22283,N_20486,N_20254);
xnor U22284 (N_22284,N_20145,N_20622);
nor U22285 (N_22285,N_20007,N_20765);
and U22286 (N_22286,N_20623,N_19730);
nand U22287 (N_22287,N_20936,N_19955);
nand U22288 (N_22288,N_19919,N_20935);
and U22289 (N_22289,N_20403,N_19843);
nand U22290 (N_22290,N_20936,N_19992);
and U22291 (N_22291,N_20379,N_20113);
nand U22292 (N_22292,N_20729,N_20318);
xnor U22293 (N_22293,N_20165,N_20353);
xnor U22294 (N_22294,N_19502,N_20262);
or U22295 (N_22295,N_19643,N_20789);
and U22296 (N_22296,N_19850,N_20299);
xor U22297 (N_22297,N_20342,N_20824);
xor U22298 (N_22298,N_20656,N_20159);
nand U22299 (N_22299,N_19887,N_20241);
xnor U22300 (N_22300,N_20785,N_19636);
nor U22301 (N_22301,N_19775,N_19954);
xnor U22302 (N_22302,N_20710,N_19814);
nand U22303 (N_22303,N_20056,N_20103);
nand U22304 (N_22304,N_20946,N_19853);
nor U22305 (N_22305,N_20947,N_20830);
or U22306 (N_22306,N_20835,N_20519);
and U22307 (N_22307,N_19917,N_19522);
or U22308 (N_22308,N_20242,N_20689);
and U22309 (N_22309,N_20691,N_20004);
nor U22310 (N_22310,N_19726,N_20087);
and U22311 (N_22311,N_19980,N_19616);
or U22312 (N_22312,N_19558,N_19634);
xnor U22313 (N_22313,N_19884,N_19656);
xor U22314 (N_22314,N_20149,N_19893);
nand U22315 (N_22315,N_20402,N_20030);
xor U22316 (N_22316,N_20100,N_20200);
nand U22317 (N_22317,N_19608,N_20607);
and U22318 (N_22318,N_20640,N_20461);
nand U22319 (N_22319,N_20025,N_20081);
nand U22320 (N_22320,N_20068,N_20993);
nor U22321 (N_22321,N_19613,N_20956);
nand U22322 (N_22322,N_19753,N_19723);
or U22323 (N_22323,N_20540,N_20259);
xor U22324 (N_22324,N_20055,N_20890);
xor U22325 (N_22325,N_20956,N_20078);
xor U22326 (N_22326,N_20206,N_19891);
nor U22327 (N_22327,N_20968,N_19629);
xnor U22328 (N_22328,N_20651,N_20547);
nand U22329 (N_22329,N_20646,N_20481);
and U22330 (N_22330,N_20698,N_19715);
and U22331 (N_22331,N_20760,N_20880);
xnor U22332 (N_22332,N_20246,N_19615);
nor U22333 (N_22333,N_20611,N_20840);
nor U22334 (N_22334,N_20962,N_20269);
xor U22335 (N_22335,N_20325,N_20613);
or U22336 (N_22336,N_20305,N_19803);
or U22337 (N_22337,N_20462,N_19577);
xor U22338 (N_22338,N_20898,N_20014);
or U22339 (N_22339,N_19579,N_19511);
nand U22340 (N_22340,N_20085,N_19822);
and U22341 (N_22341,N_20443,N_20103);
or U22342 (N_22342,N_20640,N_19554);
or U22343 (N_22343,N_20634,N_20023);
nand U22344 (N_22344,N_19581,N_19878);
and U22345 (N_22345,N_20140,N_19513);
nor U22346 (N_22346,N_19613,N_19643);
and U22347 (N_22347,N_19955,N_19545);
xor U22348 (N_22348,N_20535,N_20407);
or U22349 (N_22349,N_20631,N_19510);
or U22350 (N_22350,N_20203,N_20803);
nand U22351 (N_22351,N_20889,N_20843);
and U22352 (N_22352,N_20912,N_20858);
nor U22353 (N_22353,N_20194,N_19717);
nand U22354 (N_22354,N_20876,N_19993);
nand U22355 (N_22355,N_20576,N_20305);
and U22356 (N_22356,N_20505,N_20533);
xor U22357 (N_22357,N_19825,N_20715);
and U22358 (N_22358,N_20054,N_19846);
nor U22359 (N_22359,N_19515,N_20349);
nand U22360 (N_22360,N_19886,N_20481);
nand U22361 (N_22361,N_20587,N_20628);
or U22362 (N_22362,N_20449,N_19894);
nand U22363 (N_22363,N_19965,N_20749);
and U22364 (N_22364,N_20089,N_19563);
and U22365 (N_22365,N_20398,N_19823);
xor U22366 (N_22366,N_20380,N_19776);
nand U22367 (N_22367,N_20115,N_20683);
xnor U22368 (N_22368,N_20970,N_20983);
nor U22369 (N_22369,N_20304,N_20761);
or U22370 (N_22370,N_20531,N_20614);
xor U22371 (N_22371,N_20710,N_20259);
xnor U22372 (N_22372,N_19515,N_19533);
xor U22373 (N_22373,N_19565,N_19658);
nor U22374 (N_22374,N_19507,N_20303);
and U22375 (N_22375,N_19501,N_19592);
or U22376 (N_22376,N_20402,N_19937);
and U22377 (N_22377,N_20718,N_20810);
or U22378 (N_22378,N_20754,N_19681);
and U22379 (N_22379,N_20783,N_20606);
nand U22380 (N_22380,N_19709,N_20032);
or U22381 (N_22381,N_19897,N_19513);
xnor U22382 (N_22382,N_20435,N_19563);
or U22383 (N_22383,N_20415,N_19726);
nand U22384 (N_22384,N_20458,N_20375);
nand U22385 (N_22385,N_20123,N_19787);
and U22386 (N_22386,N_19924,N_20592);
or U22387 (N_22387,N_19823,N_20092);
xor U22388 (N_22388,N_19819,N_20512);
nor U22389 (N_22389,N_19988,N_20541);
nor U22390 (N_22390,N_20151,N_19733);
xor U22391 (N_22391,N_19779,N_20984);
nand U22392 (N_22392,N_19801,N_20177);
nor U22393 (N_22393,N_19990,N_19668);
xnor U22394 (N_22394,N_20964,N_20684);
nand U22395 (N_22395,N_19659,N_20154);
or U22396 (N_22396,N_20429,N_20821);
or U22397 (N_22397,N_19531,N_19598);
nand U22398 (N_22398,N_20380,N_20824);
nor U22399 (N_22399,N_20817,N_20499);
or U22400 (N_22400,N_20485,N_20834);
xnor U22401 (N_22401,N_19540,N_20793);
nor U22402 (N_22402,N_20321,N_19902);
xor U22403 (N_22403,N_20190,N_20063);
or U22404 (N_22404,N_20800,N_20454);
and U22405 (N_22405,N_19879,N_20711);
nor U22406 (N_22406,N_20709,N_20982);
nor U22407 (N_22407,N_19630,N_19998);
or U22408 (N_22408,N_20407,N_20121);
nor U22409 (N_22409,N_20287,N_20692);
xnor U22410 (N_22410,N_20726,N_20958);
and U22411 (N_22411,N_19982,N_19838);
and U22412 (N_22412,N_19869,N_20286);
nor U22413 (N_22413,N_20490,N_19528);
and U22414 (N_22414,N_20003,N_19960);
xnor U22415 (N_22415,N_19865,N_20754);
nand U22416 (N_22416,N_19598,N_19907);
or U22417 (N_22417,N_20017,N_20487);
and U22418 (N_22418,N_20572,N_20019);
or U22419 (N_22419,N_20553,N_19889);
nor U22420 (N_22420,N_20290,N_20125);
nand U22421 (N_22421,N_19574,N_19775);
xnor U22422 (N_22422,N_19780,N_20928);
xnor U22423 (N_22423,N_19653,N_20052);
or U22424 (N_22424,N_19827,N_19882);
xor U22425 (N_22425,N_20978,N_19925);
nand U22426 (N_22426,N_20331,N_20211);
and U22427 (N_22427,N_20676,N_20509);
nand U22428 (N_22428,N_19886,N_19716);
nor U22429 (N_22429,N_19920,N_20271);
and U22430 (N_22430,N_20192,N_20678);
xor U22431 (N_22431,N_20735,N_20448);
xnor U22432 (N_22432,N_19631,N_19666);
xor U22433 (N_22433,N_20322,N_20098);
xnor U22434 (N_22434,N_20501,N_20658);
xor U22435 (N_22435,N_19517,N_19885);
xnor U22436 (N_22436,N_20060,N_20408);
and U22437 (N_22437,N_19571,N_20371);
nand U22438 (N_22438,N_19547,N_20007);
nand U22439 (N_22439,N_20896,N_20745);
and U22440 (N_22440,N_20966,N_20298);
or U22441 (N_22441,N_20564,N_19734);
and U22442 (N_22442,N_20119,N_20768);
and U22443 (N_22443,N_20213,N_20275);
xnor U22444 (N_22444,N_20272,N_19689);
or U22445 (N_22445,N_19823,N_20279);
nand U22446 (N_22446,N_20859,N_20770);
nand U22447 (N_22447,N_20961,N_19747);
or U22448 (N_22448,N_20946,N_19516);
xor U22449 (N_22449,N_20841,N_19846);
and U22450 (N_22450,N_20927,N_20464);
xnor U22451 (N_22451,N_20218,N_19500);
and U22452 (N_22452,N_20932,N_19836);
xor U22453 (N_22453,N_19633,N_20872);
nor U22454 (N_22454,N_20527,N_19922);
xor U22455 (N_22455,N_19827,N_20055);
or U22456 (N_22456,N_20206,N_20429);
or U22457 (N_22457,N_20094,N_20414);
or U22458 (N_22458,N_20737,N_19974);
xnor U22459 (N_22459,N_20493,N_20360);
nand U22460 (N_22460,N_20631,N_20180);
nor U22461 (N_22461,N_20672,N_19894);
nand U22462 (N_22462,N_19910,N_20647);
or U22463 (N_22463,N_19828,N_20069);
and U22464 (N_22464,N_20613,N_20588);
nor U22465 (N_22465,N_20066,N_19882);
nand U22466 (N_22466,N_20160,N_19738);
xnor U22467 (N_22467,N_19775,N_19704);
and U22468 (N_22468,N_20045,N_19569);
and U22469 (N_22469,N_19661,N_19837);
and U22470 (N_22470,N_20187,N_20332);
xnor U22471 (N_22471,N_19630,N_20020);
nor U22472 (N_22472,N_20022,N_20167);
nor U22473 (N_22473,N_20501,N_19558);
xnor U22474 (N_22474,N_19877,N_20255);
nor U22475 (N_22475,N_20088,N_19789);
and U22476 (N_22476,N_20604,N_20524);
nor U22477 (N_22477,N_20226,N_20516);
nand U22478 (N_22478,N_20664,N_19882);
nand U22479 (N_22479,N_20499,N_19536);
nand U22480 (N_22480,N_20686,N_20747);
nor U22481 (N_22481,N_19504,N_20533);
and U22482 (N_22482,N_20134,N_20678);
and U22483 (N_22483,N_20590,N_20007);
or U22484 (N_22484,N_19679,N_19915);
nand U22485 (N_22485,N_20708,N_20910);
nor U22486 (N_22486,N_20541,N_20915);
nand U22487 (N_22487,N_20556,N_19750);
nor U22488 (N_22488,N_20668,N_20310);
nand U22489 (N_22489,N_20297,N_20449);
or U22490 (N_22490,N_20401,N_20478);
nand U22491 (N_22491,N_20458,N_19545);
nor U22492 (N_22492,N_19740,N_19530);
nor U22493 (N_22493,N_19742,N_19818);
and U22494 (N_22494,N_20339,N_19914);
or U22495 (N_22495,N_20794,N_20696);
nand U22496 (N_22496,N_20226,N_20890);
xnor U22497 (N_22497,N_19933,N_20240);
or U22498 (N_22498,N_20490,N_19521);
nand U22499 (N_22499,N_19945,N_20443);
and U22500 (N_22500,N_22220,N_22370);
xor U22501 (N_22501,N_21718,N_22210);
or U22502 (N_22502,N_21310,N_21287);
or U22503 (N_22503,N_22386,N_21578);
and U22504 (N_22504,N_21436,N_21676);
or U22505 (N_22505,N_21738,N_22408);
nor U22506 (N_22506,N_22372,N_21284);
nand U22507 (N_22507,N_22481,N_21566);
xnor U22508 (N_22508,N_21082,N_22230);
or U22509 (N_22509,N_22318,N_22018);
nand U22510 (N_22510,N_22187,N_22056);
nand U22511 (N_22511,N_21120,N_21489);
xor U22512 (N_22512,N_22200,N_22222);
nand U22513 (N_22513,N_21755,N_22265);
nand U22514 (N_22514,N_22027,N_21129);
and U22515 (N_22515,N_21325,N_21753);
and U22516 (N_22516,N_21801,N_21869);
and U22517 (N_22517,N_22344,N_21092);
and U22518 (N_22518,N_21172,N_21587);
nor U22519 (N_22519,N_22353,N_21192);
or U22520 (N_22520,N_21953,N_22239);
or U22521 (N_22521,N_21593,N_22463);
xnor U22522 (N_22522,N_22270,N_21889);
nand U22523 (N_22523,N_21087,N_21634);
nor U22524 (N_22524,N_21452,N_21317);
and U22525 (N_22525,N_21212,N_21659);
or U22526 (N_22526,N_22392,N_22449);
or U22527 (N_22527,N_21205,N_22469);
or U22528 (N_22528,N_22020,N_21012);
or U22529 (N_22529,N_21565,N_21077);
nand U22530 (N_22530,N_21181,N_21496);
nor U22531 (N_22531,N_21562,N_21846);
nand U22532 (N_22532,N_21538,N_21184);
xor U22533 (N_22533,N_21219,N_22458);
nand U22534 (N_22534,N_21180,N_21653);
and U22535 (N_22535,N_22231,N_21467);
or U22536 (N_22536,N_21732,N_21655);
nand U22537 (N_22537,N_21335,N_21878);
xnor U22538 (N_22538,N_21369,N_21473);
nor U22539 (N_22539,N_21556,N_21690);
and U22540 (N_22540,N_21057,N_21855);
nor U22541 (N_22541,N_21966,N_21618);
nor U22542 (N_22542,N_21961,N_22323);
xor U22543 (N_22543,N_22155,N_22066);
nand U22544 (N_22544,N_22117,N_21071);
xnor U22545 (N_22545,N_21045,N_21863);
nand U22546 (N_22546,N_22436,N_21886);
nand U22547 (N_22547,N_21599,N_22075);
nand U22548 (N_22548,N_21629,N_21602);
xnor U22549 (N_22549,N_22476,N_21227);
nand U22550 (N_22550,N_22193,N_21487);
or U22551 (N_22551,N_21145,N_21568);
nand U22552 (N_22552,N_21713,N_22226);
or U22553 (N_22553,N_22329,N_22494);
or U22554 (N_22554,N_22065,N_21802);
xor U22555 (N_22555,N_21925,N_21897);
xnor U22556 (N_22556,N_21028,N_22433);
nand U22557 (N_22557,N_21497,N_22090);
nor U22558 (N_22558,N_21196,N_21788);
nand U22559 (N_22559,N_22198,N_22424);
and U22560 (N_22560,N_21503,N_22406);
xor U22561 (N_22561,N_22173,N_22477);
nor U22562 (N_22562,N_21262,N_21164);
nor U22563 (N_22563,N_22307,N_22276);
and U22564 (N_22564,N_21030,N_21934);
xor U22565 (N_22565,N_21074,N_22109);
and U22566 (N_22566,N_21331,N_21620);
nand U22567 (N_22567,N_21548,N_22261);
xnor U22568 (N_22568,N_21533,N_21281);
or U22569 (N_22569,N_21792,N_21063);
nand U22570 (N_22570,N_22060,N_21509);
nor U22571 (N_22571,N_21600,N_22175);
and U22572 (N_22572,N_21131,N_22237);
xor U22573 (N_22573,N_22167,N_22029);
or U22574 (N_22574,N_21787,N_21817);
nand U22575 (N_22575,N_21661,N_21151);
or U22576 (N_22576,N_21737,N_21011);
nand U22577 (N_22577,N_22396,N_21770);
nand U22578 (N_22578,N_21988,N_22205);
nand U22579 (N_22579,N_21607,N_21336);
nand U22580 (N_22580,N_21564,N_21025);
or U22581 (N_22581,N_22233,N_22467);
or U22582 (N_22582,N_22023,N_22267);
nand U22583 (N_22583,N_21899,N_21757);
or U22584 (N_22584,N_22331,N_22111);
nor U22585 (N_22585,N_22213,N_21141);
xnor U22586 (N_22586,N_21308,N_22209);
xnor U22587 (N_22587,N_21266,N_21225);
xor U22588 (N_22588,N_22119,N_22382);
nand U22589 (N_22589,N_22201,N_21734);
nor U22590 (N_22590,N_21039,N_21637);
and U22591 (N_22591,N_22168,N_22170);
and U22592 (N_22592,N_22364,N_22328);
xor U22593 (N_22593,N_21384,N_22037);
and U22594 (N_22594,N_21032,N_21278);
xnor U22595 (N_22595,N_21409,N_21823);
nor U22596 (N_22596,N_21407,N_21230);
and U22597 (N_22597,N_22212,N_21260);
and U22598 (N_22598,N_21632,N_21270);
or U22599 (N_22599,N_22019,N_21550);
nor U22600 (N_22600,N_22339,N_21847);
or U22601 (N_22601,N_21860,N_22369);
nor U22602 (N_22602,N_21264,N_22437);
nor U22603 (N_22603,N_21622,N_21474);
and U22604 (N_22604,N_22289,N_22256);
nand U22605 (N_22605,N_21315,N_21983);
and U22606 (N_22606,N_21505,N_21457);
nor U22607 (N_22607,N_21932,N_22482);
nand U22608 (N_22608,N_21610,N_21882);
or U22609 (N_22609,N_21162,N_21495);
nor U22610 (N_22610,N_21206,N_22462);
nor U22611 (N_22611,N_22346,N_21640);
nand U22612 (N_22612,N_22208,N_22082);
nor U22613 (N_22613,N_21088,N_21099);
nor U22614 (N_22614,N_21643,N_21534);
and U22615 (N_22615,N_21084,N_21042);
or U22616 (N_22616,N_22043,N_22079);
and U22617 (N_22617,N_21651,N_21746);
nor U22618 (N_22618,N_21105,N_21909);
or U22619 (N_22619,N_22286,N_21806);
and U22620 (N_22620,N_21774,N_21217);
xor U22621 (N_22621,N_22185,N_21322);
or U22622 (N_22622,N_21856,N_21586);
and U22623 (N_22623,N_21916,N_21330);
or U22624 (N_22624,N_21437,N_22073);
and U22625 (N_22625,N_21765,N_21530);
or U22626 (N_22626,N_22127,N_21572);
or U22627 (N_22627,N_21874,N_21938);
or U22628 (N_22628,N_22247,N_21689);
nor U22629 (N_22629,N_21234,N_21933);
xor U22630 (N_22630,N_21694,N_21019);
nor U22631 (N_22631,N_21880,N_21604);
or U22632 (N_22632,N_22045,N_22496);
xnor U22633 (N_22633,N_22016,N_21744);
or U22634 (N_22634,N_21958,N_21388);
xnor U22635 (N_22635,N_22076,N_21175);
nor U22636 (N_22636,N_21229,N_21290);
nand U22637 (N_22637,N_21853,N_22257);
nand U22638 (N_22638,N_22225,N_21213);
xnor U22639 (N_22639,N_21567,N_21829);
xnor U22640 (N_22640,N_21244,N_21132);
xnor U22641 (N_22641,N_21392,N_22316);
xor U22642 (N_22642,N_21512,N_22394);
nor U22643 (N_22643,N_21571,N_22250);
xnor U22644 (N_22644,N_21100,N_22093);
and U22645 (N_22645,N_22492,N_21908);
xnor U22646 (N_22646,N_22218,N_22010);
xnor U22647 (N_22647,N_21528,N_21173);
nor U22648 (N_22648,N_22303,N_21349);
nor U22649 (N_22649,N_22030,N_21545);
nor U22650 (N_22650,N_21472,N_21768);
or U22651 (N_22651,N_22260,N_22374);
nor U22652 (N_22652,N_21194,N_21759);
or U22653 (N_22653,N_21096,N_21666);
and U22654 (N_22654,N_21361,N_21047);
nand U22655 (N_22655,N_21769,N_21685);
and U22656 (N_22656,N_22480,N_22135);
nand U22657 (N_22657,N_22129,N_21803);
xnor U22658 (N_22658,N_21379,N_21884);
and U22659 (N_22659,N_21269,N_21558);
nor U22660 (N_22660,N_21805,N_22332);
and U22661 (N_22661,N_21647,N_22269);
nand U22662 (N_22662,N_21560,N_22409);
nor U22663 (N_22663,N_22086,N_22297);
or U22664 (N_22664,N_21553,N_21780);
xor U22665 (N_22665,N_21646,N_22262);
or U22666 (N_22666,N_21917,N_22485);
or U22667 (N_22667,N_21292,N_21453);
or U22668 (N_22668,N_21671,N_22348);
nor U22669 (N_22669,N_22004,N_21594);
or U22670 (N_22670,N_22244,N_21059);
and U22671 (N_22671,N_21037,N_22191);
xnor U22672 (N_22672,N_21477,N_22491);
or U22673 (N_22673,N_22371,N_21169);
xnor U22674 (N_22674,N_22089,N_21395);
nor U22675 (N_22675,N_21420,N_22055);
nor U22676 (N_22676,N_21050,N_22301);
nor U22677 (N_22677,N_21464,N_21060);
xnor U22678 (N_22678,N_21771,N_22162);
and U22679 (N_22679,N_21524,N_21081);
nor U22680 (N_22680,N_21009,N_22497);
nand U22681 (N_22681,N_21963,N_21842);
nor U22682 (N_22682,N_22121,N_21750);
and U22683 (N_22683,N_22039,N_21910);
nor U22684 (N_22684,N_22139,N_22042);
or U22685 (N_22685,N_21589,N_22499);
or U22686 (N_22686,N_21258,N_21176);
nand U22687 (N_22687,N_21525,N_21121);
xnor U22688 (N_22688,N_21809,N_22221);
nor U22689 (N_22689,N_22182,N_22280);
xor U22690 (N_22690,N_21228,N_21949);
or U22691 (N_22691,N_22118,N_21535);
nor U22692 (N_22692,N_21752,N_21764);
nand U22693 (N_22693,N_21135,N_21575);
or U22694 (N_22694,N_21118,N_22398);
nor U22695 (N_22695,N_22115,N_21365);
and U22696 (N_22696,N_21945,N_21285);
nor U22697 (N_22697,N_22390,N_21998);
and U22698 (N_22698,N_21796,N_21102);
nand U22699 (N_22699,N_22425,N_21968);
and U22700 (N_22700,N_22405,N_22421);
or U22701 (N_22701,N_21631,N_21171);
xnor U22702 (N_22702,N_21499,N_22298);
nand U22703 (N_22703,N_21872,N_21203);
xnor U22704 (N_22704,N_22308,N_21888);
nor U22705 (N_22705,N_22204,N_21990);
nand U22706 (N_22706,N_21763,N_21611);
or U22707 (N_22707,N_22181,N_21098);
nor U22708 (N_22708,N_22271,N_21893);
nor U22709 (N_22709,N_21581,N_21526);
nand U22710 (N_22710,N_21928,N_21914);
xnor U22711 (N_22711,N_22157,N_22051);
or U22712 (N_22712,N_21065,N_21166);
nor U22713 (N_22713,N_22203,N_21895);
xor U22714 (N_22714,N_22116,N_21023);
nand U22715 (N_22715,N_21896,N_22196);
nor U22716 (N_22716,N_21149,N_21106);
xnor U22717 (N_22717,N_21426,N_21912);
or U22718 (N_22718,N_21049,N_21439);
and U22719 (N_22719,N_21351,N_21391);
nor U22720 (N_22720,N_21017,N_22363);
and U22721 (N_22721,N_21339,N_21320);
nor U22722 (N_22722,N_21044,N_21861);
xor U22723 (N_22723,N_21577,N_21724);
nor U22724 (N_22724,N_21306,N_21731);
or U22725 (N_22725,N_21279,N_21356);
nor U22726 (N_22726,N_21137,N_21662);
nor U22727 (N_22727,N_21479,N_21703);
nor U22728 (N_22728,N_21794,N_21202);
or U22729 (N_22729,N_21508,N_22466);
and U22730 (N_22730,N_22327,N_21546);
or U22731 (N_22731,N_21109,N_22341);
and U22732 (N_22732,N_21348,N_21877);
xor U22733 (N_22733,N_21642,N_21778);
xnor U22734 (N_22734,N_21143,N_21160);
nor U22735 (N_22735,N_21779,N_21201);
nor U22736 (N_22736,N_21412,N_21127);
xor U22737 (N_22737,N_21969,N_21943);
or U22738 (N_22738,N_21022,N_21165);
and U22739 (N_22739,N_22351,N_22317);
nand U22740 (N_22740,N_21040,N_21862);
and U22741 (N_22741,N_21729,N_21529);
or U22742 (N_22742,N_21431,N_21274);
xnor U22743 (N_22743,N_22160,N_22350);
xor U22744 (N_22744,N_21403,N_21454);
nor U22745 (N_22745,N_21584,N_22136);
nand U22746 (N_22746,N_21507,N_21490);
nand U22747 (N_22747,N_22024,N_21235);
or U22748 (N_22748,N_22154,N_21960);
or U22749 (N_22749,N_22202,N_21232);
or U22750 (N_22750,N_22373,N_21543);
or U22751 (N_22751,N_21657,N_21520);
nor U22752 (N_22752,N_21785,N_21691);
and U22753 (N_22753,N_21328,N_21375);
nand U22754 (N_22754,N_21965,N_21277);
or U22755 (N_22755,N_21980,N_21563);
xnor U22756 (N_22756,N_22413,N_22284);
or U22757 (N_22757,N_21876,N_22197);
xnor U22758 (N_22758,N_21302,N_21210);
xnor U22759 (N_22759,N_22368,N_21043);
nand U22760 (N_22760,N_21372,N_21513);
xor U22761 (N_22761,N_21033,N_22358);
xnor U22762 (N_22762,N_21170,N_21838);
and U22763 (N_22763,N_22444,N_21273);
xnor U22764 (N_22764,N_22391,N_21001);
or U22765 (N_22765,N_22147,N_22465);
or U22766 (N_22766,N_21163,N_21830);
xnor U22767 (N_22767,N_21465,N_21821);
and U22768 (N_22768,N_22451,N_22091);
xor U22769 (N_22769,N_21854,N_22385);
xor U22770 (N_22770,N_21839,N_21826);
nor U22771 (N_22771,N_21214,N_22174);
and U22772 (N_22772,N_22335,N_21153);
nand U22773 (N_22773,N_21382,N_21185);
and U22774 (N_22774,N_22132,N_21784);
nor U22775 (N_22775,N_21720,N_21374);
and U22776 (N_22776,N_21051,N_21034);
and U22777 (N_22777,N_22285,N_22140);
or U22778 (N_22778,N_22375,N_21946);
and U22779 (N_22779,N_21075,N_21745);
xor U22780 (N_22780,N_21405,N_21378);
or U22781 (N_22781,N_21549,N_21195);
or U22782 (N_22782,N_21812,N_21608);
xor U22783 (N_22783,N_21068,N_21673);
nor U22784 (N_22784,N_21000,N_21038);
nand U22785 (N_22785,N_22067,N_21362);
and U22786 (N_22786,N_21404,N_21677);
nor U22787 (N_22787,N_21427,N_21698);
and U22788 (N_22788,N_21641,N_21444);
or U22789 (N_22789,N_21865,N_21159);
or U22790 (N_22790,N_21303,N_21580);
nor U22791 (N_22791,N_21819,N_21644);
nand U22792 (N_22792,N_22028,N_21761);
nand U22793 (N_22793,N_21289,N_21255);
or U22794 (N_22794,N_22435,N_22282);
xor U22795 (N_22795,N_21712,N_21951);
xnor U22796 (N_22796,N_22044,N_21389);
nor U22797 (N_22797,N_21240,N_21552);
nand U22798 (N_22798,N_21332,N_21236);
xor U22799 (N_22799,N_21055,N_21337);
and U22800 (N_22800,N_21523,N_22235);
nand U22801 (N_22801,N_21625,N_21613);
or U22802 (N_22802,N_21144,N_21539);
or U22803 (N_22803,N_22041,N_21590);
or U22804 (N_22804,N_21340,N_21595);
or U22805 (N_22805,N_21736,N_21476);
xor U22806 (N_22806,N_21238,N_22080);
or U22807 (N_22807,N_21808,N_21841);
or U22808 (N_22808,N_22078,N_22493);
or U22809 (N_22809,N_21247,N_21748);
nand U22810 (N_22810,N_22326,N_21293);
nor U22811 (N_22811,N_21198,N_21518);
nand U22812 (N_22812,N_21996,N_22410);
nor U22813 (N_22813,N_22443,N_22001);
nor U22814 (N_22814,N_21422,N_21664);
and U22815 (N_22815,N_21492,N_21015);
or U22816 (N_22816,N_22272,N_21130);
and U22817 (N_22817,N_21681,N_22402);
xor U22818 (N_22818,N_21972,N_21605);
and U22819 (N_22819,N_21758,N_21128);
and U22820 (N_22820,N_22486,N_22074);
xnor U22821 (N_22821,N_21443,N_21502);
or U22822 (N_22822,N_21663,N_21253);
and U22823 (N_22823,N_21221,N_21209);
or U22824 (N_22824,N_22330,N_21716);
and U22825 (N_22825,N_21923,N_22143);
nand U22826 (N_22826,N_22022,N_21386);
xor U22827 (N_22827,N_21101,N_21211);
or U22828 (N_22828,N_21463,N_22014);
and U22829 (N_22829,N_22487,N_21656);
or U22830 (N_22830,N_21814,N_21527);
nand U22831 (N_22831,N_22114,N_22274);
nor U22832 (N_22832,N_22321,N_21466);
and U22833 (N_22833,N_22283,N_21927);
or U22834 (N_22834,N_21275,N_21762);
nor U22835 (N_22835,N_21344,N_21596);
or U22836 (N_22836,N_21080,N_21993);
nor U22837 (N_22837,N_22429,N_22069);
and U22838 (N_22838,N_22428,N_21125);
nor U22839 (N_22839,N_21094,N_21591);
xnor U22840 (N_22840,N_21189,N_21682);
nor U22841 (N_22841,N_21760,N_21418);
xor U22842 (N_22842,N_21743,N_22038);
nor U22843 (N_22843,N_21633,N_21058);
nand U22844 (N_22844,N_22367,N_21767);
nand U22845 (N_22845,N_21183,N_21323);
or U22846 (N_22846,N_21157,N_22259);
xnor U22847 (N_22847,N_21727,N_21924);
nor U22848 (N_22848,N_22365,N_22159);
or U22849 (N_22849,N_21450,N_21083);
or U22850 (N_22850,N_21462,N_21178);
xor U22851 (N_22851,N_21956,N_21749);
and U22852 (N_22852,N_22054,N_22357);
nand U22853 (N_22853,N_21222,N_21926);
and U22854 (N_22854,N_21635,N_21062);
or U22855 (N_22855,N_22474,N_21008);
and U22856 (N_22856,N_21967,N_21031);
and U22857 (N_22857,N_22387,N_21954);
nand U22858 (N_22858,N_22062,N_22034);
nor U22859 (N_22859,N_21460,N_21286);
or U22860 (N_22860,N_21035,N_21188);
or U22861 (N_22861,N_21791,N_21305);
nor U22862 (N_22862,N_21367,N_21112);
or U22863 (N_22863,N_22223,N_21588);
and U22864 (N_22864,N_22112,N_21123);
nor U22865 (N_22865,N_21321,N_21020);
xnor U22866 (N_22866,N_21606,N_21992);
xnor U22867 (N_22867,N_21840,N_22227);
nor U22868 (N_22868,N_22313,N_22009);
nor U22869 (N_22869,N_21517,N_21021);
xnor U22870 (N_22870,N_21789,N_21674);
nand U22871 (N_22871,N_21532,N_21848);
xnor U22872 (N_22872,N_22059,N_21069);
and U22873 (N_22873,N_22412,N_22025);
and U22874 (N_22874,N_21799,N_21559);
xor U22875 (N_22875,N_22411,N_22013);
nand U22876 (N_22876,N_21696,N_21061);
nand U22877 (N_22877,N_21156,N_21239);
and U22878 (N_22878,N_21393,N_21981);
xnor U22879 (N_22879,N_21702,N_21781);
or U22880 (N_22880,N_22300,N_21246);
and U22881 (N_22881,N_21824,N_21493);
nand U22882 (N_22882,N_21510,N_22420);
or U22883 (N_22883,N_22229,N_21612);
and U22884 (N_22884,N_21024,N_22058);
nand U22885 (N_22885,N_21944,N_21747);
nand U22886 (N_22886,N_22113,N_22319);
xor U22887 (N_22887,N_21377,N_21288);
or U22888 (N_22888,N_21215,N_21003);
nor U22889 (N_22889,N_21579,N_22295);
xnor U22890 (N_22890,N_22254,N_21997);
nand U22891 (N_22891,N_21133,N_21086);
or U22892 (N_22892,N_22234,N_22057);
or U22893 (N_22893,N_21347,N_21027);
or U22894 (N_22894,N_21999,N_21470);
nand U22895 (N_22895,N_21807,N_21231);
or U22896 (N_22896,N_21147,N_21371);
nand U22897 (N_22897,N_21397,N_22468);
xor U22898 (N_22898,N_21906,N_21354);
and U22899 (N_22899,N_21313,N_21864);
xnor U22900 (N_22900,N_22361,N_22071);
nand U22901 (N_22901,N_21708,N_21658);
or U22902 (N_22902,N_21811,N_22224);
or U22903 (N_22903,N_21511,N_21725);
nand U22904 (N_22904,N_22108,N_22153);
xor U22905 (N_22905,N_21915,N_22354);
or U22906 (N_22906,N_22249,N_21717);
or U22907 (N_22907,N_21079,N_21394);
xnor U22908 (N_22908,N_22158,N_21675);
or U22909 (N_22909,N_22453,N_21973);
nor U22910 (N_22910,N_21155,N_21428);
xor U22911 (N_22911,N_21783,N_21570);
nor U22912 (N_22912,N_21091,N_21174);
nor U22913 (N_22913,N_21433,N_21687);
nand U22914 (N_22914,N_22008,N_22096);
or U22915 (N_22915,N_21547,N_21208);
xor U22916 (N_22916,N_22452,N_21268);
nor U22917 (N_22917,N_21707,N_21186);
and U22918 (N_22918,N_22434,N_21073);
xnor U22919 (N_22919,N_21728,N_21684);
and U22920 (N_22920,N_21341,N_22377);
nand U22921 (N_22921,N_21937,N_21935);
or U22922 (N_22922,N_21381,N_21124);
nor U22923 (N_22923,N_22000,N_21256);
xor U22924 (N_22924,N_22048,N_21134);
nor U22925 (N_22925,N_22347,N_21913);
and U22926 (N_22926,N_21252,N_21786);
nor U22927 (N_22927,N_22142,N_22356);
and U22928 (N_22928,N_22026,N_21432);
nand U22929 (N_22929,N_21199,N_21297);
or U22930 (N_22930,N_21795,N_22178);
nand U22931 (N_22931,N_21498,N_21522);
xor U22932 (N_22932,N_22128,N_21670);
nor U22933 (N_22933,N_21892,N_21434);
xor U22934 (N_22934,N_21346,N_21064);
and U22935 (N_22935,N_22176,N_22475);
xnor U22936 (N_22936,N_22456,N_22287);
and U22937 (N_22937,N_21977,N_22094);
nand U22938 (N_22938,N_21645,N_21929);
and U22939 (N_22939,N_21154,N_22349);
or U22940 (N_22940,N_22156,N_22012);
and U22941 (N_22941,N_22432,N_21881);
xor U22942 (N_22942,N_21013,N_21701);
xor U22943 (N_22943,N_21480,N_21364);
and U22944 (N_22944,N_22273,N_22376);
or U22945 (N_22945,N_22302,N_21318);
xnor U22946 (N_22946,N_21089,N_21216);
and U22947 (N_22947,N_22459,N_21329);
or U22948 (N_22948,N_22455,N_22061);
xor U22949 (N_22949,N_22002,N_21669);
xnor U22950 (N_22950,N_22166,N_21220);
xnor U22951 (N_22951,N_22315,N_21387);
xnor U22952 (N_22952,N_22438,N_21085);
nor U22953 (N_22953,N_21551,N_21773);
and U22954 (N_22954,N_22092,N_21751);
nand U22955 (N_22955,N_22240,N_22495);
or U22956 (N_22956,N_22097,N_21048);
or U22957 (N_22957,N_21350,N_22415);
or U22958 (N_22958,N_21905,N_22278);
xnor U22959 (N_22959,N_21046,N_21282);
and U22960 (N_22960,N_22035,N_21424);
nor U22961 (N_22961,N_21114,N_21800);
nand U22962 (N_22962,N_22407,N_22484);
nor U22963 (N_22963,N_21628,N_21723);
or U22964 (N_22964,N_22401,N_21119);
or U22965 (N_22965,N_21415,N_22011);
nor U22966 (N_22966,N_22106,N_21456);
and U22967 (N_22967,N_22255,N_21316);
nor U22968 (N_22968,N_21804,N_21398);
and U22969 (N_22969,N_22084,N_21093);
nand U22970 (N_22970,N_21385,N_22184);
xor U22971 (N_22971,N_21867,N_21609);
or U22972 (N_22972,N_22188,N_21782);
xnor U22973 (N_22973,N_22161,N_21002);
nand U22974 (N_22974,N_22151,N_21904);
or U22975 (N_22975,N_21014,N_21076);
or U22976 (N_22976,N_22228,N_21544);
and U22977 (N_22977,N_21104,N_21485);
xnor U22978 (N_22978,N_21561,N_22126);
nor U22979 (N_22979,N_21798,N_21831);
or U22980 (N_22980,N_22088,N_21531);
xnor U22981 (N_22981,N_22100,N_21446);
nor U22982 (N_22982,N_21078,N_22216);
xor U22983 (N_22983,N_21891,N_21936);
nor U22984 (N_22984,N_21029,N_22130);
nor U22985 (N_22985,N_21376,N_21621);
or U22986 (N_22986,N_21857,N_22125);
nand U22987 (N_22987,N_21408,N_21307);
nand U22988 (N_22988,N_21627,N_21224);
xnor U22989 (N_22989,N_22345,N_21484);
nor U22990 (N_22990,N_21686,N_21585);
and U22991 (N_22991,N_22416,N_22052);
nor U22992 (N_22992,N_21665,N_21352);
xnor U22993 (N_22993,N_21486,N_22426);
xnor U22994 (N_22994,N_21167,N_22460);
xor U22995 (N_22995,N_21521,N_22186);
or U22996 (N_22996,N_21870,N_21006);
nor U22997 (N_22997,N_21468,N_21257);
nor U22998 (N_22998,N_21056,N_21693);
nand U22999 (N_22999,N_22422,N_21836);
and U23000 (N_23000,N_21898,N_22266);
xor U23001 (N_23001,N_21837,N_21710);
or U23002 (N_23002,N_21298,N_22404);
nand U23003 (N_23003,N_21541,N_22245);
nor U23004 (N_23004,N_22473,N_21358);
nor U23005 (N_23005,N_21601,N_21138);
xor U23006 (N_23006,N_21413,N_21343);
or U23007 (N_23007,N_21342,N_21401);
xor U23008 (N_23008,N_21311,N_21950);
nor U23009 (N_23009,N_21324,N_21276);
or U23010 (N_23010,N_22448,N_21226);
nand U23011 (N_23011,N_21721,N_21380);
nor U23012 (N_23012,N_21471,N_21903);
nor U23013 (N_23013,N_21797,N_21974);
xor U23014 (N_23014,N_21067,N_21639);
or U23015 (N_23015,N_21430,N_21416);
or U23016 (N_23016,N_22081,N_21249);
and U23017 (N_23017,N_22479,N_21140);
and U23018 (N_23018,N_22040,N_21948);
xor U23019 (N_23019,N_22164,N_22033);
xor U23020 (N_23020,N_21197,N_21304);
nor U23021 (N_23021,N_21360,N_21248);
nor U23022 (N_23022,N_21319,N_21955);
and U23023 (N_23023,N_22177,N_21126);
and U23024 (N_23024,N_22258,N_22217);
and U23025 (N_23025,N_21756,N_21383);
and U23026 (N_23026,N_22360,N_22122);
xor U23027 (N_23027,N_21740,N_21569);
or U23028 (N_23028,N_22311,N_21187);
nor U23029 (N_23029,N_22293,N_21295);
or U23030 (N_23030,N_21237,N_22461);
or U23031 (N_23031,N_22400,N_21103);
nor U23032 (N_23032,N_22355,N_22277);
xnor U23033 (N_23033,N_21449,N_21148);
xor U23034 (N_23034,N_22290,N_22248);
or U23035 (N_23035,N_21883,N_22306);
and U23036 (N_23036,N_22104,N_21300);
xnor U23037 (N_23037,N_21514,N_21190);
or U23038 (N_23038,N_22288,N_22464);
nand U23039 (N_23039,N_22389,N_21117);
nand U23040 (N_23040,N_22336,N_22430);
nor U23041 (N_23041,N_21931,N_21979);
or U23042 (N_23042,N_21245,N_21871);
nand U23043 (N_23043,N_21461,N_21576);
and U23044 (N_23044,N_21223,N_21250);
nor U23045 (N_23045,N_21825,N_21850);
nand U23046 (N_23046,N_21894,N_21090);
nor U23047 (N_23047,N_22343,N_22446);
and U23048 (N_23048,N_21868,N_21271);
and U23049 (N_23049,N_22309,N_21004);
nor U23050 (N_23050,N_22165,N_22470);
and U23051 (N_23051,N_21741,N_22146);
nand U23052 (N_23052,N_21650,N_21709);
and U23053 (N_23053,N_21353,N_21557);
or U23054 (N_23054,N_21978,N_22325);
and U23055 (N_23055,N_21697,N_21678);
and U23056 (N_23056,N_21614,N_22215);
or U23057 (N_23057,N_21793,N_22378);
and U23058 (N_23058,N_22397,N_21506);
xnor U23059 (N_23059,N_22015,N_22324);
nand U23060 (N_23060,N_22242,N_21491);
and U23061 (N_23061,N_21327,N_21097);
nand U23062 (N_23062,N_21158,N_22144);
nor U23063 (N_23063,N_22032,N_21207);
xnor U23064 (N_23064,N_22124,N_21254);
and U23065 (N_23065,N_21879,N_22450);
nor U23066 (N_23066,N_22206,N_21885);
and U23067 (N_23067,N_21739,N_21615);
and U23068 (N_23068,N_21459,N_22207);
nand U23069 (N_23069,N_21930,N_22291);
nor U23070 (N_23070,N_21772,N_22388);
or U23071 (N_23071,N_21901,N_21982);
nand U23072 (N_23072,N_21679,N_21373);
nand U23073 (N_23073,N_21939,N_21241);
xor U23074 (N_23074,N_21922,N_22087);
xor U23075 (N_23075,N_21555,N_21952);
nand U23076 (N_23076,N_22172,N_22107);
nor U23077 (N_23077,N_22380,N_21827);
and U23078 (N_23078,N_21719,N_21700);
nor U23079 (N_23079,N_21624,N_22304);
nor U23080 (N_23080,N_21168,N_21442);
xor U23081 (N_23081,N_21072,N_21907);
nor U23082 (N_23082,N_21406,N_21242);
nand U23083 (N_23083,N_22403,N_22134);
and U23084 (N_23084,N_21475,N_21699);
nand U23085 (N_23085,N_21704,N_22431);
nand U23086 (N_23086,N_21660,N_21357);
nor U23087 (N_23087,N_22314,N_22085);
and U23088 (N_23088,N_21845,N_21469);
xnor U23089 (N_23089,N_21947,N_21890);
or U23090 (N_23090,N_22322,N_21054);
nor U23091 (N_23091,N_22145,N_21294);
and U23092 (N_23092,N_21730,N_22299);
or U23093 (N_23093,N_22102,N_21280);
and U23094 (N_23094,N_22098,N_21991);
xor U23095 (N_23095,N_21985,N_22292);
nor U23096 (N_23096,N_21441,N_21494);
nand U23097 (N_23097,N_21243,N_22471);
nand U23098 (N_23098,N_22036,N_21488);
nor U23099 (N_23099,N_21333,N_21363);
or U23100 (N_23100,N_21326,N_21007);
nand U23101 (N_23101,N_21478,N_22419);
or U23102 (N_23102,N_21813,N_22279);
xor U23103 (N_23103,N_21722,N_22005);
nand U23104 (N_23104,N_22454,N_22214);
xnor U23105 (N_23105,N_21423,N_21667);
and U23106 (N_23106,N_21182,N_21152);
and U23107 (N_23107,N_22393,N_22171);
nor U23108 (N_23108,N_22488,N_22275);
nand U23109 (N_23109,N_21976,N_21995);
nand U23110 (N_23110,N_21396,N_22320);
or U23111 (N_23111,N_21161,N_22099);
xor U23112 (N_23112,N_21706,N_21994);
or U23113 (N_23113,N_21052,N_21108);
xnor U23114 (N_23114,N_22296,N_22447);
xnor U23115 (N_23115,N_22199,N_22137);
nand U23116 (N_23116,N_22072,N_21957);
nand U23117 (N_23117,N_21536,N_22359);
nor U23118 (N_23118,N_21619,N_22006);
or U23119 (N_23119,N_21481,N_21766);
xnor U23120 (N_23120,N_21554,N_21445);
and U23121 (N_23121,N_21733,N_21636);
xnor U23122 (N_23122,N_22021,N_22031);
nand U23123 (N_23123,N_21438,N_22152);
and U23124 (N_23124,N_22241,N_22138);
xnor U23125 (N_23125,N_21010,N_21695);
nor U23126 (N_23126,N_21654,N_21036);
and U23127 (N_23127,N_21574,N_21616);
nor U23128 (N_23128,N_21334,N_22457);
and U23129 (N_23129,N_21984,N_22333);
nor U23130 (N_23130,N_22183,N_21941);
nand U23131 (N_23131,N_21267,N_21828);
xor U23132 (N_23132,N_21648,N_21146);
nand U23133 (N_23133,N_22163,N_21858);
and U23134 (N_23134,N_22068,N_22133);
nor U23135 (N_23135,N_21668,N_21962);
and U23136 (N_23136,N_21314,N_21986);
or U23137 (N_23137,N_21410,N_21680);
nand U23138 (N_23138,N_21911,N_22253);
and U23139 (N_23139,N_22243,N_21259);
and U23140 (N_23140,N_22211,N_21113);
or U23141 (N_23141,N_21726,N_21272);
nor U23142 (N_23142,N_21414,N_22131);
nand U23143 (N_23143,N_21016,N_21638);
nor U23144 (N_23144,N_21301,N_21940);
and U23145 (N_23145,N_21283,N_21843);
and U23146 (N_23146,N_22017,N_22063);
or U23147 (N_23147,N_21970,N_21818);
and U23148 (N_23148,N_22101,N_21309);
and U23149 (N_23149,N_21455,N_21688);
nor U23150 (N_23150,N_21921,N_21583);
or U23151 (N_23151,N_22294,N_22263);
nor U23152 (N_23152,N_21504,N_21026);
or U23153 (N_23153,N_21652,N_21419);
and U23154 (N_23154,N_21053,N_21735);
nor U23155 (N_23155,N_22141,N_21834);
xnor U23156 (N_23156,N_21815,N_21754);
xor U23157 (N_23157,N_21835,N_21263);
xor U23158 (N_23158,N_21777,N_22046);
and U23159 (N_23159,N_22442,N_22047);
nor U23160 (N_23160,N_21875,N_21296);
nor U23161 (N_23161,N_21107,N_21417);
nor U23162 (N_23162,N_21964,N_22264);
xor U23163 (N_23163,N_21425,N_21122);
xnor U23164 (N_23164,N_21018,N_22251);
nand U23165 (N_23165,N_22003,N_22236);
and U23166 (N_23166,N_22095,N_22064);
xor U23167 (N_23167,N_22498,N_22312);
or U23168 (N_23168,N_21447,N_21136);
xor U23169 (N_23169,N_21355,N_21775);
nor U23170 (N_23170,N_21844,N_21368);
xnor U23171 (N_23171,N_21692,N_22340);
or U23172 (N_23172,N_21816,N_21920);
nand U23173 (N_23173,N_21597,N_22439);
or U23174 (N_23174,N_21672,N_21711);
xnor U23175 (N_23175,N_21598,N_21429);
xor U23176 (N_23176,N_22105,N_21440);
or U23177 (N_23177,N_21542,N_21370);
xnor U23178 (N_23178,N_22445,N_21715);
nand U23179 (N_23179,N_22384,N_21421);
nand U23180 (N_23180,N_21971,N_21116);
or U23181 (N_23181,N_21359,N_21458);
nand U23182 (N_23182,N_21041,N_22246);
or U23183 (N_23183,N_21873,N_21177);
and U23184 (N_23184,N_22472,N_22195);
nor U23185 (N_23185,N_21482,N_21435);
nand U23186 (N_23186,N_21851,N_22252);
xor U23187 (N_23187,N_21833,N_22050);
nand U23188 (N_23188,N_21942,N_21975);
and U23189 (N_23189,N_21265,N_21402);
and U23190 (N_23190,N_22381,N_22362);
nand U23191 (N_23191,N_22379,N_21832);
xor U23192 (N_23192,N_21626,N_21448);
nor U23193 (N_23193,N_21918,N_22238);
and U23194 (N_23194,N_21312,N_22310);
or U23195 (N_23195,N_21400,N_21204);
or U23196 (N_23196,N_22053,N_21291);
and U23197 (N_23197,N_22192,N_22305);
nor U23198 (N_23198,N_22489,N_22179);
xor U23199 (N_23199,N_21592,N_21866);
nand U23200 (N_23200,N_21776,N_21345);
nand U23201 (N_23201,N_22070,N_22149);
and U23202 (N_23202,N_22049,N_22148);
or U23203 (N_23203,N_21390,N_21501);
or U23204 (N_23204,N_22103,N_22268);
xor U23205 (N_23205,N_21366,N_22169);
or U23206 (N_23206,N_21251,N_22414);
nor U23207 (N_23207,N_21630,N_21649);
or U23208 (N_23208,N_21822,N_22417);
nand U23209 (N_23209,N_21516,N_21617);
nor U23210 (N_23210,N_21537,N_22337);
and U23211 (N_23211,N_21500,N_21150);
xor U23212 (N_23212,N_21849,N_21399);
and U23213 (N_23213,N_22083,N_22423);
or U23214 (N_23214,N_21887,N_22427);
nor U23215 (N_23215,N_22440,N_21005);
or U23216 (N_23216,N_21261,N_22123);
nor U23217 (N_23217,N_22490,N_21111);
and U23218 (N_23218,N_21179,N_22352);
nor U23219 (N_23219,N_22399,N_22418);
nor U23220 (N_23220,N_21193,N_21705);
or U23221 (N_23221,N_22189,N_22110);
nand U23222 (N_23222,N_22334,N_21233);
xnor U23223 (N_23223,N_21919,N_21540);
nand U23224 (N_23224,N_22441,N_22281);
xor U23225 (N_23225,N_22366,N_22338);
nand U23226 (N_23226,N_21066,N_21852);
or U23227 (N_23227,N_21582,N_22478);
nor U23228 (N_23228,N_21820,N_22180);
and U23229 (N_23229,N_22342,N_21218);
xnor U23230 (N_23230,N_22077,N_21959);
nand U23231 (N_23231,N_21900,N_21987);
or U23232 (N_23232,N_22232,N_21483);
nor U23233 (N_23233,N_21191,N_21859);
xor U23234 (N_23234,N_22150,N_21338);
and U23235 (N_23235,N_21714,N_21110);
and U23236 (N_23236,N_21519,N_21142);
xor U23237 (N_23237,N_22194,N_22219);
xor U23238 (N_23238,N_21623,N_21451);
or U23239 (N_23239,N_21411,N_21573);
or U23240 (N_23240,N_21810,N_21902);
and U23241 (N_23241,N_21515,N_22007);
nor U23242 (N_23242,N_22483,N_22395);
nor U23243 (N_23243,N_21989,N_21070);
xnor U23244 (N_23244,N_21603,N_22120);
or U23245 (N_23245,N_21742,N_21095);
xor U23246 (N_23246,N_21200,N_21115);
and U23247 (N_23247,N_21139,N_21790);
nor U23248 (N_23248,N_21299,N_21683);
xor U23249 (N_23249,N_22383,N_22190);
nor U23250 (N_23250,N_21396,N_21741);
xnor U23251 (N_23251,N_22026,N_22055);
nor U23252 (N_23252,N_21049,N_22032);
nand U23253 (N_23253,N_21974,N_22290);
nand U23254 (N_23254,N_21382,N_21371);
nand U23255 (N_23255,N_22150,N_22443);
and U23256 (N_23256,N_21851,N_21224);
nand U23257 (N_23257,N_22142,N_21693);
or U23258 (N_23258,N_21396,N_22081);
nand U23259 (N_23259,N_21228,N_21272);
and U23260 (N_23260,N_22442,N_21212);
xnor U23261 (N_23261,N_22209,N_21239);
xor U23262 (N_23262,N_21087,N_22344);
nor U23263 (N_23263,N_21250,N_21616);
nor U23264 (N_23264,N_22288,N_22281);
and U23265 (N_23265,N_21044,N_21437);
nor U23266 (N_23266,N_21517,N_21960);
or U23267 (N_23267,N_21678,N_22443);
nand U23268 (N_23268,N_22207,N_21690);
nor U23269 (N_23269,N_21441,N_21177);
xor U23270 (N_23270,N_21421,N_21536);
nand U23271 (N_23271,N_21482,N_22215);
or U23272 (N_23272,N_21842,N_21077);
or U23273 (N_23273,N_21945,N_21630);
and U23274 (N_23274,N_21151,N_21139);
nand U23275 (N_23275,N_21489,N_22491);
xor U23276 (N_23276,N_21661,N_21427);
and U23277 (N_23277,N_21035,N_21487);
nand U23278 (N_23278,N_21717,N_22386);
and U23279 (N_23279,N_22027,N_22031);
or U23280 (N_23280,N_21918,N_22376);
nor U23281 (N_23281,N_21733,N_21270);
xor U23282 (N_23282,N_21835,N_22104);
nand U23283 (N_23283,N_21612,N_22005);
and U23284 (N_23284,N_21753,N_21591);
or U23285 (N_23285,N_21702,N_21244);
xnor U23286 (N_23286,N_21779,N_22316);
xnor U23287 (N_23287,N_21192,N_21634);
nand U23288 (N_23288,N_21347,N_21326);
xor U23289 (N_23289,N_21181,N_22426);
nor U23290 (N_23290,N_21855,N_21451);
xor U23291 (N_23291,N_21646,N_21636);
xor U23292 (N_23292,N_22366,N_21803);
nor U23293 (N_23293,N_22098,N_21434);
and U23294 (N_23294,N_22288,N_22225);
or U23295 (N_23295,N_21742,N_21901);
and U23296 (N_23296,N_22427,N_21563);
xor U23297 (N_23297,N_21698,N_21611);
xnor U23298 (N_23298,N_21824,N_21321);
or U23299 (N_23299,N_21778,N_21785);
nand U23300 (N_23300,N_21765,N_21016);
or U23301 (N_23301,N_22412,N_21039);
nor U23302 (N_23302,N_21816,N_22007);
or U23303 (N_23303,N_21296,N_21522);
nand U23304 (N_23304,N_22195,N_21029);
xnor U23305 (N_23305,N_21494,N_22181);
nand U23306 (N_23306,N_21495,N_21323);
nand U23307 (N_23307,N_22088,N_21150);
xor U23308 (N_23308,N_21155,N_22499);
nand U23309 (N_23309,N_21027,N_22311);
and U23310 (N_23310,N_21143,N_21471);
nor U23311 (N_23311,N_21030,N_21067);
xnor U23312 (N_23312,N_21036,N_22093);
nand U23313 (N_23313,N_22338,N_22471);
xor U23314 (N_23314,N_21027,N_21534);
nor U23315 (N_23315,N_21021,N_21291);
xor U23316 (N_23316,N_22375,N_21149);
xnor U23317 (N_23317,N_21015,N_21014);
nor U23318 (N_23318,N_22461,N_21263);
or U23319 (N_23319,N_21966,N_21997);
nor U23320 (N_23320,N_22140,N_21176);
and U23321 (N_23321,N_22362,N_21201);
nor U23322 (N_23322,N_21626,N_22222);
nand U23323 (N_23323,N_21450,N_22119);
xnor U23324 (N_23324,N_21057,N_21761);
and U23325 (N_23325,N_21135,N_22254);
and U23326 (N_23326,N_21213,N_21818);
and U23327 (N_23327,N_21626,N_22170);
nand U23328 (N_23328,N_22209,N_22388);
or U23329 (N_23329,N_21575,N_21451);
and U23330 (N_23330,N_22205,N_22491);
and U23331 (N_23331,N_22227,N_21216);
nor U23332 (N_23332,N_22229,N_22318);
and U23333 (N_23333,N_22407,N_21190);
nor U23334 (N_23334,N_21511,N_21537);
nand U23335 (N_23335,N_21645,N_21949);
nand U23336 (N_23336,N_22320,N_21486);
xnor U23337 (N_23337,N_21684,N_22297);
nor U23338 (N_23338,N_22463,N_22114);
nand U23339 (N_23339,N_22404,N_21391);
and U23340 (N_23340,N_21332,N_21244);
xor U23341 (N_23341,N_21048,N_21669);
nand U23342 (N_23342,N_22324,N_21743);
or U23343 (N_23343,N_22070,N_21232);
or U23344 (N_23344,N_22381,N_22003);
and U23345 (N_23345,N_21062,N_21969);
nand U23346 (N_23346,N_21106,N_22013);
and U23347 (N_23347,N_22286,N_21436);
nand U23348 (N_23348,N_21829,N_21585);
nor U23349 (N_23349,N_21199,N_21078);
nor U23350 (N_23350,N_22008,N_21105);
or U23351 (N_23351,N_21410,N_21161);
nand U23352 (N_23352,N_21518,N_22268);
and U23353 (N_23353,N_21041,N_21076);
nor U23354 (N_23354,N_21110,N_21581);
nand U23355 (N_23355,N_21990,N_21246);
and U23356 (N_23356,N_21739,N_22009);
xnor U23357 (N_23357,N_21204,N_21098);
xor U23358 (N_23358,N_22158,N_21148);
or U23359 (N_23359,N_21892,N_21646);
and U23360 (N_23360,N_21494,N_21269);
nor U23361 (N_23361,N_22396,N_21876);
nand U23362 (N_23362,N_21203,N_21100);
xnor U23363 (N_23363,N_22251,N_21662);
or U23364 (N_23364,N_21876,N_22319);
nand U23365 (N_23365,N_22069,N_21077);
xor U23366 (N_23366,N_21928,N_21071);
xor U23367 (N_23367,N_21048,N_21873);
nand U23368 (N_23368,N_21933,N_21427);
or U23369 (N_23369,N_21073,N_21618);
and U23370 (N_23370,N_21514,N_21670);
and U23371 (N_23371,N_21286,N_22257);
and U23372 (N_23372,N_22319,N_22269);
nor U23373 (N_23373,N_22457,N_21233);
or U23374 (N_23374,N_21170,N_21749);
and U23375 (N_23375,N_21539,N_21791);
nand U23376 (N_23376,N_21851,N_21314);
nor U23377 (N_23377,N_22453,N_21925);
nand U23378 (N_23378,N_22492,N_22381);
nor U23379 (N_23379,N_22219,N_21160);
or U23380 (N_23380,N_22109,N_22004);
nor U23381 (N_23381,N_21422,N_22306);
xor U23382 (N_23382,N_21730,N_22287);
xor U23383 (N_23383,N_21114,N_21072);
or U23384 (N_23384,N_21032,N_22323);
xnor U23385 (N_23385,N_22476,N_21733);
nor U23386 (N_23386,N_22079,N_21182);
xor U23387 (N_23387,N_21325,N_21354);
or U23388 (N_23388,N_22337,N_21939);
nand U23389 (N_23389,N_22404,N_21295);
xnor U23390 (N_23390,N_21352,N_22100);
nand U23391 (N_23391,N_21462,N_21514);
nand U23392 (N_23392,N_21218,N_21191);
or U23393 (N_23393,N_22456,N_22029);
nor U23394 (N_23394,N_22114,N_22107);
xor U23395 (N_23395,N_21019,N_21511);
nand U23396 (N_23396,N_21567,N_21375);
xnor U23397 (N_23397,N_21877,N_22398);
or U23398 (N_23398,N_21936,N_21439);
and U23399 (N_23399,N_22155,N_22325);
and U23400 (N_23400,N_21734,N_22249);
or U23401 (N_23401,N_21755,N_21161);
nor U23402 (N_23402,N_21850,N_21268);
nor U23403 (N_23403,N_22031,N_21606);
nand U23404 (N_23404,N_22499,N_21361);
and U23405 (N_23405,N_22219,N_22084);
nor U23406 (N_23406,N_21273,N_21040);
xor U23407 (N_23407,N_22016,N_22215);
nor U23408 (N_23408,N_21403,N_21789);
nor U23409 (N_23409,N_22413,N_21337);
nor U23410 (N_23410,N_21460,N_21557);
nand U23411 (N_23411,N_21357,N_21906);
and U23412 (N_23412,N_22198,N_22323);
or U23413 (N_23413,N_21587,N_21910);
or U23414 (N_23414,N_22092,N_21562);
xor U23415 (N_23415,N_21169,N_21423);
and U23416 (N_23416,N_22239,N_21872);
nor U23417 (N_23417,N_21261,N_21470);
nor U23418 (N_23418,N_22373,N_21686);
or U23419 (N_23419,N_21659,N_21943);
xnor U23420 (N_23420,N_22260,N_22428);
and U23421 (N_23421,N_21358,N_21958);
nor U23422 (N_23422,N_21604,N_21572);
and U23423 (N_23423,N_22421,N_21755);
and U23424 (N_23424,N_22298,N_22026);
and U23425 (N_23425,N_21461,N_22036);
or U23426 (N_23426,N_21662,N_21876);
nor U23427 (N_23427,N_21927,N_22333);
nand U23428 (N_23428,N_22122,N_22232);
and U23429 (N_23429,N_21262,N_21175);
xor U23430 (N_23430,N_21889,N_21753);
or U23431 (N_23431,N_22098,N_22286);
xnor U23432 (N_23432,N_21517,N_21830);
nor U23433 (N_23433,N_21828,N_21026);
nand U23434 (N_23434,N_22328,N_22429);
nor U23435 (N_23435,N_21308,N_21683);
nand U23436 (N_23436,N_22008,N_22076);
and U23437 (N_23437,N_22460,N_21712);
and U23438 (N_23438,N_22100,N_21265);
and U23439 (N_23439,N_21258,N_21162);
nand U23440 (N_23440,N_22104,N_21925);
nor U23441 (N_23441,N_21443,N_21035);
xor U23442 (N_23442,N_21997,N_21243);
xor U23443 (N_23443,N_21638,N_21308);
or U23444 (N_23444,N_21314,N_21422);
or U23445 (N_23445,N_21789,N_21573);
nand U23446 (N_23446,N_21986,N_21384);
and U23447 (N_23447,N_21495,N_21543);
nand U23448 (N_23448,N_22169,N_21038);
nand U23449 (N_23449,N_22123,N_21776);
and U23450 (N_23450,N_21313,N_21986);
xor U23451 (N_23451,N_21834,N_21683);
xnor U23452 (N_23452,N_22067,N_21671);
xor U23453 (N_23453,N_21499,N_21227);
xor U23454 (N_23454,N_21925,N_21929);
nor U23455 (N_23455,N_21972,N_21384);
and U23456 (N_23456,N_22262,N_21707);
and U23457 (N_23457,N_21243,N_21603);
nor U23458 (N_23458,N_21325,N_21875);
xnor U23459 (N_23459,N_21692,N_21629);
xor U23460 (N_23460,N_21156,N_22017);
or U23461 (N_23461,N_21004,N_22361);
and U23462 (N_23462,N_21220,N_21125);
nor U23463 (N_23463,N_21547,N_21024);
nor U23464 (N_23464,N_22144,N_21950);
nand U23465 (N_23465,N_21004,N_22303);
nand U23466 (N_23466,N_22350,N_22190);
xnor U23467 (N_23467,N_22241,N_21154);
xnor U23468 (N_23468,N_21848,N_21374);
xor U23469 (N_23469,N_21809,N_21046);
and U23470 (N_23470,N_21050,N_21435);
xnor U23471 (N_23471,N_21398,N_21537);
nand U23472 (N_23472,N_21672,N_21802);
nor U23473 (N_23473,N_21391,N_21833);
or U23474 (N_23474,N_21501,N_21015);
nor U23475 (N_23475,N_21912,N_21827);
nor U23476 (N_23476,N_21148,N_21263);
nor U23477 (N_23477,N_21295,N_22369);
nor U23478 (N_23478,N_21146,N_21140);
nor U23479 (N_23479,N_21139,N_21362);
and U23480 (N_23480,N_21815,N_21451);
or U23481 (N_23481,N_21161,N_21564);
xor U23482 (N_23482,N_21639,N_21156);
or U23483 (N_23483,N_21599,N_21865);
nor U23484 (N_23484,N_21393,N_22049);
nand U23485 (N_23485,N_21070,N_21183);
xor U23486 (N_23486,N_22317,N_21919);
nor U23487 (N_23487,N_22010,N_21106);
nor U23488 (N_23488,N_22262,N_21766);
nand U23489 (N_23489,N_21913,N_21637);
nor U23490 (N_23490,N_21592,N_21415);
nand U23491 (N_23491,N_22326,N_21656);
nor U23492 (N_23492,N_21229,N_22236);
nand U23493 (N_23493,N_21475,N_21618);
or U23494 (N_23494,N_22150,N_22077);
nor U23495 (N_23495,N_21885,N_21749);
and U23496 (N_23496,N_21841,N_22399);
xor U23497 (N_23497,N_22383,N_22255);
or U23498 (N_23498,N_21018,N_22375);
nor U23499 (N_23499,N_21955,N_21669);
nand U23500 (N_23500,N_21470,N_21452);
and U23501 (N_23501,N_21091,N_21100);
and U23502 (N_23502,N_21468,N_22256);
xor U23503 (N_23503,N_21980,N_22434);
nand U23504 (N_23504,N_22090,N_22381);
xor U23505 (N_23505,N_21153,N_21674);
nor U23506 (N_23506,N_21492,N_22036);
xnor U23507 (N_23507,N_21620,N_22138);
nor U23508 (N_23508,N_21597,N_21746);
or U23509 (N_23509,N_22364,N_21888);
xor U23510 (N_23510,N_21794,N_21483);
xor U23511 (N_23511,N_21962,N_21863);
and U23512 (N_23512,N_21549,N_21681);
or U23513 (N_23513,N_22259,N_21281);
or U23514 (N_23514,N_22279,N_21594);
xnor U23515 (N_23515,N_21075,N_21408);
nand U23516 (N_23516,N_22412,N_22011);
and U23517 (N_23517,N_21817,N_22293);
xnor U23518 (N_23518,N_21231,N_22285);
or U23519 (N_23519,N_21846,N_21070);
or U23520 (N_23520,N_21998,N_21881);
nand U23521 (N_23521,N_21439,N_21768);
and U23522 (N_23522,N_21173,N_21134);
xor U23523 (N_23523,N_21586,N_22111);
and U23524 (N_23524,N_22480,N_21396);
and U23525 (N_23525,N_21103,N_22456);
nor U23526 (N_23526,N_21671,N_22021);
nand U23527 (N_23527,N_22142,N_21907);
nor U23528 (N_23528,N_21408,N_22036);
nor U23529 (N_23529,N_21126,N_21849);
and U23530 (N_23530,N_22477,N_22384);
nor U23531 (N_23531,N_21080,N_22298);
xnor U23532 (N_23532,N_21853,N_21241);
nand U23533 (N_23533,N_21955,N_22413);
nor U23534 (N_23534,N_21978,N_21727);
xnor U23535 (N_23535,N_22319,N_21375);
nor U23536 (N_23536,N_21578,N_21419);
or U23537 (N_23537,N_22164,N_21503);
xor U23538 (N_23538,N_21489,N_21091);
or U23539 (N_23539,N_21544,N_21717);
nand U23540 (N_23540,N_21681,N_21845);
nor U23541 (N_23541,N_21640,N_21170);
or U23542 (N_23542,N_22133,N_21626);
xnor U23543 (N_23543,N_21571,N_22485);
or U23544 (N_23544,N_21029,N_21995);
xnor U23545 (N_23545,N_21370,N_21491);
and U23546 (N_23546,N_21965,N_22184);
xor U23547 (N_23547,N_21679,N_22316);
and U23548 (N_23548,N_21445,N_21034);
xor U23549 (N_23549,N_21597,N_22052);
or U23550 (N_23550,N_22321,N_21123);
nor U23551 (N_23551,N_21935,N_21030);
and U23552 (N_23552,N_21976,N_22472);
nand U23553 (N_23553,N_22181,N_21973);
and U23554 (N_23554,N_21986,N_21537);
and U23555 (N_23555,N_22467,N_21600);
nor U23556 (N_23556,N_22027,N_21653);
nor U23557 (N_23557,N_21544,N_21890);
or U23558 (N_23558,N_21316,N_21225);
or U23559 (N_23559,N_21745,N_22271);
and U23560 (N_23560,N_22027,N_22364);
nor U23561 (N_23561,N_22104,N_22458);
nand U23562 (N_23562,N_21031,N_22204);
and U23563 (N_23563,N_21084,N_22009);
nor U23564 (N_23564,N_21763,N_22455);
nand U23565 (N_23565,N_22294,N_21239);
nor U23566 (N_23566,N_21079,N_22301);
and U23567 (N_23567,N_21580,N_21953);
nor U23568 (N_23568,N_21218,N_21841);
nand U23569 (N_23569,N_21426,N_22267);
nor U23570 (N_23570,N_21556,N_22012);
or U23571 (N_23571,N_22178,N_21956);
nand U23572 (N_23572,N_21239,N_21812);
nor U23573 (N_23573,N_21579,N_21068);
xor U23574 (N_23574,N_21979,N_21570);
nand U23575 (N_23575,N_21501,N_21486);
or U23576 (N_23576,N_21129,N_21411);
or U23577 (N_23577,N_21375,N_21388);
and U23578 (N_23578,N_21546,N_22457);
xnor U23579 (N_23579,N_21660,N_21517);
nor U23580 (N_23580,N_21280,N_22174);
or U23581 (N_23581,N_21006,N_21860);
nor U23582 (N_23582,N_21256,N_22416);
nor U23583 (N_23583,N_21010,N_21103);
nand U23584 (N_23584,N_22325,N_21320);
nor U23585 (N_23585,N_21462,N_21834);
xnor U23586 (N_23586,N_22141,N_21796);
or U23587 (N_23587,N_21073,N_21932);
nand U23588 (N_23588,N_22296,N_21176);
nand U23589 (N_23589,N_22437,N_21486);
and U23590 (N_23590,N_22395,N_21588);
nor U23591 (N_23591,N_22187,N_21997);
nand U23592 (N_23592,N_21443,N_21458);
nand U23593 (N_23593,N_21805,N_21372);
xnor U23594 (N_23594,N_22002,N_22187);
nand U23595 (N_23595,N_21630,N_21308);
nor U23596 (N_23596,N_21115,N_21970);
and U23597 (N_23597,N_21672,N_21911);
nor U23598 (N_23598,N_21685,N_21570);
nand U23599 (N_23599,N_21786,N_21628);
nand U23600 (N_23600,N_21324,N_21046);
xnor U23601 (N_23601,N_21056,N_22154);
nor U23602 (N_23602,N_21112,N_22202);
nor U23603 (N_23603,N_21556,N_21345);
xnor U23604 (N_23604,N_21768,N_21689);
xnor U23605 (N_23605,N_22033,N_21482);
and U23606 (N_23606,N_22100,N_22348);
nand U23607 (N_23607,N_21976,N_22017);
xor U23608 (N_23608,N_22461,N_22011);
nor U23609 (N_23609,N_21550,N_21887);
xnor U23610 (N_23610,N_21133,N_21474);
and U23611 (N_23611,N_21268,N_21831);
nor U23612 (N_23612,N_21141,N_21765);
and U23613 (N_23613,N_21911,N_21217);
nor U23614 (N_23614,N_22294,N_21453);
xnor U23615 (N_23615,N_21632,N_21313);
and U23616 (N_23616,N_21440,N_21910);
nand U23617 (N_23617,N_21715,N_21659);
or U23618 (N_23618,N_22071,N_22005);
nor U23619 (N_23619,N_21668,N_21928);
or U23620 (N_23620,N_21781,N_21434);
or U23621 (N_23621,N_22421,N_21476);
nor U23622 (N_23622,N_21057,N_21933);
nor U23623 (N_23623,N_22185,N_22442);
or U23624 (N_23624,N_21520,N_21687);
or U23625 (N_23625,N_21807,N_22350);
nor U23626 (N_23626,N_21659,N_22017);
nor U23627 (N_23627,N_21276,N_21029);
and U23628 (N_23628,N_21629,N_22335);
xnor U23629 (N_23629,N_22490,N_21141);
nor U23630 (N_23630,N_21996,N_21231);
nor U23631 (N_23631,N_21143,N_21107);
and U23632 (N_23632,N_21782,N_21224);
nor U23633 (N_23633,N_22119,N_21009);
xor U23634 (N_23634,N_21549,N_21450);
and U23635 (N_23635,N_21572,N_22368);
or U23636 (N_23636,N_22297,N_21303);
xnor U23637 (N_23637,N_22073,N_21802);
or U23638 (N_23638,N_21265,N_21476);
nor U23639 (N_23639,N_21004,N_22403);
and U23640 (N_23640,N_21825,N_22067);
nand U23641 (N_23641,N_21602,N_21333);
and U23642 (N_23642,N_22148,N_22307);
nor U23643 (N_23643,N_21162,N_21987);
xor U23644 (N_23644,N_21663,N_21391);
nand U23645 (N_23645,N_22069,N_21046);
or U23646 (N_23646,N_22429,N_22254);
nand U23647 (N_23647,N_21806,N_21509);
nand U23648 (N_23648,N_21772,N_21059);
nor U23649 (N_23649,N_21245,N_22076);
nand U23650 (N_23650,N_21551,N_21681);
nand U23651 (N_23651,N_21831,N_22434);
xnor U23652 (N_23652,N_21624,N_22146);
or U23653 (N_23653,N_22408,N_21957);
nand U23654 (N_23654,N_21508,N_22077);
nand U23655 (N_23655,N_21768,N_21161);
xor U23656 (N_23656,N_21480,N_22053);
nor U23657 (N_23657,N_21979,N_21130);
or U23658 (N_23658,N_21918,N_21091);
nor U23659 (N_23659,N_21097,N_21851);
xor U23660 (N_23660,N_21392,N_21751);
or U23661 (N_23661,N_21890,N_21052);
or U23662 (N_23662,N_21721,N_22181);
or U23663 (N_23663,N_21518,N_21243);
nor U23664 (N_23664,N_21486,N_21146);
nor U23665 (N_23665,N_22100,N_21748);
xnor U23666 (N_23666,N_22020,N_21984);
and U23667 (N_23667,N_21107,N_21965);
nor U23668 (N_23668,N_22441,N_22134);
nor U23669 (N_23669,N_21371,N_21146);
and U23670 (N_23670,N_22345,N_21040);
nand U23671 (N_23671,N_21729,N_22095);
or U23672 (N_23672,N_21951,N_21284);
nor U23673 (N_23673,N_21720,N_21054);
nand U23674 (N_23674,N_21184,N_21537);
xor U23675 (N_23675,N_21583,N_21101);
nor U23676 (N_23676,N_22250,N_21286);
and U23677 (N_23677,N_22280,N_21318);
or U23678 (N_23678,N_21757,N_21238);
or U23679 (N_23679,N_22414,N_22027);
or U23680 (N_23680,N_21575,N_21352);
xor U23681 (N_23681,N_22386,N_21728);
nand U23682 (N_23682,N_21786,N_21228);
nor U23683 (N_23683,N_21739,N_21659);
nand U23684 (N_23684,N_21435,N_21356);
or U23685 (N_23685,N_22305,N_22297);
or U23686 (N_23686,N_21239,N_21538);
nand U23687 (N_23687,N_21089,N_22314);
and U23688 (N_23688,N_21190,N_21841);
and U23689 (N_23689,N_22038,N_21795);
xor U23690 (N_23690,N_21213,N_21965);
and U23691 (N_23691,N_21580,N_21400);
xor U23692 (N_23692,N_22302,N_21656);
xnor U23693 (N_23693,N_21944,N_21312);
xnor U23694 (N_23694,N_22332,N_21400);
and U23695 (N_23695,N_21079,N_22123);
nor U23696 (N_23696,N_21364,N_21398);
nor U23697 (N_23697,N_22495,N_21525);
and U23698 (N_23698,N_21873,N_21734);
or U23699 (N_23699,N_21436,N_22472);
or U23700 (N_23700,N_21648,N_21383);
nand U23701 (N_23701,N_22171,N_22249);
nand U23702 (N_23702,N_21833,N_21430);
nor U23703 (N_23703,N_21434,N_21320);
nor U23704 (N_23704,N_22166,N_22395);
nor U23705 (N_23705,N_21403,N_22105);
nand U23706 (N_23706,N_22217,N_21437);
nand U23707 (N_23707,N_21841,N_22270);
and U23708 (N_23708,N_22432,N_21709);
xnor U23709 (N_23709,N_22290,N_21746);
or U23710 (N_23710,N_21746,N_22163);
or U23711 (N_23711,N_22496,N_22445);
and U23712 (N_23712,N_21664,N_21648);
xor U23713 (N_23713,N_22464,N_22113);
nand U23714 (N_23714,N_22364,N_21668);
or U23715 (N_23715,N_21334,N_21996);
nor U23716 (N_23716,N_21548,N_21259);
nor U23717 (N_23717,N_21647,N_21284);
and U23718 (N_23718,N_22169,N_21876);
and U23719 (N_23719,N_21840,N_21013);
nand U23720 (N_23720,N_21667,N_21697);
nor U23721 (N_23721,N_21424,N_21094);
nand U23722 (N_23722,N_21470,N_21094);
or U23723 (N_23723,N_21932,N_21337);
xnor U23724 (N_23724,N_22423,N_21470);
and U23725 (N_23725,N_22009,N_22049);
or U23726 (N_23726,N_22094,N_21251);
and U23727 (N_23727,N_21708,N_21623);
xor U23728 (N_23728,N_22048,N_22493);
nand U23729 (N_23729,N_21540,N_22436);
or U23730 (N_23730,N_22495,N_22168);
or U23731 (N_23731,N_21654,N_22028);
and U23732 (N_23732,N_21381,N_21614);
and U23733 (N_23733,N_21278,N_22455);
or U23734 (N_23734,N_21357,N_21095);
or U23735 (N_23735,N_21010,N_22050);
or U23736 (N_23736,N_21089,N_21017);
nand U23737 (N_23737,N_22321,N_21091);
nor U23738 (N_23738,N_21701,N_22237);
xor U23739 (N_23739,N_22349,N_21976);
and U23740 (N_23740,N_21761,N_22194);
xor U23741 (N_23741,N_21854,N_22115);
nor U23742 (N_23742,N_21437,N_21483);
nand U23743 (N_23743,N_21943,N_21781);
nor U23744 (N_23744,N_22295,N_22048);
and U23745 (N_23745,N_21695,N_22060);
nand U23746 (N_23746,N_21300,N_21607);
or U23747 (N_23747,N_21447,N_22474);
xor U23748 (N_23748,N_22219,N_21916);
nor U23749 (N_23749,N_21238,N_21440);
and U23750 (N_23750,N_21326,N_22029);
nor U23751 (N_23751,N_21170,N_22444);
or U23752 (N_23752,N_22302,N_22349);
and U23753 (N_23753,N_22254,N_21729);
nor U23754 (N_23754,N_21869,N_21586);
and U23755 (N_23755,N_21071,N_22050);
and U23756 (N_23756,N_22010,N_21031);
and U23757 (N_23757,N_21321,N_21279);
and U23758 (N_23758,N_21206,N_22068);
nor U23759 (N_23759,N_22330,N_21827);
xor U23760 (N_23760,N_21962,N_21307);
or U23761 (N_23761,N_22261,N_21513);
or U23762 (N_23762,N_21737,N_21645);
nand U23763 (N_23763,N_21922,N_21909);
nand U23764 (N_23764,N_21886,N_21299);
nand U23765 (N_23765,N_21787,N_21805);
xnor U23766 (N_23766,N_22167,N_22071);
nor U23767 (N_23767,N_21218,N_21968);
nor U23768 (N_23768,N_21671,N_22224);
and U23769 (N_23769,N_21530,N_21040);
nand U23770 (N_23770,N_21168,N_21692);
or U23771 (N_23771,N_21697,N_22114);
nor U23772 (N_23772,N_21403,N_21644);
nand U23773 (N_23773,N_21128,N_21214);
nand U23774 (N_23774,N_21208,N_21429);
xnor U23775 (N_23775,N_21614,N_21582);
nor U23776 (N_23776,N_22081,N_21182);
nor U23777 (N_23777,N_21352,N_21363);
nand U23778 (N_23778,N_21615,N_22124);
and U23779 (N_23779,N_21523,N_21117);
or U23780 (N_23780,N_22479,N_21210);
and U23781 (N_23781,N_22338,N_21802);
nor U23782 (N_23782,N_22077,N_22146);
or U23783 (N_23783,N_21374,N_22001);
or U23784 (N_23784,N_21021,N_21553);
and U23785 (N_23785,N_21663,N_21341);
and U23786 (N_23786,N_21514,N_21652);
xnor U23787 (N_23787,N_21595,N_21161);
nand U23788 (N_23788,N_21403,N_21278);
xnor U23789 (N_23789,N_21752,N_21497);
nand U23790 (N_23790,N_22025,N_21123);
or U23791 (N_23791,N_21749,N_21444);
nand U23792 (N_23792,N_22076,N_21310);
nor U23793 (N_23793,N_22078,N_21694);
and U23794 (N_23794,N_22351,N_21226);
xor U23795 (N_23795,N_22467,N_22322);
xnor U23796 (N_23796,N_22038,N_21133);
and U23797 (N_23797,N_22138,N_21911);
nand U23798 (N_23798,N_22180,N_21837);
xnor U23799 (N_23799,N_21293,N_22481);
nand U23800 (N_23800,N_21060,N_21639);
nor U23801 (N_23801,N_22133,N_22247);
and U23802 (N_23802,N_21290,N_21019);
nand U23803 (N_23803,N_21648,N_21127);
nand U23804 (N_23804,N_21844,N_21980);
nor U23805 (N_23805,N_21886,N_21432);
nor U23806 (N_23806,N_21567,N_21690);
xnor U23807 (N_23807,N_21250,N_22240);
nor U23808 (N_23808,N_21671,N_21496);
or U23809 (N_23809,N_21092,N_22326);
xnor U23810 (N_23810,N_21544,N_21374);
or U23811 (N_23811,N_21500,N_22170);
or U23812 (N_23812,N_22120,N_21027);
xnor U23813 (N_23813,N_21561,N_21782);
xnor U23814 (N_23814,N_21620,N_21774);
or U23815 (N_23815,N_21625,N_21040);
or U23816 (N_23816,N_22397,N_22041);
or U23817 (N_23817,N_21685,N_22001);
or U23818 (N_23818,N_21495,N_21380);
nor U23819 (N_23819,N_21406,N_21728);
and U23820 (N_23820,N_21071,N_21095);
xor U23821 (N_23821,N_21868,N_21925);
xor U23822 (N_23822,N_21566,N_21544);
nand U23823 (N_23823,N_21216,N_21407);
and U23824 (N_23824,N_21503,N_22063);
nand U23825 (N_23825,N_21502,N_21460);
nand U23826 (N_23826,N_22017,N_22024);
nor U23827 (N_23827,N_21961,N_22452);
or U23828 (N_23828,N_21645,N_21126);
and U23829 (N_23829,N_21728,N_22383);
nor U23830 (N_23830,N_22488,N_21914);
nand U23831 (N_23831,N_21900,N_21384);
and U23832 (N_23832,N_22485,N_22227);
or U23833 (N_23833,N_21575,N_21560);
xor U23834 (N_23834,N_22342,N_22196);
and U23835 (N_23835,N_21953,N_21626);
nor U23836 (N_23836,N_22287,N_22059);
xnor U23837 (N_23837,N_21706,N_21522);
nor U23838 (N_23838,N_22410,N_22042);
or U23839 (N_23839,N_21529,N_21494);
nor U23840 (N_23840,N_22092,N_21988);
or U23841 (N_23841,N_22133,N_22378);
nand U23842 (N_23842,N_21188,N_21980);
nor U23843 (N_23843,N_21339,N_22169);
or U23844 (N_23844,N_21935,N_22449);
nand U23845 (N_23845,N_21408,N_22341);
xor U23846 (N_23846,N_21751,N_21246);
xor U23847 (N_23847,N_21964,N_21191);
xor U23848 (N_23848,N_22462,N_21556);
nor U23849 (N_23849,N_21534,N_21749);
nor U23850 (N_23850,N_22338,N_22438);
nand U23851 (N_23851,N_21691,N_22103);
and U23852 (N_23852,N_21169,N_21443);
nand U23853 (N_23853,N_21498,N_21287);
and U23854 (N_23854,N_22145,N_21894);
or U23855 (N_23855,N_22378,N_21225);
or U23856 (N_23856,N_21499,N_22124);
xor U23857 (N_23857,N_21475,N_22327);
xnor U23858 (N_23858,N_21881,N_21693);
nand U23859 (N_23859,N_21185,N_21226);
or U23860 (N_23860,N_21360,N_21166);
xor U23861 (N_23861,N_22133,N_22358);
and U23862 (N_23862,N_21848,N_22219);
nand U23863 (N_23863,N_22094,N_22282);
and U23864 (N_23864,N_21294,N_21422);
nand U23865 (N_23865,N_22105,N_21874);
or U23866 (N_23866,N_22039,N_21079);
nor U23867 (N_23867,N_22441,N_21986);
or U23868 (N_23868,N_21048,N_22151);
or U23869 (N_23869,N_21803,N_21530);
and U23870 (N_23870,N_22356,N_22017);
nand U23871 (N_23871,N_21161,N_22166);
nand U23872 (N_23872,N_21238,N_22023);
nand U23873 (N_23873,N_21232,N_21272);
and U23874 (N_23874,N_21147,N_21907);
nor U23875 (N_23875,N_21081,N_21761);
nand U23876 (N_23876,N_22352,N_22493);
nand U23877 (N_23877,N_21515,N_21315);
xor U23878 (N_23878,N_21942,N_22472);
xnor U23879 (N_23879,N_22187,N_22403);
xor U23880 (N_23880,N_21641,N_21083);
xor U23881 (N_23881,N_22338,N_21013);
and U23882 (N_23882,N_21154,N_21823);
nand U23883 (N_23883,N_21765,N_21690);
or U23884 (N_23884,N_21510,N_21409);
nor U23885 (N_23885,N_21924,N_22134);
xnor U23886 (N_23886,N_21128,N_21223);
xor U23887 (N_23887,N_21554,N_21654);
nand U23888 (N_23888,N_21178,N_21561);
or U23889 (N_23889,N_21955,N_21234);
and U23890 (N_23890,N_21772,N_22098);
nor U23891 (N_23891,N_21513,N_21435);
xnor U23892 (N_23892,N_21452,N_21708);
xor U23893 (N_23893,N_21788,N_22226);
or U23894 (N_23894,N_22238,N_22486);
and U23895 (N_23895,N_21902,N_21906);
nor U23896 (N_23896,N_22412,N_22279);
nor U23897 (N_23897,N_21182,N_22044);
xnor U23898 (N_23898,N_21284,N_21138);
nand U23899 (N_23899,N_22223,N_22069);
nand U23900 (N_23900,N_21116,N_21480);
and U23901 (N_23901,N_21773,N_21918);
xor U23902 (N_23902,N_21479,N_21990);
nor U23903 (N_23903,N_21001,N_22327);
and U23904 (N_23904,N_21466,N_21317);
nor U23905 (N_23905,N_21178,N_22345);
and U23906 (N_23906,N_21618,N_22326);
xnor U23907 (N_23907,N_21524,N_22285);
and U23908 (N_23908,N_21216,N_21886);
nand U23909 (N_23909,N_21150,N_21719);
or U23910 (N_23910,N_21624,N_21954);
and U23911 (N_23911,N_22269,N_22359);
nand U23912 (N_23912,N_21357,N_21462);
xor U23913 (N_23913,N_22265,N_21537);
nor U23914 (N_23914,N_22199,N_21252);
nand U23915 (N_23915,N_21889,N_21941);
nor U23916 (N_23916,N_22368,N_21265);
and U23917 (N_23917,N_21164,N_21040);
nor U23918 (N_23918,N_21270,N_22217);
nor U23919 (N_23919,N_22355,N_21964);
nor U23920 (N_23920,N_21494,N_21134);
nand U23921 (N_23921,N_22230,N_22424);
and U23922 (N_23922,N_21642,N_22497);
or U23923 (N_23923,N_22161,N_21539);
or U23924 (N_23924,N_21054,N_21969);
nand U23925 (N_23925,N_21201,N_21126);
nand U23926 (N_23926,N_21364,N_21943);
nand U23927 (N_23927,N_21873,N_21206);
or U23928 (N_23928,N_21076,N_22076);
or U23929 (N_23929,N_22034,N_22162);
nand U23930 (N_23930,N_22128,N_21149);
nor U23931 (N_23931,N_22264,N_21234);
and U23932 (N_23932,N_22355,N_22370);
and U23933 (N_23933,N_21569,N_22349);
nand U23934 (N_23934,N_22249,N_21855);
nand U23935 (N_23935,N_21235,N_22277);
nand U23936 (N_23936,N_21667,N_21845);
nor U23937 (N_23937,N_21317,N_21081);
nand U23938 (N_23938,N_21740,N_21504);
xor U23939 (N_23939,N_21424,N_21776);
nor U23940 (N_23940,N_21774,N_21858);
nor U23941 (N_23941,N_21305,N_21989);
or U23942 (N_23942,N_21901,N_21070);
xnor U23943 (N_23943,N_22398,N_21429);
xnor U23944 (N_23944,N_21186,N_22413);
or U23945 (N_23945,N_22381,N_21138);
and U23946 (N_23946,N_21675,N_22412);
xnor U23947 (N_23947,N_21715,N_21205);
and U23948 (N_23948,N_22319,N_21606);
nor U23949 (N_23949,N_21357,N_22085);
nand U23950 (N_23950,N_21290,N_21754);
xor U23951 (N_23951,N_22168,N_22429);
nand U23952 (N_23952,N_22105,N_21357);
nor U23953 (N_23953,N_21775,N_21423);
nor U23954 (N_23954,N_21965,N_21253);
or U23955 (N_23955,N_21252,N_22106);
or U23956 (N_23956,N_21441,N_22113);
nand U23957 (N_23957,N_21435,N_21772);
or U23958 (N_23958,N_22092,N_21513);
and U23959 (N_23959,N_22159,N_21997);
nand U23960 (N_23960,N_21451,N_21930);
nand U23961 (N_23961,N_21331,N_22266);
xor U23962 (N_23962,N_22191,N_21873);
and U23963 (N_23963,N_22259,N_22405);
and U23964 (N_23964,N_21641,N_21283);
xor U23965 (N_23965,N_21093,N_21000);
nand U23966 (N_23966,N_21086,N_21359);
and U23967 (N_23967,N_21827,N_22488);
and U23968 (N_23968,N_22385,N_21053);
xnor U23969 (N_23969,N_22432,N_22359);
nor U23970 (N_23970,N_21161,N_22420);
or U23971 (N_23971,N_21962,N_21041);
xor U23972 (N_23972,N_22430,N_21389);
nor U23973 (N_23973,N_22091,N_22175);
and U23974 (N_23974,N_21635,N_21868);
or U23975 (N_23975,N_21548,N_21434);
nor U23976 (N_23976,N_22301,N_21058);
and U23977 (N_23977,N_22414,N_21260);
or U23978 (N_23978,N_21422,N_22215);
nor U23979 (N_23979,N_22318,N_22268);
or U23980 (N_23980,N_21713,N_21651);
nand U23981 (N_23981,N_22089,N_21838);
and U23982 (N_23982,N_21627,N_21732);
nand U23983 (N_23983,N_22057,N_21861);
and U23984 (N_23984,N_22047,N_22335);
or U23985 (N_23985,N_21714,N_22023);
nor U23986 (N_23986,N_21850,N_21744);
and U23987 (N_23987,N_21747,N_22251);
nor U23988 (N_23988,N_22420,N_21954);
nand U23989 (N_23989,N_22110,N_21041);
and U23990 (N_23990,N_21619,N_22267);
nor U23991 (N_23991,N_22270,N_21747);
nor U23992 (N_23992,N_21689,N_21159);
xor U23993 (N_23993,N_21318,N_22496);
nor U23994 (N_23994,N_21284,N_21362);
nand U23995 (N_23995,N_21932,N_21199);
nand U23996 (N_23996,N_22029,N_21415);
or U23997 (N_23997,N_21029,N_21303);
and U23998 (N_23998,N_22016,N_21790);
xnor U23999 (N_23999,N_21384,N_21211);
and U24000 (N_24000,N_23188,N_22889);
nand U24001 (N_24001,N_23185,N_22568);
and U24002 (N_24002,N_22571,N_23651);
nand U24003 (N_24003,N_22550,N_23194);
and U24004 (N_24004,N_23431,N_23634);
and U24005 (N_24005,N_23725,N_23496);
and U24006 (N_24006,N_22519,N_22749);
nand U24007 (N_24007,N_23518,N_23277);
or U24008 (N_24008,N_23937,N_23543);
nand U24009 (N_24009,N_22986,N_22899);
nor U24010 (N_24010,N_23285,N_23141);
xnor U24011 (N_24011,N_23839,N_23921);
nor U24012 (N_24012,N_23763,N_22837);
nand U24013 (N_24013,N_22699,N_23843);
xor U24014 (N_24014,N_22637,N_23758);
or U24015 (N_24015,N_23583,N_22799);
and U24016 (N_24016,N_23816,N_23177);
and U24017 (N_24017,N_22835,N_22760);
xor U24018 (N_24018,N_23638,N_23125);
or U24019 (N_24019,N_23786,N_22911);
xor U24020 (N_24020,N_23942,N_22654);
nor U24021 (N_24021,N_23525,N_22668);
and U24022 (N_24022,N_22732,N_23392);
or U24023 (N_24023,N_22578,N_23881);
and U24024 (N_24024,N_22703,N_22791);
nor U24025 (N_24025,N_22562,N_23421);
nor U24026 (N_24026,N_23098,N_23293);
nor U24027 (N_24027,N_23913,N_23570);
or U24028 (N_24028,N_22815,N_23642);
nand U24029 (N_24029,N_23924,N_22647);
nand U24030 (N_24030,N_22782,N_23727);
and U24031 (N_24031,N_23626,N_23990);
or U24032 (N_24032,N_23756,N_22591);
xor U24033 (N_24033,N_23814,N_23487);
xnor U24034 (N_24034,N_22962,N_23492);
nand U24035 (N_24035,N_22661,N_23273);
nand U24036 (N_24036,N_23464,N_22956);
and U24037 (N_24037,N_23797,N_23472);
nand U24038 (N_24038,N_23210,N_23710);
xor U24039 (N_24039,N_23289,N_23987);
or U24040 (N_24040,N_22810,N_22579);
nor U24041 (N_24041,N_23984,N_23555);
xor U24042 (N_24042,N_23803,N_23728);
nor U24043 (N_24043,N_23902,N_22722);
nand U24044 (N_24044,N_22786,N_22869);
nand U24045 (N_24045,N_23589,N_23065);
xor U24046 (N_24046,N_22714,N_22763);
nor U24047 (N_24047,N_23844,N_23788);
xnor U24048 (N_24048,N_23478,N_23215);
nor U24049 (N_24049,N_23485,N_23676);
or U24050 (N_24050,N_23977,N_23039);
nand U24051 (N_24051,N_23313,N_23545);
nand U24052 (N_24052,N_23407,N_22857);
nor U24053 (N_24053,N_22942,N_23140);
or U24054 (N_24054,N_23938,N_23052);
nor U24055 (N_24055,N_23375,N_23195);
nor U24056 (N_24056,N_22943,N_22887);
nand U24057 (N_24057,N_23948,N_23677);
nand U24058 (N_24058,N_23418,N_23227);
or U24059 (N_24059,N_23353,N_23197);
or U24060 (N_24060,N_22831,N_22643);
nor U24061 (N_24061,N_23240,N_23712);
xnor U24062 (N_24062,N_22853,N_22950);
nor U24063 (N_24063,N_23877,N_23272);
or U24064 (N_24064,N_23862,N_23494);
or U24065 (N_24065,N_23480,N_23341);
nor U24066 (N_24066,N_23900,N_23701);
nand U24067 (N_24067,N_23323,N_22707);
or U24068 (N_24068,N_23889,N_23696);
nand U24069 (N_24069,N_23654,N_23815);
nand U24070 (N_24070,N_22925,N_23151);
or U24071 (N_24071,N_23196,N_23427);
and U24072 (N_24072,N_23517,N_23688);
nand U24073 (N_24073,N_22616,N_23025);
and U24074 (N_24074,N_23904,N_23908);
nor U24075 (N_24075,N_23069,N_22548);
nor U24076 (N_24076,N_22599,N_23707);
nor U24077 (N_24077,N_22854,N_23952);
or U24078 (N_24078,N_23137,N_23505);
xnor U24079 (N_24079,N_23886,N_23153);
nand U24080 (N_24080,N_22514,N_22987);
nor U24081 (N_24081,N_23829,N_23306);
nor U24082 (N_24082,N_23250,N_23602);
or U24083 (N_24083,N_23001,N_22803);
nor U24084 (N_24084,N_23563,N_23523);
nor U24085 (N_24085,N_22762,N_23493);
xnor U24086 (N_24086,N_23567,N_23876);
and U24087 (N_24087,N_22759,N_23174);
xor U24088 (N_24088,N_23686,N_23930);
xor U24089 (N_24089,N_23777,N_22862);
nand U24090 (N_24090,N_22744,N_23510);
and U24091 (N_24091,N_23871,N_23484);
nand U24092 (N_24092,N_23429,N_23693);
or U24093 (N_24093,N_23733,N_22967);
nor U24094 (N_24094,N_22990,N_23056);
nand U24095 (N_24095,N_22752,N_22560);
nand U24096 (N_24096,N_22503,N_22684);
or U24097 (N_24097,N_23695,N_23507);
and U24098 (N_24098,N_23334,N_22965);
xor U24099 (N_24099,N_23382,N_23622);
nand U24100 (N_24100,N_23000,N_22918);
nor U24101 (N_24101,N_23437,N_23827);
nand U24102 (N_24102,N_23956,N_22634);
and U24103 (N_24103,N_23312,N_23633);
nand U24104 (N_24104,N_23625,N_23818);
and U24105 (N_24105,N_23776,N_22932);
xor U24106 (N_24106,N_22743,N_23524);
nand U24107 (N_24107,N_23536,N_22811);
or U24108 (N_24108,N_23417,N_23586);
and U24109 (N_24109,N_22961,N_23286);
or U24110 (N_24110,N_22745,N_23561);
xnor U24111 (N_24111,N_23389,N_22522);
or U24112 (N_24112,N_23853,N_23859);
nor U24113 (N_24113,N_22711,N_23093);
nor U24114 (N_24114,N_23087,N_22630);
nand U24115 (N_24115,N_22721,N_22690);
nor U24116 (N_24116,N_23176,N_23370);
nor U24117 (N_24117,N_22641,N_23038);
nand U24118 (N_24118,N_23404,N_22608);
xor U24119 (N_24119,N_23996,N_23729);
and U24120 (N_24120,N_23112,N_22597);
nand U24121 (N_24121,N_23340,N_22793);
and U24122 (N_24122,N_22993,N_22806);
and U24123 (N_24123,N_23857,N_23730);
xnor U24124 (N_24124,N_23363,N_22547);
nor U24125 (N_24125,N_23690,N_23079);
xnor U24126 (N_24126,N_22674,N_22555);
and U24127 (N_24127,N_23755,N_23752);
xor U24128 (N_24128,N_23444,N_23754);
nand U24129 (N_24129,N_22895,N_22559);
and U24130 (N_24130,N_23491,N_23806);
xnor U24131 (N_24131,N_23869,N_23648);
and U24132 (N_24132,N_23088,N_22733);
xnor U24133 (N_24133,N_23934,N_23047);
or U24134 (N_24134,N_22681,N_23413);
nor U24135 (N_24135,N_23587,N_23299);
and U24136 (N_24136,N_23894,N_23405);
and U24137 (N_24137,N_22748,N_23978);
and U24138 (N_24138,N_23322,N_23258);
and U24139 (N_24139,N_22800,N_23577);
xnor U24140 (N_24140,N_23106,N_22881);
nor U24141 (N_24141,N_23771,N_22841);
xnor U24142 (N_24142,N_22628,N_22888);
nand U24143 (N_24143,N_23424,N_22808);
or U24144 (N_24144,N_23539,N_22671);
nor U24145 (N_24145,N_22713,N_23330);
and U24146 (N_24146,N_23640,N_23346);
and U24147 (N_24147,N_23706,N_23320);
nor U24148 (N_24148,N_22670,N_23458);
xor U24149 (N_24149,N_23588,N_23476);
and U24150 (N_24150,N_23135,N_23747);
nand U24151 (N_24151,N_23451,N_23506);
and U24152 (N_24152,N_23048,N_23678);
and U24153 (N_24153,N_23211,N_23339);
nor U24154 (N_24154,N_23898,N_23874);
xor U24155 (N_24155,N_22664,N_23782);
nand U24156 (N_24156,N_23373,N_23946);
nand U24157 (N_24157,N_23745,N_23265);
nand U24158 (N_24158,N_22886,N_23888);
or U24159 (N_24159,N_23275,N_22790);
nor U24160 (N_24160,N_23832,N_23049);
nor U24161 (N_24161,N_23007,N_22873);
nor U24162 (N_24162,N_23580,N_23576);
and U24163 (N_24163,N_23593,N_22650);
xor U24164 (N_24164,N_22566,N_23855);
nand U24165 (N_24165,N_23719,N_22700);
nor U24166 (N_24166,N_23138,N_23055);
nand U24167 (N_24167,N_22813,N_22532);
nand U24168 (N_24168,N_22601,N_23830);
and U24169 (N_24169,N_23011,N_22594);
nand U24170 (N_24170,N_23142,N_22586);
or U24171 (N_24171,N_23896,N_23623);
xnor U24172 (N_24172,N_23213,N_23994);
xor U24173 (N_24173,N_22850,N_23632);
nand U24174 (N_24174,N_23915,N_23919);
xor U24175 (N_24175,N_22820,N_23222);
xor U24176 (N_24176,N_23269,N_23344);
nor U24177 (N_24177,N_23027,N_23460);
nand U24178 (N_24178,N_23336,N_23445);
nor U24179 (N_24179,N_23498,N_22516);
nor U24180 (N_24180,N_22880,N_23531);
and U24181 (N_24181,N_22705,N_22504);
nand U24182 (N_24182,N_23294,N_23720);
and U24183 (N_24183,N_23081,N_23973);
nand U24184 (N_24184,N_23226,N_23152);
or U24185 (N_24185,N_23159,N_22600);
nor U24186 (N_24186,N_22890,N_23267);
xor U24187 (N_24187,N_23601,N_23256);
and U24188 (N_24188,N_22912,N_23452);
xnor U24189 (N_24189,N_22777,N_22679);
nor U24190 (N_24190,N_23718,N_23558);
xnor U24191 (N_24191,N_23599,N_22604);
or U24192 (N_24192,N_23129,N_23909);
nand U24193 (N_24193,N_23997,N_23940);
nor U24194 (N_24194,N_23395,N_23109);
and U24195 (N_24195,N_23333,N_22821);
or U24196 (N_24196,N_22917,N_22913);
nand U24197 (N_24197,N_23483,N_22908);
xor U24198 (N_24198,N_23689,N_22875);
nor U24199 (N_24199,N_22794,N_23682);
nor U24200 (N_24200,N_23732,N_22620);
or U24201 (N_24201,N_23050,N_23641);
and U24202 (N_24202,N_23772,N_23958);
nand U24203 (N_24203,N_22994,N_22618);
or U24204 (N_24204,N_22610,N_22855);
nand U24205 (N_24205,N_23063,N_23017);
and U24206 (N_24206,N_23746,N_23652);
and U24207 (N_24207,N_22948,N_23073);
nand U24208 (N_24208,N_23166,N_22682);
xnor U24209 (N_24209,N_22500,N_23590);
nand U24210 (N_24210,N_23804,N_23709);
and U24211 (N_24211,N_23883,N_23402);
xnor U24212 (N_24212,N_23846,N_22904);
nand U24213 (N_24213,N_23530,N_23032);
or U24214 (N_24214,N_22551,N_22509);
xnor U24215 (N_24215,N_23446,N_23840);
nand U24216 (N_24216,N_22901,N_23509);
xnor U24217 (N_24217,N_23110,N_23995);
nand U24218 (N_24218,N_23813,N_23516);
nand U24219 (N_24219,N_23596,N_23559);
or U24220 (N_24220,N_23180,N_23557);
and U24221 (N_24221,N_23271,N_23260);
xor U24222 (N_24222,N_23669,N_22642);
and U24223 (N_24223,N_23443,N_23310);
xor U24224 (N_24224,N_22879,N_23753);
nand U24225 (N_24225,N_22561,N_23121);
or U24226 (N_24226,N_23699,N_23532);
xnor U24227 (N_24227,N_22572,N_23992);
or U24228 (N_24228,N_23597,N_22755);
nand U24229 (N_24229,N_22845,N_23118);
and U24230 (N_24230,N_22718,N_23584);
xor U24231 (N_24231,N_23008,N_23094);
nand U24232 (N_24232,N_22979,N_22867);
nor U24233 (N_24233,N_23108,N_22613);
nor U24234 (N_24234,N_22724,N_22525);
and U24235 (N_24235,N_23671,N_23964);
nor U24236 (N_24236,N_23887,N_22852);
and U24237 (N_24237,N_23820,N_23084);
nor U24238 (N_24238,N_23895,N_22840);
nand U24239 (N_24239,N_22656,N_23158);
and U24240 (N_24240,N_23867,N_23658);
nor U24241 (N_24241,N_23100,N_22667);
nand U24242 (N_24242,N_23014,N_23352);
xor U24243 (N_24243,N_23033,N_22691);
and U24244 (N_24244,N_23960,N_23242);
nand U24245 (N_24245,N_23342,N_23629);
xnor U24246 (N_24246,N_23947,N_22937);
xor U24247 (N_24247,N_23091,N_23348);
and U24248 (N_24248,N_22697,N_23660);
nor U24249 (N_24249,N_22717,N_23343);
and U24250 (N_24250,N_22751,N_23662);
and U24251 (N_24251,N_23740,N_22940);
nor U24252 (N_24252,N_22617,N_23912);
nand U24253 (N_24253,N_23010,N_22902);
and U24254 (N_24254,N_23283,N_22527);
and U24255 (N_24255,N_23082,N_23790);
nand U24256 (N_24256,N_23120,N_22534);
nand U24257 (N_24257,N_22952,N_23086);
nor U24258 (N_24258,N_22982,N_22740);
nand U24259 (N_24259,N_23154,N_23891);
and U24260 (N_24260,N_22891,N_22784);
and U24261 (N_24261,N_23779,N_22685);
nor U24262 (N_24262,N_23274,N_23526);
xnor U24263 (N_24263,N_23655,N_22624);
and U24264 (N_24264,N_22927,N_23991);
or U24265 (N_24265,N_23009,N_23833);
nand U24266 (N_24266,N_23512,N_23369);
nand U24267 (N_24267,N_23624,N_22788);
or U24268 (N_24268,N_22676,N_23611);
or U24269 (N_24269,N_23351,N_23036);
nand U24270 (N_24270,N_23618,N_22557);
or U24271 (N_24271,N_22771,N_23467);
nor U24272 (N_24272,N_23354,N_22539);
or U24273 (N_24273,N_23954,N_22916);
and U24274 (N_24274,N_22645,N_22569);
nand U24275 (N_24275,N_23026,N_23311);
xor U24276 (N_24276,N_23305,N_23550);
or U24277 (N_24277,N_22828,N_23999);
nor U24278 (N_24278,N_22692,N_23600);
nor U24279 (N_24279,N_23714,N_23836);
or U24280 (N_24280,N_22836,N_23778);
and U24281 (N_24281,N_22686,N_22541);
or U24282 (N_24282,N_23982,N_22621);
and U24283 (N_24283,N_23132,N_22866);
nor U24284 (N_24284,N_23656,N_23674);
and U24285 (N_24285,N_23966,N_23594);
nor U24286 (N_24286,N_23278,N_22985);
xnor U24287 (N_24287,N_23917,N_22629);
xor U24288 (N_24288,N_23922,N_23303);
nor U24289 (N_24289,N_23308,N_22672);
xnor U24290 (N_24290,N_23416,N_23479);
and U24291 (N_24291,N_23554,N_23649);
and U24292 (N_24292,N_23528,N_23168);
and U24293 (N_24293,N_22535,N_23681);
xnor U24294 (N_24294,N_23276,N_22930);
or U24295 (N_24295,N_23015,N_22678);
xor U24296 (N_24296,N_23178,N_22801);
or U24297 (N_24297,N_23565,N_23173);
and U24298 (N_24298,N_23762,N_23092);
nand U24299 (N_24299,N_23075,N_22577);
xnor U24300 (N_24300,N_23616,N_23175);
nand U24301 (N_24301,N_23668,N_23372);
or U24302 (N_24302,N_23514,N_23713);
nor U24303 (N_24303,N_23787,N_23998);
nand U24304 (N_24304,N_23233,N_23238);
nand U24305 (N_24305,N_23780,N_23606);
and U24306 (N_24306,N_23513,N_23979);
and U24307 (N_24307,N_22812,N_23608);
or U24308 (N_24308,N_23281,N_23521);
xnor U24309 (N_24309,N_23944,N_22689);
or U24310 (N_24310,N_22896,N_23139);
xor U24311 (N_24311,N_23737,N_23302);
nor U24312 (N_24312,N_23819,N_23077);
xnor U24313 (N_24313,N_23184,N_22919);
nand U24314 (N_24314,N_22998,N_23500);
nand U24315 (N_24315,N_22530,N_23926);
nand U24316 (N_24316,N_23237,N_23414);
xor U24317 (N_24317,N_23214,N_22960);
and U24318 (N_24318,N_23230,N_23556);
and U24319 (N_24319,N_23542,N_22508);
and U24320 (N_24320,N_23918,N_23198);
nand U24321 (N_24321,N_23186,N_23143);
nand U24322 (N_24322,N_23469,N_23735);
or U24323 (N_24323,N_23906,N_22615);
or U24324 (N_24324,N_22770,N_22526);
and U24325 (N_24325,N_22649,N_23287);
xor U24326 (N_24326,N_23663,N_23058);
or U24327 (N_24327,N_23134,N_23865);
nand U24328 (N_24328,N_23468,N_22978);
nand U24329 (N_24329,N_23983,N_22646);
and U24330 (N_24330,N_22658,N_23604);
nand U24331 (N_24331,N_23993,N_22847);
nand U24332 (N_24332,N_22505,N_23204);
xor U24333 (N_24333,N_22719,N_22622);
nand U24334 (N_24334,N_22570,N_23419);
or U24335 (N_24335,N_22623,N_23957);
nor U24336 (N_24336,N_22593,N_23164);
or U24337 (N_24337,N_23868,N_23817);
xor U24338 (N_24338,N_23029,N_22644);
and U24339 (N_24339,N_23962,N_23264);
nor U24340 (N_24340,N_23552,N_23761);
xor U24341 (N_24341,N_23775,N_23808);
nand U24342 (N_24342,N_23060,N_23872);
xnor U24343 (N_24343,N_22580,N_23639);
or U24344 (N_24344,N_23356,N_23717);
xnor U24345 (N_24345,N_22728,N_22709);
xor U24346 (N_24346,N_22710,N_22627);
nand U24347 (N_24347,N_22991,N_22614);
xor U24348 (N_24348,N_23793,N_23935);
or U24349 (N_24349,N_23628,N_23440);
or U24350 (N_24350,N_22783,N_22903);
nand U24351 (N_24351,N_23329,N_22951);
nor U24352 (N_24352,N_23534,N_23850);
xor U24353 (N_24353,N_23792,N_23241);
nand U24354 (N_24354,N_22753,N_23743);
nor U24355 (N_24355,N_22585,N_22727);
nor U24356 (N_24356,N_23384,N_23378);
or U24357 (N_24357,N_23080,N_23163);
nand U24358 (N_24358,N_22772,N_23062);
and U24359 (N_24359,N_22575,N_23548);
nor U24360 (N_24360,N_22941,N_23057);
xor U24361 (N_24361,N_23202,N_23497);
nand U24362 (N_24362,N_23337,N_23428);
nand U24363 (N_24363,N_22934,N_22935);
or U24364 (N_24364,N_23236,N_22553);
xnor U24365 (N_24365,N_22677,N_23268);
and U24366 (N_24366,N_23074,N_22652);
xor U24367 (N_24367,N_23595,N_23635);
nor U24368 (N_24368,N_22859,N_23653);
nand U24369 (N_24369,N_22730,N_23379);
nand U24370 (N_24370,N_23679,N_23905);
and U24371 (N_24371,N_23107,N_22716);
nand U24372 (N_24372,N_23931,N_23711);
nor U24373 (N_24373,N_22830,N_22984);
nor U24374 (N_24374,N_22832,N_22757);
nand U24375 (N_24375,N_23078,N_23335);
and U24376 (N_24376,N_23441,N_23579);
xnor U24377 (N_24377,N_22878,N_22885);
nor U24378 (N_24378,N_22877,N_23436);
nor U24379 (N_24379,N_22531,N_23412);
nor U24380 (N_24380,N_23099,N_23400);
or U24381 (N_24381,N_22523,N_22910);
nor U24382 (N_24382,N_23798,N_23704);
nand U24383 (N_24383,N_22513,N_22660);
or U24384 (N_24384,N_22704,N_22737);
nor U24385 (N_24385,N_22981,N_22779);
or U24386 (N_24386,N_23433,N_22512);
and U24387 (N_24387,N_23396,N_22928);
nor U24388 (N_24388,N_23591,N_23040);
nor U24389 (N_24389,N_23249,N_23376);
nand U24390 (N_24390,N_22795,N_22708);
nand U24391 (N_24391,N_23083,N_23206);
and U24392 (N_24392,N_22839,N_22816);
or U24393 (N_24393,N_23592,N_22706);
nor U24394 (N_24394,N_22818,N_23187);
xor U24395 (N_24395,N_23785,N_23279);
nor U24396 (N_24396,N_23362,N_22576);
nand U24397 (N_24397,N_23609,N_22846);
nor U24398 (N_24398,N_23582,N_23316);
nor U24399 (N_24399,N_22796,N_23051);
or U24400 (N_24400,N_22931,N_23013);
or U24401 (N_24401,N_23116,N_23928);
or U24402 (N_24402,N_23927,N_23899);
nor U24403 (N_24403,N_22590,N_22696);
nor U24404 (N_24404,N_22785,N_22653);
nand U24405 (N_24405,N_23828,N_23324);
or U24406 (N_24406,N_23612,N_23231);
and U24407 (N_24407,N_23224,N_23355);
and U24408 (N_24408,N_22922,N_23630);
nor U24409 (N_24409,N_22675,N_23315);
nor U24410 (N_24410,N_22976,N_22870);
xnor U24411 (N_24411,N_23810,N_22814);
and U24412 (N_24412,N_23466,N_22871);
nand U24413 (N_24413,N_23035,N_23636);
xor U24414 (N_24414,N_22666,N_22524);
nor U24415 (N_24415,N_22804,N_23959);
and U24416 (N_24416,N_22974,N_23541);
or U24417 (N_24417,N_23546,N_23457);
nor U24418 (N_24418,N_23823,N_22972);
and U24419 (N_24419,N_22809,N_23607);
and U24420 (N_24420,N_23255,N_23349);
xor U24421 (N_24421,N_23037,N_23698);
nand U24422 (N_24422,N_22778,N_23482);
and U24423 (N_24423,N_23115,N_23071);
or U24424 (N_24424,N_23162,N_23119);
and U24425 (N_24425,N_23739,N_23368);
and U24426 (N_24426,N_23208,N_23860);
nand U24427 (N_24427,N_23390,N_23085);
xor U24428 (N_24428,N_23410,N_23061);
or U24429 (N_24429,N_22549,N_23005);
nand U24430 (N_24430,N_23200,N_23165);
and U24431 (N_24431,N_22720,N_22537);
or U24432 (N_24432,N_23420,N_23105);
nor U24433 (N_24433,N_23708,N_23095);
xor U24434 (N_24434,N_22723,N_23430);
or U24435 (N_24435,N_23199,N_22874);
nor U24436 (N_24436,N_23246,N_23511);
nor U24437 (N_24437,N_22781,N_23974);
xnor U24438 (N_24438,N_23114,N_23533);
xor U24439 (N_24439,N_23650,N_23884);
nor U24440 (N_24440,N_23923,N_23892);
nor U24441 (N_24441,N_23967,N_23981);
nand U24442 (N_24442,N_23314,N_23873);
and U24443 (N_24443,N_23975,N_22838);
xor U24444 (N_24444,N_23723,N_23189);
or U24445 (N_24445,N_22834,N_23619);
or U24446 (N_24446,N_22533,N_23123);
nor U24447 (N_24447,N_22611,N_23325);
and U24448 (N_24448,N_23789,N_23284);
or U24449 (N_24449,N_23366,N_23985);
nor U24450 (N_24450,N_23220,N_22921);
xor U24451 (N_24451,N_22872,N_23691);
nand U24452 (N_24452,N_22702,N_23435);
nor U24453 (N_24453,N_23462,N_23757);
or U24454 (N_24454,N_22926,N_23705);
nand U24455 (N_24455,N_23796,N_23364);
and U24456 (N_24456,N_23282,N_22829);
or U24457 (N_24457,N_23191,N_23538);
or U24458 (N_24458,N_23673,N_23659);
nor U24459 (N_24459,N_23508,N_22588);
and U24460 (N_24460,N_23434,N_22598);
or U24461 (N_24461,N_22683,N_22635);
or U24462 (N_24462,N_22564,N_23053);
xor U24463 (N_24463,N_23358,N_23615);
and U24464 (N_24464,N_23454,N_22659);
and U24465 (N_24465,N_23614,N_23328);
and U24466 (N_24466,N_23031,N_22955);
nor U24467 (N_24467,N_23784,N_23527);
and U24468 (N_24468,N_23627,N_22989);
nand U24469 (N_24469,N_22750,N_22558);
nor U24470 (N_24470,N_23111,N_22758);
or U24471 (N_24471,N_22583,N_23742);
xnor U24472 (N_24472,N_23826,N_23951);
nor U24473 (N_24473,N_22693,N_23972);
nand U24474 (N_24474,N_23104,N_22606);
and U24475 (N_24475,N_23744,N_23759);
and U24476 (N_24476,N_22520,N_23741);
and U24477 (N_24477,N_23398,N_22968);
nor U24478 (N_24478,N_23799,N_22946);
xor U24479 (N_24479,N_22954,N_23350);
nor U24480 (N_24480,N_23181,N_23549);
and U24481 (N_24481,N_23386,N_23232);
xnor U24482 (N_24482,N_23461,N_22712);
and U24483 (N_24483,N_23644,N_23722);
nor U24484 (N_24484,N_23296,N_22738);
and U24485 (N_24485,N_22736,N_23393);
nor U24486 (N_24486,N_23878,N_23495);
and U24487 (N_24487,N_23183,N_22529);
xnor U24488 (N_24488,N_22544,N_23683);
and U24489 (N_24489,N_23553,N_23374);
nand U24490 (N_24490,N_23387,N_23295);
xnor U24491 (N_24491,N_23687,N_22966);
nor U24492 (N_24492,N_22701,N_23243);
xor U24493 (N_24493,N_23447,N_23502);
or U24494 (N_24494,N_23613,N_23901);
and U24495 (N_24495,N_22900,N_22636);
nor U24496 (N_24496,N_23760,N_23147);
nor U24497 (N_24497,N_23721,N_23551);
nor U24498 (N_24498,N_23903,N_23643);
xor U24499 (N_24499,N_23573,N_23045);
and U24500 (N_24500,N_23298,N_22766);
and U24501 (N_24501,N_23807,N_23945);
nor U24502 (N_24502,N_23968,N_23422);
nand U24503 (N_24503,N_23925,N_23961);
or U24504 (N_24504,N_23515,N_22596);
and U24505 (N_24505,N_23043,N_22742);
or U24506 (N_24506,N_23235,N_23270);
nor U24507 (N_24507,N_23297,N_23939);
nor U24508 (N_24508,N_22780,N_23875);
xnor U24509 (N_24509,N_23637,N_23499);
or U24510 (N_24510,N_23207,N_23598);
nand U24511 (N_24511,N_22545,N_23971);
nor U24512 (N_24512,N_23361,N_23169);
or U24513 (N_24513,N_23453,N_23716);
nor U24514 (N_24514,N_22538,N_22536);
and U24515 (N_24515,N_23851,N_23347);
xnor U24516 (N_24516,N_23501,N_22574);
and U24517 (N_24517,N_22933,N_23835);
nand U24518 (N_24518,N_23423,N_23822);
nor U24519 (N_24519,N_23578,N_23406);
nor U24520 (N_24520,N_22521,N_22639);
nor U24521 (N_24521,N_23380,N_23692);
nor U24522 (N_24522,N_23450,N_23879);
or U24523 (N_24523,N_22848,N_23764);
or U24524 (N_24524,N_22851,N_22980);
nand U24525 (N_24525,N_23090,N_22924);
nand U24526 (N_24526,N_22923,N_23970);
nand U24527 (N_24527,N_23113,N_22655);
nor U24528 (N_24528,N_23471,N_22970);
or U24529 (N_24529,N_23749,N_22929);
xor U24530 (N_24530,N_22631,N_23474);
nand U24531 (N_24531,N_23367,N_22775);
nor U24532 (N_24532,N_22997,N_23473);
nor U24533 (N_24533,N_23617,N_23519);
or U24534 (N_24534,N_23345,N_23253);
nor U24535 (N_24535,N_22849,N_22698);
and U24536 (N_24536,N_23216,N_22543);
or U24537 (N_24537,N_23317,N_23046);
or U24538 (N_24538,N_23127,N_23914);
xor U24539 (N_24539,N_23503,N_23897);
nand U24540 (N_24540,N_23067,N_22953);
nand U24541 (N_24541,N_23149,N_22843);
xor U24542 (N_24542,N_23861,N_22938);
nand U24543 (N_24543,N_23988,N_22626);
nand U24544 (N_24544,N_23963,N_22947);
or U24545 (N_24545,N_23397,N_23321);
nor U24546 (N_24546,N_23694,N_23470);
nor U24547 (N_24547,N_23409,N_22587);
and U24548 (N_24548,N_23024,N_22552);
nor U24549 (N_24549,N_22876,N_22893);
or U24550 (N_24550,N_23566,N_23403);
and U24551 (N_24551,N_23781,N_23529);
nor U24552 (N_24552,N_22633,N_22695);
and U24553 (N_24553,N_23547,N_22819);
or U24554 (N_24554,N_23338,N_22897);
or U24555 (N_24555,N_23304,N_23560);
xnor U24556 (N_24556,N_22964,N_23929);
xor U24557 (N_24557,N_23481,N_22936);
and U24558 (N_24558,N_22663,N_23522);
and U24559 (N_24559,N_23371,N_23203);
and U24560 (N_24560,N_23751,N_23941);
nor U24561 (N_24561,N_23670,N_23574);
xor U24562 (N_24562,N_23750,N_22657);
and U24563 (N_24563,N_22607,N_23748);
nand U24564 (N_24564,N_22735,N_22612);
nand U24565 (N_24565,N_22715,N_22511);
xor U24566 (N_24566,N_22858,N_23535);
xnor U24567 (N_24567,N_22898,N_23911);
or U24568 (N_24568,N_23442,N_23044);
nand U24569 (N_24569,N_22510,N_22973);
or U24570 (N_24570,N_22638,N_22971);
nand U24571 (N_24571,N_23097,N_23234);
and U24572 (N_24572,N_23890,N_22602);
xor U24573 (N_24573,N_23266,N_23581);
and U24574 (N_24574,N_23932,N_22996);
nand U24575 (N_24575,N_23842,N_23802);
nand U24576 (N_24576,N_23059,N_23006);
nand U24577 (N_24577,N_22595,N_23965);
and U24578 (N_24578,N_23920,N_23465);
nor U24579 (N_24579,N_22905,N_23585);
xnor U24580 (N_24580,N_22975,N_23292);
or U24581 (N_24581,N_23170,N_22662);
nand U24582 (N_24582,N_23791,N_23205);
or U24583 (N_24583,N_23300,N_23425);
or U24584 (N_24584,N_23620,N_23540);
xnor U24585 (N_24585,N_23805,N_23936);
xnor U24586 (N_24586,N_23193,N_22909);
nor U24587 (N_24587,N_23016,N_23076);
xnor U24588 (N_24588,N_23858,N_23018);
or U24589 (N_24589,N_23225,N_22865);
nand U24590 (N_24590,N_22603,N_22817);
or U24591 (N_24591,N_23675,N_23774);
xor U24592 (N_24592,N_23021,N_22864);
nand U24593 (N_24593,N_23212,N_23223);
nand U24594 (N_24594,N_23773,N_23172);
or U24595 (N_24595,N_22827,N_23724);
or U24596 (N_24596,N_23391,N_22999);
xnor U24597 (N_24597,N_22860,N_23319);
xnor U24598 (N_24598,N_22825,N_23767);
and U24599 (N_24599,N_22741,N_22949);
xor U24600 (N_24600,N_22694,N_23318);
and U24601 (N_24601,N_22725,N_22563);
nor U24602 (N_24602,N_23603,N_22944);
nand U24603 (N_24603,N_23800,N_23809);
nor U24604 (N_24604,N_23103,N_23280);
nand U24605 (N_24605,N_23101,N_23003);
nand U24606 (N_24606,N_23537,N_22995);
or U24607 (N_24607,N_23488,N_22826);
or U24608 (N_24608,N_22507,N_22833);
and U24609 (N_24609,N_23989,N_23845);
and U24610 (N_24610,N_22992,N_23201);
and U24611 (N_24611,N_23426,N_23955);
and U24612 (N_24612,N_23157,N_23432);
xnor U24613 (N_24613,N_23811,N_23089);
nor U24614 (N_24614,N_23852,N_23459);
or U24615 (N_24615,N_23102,N_23054);
or U24616 (N_24616,N_23893,N_22625);
xor U24617 (N_24617,N_23122,N_23179);
nand U24618 (N_24618,N_23834,N_22673);
xnor U24619 (N_24619,N_23449,N_22573);
xor U24620 (N_24620,N_23332,N_23765);
xor U24621 (N_24621,N_22518,N_23217);
and U24622 (N_24622,N_22842,N_23980);
nand U24623 (N_24623,N_23475,N_22747);
and U24624 (N_24624,N_22983,N_23863);
nor U24625 (N_24625,N_22605,N_22807);
nor U24626 (N_24626,N_23680,N_22945);
or U24627 (N_24627,N_22767,N_23672);
and U24628 (N_24628,N_23288,N_22517);
nand U24629 (N_24629,N_23219,N_23070);
and U24630 (N_24630,N_23953,N_23976);
and U24631 (N_24631,N_23801,N_23824);
or U24632 (N_24632,N_23463,N_23455);
or U24633 (N_24633,N_22632,N_23504);
nor U24634 (N_24634,N_23794,N_23130);
xnor U24635 (N_24635,N_23986,N_23259);
nor U24636 (N_24636,N_22768,N_23568);
xnor U24637 (N_24637,N_23700,N_23882);
xor U24638 (N_24638,N_23126,N_22756);
nand U24639 (N_24639,N_23262,N_23731);
nand U24640 (N_24640,N_22787,N_22687);
and U24641 (N_24641,N_22805,N_23161);
nand U24642 (N_24642,N_22546,N_22764);
or U24643 (N_24643,N_23381,N_22688);
nor U24644 (N_24644,N_23360,N_22823);
and U24645 (N_24645,N_22977,N_22761);
xnor U24646 (N_24646,N_22501,N_22969);
xnor U24647 (N_24647,N_23950,N_23610);
xnor U24648 (N_24648,N_22565,N_23697);
nand U24649 (N_24649,N_23438,N_23252);
xor U24650 (N_24650,N_23096,N_22883);
nand U24651 (N_24651,N_23020,N_22609);
xor U24652 (N_24652,N_23171,N_23192);
nor U24653 (N_24653,N_23002,N_23066);
and U24654 (N_24654,N_23664,N_23969);
nor U24655 (N_24655,N_22856,N_23880);
nor U24656 (N_24656,N_22540,N_23385);
nor U24657 (N_24657,N_22906,N_22959);
or U24658 (N_24658,N_23770,N_23661);
and U24659 (N_24659,N_23562,N_23667);
or U24660 (N_24660,N_23685,N_23327);
or U24661 (N_24661,N_23703,N_23209);
xnor U24662 (N_24662,N_23257,N_23854);
xor U24663 (N_24663,N_22665,N_22957);
nor U24664 (N_24664,N_23408,N_23736);
nor U24665 (N_24665,N_23702,N_22915);
or U24666 (N_24666,N_22776,N_22963);
nand U24667 (N_24667,N_23190,N_22515);
and U24668 (N_24668,N_22769,N_23155);
nand U24669 (N_24669,N_23448,N_23144);
xor U24670 (N_24670,N_22582,N_23133);
nand U24671 (N_24671,N_23156,N_22797);
and U24672 (N_24672,N_23377,N_23856);
nand U24673 (N_24673,N_23621,N_23064);
nand U24674 (N_24674,N_23022,N_23572);
and U24675 (N_24675,N_23028,N_22939);
and U24676 (N_24676,N_22861,N_23657);
nand U24677 (N_24677,N_23124,N_23247);
nor U24678 (N_24678,N_23251,N_23150);
nor U24679 (N_24679,N_22892,N_23821);
nand U24680 (N_24680,N_23738,N_22746);
or U24681 (N_24681,N_23486,N_23004);
nor U24682 (N_24682,N_22792,N_22581);
xnor U24683 (N_24683,N_23837,N_23254);
and U24684 (N_24684,N_23575,N_23715);
or U24685 (N_24685,N_23907,N_23864);
xor U24686 (N_24686,N_23290,N_22754);
nand U24687 (N_24687,N_23182,N_23012);
xor U24688 (N_24688,N_23943,N_23795);
or U24689 (N_24689,N_23866,N_23019);
nor U24690 (N_24690,N_22863,N_23030);
xnor U24691 (N_24691,N_23666,N_23221);
nand U24692 (N_24692,N_23229,N_23383);
or U24693 (N_24693,N_22669,N_23415);
nor U24694 (N_24694,N_23477,N_22542);
or U24695 (N_24695,N_22894,N_23041);
xnor U24696 (N_24696,N_22648,N_22824);
nand U24697 (N_24697,N_23228,N_23148);
and U24698 (N_24698,N_23136,N_23847);
or U24699 (N_24699,N_22844,N_23783);
and U24700 (N_24700,N_22554,N_23665);
and U24701 (N_24701,N_23849,N_23394);
nor U24702 (N_24702,N_22739,N_22765);
xnor U24703 (N_24703,N_23301,N_22822);
xnor U24704 (N_24704,N_23734,N_22567);
nand U24705 (N_24705,N_23248,N_23042);
nand U24706 (N_24706,N_23359,N_22619);
nor U24707 (N_24707,N_23769,N_23439);
xnor U24708 (N_24708,N_22774,N_23218);
xor U24709 (N_24709,N_23239,N_23331);
nor U24710 (N_24710,N_23146,N_23933);
xnor U24711 (N_24711,N_23131,N_23401);
xnor U24712 (N_24712,N_23489,N_23726);
xor U24713 (N_24713,N_23831,N_23309);
xor U24714 (N_24714,N_22773,N_23068);
nand U24715 (N_24715,N_23160,N_23645);
nand U24716 (N_24716,N_23631,N_23848);
nand U24717 (N_24717,N_22680,N_22798);
nor U24718 (N_24718,N_23838,N_22506);
nor U24719 (N_24719,N_23569,N_22651);
xnor U24720 (N_24720,N_23841,N_23365);
nand U24721 (N_24721,N_23910,N_23605);
and U24722 (N_24722,N_23023,N_22592);
xnor U24723 (N_24723,N_23261,N_22988);
or U24724 (N_24724,N_23684,N_23167);
or U24725 (N_24725,N_23357,N_22726);
xor U24726 (N_24726,N_23490,N_22556);
nand U24727 (N_24727,N_22528,N_23117);
xnor U24728 (N_24728,N_22914,N_22734);
nand U24729 (N_24729,N_22920,N_22882);
and U24730 (N_24730,N_22789,N_23291);
nor U24731 (N_24731,N_23564,N_23646);
nor U24732 (N_24732,N_23411,N_22584);
or U24733 (N_24733,N_22907,N_23768);
xnor U24734 (N_24734,N_22868,N_23949);
or U24735 (N_24735,N_23520,N_22729);
or U24736 (N_24736,N_23128,N_22802);
nand U24737 (N_24737,N_23034,N_23244);
and U24738 (N_24738,N_23388,N_23456);
and U24739 (N_24739,N_22958,N_23647);
or U24740 (N_24740,N_23544,N_23245);
nand U24741 (N_24741,N_23885,N_23145);
and U24742 (N_24742,N_23399,N_23916);
nand U24743 (N_24743,N_23326,N_23072);
xnor U24744 (N_24744,N_22640,N_23766);
nand U24745 (N_24745,N_23870,N_22589);
and U24746 (N_24746,N_23307,N_22731);
nand U24747 (N_24747,N_23825,N_22884);
and U24748 (N_24748,N_23571,N_23263);
xnor U24749 (N_24749,N_23812,N_22502);
or U24750 (N_24750,N_23943,N_22564);
or U24751 (N_24751,N_22982,N_23012);
nor U24752 (N_24752,N_23175,N_23679);
nand U24753 (N_24753,N_22753,N_23781);
or U24754 (N_24754,N_23495,N_23967);
and U24755 (N_24755,N_23167,N_23436);
nand U24756 (N_24756,N_22913,N_23830);
and U24757 (N_24757,N_22520,N_22566);
and U24758 (N_24758,N_23189,N_23948);
or U24759 (N_24759,N_23046,N_23660);
nor U24760 (N_24760,N_23010,N_23868);
xor U24761 (N_24761,N_23654,N_22629);
or U24762 (N_24762,N_23948,N_23454);
or U24763 (N_24763,N_22663,N_23424);
or U24764 (N_24764,N_23055,N_23620);
nand U24765 (N_24765,N_23254,N_22993);
or U24766 (N_24766,N_23569,N_23346);
xnor U24767 (N_24767,N_23243,N_22574);
nand U24768 (N_24768,N_23958,N_23093);
xor U24769 (N_24769,N_22737,N_22801);
nand U24770 (N_24770,N_22838,N_22710);
and U24771 (N_24771,N_23226,N_23701);
and U24772 (N_24772,N_23943,N_23771);
or U24773 (N_24773,N_23080,N_22600);
nand U24774 (N_24774,N_22598,N_22665);
and U24775 (N_24775,N_22633,N_23483);
xor U24776 (N_24776,N_23519,N_22860);
or U24777 (N_24777,N_22807,N_23034);
xnor U24778 (N_24778,N_23243,N_23755);
nor U24779 (N_24779,N_23944,N_22597);
nand U24780 (N_24780,N_23086,N_23739);
and U24781 (N_24781,N_23093,N_23997);
or U24782 (N_24782,N_23190,N_22755);
xnor U24783 (N_24783,N_23340,N_23687);
and U24784 (N_24784,N_23680,N_22992);
xnor U24785 (N_24785,N_23544,N_23832);
xnor U24786 (N_24786,N_23511,N_23974);
xor U24787 (N_24787,N_23090,N_22705);
or U24788 (N_24788,N_23043,N_23291);
nor U24789 (N_24789,N_23619,N_23955);
xnor U24790 (N_24790,N_22905,N_23057);
xor U24791 (N_24791,N_23882,N_22642);
nor U24792 (N_24792,N_23445,N_22859);
nand U24793 (N_24793,N_22699,N_23748);
xnor U24794 (N_24794,N_23054,N_22877);
or U24795 (N_24795,N_23776,N_22648);
nand U24796 (N_24796,N_22660,N_22881);
nor U24797 (N_24797,N_22561,N_22862);
or U24798 (N_24798,N_23920,N_22533);
or U24799 (N_24799,N_23818,N_23391);
xnor U24800 (N_24800,N_22783,N_22795);
nor U24801 (N_24801,N_22833,N_23546);
nand U24802 (N_24802,N_23874,N_22851);
xor U24803 (N_24803,N_22941,N_22670);
xnor U24804 (N_24804,N_23753,N_23411);
nor U24805 (N_24805,N_22724,N_23556);
nor U24806 (N_24806,N_22554,N_23660);
nor U24807 (N_24807,N_23501,N_23202);
and U24808 (N_24808,N_22719,N_23556);
nor U24809 (N_24809,N_22630,N_22701);
or U24810 (N_24810,N_23128,N_23319);
and U24811 (N_24811,N_23750,N_23124);
nor U24812 (N_24812,N_23204,N_23176);
nor U24813 (N_24813,N_23336,N_23166);
and U24814 (N_24814,N_23421,N_23642);
or U24815 (N_24815,N_22831,N_23193);
or U24816 (N_24816,N_23251,N_23382);
nor U24817 (N_24817,N_22512,N_22729);
xor U24818 (N_24818,N_23238,N_22645);
or U24819 (N_24819,N_22735,N_23484);
nand U24820 (N_24820,N_23654,N_23401);
or U24821 (N_24821,N_23256,N_23695);
and U24822 (N_24822,N_23421,N_23186);
nand U24823 (N_24823,N_23977,N_22638);
nand U24824 (N_24824,N_23323,N_22999);
nand U24825 (N_24825,N_23451,N_22895);
and U24826 (N_24826,N_22818,N_22755);
nand U24827 (N_24827,N_23926,N_23315);
xnor U24828 (N_24828,N_23900,N_23619);
nand U24829 (N_24829,N_23523,N_23188);
and U24830 (N_24830,N_23693,N_22919);
nor U24831 (N_24831,N_22954,N_23182);
and U24832 (N_24832,N_23440,N_22746);
nor U24833 (N_24833,N_23293,N_22818);
or U24834 (N_24834,N_23438,N_23180);
and U24835 (N_24835,N_23478,N_23064);
nor U24836 (N_24836,N_23625,N_22652);
and U24837 (N_24837,N_23634,N_22773);
xnor U24838 (N_24838,N_22728,N_23863);
nand U24839 (N_24839,N_23261,N_23484);
nor U24840 (N_24840,N_23278,N_23304);
and U24841 (N_24841,N_23364,N_23522);
and U24842 (N_24842,N_23786,N_23587);
nand U24843 (N_24843,N_23247,N_23286);
xnor U24844 (N_24844,N_22725,N_23961);
or U24845 (N_24845,N_23084,N_22988);
nor U24846 (N_24846,N_23377,N_23518);
nand U24847 (N_24847,N_23363,N_23406);
nand U24848 (N_24848,N_23868,N_23379);
and U24849 (N_24849,N_23959,N_23093);
and U24850 (N_24850,N_23385,N_22932);
nand U24851 (N_24851,N_22789,N_23785);
xor U24852 (N_24852,N_23593,N_22504);
and U24853 (N_24853,N_22523,N_23700);
and U24854 (N_24854,N_22620,N_23675);
nand U24855 (N_24855,N_23627,N_23149);
xor U24856 (N_24856,N_22835,N_22941);
nor U24857 (N_24857,N_23123,N_23413);
nand U24858 (N_24858,N_23658,N_23064);
and U24859 (N_24859,N_23686,N_23862);
or U24860 (N_24860,N_23821,N_23008);
or U24861 (N_24861,N_23501,N_23773);
or U24862 (N_24862,N_23652,N_22531);
nor U24863 (N_24863,N_23012,N_22569);
xnor U24864 (N_24864,N_23884,N_23147);
nand U24865 (N_24865,N_22629,N_23729);
or U24866 (N_24866,N_23761,N_23250);
nand U24867 (N_24867,N_22694,N_23128);
nor U24868 (N_24868,N_22796,N_23309);
nor U24869 (N_24869,N_23382,N_23359);
xor U24870 (N_24870,N_22637,N_22757);
nand U24871 (N_24871,N_23191,N_22882);
or U24872 (N_24872,N_23727,N_22646);
nand U24873 (N_24873,N_23771,N_23774);
xnor U24874 (N_24874,N_22846,N_23604);
xor U24875 (N_24875,N_23594,N_23141);
nor U24876 (N_24876,N_22553,N_23100);
and U24877 (N_24877,N_23237,N_23069);
or U24878 (N_24878,N_23885,N_23262);
or U24879 (N_24879,N_22577,N_22560);
nor U24880 (N_24880,N_23010,N_23906);
nand U24881 (N_24881,N_23223,N_23391);
xor U24882 (N_24882,N_22683,N_23663);
xnor U24883 (N_24883,N_23957,N_23870);
and U24884 (N_24884,N_23871,N_22658);
nor U24885 (N_24885,N_23009,N_22820);
nor U24886 (N_24886,N_23386,N_23415);
xnor U24887 (N_24887,N_23591,N_23005);
or U24888 (N_24888,N_23091,N_23594);
and U24889 (N_24889,N_23920,N_23600);
nand U24890 (N_24890,N_22500,N_23467);
or U24891 (N_24891,N_22501,N_23647);
nor U24892 (N_24892,N_22543,N_23546);
nand U24893 (N_24893,N_22858,N_23081);
or U24894 (N_24894,N_23084,N_23294);
nand U24895 (N_24895,N_23128,N_23059);
and U24896 (N_24896,N_23253,N_22529);
or U24897 (N_24897,N_22513,N_22692);
nand U24898 (N_24898,N_23399,N_22971);
nand U24899 (N_24899,N_22933,N_23132);
or U24900 (N_24900,N_23441,N_23717);
and U24901 (N_24901,N_22596,N_23551);
nor U24902 (N_24902,N_23091,N_23285);
nand U24903 (N_24903,N_23274,N_23072);
nor U24904 (N_24904,N_22538,N_22562);
nand U24905 (N_24905,N_23181,N_23335);
nor U24906 (N_24906,N_23092,N_23191);
nor U24907 (N_24907,N_23331,N_23406);
or U24908 (N_24908,N_23469,N_23086);
or U24909 (N_24909,N_22668,N_23667);
nor U24910 (N_24910,N_23027,N_22506);
nand U24911 (N_24911,N_23561,N_23650);
nand U24912 (N_24912,N_23279,N_23036);
and U24913 (N_24913,N_22847,N_23655);
xor U24914 (N_24914,N_22897,N_23898);
nand U24915 (N_24915,N_23302,N_23553);
xnor U24916 (N_24916,N_23420,N_23894);
nor U24917 (N_24917,N_22876,N_22582);
and U24918 (N_24918,N_23537,N_23016);
and U24919 (N_24919,N_23618,N_22521);
nand U24920 (N_24920,N_23028,N_22808);
or U24921 (N_24921,N_23738,N_23481);
xnor U24922 (N_24922,N_23969,N_22878);
xor U24923 (N_24923,N_23330,N_23501);
nor U24924 (N_24924,N_23304,N_23200);
nand U24925 (N_24925,N_23251,N_23330);
nand U24926 (N_24926,N_22996,N_22960);
or U24927 (N_24927,N_23083,N_23568);
nand U24928 (N_24928,N_23573,N_22699);
xor U24929 (N_24929,N_23165,N_23148);
and U24930 (N_24930,N_23136,N_22696);
nand U24931 (N_24931,N_23640,N_23730);
xnor U24932 (N_24932,N_23692,N_23654);
and U24933 (N_24933,N_22937,N_22827);
nor U24934 (N_24934,N_23859,N_23647);
xnor U24935 (N_24935,N_23915,N_23567);
nand U24936 (N_24936,N_23825,N_23705);
nand U24937 (N_24937,N_22701,N_22827);
or U24938 (N_24938,N_23113,N_22684);
and U24939 (N_24939,N_23038,N_23445);
and U24940 (N_24940,N_23043,N_22540);
or U24941 (N_24941,N_23618,N_23227);
nand U24942 (N_24942,N_22787,N_23599);
nor U24943 (N_24943,N_23411,N_22826);
nor U24944 (N_24944,N_23095,N_23103);
nand U24945 (N_24945,N_23353,N_23662);
and U24946 (N_24946,N_23665,N_22594);
nand U24947 (N_24947,N_22837,N_23609);
nor U24948 (N_24948,N_22985,N_23223);
xnor U24949 (N_24949,N_22625,N_22556);
nand U24950 (N_24950,N_23436,N_23281);
or U24951 (N_24951,N_23726,N_23103);
and U24952 (N_24952,N_23914,N_22539);
or U24953 (N_24953,N_23518,N_23527);
xnor U24954 (N_24954,N_23080,N_23409);
or U24955 (N_24955,N_23697,N_23943);
nor U24956 (N_24956,N_23009,N_23702);
or U24957 (N_24957,N_23748,N_23726);
nand U24958 (N_24958,N_23058,N_23738);
xor U24959 (N_24959,N_23656,N_22804);
or U24960 (N_24960,N_23293,N_23511);
nand U24961 (N_24961,N_23001,N_23891);
nor U24962 (N_24962,N_23207,N_23351);
xor U24963 (N_24963,N_22877,N_23501);
or U24964 (N_24964,N_23754,N_22512);
nor U24965 (N_24965,N_22920,N_23134);
and U24966 (N_24966,N_22703,N_22999);
or U24967 (N_24967,N_23179,N_22705);
or U24968 (N_24968,N_22990,N_23819);
nor U24969 (N_24969,N_23579,N_23569);
and U24970 (N_24970,N_22771,N_22701);
or U24971 (N_24971,N_23384,N_23574);
and U24972 (N_24972,N_22920,N_23672);
or U24973 (N_24973,N_22670,N_22748);
xnor U24974 (N_24974,N_23813,N_23953);
nor U24975 (N_24975,N_22560,N_22952);
nor U24976 (N_24976,N_22777,N_22948);
nor U24977 (N_24977,N_23174,N_22585);
xnor U24978 (N_24978,N_22705,N_23143);
nor U24979 (N_24979,N_23995,N_22848);
xnor U24980 (N_24980,N_22544,N_23774);
and U24981 (N_24981,N_22828,N_23268);
or U24982 (N_24982,N_23871,N_22944);
or U24983 (N_24983,N_22839,N_23951);
and U24984 (N_24984,N_22787,N_23043);
and U24985 (N_24985,N_22648,N_23145);
and U24986 (N_24986,N_23215,N_23261);
nor U24987 (N_24987,N_22787,N_22864);
nand U24988 (N_24988,N_23979,N_22544);
and U24989 (N_24989,N_23527,N_23912);
xnor U24990 (N_24990,N_23131,N_23846);
and U24991 (N_24991,N_22729,N_22583);
nor U24992 (N_24992,N_22987,N_23161);
and U24993 (N_24993,N_22836,N_23504);
nand U24994 (N_24994,N_22896,N_22750);
and U24995 (N_24995,N_23184,N_22628);
or U24996 (N_24996,N_22638,N_23551);
and U24997 (N_24997,N_22946,N_23089);
nand U24998 (N_24998,N_23666,N_23116);
nor U24999 (N_24999,N_22670,N_22855);
and U25000 (N_25000,N_23506,N_22784);
nor U25001 (N_25001,N_22550,N_23453);
xnor U25002 (N_25002,N_23720,N_23062);
nand U25003 (N_25003,N_22869,N_22882);
nand U25004 (N_25004,N_23188,N_23409);
nand U25005 (N_25005,N_23198,N_22628);
nand U25006 (N_25006,N_23999,N_22883);
xor U25007 (N_25007,N_22525,N_23879);
xor U25008 (N_25008,N_22637,N_22996);
and U25009 (N_25009,N_23993,N_23424);
and U25010 (N_25010,N_22534,N_22585);
nand U25011 (N_25011,N_23046,N_23301);
and U25012 (N_25012,N_23293,N_23046);
xnor U25013 (N_25013,N_22864,N_23965);
or U25014 (N_25014,N_22957,N_22590);
nor U25015 (N_25015,N_23598,N_23035);
or U25016 (N_25016,N_23720,N_23403);
and U25017 (N_25017,N_23569,N_23884);
and U25018 (N_25018,N_22594,N_23455);
nor U25019 (N_25019,N_23493,N_23450);
xor U25020 (N_25020,N_23913,N_23731);
xor U25021 (N_25021,N_23485,N_22636);
or U25022 (N_25022,N_23780,N_23031);
xnor U25023 (N_25023,N_22770,N_23343);
or U25024 (N_25024,N_23485,N_23603);
and U25025 (N_25025,N_23666,N_23473);
nor U25026 (N_25026,N_23249,N_23407);
xor U25027 (N_25027,N_22691,N_23871);
or U25028 (N_25028,N_22795,N_23316);
or U25029 (N_25029,N_23242,N_23411);
and U25030 (N_25030,N_23254,N_23030);
and U25031 (N_25031,N_23895,N_23964);
nand U25032 (N_25032,N_23004,N_23505);
nor U25033 (N_25033,N_22885,N_23078);
nand U25034 (N_25034,N_22763,N_23383);
or U25035 (N_25035,N_23659,N_23188);
and U25036 (N_25036,N_22896,N_23397);
nand U25037 (N_25037,N_23562,N_23731);
nand U25038 (N_25038,N_23329,N_23264);
nor U25039 (N_25039,N_23118,N_23392);
xnor U25040 (N_25040,N_22624,N_23870);
nor U25041 (N_25041,N_23830,N_23442);
xnor U25042 (N_25042,N_22872,N_23022);
xor U25043 (N_25043,N_23089,N_23785);
xnor U25044 (N_25044,N_23948,N_23778);
xor U25045 (N_25045,N_22921,N_22852);
nand U25046 (N_25046,N_23345,N_22531);
and U25047 (N_25047,N_22883,N_23691);
nor U25048 (N_25048,N_23478,N_22801);
nand U25049 (N_25049,N_22921,N_23994);
and U25050 (N_25050,N_22767,N_22949);
and U25051 (N_25051,N_22646,N_22832);
nor U25052 (N_25052,N_23673,N_22522);
nand U25053 (N_25053,N_23695,N_22675);
nand U25054 (N_25054,N_23852,N_23235);
and U25055 (N_25055,N_23482,N_23687);
nand U25056 (N_25056,N_23426,N_22672);
nand U25057 (N_25057,N_22756,N_23185);
nand U25058 (N_25058,N_23127,N_23762);
xnor U25059 (N_25059,N_23633,N_22770);
and U25060 (N_25060,N_23602,N_23044);
xor U25061 (N_25061,N_22549,N_23654);
nand U25062 (N_25062,N_22887,N_23697);
xnor U25063 (N_25063,N_23735,N_23353);
and U25064 (N_25064,N_22626,N_23089);
xor U25065 (N_25065,N_23863,N_22605);
nor U25066 (N_25066,N_23999,N_23341);
nand U25067 (N_25067,N_23695,N_23146);
nor U25068 (N_25068,N_23413,N_22980);
nand U25069 (N_25069,N_23967,N_23758);
xnor U25070 (N_25070,N_23461,N_22683);
nor U25071 (N_25071,N_23458,N_23557);
nor U25072 (N_25072,N_23349,N_23478);
xnor U25073 (N_25073,N_22985,N_23023);
nor U25074 (N_25074,N_23651,N_22585);
or U25075 (N_25075,N_23050,N_22831);
and U25076 (N_25076,N_23062,N_23573);
and U25077 (N_25077,N_23759,N_23895);
and U25078 (N_25078,N_23659,N_22714);
nand U25079 (N_25079,N_23767,N_23242);
and U25080 (N_25080,N_23970,N_22778);
xnor U25081 (N_25081,N_23336,N_23274);
nand U25082 (N_25082,N_23294,N_22731);
nor U25083 (N_25083,N_22532,N_22683);
nand U25084 (N_25084,N_22994,N_23778);
nand U25085 (N_25085,N_23045,N_23231);
nor U25086 (N_25086,N_23925,N_23811);
nor U25087 (N_25087,N_23750,N_23777);
nand U25088 (N_25088,N_23482,N_23386);
and U25089 (N_25089,N_22722,N_23285);
and U25090 (N_25090,N_23374,N_23464);
xor U25091 (N_25091,N_23393,N_23909);
xor U25092 (N_25092,N_23423,N_23019);
nor U25093 (N_25093,N_22667,N_22585);
and U25094 (N_25094,N_23543,N_22539);
nand U25095 (N_25095,N_23632,N_23705);
nand U25096 (N_25096,N_23575,N_22718);
nor U25097 (N_25097,N_23408,N_22719);
nand U25098 (N_25098,N_23155,N_23765);
and U25099 (N_25099,N_22538,N_23869);
nand U25100 (N_25100,N_22583,N_23248);
and U25101 (N_25101,N_23576,N_22746);
nand U25102 (N_25102,N_22653,N_23330);
and U25103 (N_25103,N_23913,N_23961);
and U25104 (N_25104,N_22803,N_23186);
nand U25105 (N_25105,N_23928,N_23591);
nand U25106 (N_25106,N_23320,N_23492);
nand U25107 (N_25107,N_23095,N_23577);
nand U25108 (N_25108,N_22569,N_23358);
xnor U25109 (N_25109,N_22928,N_23293);
nor U25110 (N_25110,N_23231,N_23184);
nand U25111 (N_25111,N_22607,N_22996);
xor U25112 (N_25112,N_22645,N_23720);
xor U25113 (N_25113,N_22769,N_23356);
xnor U25114 (N_25114,N_23685,N_23126);
nand U25115 (N_25115,N_23109,N_22783);
nand U25116 (N_25116,N_23203,N_23706);
xnor U25117 (N_25117,N_23109,N_22911);
and U25118 (N_25118,N_23722,N_23797);
nor U25119 (N_25119,N_23826,N_22931);
nor U25120 (N_25120,N_23554,N_23640);
nor U25121 (N_25121,N_22654,N_22624);
and U25122 (N_25122,N_22951,N_22679);
nor U25123 (N_25123,N_23417,N_22627);
xor U25124 (N_25124,N_23801,N_22827);
nand U25125 (N_25125,N_23777,N_22955);
and U25126 (N_25126,N_23103,N_23249);
nand U25127 (N_25127,N_23286,N_23201);
xnor U25128 (N_25128,N_22946,N_23438);
nor U25129 (N_25129,N_22790,N_22783);
nor U25130 (N_25130,N_22695,N_22855);
xor U25131 (N_25131,N_22757,N_23069);
or U25132 (N_25132,N_23998,N_22516);
nand U25133 (N_25133,N_22579,N_23729);
or U25134 (N_25134,N_23224,N_22967);
xnor U25135 (N_25135,N_23987,N_23228);
nand U25136 (N_25136,N_22527,N_22628);
nand U25137 (N_25137,N_23519,N_23207);
nor U25138 (N_25138,N_22943,N_22870);
nor U25139 (N_25139,N_23486,N_22989);
and U25140 (N_25140,N_23135,N_22518);
xnor U25141 (N_25141,N_22887,N_22989);
xor U25142 (N_25142,N_22802,N_23897);
or U25143 (N_25143,N_23322,N_23937);
nor U25144 (N_25144,N_23696,N_22744);
nand U25145 (N_25145,N_23731,N_22995);
nand U25146 (N_25146,N_22645,N_23968);
and U25147 (N_25147,N_22787,N_23065);
or U25148 (N_25148,N_23768,N_23718);
xor U25149 (N_25149,N_23800,N_22948);
and U25150 (N_25150,N_22878,N_23026);
or U25151 (N_25151,N_23134,N_22861);
xor U25152 (N_25152,N_23876,N_23504);
xnor U25153 (N_25153,N_22979,N_23120);
nor U25154 (N_25154,N_23579,N_22990);
xnor U25155 (N_25155,N_22736,N_23239);
xor U25156 (N_25156,N_22567,N_22609);
xnor U25157 (N_25157,N_23732,N_23376);
xnor U25158 (N_25158,N_22941,N_23952);
and U25159 (N_25159,N_23744,N_22763);
nand U25160 (N_25160,N_23273,N_23219);
or U25161 (N_25161,N_22712,N_22608);
and U25162 (N_25162,N_23469,N_22740);
nand U25163 (N_25163,N_23479,N_23897);
nor U25164 (N_25164,N_23840,N_23958);
or U25165 (N_25165,N_23938,N_22531);
xor U25166 (N_25166,N_23732,N_23779);
xor U25167 (N_25167,N_22926,N_23405);
or U25168 (N_25168,N_22665,N_23150);
or U25169 (N_25169,N_22668,N_23018);
nor U25170 (N_25170,N_23246,N_23398);
xor U25171 (N_25171,N_22827,N_23222);
nor U25172 (N_25172,N_22783,N_23885);
nand U25173 (N_25173,N_22928,N_23739);
nor U25174 (N_25174,N_23860,N_23659);
nand U25175 (N_25175,N_23257,N_22668);
nand U25176 (N_25176,N_22994,N_23078);
or U25177 (N_25177,N_23979,N_23903);
nor U25178 (N_25178,N_23341,N_22884);
nand U25179 (N_25179,N_22954,N_23521);
nor U25180 (N_25180,N_23132,N_22581);
or U25181 (N_25181,N_22766,N_23249);
nand U25182 (N_25182,N_22981,N_23429);
nor U25183 (N_25183,N_23537,N_23174);
xnor U25184 (N_25184,N_23610,N_23358);
or U25185 (N_25185,N_23634,N_23104);
xor U25186 (N_25186,N_22905,N_23344);
xor U25187 (N_25187,N_23523,N_23612);
nor U25188 (N_25188,N_23693,N_23402);
or U25189 (N_25189,N_22952,N_23490);
xor U25190 (N_25190,N_22900,N_23031);
or U25191 (N_25191,N_22667,N_23974);
xor U25192 (N_25192,N_23690,N_23832);
xor U25193 (N_25193,N_22554,N_23807);
or U25194 (N_25194,N_23262,N_23027);
xnor U25195 (N_25195,N_23206,N_23151);
and U25196 (N_25196,N_23248,N_22793);
xnor U25197 (N_25197,N_23015,N_23456);
and U25198 (N_25198,N_23786,N_23110);
nor U25199 (N_25199,N_23673,N_23628);
nor U25200 (N_25200,N_23103,N_23083);
xor U25201 (N_25201,N_23144,N_22790);
or U25202 (N_25202,N_23424,N_22608);
or U25203 (N_25203,N_23207,N_22830);
nand U25204 (N_25204,N_22650,N_23001);
nor U25205 (N_25205,N_22746,N_22782);
or U25206 (N_25206,N_22705,N_23413);
and U25207 (N_25207,N_23726,N_23212);
nand U25208 (N_25208,N_22732,N_23848);
xor U25209 (N_25209,N_23423,N_22607);
nand U25210 (N_25210,N_22571,N_23372);
or U25211 (N_25211,N_22501,N_22934);
nor U25212 (N_25212,N_23707,N_23599);
nand U25213 (N_25213,N_22965,N_23948);
xor U25214 (N_25214,N_22781,N_23447);
and U25215 (N_25215,N_22753,N_22632);
or U25216 (N_25216,N_23756,N_23468);
nor U25217 (N_25217,N_22719,N_23343);
and U25218 (N_25218,N_23915,N_23736);
nor U25219 (N_25219,N_22766,N_23339);
xnor U25220 (N_25220,N_23479,N_23405);
nor U25221 (N_25221,N_23539,N_23622);
xnor U25222 (N_25222,N_23029,N_23137);
nand U25223 (N_25223,N_23762,N_22607);
xor U25224 (N_25224,N_23292,N_23059);
nand U25225 (N_25225,N_22871,N_23153);
or U25226 (N_25226,N_23569,N_22977);
xor U25227 (N_25227,N_23868,N_22680);
or U25228 (N_25228,N_23162,N_23499);
or U25229 (N_25229,N_22879,N_23056);
or U25230 (N_25230,N_22860,N_23655);
nand U25231 (N_25231,N_23575,N_23646);
nand U25232 (N_25232,N_23243,N_22873);
nand U25233 (N_25233,N_23649,N_23941);
xnor U25234 (N_25234,N_22903,N_23262);
nand U25235 (N_25235,N_23198,N_23331);
nor U25236 (N_25236,N_23234,N_22740);
and U25237 (N_25237,N_23953,N_23241);
or U25238 (N_25238,N_22808,N_22866);
and U25239 (N_25239,N_22516,N_23208);
xnor U25240 (N_25240,N_23608,N_23005);
nand U25241 (N_25241,N_23984,N_23239);
xnor U25242 (N_25242,N_22634,N_23587);
xnor U25243 (N_25243,N_23550,N_23138);
xor U25244 (N_25244,N_23420,N_23206);
or U25245 (N_25245,N_22960,N_23491);
nor U25246 (N_25246,N_23523,N_22728);
or U25247 (N_25247,N_23284,N_23794);
xnor U25248 (N_25248,N_22732,N_22875);
nor U25249 (N_25249,N_23139,N_23932);
nor U25250 (N_25250,N_23055,N_22572);
nor U25251 (N_25251,N_22622,N_23225);
or U25252 (N_25252,N_23572,N_23903);
and U25253 (N_25253,N_23800,N_23407);
nand U25254 (N_25254,N_23634,N_23879);
nand U25255 (N_25255,N_23064,N_23893);
and U25256 (N_25256,N_23156,N_23161);
nand U25257 (N_25257,N_23706,N_23525);
xnor U25258 (N_25258,N_23843,N_22689);
nor U25259 (N_25259,N_22623,N_23136);
and U25260 (N_25260,N_23524,N_23823);
xnor U25261 (N_25261,N_23470,N_23480);
xor U25262 (N_25262,N_22684,N_22961);
nor U25263 (N_25263,N_22998,N_23589);
nor U25264 (N_25264,N_23403,N_23378);
xnor U25265 (N_25265,N_23238,N_23431);
nor U25266 (N_25266,N_23918,N_23186);
and U25267 (N_25267,N_23321,N_22657);
or U25268 (N_25268,N_22549,N_22627);
nand U25269 (N_25269,N_23414,N_23914);
and U25270 (N_25270,N_23393,N_22750);
or U25271 (N_25271,N_23011,N_22997);
nand U25272 (N_25272,N_22518,N_23085);
and U25273 (N_25273,N_23891,N_22754);
nand U25274 (N_25274,N_22689,N_23049);
and U25275 (N_25275,N_23959,N_22577);
nand U25276 (N_25276,N_23190,N_23544);
nand U25277 (N_25277,N_22879,N_23066);
or U25278 (N_25278,N_23929,N_23138);
xor U25279 (N_25279,N_23659,N_23546);
or U25280 (N_25280,N_23546,N_23728);
or U25281 (N_25281,N_22941,N_22818);
or U25282 (N_25282,N_23609,N_22617);
or U25283 (N_25283,N_23989,N_22690);
nand U25284 (N_25284,N_23448,N_22515);
nand U25285 (N_25285,N_23270,N_22863);
and U25286 (N_25286,N_23759,N_23393);
or U25287 (N_25287,N_22961,N_23786);
xor U25288 (N_25288,N_23385,N_22514);
nand U25289 (N_25289,N_22842,N_23472);
xor U25290 (N_25290,N_23875,N_22812);
xor U25291 (N_25291,N_23799,N_23515);
nor U25292 (N_25292,N_23750,N_22747);
xor U25293 (N_25293,N_23614,N_23122);
xnor U25294 (N_25294,N_23326,N_22558);
nor U25295 (N_25295,N_23239,N_23738);
xnor U25296 (N_25296,N_23152,N_23659);
nand U25297 (N_25297,N_23229,N_23692);
nor U25298 (N_25298,N_23839,N_23014);
and U25299 (N_25299,N_23659,N_23667);
or U25300 (N_25300,N_23692,N_23502);
xnor U25301 (N_25301,N_22915,N_23489);
nand U25302 (N_25302,N_23339,N_23520);
nand U25303 (N_25303,N_22765,N_22724);
nand U25304 (N_25304,N_23737,N_22940);
nand U25305 (N_25305,N_23731,N_22893);
or U25306 (N_25306,N_23084,N_22970);
xor U25307 (N_25307,N_23217,N_23465);
nand U25308 (N_25308,N_23571,N_22795);
xor U25309 (N_25309,N_23928,N_22821);
nor U25310 (N_25310,N_22995,N_22637);
nor U25311 (N_25311,N_23281,N_22975);
and U25312 (N_25312,N_23526,N_23719);
nand U25313 (N_25313,N_22695,N_22685);
and U25314 (N_25314,N_23177,N_22659);
and U25315 (N_25315,N_23067,N_23950);
or U25316 (N_25316,N_23554,N_23970);
nand U25317 (N_25317,N_22699,N_23726);
nand U25318 (N_25318,N_22626,N_22812);
nand U25319 (N_25319,N_22683,N_23258);
xnor U25320 (N_25320,N_23178,N_23722);
or U25321 (N_25321,N_23889,N_22966);
nand U25322 (N_25322,N_23197,N_23358);
and U25323 (N_25323,N_22754,N_23246);
xnor U25324 (N_25324,N_23638,N_23226);
and U25325 (N_25325,N_23961,N_23126);
xnor U25326 (N_25326,N_22543,N_23365);
xor U25327 (N_25327,N_23560,N_23422);
or U25328 (N_25328,N_23351,N_23717);
nor U25329 (N_25329,N_23457,N_22768);
and U25330 (N_25330,N_23137,N_23948);
or U25331 (N_25331,N_23287,N_22842);
or U25332 (N_25332,N_22568,N_22811);
nor U25333 (N_25333,N_23395,N_23477);
or U25334 (N_25334,N_22738,N_23790);
and U25335 (N_25335,N_22960,N_23502);
nand U25336 (N_25336,N_22853,N_23930);
or U25337 (N_25337,N_22596,N_23200);
and U25338 (N_25338,N_22734,N_23719);
nor U25339 (N_25339,N_23774,N_23312);
or U25340 (N_25340,N_22799,N_23419);
nand U25341 (N_25341,N_23184,N_22539);
xor U25342 (N_25342,N_22597,N_23591);
xor U25343 (N_25343,N_22701,N_23112);
nor U25344 (N_25344,N_23414,N_23991);
nor U25345 (N_25345,N_23968,N_22649);
nor U25346 (N_25346,N_22538,N_22782);
and U25347 (N_25347,N_22835,N_22575);
nand U25348 (N_25348,N_22608,N_23405);
or U25349 (N_25349,N_23408,N_23348);
nor U25350 (N_25350,N_23251,N_23340);
and U25351 (N_25351,N_23197,N_23716);
nor U25352 (N_25352,N_23341,N_23644);
nand U25353 (N_25353,N_22758,N_23401);
nor U25354 (N_25354,N_23372,N_22582);
xor U25355 (N_25355,N_22628,N_23518);
and U25356 (N_25356,N_23589,N_23828);
xor U25357 (N_25357,N_22683,N_23766);
xnor U25358 (N_25358,N_23384,N_23538);
and U25359 (N_25359,N_22957,N_23773);
xor U25360 (N_25360,N_23921,N_22796);
nor U25361 (N_25361,N_23538,N_23438);
xor U25362 (N_25362,N_23612,N_23342);
nor U25363 (N_25363,N_23475,N_23574);
nand U25364 (N_25364,N_23059,N_23640);
nand U25365 (N_25365,N_23618,N_23168);
or U25366 (N_25366,N_23875,N_23859);
xor U25367 (N_25367,N_23243,N_22520);
xor U25368 (N_25368,N_23891,N_23028);
nor U25369 (N_25369,N_23816,N_22793);
xor U25370 (N_25370,N_23560,N_22858);
nor U25371 (N_25371,N_23639,N_23158);
or U25372 (N_25372,N_23358,N_22882);
nand U25373 (N_25373,N_23490,N_23774);
or U25374 (N_25374,N_23488,N_23714);
or U25375 (N_25375,N_23225,N_22746);
nand U25376 (N_25376,N_23265,N_22624);
xor U25377 (N_25377,N_23294,N_23303);
or U25378 (N_25378,N_22803,N_23426);
or U25379 (N_25379,N_23364,N_23714);
and U25380 (N_25380,N_23976,N_23403);
nor U25381 (N_25381,N_22860,N_23800);
xnor U25382 (N_25382,N_22757,N_22627);
and U25383 (N_25383,N_23955,N_22512);
and U25384 (N_25384,N_23058,N_23317);
nand U25385 (N_25385,N_22533,N_22821);
and U25386 (N_25386,N_23505,N_23824);
nand U25387 (N_25387,N_23808,N_23181);
nor U25388 (N_25388,N_23725,N_22912);
xor U25389 (N_25389,N_22892,N_23666);
xnor U25390 (N_25390,N_23432,N_22797);
or U25391 (N_25391,N_23028,N_23871);
or U25392 (N_25392,N_22612,N_23743);
nor U25393 (N_25393,N_23731,N_22942);
nor U25394 (N_25394,N_23938,N_23773);
nand U25395 (N_25395,N_23046,N_22671);
xor U25396 (N_25396,N_23595,N_23513);
and U25397 (N_25397,N_23774,N_23975);
nand U25398 (N_25398,N_23473,N_23611);
xor U25399 (N_25399,N_23619,N_23804);
or U25400 (N_25400,N_23471,N_22577);
nor U25401 (N_25401,N_23696,N_22696);
or U25402 (N_25402,N_22957,N_22631);
and U25403 (N_25403,N_23666,N_23874);
xnor U25404 (N_25404,N_23594,N_23622);
nand U25405 (N_25405,N_22763,N_23568);
xor U25406 (N_25406,N_22558,N_23690);
and U25407 (N_25407,N_22712,N_23749);
nor U25408 (N_25408,N_23992,N_23186);
nand U25409 (N_25409,N_23756,N_22752);
or U25410 (N_25410,N_22544,N_23980);
nand U25411 (N_25411,N_22765,N_22894);
or U25412 (N_25412,N_23452,N_22682);
nor U25413 (N_25413,N_23166,N_22649);
nor U25414 (N_25414,N_23845,N_23502);
or U25415 (N_25415,N_23574,N_22700);
or U25416 (N_25416,N_23587,N_22772);
and U25417 (N_25417,N_23889,N_23044);
nor U25418 (N_25418,N_22755,N_23076);
nand U25419 (N_25419,N_22597,N_23608);
xor U25420 (N_25420,N_23086,N_22653);
nand U25421 (N_25421,N_22889,N_23828);
and U25422 (N_25422,N_23000,N_23424);
or U25423 (N_25423,N_23550,N_23758);
nor U25424 (N_25424,N_23821,N_23212);
xnor U25425 (N_25425,N_22807,N_23017);
xnor U25426 (N_25426,N_23049,N_23034);
nand U25427 (N_25427,N_23365,N_23078);
nor U25428 (N_25428,N_23355,N_22797);
and U25429 (N_25429,N_23328,N_23385);
and U25430 (N_25430,N_22565,N_23920);
and U25431 (N_25431,N_23931,N_23542);
and U25432 (N_25432,N_23676,N_23475);
and U25433 (N_25433,N_23493,N_22851);
nand U25434 (N_25434,N_23843,N_23669);
nand U25435 (N_25435,N_23015,N_23724);
nand U25436 (N_25436,N_22820,N_22544);
xnor U25437 (N_25437,N_22972,N_23231);
nand U25438 (N_25438,N_23884,N_23069);
and U25439 (N_25439,N_22880,N_23329);
and U25440 (N_25440,N_23756,N_23629);
nor U25441 (N_25441,N_23754,N_23139);
xnor U25442 (N_25442,N_23229,N_22820);
nor U25443 (N_25443,N_22514,N_22645);
nand U25444 (N_25444,N_22893,N_23225);
and U25445 (N_25445,N_23370,N_22513);
nor U25446 (N_25446,N_23427,N_23646);
and U25447 (N_25447,N_23156,N_22983);
and U25448 (N_25448,N_22677,N_22960);
or U25449 (N_25449,N_23669,N_23774);
xnor U25450 (N_25450,N_23446,N_23968);
or U25451 (N_25451,N_22719,N_22977);
nor U25452 (N_25452,N_23748,N_22595);
xnor U25453 (N_25453,N_23641,N_23334);
xor U25454 (N_25454,N_23981,N_22752);
xor U25455 (N_25455,N_23331,N_22853);
xor U25456 (N_25456,N_23027,N_23543);
nor U25457 (N_25457,N_23254,N_23404);
xnor U25458 (N_25458,N_22756,N_23965);
or U25459 (N_25459,N_23512,N_22963);
nor U25460 (N_25460,N_22765,N_22821);
xor U25461 (N_25461,N_23402,N_23285);
xnor U25462 (N_25462,N_23189,N_23646);
or U25463 (N_25463,N_23072,N_23160);
or U25464 (N_25464,N_23501,N_23913);
nor U25465 (N_25465,N_23949,N_23943);
nand U25466 (N_25466,N_23081,N_23234);
nand U25467 (N_25467,N_23172,N_23383);
xnor U25468 (N_25468,N_22925,N_23358);
or U25469 (N_25469,N_22730,N_22658);
or U25470 (N_25470,N_22959,N_23150);
xor U25471 (N_25471,N_23975,N_22764);
nor U25472 (N_25472,N_22574,N_23577);
nor U25473 (N_25473,N_23338,N_22679);
nand U25474 (N_25474,N_22671,N_23866);
nand U25475 (N_25475,N_22943,N_23717);
xnor U25476 (N_25476,N_23799,N_23986);
xnor U25477 (N_25477,N_22611,N_22875);
nor U25478 (N_25478,N_23662,N_22806);
or U25479 (N_25479,N_23556,N_22676);
or U25480 (N_25480,N_23914,N_23910);
and U25481 (N_25481,N_23623,N_22517);
nor U25482 (N_25482,N_23829,N_23182);
nand U25483 (N_25483,N_23036,N_23195);
or U25484 (N_25484,N_23030,N_22727);
nand U25485 (N_25485,N_23810,N_23489);
or U25486 (N_25486,N_23980,N_23577);
and U25487 (N_25487,N_22965,N_22986);
or U25488 (N_25488,N_23506,N_23635);
and U25489 (N_25489,N_23002,N_22500);
xor U25490 (N_25490,N_23729,N_23128);
xnor U25491 (N_25491,N_23841,N_23493);
xnor U25492 (N_25492,N_23321,N_23458);
xnor U25493 (N_25493,N_23432,N_23846);
and U25494 (N_25494,N_22901,N_22540);
nor U25495 (N_25495,N_23740,N_23353);
or U25496 (N_25496,N_23350,N_23223);
nor U25497 (N_25497,N_23991,N_23816);
and U25498 (N_25498,N_23422,N_23024);
and U25499 (N_25499,N_22867,N_22656);
nand U25500 (N_25500,N_25023,N_25103);
nand U25501 (N_25501,N_24664,N_24087);
and U25502 (N_25502,N_25395,N_24885);
nand U25503 (N_25503,N_24868,N_24118);
nand U25504 (N_25504,N_25481,N_24147);
and U25505 (N_25505,N_25078,N_24520);
or U25506 (N_25506,N_24004,N_25175);
or U25507 (N_25507,N_25096,N_24609);
or U25508 (N_25508,N_24494,N_25032);
or U25509 (N_25509,N_25012,N_24600);
xor U25510 (N_25510,N_24020,N_24248);
or U25511 (N_25511,N_25225,N_25014);
and U25512 (N_25512,N_25140,N_24431);
nand U25513 (N_25513,N_25290,N_24576);
and U25514 (N_25514,N_24077,N_25455);
nand U25515 (N_25515,N_24218,N_24000);
nand U25516 (N_25516,N_24382,N_25322);
nand U25517 (N_25517,N_24303,N_24247);
nor U25518 (N_25518,N_24794,N_25282);
or U25519 (N_25519,N_25362,N_24357);
nor U25520 (N_25520,N_24737,N_25198);
xor U25521 (N_25521,N_24208,N_24710);
nor U25522 (N_25522,N_25356,N_24030);
xor U25523 (N_25523,N_24254,N_24489);
xor U25524 (N_25524,N_24286,N_25399);
nor U25525 (N_25525,N_25240,N_24597);
xnor U25526 (N_25526,N_24916,N_24844);
and U25527 (N_25527,N_25365,N_24073);
or U25528 (N_25528,N_24728,N_24646);
xnor U25529 (N_25529,N_25045,N_24793);
and U25530 (N_25530,N_24134,N_25107);
xor U25531 (N_25531,N_24581,N_24864);
and U25532 (N_25532,N_24309,N_24536);
or U25533 (N_25533,N_25017,N_24679);
nor U25534 (N_25534,N_24585,N_24858);
and U25535 (N_25535,N_25200,N_25030);
nand U25536 (N_25536,N_25304,N_24946);
or U25537 (N_25537,N_24748,N_24805);
xnor U25538 (N_25538,N_24818,N_24525);
xor U25539 (N_25539,N_25446,N_25047);
xnor U25540 (N_25540,N_24194,N_24475);
and U25541 (N_25541,N_25011,N_24156);
xor U25542 (N_25542,N_24468,N_24275);
or U25543 (N_25543,N_24028,N_24908);
and U25544 (N_25544,N_24022,N_24438);
nor U25545 (N_25545,N_25280,N_24036);
nor U25546 (N_25546,N_25270,N_25217);
or U25547 (N_25547,N_24097,N_25154);
or U25548 (N_25548,N_24562,N_25005);
nand U25549 (N_25549,N_24932,N_25233);
or U25550 (N_25550,N_25347,N_25434);
xnor U25551 (N_25551,N_24522,N_25123);
or U25552 (N_25552,N_25259,N_24950);
nand U25553 (N_25553,N_24310,N_24974);
or U25554 (N_25554,N_24219,N_24680);
xor U25555 (N_25555,N_25401,N_24855);
nor U25556 (N_25556,N_24010,N_24406);
nand U25557 (N_25557,N_24682,N_24377);
nand U25558 (N_25558,N_24743,N_24298);
and U25559 (N_25559,N_24344,N_25264);
nand U25560 (N_25560,N_24982,N_24207);
or U25561 (N_25561,N_24258,N_25367);
nor U25562 (N_25562,N_24435,N_24112);
xnor U25563 (N_25563,N_25036,N_24952);
or U25564 (N_25564,N_24083,N_24658);
nor U25565 (N_25565,N_25316,N_25223);
and U25566 (N_25566,N_24423,N_25370);
and U25567 (N_25567,N_25176,N_25432);
nor U25568 (N_25568,N_25443,N_24325);
nor U25569 (N_25569,N_24441,N_24553);
and U25570 (N_25570,N_25102,N_25268);
nand U25571 (N_25571,N_25160,N_24933);
nand U25572 (N_25572,N_24662,N_25207);
or U25573 (N_25573,N_25188,N_24740);
or U25574 (N_25574,N_25345,N_25049);
and U25575 (N_25575,N_25374,N_24398);
nor U25576 (N_25576,N_24356,N_25413);
or U25577 (N_25577,N_24718,N_24419);
nor U25578 (N_25578,N_25122,N_25069);
xor U25579 (N_25579,N_24867,N_24162);
nand U25580 (N_25580,N_24615,N_24428);
xnor U25581 (N_25581,N_24695,N_24798);
nor U25582 (N_25582,N_24947,N_24624);
xor U25583 (N_25583,N_25380,N_24394);
and U25584 (N_25584,N_25031,N_24215);
and U25585 (N_25585,N_24098,N_25189);
xnor U25586 (N_25586,N_24365,N_24928);
and U25587 (N_25587,N_24267,N_25174);
and U25588 (N_25588,N_25281,N_25241);
or U25589 (N_25589,N_24584,N_24314);
and U25590 (N_25590,N_24560,N_24359);
xor U25591 (N_25591,N_24980,N_25468);
nand U25592 (N_25592,N_24274,N_25085);
or U25593 (N_25593,N_24951,N_24228);
and U25594 (N_25594,N_25067,N_24111);
nand U25595 (N_25595,N_24271,N_24660);
xor U25596 (N_25596,N_24404,N_24455);
xnor U25597 (N_25597,N_24734,N_24973);
xor U25598 (N_25598,N_25495,N_24461);
xnor U25599 (N_25599,N_24556,N_24714);
nand U25600 (N_25600,N_24319,N_24145);
xnor U25601 (N_25601,N_25035,N_24711);
xnor U25602 (N_25602,N_25235,N_24211);
and U25603 (N_25603,N_25063,N_24586);
or U25604 (N_25604,N_25405,N_24893);
xor U25605 (N_25605,N_24446,N_25295);
nand U25606 (N_25606,N_24549,N_25192);
nor U25607 (N_25607,N_25210,N_25263);
or U25608 (N_25608,N_25283,N_24239);
nor U25609 (N_25609,N_25288,N_25287);
nor U25610 (N_25610,N_24393,N_24306);
or U25611 (N_25611,N_25289,N_24003);
nand U25612 (N_25612,N_24488,N_24392);
and U25613 (N_25613,N_24834,N_25279);
xor U25614 (N_25614,N_24639,N_25359);
nand U25615 (N_25615,N_24074,N_24625);
or U25616 (N_25616,N_24535,N_24548);
nor U25617 (N_25617,N_24065,N_24216);
xnor U25618 (N_25618,N_24311,N_25179);
xor U25619 (N_25619,N_25342,N_24316);
nand U25620 (N_25620,N_24617,N_24371);
xor U25621 (N_25621,N_24029,N_25084);
nor U25622 (N_25622,N_24882,N_24731);
nor U25623 (N_25623,N_25002,N_25144);
nand U25624 (N_25624,N_24913,N_24761);
nand U25625 (N_25625,N_25054,N_24294);
nand U25626 (N_25626,N_25185,N_25250);
nand U25627 (N_25627,N_24165,N_24315);
or U25628 (N_25628,N_24747,N_25056);
and U25629 (N_25629,N_25389,N_25204);
and U25630 (N_25630,N_24607,N_24861);
nor U25631 (N_25631,N_24395,N_24039);
nand U25632 (N_25632,N_25350,N_25007);
nand U25633 (N_25633,N_24801,N_24860);
and U25634 (N_25634,N_24160,N_24230);
nor U25635 (N_25635,N_24440,N_24132);
or U25636 (N_25636,N_24785,N_24757);
and U25637 (N_25637,N_25046,N_24895);
xnor U25638 (N_25638,N_24719,N_24199);
xnor U25639 (N_25639,N_24119,N_25221);
nand U25640 (N_25640,N_25034,N_24340);
or U25641 (N_25641,N_24724,N_24846);
nand U25642 (N_25642,N_24222,N_24091);
xor U25643 (N_25643,N_25141,N_24811);
or U25644 (N_25644,N_25145,N_25499);
nand U25645 (N_25645,N_25152,N_25465);
or U25646 (N_25646,N_24102,N_25022);
and U25647 (N_25647,N_24852,N_24399);
xor U25648 (N_25648,N_25497,N_24405);
and U25649 (N_25649,N_25454,N_24715);
or U25650 (N_25650,N_24642,N_24063);
nor U25651 (N_25651,N_25134,N_25202);
xor U25652 (N_25652,N_25422,N_24959);
nor U25653 (N_25653,N_24587,N_24764);
and U25654 (N_25654,N_25068,N_25383);
and U25655 (N_25655,N_24904,N_25110);
nand U25656 (N_25656,N_24583,N_24327);
or U25657 (N_25657,N_25000,N_24690);
and U25658 (N_25658,N_25149,N_24200);
and U25659 (N_25659,N_24277,N_24804);
or U25660 (N_25660,N_24100,N_24031);
nand U25661 (N_25661,N_24700,N_25494);
and U25662 (N_25662,N_24550,N_24927);
or U25663 (N_25663,N_24850,N_24246);
xnor U25664 (N_25664,N_25245,N_25199);
nand U25665 (N_25665,N_24055,N_24923);
nor U25666 (N_25666,N_24040,N_24839);
xnor U25667 (N_25667,N_24188,N_25273);
nor U25668 (N_25668,N_24092,N_24786);
nor U25669 (N_25669,N_24061,N_25037);
and U25670 (N_25670,N_24444,N_24921);
xor U25671 (N_25671,N_24348,N_24568);
nor U25672 (N_25672,N_25331,N_24762);
xor U25673 (N_25673,N_24414,N_25246);
nor U25674 (N_25674,N_24108,N_25244);
and U25675 (N_25675,N_25412,N_25206);
xor U25676 (N_25676,N_24606,N_25150);
or U25677 (N_25677,N_25409,N_25439);
nand U25678 (N_25678,N_24857,N_25253);
nor U25679 (N_25679,N_24524,N_24631);
xnor U25680 (N_25680,N_25087,N_24621);
and U25681 (N_25681,N_24675,N_24209);
xnor U25682 (N_25682,N_24692,N_25423);
nand U25683 (N_25683,N_24351,N_24840);
nand U25684 (N_25684,N_25033,N_25449);
and U25685 (N_25685,N_24129,N_24096);
nand U25686 (N_25686,N_24025,N_24939);
nor U25687 (N_25687,N_25469,N_24139);
xnor U25688 (N_25688,N_24047,N_25417);
and U25689 (N_25689,N_24683,N_24221);
nor U25690 (N_25690,N_24969,N_25301);
or U25691 (N_25691,N_25187,N_24744);
xor U25692 (N_25692,N_25115,N_24835);
xnor U25693 (N_25693,N_24516,N_25095);
xnor U25694 (N_25694,N_24523,N_24323);
or U25695 (N_25695,N_25209,N_24305);
and U25696 (N_25696,N_24645,N_25062);
nand U25697 (N_25697,N_24802,N_24651);
xor U25698 (N_25698,N_24978,N_24957);
and U25699 (N_25699,N_24270,N_24842);
or U25700 (N_25700,N_24579,N_25184);
xor U25701 (N_25701,N_24128,N_24300);
or U25702 (N_25702,N_25232,N_25489);
xnor U25703 (N_25703,N_25111,N_24693);
nor U25704 (N_25704,N_24497,N_24499);
and U25705 (N_25705,N_24429,N_24241);
nand U25706 (N_25706,N_25003,N_24865);
and U25707 (N_25707,N_25091,N_24322);
nand U25708 (N_25708,N_25013,N_24886);
nor U25709 (N_25709,N_25008,N_25298);
nand U25710 (N_25710,N_25098,N_24292);
and U25711 (N_25711,N_24563,N_24380);
xor U25712 (N_25712,N_24157,N_24276);
nor U25713 (N_25713,N_24436,N_25071);
xnor U25714 (N_25714,N_24237,N_25226);
or U25715 (N_25715,N_25337,N_25112);
and U25716 (N_25716,N_25137,N_24821);
and U25717 (N_25717,N_24295,N_25219);
nand U25718 (N_25718,N_24832,N_24005);
and U25719 (N_25719,N_25349,N_24827);
and U25720 (N_25720,N_25048,N_24756);
nand U25721 (N_25721,N_24674,N_24140);
nand U25722 (N_25722,N_24984,N_24390);
or U25723 (N_25723,N_24605,N_25324);
nand U25724 (N_25724,N_25478,N_24647);
or U25725 (N_25725,N_24396,N_24822);
nor U25726 (N_25726,N_24830,N_24352);
or U25727 (N_25727,N_24153,N_24224);
nor U25728 (N_25728,N_24686,N_24954);
nand U25729 (N_25729,N_25116,N_24771);
nand U25730 (N_25730,N_24925,N_25173);
xor U25731 (N_25731,N_24596,N_24926);
and U25732 (N_25732,N_25101,N_24593);
or U25733 (N_25733,N_25404,N_25220);
or U25734 (N_25734,N_24511,N_25428);
or U25735 (N_25735,N_24993,N_24462);
nor U25736 (N_25736,N_24349,N_24866);
and U25737 (N_25737,N_25211,N_24767);
nor U25738 (N_25738,N_24777,N_24180);
nand U25739 (N_25739,N_24825,N_25089);
nor U25740 (N_25740,N_24759,N_25234);
or U25741 (N_25741,N_24149,N_24387);
xnor U25742 (N_25742,N_24612,N_24899);
or U25743 (N_25743,N_24198,N_25159);
or U25744 (N_25744,N_24565,N_24317);
nand U25745 (N_25745,N_24027,N_25208);
nor U25746 (N_25746,N_25132,N_25320);
nand U25747 (N_25747,N_24422,N_24884);
nor U25748 (N_25748,N_25402,N_25213);
nor U25749 (N_25749,N_25484,N_24705);
nand U25750 (N_25750,N_25010,N_25332);
nor U25751 (N_25751,N_24929,N_25238);
nand U25752 (N_25752,N_25090,N_25334);
nor U25753 (N_25753,N_24673,N_25124);
nor U25754 (N_25754,N_25027,N_24726);
nand U25755 (N_25755,N_25265,N_24150);
xor U25756 (N_25756,N_25450,N_25178);
xor U25757 (N_25757,N_25127,N_24809);
nand U25758 (N_25758,N_24910,N_24467);
or U25759 (N_25759,N_24637,N_25104);
nor U25760 (N_25760,N_24226,N_25488);
nor U25761 (N_25761,N_24813,N_25269);
or U25762 (N_25762,N_25292,N_24350);
nand U25763 (N_25763,N_24629,N_24627);
nand U25764 (N_25764,N_25351,N_24722);
nand U25765 (N_25765,N_25128,N_24236);
nor U25766 (N_25766,N_24936,N_24883);
or U25767 (N_25767,N_24273,N_25146);
and U25768 (N_25768,N_25165,N_25181);
or U25769 (N_25769,N_25384,N_24244);
and U25770 (N_25770,N_25352,N_25336);
nand U25771 (N_25771,N_25305,N_24554);
nor U25772 (N_25772,N_25406,N_25441);
nand U25773 (N_25773,N_25314,N_25415);
xor U25774 (N_25774,N_24545,N_24375);
xor U25775 (N_25775,N_24477,N_24965);
and U25776 (N_25776,N_24113,N_24580);
or U25777 (N_25777,N_24427,N_24183);
and U25778 (N_25778,N_24931,N_24019);
or U25779 (N_25779,N_24082,N_24308);
or U25780 (N_25780,N_24388,N_24824);
or U25781 (N_25781,N_25474,N_24613);
nor U25782 (N_25782,N_24173,N_24033);
and U25783 (N_25783,N_24589,N_24355);
nor U25784 (N_25784,N_24291,N_24512);
xnor U25785 (N_25785,N_24502,N_24796);
nand U25786 (N_25786,N_25106,N_25135);
nor U25787 (N_25787,N_25471,N_24127);
or U25788 (N_25788,N_25074,N_25133);
and U25789 (N_25789,N_24848,N_24900);
xnor U25790 (N_25790,N_24217,N_24665);
nor U25791 (N_25791,N_24815,N_24363);
and U25792 (N_25792,N_24603,N_24206);
or U25793 (N_25793,N_25311,N_24329);
and U25794 (N_25794,N_24555,N_24820);
nand U25795 (N_25795,N_24046,N_24810);
xor U25796 (N_25796,N_24358,N_24880);
or U25797 (N_25797,N_24730,N_24301);
or U25798 (N_25798,N_25357,N_24024);
nor U25799 (N_25799,N_25461,N_24540);
or U25800 (N_25800,N_24093,N_25093);
nand U25801 (N_25801,N_24197,N_25195);
or U25802 (N_25802,N_25157,N_25252);
or U25803 (N_25803,N_25437,N_25186);
nor U25804 (N_25804,N_24938,N_24590);
nand U25805 (N_25805,N_24917,N_25492);
nand U25806 (N_25806,N_24628,N_24812);
or U25807 (N_25807,N_25243,N_24470);
or U25808 (N_25808,N_24122,N_25391);
and U25809 (N_25809,N_24347,N_25343);
and U25810 (N_25810,N_24282,N_24391);
and U25811 (N_25811,N_24691,N_25438);
and U25812 (N_25812,N_24630,N_24706);
nand U25813 (N_25813,N_24038,N_24935);
and U25814 (N_25814,N_24843,N_25148);
and U25815 (N_25815,N_24752,N_25139);
or U25816 (N_25816,N_24044,N_24066);
nand U25817 (N_25817,N_24018,N_25129);
nor U25818 (N_25818,N_24459,N_25073);
nor U25819 (N_25819,N_24203,N_25042);
nor U25820 (N_25820,N_24849,N_24471);
nor U25821 (N_25821,N_24782,N_24486);
or U25822 (N_25822,N_25303,N_25327);
and U25823 (N_25823,N_25004,N_24988);
xor U25824 (N_25824,N_24790,N_24888);
xor U25825 (N_25825,N_24413,N_24775);
nor U25826 (N_25826,N_24799,N_24879);
nor U25827 (N_25827,N_24360,N_24769);
or U25828 (N_25828,N_24643,N_24177);
or U25829 (N_25829,N_25029,N_25097);
nor U25830 (N_25830,N_24465,N_24688);
xor U25831 (N_25831,N_24281,N_24896);
or U25832 (N_25832,N_24453,N_24551);
nand U25833 (N_25833,N_24725,N_24774);
or U25834 (N_25834,N_24478,N_24531);
or U25835 (N_25835,N_24434,N_25070);
nor U25836 (N_25836,N_24086,N_24169);
nor U25837 (N_25837,N_24573,N_24723);
nor U25838 (N_25838,N_24800,N_24233);
nor U25839 (N_25839,N_24614,N_24519);
and U25840 (N_25840,N_24255,N_25444);
or U25841 (N_25841,N_25118,N_24176);
and U25842 (N_25842,N_24289,N_24945);
nand U25843 (N_25843,N_25168,N_25052);
and U25844 (N_25844,N_25183,N_24015);
nor U25845 (N_25845,N_24313,N_25039);
nor U25846 (N_25846,N_24501,N_24697);
nor U25847 (N_25847,N_25020,N_24179);
xor U25848 (N_25848,N_24374,N_24669);
xor U25849 (N_25849,N_25307,N_24966);
and U25850 (N_25850,N_24163,N_24094);
or U25851 (N_25851,N_24079,N_24862);
or U25852 (N_25852,N_24016,N_24182);
xor U25853 (N_25853,N_25445,N_24114);
or U25854 (N_25854,N_24749,N_25044);
nand U25855 (N_25855,N_24681,N_24495);
or U25856 (N_25856,N_24911,N_25167);
and U25857 (N_25857,N_25256,N_24368);
or U25858 (N_25858,N_25258,N_24559);
xnor U25859 (N_25859,N_24996,N_24870);
nand U25860 (N_25860,N_24526,N_25425);
xor U25861 (N_25861,N_25486,N_25358);
nor U25862 (N_25862,N_25040,N_24212);
or U25863 (N_25863,N_24971,N_24068);
nor U25864 (N_25864,N_24223,N_25205);
xor U25865 (N_25865,N_25169,N_24956);
nor U25866 (N_25866,N_24653,N_25231);
and U25867 (N_25867,N_24123,N_24720);
nor U25868 (N_25868,N_25453,N_25296);
and U25869 (N_25869,N_24213,N_25064);
nor U25870 (N_25870,N_24460,N_25171);
or U25871 (N_25871,N_24738,N_24408);
and U25872 (N_25872,N_24085,N_24997);
xnor U25873 (N_25873,N_24121,N_24514);
or U25874 (N_25874,N_25294,N_25161);
nor U25875 (N_25875,N_24701,N_25487);
nand U25876 (N_25876,N_25328,N_24265);
xor U25877 (N_25877,N_24506,N_24443);
and U25878 (N_25878,N_24474,N_24569);
nor U25879 (N_25879,N_24369,N_24684);
nor U25880 (N_25880,N_25398,N_24527);
nand U25881 (N_25881,N_24227,N_24713);
nor U25882 (N_25882,N_24250,N_25457);
or U25883 (N_25883,N_24402,N_24411);
xnor U25884 (N_25884,N_25119,N_25431);
nand U25885 (N_25885,N_24873,N_24064);
xnor U25886 (N_25886,N_24304,N_25385);
and U25887 (N_25887,N_24937,N_24986);
or U25888 (N_25888,N_24518,N_25435);
xor U25889 (N_25889,N_24558,N_24547);
nand U25890 (N_25890,N_25251,N_25050);
nand U25891 (N_25891,N_24766,N_25051);
nor U25892 (N_25892,N_25080,N_24591);
nor U25893 (N_25893,N_24454,N_24007);
xnor U25894 (N_25894,N_25275,N_24878);
xor U25895 (N_25895,N_24906,N_24561);
nand U25896 (N_25896,N_24017,N_25429);
nand U25897 (N_25897,N_25339,N_25182);
and U25898 (N_25898,N_24135,N_24707);
xor U25899 (N_25899,N_24949,N_24205);
or U25900 (N_25900,N_24386,N_24542);
and U25901 (N_25901,N_25479,N_25255);
nor U25902 (N_25902,N_24712,N_24469);
or U25903 (N_25903,N_24253,N_24975);
and U25904 (N_25904,N_24345,N_25355);
nand U25905 (N_25905,N_24998,N_24940);
nor U25906 (N_25906,N_25392,N_24326);
nor U25907 (N_25907,N_24828,N_24159);
or U25908 (N_25908,N_24678,N_24826);
nand U25909 (N_25909,N_25079,N_24566);
nand U25910 (N_25910,N_24838,N_24034);
xor U25911 (N_25911,N_24677,N_25041);
nand U25912 (N_25912,N_24424,N_24874);
nand U25913 (N_25913,N_24795,N_24195);
and U25914 (N_25914,N_25212,N_25024);
and U25915 (N_25915,N_24171,N_24492);
and U25916 (N_25916,N_24343,N_25126);
nand U25917 (N_25917,N_25072,N_25440);
xnor U25918 (N_25918,N_24333,N_24657);
nor U25919 (N_25919,N_24238,N_25286);
or U25920 (N_25920,N_25147,N_24484);
and U25921 (N_25921,N_24190,N_24339);
or U25922 (N_25922,N_25267,N_24078);
nor U25923 (N_25923,N_24336,N_24564);
nand U25924 (N_25924,N_24192,N_25346);
nor U25925 (N_25925,N_24919,N_24042);
nor U25926 (N_25926,N_24447,N_24736);
xnor U25927 (N_25927,N_24955,N_24831);
nand U25928 (N_25928,N_24131,N_24633);
xnor U25929 (N_25929,N_24856,N_24152);
and U25930 (N_25930,N_25430,N_24417);
or U25931 (N_25931,N_25239,N_24330);
or U25932 (N_25932,N_24768,N_25153);
nand U25933 (N_25933,N_24620,N_25373);
and U25934 (N_25934,N_25081,N_25467);
nor U25935 (N_25935,N_25249,N_25170);
or U25936 (N_25936,N_24635,N_24035);
nand U25937 (N_25937,N_24403,N_24485);
nand U25938 (N_25938,N_24008,N_24505);
or U25939 (N_25939,N_24362,N_24299);
xnor U25940 (N_25940,N_24708,N_24293);
xor U25941 (N_25941,N_24186,N_24266);
nor U25942 (N_25942,N_24739,N_25361);
nor U25943 (N_25943,N_25201,N_24482);
nand U25944 (N_25944,N_24072,N_25396);
nor U25945 (N_25945,N_24918,N_24765);
nand U25946 (N_25946,N_24872,N_24136);
or U25947 (N_25947,N_24481,N_24970);
nand U25948 (N_25948,N_24151,N_24463);
and U25949 (N_25949,N_25379,N_25371);
and U25950 (N_25950,N_24806,N_24532);
nand U25951 (N_25951,N_25216,N_24797);
and U25952 (N_25952,N_24823,N_24672);
nor U25953 (N_25953,N_25242,N_24841);
and U25954 (N_25954,N_24816,N_24307);
nand U25955 (N_25955,N_24106,N_24164);
and U25956 (N_25956,N_24694,N_24280);
nand U25957 (N_25957,N_25006,N_24601);
nor U25958 (N_25958,N_24479,N_24504);
and U25959 (N_25959,N_24331,N_24490);
nand U25960 (N_25960,N_24619,N_25197);
xnor U25961 (N_25961,N_24041,N_25297);
nor U25962 (N_25962,N_24338,N_24418);
and U25963 (N_25963,N_24592,N_25448);
and U25964 (N_25964,N_24174,N_25318);
nor U25965 (N_25965,N_24451,N_24229);
nand U25966 (N_25966,N_24328,N_24269);
and U25967 (N_25967,N_24751,N_24659);
nand U25968 (N_25968,N_25407,N_24698);
and U25969 (N_25969,N_24903,N_24415);
xor U25970 (N_25970,N_24533,N_24787);
nor U25971 (N_25971,N_25366,N_24972);
or U25972 (N_25972,N_25458,N_24006);
xnor U25973 (N_25973,N_24458,N_24537);
or U25974 (N_25974,N_24450,N_24433);
or U25975 (N_25975,N_24154,N_24924);
nand U25976 (N_25976,N_25427,N_24059);
nor U25977 (N_25977,N_24480,N_25172);
or U25978 (N_25978,N_24517,N_25341);
or U25979 (N_25979,N_24622,N_25426);
and U25980 (N_25980,N_24144,N_25364);
nand U25981 (N_25981,N_25066,N_25442);
nor U25982 (N_25982,N_24148,N_24943);
or U25983 (N_25983,N_25317,N_25416);
nor U25984 (N_25984,N_25077,N_24656);
and U25985 (N_25985,N_24272,N_24220);
nor U25986 (N_25986,N_25300,N_25193);
nand U25987 (N_25987,N_25271,N_24529);
or U25988 (N_25988,N_24983,N_25100);
nor U25989 (N_25989,N_24193,N_24476);
xor U25990 (N_25990,N_24746,N_24930);
or U25991 (N_25991,N_24814,N_24753);
and U25992 (N_25992,N_24513,N_25460);
xnor U25993 (N_25993,N_24062,N_24142);
xor U25994 (N_25994,N_25121,N_24302);
xor U25995 (N_25995,N_24960,N_24168);
nor U25996 (N_25996,N_24175,N_25325);
and U25997 (N_25997,N_25310,N_25088);
nand U25998 (N_25998,N_24803,N_25376);
or U25999 (N_25999,N_25459,N_24242);
or U26000 (N_26000,N_25060,N_24668);
xnor U26001 (N_26001,N_24544,N_25333);
nor U26002 (N_26002,N_24191,N_25230);
and U26003 (N_26003,N_24709,N_24425);
nor U26004 (N_26004,N_24076,N_24161);
nor U26005 (N_26005,N_25229,N_25368);
nand U26006 (N_26006,N_25151,N_24977);
and U26007 (N_26007,N_25462,N_24324);
and U26008 (N_26008,N_24889,N_24990);
nand U26009 (N_26009,N_24717,N_24599);
or U26010 (N_26010,N_24808,N_25436);
and U26011 (N_26011,N_25109,N_25375);
and U26012 (N_26012,N_24381,N_25237);
or U26013 (N_26013,N_24011,N_24833);
nor U26014 (N_26014,N_24137,N_25018);
xor U26015 (N_26015,N_24778,N_24588);
nand U26016 (N_26016,N_24057,N_24288);
xnor U26017 (N_26017,N_24320,N_24871);
and U26018 (N_26018,N_25480,N_24721);
or U26019 (N_26019,N_24571,N_24741);
nor U26020 (N_26020,N_24378,N_24727);
xor U26021 (N_26021,N_24287,N_24618);
or U26022 (N_26022,N_24167,N_25419);
and U26023 (N_26023,N_25190,N_24948);
nand U26024 (N_26024,N_25291,N_24817);
nor U26025 (N_26025,N_24099,N_24268);
nor U26026 (N_26026,N_24979,N_24225);
or U26027 (N_26027,N_25099,N_24439);
xnor U26028 (N_26028,N_24598,N_24261);
and U26029 (N_26029,N_24354,N_25456);
nor U26030 (N_26030,N_24515,N_24941);
nor U26031 (N_26031,N_24991,N_24897);
xor U26032 (N_26032,N_25131,N_24702);
or U26033 (N_26033,N_24670,N_25177);
or U26034 (N_26034,N_24146,N_24546);
or U26035 (N_26035,N_24987,N_25248);
or U26036 (N_26036,N_24666,N_24528);
nor U26037 (N_26037,N_25156,N_24567);
xor U26038 (N_26038,N_24296,N_24962);
and U26039 (N_26039,N_24342,N_24401);
xor U26040 (N_26040,N_25490,N_24992);
and U26041 (N_26041,N_25387,N_24578);
nor U26042 (N_26042,N_24530,N_24543);
nand U26043 (N_26043,N_24854,N_25344);
or U26044 (N_26044,N_25420,N_24043);
nand U26045 (N_26045,N_24498,N_24312);
nor U26046 (N_26046,N_25266,N_25329);
nand U26047 (N_26047,N_24894,N_24915);
nand U26048 (N_26048,N_24080,N_25372);
xor U26049 (N_26049,N_24901,N_25340);
nand U26050 (N_26050,N_24689,N_25363);
nor U26051 (N_26051,N_24120,N_24012);
or U26052 (N_26052,N_24259,N_24117);
xor U26053 (N_26053,N_24389,N_24541);
or U26054 (N_26054,N_24013,N_24976);
nand U26055 (N_26055,N_24457,N_25094);
nor U26056 (N_26056,N_24101,N_24791);
and U26057 (N_26057,N_24575,N_25483);
xor U26058 (N_26058,N_24876,N_24981);
and U26059 (N_26059,N_24958,N_25261);
xnor U26060 (N_26060,N_24232,N_24650);
and U26061 (N_26061,N_25082,N_24107);
nand U26062 (N_26062,N_25397,N_24202);
and U26063 (N_26063,N_24967,N_24510);
xnor U26064 (N_26064,N_25164,N_25335);
or U26065 (N_26065,N_24557,N_25025);
and U26066 (N_26066,N_24994,N_25452);
nand U26067 (N_26067,N_24456,N_24784);
and U26068 (N_26068,N_24538,N_25299);
nor U26069 (N_26069,N_24891,N_25236);
or U26070 (N_26070,N_24400,N_24442);
nor U26071 (N_26071,N_24376,N_24341);
or U26072 (N_26072,N_24014,N_24069);
nor U26073 (N_26073,N_24172,N_25143);
nand U26074 (N_26074,N_24671,N_24507);
and U26075 (N_26075,N_24249,N_25166);
nand U26076 (N_26076,N_25158,N_25493);
or U26077 (N_26077,N_24890,N_24245);
and U26078 (N_26078,N_24370,N_24570);
nand U26079 (N_26079,N_24792,N_24133);
and U26080 (N_26080,N_25410,N_25302);
nor U26081 (N_26081,N_24054,N_24210);
xnor U26082 (N_26082,N_24110,N_24279);
xnor U26083 (N_26083,N_24750,N_24758);
and U26084 (N_26084,N_24654,N_24934);
nor U26085 (N_26085,N_25016,N_24745);
nor U26086 (N_26086,N_24851,N_24807);
nand U26087 (N_26087,N_25284,N_25309);
nor U26088 (N_26088,N_25065,N_24703);
xnor U26089 (N_26089,N_24052,N_25214);
nor U26090 (N_26090,N_25086,N_25274);
nor U26091 (N_26091,N_24508,N_24649);
or U26092 (N_26092,N_24667,N_25390);
and U26093 (N_26093,N_24361,N_24942);
nand U26094 (N_26094,N_24051,N_24262);
nor U26095 (N_26095,N_25108,N_24999);
nor U26096 (N_26096,N_25009,N_24067);
and U26097 (N_26097,N_24780,N_24115);
nand U26098 (N_26098,N_24875,N_24170);
nor U26099 (N_26099,N_24687,N_25254);
nand U26100 (N_26100,N_25138,N_24001);
nor U26101 (N_26101,N_24626,N_24779);
or U26102 (N_26102,N_24448,N_24604);
xnor U26103 (N_26103,N_24231,N_24845);
nand U26104 (N_26104,N_25473,N_24754);
xor U26105 (N_26105,N_24944,N_24539);
xnor U26106 (N_26106,N_24733,N_25218);
and U26107 (N_26107,N_25411,N_24582);
or U26108 (N_26108,N_25262,N_24260);
nor U26109 (N_26109,N_24075,N_25400);
or U26110 (N_26110,N_24185,N_24412);
xnor U26111 (N_26111,N_25191,N_24373);
nand U26112 (N_26112,N_25015,N_25382);
or U26113 (N_26113,N_24384,N_25092);
xor U26114 (N_26114,N_25491,N_24058);
nor U26115 (N_26115,N_24964,N_25498);
nand U26116 (N_26116,N_24503,N_24685);
nand U26117 (N_26117,N_25360,N_24184);
and U26118 (N_26118,N_25163,N_25194);
nand U26119 (N_26119,N_24243,N_24552);
nand U26120 (N_26120,N_25315,N_24521);
or U26121 (N_26121,N_24056,N_24125);
and U26122 (N_26122,N_24452,N_25293);
nand U26123 (N_26123,N_24187,N_25026);
and U26124 (N_26124,N_24285,N_25162);
nor U26125 (N_26125,N_25120,N_24961);
nor U26126 (N_26126,N_24155,N_25224);
and U26127 (N_26127,N_24836,N_24985);
and U26128 (N_26128,N_24632,N_24914);
nor U26129 (N_26129,N_24204,N_24060);
xor U26130 (N_26130,N_24318,N_24105);
or U26131 (N_26131,N_24922,N_25378);
and U26132 (N_26132,N_24070,N_24783);
and U26133 (N_26133,N_25058,N_24437);
nor U26134 (N_26134,N_24847,N_24853);
or U26135 (N_26135,N_25053,N_24367);
xnor U26136 (N_26136,N_24905,N_25477);
nand U26137 (N_26137,N_24863,N_24048);
nor U26138 (N_26138,N_24829,N_24346);
xnor U26139 (N_26139,N_24251,N_24735);
nand U26140 (N_26140,N_24772,N_24789);
xnor U26141 (N_26141,N_24335,N_24881);
and U26142 (N_26142,N_25136,N_24432);
xnor U26143 (N_26143,N_25338,N_25330);
and U26144 (N_26144,N_24283,N_25451);
and U26145 (N_26145,N_24364,N_25277);
or U26146 (N_26146,N_24892,N_24595);
xnor U26147 (N_26147,N_24385,N_25476);
or U26148 (N_26148,N_25403,N_24732);
nand U26149 (N_26149,N_25222,N_25319);
or U26150 (N_26150,N_24235,N_24763);
nand U26151 (N_26151,N_24773,N_24920);
xor U26152 (N_26152,N_24636,N_25272);
nor U26153 (N_26153,N_25496,N_25394);
nor U26154 (N_26154,N_25485,N_24049);
or U26155 (N_26155,N_24611,N_24334);
xor U26156 (N_26156,N_24755,N_24234);
nand U26157 (N_26157,N_24953,N_24050);
nor U26158 (N_26158,N_24634,N_24332);
and U26159 (N_26159,N_24037,N_25114);
nand U26160 (N_26160,N_24909,N_24472);
or U26161 (N_26161,N_24397,N_24877);
xor U26162 (N_26162,N_24995,N_24887);
nand U26163 (N_26163,N_25130,N_24240);
nand U26164 (N_26164,N_24989,N_25057);
nand U26165 (N_26165,N_24487,N_25019);
and U26166 (N_26166,N_25321,N_24416);
nor U26167 (N_26167,N_25043,N_25377);
and U26168 (N_26168,N_25021,N_24290);
and U26169 (N_26169,N_24869,N_25482);
nand U26170 (N_26170,N_24321,N_25028);
nor U26171 (N_26171,N_25463,N_25061);
xnor U26172 (N_26172,N_24574,N_24214);
xor U26173 (N_26173,N_24781,N_25408);
or U26174 (N_26174,N_24138,N_24509);
nor U26175 (N_26175,N_25466,N_24837);
and U26176 (N_26176,N_25203,N_25215);
nor U26177 (N_26177,N_24297,N_25312);
and U26178 (N_26178,N_25475,N_24776);
and U26179 (N_26179,N_25369,N_24032);
xor U26180 (N_26180,N_25117,N_25470);
xor U26181 (N_26181,N_24464,N_24496);
and U26182 (N_26182,N_24699,N_24383);
and U26183 (N_26183,N_25038,N_24126);
nor U26184 (N_26184,N_25227,N_24263);
xnor U26185 (N_26185,N_24103,N_24410);
nor U26186 (N_26186,N_25418,N_24081);
xnor U26187 (N_26187,N_24009,N_24178);
or U26188 (N_26188,N_25472,N_24661);
nand U26189 (N_26189,N_25260,N_24500);
and U26190 (N_26190,N_24130,N_24594);
nand U26191 (N_26191,N_24104,N_24716);
xor U26192 (N_26192,N_25348,N_24760);
nand U26193 (N_26193,N_24968,N_24638);
xnor U26194 (N_26194,N_24608,N_24379);
or U26195 (N_26195,N_25105,N_25386);
and U26196 (N_26196,N_25313,N_24704);
nor U26197 (N_26197,N_24116,N_25076);
xor U26198 (N_26198,N_24902,N_24648);
xor U26199 (N_26199,N_24655,N_24859);
and U26200 (N_26200,N_24644,N_24898);
nor U26201 (N_26201,N_24257,N_24407);
nand U26202 (N_26202,N_24181,N_24770);
and U26203 (N_26203,N_24610,N_24201);
and U26204 (N_26204,N_24158,N_24002);
xnor U26205 (N_26205,N_25257,N_24021);
xor U26206 (N_26206,N_24278,N_24420);
xnor U26207 (N_26207,N_24819,N_25306);
and U26208 (N_26208,N_25155,N_24652);
and U26209 (N_26209,N_25353,N_25276);
or U26210 (N_26210,N_25059,N_25278);
xnor U26211 (N_26211,N_24421,N_25464);
nor U26212 (N_26212,N_24907,N_24109);
xor U26213 (N_26213,N_24640,N_24663);
and U26214 (N_26214,N_24264,N_24095);
or U26215 (N_26215,N_24445,N_24141);
nor U26216 (N_26216,N_24366,N_24466);
and U26217 (N_26217,N_24641,N_25285);
xnor U26218 (N_26218,N_25083,N_25180);
xnor U26219 (N_26219,N_24491,N_24124);
or U26220 (N_26220,N_24252,N_25125);
xor U26221 (N_26221,N_24493,N_25421);
nor U26222 (N_26222,N_25308,N_24071);
nand U26223 (N_26223,N_24023,N_24409);
and U26224 (N_26224,N_25113,N_24473);
nand U26225 (N_26225,N_24143,N_25075);
or U26226 (N_26226,N_24053,N_24430);
nand U26227 (N_26227,N_24089,N_24353);
nor U26228 (N_26228,N_24166,N_24426);
and U26229 (N_26229,N_24196,N_25055);
or U26230 (N_26230,N_24483,N_24616);
xor U26231 (N_26231,N_24026,N_24623);
nor U26232 (N_26232,N_24084,N_24256);
nand U26233 (N_26233,N_24372,N_25393);
xnor U26234 (N_26234,N_24696,N_25142);
nor U26235 (N_26235,N_24602,N_24729);
or U26236 (N_26236,N_25196,N_25247);
nor U26237 (N_26237,N_25326,N_24045);
nor U26238 (N_26238,N_24088,N_24534);
xor U26239 (N_26239,N_24337,N_25381);
nand U26240 (N_26240,N_24742,N_24912);
xnor U26241 (N_26241,N_24963,N_25323);
and U26242 (N_26242,N_25001,N_24572);
or U26243 (N_26243,N_25447,N_25354);
and U26244 (N_26244,N_25424,N_25433);
nand U26245 (N_26245,N_24676,N_25414);
and U26246 (N_26246,N_24577,N_24090);
nor U26247 (N_26247,N_24189,N_24449);
nor U26248 (N_26248,N_25388,N_25228);
and U26249 (N_26249,N_24284,N_24788);
nand U26250 (N_26250,N_24437,N_24704);
nand U26251 (N_26251,N_24147,N_25271);
and U26252 (N_26252,N_24281,N_24614);
or U26253 (N_26253,N_25032,N_24943);
nor U26254 (N_26254,N_24549,N_25004);
nor U26255 (N_26255,N_25480,N_24694);
xor U26256 (N_26256,N_24573,N_24715);
xor U26257 (N_26257,N_24270,N_25295);
xnor U26258 (N_26258,N_25190,N_25316);
nand U26259 (N_26259,N_25011,N_25074);
nand U26260 (N_26260,N_25442,N_25137);
or U26261 (N_26261,N_24237,N_24629);
xor U26262 (N_26262,N_25489,N_25337);
or U26263 (N_26263,N_25350,N_25210);
and U26264 (N_26264,N_24722,N_25055);
nand U26265 (N_26265,N_24857,N_24923);
or U26266 (N_26266,N_25215,N_25252);
nand U26267 (N_26267,N_24836,N_25388);
nand U26268 (N_26268,N_24263,N_24591);
or U26269 (N_26269,N_24462,N_24433);
nand U26270 (N_26270,N_25190,N_24273);
and U26271 (N_26271,N_24307,N_24533);
xnor U26272 (N_26272,N_24820,N_25006);
xnor U26273 (N_26273,N_24087,N_24945);
nor U26274 (N_26274,N_24857,N_25202);
nand U26275 (N_26275,N_24830,N_24221);
or U26276 (N_26276,N_25263,N_24574);
and U26277 (N_26277,N_25275,N_24171);
and U26278 (N_26278,N_24236,N_24239);
xor U26279 (N_26279,N_24042,N_24021);
xnor U26280 (N_26280,N_24092,N_24764);
nor U26281 (N_26281,N_24419,N_24703);
xnor U26282 (N_26282,N_24141,N_24129);
and U26283 (N_26283,N_24542,N_24125);
xor U26284 (N_26284,N_24535,N_25072);
or U26285 (N_26285,N_25121,N_25483);
nand U26286 (N_26286,N_25060,N_24582);
xnor U26287 (N_26287,N_24020,N_24960);
xnor U26288 (N_26288,N_24599,N_25158);
nor U26289 (N_26289,N_25034,N_24277);
xnor U26290 (N_26290,N_24090,N_24510);
and U26291 (N_26291,N_24954,N_25070);
xor U26292 (N_26292,N_24797,N_24929);
or U26293 (N_26293,N_24589,N_24001);
or U26294 (N_26294,N_24841,N_24423);
nor U26295 (N_26295,N_24687,N_24366);
nand U26296 (N_26296,N_24366,N_24619);
nor U26297 (N_26297,N_25210,N_25251);
and U26298 (N_26298,N_25158,N_24519);
nand U26299 (N_26299,N_24162,N_25038);
nand U26300 (N_26300,N_25160,N_24022);
xor U26301 (N_26301,N_24707,N_24606);
or U26302 (N_26302,N_24150,N_24790);
xnor U26303 (N_26303,N_24284,N_24713);
xor U26304 (N_26304,N_24313,N_24585);
nor U26305 (N_26305,N_24586,N_24515);
nor U26306 (N_26306,N_24880,N_24881);
xor U26307 (N_26307,N_24614,N_24443);
or U26308 (N_26308,N_25135,N_24101);
xor U26309 (N_26309,N_24754,N_24175);
or U26310 (N_26310,N_25137,N_24723);
nand U26311 (N_26311,N_25424,N_25050);
and U26312 (N_26312,N_24518,N_24481);
nand U26313 (N_26313,N_25404,N_24996);
and U26314 (N_26314,N_24929,N_24134);
nor U26315 (N_26315,N_24344,N_24229);
xnor U26316 (N_26316,N_24730,N_24137);
or U26317 (N_26317,N_24474,N_24842);
nor U26318 (N_26318,N_24332,N_24889);
nand U26319 (N_26319,N_24447,N_24609);
xor U26320 (N_26320,N_24687,N_24894);
nor U26321 (N_26321,N_24276,N_25034);
nor U26322 (N_26322,N_25231,N_24757);
nand U26323 (N_26323,N_24550,N_24570);
nor U26324 (N_26324,N_24698,N_25100);
and U26325 (N_26325,N_25066,N_24631);
xnor U26326 (N_26326,N_24260,N_24237);
xor U26327 (N_26327,N_24676,N_25181);
xor U26328 (N_26328,N_25357,N_24658);
nor U26329 (N_26329,N_24773,N_24605);
nor U26330 (N_26330,N_24138,N_24244);
nor U26331 (N_26331,N_24533,N_25288);
and U26332 (N_26332,N_24475,N_24529);
or U26333 (N_26333,N_24615,N_24573);
and U26334 (N_26334,N_25472,N_24802);
xor U26335 (N_26335,N_25391,N_25429);
and U26336 (N_26336,N_25423,N_24431);
nand U26337 (N_26337,N_24359,N_24196);
xnor U26338 (N_26338,N_24970,N_24497);
nand U26339 (N_26339,N_24339,N_24474);
and U26340 (N_26340,N_25002,N_24347);
nand U26341 (N_26341,N_24480,N_25368);
nor U26342 (N_26342,N_24194,N_24670);
nor U26343 (N_26343,N_24248,N_24942);
or U26344 (N_26344,N_24465,N_24554);
xnor U26345 (N_26345,N_24258,N_25241);
or U26346 (N_26346,N_24241,N_24137);
and U26347 (N_26347,N_25251,N_24710);
xnor U26348 (N_26348,N_25499,N_24961);
nand U26349 (N_26349,N_24139,N_24092);
or U26350 (N_26350,N_25432,N_25221);
xnor U26351 (N_26351,N_24405,N_24397);
nand U26352 (N_26352,N_25242,N_25498);
nor U26353 (N_26353,N_24360,N_24572);
nor U26354 (N_26354,N_24232,N_25223);
nand U26355 (N_26355,N_25094,N_24948);
and U26356 (N_26356,N_24210,N_24666);
and U26357 (N_26357,N_24368,N_24584);
nor U26358 (N_26358,N_24385,N_24948);
nand U26359 (N_26359,N_24227,N_24143);
xnor U26360 (N_26360,N_24288,N_25092);
and U26361 (N_26361,N_24627,N_25388);
xnor U26362 (N_26362,N_24301,N_24110);
and U26363 (N_26363,N_24266,N_24582);
and U26364 (N_26364,N_24156,N_24368);
nor U26365 (N_26365,N_24632,N_24575);
and U26366 (N_26366,N_24651,N_24309);
or U26367 (N_26367,N_25114,N_24203);
xor U26368 (N_26368,N_24597,N_25055);
nand U26369 (N_26369,N_24815,N_25325);
or U26370 (N_26370,N_24020,N_24914);
nor U26371 (N_26371,N_25422,N_24673);
nor U26372 (N_26372,N_25004,N_24196);
xor U26373 (N_26373,N_25385,N_24587);
or U26374 (N_26374,N_25181,N_24845);
xor U26375 (N_26375,N_24149,N_24917);
xnor U26376 (N_26376,N_24219,N_24508);
nand U26377 (N_26377,N_24440,N_25362);
nor U26378 (N_26378,N_25494,N_24852);
nor U26379 (N_26379,N_24281,N_24432);
nand U26380 (N_26380,N_25131,N_24759);
and U26381 (N_26381,N_24401,N_25428);
or U26382 (N_26382,N_24055,N_24348);
nand U26383 (N_26383,N_24265,N_24267);
xor U26384 (N_26384,N_25143,N_24877);
nor U26385 (N_26385,N_24834,N_25320);
or U26386 (N_26386,N_24198,N_25381);
and U26387 (N_26387,N_24904,N_25239);
or U26388 (N_26388,N_24428,N_24576);
or U26389 (N_26389,N_24793,N_24539);
or U26390 (N_26390,N_24635,N_24284);
nor U26391 (N_26391,N_25237,N_24443);
nand U26392 (N_26392,N_25313,N_25224);
and U26393 (N_26393,N_25371,N_24819);
nand U26394 (N_26394,N_24696,N_24841);
xnor U26395 (N_26395,N_24212,N_24107);
xor U26396 (N_26396,N_24173,N_25077);
nand U26397 (N_26397,N_24425,N_24233);
nor U26398 (N_26398,N_25489,N_24601);
and U26399 (N_26399,N_25283,N_24352);
nor U26400 (N_26400,N_24931,N_25244);
and U26401 (N_26401,N_24896,N_24420);
nand U26402 (N_26402,N_24284,N_25366);
xnor U26403 (N_26403,N_24610,N_24657);
and U26404 (N_26404,N_24287,N_25063);
nor U26405 (N_26405,N_24597,N_24258);
nor U26406 (N_26406,N_24387,N_25283);
nand U26407 (N_26407,N_25083,N_24935);
nand U26408 (N_26408,N_25096,N_24471);
or U26409 (N_26409,N_25198,N_24703);
and U26410 (N_26410,N_24365,N_24591);
xor U26411 (N_26411,N_25473,N_24675);
nand U26412 (N_26412,N_25069,N_24803);
nor U26413 (N_26413,N_24512,N_24499);
and U26414 (N_26414,N_25136,N_25261);
nand U26415 (N_26415,N_25349,N_25177);
nand U26416 (N_26416,N_24918,N_25082);
or U26417 (N_26417,N_24434,N_24989);
or U26418 (N_26418,N_24657,N_24386);
nor U26419 (N_26419,N_25032,N_25437);
and U26420 (N_26420,N_24361,N_24423);
or U26421 (N_26421,N_25105,N_24192);
or U26422 (N_26422,N_24869,N_24670);
nand U26423 (N_26423,N_24676,N_25096);
or U26424 (N_26424,N_24154,N_24141);
nand U26425 (N_26425,N_24282,N_25071);
nand U26426 (N_26426,N_25110,N_25210);
xnor U26427 (N_26427,N_24868,N_25083);
nor U26428 (N_26428,N_24882,N_25202);
nand U26429 (N_26429,N_24139,N_24785);
nand U26430 (N_26430,N_24759,N_24977);
or U26431 (N_26431,N_24411,N_25331);
xor U26432 (N_26432,N_24157,N_25060);
or U26433 (N_26433,N_24054,N_24739);
xor U26434 (N_26434,N_24964,N_25259);
nor U26435 (N_26435,N_24128,N_24743);
nand U26436 (N_26436,N_24853,N_25487);
nor U26437 (N_26437,N_24607,N_24867);
nand U26438 (N_26438,N_24984,N_24035);
nand U26439 (N_26439,N_24536,N_25450);
nand U26440 (N_26440,N_24345,N_24945);
and U26441 (N_26441,N_25177,N_24798);
or U26442 (N_26442,N_25388,N_24378);
and U26443 (N_26443,N_24409,N_24895);
nor U26444 (N_26444,N_24778,N_24232);
nand U26445 (N_26445,N_24793,N_25208);
nand U26446 (N_26446,N_24998,N_25454);
nand U26447 (N_26447,N_25218,N_25480);
nor U26448 (N_26448,N_24414,N_24309);
nand U26449 (N_26449,N_25118,N_24428);
nand U26450 (N_26450,N_24185,N_24357);
nand U26451 (N_26451,N_24000,N_24518);
xor U26452 (N_26452,N_24217,N_24223);
xor U26453 (N_26453,N_24934,N_24017);
nand U26454 (N_26454,N_24913,N_24805);
nor U26455 (N_26455,N_25183,N_25424);
xnor U26456 (N_26456,N_25073,N_25317);
nor U26457 (N_26457,N_24479,N_24789);
xor U26458 (N_26458,N_25220,N_24056);
and U26459 (N_26459,N_24581,N_24819);
and U26460 (N_26460,N_25014,N_24791);
or U26461 (N_26461,N_25074,N_25130);
nor U26462 (N_26462,N_24886,N_25397);
and U26463 (N_26463,N_25448,N_24287);
nor U26464 (N_26464,N_25295,N_25492);
nor U26465 (N_26465,N_24305,N_24184);
and U26466 (N_26466,N_24319,N_25411);
xor U26467 (N_26467,N_25323,N_24835);
nand U26468 (N_26468,N_24970,N_24771);
nand U26469 (N_26469,N_24276,N_25176);
or U26470 (N_26470,N_24660,N_24425);
xor U26471 (N_26471,N_24049,N_25198);
and U26472 (N_26472,N_25175,N_24809);
xor U26473 (N_26473,N_24618,N_25269);
nand U26474 (N_26474,N_24840,N_24675);
nand U26475 (N_26475,N_24612,N_24902);
xnor U26476 (N_26476,N_24672,N_24158);
and U26477 (N_26477,N_25295,N_24676);
and U26478 (N_26478,N_24730,N_24778);
and U26479 (N_26479,N_24560,N_24152);
nand U26480 (N_26480,N_25030,N_24382);
nand U26481 (N_26481,N_25484,N_25321);
nor U26482 (N_26482,N_24106,N_24597);
nor U26483 (N_26483,N_24472,N_24340);
and U26484 (N_26484,N_24065,N_24640);
nand U26485 (N_26485,N_24216,N_24821);
or U26486 (N_26486,N_24722,N_24883);
or U26487 (N_26487,N_25062,N_24441);
xnor U26488 (N_26488,N_25394,N_24550);
nand U26489 (N_26489,N_24591,N_24290);
or U26490 (N_26490,N_24161,N_25071);
nand U26491 (N_26491,N_24446,N_24790);
nor U26492 (N_26492,N_24953,N_24767);
and U26493 (N_26493,N_24027,N_25265);
nor U26494 (N_26494,N_24957,N_25156);
xor U26495 (N_26495,N_24138,N_25135);
nand U26496 (N_26496,N_25197,N_24663);
or U26497 (N_26497,N_25483,N_24629);
and U26498 (N_26498,N_25092,N_24897);
xnor U26499 (N_26499,N_24979,N_25388);
or U26500 (N_26500,N_25387,N_24515);
and U26501 (N_26501,N_24282,N_24797);
xnor U26502 (N_26502,N_25089,N_24316);
nand U26503 (N_26503,N_24695,N_24978);
and U26504 (N_26504,N_24066,N_25224);
xor U26505 (N_26505,N_25389,N_24308);
nand U26506 (N_26506,N_25003,N_24648);
or U26507 (N_26507,N_24587,N_24629);
and U26508 (N_26508,N_24755,N_24407);
xor U26509 (N_26509,N_25159,N_24845);
nor U26510 (N_26510,N_24670,N_24221);
nand U26511 (N_26511,N_25164,N_25418);
and U26512 (N_26512,N_24049,N_24498);
nand U26513 (N_26513,N_24647,N_24994);
or U26514 (N_26514,N_24935,N_24810);
xor U26515 (N_26515,N_24560,N_25390);
or U26516 (N_26516,N_25411,N_25144);
and U26517 (N_26517,N_24268,N_24124);
xnor U26518 (N_26518,N_24256,N_25183);
nor U26519 (N_26519,N_25219,N_25152);
and U26520 (N_26520,N_24510,N_24665);
nand U26521 (N_26521,N_24008,N_24495);
xor U26522 (N_26522,N_24492,N_24531);
and U26523 (N_26523,N_24257,N_24296);
or U26524 (N_26524,N_24958,N_25219);
nand U26525 (N_26525,N_24800,N_24496);
or U26526 (N_26526,N_24784,N_25397);
nand U26527 (N_26527,N_24474,N_25192);
or U26528 (N_26528,N_24821,N_24656);
or U26529 (N_26529,N_24471,N_25255);
and U26530 (N_26530,N_24494,N_25458);
nand U26531 (N_26531,N_25181,N_24415);
or U26532 (N_26532,N_24671,N_24327);
and U26533 (N_26533,N_24206,N_24202);
or U26534 (N_26534,N_24486,N_25381);
nor U26535 (N_26535,N_24652,N_24019);
xor U26536 (N_26536,N_25157,N_24401);
nand U26537 (N_26537,N_25183,N_24240);
nand U26538 (N_26538,N_25249,N_24398);
and U26539 (N_26539,N_24976,N_24943);
nand U26540 (N_26540,N_25428,N_24857);
and U26541 (N_26541,N_24073,N_25356);
xor U26542 (N_26542,N_25022,N_25260);
nor U26543 (N_26543,N_25160,N_24369);
and U26544 (N_26544,N_24463,N_24159);
nor U26545 (N_26545,N_24850,N_24005);
nand U26546 (N_26546,N_24567,N_24154);
xor U26547 (N_26547,N_24983,N_24677);
xnor U26548 (N_26548,N_25183,N_25389);
nor U26549 (N_26549,N_25418,N_24949);
xnor U26550 (N_26550,N_25371,N_24668);
nor U26551 (N_26551,N_24335,N_24679);
and U26552 (N_26552,N_25109,N_25314);
and U26553 (N_26553,N_24449,N_24377);
nand U26554 (N_26554,N_24500,N_24911);
nand U26555 (N_26555,N_25276,N_24214);
xor U26556 (N_26556,N_25306,N_24561);
nand U26557 (N_26557,N_25050,N_24605);
nor U26558 (N_26558,N_25011,N_25433);
nor U26559 (N_26559,N_25430,N_24648);
nor U26560 (N_26560,N_25151,N_25419);
xor U26561 (N_26561,N_24799,N_25323);
nor U26562 (N_26562,N_24938,N_24688);
nand U26563 (N_26563,N_24385,N_24222);
or U26564 (N_26564,N_25364,N_24701);
nor U26565 (N_26565,N_25115,N_24271);
or U26566 (N_26566,N_25389,N_24980);
xnor U26567 (N_26567,N_25491,N_24505);
xnor U26568 (N_26568,N_25472,N_24233);
and U26569 (N_26569,N_24286,N_24376);
nand U26570 (N_26570,N_25319,N_24781);
nand U26571 (N_26571,N_24005,N_25300);
xor U26572 (N_26572,N_24561,N_24197);
nor U26573 (N_26573,N_24430,N_24114);
xnor U26574 (N_26574,N_24382,N_25356);
nand U26575 (N_26575,N_24996,N_24386);
xnor U26576 (N_26576,N_24577,N_25305);
nand U26577 (N_26577,N_24434,N_24840);
nor U26578 (N_26578,N_25405,N_25086);
and U26579 (N_26579,N_24522,N_24031);
nor U26580 (N_26580,N_24207,N_24816);
nand U26581 (N_26581,N_24557,N_25070);
and U26582 (N_26582,N_24070,N_24490);
and U26583 (N_26583,N_25194,N_24481);
and U26584 (N_26584,N_24960,N_24732);
xor U26585 (N_26585,N_24957,N_25033);
and U26586 (N_26586,N_24837,N_25162);
and U26587 (N_26587,N_24371,N_24150);
and U26588 (N_26588,N_24350,N_25173);
or U26589 (N_26589,N_24665,N_25142);
nand U26590 (N_26590,N_25376,N_24681);
nand U26591 (N_26591,N_24255,N_24904);
nor U26592 (N_26592,N_25219,N_25436);
or U26593 (N_26593,N_24098,N_24264);
xor U26594 (N_26594,N_24886,N_24049);
nand U26595 (N_26595,N_25267,N_25140);
or U26596 (N_26596,N_24774,N_24482);
or U26597 (N_26597,N_25043,N_24949);
and U26598 (N_26598,N_24139,N_25430);
nor U26599 (N_26599,N_25088,N_24021);
and U26600 (N_26600,N_24462,N_24691);
or U26601 (N_26601,N_25304,N_24651);
nor U26602 (N_26602,N_24375,N_25133);
and U26603 (N_26603,N_24299,N_25423);
or U26604 (N_26604,N_24378,N_24837);
and U26605 (N_26605,N_24122,N_24354);
and U26606 (N_26606,N_24402,N_24756);
or U26607 (N_26607,N_24907,N_24782);
nor U26608 (N_26608,N_24979,N_24355);
nor U26609 (N_26609,N_24074,N_24663);
or U26610 (N_26610,N_24169,N_24408);
nand U26611 (N_26611,N_25003,N_24314);
and U26612 (N_26612,N_24500,N_25065);
nand U26613 (N_26613,N_24092,N_25274);
and U26614 (N_26614,N_24633,N_24456);
nand U26615 (N_26615,N_25439,N_25402);
nand U26616 (N_26616,N_24073,N_25441);
nand U26617 (N_26617,N_24881,N_25261);
nand U26618 (N_26618,N_25139,N_25096);
xnor U26619 (N_26619,N_25087,N_24284);
nand U26620 (N_26620,N_24153,N_24861);
or U26621 (N_26621,N_24436,N_24320);
xor U26622 (N_26622,N_25158,N_24101);
or U26623 (N_26623,N_24817,N_25375);
nor U26624 (N_26624,N_24983,N_24841);
or U26625 (N_26625,N_24533,N_24414);
nand U26626 (N_26626,N_25371,N_24315);
nand U26627 (N_26627,N_24430,N_24658);
and U26628 (N_26628,N_24111,N_25014);
xor U26629 (N_26629,N_25057,N_24977);
nor U26630 (N_26630,N_24484,N_24235);
and U26631 (N_26631,N_24301,N_24094);
nor U26632 (N_26632,N_24063,N_24625);
and U26633 (N_26633,N_25466,N_25143);
xor U26634 (N_26634,N_25276,N_24777);
or U26635 (N_26635,N_24481,N_24536);
nor U26636 (N_26636,N_24371,N_24886);
nand U26637 (N_26637,N_24794,N_24823);
and U26638 (N_26638,N_24822,N_24554);
xnor U26639 (N_26639,N_24613,N_24394);
nor U26640 (N_26640,N_24879,N_25173);
and U26641 (N_26641,N_24618,N_25034);
and U26642 (N_26642,N_24710,N_24775);
xnor U26643 (N_26643,N_24851,N_24008);
xor U26644 (N_26644,N_25217,N_24945);
and U26645 (N_26645,N_24124,N_24769);
xor U26646 (N_26646,N_24948,N_24370);
and U26647 (N_26647,N_24816,N_25120);
or U26648 (N_26648,N_25473,N_25281);
xnor U26649 (N_26649,N_24994,N_24517);
xor U26650 (N_26650,N_24682,N_24408);
nor U26651 (N_26651,N_24256,N_24417);
or U26652 (N_26652,N_25052,N_24774);
nor U26653 (N_26653,N_24045,N_24812);
and U26654 (N_26654,N_25244,N_24246);
nand U26655 (N_26655,N_25370,N_24417);
or U26656 (N_26656,N_24341,N_24206);
and U26657 (N_26657,N_24339,N_24680);
xor U26658 (N_26658,N_25234,N_25449);
nand U26659 (N_26659,N_24123,N_24690);
nand U26660 (N_26660,N_24571,N_24301);
nor U26661 (N_26661,N_24332,N_25227);
nor U26662 (N_26662,N_24333,N_24211);
nand U26663 (N_26663,N_24221,N_25248);
or U26664 (N_26664,N_24280,N_24996);
nor U26665 (N_26665,N_24477,N_24507);
or U26666 (N_26666,N_25286,N_25382);
xnor U26667 (N_26667,N_24788,N_25390);
and U26668 (N_26668,N_24694,N_24597);
nor U26669 (N_26669,N_24801,N_24779);
or U26670 (N_26670,N_24086,N_24923);
and U26671 (N_26671,N_24772,N_24295);
nor U26672 (N_26672,N_25271,N_24177);
xnor U26673 (N_26673,N_25123,N_24615);
nand U26674 (N_26674,N_24856,N_24717);
and U26675 (N_26675,N_24198,N_24344);
nand U26676 (N_26676,N_24029,N_24192);
and U26677 (N_26677,N_24274,N_24819);
xnor U26678 (N_26678,N_24397,N_25074);
and U26679 (N_26679,N_24976,N_24502);
xor U26680 (N_26680,N_24335,N_24271);
nand U26681 (N_26681,N_24892,N_24755);
and U26682 (N_26682,N_24030,N_24089);
nor U26683 (N_26683,N_24638,N_24000);
nor U26684 (N_26684,N_24541,N_25366);
or U26685 (N_26685,N_24352,N_25389);
or U26686 (N_26686,N_24870,N_24337);
nand U26687 (N_26687,N_24636,N_24040);
xor U26688 (N_26688,N_24783,N_24268);
or U26689 (N_26689,N_24005,N_24337);
and U26690 (N_26690,N_24063,N_25101);
and U26691 (N_26691,N_24710,N_24055);
and U26692 (N_26692,N_24905,N_24930);
or U26693 (N_26693,N_25253,N_25318);
nand U26694 (N_26694,N_24399,N_25406);
nor U26695 (N_26695,N_24194,N_25439);
and U26696 (N_26696,N_24731,N_25062);
and U26697 (N_26697,N_24056,N_24495);
or U26698 (N_26698,N_24471,N_24174);
or U26699 (N_26699,N_24730,N_25223);
nand U26700 (N_26700,N_25212,N_24105);
or U26701 (N_26701,N_25023,N_24418);
nor U26702 (N_26702,N_24159,N_25164);
nor U26703 (N_26703,N_24168,N_24847);
nand U26704 (N_26704,N_24130,N_24898);
nor U26705 (N_26705,N_25139,N_24531);
or U26706 (N_26706,N_24047,N_24572);
or U26707 (N_26707,N_24421,N_25216);
or U26708 (N_26708,N_24029,N_24352);
and U26709 (N_26709,N_24074,N_24850);
and U26710 (N_26710,N_24108,N_25367);
and U26711 (N_26711,N_25402,N_24101);
nor U26712 (N_26712,N_24131,N_25429);
xnor U26713 (N_26713,N_24040,N_25472);
or U26714 (N_26714,N_25112,N_24616);
nand U26715 (N_26715,N_24616,N_24262);
nand U26716 (N_26716,N_24526,N_24127);
nand U26717 (N_26717,N_25073,N_25204);
nor U26718 (N_26718,N_24468,N_24910);
nor U26719 (N_26719,N_24299,N_24220);
or U26720 (N_26720,N_24225,N_24692);
xnor U26721 (N_26721,N_24334,N_24442);
nand U26722 (N_26722,N_24361,N_24299);
nand U26723 (N_26723,N_24537,N_24673);
xor U26724 (N_26724,N_24167,N_24153);
or U26725 (N_26725,N_24749,N_24395);
and U26726 (N_26726,N_24109,N_25174);
or U26727 (N_26727,N_24017,N_24804);
xor U26728 (N_26728,N_24381,N_25186);
nor U26729 (N_26729,N_24432,N_25132);
nor U26730 (N_26730,N_24192,N_25361);
xnor U26731 (N_26731,N_24924,N_24121);
and U26732 (N_26732,N_25347,N_25455);
nand U26733 (N_26733,N_24318,N_25359);
nand U26734 (N_26734,N_24554,N_24143);
and U26735 (N_26735,N_25445,N_24878);
nand U26736 (N_26736,N_24662,N_24456);
xor U26737 (N_26737,N_25307,N_24266);
xnor U26738 (N_26738,N_24213,N_25390);
nand U26739 (N_26739,N_25130,N_25412);
and U26740 (N_26740,N_24624,N_24959);
nand U26741 (N_26741,N_24402,N_24384);
and U26742 (N_26742,N_24127,N_25432);
nor U26743 (N_26743,N_24039,N_24661);
and U26744 (N_26744,N_24436,N_24328);
nand U26745 (N_26745,N_25257,N_25046);
nand U26746 (N_26746,N_25457,N_24043);
nor U26747 (N_26747,N_24019,N_25439);
nand U26748 (N_26748,N_24691,N_24957);
or U26749 (N_26749,N_24727,N_24892);
xnor U26750 (N_26750,N_24803,N_24026);
and U26751 (N_26751,N_24469,N_25391);
xnor U26752 (N_26752,N_24143,N_24841);
or U26753 (N_26753,N_25226,N_24984);
xnor U26754 (N_26754,N_24033,N_24714);
or U26755 (N_26755,N_24770,N_25064);
or U26756 (N_26756,N_24874,N_25049);
xnor U26757 (N_26757,N_24883,N_24885);
xnor U26758 (N_26758,N_24528,N_24158);
or U26759 (N_26759,N_25060,N_24831);
xnor U26760 (N_26760,N_24329,N_25250);
or U26761 (N_26761,N_24777,N_24893);
nand U26762 (N_26762,N_25455,N_24907);
xnor U26763 (N_26763,N_24832,N_25013);
nand U26764 (N_26764,N_24055,N_25123);
nor U26765 (N_26765,N_25071,N_25002);
or U26766 (N_26766,N_25087,N_24489);
nor U26767 (N_26767,N_24441,N_24307);
xor U26768 (N_26768,N_25351,N_24448);
nand U26769 (N_26769,N_24908,N_25036);
and U26770 (N_26770,N_24324,N_24932);
and U26771 (N_26771,N_25080,N_24975);
or U26772 (N_26772,N_24704,N_24601);
nand U26773 (N_26773,N_24906,N_25247);
or U26774 (N_26774,N_25446,N_24444);
and U26775 (N_26775,N_24903,N_24015);
nor U26776 (N_26776,N_24043,N_24796);
and U26777 (N_26777,N_25320,N_25080);
nor U26778 (N_26778,N_24610,N_24644);
xnor U26779 (N_26779,N_25426,N_24837);
xnor U26780 (N_26780,N_25237,N_24877);
nor U26781 (N_26781,N_25006,N_24694);
or U26782 (N_26782,N_25365,N_24108);
and U26783 (N_26783,N_24190,N_24262);
nor U26784 (N_26784,N_25030,N_24808);
or U26785 (N_26785,N_25361,N_25400);
xnor U26786 (N_26786,N_24547,N_24276);
or U26787 (N_26787,N_24808,N_25217);
nand U26788 (N_26788,N_24649,N_24014);
nor U26789 (N_26789,N_25305,N_24423);
xor U26790 (N_26790,N_25395,N_25333);
or U26791 (N_26791,N_25007,N_24706);
or U26792 (N_26792,N_25228,N_24984);
or U26793 (N_26793,N_25235,N_24398);
nor U26794 (N_26794,N_25371,N_24158);
xor U26795 (N_26795,N_24195,N_24491);
xnor U26796 (N_26796,N_24148,N_24166);
nor U26797 (N_26797,N_24767,N_24726);
nor U26798 (N_26798,N_24228,N_25159);
xor U26799 (N_26799,N_25348,N_24639);
xnor U26800 (N_26800,N_24986,N_24600);
nor U26801 (N_26801,N_24378,N_24585);
nor U26802 (N_26802,N_25038,N_24539);
nor U26803 (N_26803,N_25438,N_24573);
xnor U26804 (N_26804,N_24520,N_24227);
nor U26805 (N_26805,N_24974,N_24383);
and U26806 (N_26806,N_25234,N_24757);
nor U26807 (N_26807,N_24124,N_25223);
or U26808 (N_26808,N_24226,N_24005);
or U26809 (N_26809,N_24769,N_24167);
nor U26810 (N_26810,N_25077,N_24797);
or U26811 (N_26811,N_24950,N_24615);
xor U26812 (N_26812,N_24377,N_24066);
or U26813 (N_26813,N_24539,N_24912);
nor U26814 (N_26814,N_25469,N_25365);
nor U26815 (N_26815,N_25253,N_24131);
and U26816 (N_26816,N_24624,N_25080);
nor U26817 (N_26817,N_24642,N_24689);
nand U26818 (N_26818,N_24147,N_24808);
and U26819 (N_26819,N_25058,N_25104);
and U26820 (N_26820,N_25460,N_24136);
xor U26821 (N_26821,N_24595,N_24078);
xnor U26822 (N_26822,N_24066,N_24457);
and U26823 (N_26823,N_25319,N_25461);
nor U26824 (N_26824,N_24537,N_25408);
and U26825 (N_26825,N_24920,N_25002);
and U26826 (N_26826,N_24391,N_24721);
or U26827 (N_26827,N_24930,N_24898);
or U26828 (N_26828,N_25074,N_24633);
and U26829 (N_26829,N_24192,N_24326);
xnor U26830 (N_26830,N_24329,N_24034);
or U26831 (N_26831,N_25213,N_25356);
or U26832 (N_26832,N_24878,N_24315);
and U26833 (N_26833,N_24834,N_25352);
nand U26834 (N_26834,N_24048,N_24525);
xnor U26835 (N_26835,N_24230,N_24465);
nor U26836 (N_26836,N_24814,N_24360);
xor U26837 (N_26837,N_24543,N_24898);
and U26838 (N_26838,N_24596,N_24192);
nand U26839 (N_26839,N_25236,N_24219);
nor U26840 (N_26840,N_24955,N_25348);
xnor U26841 (N_26841,N_25040,N_24614);
or U26842 (N_26842,N_24092,N_24124);
and U26843 (N_26843,N_24548,N_25159);
or U26844 (N_26844,N_24451,N_24460);
nand U26845 (N_26845,N_24678,N_25316);
xor U26846 (N_26846,N_24582,N_24694);
nor U26847 (N_26847,N_24968,N_25238);
nand U26848 (N_26848,N_24800,N_24674);
xor U26849 (N_26849,N_25111,N_25384);
nand U26850 (N_26850,N_25320,N_24479);
or U26851 (N_26851,N_25350,N_24761);
nand U26852 (N_26852,N_24686,N_24646);
xor U26853 (N_26853,N_24117,N_24451);
nor U26854 (N_26854,N_24859,N_24438);
and U26855 (N_26855,N_24139,N_24905);
nand U26856 (N_26856,N_24942,N_24866);
or U26857 (N_26857,N_24246,N_24432);
or U26858 (N_26858,N_25372,N_24038);
xnor U26859 (N_26859,N_24750,N_25085);
or U26860 (N_26860,N_24246,N_25093);
nand U26861 (N_26861,N_24025,N_24640);
and U26862 (N_26862,N_24893,N_24852);
nand U26863 (N_26863,N_24171,N_24179);
or U26864 (N_26864,N_25092,N_24260);
or U26865 (N_26865,N_24949,N_24479);
xnor U26866 (N_26866,N_24327,N_24464);
nor U26867 (N_26867,N_24882,N_25183);
or U26868 (N_26868,N_25261,N_24540);
and U26869 (N_26869,N_24306,N_24354);
or U26870 (N_26870,N_24547,N_24009);
nand U26871 (N_26871,N_24426,N_25481);
and U26872 (N_26872,N_24971,N_25429);
nor U26873 (N_26873,N_25411,N_24396);
nor U26874 (N_26874,N_24346,N_25365);
xor U26875 (N_26875,N_24277,N_24955);
and U26876 (N_26876,N_24185,N_24007);
and U26877 (N_26877,N_24312,N_24715);
nand U26878 (N_26878,N_25026,N_25265);
xnor U26879 (N_26879,N_24393,N_24955);
xor U26880 (N_26880,N_24288,N_24893);
or U26881 (N_26881,N_24973,N_25064);
or U26882 (N_26882,N_25312,N_24007);
nor U26883 (N_26883,N_25309,N_25232);
nand U26884 (N_26884,N_25376,N_25487);
nor U26885 (N_26885,N_24954,N_24643);
nand U26886 (N_26886,N_24037,N_25087);
xor U26887 (N_26887,N_24418,N_24429);
or U26888 (N_26888,N_24305,N_24520);
nand U26889 (N_26889,N_25009,N_25325);
nor U26890 (N_26890,N_24623,N_24892);
nor U26891 (N_26891,N_25093,N_25358);
xor U26892 (N_26892,N_24125,N_25083);
xnor U26893 (N_26893,N_24683,N_24488);
nand U26894 (N_26894,N_24618,N_25175);
nor U26895 (N_26895,N_25468,N_24900);
or U26896 (N_26896,N_24236,N_24813);
and U26897 (N_26897,N_24204,N_24172);
or U26898 (N_26898,N_25101,N_24555);
nand U26899 (N_26899,N_24394,N_24548);
nand U26900 (N_26900,N_25052,N_25050);
nand U26901 (N_26901,N_24633,N_25318);
and U26902 (N_26902,N_24116,N_24373);
nor U26903 (N_26903,N_24771,N_24688);
nor U26904 (N_26904,N_24215,N_25161);
and U26905 (N_26905,N_24504,N_24462);
nand U26906 (N_26906,N_24948,N_24665);
and U26907 (N_26907,N_24705,N_24183);
nand U26908 (N_26908,N_24029,N_25083);
and U26909 (N_26909,N_24260,N_25343);
and U26910 (N_26910,N_25382,N_25171);
nand U26911 (N_26911,N_24427,N_25157);
and U26912 (N_26912,N_24308,N_24866);
and U26913 (N_26913,N_24469,N_24798);
or U26914 (N_26914,N_25242,N_24516);
nand U26915 (N_26915,N_24547,N_25018);
nor U26916 (N_26916,N_25218,N_24990);
xnor U26917 (N_26917,N_24288,N_25298);
or U26918 (N_26918,N_24014,N_25347);
nor U26919 (N_26919,N_24721,N_25016);
nand U26920 (N_26920,N_25314,N_24340);
nor U26921 (N_26921,N_24653,N_24136);
nand U26922 (N_26922,N_24046,N_24088);
or U26923 (N_26923,N_25104,N_24589);
xnor U26924 (N_26924,N_24114,N_25211);
nor U26925 (N_26925,N_25461,N_24287);
and U26926 (N_26926,N_25438,N_25029);
and U26927 (N_26927,N_24394,N_25304);
and U26928 (N_26928,N_25374,N_24083);
and U26929 (N_26929,N_25147,N_24695);
or U26930 (N_26930,N_24212,N_24434);
or U26931 (N_26931,N_25457,N_24638);
or U26932 (N_26932,N_25296,N_24870);
xor U26933 (N_26933,N_25478,N_24034);
or U26934 (N_26934,N_24731,N_24003);
xor U26935 (N_26935,N_24843,N_24870);
nor U26936 (N_26936,N_24361,N_24160);
or U26937 (N_26937,N_24554,N_24284);
xor U26938 (N_26938,N_25373,N_24986);
or U26939 (N_26939,N_24875,N_24006);
xnor U26940 (N_26940,N_24938,N_24736);
nand U26941 (N_26941,N_24820,N_24355);
and U26942 (N_26942,N_25105,N_24433);
nand U26943 (N_26943,N_24925,N_24295);
or U26944 (N_26944,N_24037,N_25203);
nand U26945 (N_26945,N_24571,N_24097);
xnor U26946 (N_26946,N_24310,N_24223);
nand U26947 (N_26947,N_24577,N_24946);
and U26948 (N_26948,N_25120,N_24586);
nor U26949 (N_26949,N_24914,N_24278);
xor U26950 (N_26950,N_24849,N_24394);
and U26951 (N_26951,N_24047,N_25373);
or U26952 (N_26952,N_24504,N_25263);
and U26953 (N_26953,N_24847,N_24771);
or U26954 (N_26954,N_24753,N_25216);
nor U26955 (N_26955,N_24202,N_24338);
xnor U26956 (N_26956,N_24127,N_24373);
and U26957 (N_26957,N_25372,N_24680);
and U26958 (N_26958,N_25102,N_24310);
nor U26959 (N_26959,N_25331,N_24724);
nand U26960 (N_26960,N_24050,N_24389);
nand U26961 (N_26961,N_25476,N_24595);
nor U26962 (N_26962,N_25464,N_25215);
xor U26963 (N_26963,N_24706,N_24707);
or U26964 (N_26964,N_25102,N_24702);
and U26965 (N_26965,N_25038,N_25239);
and U26966 (N_26966,N_25446,N_25456);
nor U26967 (N_26967,N_24097,N_24895);
nand U26968 (N_26968,N_25315,N_24763);
nor U26969 (N_26969,N_25053,N_24991);
xor U26970 (N_26970,N_24941,N_24678);
nand U26971 (N_26971,N_25317,N_25270);
nor U26972 (N_26972,N_25308,N_24626);
and U26973 (N_26973,N_25388,N_24153);
nor U26974 (N_26974,N_25216,N_24235);
xnor U26975 (N_26975,N_25131,N_25175);
nand U26976 (N_26976,N_24104,N_24070);
nand U26977 (N_26977,N_24783,N_24945);
or U26978 (N_26978,N_24387,N_24956);
xor U26979 (N_26979,N_25497,N_25283);
nand U26980 (N_26980,N_24682,N_25086);
or U26981 (N_26981,N_24408,N_24089);
or U26982 (N_26982,N_25113,N_25450);
or U26983 (N_26983,N_24158,N_24588);
nand U26984 (N_26984,N_25314,N_24172);
or U26985 (N_26985,N_24928,N_24878);
xnor U26986 (N_26986,N_24104,N_24167);
and U26987 (N_26987,N_24687,N_25282);
and U26988 (N_26988,N_24248,N_24281);
nand U26989 (N_26989,N_24312,N_24472);
xor U26990 (N_26990,N_24975,N_24427);
nor U26991 (N_26991,N_24329,N_24212);
xor U26992 (N_26992,N_24321,N_25046);
xnor U26993 (N_26993,N_24172,N_25100);
nand U26994 (N_26994,N_24833,N_24132);
nor U26995 (N_26995,N_25063,N_24165);
nand U26996 (N_26996,N_25294,N_24406);
nand U26997 (N_26997,N_24678,N_25482);
nand U26998 (N_26998,N_24989,N_24296);
nor U26999 (N_26999,N_25174,N_24248);
nand U27000 (N_27000,N_26163,N_26614);
and U27001 (N_27001,N_26102,N_25884);
or U27002 (N_27002,N_26397,N_25876);
nor U27003 (N_27003,N_26269,N_26564);
nor U27004 (N_27004,N_26537,N_26446);
xor U27005 (N_27005,N_26516,N_25956);
or U27006 (N_27006,N_26636,N_25631);
and U27007 (N_27007,N_25777,N_26245);
nand U27008 (N_27008,N_26070,N_26903);
xnor U27009 (N_27009,N_26561,N_26222);
nand U27010 (N_27010,N_26525,N_26773);
nor U27011 (N_27011,N_26183,N_25549);
and U27012 (N_27012,N_26557,N_25961);
nand U27013 (N_27013,N_26615,N_25521);
and U27014 (N_27014,N_26059,N_26954);
or U27015 (N_27015,N_25730,N_26483);
nor U27016 (N_27016,N_26191,N_26410);
nand U27017 (N_27017,N_26423,N_26385);
or U27018 (N_27018,N_25656,N_26538);
or U27019 (N_27019,N_25909,N_26902);
or U27020 (N_27020,N_26644,N_25646);
and U27021 (N_27021,N_26330,N_25558);
nand U27022 (N_27022,N_26719,N_26379);
and U27023 (N_27023,N_26603,N_25654);
nor U27024 (N_27024,N_26608,N_26599);
nand U27025 (N_27025,N_26866,N_25574);
xor U27026 (N_27026,N_26002,N_26743);
xor U27027 (N_27027,N_26343,N_26863);
nor U27028 (N_27028,N_26649,N_26710);
nand U27029 (N_27029,N_26154,N_25515);
xor U27030 (N_27030,N_26577,N_26788);
xnor U27031 (N_27031,N_26237,N_26306);
nor U27032 (N_27032,N_26654,N_25893);
nor U27033 (N_27033,N_26819,N_26852);
xnor U27034 (N_27034,N_25925,N_25670);
and U27035 (N_27035,N_26873,N_25568);
nor U27036 (N_27036,N_26856,N_25946);
nor U27037 (N_27037,N_26673,N_26253);
nor U27038 (N_27038,N_26075,N_26167);
and U27039 (N_27039,N_26161,N_26254);
or U27040 (N_27040,N_26030,N_26203);
nor U27041 (N_27041,N_26581,N_25921);
nand U27042 (N_27042,N_26575,N_26045);
nand U27043 (N_27043,N_26079,N_26211);
nand U27044 (N_27044,N_25836,N_26630);
and U27045 (N_27045,N_26833,N_26309);
and U27046 (N_27046,N_25958,N_26929);
or U27047 (N_27047,N_26701,N_25557);
and U27048 (N_27048,N_25570,N_26052);
or U27049 (N_27049,N_26248,N_25583);
or U27050 (N_27050,N_26946,N_25600);
xnor U27051 (N_27051,N_26375,N_26150);
nand U27052 (N_27052,N_26486,N_26541);
xor U27053 (N_27053,N_25529,N_26996);
or U27054 (N_27054,N_26641,N_25863);
or U27055 (N_27055,N_25704,N_26249);
and U27056 (N_27056,N_25805,N_25639);
nand U27057 (N_27057,N_26590,N_26979);
or U27058 (N_27058,N_25957,N_25765);
xor U27059 (N_27059,N_26421,N_26126);
or U27060 (N_27060,N_26589,N_25533);
and U27061 (N_27061,N_26036,N_25724);
and U27062 (N_27062,N_26029,N_25636);
nand U27063 (N_27063,N_25688,N_26048);
and U27064 (N_27064,N_26889,N_25546);
and U27065 (N_27065,N_26470,N_25959);
nor U27066 (N_27066,N_25771,N_26548);
nor U27067 (N_27067,N_25865,N_25717);
and U27068 (N_27068,N_26677,N_26143);
and U27069 (N_27069,N_25618,N_25752);
nor U27070 (N_27070,N_25617,N_25622);
nand U27071 (N_27071,N_26617,N_25855);
nand U27072 (N_27072,N_26879,N_26999);
nor U27073 (N_27073,N_26145,N_25862);
or U27074 (N_27074,N_26228,N_26857);
nor U27075 (N_27075,N_25503,N_25810);
or U27076 (N_27076,N_26393,N_25530);
nand U27077 (N_27077,N_26521,N_25534);
nand U27078 (N_27078,N_25536,N_25633);
and U27079 (N_27079,N_26319,N_26207);
or U27080 (N_27080,N_25612,N_26655);
or U27081 (N_27081,N_26982,N_26128);
or U27082 (N_27082,N_26696,N_26164);
nor U27083 (N_27083,N_25507,N_26199);
nand U27084 (N_27084,N_26756,N_26116);
or U27085 (N_27085,N_26439,N_25755);
and U27086 (N_27086,N_25516,N_26204);
nand U27087 (N_27087,N_26598,N_25861);
and U27088 (N_27088,N_26332,N_26298);
nor U27089 (N_27089,N_25852,N_25760);
nand U27090 (N_27090,N_26777,N_26514);
nand U27091 (N_27091,N_25860,N_26813);
nand U27092 (N_27092,N_25750,N_25713);
and U27093 (N_27093,N_26606,N_26736);
or U27094 (N_27094,N_26078,N_25910);
and U27095 (N_27095,N_26612,N_26702);
xor U27096 (N_27096,N_26661,N_26988);
and U27097 (N_27097,N_26342,N_25596);
or U27098 (N_27098,N_26651,N_26600);
nor U27099 (N_27099,N_25814,N_26270);
and U27100 (N_27100,N_26454,N_26014);
or U27101 (N_27101,N_26295,N_26355);
xnor U27102 (N_27102,N_26361,N_26482);
or U27103 (N_27103,N_26318,N_25651);
and U27104 (N_27104,N_26433,N_26132);
or U27105 (N_27105,N_25671,N_26042);
or U27106 (N_27106,N_26877,N_26658);
and U27107 (N_27107,N_26678,N_26668);
and U27108 (N_27108,N_26186,N_26530);
xnor U27109 (N_27109,N_26955,N_26665);
or U27110 (N_27110,N_25877,N_26149);
nor U27111 (N_27111,N_26290,N_26113);
and U27112 (N_27112,N_26631,N_26261);
xnor U27113 (N_27113,N_26384,N_26383);
nor U27114 (N_27114,N_26837,N_25787);
and U27115 (N_27115,N_25912,N_25812);
and U27116 (N_27116,N_26939,N_25822);
and U27117 (N_27117,N_26314,N_26560);
nor U27118 (N_27118,N_25914,N_26452);
or U27119 (N_27119,N_26604,N_25984);
or U27120 (N_27120,N_26300,N_26185);
nand U27121 (N_27121,N_26110,N_25510);
nand U27122 (N_27122,N_25624,N_25916);
or U27123 (N_27123,N_26353,N_26583);
xnor U27124 (N_27124,N_26931,N_25842);
nand U27125 (N_27125,N_26974,N_26305);
nand U27126 (N_27126,N_25584,N_26418);
or U27127 (N_27127,N_25757,N_26925);
or U27128 (N_27128,N_25819,N_26120);
xnor U27129 (N_27129,N_25872,N_25758);
and U27130 (N_27130,N_25532,N_26840);
nor U27131 (N_27131,N_25663,N_26966);
xnor U27132 (N_27132,N_26947,N_26209);
xnor U27133 (N_27133,N_25785,N_26748);
or U27134 (N_27134,N_26061,N_25885);
xnor U27135 (N_27135,N_26189,N_26755);
nand U27136 (N_27136,N_26474,N_26758);
xor U27137 (N_27137,N_26354,N_26591);
or U27138 (N_27138,N_25791,N_26805);
nor U27139 (N_27139,N_26559,N_25563);
nor U27140 (N_27140,N_25832,N_26394);
or U27141 (N_27141,N_25638,N_25513);
nor U27142 (N_27142,N_26247,N_26089);
and U27143 (N_27143,N_26401,N_26056);
and U27144 (N_27144,N_26734,N_25517);
and U27145 (N_27145,N_25733,N_25774);
xor U27146 (N_27146,N_26607,N_26739);
nand U27147 (N_27147,N_26366,N_26676);
or U27148 (N_27148,N_26028,N_26843);
and U27149 (N_27149,N_25608,N_26964);
nor U27150 (N_27150,N_25548,N_25705);
xor U27151 (N_27151,N_25601,N_26798);
nor U27152 (N_27152,N_26887,N_25944);
nor U27153 (N_27153,N_26674,N_26069);
and U27154 (N_27154,N_26706,N_26810);
nor U27155 (N_27155,N_26271,N_26007);
nor U27156 (N_27156,N_26451,N_26460);
xnor U27157 (N_27157,N_26333,N_26420);
xnor U27158 (N_27158,N_26808,N_26860);
and U27159 (N_27159,N_25888,N_26223);
and U27160 (N_27160,N_25880,N_26595);
nand U27161 (N_27161,N_25841,N_26416);
xnor U27162 (N_27162,N_26147,N_26422);
xnor U27163 (N_27163,N_26171,N_25715);
or U27164 (N_27164,N_26304,N_25696);
or U27165 (N_27165,N_26005,N_26831);
nand U27166 (N_27166,N_25985,N_26832);
xor U27167 (N_27167,N_26259,N_25784);
xor U27168 (N_27168,N_25859,N_26090);
and U27169 (N_27169,N_25905,N_26198);
or U27170 (N_27170,N_26442,N_25960);
and U27171 (N_27171,N_26096,N_26691);
nand U27172 (N_27172,N_26667,N_26475);
or U27173 (N_27173,N_26368,N_26727);
or U27174 (N_27174,N_26277,N_26724);
nor U27175 (N_27175,N_26571,N_25829);
or U27176 (N_27176,N_25918,N_25967);
nand U27177 (N_27177,N_26313,N_25751);
and U27178 (N_27178,N_26461,N_26448);
xor U27179 (N_27179,N_26910,N_26820);
or U27180 (N_27180,N_25500,N_25703);
or U27181 (N_27181,N_26455,N_25900);
and U27182 (N_27182,N_25552,N_26034);
and U27183 (N_27183,N_26001,N_25736);
or U27184 (N_27184,N_25709,N_25502);
nand U27185 (N_27185,N_26757,N_26515);
or U27186 (N_27186,N_26205,N_26823);
or U27187 (N_27187,N_25556,N_26875);
xor U27188 (N_27188,N_26990,N_25658);
or U27189 (N_27189,N_26387,N_25538);
xnor U27190 (N_27190,N_26103,N_25613);
or U27191 (N_27191,N_26664,N_25664);
xnor U27192 (N_27192,N_25924,N_26834);
or U27193 (N_27193,N_25948,N_25678);
and U27194 (N_27194,N_25920,N_26338);
and U27195 (N_27195,N_26493,N_26502);
nor U27196 (N_27196,N_26322,N_26650);
and U27197 (N_27197,N_25565,N_26913);
and U27198 (N_27198,N_25780,N_26490);
xor U27199 (N_27199,N_26647,N_26158);
xor U27200 (N_27200,N_26170,N_25588);
xor U27201 (N_27201,N_25630,N_26278);
and U27202 (N_27202,N_26723,N_26792);
nand U27203 (N_27203,N_26582,N_26895);
nor U27204 (N_27204,N_25772,N_25953);
xor U27205 (N_27205,N_26711,N_26473);
or U27206 (N_27206,N_26071,N_26534);
nand U27207 (N_27207,N_26180,N_26826);
nand U27208 (N_27208,N_26732,N_26836);
nand U27209 (N_27209,N_25520,N_26081);
or U27210 (N_27210,N_25566,N_26326);
nand U27211 (N_27211,N_26662,N_26297);
nand U27212 (N_27212,N_26025,N_26276);
nand U27213 (N_27213,N_26566,N_26489);
and U27214 (N_27214,N_25779,N_26496);
nand U27215 (N_27215,N_26218,N_26426);
or U27216 (N_27216,N_25615,N_25782);
nor U27217 (N_27217,N_26262,N_25952);
nand U27218 (N_27218,N_26082,N_25629);
nand U27219 (N_27219,N_26003,N_26424);
and U27220 (N_27220,N_26264,N_26842);
nand U27221 (N_27221,N_26994,N_25699);
nor U27222 (N_27222,N_25831,N_25700);
xnor U27223 (N_27223,N_26928,N_25881);
or U27224 (N_27224,N_26299,N_25839);
and U27225 (N_27225,N_26803,N_25587);
or U27226 (N_27226,N_25874,N_25845);
and U27227 (N_27227,N_25828,N_26553);
and U27228 (N_27228,N_25564,N_25786);
xnor U27229 (N_27229,N_26152,N_25943);
nor U27230 (N_27230,N_26233,N_26317);
nor U27231 (N_27231,N_26425,N_26478);
xor U27232 (N_27232,N_25825,N_26640);
xor U27233 (N_27233,N_26714,N_26301);
and U27234 (N_27234,N_25727,N_26550);
nand U27235 (N_27235,N_26980,N_25580);
or U27236 (N_27236,N_26572,N_26688);
nor U27237 (N_27237,N_26142,N_26848);
or U27238 (N_27238,N_26337,N_25763);
xnor U27239 (N_27239,N_26196,N_26894);
xnor U27240 (N_27240,N_25793,N_26869);
or U27241 (N_27241,N_26224,N_26221);
and U27242 (N_27242,N_26588,N_26184);
xnor U27243 (N_27243,N_25795,N_26457);
nor U27244 (N_27244,N_26844,N_26445);
and U27245 (N_27245,N_26526,N_26616);
and U27246 (N_27246,N_26471,N_26408);
xnor U27247 (N_27247,N_26830,N_25853);
or U27248 (N_27248,N_26914,N_26621);
nand U27249 (N_27249,N_25537,N_26498);
nand U27250 (N_27250,N_26829,N_26684);
nor U27251 (N_27251,N_26957,N_26699);
or U27252 (N_27252,N_26510,N_26362);
or U27253 (N_27253,N_26243,N_26043);
nand U27254 (N_27254,N_26970,N_26363);
and U27255 (N_27255,N_26374,N_26121);
and U27256 (N_27256,N_26086,N_26632);
and U27257 (N_27257,N_26372,N_26329);
and U27258 (N_27258,N_25672,N_25933);
and U27259 (N_27259,N_26033,N_25955);
nand U27260 (N_27260,N_25954,N_26791);
or U27261 (N_27261,N_26663,N_26462);
nand U27262 (N_27262,N_25968,N_25682);
xor U27263 (N_27263,N_25525,N_26943);
nand U27264 (N_27264,N_26975,N_25575);
and U27265 (N_27265,N_25505,N_25640);
nor U27266 (N_27266,N_26407,N_26799);
nor U27267 (N_27267,N_25514,N_26108);
nor U27268 (N_27268,N_25906,N_25708);
nand U27269 (N_27269,N_25858,N_26924);
or U27270 (N_27270,N_25983,N_26019);
nand U27271 (N_27271,N_26853,N_26117);
xor U27272 (N_27272,N_25634,N_26468);
or U27273 (N_27273,N_26992,N_26215);
nor U27274 (N_27274,N_26404,N_25710);
xor U27275 (N_27275,N_26718,N_25898);
nand U27276 (N_27276,N_26740,N_26923);
nor U27277 (N_27277,N_25972,N_25643);
or U27278 (N_27278,N_26870,N_26279);
and U27279 (N_27279,N_25610,N_26963);
or U27280 (N_27280,N_26517,N_26623);
xnor U27281 (N_27281,N_25674,N_26513);
xnor U27282 (N_27282,N_26596,N_26016);
or U27283 (N_27283,N_25691,N_26356);
nor U27284 (N_27284,N_26181,N_25676);
nand U27285 (N_27285,N_26785,N_26341);
xor U27286 (N_27286,N_26027,N_26359);
and U27287 (N_27287,N_26491,N_26746);
or U27288 (N_27288,N_26111,N_26340);
xnor U27289 (N_27289,N_25649,N_26563);
or U27290 (N_27290,N_25947,N_25623);
nand U27291 (N_27291,N_25753,N_25759);
and U27292 (N_27292,N_25581,N_26694);
or U27293 (N_27293,N_26272,N_25962);
nand U27294 (N_27294,N_26953,N_26783);
or U27295 (N_27295,N_25927,N_25789);
nor U27296 (N_27296,N_26993,N_25975);
or U27297 (N_27297,N_25645,N_26365);
and U27298 (N_27298,N_26965,N_26680);
nand U27299 (N_27299,N_26692,N_26213);
or U27300 (N_27300,N_26610,N_26432);
or U27301 (N_27301,N_25873,N_26084);
and U27302 (N_27302,N_26554,N_26715);
xor U27303 (N_27303,N_25808,N_26722);
or U27304 (N_27304,N_25802,N_26916);
nand U27305 (N_27305,N_26465,N_26527);
nor U27306 (N_27306,N_26088,N_26073);
nand U27307 (N_27307,N_25641,N_26760);
or U27308 (N_27308,N_25578,N_26753);
and U27309 (N_27309,N_25847,N_26789);
or U27310 (N_27310,N_25569,N_26580);
and U27311 (N_27311,N_25868,N_25796);
and U27312 (N_27312,N_25616,N_25598);
and U27313 (N_27313,N_26771,N_25550);
or U27314 (N_27314,N_26961,N_26360);
nor U27315 (N_27315,N_25942,N_25941);
nor U27316 (N_27316,N_25642,N_26179);
xor U27317 (N_27317,N_26744,N_26921);
nand U27318 (N_27318,N_25685,N_26060);
and U27319 (N_27319,N_26006,N_25965);
xnor U27320 (N_27320,N_26689,N_25949);
and U27321 (N_27321,N_26900,N_26519);
or U27322 (N_27322,N_25897,N_25895);
xnor U27323 (N_27323,N_26818,N_25887);
or U27324 (N_27324,N_25989,N_26584);
or U27325 (N_27325,N_25800,N_25693);
nand U27326 (N_27326,N_26841,N_25982);
xor U27327 (N_27327,N_25837,N_25997);
or U27328 (N_27328,N_26940,N_26021);
nand U27329 (N_27329,N_26687,N_26653);
nor U27330 (N_27330,N_26055,N_26488);
and U27331 (N_27331,N_25501,N_25716);
or U27332 (N_27332,N_26188,N_26484);
or U27333 (N_27333,N_26373,N_26944);
xor U27334 (N_27334,N_26700,N_26804);
xor U27335 (N_27335,N_25922,N_26666);
nand U27336 (N_27336,N_25720,N_26010);
nor U27337 (N_27337,N_26811,N_26011);
or U27338 (N_27338,N_26893,N_26670);
nand U27339 (N_27339,N_25687,N_25977);
nand U27340 (N_27340,N_26172,N_26720);
or U27341 (N_27341,N_26735,N_26315);
xor U27342 (N_27342,N_25749,N_25813);
nor U27343 (N_27343,N_25519,N_26637);
nand U27344 (N_27344,N_26660,N_26112);
nor U27345 (N_27345,N_25614,N_25970);
and U27346 (N_27346,N_26948,N_26035);
xnor U27347 (N_27347,N_26477,N_25635);
nand U27348 (N_27348,N_26729,N_26101);
and U27349 (N_27349,N_26569,N_26242);
nor U27350 (N_27350,N_25934,N_26072);
xnor U27351 (N_27351,N_25665,N_26386);
xnor U27352 (N_27352,N_25653,N_26447);
nand U27353 (N_27353,N_26124,N_26392);
nand U27354 (N_27354,N_26436,N_26570);
nor U27355 (N_27355,N_26952,N_26533);
and U27356 (N_27356,N_26801,N_26251);
xor U27357 (N_27357,N_26645,N_25930);
nand U27358 (N_27358,N_26772,N_26358);
or U27359 (N_27359,N_26802,N_25527);
xor U27360 (N_27360,N_26926,N_25597);
and U27361 (N_27361,N_26138,N_26765);
xor U27362 (N_27362,N_25824,N_26155);
nor U27363 (N_27363,N_25999,N_26009);
and U27364 (N_27364,N_26347,N_26969);
nand U27365 (N_27365,N_26268,N_26012);
xnor U27366 (N_27366,N_26817,N_26068);
nand U27367 (N_27367,N_26463,N_26370);
or U27368 (N_27368,N_26265,N_26639);
nor U27369 (N_27369,N_26396,N_26872);
xnor U27370 (N_27370,N_25823,N_26741);
xor U27371 (N_27371,N_25695,N_26414);
or U27372 (N_27372,N_26859,N_26291);
nor U27373 (N_27373,N_25611,N_26897);
or U27374 (N_27374,N_26750,N_25939);
or U27375 (N_27375,N_26985,N_26160);
and U27376 (N_27376,N_26194,N_26695);
nor U27377 (N_27377,N_25506,N_25871);
and U27378 (N_27378,N_25988,N_26503);
or U27379 (N_27379,N_26881,N_25804);
or U27380 (N_27380,N_25744,N_25756);
or U27381 (N_27381,N_26367,N_26814);
or U27382 (N_27382,N_25973,N_26310);
nor U27383 (N_27383,N_26991,N_26178);
nand U27384 (N_27384,N_26945,N_25951);
nor U27385 (N_27385,N_25652,N_26917);
and U27386 (N_27386,N_26769,N_25738);
or U27387 (N_27387,N_26922,N_26031);
nand U27388 (N_27388,N_25821,N_26087);
xor U27389 (N_27389,N_26850,N_26284);
nand U27390 (N_27390,N_26638,N_26747);
nor U27391 (N_27391,N_26100,N_26467);
and U27392 (N_27392,N_25915,N_25748);
nand U27393 (N_27393,N_26316,N_26539);
nor U27394 (N_27394,N_26908,N_25883);
xor U27395 (N_27395,N_26997,N_25761);
and U27396 (N_27396,N_25541,N_26976);
and U27397 (N_27397,N_25929,N_26642);
nand U27398 (N_27398,N_26444,N_25840);
and U27399 (N_27399,N_25686,N_25628);
nor U27400 (N_27400,N_25864,N_26371);
or U27401 (N_27401,N_25667,N_25806);
and U27402 (N_27402,N_25559,N_26998);
or U27403 (N_27403,N_25950,N_25741);
or U27404 (N_27404,N_25743,N_26529);
nor U27405 (N_27405,N_26611,N_26476);
nor U27406 (N_27406,N_26793,N_26568);
and U27407 (N_27407,N_25798,N_25567);
nor U27408 (N_27408,N_25990,N_25963);
xnor U27409 (N_27409,N_26544,N_25544);
and U27410 (N_27410,N_26778,N_25899);
or U27411 (N_27411,N_25586,N_25627);
xnor U27412 (N_27412,N_25702,N_25560);
xor U27413 (N_27413,N_25603,N_26459);
nor U27414 (N_27414,N_26531,N_26522);
nand U27415 (N_27415,N_26144,N_25856);
or U27416 (N_27416,N_25935,N_26505);
and U27417 (N_27417,N_26325,N_25894);
xor U27418 (N_27418,N_25995,N_26201);
xnor U27419 (N_27419,N_26252,N_26780);
and U27420 (N_27420,N_25683,N_25599);
xor U27421 (N_27421,N_25783,N_25827);
and U27422 (N_27422,N_26738,N_26594);
xnor U27423 (N_27423,N_26862,N_25620);
xor U27424 (N_27424,N_26429,N_25669);
and U27425 (N_27425,N_26311,N_25773);
nor U27426 (N_27426,N_25731,N_26709);
or U27427 (N_27427,N_25659,N_26232);
xor U27428 (N_27428,N_26770,N_26919);
xnor U27429 (N_27429,N_26936,N_26984);
nor U27430 (N_27430,N_26937,N_25706);
or U27431 (N_27431,N_26697,N_25980);
xnor U27432 (N_27432,N_26652,N_26308);
xnor U27433 (N_27433,N_26066,N_25666);
nor U27434 (N_27434,N_25673,N_26573);
nor U27435 (N_27435,N_25797,N_25911);
xor U27436 (N_27436,N_26828,N_26849);
and U27437 (N_27437,N_25826,N_25843);
or U27438 (N_27438,N_26419,N_26409);
nand U27439 (N_27439,N_25572,N_26125);
xnor U27440 (N_27440,N_26960,N_25735);
nor U27441 (N_27441,N_25834,N_25680);
xor U27442 (N_27442,N_26752,N_26044);
nand U27443 (N_27443,N_26469,N_26107);
and U27444 (N_27444,N_26492,N_25625);
or U27445 (N_27445,N_25992,N_25732);
xnor U27446 (N_27446,N_26399,N_26274);
or U27447 (N_27447,N_25681,N_26884);
nand U27448 (N_27448,N_26549,N_26962);
nor U27449 (N_27449,N_26114,N_26256);
xor U27450 (N_27450,N_26208,N_26950);
nand U27451 (N_27451,N_26620,N_25936);
xnor U27452 (N_27452,N_26888,N_25794);
nor U27453 (N_27453,N_26255,N_26507);
and U27454 (N_27454,N_26400,N_25555);
nor U27455 (N_27455,N_26846,N_25820);
xor U27456 (N_27456,N_26156,N_25582);
xor U27457 (N_27457,N_26518,N_26495);
or U27458 (N_27458,N_25974,N_26593);
or U27459 (N_27459,N_26219,N_26046);
or U27460 (N_27460,N_26708,N_26239);
nor U27461 (N_27461,N_26200,N_25590);
nor U27462 (N_27462,N_26391,N_25504);
and U27463 (N_27463,N_26402,N_26312);
xor U27464 (N_27464,N_26892,N_26812);
and U27465 (N_27465,N_26682,N_26324);
xor U27466 (N_27466,N_26520,N_25661);
and U27467 (N_27467,N_25721,N_26733);
xnor U27468 (N_27468,N_25609,N_25937);
or U27469 (N_27469,N_25531,N_26349);
xnor U27470 (N_27470,N_26092,N_26464);
and U27471 (N_27471,N_26958,N_25714);
xnor U27472 (N_27472,N_26501,N_26435);
xor U27473 (N_27473,N_26567,N_26899);
nand U27474 (N_27474,N_26104,N_26774);
xnor U27475 (N_27475,N_25901,N_26624);
or U27476 (N_27476,N_25846,N_25737);
xor U27477 (N_27477,N_26438,N_26146);
nor U27478 (N_27478,N_26118,N_26041);
nor U27479 (N_27479,N_26093,N_26634);
xnor U27480 (N_27480,N_26450,N_26094);
or U27481 (N_27481,N_26885,N_25592);
xor U27482 (N_27482,N_26807,N_26855);
or U27483 (N_27483,N_26726,N_26364);
or U27484 (N_27484,N_25769,N_26795);
nor U27485 (N_27485,N_26809,N_25913);
nand U27486 (N_27486,N_26260,N_26499);
nor U27487 (N_27487,N_26134,N_26911);
nand U27488 (N_27488,N_25790,N_26428);
nor U27489 (N_27489,N_26972,N_26956);
or U27490 (N_27490,N_26024,N_25844);
nand U27491 (N_27491,N_26690,N_25931);
xor U27492 (N_27492,N_26267,N_26390);
or U27493 (N_27493,N_25711,N_26321);
and U27494 (N_27494,N_26320,N_25745);
nand U27495 (N_27495,N_25904,N_26263);
xor U27496 (N_27496,N_25996,N_25889);
nor U27497 (N_27497,N_26685,N_26825);
or U27498 (N_27498,N_26764,N_26346);
and U27499 (N_27499,N_26742,N_25542);
and U27500 (N_27500,N_26861,N_25632);
or U27501 (N_27501,N_26415,N_25554);
or U27502 (N_27502,N_25928,N_25747);
nand U27503 (N_27503,N_25619,N_26656);
xor U27504 (N_27504,N_26905,N_26851);
nand U27505 (N_27505,N_25734,N_25762);
nor U27506 (N_27506,N_26989,N_25770);
and U27507 (N_27507,N_25518,N_26456);
or U27508 (N_27508,N_26904,N_25522);
xor U27509 (N_27509,N_25766,N_26730);
nand U27510 (N_27510,N_25606,N_26901);
nor U27511 (N_27511,N_25723,N_26717);
and U27512 (N_27512,N_25677,N_25768);
xnor U27513 (N_27513,N_26136,N_25857);
or U27514 (N_27514,N_26906,N_25867);
nor U27515 (N_27515,N_26648,N_26336);
xnor U27516 (N_27516,N_26628,N_25807);
nor U27517 (N_27517,N_26106,N_25879);
or U27518 (N_27518,N_26725,N_25903);
or U27519 (N_27519,N_26890,N_26763);
or U27520 (N_27520,N_26497,N_26977);
xor U27521 (N_27521,N_26597,N_26657);
xnor U27522 (N_27522,N_25932,N_26821);
or U27523 (N_27523,N_26197,N_26229);
xor U27524 (N_27524,N_26775,N_26886);
nor U27525 (N_27525,N_25792,N_26091);
or U27526 (N_27526,N_26679,N_26816);
xnor U27527 (N_27527,N_26040,N_26225);
nor U27528 (N_27528,N_26175,N_26779);
xor U27529 (N_27529,N_25579,N_25662);
xor U27530 (N_27530,N_25781,N_26037);
or U27531 (N_27531,N_25589,N_25869);
nor U27532 (N_27532,N_26506,N_26095);
nand U27533 (N_27533,N_26800,N_25994);
xor U27534 (N_27534,N_25971,N_26659);
or U27535 (N_27535,N_26097,N_26500);
or U27536 (N_27536,N_26017,N_26576);
xnor U27537 (N_27537,N_26099,N_26938);
nand U27538 (N_27538,N_26369,N_26411);
or U27539 (N_27539,N_26797,N_26202);
nor U27540 (N_27540,N_26405,N_25712);
nor U27541 (N_27541,N_26441,N_26703);
nand U27542 (N_27542,N_25775,N_25896);
nand U27543 (N_27543,N_26686,N_26074);
and U27544 (N_27544,N_25650,N_25866);
and U27545 (N_27545,N_26512,N_26289);
and U27546 (N_27546,N_26983,N_26586);
or U27547 (N_27547,N_26288,N_25809);
nor U27548 (N_27548,N_26226,N_26671);
xnor U27549 (N_27549,N_26480,N_26508);
or U27550 (N_27550,N_26935,N_25870);
nand U27551 (N_27551,N_25698,N_25707);
nor U27552 (N_27552,N_26934,N_26151);
and U27553 (N_27553,N_26238,N_26978);
nor U27554 (N_27554,N_26077,N_26054);
and U27555 (N_27555,N_26176,N_26669);
nand U27556 (N_27556,N_26382,N_25799);
or U27557 (N_27557,N_26214,N_26453);
and U27558 (N_27558,N_26351,N_26891);
nor U27559 (N_27559,N_26334,N_26835);
or U27560 (N_27560,N_26323,N_25657);
and U27561 (N_27561,N_26443,N_26587);
or U27562 (N_27562,N_26406,N_26562);
nor U27563 (N_27563,N_25815,N_26173);
nor U27564 (N_27564,N_26302,N_26004);
xor U27565 (N_27565,N_26206,N_26472);
nor U27566 (N_27566,N_26352,N_26240);
or U27567 (N_27567,N_25605,N_26427);
and U27568 (N_27568,N_26784,N_26681);
nand U27569 (N_27569,N_26845,N_26137);
nand U27570 (N_27570,N_26592,N_26629);
xor U27571 (N_27571,N_26182,N_26838);
or U27572 (N_27572,N_25803,N_26235);
xnor U27573 (N_27573,N_25689,N_25969);
and U27574 (N_27574,N_26287,N_26918);
nand U27575 (N_27575,N_26293,N_26280);
nor U27576 (N_27576,N_25547,N_26487);
nor U27577 (N_27577,N_25978,N_26051);
and U27578 (N_27578,N_25838,N_26412);
and U27579 (N_27579,N_25851,N_25595);
nor U27580 (N_27580,N_26130,N_26047);
and U27581 (N_27581,N_26015,N_26602);
and U27582 (N_27582,N_26285,N_25593);
and U27583 (N_27583,N_26675,N_26273);
nand U27584 (N_27584,N_26858,N_26139);
and U27585 (N_27585,N_26766,N_26920);
and U27586 (N_27586,N_26941,N_26348);
or U27587 (N_27587,N_26552,N_25508);
nand U27588 (N_27588,N_26909,N_26528);
or U27589 (N_27589,N_26794,N_26827);
nand U27590 (N_27590,N_25535,N_26880);
nor U27591 (N_27591,N_25979,N_25692);
nor U27592 (N_27592,N_25528,N_26731);
xnor U27593 (N_27593,N_26523,N_26195);
or U27594 (N_27594,N_26951,N_26398);
nand U27595 (N_27595,N_26413,N_25602);
xor U27596 (N_27596,N_26545,N_26008);
xnor U27597 (N_27597,N_26292,N_26234);
or U27598 (N_27598,N_26098,N_26968);
nor U27599 (N_27599,N_25854,N_26357);
and U27600 (N_27600,N_26032,N_26762);
nor U27601 (N_27601,N_26257,N_26555);
nand U27602 (N_27602,N_25585,N_26135);
or U27603 (N_27603,N_26896,N_25573);
and U27604 (N_27604,N_26064,N_26822);
and U27605 (N_27605,N_26129,N_26395);
or U27606 (N_27606,N_26898,N_26754);
nor U27607 (N_27607,N_26787,N_26839);
xnor U27608 (N_27608,N_26626,N_26166);
and U27609 (N_27609,N_25964,N_26786);
nand U27610 (N_27610,N_26458,N_25833);
or U27611 (N_27611,N_26083,N_26057);
or U27612 (N_27612,N_26546,N_26350);
xor U27613 (N_27613,N_26759,N_26782);
xor U27614 (N_27614,N_26930,N_26721);
and U27615 (N_27615,N_26633,N_25594);
or U27616 (N_27616,N_26745,N_26296);
or U27617 (N_27617,N_26551,N_26430);
nor U27618 (N_27618,N_26967,N_25684);
or U27619 (N_27619,N_26622,N_25945);
nor U27620 (N_27620,N_26065,N_26115);
nand U27621 (N_27621,N_26707,N_26981);
nand U27622 (N_27622,N_25966,N_26080);
xor U27623 (N_27623,N_26524,N_25890);
nand U27624 (N_27624,N_26693,N_25694);
nand U27625 (N_27625,N_26062,N_26449);
nand U27626 (N_27626,N_26389,N_25981);
or U27627 (N_27627,N_26574,N_25801);
xor U27628 (N_27628,N_25991,N_26380);
nor U27629 (N_27629,N_25526,N_26403);
nand U27630 (N_27630,N_25778,N_26713);
nand U27631 (N_27631,N_25509,N_26241);
or U27632 (N_27632,N_25848,N_26927);
or U27633 (N_27633,N_25718,N_26646);
nor U27634 (N_27634,N_26876,N_25923);
nor U27635 (N_27635,N_26327,N_26067);
nor U27636 (N_27636,N_26038,N_25675);
or U27637 (N_27637,N_26704,N_26258);
xor U27638 (N_27638,N_25882,N_26131);
xnor U27639 (N_27639,N_26345,N_26210);
or U27640 (N_27640,N_26749,N_26986);
xnor U27641 (N_27641,N_26417,N_26344);
nand U27642 (N_27642,N_26230,N_25725);
xnor U27643 (N_27643,N_26169,N_26246);
xor U27644 (N_27644,N_26039,N_25976);
nand U27645 (N_27645,N_25697,N_25739);
or U27646 (N_27646,N_26023,N_26705);
or U27647 (N_27647,N_26018,N_26540);
xor U27648 (N_27648,N_25754,N_26381);
nor U27649 (N_27649,N_26535,N_26806);
xnor U27650 (N_27650,N_26109,N_26971);
nand U27651 (N_27651,N_26824,N_26153);
and U27652 (N_27652,N_25987,N_25644);
and U27653 (N_27653,N_26388,N_26737);
or U27654 (N_27654,N_26140,N_26466);
nor U27655 (N_27655,N_26556,N_25835);
or U27656 (N_27656,N_26543,N_26227);
xor U27657 (N_27657,N_26781,N_26376);
and U27658 (N_27658,N_25690,N_26761);
xnor U27659 (N_27659,N_26932,N_26049);
xnor U27660 (N_27660,N_26434,N_25722);
and U27661 (N_27661,N_25919,N_26959);
nor U27662 (N_27662,N_25607,N_25728);
and U27663 (N_27663,N_25577,N_26878);
nor U27664 (N_27664,N_26796,N_25818);
nor U27665 (N_27665,N_25740,N_25907);
xor U27666 (N_27666,N_26123,N_26867);
nor U27667 (N_27667,N_26168,N_26294);
nor U27668 (N_27668,N_26058,N_26286);
nor U27669 (N_27669,N_26987,N_26494);
xor U27670 (N_27670,N_26912,N_26127);
or U27671 (N_27671,N_25553,N_26187);
xor U27672 (N_27672,N_26050,N_26728);
xor U27673 (N_27673,N_25908,N_25830);
or U27674 (N_27674,N_26177,N_26133);
or U27675 (N_27675,N_26915,N_26331);
or U27676 (N_27676,N_26174,N_26378);
and U27677 (N_27677,N_26618,N_25998);
nor U27678 (N_27678,N_26119,N_26000);
or U27679 (N_27679,N_26683,N_26613);
and U27680 (N_27680,N_25986,N_26159);
xnor U27681 (N_27681,N_26942,N_26874);
nor U27682 (N_27682,N_25742,N_26565);
and U27683 (N_27683,N_25764,N_25545);
nand U27684 (N_27684,N_26193,N_26244);
or U27685 (N_27685,N_26716,N_26485);
nor U27686 (N_27686,N_25891,N_25892);
xnor U27687 (N_27687,N_25878,N_26712);
nor U27688 (N_27688,N_26547,N_26973);
nand U27689 (N_27689,N_25902,N_26536);
or U27690 (N_27690,N_25719,N_25849);
nand U27691 (N_27691,N_26847,N_26643);
nor U27692 (N_27692,N_26162,N_25637);
and U27693 (N_27693,N_26085,N_26511);
and U27694 (N_27694,N_26437,N_25512);
and U27695 (N_27695,N_26281,N_26212);
nor U27696 (N_27696,N_26479,N_25917);
and U27697 (N_27697,N_26063,N_26865);
xnor U27698 (N_27698,N_26933,N_25540);
and U27699 (N_27699,N_25660,N_26190);
xnor U27700 (N_27700,N_26148,N_26282);
and U27701 (N_27701,N_26220,N_25571);
and U27702 (N_27702,N_26542,N_26579);
xor U27703 (N_27703,N_25523,N_26053);
nor U27704 (N_27704,N_26303,N_26698);
and U27705 (N_27705,N_26250,N_26481);
nor U27706 (N_27706,N_26864,N_25746);
nand U27707 (N_27707,N_26335,N_26105);
or U27708 (N_27708,N_26605,N_25679);
or U27709 (N_27709,N_25726,N_26627);
xnor U27710 (N_27710,N_25576,N_25626);
nor U27711 (N_27711,N_25940,N_26635);
nor U27712 (N_27712,N_25561,N_26157);
nand U27713 (N_27713,N_26578,N_25648);
or U27714 (N_27714,N_26231,N_26751);
xor U27715 (N_27715,N_26236,N_26619);
xor U27716 (N_27716,N_26871,N_26776);
xor U27717 (N_27717,N_25811,N_26440);
or U27718 (N_27718,N_26122,N_26283);
or U27719 (N_27719,N_25850,N_25993);
xor U27720 (N_27720,N_26266,N_26431);
xor U27721 (N_27721,N_25551,N_25701);
or U27722 (N_27722,N_26020,N_25767);
xnor U27723 (N_27723,N_26767,N_25524);
nand U27724 (N_27724,N_26907,N_26768);
nor U27725 (N_27725,N_26883,N_26013);
xor U27726 (N_27726,N_25788,N_25926);
nand U27727 (N_27727,N_26672,N_26026);
nand U27728 (N_27728,N_25668,N_26022);
or U27729 (N_27729,N_26601,N_26307);
or U27730 (N_27730,N_26192,N_26509);
and U27731 (N_27731,N_26165,N_25543);
nand U27732 (N_27732,N_25511,N_26868);
nand U27733 (N_27733,N_25816,N_26141);
nand U27734 (N_27734,N_26275,N_25886);
and U27735 (N_27735,N_25938,N_25655);
nand U27736 (N_27736,N_25817,N_26328);
and U27737 (N_27737,N_26995,N_26854);
nand U27738 (N_27738,N_26076,N_25604);
xor U27739 (N_27739,N_26217,N_26558);
xnor U27740 (N_27740,N_26532,N_25591);
xnor U27741 (N_27741,N_25562,N_26790);
nand U27742 (N_27742,N_25621,N_25539);
and U27743 (N_27743,N_26504,N_26815);
nor U27744 (N_27744,N_26949,N_26377);
nand U27745 (N_27745,N_25875,N_25647);
or U27746 (N_27746,N_26882,N_26339);
nand U27747 (N_27747,N_26585,N_26609);
and U27748 (N_27748,N_25776,N_25729);
nor U27749 (N_27749,N_26625,N_26216);
and U27750 (N_27750,N_26829,N_26118);
nand U27751 (N_27751,N_26338,N_25680);
and U27752 (N_27752,N_26416,N_25565);
xnor U27753 (N_27753,N_25879,N_25866);
nor U27754 (N_27754,N_25932,N_26114);
or U27755 (N_27755,N_25778,N_26737);
xor U27756 (N_27756,N_26439,N_26092);
nand U27757 (N_27757,N_26496,N_26856);
or U27758 (N_27758,N_26198,N_26276);
xnor U27759 (N_27759,N_25610,N_26007);
nor U27760 (N_27760,N_26030,N_26894);
or U27761 (N_27761,N_25610,N_26650);
and U27762 (N_27762,N_25757,N_26287);
and U27763 (N_27763,N_25877,N_25975);
or U27764 (N_27764,N_26237,N_25997);
nor U27765 (N_27765,N_25868,N_25658);
nand U27766 (N_27766,N_26024,N_26460);
and U27767 (N_27767,N_25838,N_25572);
or U27768 (N_27768,N_26992,N_26476);
and U27769 (N_27769,N_26077,N_26148);
nand U27770 (N_27770,N_25705,N_26469);
or U27771 (N_27771,N_25869,N_25777);
nor U27772 (N_27772,N_26748,N_26023);
nand U27773 (N_27773,N_26165,N_26568);
nor U27774 (N_27774,N_25568,N_25774);
xor U27775 (N_27775,N_26927,N_25839);
or U27776 (N_27776,N_26588,N_25719);
and U27777 (N_27777,N_25625,N_25831);
or U27778 (N_27778,N_26765,N_25962);
xnor U27779 (N_27779,N_26121,N_26023);
xor U27780 (N_27780,N_26225,N_26529);
nand U27781 (N_27781,N_26798,N_25940);
or U27782 (N_27782,N_26400,N_26711);
and U27783 (N_27783,N_26115,N_25986);
xnor U27784 (N_27784,N_25907,N_25617);
nand U27785 (N_27785,N_26003,N_26681);
and U27786 (N_27786,N_26676,N_25927);
xnor U27787 (N_27787,N_26737,N_25595);
nand U27788 (N_27788,N_25722,N_26988);
nor U27789 (N_27789,N_26281,N_26783);
and U27790 (N_27790,N_26008,N_26893);
nand U27791 (N_27791,N_26961,N_26161);
xor U27792 (N_27792,N_26477,N_26884);
nor U27793 (N_27793,N_25656,N_26323);
and U27794 (N_27794,N_25678,N_26036);
and U27795 (N_27795,N_26317,N_26032);
or U27796 (N_27796,N_26827,N_26883);
nand U27797 (N_27797,N_25907,N_26602);
nor U27798 (N_27798,N_26404,N_26116);
or U27799 (N_27799,N_26708,N_25700);
xor U27800 (N_27800,N_26559,N_25542);
nor U27801 (N_27801,N_26856,N_26602);
xnor U27802 (N_27802,N_26237,N_26248);
nor U27803 (N_27803,N_26670,N_26068);
and U27804 (N_27804,N_26356,N_26074);
and U27805 (N_27805,N_26503,N_26070);
xnor U27806 (N_27806,N_26865,N_26179);
nor U27807 (N_27807,N_26691,N_26786);
nor U27808 (N_27808,N_26587,N_25625);
xnor U27809 (N_27809,N_26159,N_26012);
xor U27810 (N_27810,N_26095,N_26227);
nor U27811 (N_27811,N_25998,N_25879);
nor U27812 (N_27812,N_25531,N_25987);
and U27813 (N_27813,N_26357,N_25707);
nor U27814 (N_27814,N_25522,N_26345);
nand U27815 (N_27815,N_26023,N_26139);
and U27816 (N_27816,N_25811,N_26092);
and U27817 (N_27817,N_26558,N_26341);
nand U27818 (N_27818,N_26521,N_26974);
or U27819 (N_27819,N_26623,N_25722);
and U27820 (N_27820,N_25688,N_25993);
nand U27821 (N_27821,N_26104,N_25851);
or U27822 (N_27822,N_26039,N_25811);
and U27823 (N_27823,N_26830,N_26660);
nor U27824 (N_27824,N_26061,N_26534);
or U27825 (N_27825,N_26237,N_26724);
nor U27826 (N_27826,N_26361,N_26225);
or U27827 (N_27827,N_25548,N_26855);
or U27828 (N_27828,N_26444,N_26229);
and U27829 (N_27829,N_26983,N_26298);
xnor U27830 (N_27830,N_26127,N_25826);
nand U27831 (N_27831,N_26685,N_25937);
and U27832 (N_27832,N_26637,N_26097);
nor U27833 (N_27833,N_25951,N_25914);
and U27834 (N_27834,N_25869,N_26161);
and U27835 (N_27835,N_26049,N_26226);
nand U27836 (N_27836,N_26310,N_26270);
and U27837 (N_27837,N_25711,N_26815);
and U27838 (N_27838,N_26056,N_25618);
nor U27839 (N_27839,N_26911,N_25711);
nand U27840 (N_27840,N_26299,N_25965);
nand U27841 (N_27841,N_25880,N_25584);
nor U27842 (N_27842,N_26168,N_26483);
nand U27843 (N_27843,N_26317,N_26210);
nor U27844 (N_27844,N_26141,N_26337);
nand U27845 (N_27845,N_26215,N_26208);
xor U27846 (N_27846,N_26898,N_26434);
and U27847 (N_27847,N_26324,N_26967);
nand U27848 (N_27848,N_25640,N_26581);
and U27849 (N_27849,N_25888,N_25910);
xor U27850 (N_27850,N_25545,N_25660);
and U27851 (N_27851,N_25808,N_25977);
xor U27852 (N_27852,N_26448,N_26926);
nand U27853 (N_27853,N_26409,N_26518);
or U27854 (N_27854,N_26051,N_25852);
nor U27855 (N_27855,N_26350,N_25550);
nor U27856 (N_27856,N_26555,N_25726);
and U27857 (N_27857,N_26500,N_26387);
or U27858 (N_27858,N_25774,N_26743);
or U27859 (N_27859,N_25738,N_26424);
nand U27860 (N_27860,N_26318,N_25933);
and U27861 (N_27861,N_26004,N_25523);
nor U27862 (N_27862,N_26175,N_25853);
nor U27863 (N_27863,N_26901,N_25873);
or U27864 (N_27864,N_25969,N_26404);
or U27865 (N_27865,N_25520,N_26711);
and U27866 (N_27866,N_26175,N_26028);
nor U27867 (N_27867,N_25886,N_25990);
and U27868 (N_27868,N_26399,N_26203);
nor U27869 (N_27869,N_26485,N_26314);
and U27870 (N_27870,N_26883,N_25742);
nor U27871 (N_27871,N_26031,N_26039);
nand U27872 (N_27872,N_25844,N_26301);
nand U27873 (N_27873,N_26856,N_26322);
and U27874 (N_27874,N_26810,N_25652);
xnor U27875 (N_27875,N_25676,N_26862);
nand U27876 (N_27876,N_25579,N_26947);
nand U27877 (N_27877,N_26216,N_26764);
nor U27878 (N_27878,N_25730,N_25955);
nand U27879 (N_27879,N_26388,N_26090);
or U27880 (N_27880,N_26114,N_26163);
and U27881 (N_27881,N_26137,N_26841);
xnor U27882 (N_27882,N_26888,N_26235);
or U27883 (N_27883,N_25533,N_26282);
or U27884 (N_27884,N_25522,N_26757);
or U27885 (N_27885,N_26254,N_25821);
and U27886 (N_27886,N_25749,N_26250);
or U27887 (N_27887,N_25770,N_26124);
xor U27888 (N_27888,N_25912,N_26255);
xor U27889 (N_27889,N_26697,N_26133);
xnor U27890 (N_27890,N_25801,N_26700);
and U27891 (N_27891,N_25523,N_26003);
nand U27892 (N_27892,N_26897,N_25663);
or U27893 (N_27893,N_25682,N_26919);
xnor U27894 (N_27894,N_26312,N_25626);
and U27895 (N_27895,N_25694,N_25895);
and U27896 (N_27896,N_26779,N_26931);
or U27897 (N_27897,N_25895,N_25560);
xnor U27898 (N_27898,N_26653,N_25804);
xnor U27899 (N_27899,N_26086,N_25794);
nand U27900 (N_27900,N_25717,N_25948);
nor U27901 (N_27901,N_26139,N_25705);
xnor U27902 (N_27902,N_25602,N_26969);
or U27903 (N_27903,N_25913,N_25524);
nor U27904 (N_27904,N_25762,N_26797);
nor U27905 (N_27905,N_26632,N_26108);
xnor U27906 (N_27906,N_25509,N_25752);
xor U27907 (N_27907,N_26211,N_26621);
xor U27908 (N_27908,N_25583,N_25958);
or U27909 (N_27909,N_26217,N_25836);
and U27910 (N_27910,N_26701,N_25988);
and U27911 (N_27911,N_25632,N_26065);
nor U27912 (N_27912,N_26189,N_26663);
nand U27913 (N_27913,N_26761,N_25595);
or U27914 (N_27914,N_26122,N_25987);
nand U27915 (N_27915,N_26013,N_26981);
or U27916 (N_27916,N_26641,N_25510);
xnor U27917 (N_27917,N_25626,N_25709);
nor U27918 (N_27918,N_25877,N_26802);
nand U27919 (N_27919,N_26279,N_26592);
nand U27920 (N_27920,N_26717,N_26774);
nand U27921 (N_27921,N_26741,N_25855);
nor U27922 (N_27922,N_25541,N_26841);
nor U27923 (N_27923,N_26000,N_26089);
or U27924 (N_27924,N_26292,N_25628);
and U27925 (N_27925,N_26390,N_26174);
nand U27926 (N_27926,N_26368,N_26462);
and U27927 (N_27927,N_25758,N_26956);
and U27928 (N_27928,N_25842,N_25575);
nand U27929 (N_27929,N_26892,N_25968);
xor U27930 (N_27930,N_25784,N_25857);
and U27931 (N_27931,N_26683,N_26087);
nor U27932 (N_27932,N_26741,N_26988);
xor U27933 (N_27933,N_26645,N_26769);
xnor U27934 (N_27934,N_26901,N_25801);
xor U27935 (N_27935,N_26062,N_26574);
and U27936 (N_27936,N_25704,N_25665);
nand U27937 (N_27937,N_26251,N_25869);
and U27938 (N_27938,N_26775,N_26757);
xor U27939 (N_27939,N_25610,N_25929);
xor U27940 (N_27940,N_26526,N_25767);
nand U27941 (N_27941,N_26098,N_26736);
or U27942 (N_27942,N_25819,N_25522);
xor U27943 (N_27943,N_26067,N_25849);
xor U27944 (N_27944,N_26228,N_26782);
or U27945 (N_27945,N_26819,N_26091);
or U27946 (N_27946,N_26338,N_25877);
and U27947 (N_27947,N_25960,N_25999);
and U27948 (N_27948,N_25815,N_26468);
or U27949 (N_27949,N_26727,N_25968);
and U27950 (N_27950,N_25991,N_26474);
xnor U27951 (N_27951,N_25776,N_26678);
nor U27952 (N_27952,N_25894,N_25697);
nand U27953 (N_27953,N_26535,N_26782);
nand U27954 (N_27954,N_25917,N_25741);
and U27955 (N_27955,N_26177,N_26531);
nor U27956 (N_27956,N_26499,N_25858);
or U27957 (N_27957,N_26639,N_25835);
or U27958 (N_27958,N_26709,N_25784);
xor U27959 (N_27959,N_25608,N_25684);
and U27960 (N_27960,N_26392,N_26998);
xor U27961 (N_27961,N_26292,N_26457);
or U27962 (N_27962,N_25883,N_26347);
and U27963 (N_27963,N_25862,N_26335);
or U27964 (N_27964,N_25619,N_26865);
nor U27965 (N_27965,N_26536,N_26665);
or U27966 (N_27966,N_25603,N_26710);
nor U27967 (N_27967,N_26871,N_26813);
nand U27968 (N_27968,N_25694,N_25768);
nor U27969 (N_27969,N_26183,N_26801);
nor U27970 (N_27970,N_26891,N_25512);
nand U27971 (N_27971,N_26962,N_26006);
nor U27972 (N_27972,N_25643,N_25571);
xnor U27973 (N_27973,N_26826,N_25525);
xor U27974 (N_27974,N_26245,N_25920);
nor U27975 (N_27975,N_25942,N_26283);
xnor U27976 (N_27976,N_26222,N_26491);
or U27977 (N_27977,N_25695,N_26893);
or U27978 (N_27978,N_26496,N_26568);
or U27979 (N_27979,N_26107,N_26034);
nand U27980 (N_27980,N_25702,N_26369);
or U27981 (N_27981,N_26502,N_25923);
and U27982 (N_27982,N_26939,N_26748);
or U27983 (N_27983,N_26699,N_26337);
and U27984 (N_27984,N_26708,N_26745);
xor U27985 (N_27985,N_26133,N_25812);
xnor U27986 (N_27986,N_26558,N_26333);
nor U27987 (N_27987,N_26668,N_25732);
nor U27988 (N_27988,N_25984,N_26076);
nor U27989 (N_27989,N_26191,N_26400);
nor U27990 (N_27990,N_26786,N_25620);
nor U27991 (N_27991,N_26976,N_25503);
nand U27992 (N_27992,N_26905,N_26691);
nor U27993 (N_27993,N_26529,N_25887);
nand U27994 (N_27994,N_26015,N_26167);
or U27995 (N_27995,N_26586,N_25599);
and U27996 (N_27996,N_25588,N_26106);
nand U27997 (N_27997,N_26907,N_26303);
xor U27998 (N_27998,N_26674,N_26839);
and U27999 (N_27999,N_26016,N_25565);
nand U28000 (N_28000,N_25752,N_26412);
and U28001 (N_28001,N_26449,N_26081);
xnor U28002 (N_28002,N_25893,N_26637);
nor U28003 (N_28003,N_26431,N_26781);
nor U28004 (N_28004,N_25565,N_25981);
and U28005 (N_28005,N_25736,N_26674);
nor U28006 (N_28006,N_26934,N_26259);
xor U28007 (N_28007,N_25684,N_26404);
nor U28008 (N_28008,N_25643,N_26833);
and U28009 (N_28009,N_25760,N_26168);
xor U28010 (N_28010,N_25527,N_26459);
or U28011 (N_28011,N_26693,N_25536);
or U28012 (N_28012,N_25927,N_25855);
and U28013 (N_28013,N_26470,N_26827);
xor U28014 (N_28014,N_25668,N_26210);
nand U28015 (N_28015,N_26657,N_25629);
xor U28016 (N_28016,N_25772,N_26088);
or U28017 (N_28017,N_25917,N_26678);
or U28018 (N_28018,N_25807,N_25986);
or U28019 (N_28019,N_25780,N_26981);
and U28020 (N_28020,N_25774,N_25621);
nor U28021 (N_28021,N_26844,N_25683);
xnor U28022 (N_28022,N_26420,N_26547);
nor U28023 (N_28023,N_26882,N_26088);
or U28024 (N_28024,N_26860,N_26116);
nand U28025 (N_28025,N_25624,N_25597);
nand U28026 (N_28026,N_26012,N_26772);
or U28027 (N_28027,N_25556,N_26898);
nand U28028 (N_28028,N_25645,N_26031);
xor U28029 (N_28029,N_25583,N_26743);
nand U28030 (N_28030,N_26078,N_25942);
xnor U28031 (N_28031,N_25750,N_26579);
nand U28032 (N_28032,N_26709,N_25832);
nor U28033 (N_28033,N_26464,N_25917);
xnor U28034 (N_28034,N_25567,N_26234);
nor U28035 (N_28035,N_26310,N_26885);
xor U28036 (N_28036,N_26588,N_26081);
or U28037 (N_28037,N_26870,N_26200);
xor U28038 (N_28038,N_25925,N_26317);
or U28039 (N_28039,N_25647,N_25765);
nand U28040 (N_28040,N_26689,N_26814);
and U28041 (N_28041,N_26456,N_26719);
nor U28042 (N_28042,N_25863,N_26628);
or U28043 (N_28043,N_26538,N_26519);
and U28044 (N_28044,N_26119,N_25720);
or U28045 (N_28045,N_26805,N_25621);
nand U28046 (N_28046,N_26108,N_26216);
nand U28047 (N_28047,N_26421,N_26026);
nor U28048 (N_28048,N_26715,N_25733);
nand U28049 (N_28049,N_26732,N_26710);
nor U28050 (N_28050,N_26769,N_26013);
nand U28051 (N_28051,N_26379,N_26771);
nor U28052 (N_28052,N_26021,N_26162);
or U28053 (N_28053,N_26908,N_25635);
and U28054 (N_28054,N_26207,N_26070);
and U28055 (N_28055,N_25559,N_26964);
xnor U28056 (N_28056,N_26896,N_26673);
nor U28057 (N_28057,N_25840,N_26484);
nor U28058 (N_28058,N_26898,N_26011);
nor U28059 (N_28059,N_25631,N_25776);
nor U28060 (N_28060,N_26872,N_26400);
nor U28061 (N_28061,N_26729,N_26630);
or U28062 (N_28062,N_26107,N_26106);
xor U28063 (N_28063,N_26776,N_26794);
or U28064 (N_28064,N_26110,N_25700);
nand U28065 (N_28065,N_26023,N_26300);
nand U28066 (N_28066,N_26611,N_26661);
nand U28067 (N_28067,N_26328,N_26699);
or U28068 (N_28068,N_25960,N_25519);
nand U28069 (N_28069,N_25841,N_25519);
nor U28070 (N_28070,N_26045,N_26437);
and U28071 (N_28071,N_26767,N_25640);
or U28072 (N_28072,N_26087,N_26498);
and U28073 (N_28073,N_26965,N_26556);
or U28074 (N_28074,N_25861,N_25987);
nor U28075 (N_28075,N_25542,N_26429);
or U28076 (N_28076,N_26284,N_26431);
xnor U28077 (N_28077,N_26502,N_25705);
xor U28078 (N_28078,N_26771,N_26557);
and U28079 (N_28079,N_25985,N_26391);
nor U28080 (N_28080,N_26181,N_26758);
nand U28081 (N_28081,N_25909,N_26878);
and U28082 (N_28082,N_26378,N_26549);
xnor U28083 (N_28083,N_26939,N_26894);
nand U28084 (N_28084,N_25823,N_25557);
and U28085 (N_28085,N_26963,N_25851);
and U28086 (N_28086,N_26938,N_26491);
nor U28087 (N_28087,N_25576,N_26399);
and U28088 (N_28088,N_25663,N_25963);
or U28089 (N_28089,N_26254,N_26504);
nor U28090 (N_28090,N_25608,N_26040);
and U28091 (N_28091,N_26686,N_26467);
xnor U28092 (N_28092,N_26861,N_25815);
or U28093 (N_28093,N_25827,N_26727);
nor U28094 (N_28094,N_26924,N_26428);
and U28095 (N_28095,N_26286,N_26702);
nor U28096 (N_28096,N_26086,N_25944);
and U28097 (N_28097,N_26124,N_26351);
nor U28098 (N_28098,N_25772,N_26588);
xnor U28099 (N_28099,N_26202,N_26455);
xor U28100 (N_28100,N_26843,N_25782);
and U28101 (N_28101,N_26485,N_26794);
xnor U28102 (N_28102,N_26324,N_25955);
and U28103 (N_28103,N_26536,N_26892);
xor U28104 (N_28104,N_26571,N_26368);
xor U28105 (N_28105,N_26225,N_25751);
or U28106 (N_28106,N_25999,N_25857);
nor U28107 (N_28107,N_25787,N_26336);
nand U28108 (N_28108,N_25748,N_26331);
and U28109 (N_28109,N_26840,N_26686);
nor U28110 (N_28110,N_26583,N_26371);
xnor U28111 (N_28111,N_26896,N_26642);
nor U28112 (N_28112,N_26641,N_26336);
xor U28113 (N_28113,N_26291,N_26989);
nand U28114 (N_28114,N_25855,N_25723);
xor U28115 (N_28115,N_26212,N_25519);
nor U28116 (N_28116,N_26615,N_26315);
or U28117 (N_28117,N_25894,N_25575);
nor U28118 (N_28118,N_26940,N_26546);
or U28119 (N_28119,N_25829,N_25967);
nand U28120 (N_28120,N_26186,N_25744);
or U28121 (N_28121,N_26745,N_26057);
xor U28122 (N_28122,N_26224,N_26751);
nand U28123 (N_28123,N_26378,N_26160);
nand U28124 (N_28124,N_26609,N_26817);
or U28125 (N_28125,N_25922,N_26999);
and U28126 (N_28126,N_26230,N_26393);
xor U28127 (N_28127,N_25905,N_26633);
nor U28128 (N_28128,N_26877,N_25527);
nor U28129 (N_28129,N_26495,N_26705);
and U28130 (N_28130,N_26339,N_25971);
nor U28131 (N_28131,N_26252,N_26466);
or U28132 (N_28132,N_26117,N_25968);
nand U28133 (N_28133,N_26335,N_26504);
or U28134 (N_28134,N_25767,N_26611);
and U28135 (N_28135,N_26546,N_26277);
xnor U28136 (N_28136,N_25723,N_26333);
nand U28137 (N_28137,N_25586,N_26664);
xor U28138 (N_28138,N_26416,N_26418);
nand U28139 (N_28139,N_25547,N_25736);
nand U28140 (N_28140,N_25866,N_26054);
or U28141 (N_28141,N_26278,N_26314);
and U28142 (N_28142,N_25546,N_26159);
or U28143 (N_28143,N_25937,N_25964);
nand U28144 (N_28144,N_26204,N_26767);
xor U28145 (N_28145,N_26322,N_26230);
and U28146 (N_28146,N_25692,N_26199);
and U28147 (N_28147,N_26863,N_26777);
nor U28148 (N_28148,N_25866,N_26756);
or U28149 (N_28149,N_26149,N_25634);
and U28150 (N_28150,N_26322,N_25953);
nor U28151 (N_28151,N_26337,N_26793);
xor U28152 (N_28152,N_26027,N_25980);
and U28153 (N_28153,N_26818,N_25941);
nor U28154 (N_28154,N_26821,N_26192);
and U28155 (N_28155,N_26951,N_25682);
nand U28156 (N_28156,N_25996,N_26912);
and U28157 (N_28157,N_26278,N_26977);
or U28158 (N_28158,N_25815,N_26333);
nor U28159 (N_28159,N_26284,N_26922);
xor U28160 (N_28160,N_25933,N_26562);
xor U28161 (N_28161,N_26248,N_26198);
and U28162 (N_28162,N_26001,N_26369);
xnor U28163 (N_28163,N_25881,N_25537);
and U28164 (N_28164,N_26587,N_26061);
nor U28165 (N_28165,N_26946,N_25655);
xnor U28166 (N_28166,N_26230,N_26130);
or U28167 (N_28167,N_26172,N_25547);
and U28168 (N_28168,N_26130,N_26564);
xnor U28169 (N_28169,N_25581,N_25936);
or U28170 (N_28170,N_26496,N_26155);
nand U28171 (N_28171,N_26087,N_26186);
nor U28172 (N_28172,N_26790,N_26091);
or U28173 (N_28173,N_26529,N_25502);
or U28174 (N_28174,N_26918,N_25902);
xor U28175 (N_28175,N_25633,N_25783);
nor U28176 (N_28176,N_25800,N_25656);
and U28177 (N_28177,N_26554,N_25816);
and U28178 (N_28178,N_26348,N_26804);
or U28179 (N_28179,N_25655,N_25851);
nor U28180 (N_28180,N_26196,N_25956);
and U28181 (N_28181,N_25598,N_26520);
nand U28182 (N_28182,N_26652,N_26797);
nand U28183 (N_28183,N_26460,N_25622);
and U28184 (N_28184,N_26063,N_26669);
and U28185 (N_28185,N_25924,N_25630);
and U28186 (N_28186,N_26475,N_26450);
nand U28187 (N_28187,N_26468,N_26805);
nand U28188 (N_28188,N_26837,N_26771);
nand U28189 (N_28189,N_26407,N_26026);
and U28190 (N_28190,N_26955,N_26296);
xor U28191 (N_28191,N_26497,N_26981);
or U28192 (N_28192,N_26279,N_26260);
or U28193 (N_28193,N_25544,N_26940);
nand U28194 (N_28194,N_25721,N_26826);
xor U28195 (N_28195,N_26632,N_26851);
and U28196 (N_28196,N_26798,N_25516);
or U28197 (N_28197,N_26391,N_25873);
or U28198 (N_28198,N_25751,N_26016);
nand U28199 (N_28199,N_25500,N_26146);
nor U28200 (N_28200,N_26728,N_26112);
nand U28201 (N_28201,N_26152,N_25656);
and U28202 (N_28202,N_25915,N_26120);
nor U28203 (N_28203,N_26338,N_26025);
nand U28204 (N_28204,N_25530,N_26726);
xnor U28205 (N_28205,N_26689,N_26646);
xnor U28206 (N_28206,N_25800,N_25573);
or U28207 (N_28207,N_25842,N_25655);
xnor U28208 (N_28208,N_26223,N_26758);
and U28209 (N_28209,N_25507,N_26564);
or U28210 (N_28210,N_25690,N_25759);
or U28211 (N_28211,N_26987,N_26687);
or U28212 (N_28212,N_25556,N_26643);
or U28213 (N_28213,N_26016,N_25726);
nor U28214 (N_28214,N_26653,N_25851);
nand U28215 (N_28215,N_25912,N_26941);
and U28216 (N_28216,N_25897,N_26197);
nor U28217 (N_28217,N_26443,N_26920);
nor U28218 (N_28218,N_25693,N_25852);
and U28219 (N_28219,N_25968,N_26122);
or U28220 (N_28220,N_26642,N_26672);
xnor U28221 (N_28221,N_26264,N_26448);
nor U28222 (N_28222,N_26938,N_26036);
nand U28223 (N_28223,N_26505,N_25836);
and U28224 (N_28224,N_26602,N_26502);
nor U28225 (N_28225,N_26719,N_26797);
and U28226 (N_28226,N_26308,N_26370);
nor U28227 (N_28227,N_26419,N_26534);
and U28228 (N_28228,N_26840,N_26084);
nand U28229 (N_28229,N_26949,N_25928);
xor U28230 (N_28230,N_26336,N_26487);
nor U28231 (N_28231,N_26116,N_25802);
xnor U28232 (N_28232,N_26381,N_26719);
nand U28233 (N_28233,N_26063,N_26970);
xor U28234 (N_28234,N_26856,N_26079);
nand U28235 (N_28235,N_26032,N_26741);
nor U28236 (N_28236,N_26114,N_26586);
and U28237 (N_28237,N_26652,N_26733);
nor U28238 (N_28238,N_26847,N_25552);
or U28239 (N_28239,N_26729,N_26134);
and U28240 (N_28240,N_25974,N_25979);
xor U28241 (N_28241,N_26609,N_25848);
nand U28242 (N_28242,N_26367,N_26589);
xor U28243 (N_28243,N_25574,N_26173);
xnor U28244 (N_28244,N_25577,N_26724);
nand U28245 (N_28245,N_25953,N_25884);
nand U28246 (N_28246,N_26628,N_26789);
or U28247 (N_28247,N_26630,N_26551);
nand U28248 (N_28248,N_26805,N_25817);
or U28249 (N_28249,N_25660,N_26818);
or U28250 (N_28250,N_26576,N_26423);
or U28251 (N_28251,N_25532,N_26538);
and U28252 (N_28252,N_25632,N_26836);
nand U28253 (N_28253,N_26695,N_26941);
nor U28254 (N_28254,N_26689,N_26300);
nor U28255 (N_28255,N_26442,N_26478);
or U28256 (N_28256,N_26285,N_25732);
nor U28257 (N_28257,N_26040,N_26075);
or U28258 (N_28258,N_26536,N_25820);
nand U28259 (N_28259,N_25620,N_26029);
xor U28260 (N_28260,N_26316,N_26771);
and U28261 (N_28261,N_26078,N_25680);
and U28262 (N_28262,N_26893,N_26984);
xnor U28263 (N_28263,N_25749,N_26427);
or U28264 (N_28264,N_25857,N_26946);
or U28265 (N_28265,N_26221,N_26323);
and U28266 (N_28266,N_26708,N_26910);
or U28267 (N_28267,N_26765,N_25891);
or U28268 (N_28268,N_26758,N_26386);
or U28269 (N_28269,N_25833,N_26424);
nand U28270 (N_28270,N_25992,N_26594);
nand U28271 (N_28271,N_26971,N_26290);
or U28272 (N_28272,N_25852,N_25525);
nand U28273 (N_28273,N_26715,N_26954);
nand U28274 (N_28274,N_25731,N_26587);
nor U28275 (N_28275,N_26086,N_25880);
or U28276 (N_28276,N_26201,N_25699);
or U28277 (N_28277,N_26458,N_26843);
or U28278 (N_28278,N_25569,N_26672);
xnor U28279 (N_28279,N_26460,N_25811);
and U28280 (N_28280,N_25599,N_26833);
xnor U28281 (N_28281,N_25797,N_26253);
nand U28282 (N_28282,N_26717,N_26849);
or U28283 (N_28283,N_26969,N_26339);
nor U28284 (N_28284,N_25535,N_26064);
or U28285 (N_28285,N_26592,N_26839);
nor U28286 (N_28286,N_25839,N_26517);
and U28287 (N_28287,N_26695,N_25729);
nand U28288 (N_28288,N_26179,N_26528);
and U28289 (N_28289,N_26098,N_25669);
or U28290 (N_28290,N_26757,N_25564);
or U28291 (N_28291,N_25840,N_26338);
nor U28292 (N_28292,N_25698,N_25800);
xnor U28293 (N_28293,N_25509,N_26987);
or U28294 (N_28294,N_26069,N_26075);
or U28295 (N_28295,N_26109,N_26564);
or U28296 (N_28296,N_25876,N_26167);
and U28297 (N_28297,N_25721,N_26236);
nand U28298 (N_28298,N_26694,N_25665);
or U28299 (N_28299,N_26634,N_25838);
nor U28300 (N_28300,N_26247,N_25804);
or U28301 (N_28301,N_26676,N_26733);
xor U28302 (N_28302,N_26424,N_25933);
nand U28303 (N_28303,N_25916,N_26248);
and U28304 (N_28304,N_26324,N_26860);
and U28305 (N_28305,N_25917,N_26350);
nand U28306 (N_28306,N_26132,N_26670);
nor U28307 (N_28307,N_25664,N_26665);
nor U28308 (N_28308,N_26878,N_26292);
nand U28309 (N_28309,N_26214,N_26301);
or U28310 (N_28310,N_26124,N_26978);
and U28311 (N_28311,N_26326,N_26333);
nand U28312 (N_28312,N_26421,N_26977);
nor U28313 (N_28313,N_25612,N_25956);
nand U28314 (N_28314,N_26396,N_26860);
xnor U28315 (N_28315,N_26804,N_25561);
nand U28316 (N_28316,N_26407,N_26319);
or U28317 (N_28317,N_26001,N_26411);
nand U28318 (N_28318,N_26938,N_25857);
and U28319 (N_28319,N_25699,N_26968);
xnor U28320 (N_28320,N_26914,N_26898);
and U28321 (N_28321,N_25894,N_26974);
nor U28322 (N_28322,N_26501,N_26513);
and U28323 (N_28323,N_26774,N_26287);
and U28324 (N_28324,N_26620,N_26211);
or U28325 (N_28325,N_26629,N_26185);
and U28326 (N_28326,N_26170,N_26617);
nor U28327 (N_28327,N_26550,N_26551);
xnor U28328 (N_28328,N_26275,N_25728);
xor U28329 (N_28329,N_26196,N_26002);
nand U28330 (N_28330,N_25723,N_25542);
xor U28331 (N_28331,N_26432,N_26569);
and U28332 (N_28332,N_25593,N_25912);
nand U28333 (N_28333,N_25686,N_25702);
nand U28334 (N_28334,N_25696,N_26551);
or U28335 (N_28335,N_26696,N_25995);
nand U28336 (N_28336,N_26059,N_25629);
nor U28337 (N_28337,N_26014,N_25681);
and U28338 (N_28338,N_26027,N_25765);
nor U28339 (N_28339,N_25863,N_26768);
xnor U28340 (N_28340,N_26898,N_26154);
xnor U28341 (N_28341,N_25884,N_26191);
or U28342 (N_28342,N_25850,N_25918);
nor U28343 (N_28343,N_26985,N_26336);
and U28344 (N_28344,N_26889,N_25559);
nor U28345 (N_28345,N_25900,N_26903);
and U28346 (N_28346,N_25777,N_26992);
or U28347 (N_28347,N_26060,N_25749);
and U28348 (N_28348,N_26939,N_26201);
nand U28349 (N_28349,N_25584,N_26165);
nand U28350 (N_28350,N_25612,N_25782);
nand U28351 (N_28351,N_26502,N_26103);
nor U28352 (N_28352,N_26168,N_26037);
xor U28353 (N_28353,N_26124,N_25821);
xnor U28354 (N_28354,N_26513,N_26379);
or U28355 (N_28355,N_25851,N_26220);
xor U28356 (N_28356,N_25654,N_25981);
and U28357 (N_28357,N_26016,N_26484);
and U28358 (N_28358,N_26078,N_25884);
and U28359 (N_28359,N_26893,N_26475);
nor U28360 (N_28360,N_25649,N_25665);
or U28361 (N_28361,N_25621,N_26323);
nor U28362 (N_28362,N_26227,N_26591);
nand U28363 (N_28363,N_26832,N_25772);
or U28364 (N_28364,N_26197,N_26438);
xor U28365 (N_28365,N_26008,N_26968);
or U28366 (N_28366,N_26895,N_26764);
xor U28367 (N_28367,N_26230,N_25966);
nand U28368 (N_28368,N_25675,N_26347);
xor U28369 (N_28369,N_26901,N_25665);
nor U28370 (N_28370,N_25778,N_25583);
and U28371 (N_28371,N_26931,N_26923);
xnor U28372 (N_28372,N_26153,N_26689);
nor U28373 (N_28373,N_26366,N_25751);
nand U28374 (N_28374,N_26357,N_25833);
or U28375 (N_28375,N_25611,N_25938);
and U28376 (N_28376,N_25758,N_25875);
xor U28377 (N_28377,N_25981,N_25761);
nand U28378 (N_28378,N_26792,N_26884);
xor U28379 (N_28379,N_26220,N_26498);
and U28380 (N_28380,N_26006,N_25613);
nor U28381 (N_28381,N_26337,N_26326);
nor U28382 (N_28382,N_26918,N_26926);
or U28383 (N_28383,N_26895,N_25923);
nand U28384 (N_28384,N_26643,N_26379);
xnor U28385 (N_28385,N_25537,N_26350);
nand U28386 (N_28386,N_25942,N_26478);
and U28387 (N_28387,N_25978,N_26197);
nand U28388 (N_28388,N_26696,N_26981);
nand U28389 (N_28389,N_25919,N_25883);
and U28390 (N_28390,N_26369,N_26086);
nor U28391 (N_28391,N_26892,N_25826);
xor U28392 (N_28392,N_26146,N_26073);
or U28393 (N_28393,N_26561,N_26949);
or U28394 (N_28394,N_25745,N_26892);
nor U28395 (N_28395,N_25825,N_25505);
nand U28396 (N_28396,N_25789,N_26854);
nor U28397 (N_28397,N_26149,N_26802);
nand U28398 (N_28398,N_26964,N_26218);
xnor U28399 (N_28399,N_26278,N_26162);
nand U28400 (N_28400,N_26678,N_26104);
and U28401 (N_28401,N_26819,N_26673);
nand U28402 (N_28402,N_26284,N_26994);
and U28403 (N_28403,N_25719,N_26205);
or U28404 (N_28404,N_25576,N_26589);
or U28405 (N_28405,N_26991,N_25694);
nand U28406 (N_28406,N_26620,N_26161);
nor U28407 (N_28407,N_26486,N_26816);
and U28408 (N_28408,N_26276,N_25708);
nor U28409 (N_28409,N_25721,N_26547);
and U28410 (N_28410,N_25598,N_25680);
xnor U28411 (N_28411,N_26624,N_25547);
nand U28412 (N_28412,N_25701,N_26846);
xor U28413 (N_28413,N_25685,N_26283);
or U28414 (N_28414,N_26621,N_26278);
or U28415 (N_28415,N_26039,N_26898);
nand U28416 (N_28416,N_26516,N_26544);
nor U28417 (N_28417,N_25758,N_26962);
xnor U28418 (N_28418,N_26555,N_26494);
nor U28419 (N_28419,N_26455,N_26163);
xor U28420 (N_28420,N_25604,N_25556);
and U28421 (N_28421,N_26491,N_26116);
nor U28422 (N_28422,N_26902,N_26369);
nor U28423 (N_28423,N_26956,N_25587);
or U28424 (N_28424,N_26749,N_26112);
or U28425 (N_28425,N_25871,N_26011);
xor U28426 (N_28426,N_26459,N_26546);
and U28427 (N_28427,N_26324,N_25961);
nor U28428 (N_28428,N_25628,N_26121);
xnor U28429 (N_28429,N_25728,N_26627);
and U28430 (N_28430,N_26232,N_25557);
nand U28431 (N_28431,N_26010,N_25876);
nor U28432 (N_28432,N_26790,N_26090);
or U28433 (N_28433,N_25999,N_25965);
nor U28434 (N_28434,N_26906,N_25684);
and U28435 (N_28435,N_26241,N_25565);
xnor U28436 (N_28436,N_26469,N_25688);
or U28437 (N_28437,N_26824,N_25982);
or U28438 (N_28438,N_25968,N_26550);
nand U28439 (N_28439,N_25853,N_26484);
nand U28440 (N_28440,N_25960,N_26891);
nand U28441 (N_28441,N_26026,N_26093);
nor U28442 (N_28442,N_25873,N_25943);
nor U28443 (N_28443,N_26139,N_26834);
and U28444 (N_28444,N_26384,N_26088);
nor U28445 (N_28445,N_26243,N_26315);
or U28446 (N_28446,N_26410,N_25677);
and U28447 (N_28447,N_26587,N_26491);
or U28448 (N_28448,N_26830,N_26885);
or U28449 (N_28449,N_26719,N_26700);
nand U28450 (N_28450,N_25858,N_25919);
nand U28451 (N_28451,N_26959,N_26448);
xor U28452 (N_28452,N_26973,N_26631);
nand U28453 (N_28453,N_26420,N_26417);
nand U28454 (N_28454,N_25531,N_26009);
and U28455 (N_28455,N_26298,N_26151);
or U28456 (N_28456,N_26692,N_25688);
or U28457 (N_28457,N_25629,N_25572);
and U28458 (N_28458,N_26847,N_25695);
nand U28459 (N_28459,N_25896,N_26141);
xnor U28460 (N_28460,N_26887,N_26066);
xnor U28461 (N_28461,N_25826,N_26898);
nand U28462 (N_28462,N_26066,N_26858);
and U28463 (N_28463,N_26603,N_26935);
nand U28464 (N_28464,N_26454,N_26252);
and U28465 (N_28465,N_26625,N_26915);
xnor U28466 (N_28466,N_26438,N_25926);
xor U28467 (N_28467,N_25595,N_26040);
and U28468 (N_28468,N_25510,N_25952);
or U28469 (N_28469,N_25524,N_25705);
xor U28470 (N_28470,N_26080,N_26323);
and U28471 (N_28471,N_26581,N_26589);
nor U28472 (N_28472,N_25659,N_26870);
and U28473 (N_28473,N_26118,N_26827);
xnor U28474 (N_28474,N_25982,N_25535);
nor U28475 (N_28475,N_26129,N_26773);
xor U28476 (N_28476,N_26214,N_26138);
or U28477 (N_28477,N_26612,N_25941);
nand U28478 (N_28478,N_26409,N_25518);
xnor U28479 (N_28479,N_25550,N_26305);
or U28480 (N_28480,N_25696,N_25688);
xnor U28481 (N_28481,N_26838,N_25992);
nor U28482 (N_28482,N_25749,N_25911);
xnor U28483 (N_28483,N_25534,N_26939);
nor U28484 (N_28484,N_26037,N_26817);
nor U28485 (N_28485,N_25509,N_26023);
nand U28486 (N_28486,N_26896,N_26380);
or U28487 (N_28487,N_25756,N_26440);
and U28488 (N_28488,N_26808,N_25590);
nand U28489 (N_28489,N_26559,N_25689);
or U28490 (N_28490,N_26717,N_26674);
nand U28491 (N_28491,N_26803,N_26035);
and U28492 (N_28492,N_26761,N_26210);
and U28493 (N_28493,N_26677,N_26478);
or U28494 (N_28494,N_26785,N_26542);
xnor U28495 (N_28495,N_26284,N_26398);
nor U28496 (N_28496,N_26943,N_25857);
and U28497 (N_28497,N_26380,N_25965);
or U28498 (N_28498,N_26318,N_26550);
xor U28499 (N_28499,N_26657,N_25869);
nor U28500 (N_28500,N_28261,N_28425);
or U28501 (N_28501,N_27039,N_28436);
nor U28502 (N_28502,N_27352,N_27622);
nand U28503 (N_28503,N_27569,N_28259);
xor U28504 (N_28504,N_27477,N_27858);
xnor U28505 (N_28505,N_27925,N_28050);
xor U28506 (N_28506,N_27889,N_27559);
or U28507 (N_28507,N_27608,N_27680);
xor U28508 (N_28508,N_28208,N_27376);
and U28509 (N_28509,N_27076,N_28032);
xnor U28510 (N_28510,N_27388,N_27068);
nor U28511 (N_28511,N_27747,N_28122);
and U28512 (N_28512,N_28056,N_28090);
nor U28513 (N_28513,N_27755,N_27854);
and U28514 (N_28514,N_27651,N_27861);
and U28515 (N_28515,N_27379,N_28179);
or U28516 (N_28516,N_27247,N_27494);
nand U28517 (N_28517,N_27804,N_28166);
xor U28518 (N_28518,N_28458,N_27879);
xnor U28519 (N_28519,N_27295,N_27079);
nor U28520 (N_28520,N_27703,N_28428);
and U28521 (N_28521,N_27705,N_28117);
and U28522 (N_28522,N_28078,N_27081);
nand U28523 (N_28523,N_28235,N_28393);
nand U28524 (N_28524,N_27003,N_27387);
and U28525 (N_28525,N_27899,N_27211);
xnor U28526 (N_28526,N_27083,N_27772);
or U28527 (N_28527,N_27245,N_27360);
nand U28528 (N_28528,N_27226,N_28073);
nor U28529 (N_28529,N_28465,N_28402);
xnor U28530 (N_28530,N_28283,N_27687);
nor U28531 (N_28531,N_27600,N_28102);
nand U28532 (N_28532,N_27582,N_28316);
nor U28533 (N_28533,N_28471,N_28332);
nor U28534 (N_28534,N_28443,N_28497);
or U28535 (N_28535,N_27575,N_27759);
or U28536 (N_28536,N_28315,N_27048);
and U28537 (N_28537,N_28192,N_28335);
or U28538 (N_28538,N_27589,N_27908);
or U28539 (N_28539,N_27669,N_27035);
and U28540 (N_28540,N_27512,N_27056);
xnor U28541 (N_28541,N_27993,N_27746);
nor U28542 (N_28542,N_28293,N_27710);
and U28543 (N_28543,N_28416,N_27002);
xor U28544 (N_28544,N_27151,N_28387);
xor U28545 (N_28545,N_27796,N_28077);
xnor U28546 (N_28546,N_27124,N_27317);
nor U28547 (N_28547,N_28152,N_27574);
nor U28548 (N_28548,N_28239,N_27538);
or U28549 (N_28549,N_27610,N_27536);
or U28550 (N_28550,N_28210,N_27163);
xor U28551 (N_28551,N_27458,N_28388);
nor U28552 (N_28552,N_27541,N_28064);
or U28553 (N_28553,N_28414,N_27122);
and U28554 (N_28554,N_28009,N_27304);
xnor U28555 (N_28555,N_27970,N_28422);
and U28556 (N_28556,N_27135,N_27094);
xor U28557 (N_28557,N_27902,N_28184);
or U28558 (N_28558,N_27969,N_28492);
xor U28559 (N_28559,N_28437,N_28108);
xnor U28560 (N_28560,N_27773,N_28014);
xor U28561 (N_28561,N_27121,N_28251);
or U28562 (N_28562,N_27229,N_27040);
or U28563 (N_28563,N_28389,N_28035);
and U28564 (N_28564,N_27242,N_27402);
nand U28565 (N_28565,N_27797,N_27867);
nor U28566 (N_28566,N_27486,N_27767);
and U28567 (N_28567,N_27639,N_28361);
and U28568 (N_28568,N_28027,N_27953);
xor U28569 (N_28569,N_27143,N_27614);
xor U28570 (N_28570,N_27333,N_28354);
and U28571 (N_28571,N_28325,N_28442);
xor U28572 (N_28572,N_28131,N_27105);
nor U28573 (N_28573,N_27375,N_28397);
and U28574 (N_28574,N_27307,N_28198);
and U28575 (N_28575,N_27633,N_27434);
nand U28576 (N_28576,N_27848,N_27213);
nand U28577 (N_28577,N_28417,N_28299);
and U28578 (N_28578,N_27413,N_27373);
nor U28579 (N_28579,N_27996,N_28226);
nand U28580 (N_28580,N_27266,N_27482);
xnor U28581 (N_28581,N_27252,N_27337);
nor U28582 (N_28582,N_27189,N_27812);
and U28583 (N_28583,N_27906,N_27236);
nand U28584 (N_28584,N_27133,N_28341);
xnor U28585 (N_28585,N_28279,N_28182);
or U28586 (N_28586,N_28106,N_27684);
xnor U28587 (N_28587,N_28221,N_27273);
and U28588 (N_28588,N_27297,N_27693);
nand U28589 (N_28589,N_27112,N_27845);
xor U28590 (N_28590,N_28395,N_27876);
nor U28591 (N_28591,N_28323,N_27829);
xor U28592 (N_28592,N_27464,N_27734);
nand U28593 (N_28593,N_28159,N_27285);
xnor U28594 (N_28594,N_27038,N_27983);
nor U28595 (N_28595,N_27393,N_27731);
and U28596 (N_28596,N_27543,N_27186);
and U28597 (N_28597,N_27430,N_28476);
or U28598 (N_28598,N_27066,N_27502);
or U28599 (N_28599,N_28445,N_27480);
or U28600 (N_28600,N_28270,N_27111);
nor U28601 (N_28601,N_27517,N_27113);
nand U28602 (N_28602,N_28352,N_27706);
xnor U28603 (N_28603,N_27946,N_27564);
and U28604 (N_28604,N_28263,N_27293);
or U28605 (N_28605,N_27802,N_27863);
nand U28606 (N_28606,N_28432,N_28330);
or U28607 (N_28607,N_27271,N_27104);
and U28608 (N_28608,N_27315,N_27274);
nand U28609 (N_28609,N_27001,N_27888);
or U28610 (N_28610,N_27287,N_27780);
nand U28611 (N_28611,N_27649,N_28438);
nor U28612 (N_28612,N_28236,N_27819);
nand U28613 (N_28613,N_27859,N_27279);
and U28614 (N_28614,N_27426,N_27881);
and U28615 (N_28615,N_27585,N_28135);
or U28616 (N_28616,N_28154,N_27913);
nand U28617 (N_28617,N_27192,N_28282);
xor U28618 (N_28618,N_27688,N_27563);
or U28619 (N_28619,N_28088,N_27629);
xor U28620 (N_28620,N_27696,N_27851);
nor U28621 (N_28621,N_27220,N_27123);
xnor U28622 (N_28622,N_27624,N_27846);
and U28623 (N_28623,N_28322,N_27768);
xnor U28624 (N_28624,N_27978,N_28392);
and U28625 (N_28625,N_27074,N_28362);
nand U28626 (N_28626,N_27209,N_27644);
xnor U28627 (N_28627,N_28300,N_28136);
nor U28628 (N_28628,N_27254,N_28123);
nand U28629 (N_28629,N_27397,N_27020);
or U28630 (N_28630,N_28006,N_27514);
nand U28631 (N_28631,N_27055,N_28133);
nand U28632 (N_28632,N_27880,N_28305);
or U28633 (N_28633,N_27544,N_27325);
or U28634 (N_28634,N_28256,N_27241);
and U28635 (N_28635,N_27724,N_27518);
or U28636 (N_28636,N_27704,N_27914);
or U28637 (N_28637,N_27896,N_27436);
nor U28638 (N_28638,N_27939,N_28399);
and U28639 (N_28639,N_27128,N_28241);
and U28640 (N_28640,N_27363,N_27918);
nor U28641 (N_28641,N_27515,N_27386);
or U28642 (N_28642,N_27659,N_27184);
and U28643 (N_28643,N_27817,N_28441);
or U28644 (N_28644,N_27942,N_27948);
nor U28645 (N_28645,N_27691,N_27592);
nor U28646 (N_28646,N_27481,N_27276);
nor U28647 (N_28647,N_27096,N_27919);
or U28648 (N_28648,N_27011,N_27145);
or U28649 (N_28649,N_27374,N_27895);
nand U28650 (N_28650,N_27158,N_27818);
and U28651 (N_28651,N_27052,N_27546);
or U28652 (N_28652,N_27898,N_27806);
and U28653 (N_28653,N_28022,N_27840);
or U28654 (N_28654,N_27779,N_27057);
and U28655 (N_28655,N_27621,N_27084);
nand U28656 (N_28656,N_27162,N_27856);
or U28657 (N_28657,N_28063,N_27866);
or U28658 (N_28658,N_28118,N_27136);
nand U28659 (N_28659,N_27977,N_27770);
and U28660 (N_28660,N_27927,N_27648);
and U28661 (N_28661,N_27005,N_27487);
nand U28662 (N_28662,N_27792,N_28495);
nand U28663 (N_28663,N_27415,N_27047);
xor U28664 (N_28664,N_27171,N_28462);
xnor U28665 (N_28665,N_27492,N_27045);
and U28666 (N_28666,N_28193,N_28447);
or U28667 (N_28667,N_28273,N_27404);
nand U28668 (N_28668,N_27190,N_27666);
xnor U28669 (N_28669,N_27201,N_28306);
and U28670 (N_28670,N_28199,N_27312);
and U28671 (N_28671,N_27280,N_27460);
and U28672 (N_28672,N_27821,N_28473);
nand U28673 (N_28673,N_27412,N_27308);
and U28674 (N_28674,N_27414,N_27640);
xor U28675 (N_28675,N_27645,N_27716);
xor U28676 (N_28676,N_28150,N_27532);
xnor U28677 (N_28677,N_27922,N_28285);
nand U28678 (N_28678,N_27839,N_28294);
and U28679 (N_28679,N_27193,N_28081);
and U28680 (N_28680,N_28310,N_27316);
nor U28681 (N_28681,N_27356,N_27474);
and U28682 (N_28682,N_27445,N_27023);
and U28683 (N_28683,N_28137,N_27302);
or U28684 (N_28684,N_28217,N_27420);
or U28685 (N_28685,N_28377,N_27516);
and U28686 (N_28686,N_28291,N_27408);
or U28687 (N_28687,N_27803,N_27849);
or U28688 (N_28688,N_28260,N_27831);
nand U28689 (N_28689,N_27224,N_27638);
xnor U28690 (N_28690,N_27508,N_28195);
xnor U28691 (N_28691,N_27046,N_27417);
or U28692 (N_28692,N_27573,N_28254);
xor U28693 (N_28693,N_27173,N_28003);
nand U28694 (N_28694,N_27187,N_28091);
or U28695 (N_28695,N_27204,N_28301);
and U28696 (N_28696,N_27862,N_27222);
xor U28697 (N_28697,N_28482,N_27711);
and U28698 (N_28698,N_28052,N_27920);
or U28699 (N_28699,N_28328,N_27320);
and U28700 (N_28700,N_27957,N_27366);
and U28701 (N_28701,N_28287,N_27558);
xor U28702 (N_28702,N_27826,N_27850);
nand U28703 (N_28703,N_28204,N_27447);
and U28704 (N_28704,N_27134,N_28464);
nand U28705 (N_28705,N_27885,N_28125);
or U28706 (N_28706,N_28481,N_27115);
xnor U28707 (N_28707,N_27733,N_27399);
or U28708 (N_28708,N_27737,N_27227);
xnor U28709 (N_28709,N_28149,N_27954);
and U28710 (N_28710,N_27470,N_28066);
xor U28711 (N_28711,N_27593,N_28360);
nand U28712 (N_28712,N_27540,N_27673);
or U28713 (N_28713,N_27787,N_27678);
nor U28714 (N_28714,N_28007,N_28383);
and U28715 (N_28715,N_27736,N_27195);
nor U28716 (N_28716,N_28410,N_27342);
xor U28717 (N_28717,N_27595,N_27521);
and U28718 (N_28718,N_27409,N_27965);
nand U28719 (N_28719,N_27034,N_27994);
nand U28720 (N_28720,N_27556,N_28074);
xnor U28721 (N_28721,N_27132,N_27025);
nor U28722 (N_28722,N_28004,N_27467);
xor U28723 (N_28723,N_28181,N_27443);
xnor U28724 (N_28724,N_27567,N_27869);
or U28725 (N_28725,N_27620,N_28114);
xnor U28726 (N_28726,N_27498,N_28327);
xor U28727 (N_28727,N_28309,N_28225);
or U28728 (N_28728,N_27225,N_27500);
and U28729 (N_28729,N_27459,N_27129);
and U28730 (N_28730,N_27313,N_27798);
or U28731 (N_28731,N_27228,N_27548);
nand U28732 (N_28732,N_27479,N_28061);
nand U28733 (N_28733,N_27882,N_28034);
or U28734 (N_28734,N_27864,N_28409);
and U28735 (N_28735,N_28280,N_27923);
or U28736 (N_28736,N_28396,N_28086);
nor U28737 (N_28737,N_28185,N_27847);
xnor U28738 (N_28738,N_27533,N_27756);
xor U28739 (N_28739,N_28268,N_28304);
xor U28740 (N_28740,N_28093,N_27825);
and U28741 (N_28741,N_27208,N_28079);
or U28742 (N_28742,N_27873,N_28370);
nor U28743 (N_28743,N_27258,N_27475);
nand U28744 (N_28744,N_27658,N_27346);
and U28745 (N_28745,N_27231,N_27448);
or U28746 (N_28746,N_28071,N_28411);
nand U28747 (N_28747,N_27150,N_28250);
xnor U28748 (N_28748,N_27199,N_27631);
and U28749 (N_28749,N_27206,N_27872);
or U28750 (N_28750,N_27217,N_27809);
nor U28751 (N_28751,N_28047,N_27560);
nand U28752 (N_28752,N_27932,N_28230);
nand U28753 (N_28753,N_28049,N_27341);
and U28754 (N_28754,N_27740,N_28252);
nor U28755 (N_28755,N_27566,N_28015);
xnor U28756 (N_28756,N_27654,N_28116);
or U28757 (N_28757,N_27058,N_27000);
or U28758 (N_28758,N_27072,N_27668);
or U28759 (N_28759,N_27874,N_27067);
or U28760 (N_28760,N_28453,N_27944);
xnor U28761 (N_28761,N_27641,N_27423);
nand U28762 (N_28762,N_27371,N_28303);
xnor U28763 (N_28763,N_27332,N_27381);
xnor U28764 (N_28764,N_27086,N_27361);
nand U28765 (N_28765,N_27844,N_27701);
nand U28766 (N_28766,N_27398,N_27368);
xor U28767 (N_28767,N_27033,N_27738);
nand U28768 (N_28768,N_28058,N_28240);
nor U28769 (N_28769,N_28365,N_27114);
xor U28770 (N_28770,N_28351,N_27270);
and U28771 (N_28771,N_27147,N_28030);
xnor U28772 (N_28772,N_27955,N_27232);
xnor U28773 (N_28773,N_27877,N_27975);
nand U28774 (N_28774,N_27172,N_27577);
nand U28775 (N_28775,N_28110,N_28391);
nor U28776 (N_28776,N_27160,N_28178);
nand U28777 (N_28777,N_27249,N_27700);
nor U28778 (N_28778,N_27230,N_28324);
xnor U28779 (N_28779,N_27082,N_27269);
nand U28780 (N_28780,N_27031,N_27358);
or U28781 (N_28781,N_27251,N_27805);
nor U28782 (N_28782,N_27660,N_27466);
nor U28783 (N_28783,N_27478,N_27146);
nor U28784 (N_28784,N_28336,N_27265);
or U28785 (N_28785,N_28100,N_27424);
and U28786 (N_28786,N_27290,N_28314);
xnor U28787 (N_28787,N_27116,N_28205);
or U28788 (N_28788,N_28329,N_27557);
and U28789 (N_28789,N_27009,N_27672);
nor U28790 (N_28790,N_27551,N_27093);
xnor U28791 (N_28791,N_28223,N_27016);
and U28792 (N_28792,N_28033,N_27718);
nor U28793 (N_28793,N_27791,N_27715);
or U28794 (N_28794,N_28318,N_28194);
and U28795 (N_28795,N_28109,N_27588);
and U28796 (N_28796,N_27092,N_27581);
and U28797 (N_28797,N_28384,N_27212);
and U28798 (N_28798,N_28375,N_28054);
nor U28799 (N_28799,N_27615,N_28302);
or U28800 (N_28800,N_27783,N_27326);
or U28801 (N_28801,N_27761,N_28466);
and U28802 (N_28802,N_27690,N_27801);
nor U28803 (N_28803,N_28160,N_27156);
xnor U28804 (N_28804,N_27771,N_28474);
nor U28805 (N_28805,N_27311,N_27221);
nor U28806 (N_28806,N_28339,N_28415);
nand U28807 (N_28807,N_27396,N_27303);
nor U28808 (N_28808,N_27185,N_27766);
and U28809 (N_28809,N_28168,N_27897);
nor U28810 (N_28810,N_28094,N_28320);
xnor U28811 (N_28811,N_28068,N_28130);
nand U28812 (N_28812,N_27392,N_28143);
xnor U28813 (N_28813,N_27197,N_27743);
and U28814 (N_28814,N_27607,N_27751);
nor U28815 (N_28815,N_28098,N_28266);
xnor U28816 (N_28816,N_28147,N_27177);
or U28817 (N_28817,N_27995,N_27350);
nand U28818 (N_28818,N_27305,N_28427);
xor U28819 (N_28819,N_28317,N_27739);
or U28820 (N_28820,N_27951,N_27572);
nor U28821 (N_28821,N_27099,N_27453);
nand U28822 (N_28822,N_27627,N_28019);
or U28823 (N_28823,N_27623,N_28338);
and U28824 (N_28824,N_28060,N_28498);
and U28825 (N_28825,N_28001,N_27681);
or U28826 (N_28826,N_27142,N_27349);
or U28827 (N_28827,N_28359,N_28134);
nand U28828 (N_28828,N_27934,N_28454);
and U28829 (N_28829,N_27331,N_28475);
nor U28830 (N_28830,N_27257,N_28286);
nand U28831 (N_28831,N_27218,N_28269);
nand U28832 (N_28832,N_28343,N_28145);
xnor U28833 (N_28833,N_27833,N_27988);
nor U28834 (N_28834,N_28245,N_28346);
nor U28835 (N_28835,N_27006,N_28206);
xor U28836 (N_28836,N_27547,N_28029);
and U28837 (N_28837,N_28191,N_27561);
xor U28838 (N_28838,N_27087,N_27945);
nand U28839 (N_28839,N_28249,N_28092);
and U28840 (N_28840,N_27815,N_27059);
nor U28841 (N_28841,N_27176,N_27348);
nand U28842 (N_28842,N_27579,N_27296);
nor U28843 (N_28843,N_27022,N_27745);
and U28844 (N_28844,N_27830,N_27570);
nand U28845 (N_28845,N_28376,N_27278);
nor U28846 (N_28846,N_27857,N_27967);
xnor U28847 (N_28847,N_27871,N_28262);
or U28848 (N_28848,N_28215,N_28449);
nand U28849 (N_28849,N_27855,N_27063);
or U28850 (N_28850,N_28128,N_27793);
nand U28851 (N_28851,N_27235,N_27239);
nor U28852 (N_28852,N_27454,N_27301);
or U28853 (N_28853,N_28242,N_27894);
and U28854 (N_28854,N_27476,N_27698);
or U28855 (N_28855,N_28238,N_28369);
nor U28856 (N_28856,N_27603,N_27552);
or U28857 (N_28857,N_27319,N_27194);
xnor U28858 (N_28858,N_28307,N_27987);
xor U28859 (N_28859,N_27165,N_27246);
xnor U28860 (N_28860,N_27868,N_27741);
xnor U28861 (N_28861,N_28101,N_28451);
and U28862 (N_28862,N_28326,N_27685);
nand U28863 (N_28863,N_27655,N_27702);
xnor U28864 (N_28864,N_28386,N_27657);
nand U28865 (N_28865,N_27062,N_27354);
xnor U28866 (N_28866,N_28151,N_27904);
nor U28867 (N_28867,N_27440,N_27433);
nor U28868 (N_28868,N_27073,N_27823);
xor U28869 (N_28869,N_28175,N_28348);
or U28870 (N_28870,N_28353,N_27647);
and U28871 (N_28871,N_27463,N_27909);
and U28872 (N_28872,N_28148,N_28340);
or U28873 (N_28873,N_27154,N_27018);
xor U28874 (N_28874,N_28244,N_27723);
or U28875 (N_28875,N_28082,N_27714);
or U28876 (N_28876,N_28439,N_27910);
nor U28877 (N_28877,N_27406,N_28426);
xor U28878 (N_28878,N_28219,N_27531);
and U28879 (N_28879,N_27971,N_27140);
nand U28880 (N_28880,N_27175,N_28202);
or U28881 (N_28881,N_27891,N_27979);
nor U28882 (N_28882,N_28489,N_28042);
nor U28883 (N_28883,N_28167,N_28024);
xor U28884 (N_28884,N_28196,N_27362);
nand U28885 (N_28885,N_28434,N_27469);
xor U28886 (N_28886,N_28113,N_27837);
xor U28887 (N_28887,N_28246,N_27530);
xor U28888 (N_28888,N_28418,N_27617);
or U28889 (N_28889,N_27555,N_28440);
or U28890 (N_28890,N_27180,N_27152);
and U28891 (N_28891,N_28494,N_27071);
nor U28892 (N_28892,N_27291,N_27732);
nand U28893 (N_28893,N_27523,N_27395);
nand U28894 (N_28894,N_28382,N_28288);
nand U28895 (N_28895,N_27632,N_27277);
xnor U28896 (N_28896,N_27369,N_27437);
and U28897 (N_28897,N_27907,N_27842);
nand U28898 (N_28898,N_28161,N_27446);
nand U28899 (N_28899,N_27936,N_28124);
xnor U28900 (N_28900,N_28153,N_27200);
or U28901 (N_28901,N_28344,N_27435);
nand U28902 (N_28902,N_28321,N_27149);
nand U28903 (N_28903,N_28070,N_27628);
and U28904 (N_28904,N_27618,N_27964);
nor U28905 (N_28905,N_28097,N_27653);
xor U28906 (N_28906,N_28065,N_27338);
nor U28907 (N_28907,N_27286,N_28284);
or U28908 (N_28908,N_27400,N_28008);
and U28909 (N_28909,N_27219,N_27495);
nand U28910 (N_28910,N_27032,N_27652);
xnor U28911 (N_28911,N_27181,N_28289);
or U28912 (N_28912,N_28334,N_28163);
and U28913 (N_28913,N_27933,N_28186);
nor U28914 (N_28914,N_27989,N_27750);
xnor U28915 (N_28915,N_27088,N_27166);
nand U28916 (N_28916,N_27490,N_28190);
nand U28917 (N_28917,N_28470,N_28214);
nor U28918 (N_28918,N_27903,N_27157);
xor U28919 (N_28919,N_28132,N_28264);
nor U28920 (N_28920,N_28446,N_28028);
xnor U28921 (N_28921,N_27108,N_28156);
and U28922 (N_28922,N_28319,N_28141);
and U28923 (N_28923,N_27444,N_27428);
nor U28924 (N_28924,N_27205,N_27824);
or U28925 (N_28925,N_28278,N_27697);
nor U28926 (N_28926,N_28499,N_27507);
xnor U28927 (N_28927,N_27630,N_27816);
and U28928 (N_28928,N_28477,N_28431);
nand U28929 (N_28929,N_27359,N_27210);
nand U28930 (N_28930,N_28000,N_28350);
nand U28931 (N_28931,N_28460,N_27182);
nor U28932 (N_28932,N_27283,N_28048);
nor U28933 (N_28933,N_27125,N_27966);
xnor U28934 (N_28934,N_27800,N_28356);
nand U28935 (N_28935,N_27887,N_27259);
xor U28936 (N_28936,N_27726,N_28231);
and U28937 (N_28937,N_27497,N_28333);
xnor U28938 (N_28938,N_28227,N_27886);
xnor U28939 (N_28939,N_27238,N_27786);
nand U28940 (N_28940,N_27075,N_27748);
or U28941 (N_28941,N_28120,N_28313);
xor U28942 (N_28942,N_27519,N_27024);
xor U28943 (N_28943,N_28171,N_27095);
and U28944 (N_28944,N_28368,N_28174);
xnor U28945 (N_28945,N_27789,N_27893);
xnor U28946 (N_28946,N_27449,N_28005);
and U28947 (N_28947,N_27345,N_27214);
nor U28948 (N_28948,N_27814,N_27611);
nor U28949 (N_28949,N_27596,N_28162);
xnor U28950 (N_28950,N_27642,N_27905);
nor U28951 (N_28951,N_28095,N_27499);
and U28952 (N_28952,N_27545,N_27636);
and U28953 (N_28953,N_27416,N_28490);
and U28954 (N_28954,N_28452,N_27626);
and U28955 (N_28955,N_27976,N_27405);
xor U28956 (N_28956,N_27562,N_27130);
xor U28957 (N_28957,N_27411,N_28349);
or U28958 (N_28958,N_27758,N_27725);
nand U28959 (N_28959,N_28295,N_28059);
nor U28960 (N_28960,N_27692,N_27663);
or U28961 (N_28961,N_28013,N_28139);
xnor U28962 (N_28962,N_27537,N_27952);
or U28963 (N_28963,N_27041,N_27275);
or U28964 (N_28964,N_27949,N_27339);
or U28965 (N_28965,N_28404,N_28180);
and U28966 (N_28966,N_27139,N_28201);
nand U28967 (N_28967,N_28421,N_27527);
and U28968 (N_28968,N_28337,N_27665);
and U28969 (N_28969,N_27355,N_27991);
or U28970 (N_28970,N_28456,N_28292);
or U28971 (N_28971,N_27941,N_27675);
nand U28972 (N_28972,N_27109,N_27509);
nor U28973 (N_28973,N_28213,N_28140);
and U28974 (N_28974,N_27674,N_28450);
nand U28975 (N_28975,N_28357,N_27811);
or U28976 (N_28976,N_27535,N_27616);
or U28977 (N_28977,N_28424,N_28398);
nor U28978 (N_28978,N_27248,N_27167);
or U28979 (N_28979,N_27288,N_27314);
or U28980 (N_28980,N_28129,N_28107);
xnor U28981 (N_28981,N_28222,N_27323);
nor U28982 (N_28982,N_27306,N_27870);
nand U28983 (N_28983,N_28016,N_28155);
and U28984 (N_28984,N_27256,N_27216);
and U28985 (N_28985,N_28067,N_27106);
or U28986 (N_28986,N_27625,N_27191);
xor U28987 (N_28987,N_27026,N_28311);
and U28988 (N_28988,N_28277,N_27465);
nor U28989 (N_28989,N_27568,N_28364);
xnor U28990 (N_28990,N_28347,N_27321);
nand U28991 (N_28991,N_27968,N_27425);
or U28992 (N_28992,N_27676,N_27843);
nand U28993 (N_28993,N_27237,N_27101);
nor U28994 (N_28994,N_28111,N_27822);
or U28995 (N_28995,N_27336,N_27282);
and U28996 (N_28996,N_27300,N_28459);
xor U28997 (N_28997,N_27526,N_27524);
nand U28998 (N_28998,N_28144,N_28390);
xnor U28999 (N_28999,N_27511,N_28274);
nor U29000 (N_29000,N_27014,N_27091);
and U29001 (N_29001,N_28121,N_28038);
or U29002 (N_29002,N_27126,N_27565);
and U29003 (N_29003,N_27294,N_28243);
nand U29004 (N_29004,N_27940,N_27284);
nand U29005 (N_29005,N_28072,N_28112);
or U29006 (N_29006,N_27327,N_27462);
or U29007 (N_29007,N_28381,N_27461);
and U29008 (N_29008,N_27911,N_28138);
or U29009 (N_29009,N_27646,N_27728);
nor U29010 (N_29010,N_28430,N_27643);
nand U29011 (N_29011,N_27007,N_27921);
and U29012 (N_29012,N_27170,N_27473);
xnor U29013 (N_29013,N_27029,N_28146);
xnor U29014 (N_29014,N_27044,N_27489);
nand U29015 (N_29015,N_27442,N_27250);
and U29016 (N_29016,N_27799,N_27762);
or U29017 (N_29017,N_27089,N_27080);
or U29018 (N_29018,N_27377,N_27510);
xor U29019 (N_29019,N_27529,N_27661);
nand U29020 (N_29020,N_27322,N_28472);
nand U29021 (N_29021,N_27289,N_28037);
or U29022 (N_29022,N_28189,N_27525);
and U29023 (N_29023,N_28448,N_28413);
or U29024 (N_29024,N_27351,N_27781);
xor U29025 (N_29025,N_27883,N_27037);
xor U29026 (N_29026,N_27571,N_28420);
and U29027 (N_29027,N_27019,N_28366);
or U29028 (N_29028,N_27742,N_27912);
nand U29029 (N_29029,N_28491,N_27590);
and U29030 (N_29030,N_27118,N_28271);
nor U29031 (N_29031,N_27253,N_28363);
xnor U29032 (N_29032,N_28115,N_28308);
nand U29033 (N_29033,N_28255,N_27892);
nor U29034 (N_29034,N_27429,N_28429);
xnor U29035 (N_29035,N_28312,N_27102);
nor U29036 (N_29036,N_28200,N_27496);
nor U29037 (N_29037,N_27441,N_27491);
nand U29038 (N_29038,N_27998,N_27956);
or U29039 (N_29039,N_27835,N_27984);
and U29040 (N_29040,N_28085,N_27852);
nand U29041 (N_29041,N_27730,N_27744);
and U29042 (N_29042,N_27916,N_27778);
or U29043 (N_29043,N_27383,N_27598);
and U29044 (N_29044,N_27472,N_28444);
nand U29045 (N_29045,N_28247,N_27587);
xnor U29046 (N_29046,N_27586,N_28275);
nor U29047 (N_29047,N_27760,N_27972);
nor U29048 (N_29048,N_27343,N_27981);
xnor U29049 (N_29049,N_27503,N_27078);
nor U29050 (N_29050,N_27310,N_27597);
nor U29051 (N_29051,N_27357,N_27328);
and U29052 (N_29052,N_27309,N_27117);
nor U29053 (N_29053,N_28096,N_27353);
and U29054 (N_29054,N_28253,N_27712);
xor U29055 (N_29055,N_27553,N_28455);
or U29056 (N_29056,N_28083,N_28089);
and U29057 (N_29057,N_27161,N_27127);
or U29058 (N_29058,N_27457,N_28017);
nor U29059 (N_29059,N_27164,N_27827);
nand U29060 (N_29060,N_27997,N_27749);
nand U29061 (N_29061,N_28023,N_28104);
or U29062 (N_29062,N_27030,N_27401);
or U29063 (N_29063,N_28487,N_28212);
and U29064 (N_29064,N_27717,N_27141);
nor U29065 (N_29065,N_28457,N_28232);
nor U29066 (N_29066,N_27153,N_28371);
nor U29067 (N_29067,N_27329,N_27370);
nor U29068 (N_29068,N_27012,N_27699);
and U29069 (N_29069,N_27159,N_27656);
nand U29070 (N_29070,N_28296,N_27709);
xor U29071 (N_29071,N_28478,N_27365);
xnor U29072 (N_29072,N_28010,N_27110);
or U29073 (N_29073,N_27785,N_28031);
or U29074 (N_29074,N_27064,N_28203);
xor U29075 (N_29075,N_28290,N_27244);
nand U29076 (N_29076,N_27168,N_27722);
or U29077 (N_29077,N_27077,N_27963);
xnor U29078 (N_29078,N_27422,N_28218);
or U29079 (N_29079,N_28075,N_28105);
xnor U29080 (N_29080,N_27419,N_28176);
or U29081 (N_29081,N_28276,N_28265);
nor U29082 (N_29082,N_27060,N_27790);
xor U29083 (N_29083,N_28385,N_27810);
nor U29084 (N_29084,N_27594,N_28394);
and U29085 (N_29085,N_27421,N_27671);
and U29086 (N_29086,N_28435,N_28233);
nand U29087 (N_29087,N_28298,N_27439);
and U29088 (N_29088,N_28044,N_27884);
xnor U29089 (N_29089,N_28043,N_27344);
xnor U29090 (N_29090,N_27601,N_27982);
nand U29091 (N_29091,N_27713,N_27198);
and U29092 (N_29092,N_28401,N_27050);
xor U29093 (N_29093,N_28331,N_28036);
nor U29094 (N_29094,N_27506,N_28207);
and U29095 (N_29095,N_27943,N_28021);
xor U29096 (N_29096,N_27576,N_28493);
nor U29097 (N_29097,N_27689,N_27389);
xor U29098 (N_29098,N_27928,N_28407);
xor U29099 (N_29099,N_28379,N_28406);
nand U29100 (N_29100,N_27255,N_27427);
or U29101 (N_29101,N_28220,N_28046);
or U29102 (N_29102,N_28126,N_28183);
and U29103 (N_29103,N_27929,N_27808);
or U29104 (N_29104,N_28051,N_28234);
nand U29105 (N_29105,N_27931,N_27664);
and U29106 (N_29106,N_27407,N_27878);
xor U29107 (N_29107,N_27735,N_27021);
nand U29108 (N_29108,N_27828,N_27268);
nor U29109 (N_29109,N_27776,N_27455);
xnor U29110 (N_29110,N_27155,N_27832);
xor U29111 (N_29111,N_27049,N_27875);
nor U29112 (N_29112,N_28400,N_27765);
xnor U29113 (N_29113,N_27950,N_27438);
xnor U29114 (N_29114,N_28158,N_27522);
xor U29115 (N_29115,N_28479,N_27318);
nand U29116 (N_29116,N_28461,N_27340);
and U29117 (N_29117,N_27774,N_27719);
nor U29118 (N_29118,N_27612,N_27634);
nand U29119 (N_29119,N_28258,N_27708);
and U29120 (N_29120,N_27992,N_27662);
and U29121 (N_29121,N_27550,N_28197);
or U29122 (N_29122,N_27860,N_28372);
xor U29123 (N_29123,N_28257,N_28025);
and U29124 (N_29124,N_28488,N_27372);
and U29125 (N_29125,N_27196,N_27784);
nor U29126 (N_29126,N_27015,N_28408);
nor U29127 (N_29127,N_27682,N_27890);
xnor U29128 (N_29128,N_27720,N_27403);
and U29129 (N_29129,N_27451,N_27695);
nor U29130 (N_29130,N_28484,N_27609);
or U29131 (N_29131,N_27243,N_27452);
or U29132 (N_29132,N_27262,N_28055);
nand U29133 (N_29133,N_27324,N_27584);
nor U29134 (N_29134,N_27051,N_27938);
or U29135 (N_29135,N_28374,N_27065);
or U29136 (N_29136,N_28076,N_27378);
nor U29137 (N_29137,N_27937,N_27924);
or U29138 (N_29138,N_28169,N_27431);
nand U29139 (N_29139,N_27999,N_27962);
and U29140 (N_29140,N_27679,N_28177);
nand U29141 (N_29141,N_28480,N_27013);
nand U29142 (N_29142,N_27272,N_27390);
and U29143 (N_29143,N_27148,N_28216);
nor U29144 (N_29144,N_27042,N_27053);
nand U29145 (N_29145,N_27347,N_28002);
or U29146 (N_29146,N_28045,N_27947);
nor U29147 (N_29147,N_28469,N_28345);
nor U29148 (N_29148,N_27583,N_27820);
or U29149 (N_29149,N_27233,N_27207);
xnor U29150 (N_29150,N_28272,N_28084);
or U29151 (N_29151,N_28188,N_27410);
nor U29152 (N_29152,N_28170,N_27202);
nor U29153 (N_29153,N_27769,N_28127);
nand U29154 (N_29154,N_27838,N_28142);
nor U29155 (N_29155,N_28099,N_27418);
or U29156 (N_29156,N_27330,N_27958);
nand U29157 (N_29157,N_27070,N_27520);
nand U29158 (N_29158,N_27959,N_28467);
and U29159 (N_29159,N_27292,N_28164);
nand U29160 (N_29160,N_27795,N_27504);
nand U29161 (N_29161,N_28367,N_27004);
nor U29162 (N_29162,N_27973,N_27935);
xnor U29163 (N_29163,N_27281,N_27727);
or U29164 (N_29164,N_28267,N_28062);
nor U29165 (N_29165,N_27380,N_27179);
nor U29166 (N_29166,N_27580,N_27599);
and U29167 (N_29167,N_27493,N_28355);
or U29168 (N_29168,N_28053,N_27450);
and U29169 (N_29169,N_27223,N_27384);
and U29170 (N_29170,N_27085,N_28342);
xor U29171 (N_29171,N_27391,N_27183);
nand U29172 (N_29172,N_27394,N_27298);
nor U29173 (N_29173,N_27721,N_28224);
nand U29174 (N_29174,N_27137,N_28237);
nand U29175 (N_29175,N_28380,N_28373);
xor U29176 (N_29176,N_27534,N_28173);
nor U29177 (N_29177,N_28211,N_27915);
xnor U29178 (N_29178,N_27027,N_27686);
nor U29179 (N_29179,N_27667,N_28057);
and U29180 (N_29180,N_27528,N_27763);
or U29181 (N_29181,N_27061,N_27926);
nor U29182 (N_29182,N_27261,N_28433);
nand U29183 (N_29183,N_28468,N_27456);
and U29184 (N_29184,N_27098,N_27752);
or U29185 (N_29185,N_27036,N_27542);
nor U29186 (N_29186,N_28012,N_28041);
and U29187 (N_29187,N_27054,N_28483);
or U29188 (N_29188,N_28403,N_28026);
nand U29189 (N_29189,N_27432,N_27788);
or U29190 (N_29190,N_28496,N_27234);
and U29191 (N_29191,N_27008,N_27090);
or U29192 (N_29192,N_28405,N_27169);
and U29193 (N_29193,N_27267,N_28463);
or U29194 (N_29194,N_27960,N_27729);
or U29195 (N_29195,N_27264,N_27677);
or U29196 (N_29196,N_27602,N_28485);
nor U29197 (N_29197,N_27613,N_27694);
or U29198 (N_29198,N_28248,N_28412);
nand U29199 (N_29199,N_27103,N_27834);
or U29200 (N_29200,N_27605,N_27335);
or U29201 (N_29201,N_27468,N_28119);
nand U29202 (N_29202,N_27334,N_28018);
xnor U29203 (N_29203,N_27188,N_27484);
nand U29204 (N_29204,N_27917,N_27260);
xnor U29205 (N_29205,N_27578,N_27990);
nand U29206 (N_29206,N_27753,N_28103);
nor U29207 (N_29207,N_28423,N_28297);
and U29208 (N_29208,N_27650,N_27961);
nor U29209 (N_29209,N_27619,N_27144);
nand U29210 (N_29210,N_27986,N_28011);
and U29211 (N_29211,N_27853,N_27028);
nor U29212 (N_29212,N_27757,N_27775);
nand U29213 (N_29213,N_27707,N_27901);
xor U29214 (N_29214,N_27120,N_27930);
xnor U29215 (N_29215,N_27591,N_27501);
xor U29216 (N_29216,N_27483,N_27010);
nand U29217 (N_29217,N_27119,N_28209);
nand U29218 (N_29218,N_27174,N_27100);
or U29219 (N_29219,N_27670,N_27485);
nor U29220 (N_29220,N_27178,N_27782);
and U29221 (N_29221,N_27017,N_27382);
nand U29222 (N_29222,N_27043,N_27367);
xor U29223 (N_29223,N_27683,N_28087);
xnor U29224 (N_29224,N_27471,N_27240);
nor U29225 (N_29225,N_27263,N_28187);
nor U29226 (N_29226,N_27777,N_28486);
or U29227 (N_29227,N_27606,N_27364);
and U29228 (N_29228,N_27138,N_28069);
nand U29229 (N_29229,N_28228,N_27794);
or U29230 (N_29230,N_28378,N_27985);
and U29231 (N_29231,N_28358,N_27980);
xor U29232 (N_29232,N_27974,N_27865);
xnor U29233 (N_29233,N_27107,N_28281);
xnor U29234 (N_29234,N_28419,N_28040);
or U29235 (N_29235,N_27807,N_27754);
nor U29236 (N_29236,N_27505,N_27637);
xor U29237 (N_29237,N_27069,N_27513);
or U29238 (N_29238,N_27635,N_27539);
nor U29239 (N_29239,N_28172,N_27841);
xnor U29240 (N_29240,N_28039,N_28080);
nor U29241 (N_29241,N_28157,N_27131);
nor U29242 (N_29242,N_27549,N_27488);
and U29243 (N_29243,N_27299,N_27203);
and U29244 (N_29244,N_27813,N_27836);
and U29245 (N_29245,N_27097,N_27604);
nand U29246 (N_29246,N_28229,N_27385);
nor U29247 (N_29247,N_27554,N_27900);
nor U29248 (N_29248,N_28020,N_27764);
and U29249 (N_29249,N_27215,N_28165);
nand U29250 (N_29250,N_27470,N_27735);
or U29251 (N_29251,N_28305,N_28370);
nand U29252 (N_29252,N_27805,N_28424);
nor U29253 (N_29253,N_27389,N_28129);
and U29254 (N_29254,N_28312,N_27377);
or U29255 (N_29255,N_28483,N_28099);
and U29256 (N_29256,N_27428,N_28075);
nor U29257 (N_29257,N_28295,N_27523);
and U29258 (N_29258,N_27618,N_27274);
nor U29259 (N_29259,N_27033,N_27712);
and U29260 (N_29260,N_27768,N_27232);
or U29261 (N_29261,N_28497,N_27137);
nand U29262 (N_29262,N_28145,N_27470);
nand U29263 (N_29263,N_27334,N_27942);
or U29264 (N_29264,N_27070,N_27885);
nand U29265 (N_29265,N_28406,N_27619);
nor U29266 (N_29266,N_27583,N_27945);
nor U29267 (N_29267,N_28442,N_27780);
xnor U29268 (N_29268,N_27125,N_27916);
or U29269 (N_29269,N_27006,N_27411);
nand U29270 (N_29270,N_27129,N_28025);
and U29271 (N_29271,N_28437,N_27548);
nand U29272 (N_29272,N_27827,N_27136);
nor U29273 (N_29273,N_28467,N_27829);
or U29274 (N_29274,N_27221,N_27600);
nand U29275 (N_29275,N_27607,N_27488);
and U29276 (N_29276,N_27830,N_28044);
nor U29277 (N_29277,N_27066,N_28199);
and U29278 (N_29278,N_27502,N_27247);
nor U29279 (N_29279,N_28455,N_27581);
and U29280 (N_29280,N_27191,N_27145);
nand U29281 (N_29281,N_28484,N_28266);
and U29282 (N_29282,N_28288,N_27652);
or U29283 (N_29283,N_27395,N_28356);
nor U29284 (N_29284,N_27164,N_27933);
xor U29285 (N_29285,N_27198,N_27467);
nor U29286 (N_29286,N_27913,N_27784);
or U29287 (N_29287,N_27571,N_28369);
xor U29288 (N_29288,N_28140,N_27141);
xor U29289 (N_29289,N_27136,N_27853);
nand U29290 (N_29290,N_27336,N_28047);
nand U29291 (N_29291,N_28077,N_27923);
xor U29292 (N_29292,N_28192,N_27002);
nand U29293 (N_29293,N_28229,N_28172);
nand U29294 (N_29294,N_28012,N_28049);
xnor U29295 (N_29295,N_28090,N_28332);
or U29296 (N_29296,N_28029,N_28323);
xnor U29297 (N_29297,N_27175,N_28244);
xnor U29298 (N_29298,N_27383,N_27117);
and U29299 (N_29299,N_27407,N_27304);
or U29300 (N_29300,N_27037,N_28094);
nand U29301 (N_29301,N_27545,N_28139);
nand U29302 (N_29302,N_27354,N_27084);
nand U29303 (N_29303,N_28205,N_27541);
nand U29304 (N_29304,N_28260,N_27095);
or U29305 (N_29305,N_27727,N_28234);
nand U29306 (N_29306,N_27837,N_28111);
or U29307 (N_29307,N_27426,N_28487);
xor U29308 (N_29308,N_28448,N_28410);
nor U29309 (N_29309,N_28039,N_28373);
xnor U29310 (N_29310,N_28495,N_27366);
and U29311 (N_29311,N_27072,N_28269);
xor U29312 (N_29312,N_27235,N_27801);
nor U29313 (N_29313,N_28253,N_27144);
nor U29314 (N_29314,N_28100,N_27213);
xor U29315 (N_29315,N_27227,N_27245);
nor U29316 (N_29316,N_28327,N_27274);
nor U29317 (N_29317,N_27264,N_27843);
nor U29318 (N_29318,N_27739,N_27960);
xor U29319 (N_29319,N_27580,N_28240);
nor U29320 (N_29320,N_27192,N_28088);
xor U29321 (N_29321,N_27341,N_28207);
nand U29322 (N_29322,N_27133,N_28098);
nor U29323 (N_29323,N_27927,N_27466);
nand U29324 (N_29324,N_27820,N_27646);
nand U29325 (N_29325,N_28143,N_28159);
or U29326 (N_29326,N_27173,N_27903);
and U29327 (N_29327,N_28321,N_28119);
xor U29328 (N_29328,N_27975,N_27443);
nand U29329 (N_29329,N_27980,N_27191);
or U29330 (N_29330,N_28395,N_28189);
xnor U29331 (N_29331,N_27572,N_28233);
or U29332 (N_29332,N_28355,N_28146);
nor U29333 (N_29333,N_28496,N_28310);
nand U29334 (N_29334,N_27907,N_27299);
or U29335 (N_29335,N_27046,N_28126);
nor U29336 (N_29336,N_27796,N_28318);
xnor U29337 (N_29337,N_27075,N_28421);
nor U29338 (N_29338,N_27399,N_27028);
and U29339 (N_29339,N_27950,N_27151);
and U29340 (N_29340,N_27931,N_27775);
nand U29341 (N_29341,N_27312,N_27222);
xnor U29342 (N_29342,N_28015,N_27649);
nor U29343 (N_29343,N_28134,N_27552);
xor U29344 (N_29344,N_27369,N_27524);
and U29345 (N_29345,N_27030,N_27036);
and U29346 (N_29346,N_27814,N_27170);
nand U29347 (N_29347,N_27056,N_27032);
nor U29348 (N_29348,N_27033,N_27210);
nand U29349 (N_29349,N_27827,N_27179);
xor U29350 (N_29350,N_27225,N_27441);
xnor U29351 (N_29351,N_27594,N_27643);
or U29352 (N_29352,N_27494,N_28199);
nand U29353 (N_29353,N_27822,N_28286);
and U29354 (N_29354,N_28444,N_27909);
xnor U29355 (N_29355,N_27833,N_28302);
nor U29356 (N_29356,N_28062,N_27186);
or U29357 (N_29357,N_27934,N_27763);
and U29358 (N_29358,N_28084,N_28162);
xor U29359 (N_29359,N_28464,N_27308);
nor U29360 (N_29360,N_28477,N_27313);
or U29361 (N_29361,N_27670,N_27510);
nor U29362 (N_29362,N_27364,N_27938);
nor U29363 (N_29363,N_28098,N_27446);
or U29364 (N_29364,N_27049,N_27609);
xor U29365 (N_29365,N_27133,N_27514);
xor U29366 (N_29366,N_27948,N_27559);
nor U29367 (N_29367,N_27404,N_27580);
nor U29368 (N_29368,N_27978,N_27526);
xor U29369 (N_29369,N_28082,N_28303);
nand U29370 (N_29370,N_28249,N_27947);
or U29371 (N_29371,N_28195,N_27795);
nand U29372 (N_29372,N_27398,N_27477);
nor U29373 (N_29373,N_27243,N_28419);
nor U29374 (N_29374,N_27838,N_27493);
xor U29375 (N_29375,N_27836,N_27757);
and U29376 (N_29376,N_27101,N_27370);
xor U29377 (N_29377,N_28009,N_27698);
nand U29378 (N_29378,N_27478,N_27012);
and U29379 (N_29379,N_28356,N_27577);
and U29380 (N_29380,N_28404,N_27611);
or U29381 (N_29381,N_27812,N_27865);
nand U29382 (N_29382,N_27198,N_27954);
nand U29383 (N_29383,N_27851,N_28098);
nand U29384 (N_29384,N_27941,N_27495);
nor U29385 (N_29385,N_27046,N_28498);
nor U29386 (N_29386,N_27523,N_27912);
nor U29387 (N_29387,N_27531,N_27684);
nand U29388 (N_29388,N_27727,N_27651);
or U29389 (N_29389,N_27766,N_27166);
xnor U29390 (N_29390,N_27963,N_27629);
nor U29391 (N_29391,N_27566,N_27960);
and U29392 (N_29392,N_28366,N_28056);
xnor U29393 (N_29393,N_27295,N_28322);
nand U29394 (N_29394,N_28411,N_28169);
and U29395 (N_29395,N_27535,N_28437);
nor U29396 (N_29396,N_27140,N_27987);
or U29397 (N_29397,N_27496,N_27535);
nand U29398 (N_29398,N_28457,N_28174);
xnor U29399 (N_29399,N_27013,N_27263);
or U29400 (N_29400,N_27003,N_27090);
nand U29401 (N_29401,N_27134,N_28411);
nand U29402 (N_29402,N_27095,N_27969);
nand U29403 (N_29403,N_28066,N_28405);
nand U29404 (N_29404,N_27755,N_28027);
nand U29405 (N_29405,N_27940,N_28204);
nand U29406 (N_29406,N_27635,N_27914);
xnor U29407 (N_29407,N_27488,N_28347);
and U29408 (N_29408,N_27541,N_28485);
and U29409 (N_29409,N_27802,N_27793);
nand U29410 (N_29410,N_27110,N_27865);
and U29411 (N_29411,N_27452,N_28145);
or U29412 (N_29412,N_27242,N_28334);
and U29413 (N_29413,N_27903,N_27961);
and U29414 (N_29414,N_27185,N_27686);
nor U29415 (N_29415,N_28162,N_27618);
xor U29416 (N_29416,N_27307,N_28138);
xnor U29417 (N_29417,N_27217,N_27764);
nand U29418 (N_29418,N_28494,N_28348);
or U29419 (N_29419,N_27705,N_27667);
and U29420 (N_29420,N_27316,N_27473);
or U29421 (N_29421,N_28278,N_28142);
nand U29422 (N_29422,N_28290,N_28394);
and U29423 (N_29423,N_28048,N_28072);
nor U29424 (N_29424,N_28181,N_27993);
xor U29425 (N_29425,N_28408,N_27424);
xnor U29426 (N_29426,N_28466,N_27465);
and U29427 (N_29427,N_27441,N_28437);
xor U29428 (N_29428,N_27401,N_27051);
or U29429 (N_29429,N_27661,N_27867);
or U29430 (N_29430,N_28200,N_27804);
nor U29431 (N_29431,N_28285,N_28034);
xor U29432 (N_29432,N_27458,N_27259);
xor U29433 (N_29433,N_28183,N_28286);
and U29434 (N_29434,N_28137,N_27206);
nor U29435 (N_29435,N_28017,N_27750);
nand U29436 (N_29436,N_27499,N_27813);
or U29437 (N_29437,N_27495,N_28309);
nand U29438 (N_29438,N_27748,N_27699);
and U29439 (N_29439,N_27221,N_28488);
or U29440 (N_29440,N_27517,N_28415);
and U29441 (N_29441,N_27298,N_27511);
xnor U29442 (N_29442,N_28445,N_27483);
xor U29443 (N_29443,N_27014,N_27222);
or U29444 (N_29444,N_28341,N_28074);
nor U29445 (N_29445,N_27444,N_27064);
and U29446 (N_29446,N_27097,N_27802);
nor U29447 (N_29447,N_27829,N_28341);
xor U29448 (N_29448,N_27570,N_27657);
xnor U29449 (N_29449,N_28352,N_28450);
nand U29450 (N_29450,N_27626,N_27776);
nand U29451 (N_29451,N_27732,N_27207);
and U29452 (N_29452,N_28490,N_28195);
xor U29453 (N_29453,N_27539,N_28255);
nand U29454 (N_29454,N_27683,N_27365);
xor U29455 (N_29455,N_27311,N_27006);
nor U29456 (N_29456,N_27235,N_27052);
nand U29457 (N_29457,N_27443,N_28354);
or U29458 (N_29458,N_28096,N_27741);
and U29459 (N_29459,N_27311,N_27502);
nand U29460 (N_29460,N_27713,N_27115);
and U29461 (N_29461,N_27994,N_27178);
or U29462 (N_29462,N_27904,N_28260);
xnor U29463 (N_29463,N_27497,N_27951);
or U29464 (N_29464,N_27653,N_27274);
nor U29465 (N_29465,N_27573,N_28016);
xnor U29466 (N_29466,N_27309,N_27660);
nand U29467 (N_29467,N_27132,N_27349);
nor U29468 (N_29468,N_27813,N_27865);
and U29469 (N_29469,N_28177,N_27732);
nor U29470 (N_29470,N_28061,N_28386);
nor U29471 (N_29471,N_27502,N_28275);
xor U29472 (N_29472,N_27395,N_27700);
nor U29473 (N_29473,N_28224,N_28118);
nor U29474 (N_29474,N_27565,N_28432);
nand U29475 (N_29475,N_28422,N_28093);
and U29476 (N_29476,N_27743,N_27339);
nor U29477 (N_29477,N_27026,N_27273);
nor U29478 (N_29478,N_27917,N_27504);
nand U29479 (N_29479,N_28067,N_27296);
nor U29480 (N_29480,N_28226,N_27897);
nor U29481 (N_29481,N_27279,N_27715);
xnor U29482 (N_29482,N_27903,N_27333);
xor U29483 (N_29483,N_27933,N_28020);
nor U29484 (N_29484,N_27421,N_27022);
or U29485 (N_29485,N_27235,N_27616);
xor U29486 (N_29486,N_27569,N_28282);
nand U29487 (N_29487,N_27886,N_27940);
nor U29488 (N_29488,N_27649,N_27101);
and U29489 (N_29489,N_27159,N_27298);
xnor U29490 (N_29490,N_28178,N_28234);
xnor U29491 (N_29491,N_28408,N_27127);
nand U29492 (N_29492,N_27403,N_27447);
and U29493 (N_29493,N_27330,N_27692);
nand U29494 (N_29494,N_27428,N_28413);
xor U29495 (N_29495,N_27430,N_27973);
or U29496 (N_29496,N_27301,N_27710);
or U29497 (N_29497,N_27910,N_27566);
nand U29498 (N_29498,N_27916,N_27735);
xnor U29499 (N_29499,N_28436,N_27363);
nor U29500 (N_29500,N_28158,N_28275);
nor U29501 (N_29501,N_27125,N_28152);
and U29502 (N_29502,N_27060,N_27704);
xnor U29503 (N_29503,N_28259,N_27881);
xor U29504 (N_29504,N_28272,N_28230);
and U29505 (N_29505,N_27960,N_27957);
nand U29506 (N_29506,N_27971,N_28257);
or U29507 (N_29507,N_27112,N_27081);
nor U29508 (N_29508,N_27069,N_27665);
nor U29509 (N_29509,N_27756,N_27669);
nor U29510 (N_29510,N_27640,N_28397);
nor U29511 (N_29511,N_27958,N_27040);
or U29512 (N_29512,N_27699,N_28477);
nor U29513 (N_29513,N_27562,N_28385);
nand U29514 (N_29514,N_28312,N_27431);
or U29515 (N_29515,N_27864,N_28261);
or U29516 (N_29516,N_28345,N_28113);
and U29517 (N_29517,N_27997,N_27572);
and U29518 (N_29518,N_27086,N_28370);
xnor U29519 (N_29519,N_27529,N_28155);
nand U29520 (N_29520,N_27037,N_28216);
nor U29521 (N_29521,N_27457,N_28078);
nor U29522 (N_29522,N_27580,N_28186);
or U29523 (N_29523,N_28177,N_27871);
and U29524 (N_29524,N_28410,N_27782);
nor U29525 (N_29525,N_27957,N_27652);
and U29526 (N_29526,N_27333,N_28119);
xor U29527 (N_29527,N_27357,N_27047);
nand U29528 (N_29528,N_27130,N_28186);
or U29529 (N_29529,N_28247,N_27752);
or U29530 (N_29530,N_28094,N_27669);
xnor U29531 (N_29531,N_27716,N_27773);
nor U29532 (N_29532,N_28450,N_27761);
xnor U29533 (N_29533,N_28213,N_27582);
or U29534 (N_29534,N_27691,N_28416);
xor U29535 (N_29535,N_27025,N_27774);
nand U29536 (N_29536,N_27074,N_28461);
or U29537 (N_29537,N_27954,N_27427);
xor U29538 (N_29538,N_28348,N_28151);
or U29539 (N_29539,N_27268,N_28416);
or U29540 (N_29540,N_28014,N_27759);
and U29541 (N_29541,N_28113,N_27915);
and U29542 (N_29542,N_27289,N_28266);
and U29543 (N_29543,N_27029,N_27154);
xor U29544 (N_29544,N_27222,N_28268);
or U29545 (N_29545,N_27602,N_27905);
xor U29546 (N_29546,N_27453,N_27633);
nand U29547 (N_29547,N_28286,N_27897);
or U29548 (N_29548,N_27488,N_27899);
xor U29549 (N_29549,N_28462,N_27254);
or U29550 (N_29550,N_28094,N_27863);
or U29551 (N_29551,N_27251,N_28452);
or U29552 (N_29552,N_28347,N_28286);
nand U29553 (N_29553,N_28214,N_28002);
nor U29554 (N_29554,N_28094,N_28308);
nor U29555 (N_29555,N_27325,N_27441);
xnor U29556 (N_29556,N_28214,N_27275);
nor U29557 (N_29557,N_27001,N_28125);
and U29558 (N_29558,N_27598,N_27935);
nor U29559 (N_29559,N_28480,N_28328);
nor U29560 (N_29560,N_27913,N_27258);
xnor U29561 (N_29561,N_28103,N_28294);
xnor U29562 (N_29562,N_27772,N_27327);
nor U29563 (N_29563,N_27317,N_28461);
and U29564 (N_29564,N_28419,N_28280);
nor U29565 (N_29565,N_27527,N_27304);
nand U29566 (N_29566,N_27646,N_27807);
and U29567 (N_29567,N_27432,N_27914);
and U29568 (N_29568,N_27325,N_27978);
and U29569 (N_29569,N_28028,N_28469);
nand U29570 (N_29570,N_28291,N_27820);
and U29571 (N_29571,N_28333,N_27820);
nor U29572 (N_29572,N_27992,N_28086);
nor U29573 (N_29573,N_27581,N_27659);
nor U29574 (N_29574,N_27700,N_27028);
nor U29575 (N_29575,N_27004,N_28442);
or U29576 (N_29576,N_27650,N_27453);
nor U29577 (N_29577,N_27156,N_27544);
and U29578 (N_29578,N_27146,N_27455);
or U29579 (N_29579,N_27575,N_27275);
or U29580 (N_29580,N_28028,N_27625);
and U29581 (N_29581,N_27451,N_27838);
and U29582 (N_29582,N_27937,N_27634);
nor U29583 (N_29583,N_27516,N_28363);
and U29584 (N_29584,N_28143,N_27015);
and U29585 (N_29585,N_27917,N_27118);
nand U29586 (N_29586,N_27875,N_27195);
nor U29587 (N_29587,N_27710,N_28026);
or U29588 (N_29588,N_28119,N_27282);
and U29589 (N_29589,N_28021,N_28278);
or U29590 (N_29590,N_27542,N_27581);
xor U29591 (N_29591,N_28289,N_27410);
xnor U29592 (N_29592,N_27391,N_27894);
nor U29593 (N_29593,N_27407,N_27809);
xnor U29594 (N_29594,N_27390,N_27859);
and U29595 (N_29595,N_27170,N_27854);
or U29596 (N_29596,N_27767,N_27152);
nor U29597 (N_29597,N_28340,N_27337);
xnor U29598 (N_29598,N_28147,N_27533);
or U29599 (N_29599,N_27221,N_28232);
and U29600 (N_29600,N_28129,N_27962);
or U29601 (N_29601,N_27191,N_27492);
nand U29602 (N_29602,N_28485,N_27771);
nor U29603 (N_29603,N_28449,N_27278);
and U29604 (N_29604,N_28460,N_28301);
and U29605 (N_29605,N_27277,N_27810);
xnor U29606 (N_29606,N_28260,N_27051);
and U29607 (N_29607,N_27033,N_27517);
or U29608 (N_29608,N_27318,N_27872);
nor U29609 (N_29609,N_27912,N_27731);
nand U29610 (N_29610,N_27853,N_28125);
nand U29611 (N_29611,N_27626,N_28397);
xnor U29612 (N_29612,N_27193,N_27976);
nor U29613 (N_29613,N_28428,N_27996);
or U29614 (N_29614,N_27120,N_27747);
xor U29615 (N_29615,N_27555,N_27952);
and U29616 (N_29616,N_28399,N_28010);
and U29617 (N_29617,N_27561,N_28136);
nand U29618 (N_29618,N_27615,N_28211);
nand U29619 (N_29619,N_28283,N_27470);
nand U29620 (N_29620,N_27399,N_28087);
xnor U29621 (N_29621,N_27261,N_27577);
and U29622 (N_29622,N_28356,N_27756);
and U29623 (N_29623,N_28313,N_27074);
nand U29624 (N_29624,N_28444,N_27109);
and U29625 (N_29625,N_28243,N_27914);
xor U29626 (N_29626,N_27963,N_28115);
or U29627 (N_29627,N_27575,N_28091);
and U29628 (N_29628,N_27921,N_28032);
xor U29629 (N_29629,N_28317,N_27163);
nor U29630 (N_29630,N_27158,N_28369);
xor U29631 (N_29631,N_27073,N_27244);
nor U29632 (N_29632,N_28030,N_28253);
nand U29633 (N_29633,N_27993,N_28255);
or U29634 (N_29634,N_27606,N_28111);
xnor U29635 (N_29635,N_27308,N_27059);
xor U29636 (N_29636,N_27694,N_27182);
nor U29637 (N_29637,N_27196,N_28062);
and U29638 (N_29638,N_27248,N_28063);
nand U29639 (N_29639,N_28113,N_27394);
nor U29640 (N_29640,N_27799,N_27159);
xor U29641 (N_29641,N_28310,N_28447);
nor U29642 (N_29642,N_27909,N_27749);
or U29643 (N_29643,N_27230,N_27040);
xor U29644 (N_29644,N_27920,N_28326);
and U29645 (N_29645,N_27896,N_28007);
xor U29646 (N_29646,N_27772,N_27858);
nor U29647 (N_29647,N_27939,N_27132);
xor U29648 (N_29648,N_27225,N_27809);
xnor U29649 (N_29649,N_27808,N_28492);
xnor U29650 (N_29650,N_27592,N_27573);
or U29651 (N_29651,N_28188,N_28255);
and U29652 (N_29652,N_27251,N_27604);
nor U29653 (N_29653,N_27227,N_27817);
and U29654 (N_29654,N_27501,N_27623);
nor U29655 (N_29655,N_28409,N_27469);
xnor U29656 (N_29656,N_27095,N_27252);
nand U29657 (N_29657,N_27507,N_27280);
nand U29658 (N_29658,N_28185,N_28404);
xor U29659 (N_29659,N_27387,N_27679);
nand U29660 (N_29660,N_27307,N_28315);
and U29661 (N_29661,N_28268,N_27269);
nor U29662 (N_29662,N_27404,N_28471);
and U29663 (N_29663,N_28338,N_27563);
and U29664 (N_29664,N_28377,N_27299);
xnor U29665 (N_29665,N_27601,N_27016);
xor U29666 (N_29666,N_28351,N_28498);
nand U29667 (N_29667,N_28429,N_27118);
nand U29668 (N_29668,N_27389,N_27546);
xor U29669 (N_29669,N_27854,N_27425);
nand U29670 (N_29670,N_28013,N_27101);
and U29671 (N_29671,N_28347,N_27951);
or U29672 (N_29672,N_28336,N_27140);
xor U29673 (N_29673,N_27218,N_27142);
xor U29674 (N_29674,N_27032,N_27482);
and U29675 (N_29675,N_28476,N_27242);
and U29676 (N_29676,N_27151,N_27606);
nand U29677 (N_29677,N_27563,N_27176);
or U29678 (N_29678,N_27644,N_28039);
nand U29679 (N_29679,N_27061,N_28389);
or U29680 (N_29680,N_27462,N_27118);
nor U29681 (N_29681,N_27317,N_28362);
or U29682 (N_29682,N_27135,N_28287);
nor U29683 (N_29683,N_27616,N_28493);
and U29684 (N_29684,N_27476,N_27458);
nor U29685 (N_29685,N_28494,N_28250);
and U29686 (N_29686,N_27090,N_27784);
xnor U29687 (N_29687,N_28238,N_28125);
and U29688 (N_29688,N_28366,N_27162);
or U29689 (N_29689,N_27312,N_28464);
nand U29690 (N_29690,N_27063,N_27136);
xor U29691 (N_29691,N_28040,N_27425);
or U29692 (N_29692,N_28234,N_27864);
nand U29693 (N_29693,N_28073,N_27800);
nand U29694 (N_29694,N_28425,N_28113);
nand U29695 (N_29695,N_27044,N_28123);
nand U29696 (N_29696,N_27332,N_27411);
nor U29697 (N_29697,N_27231,N_27411);
nor U29698 (N_29698,N_27815,N_27119);
nand U29699 (N_29699,N_27576,N_28228);
and U29700 (N_29700,N_27965,N_27369);
or U29701 (N_29701,N_27418,N_27949);
nor U29702 (N_29702,N_27014,N_27337);
xnor U29703 (N_29703,N_27321,N_28153);
nor U29704 (N_29704,N_28353,N_27825);
and U29705 (N_29705,N_27968,N_27709);
or U29706 (N_29706,N_27778,N_27590);
and U29707 (N_29707,N_28059,N_28433);
and U29708 (N_29708,N_27669,N_28377);
and U29709 (N_29709,N_27087,N_27319);
nor U29710 (N_29710,N_28240,N_28417);
and U29711 (N_29711,N_28489,N_28415);
xnor U29712 (N_29712,N_27323,N_28019);
nor U29713 (N_29713,N_28054,N_27347);
or U29714 (N_29714,N_27718,N_27817);
nand U29715 (N_29715,N_28003,N_27081);
nand U29716 (N_29716,N_27942,N_27658);
nor U29717 (N_29717,N_27222,N_28033);
xnor U29718 (N_29718,N_28344,N_28056);
nand U29719 (N_29719,N_27852,N_28209);
nand U29720 (N_29720,N_27697,N_28168);
nand U29721 (N_29721,N_27811,N_27035);
and U29722 (N_29722,N_27487,N_27289);
nor U29723 (N_29723,N_27625,N_28236);
xor U29724 (N_29724,N_28179,N_27549);
xnor U29725 (N_29725,N_27094,N_27725);
nand U29726 (N_29726,N_28365,N_27108);
nor U29727 (N_29727,N_28094,N_28091);
xor U29728 (N_29728,N_27291,N_27464);
or U29729 (N_29729,N_27939,N_27517);
and U29730 (N_29730,N_27704,N_27250);
nand U29731 (N_29731,N_27505,N_28178);
xnor U29732 (N_29732,N_27899,N_27125);
nand U29733 (N_29733,N_27674,N_27577);
nor U29734 (N_29734,N_27293,N_27028);
nor U29735 (N_29735,N_27986,N_27572);
and U29736 (N_29736,N_27277,N_27664);
nand U29737 (N_29737,N_27908,N_28226);
and U29738 (N_29738,N_27283,N_27228);
xor U29739 (N_29739,N_28100,N_28013);
and U29740 (N_29740,N_27103,N_27645);
xnor U29741 (N_29741,N_27486,N_27839);
xor U29742 (N_29742,N_27640,N_27650);
nor U29743 (N_29743,N_28339,N_28326);
nor U29744 (N_29744,N_27550,N_28103);
and U29745 (N_29745,N_27701,N_27525);
xor U29746 (N_29746,N_28260,N_27386);
or U29747 (N_29747,N_27293,N_28414);
or U29748 (N_29748,N_28293,N_27188);
and U29749 (N_29749,N_28117,N_27756);
nor U29750 (N_29750,N_28098,N_28478);
xor U29751 (N_29751,N_27401,N_27717);
or U29752 (N_29752,N_27226,N_28426);
nand U29753 (N_29753,N_27986,N_27000);
or U29754 (N_29754,N_27508,N_27764);
and U29755 (N_29755,N_27922,N_27753);
or U29756 (N_29756,N_28066,N_27346);
nor U29757 (N_29757,N_28377,N_27778);
xnor U29758 (N_29758,N_27163,N_27804);
nor U29759 (N_29759,N_28012,N_27091);
and U29760 (N_29760,N_27495,N_27157);
and U29761 (N_29761,N_27651,N_28300);
nand U29762 (N_29762,N_27031,N_27400);
nand U29763 (N_29763,N_28063,N_27800);
nand U29764 (N_29764,N_27604,N_27599);
and U29765 (N_29765,N_27473,N_27040);
or U29766 (N_29766,N_28172,N_28117);
xnor U29767 (N_29767,N_27028,N_27637);
nor U29768 (N_29768,N_28234,N_28139);
or U29769 (N_29769,N_28335,N_28123);
xor U29770 (N_29770,N_28213,N_28443);
and U29771 (N_29771,N_27443,N_27022);
nand U29772 (N_29772,N_28180,N_27962);
nand U29773 (N_29773,N_28325,N_27731);
and U29774 (N_29774,N_27760,N_28206);
nor U29775 (N_29775,N_27266,N_27917);
nand U29776 (N_29776,N_27178,N_27532);
xor U29777 (N_29777,N_27368,N_28476);
nand U29778 (N_29778,N_28235,N_27137);
nand U29779 (N_29779,N_27310,N_28332);
xor U29780 (N_29780,N_27635,N_27368);
or U29781 (N_29781,N_28294,N_28107);
or U29782 (N_29782,N_27816,N_27209);
xor U29783 (N_29783,N_28037,N_27132);
nor U29784 (N_29784,N_27501,N_28443);
and U29785 (N_29785,N_28390,N_28180);
nand U29786 (N_29786,N_28381,N_28008);
xor U29787 (N_29787,N_28116,N_27119);
xnor U29788 (N_29788,N_27234,N_27187);
and U29789 (N_29789,N_27290,N_28304);
and U29790 (N_29790,N_27817,N_28455);
nor U29791 (N_29791,N_27886,N_27298);
and U29792 (N_29792,N_27533,N_27178);
nand U29793 (N_29793,N_27218,N_27521);
nor U29794 (N_29794,N_28271,N_27028);
or U29795 (N_29795,N_28022,N_27020);
nor U29796 (N_29796,N_27595,N_27242);
nand U29797 (N_29797,N_27384,N_28369);
or U29798 (N_29798,N_27105,N_27434);
nor U29799 (N_29799,N_28407,N_27540);
xor U29800 (N_29800,N_27336,N_27643);
or U29801 (N_29801,N_27739,N_28446);
xnor U29802 (N_29802,N_27926,N_28146);
nand U29803 (N_29803,N_27349,N_27690);
xnor U29804 (N_29804,N_27129,N_28155);
or U29805 (N_29805,N_27281,N_27534);
or U29806 (N_29806,N_28197,N_27462);
xor U29807 (N_29807,N_28071,N_27034);
nand U29808 (N_29808,N_27234,N_28362);
and U29809 (N_29809,N_27777,N_27171);
xnor U29810 (N_29810,N_27970,N_28378);
xnor U29811 (N_29811,N_27968,N_27243);
or U29812 (N_29812,N_27606,N_28031);
nor U29813 (N_29813,N_28333,N_27806);
nand U29814 (N_29814,N_27093,N_27779);
nand U29815 (N_29815,N_27591,N_27296);
nor U29816 (N_29816,N_27083,N_27530);
and U29817 (N_29817,N_27124,N_27686);
or U29818 (N_29818,N_27480,N_27076);
xor U29819 (N_29819,N_28200,N_28290);
nand U29820 (N_29820,N_28221,N_27020);
and U29821 (N_29821,N_27760,N_27612);
nand U29822 (N_29822,N_28249,N_27652);
and U29823 (N_29823,N_28345,N_27110);
and U29824 (N_29824,N_28194,N_27090);
or U29825 (N_29825,N_27144,N_27410);
xnor U29826 (N_29826,N_28359,N_27217);
xnor U29827 (N_29827,N_28474,N_27543);
and U29828 (N_29828,N_27564,N_28261);
or U29829 (N_29829,N_27716,N_27460);
or U29830 (N_29830,N_27564,N_27413);
xnor U29831 (N_29831,N_27479,N_27344);
nand U29832 (N_29832,N_28489,N_27609);
or U29833 (N_29833,N_27247,N_27193);
xor U29834 (N_29834,N_27750,N_27078);
xnor U29835 (N_29835,N_28271,N_28000);
xor U29836 (N_29836,N_27796,N_27247);
and U29837 (N_29837,N_28208,N_27351);
or U29838 (N_29838,N_27036,N_27238);
xor U29839 (N_29839,N_27511,N_28113);
nor U29840 (N_29840,N_27549,N_28289);
and U29841 (N_29841,N_28459,N_27871);
nand U29842 (N_29842,N_27683,N_27513);
nand U29843 (N_29843,N_27672,N_27596);
or U29844 (N_29844,N_28239,N_28166);
xor U29845 (N_29845,N_28384,N_27996);
xor U29846 (N_29846,N_27599,N_27870);
or U29847 (N_29847,N_28483,N_28217);
nor U29848 (N_29848,N_27794,N_27549);
or U29849 (N_29849,N_27092,N_28386);
xor U29850 (N_29850,N_28174,N_28208);
xor U29851 (N_29851,N_28324,N_27631);
nor U29852 (N_29852,N_27957,N_28085);
or U29853 (N_29853,N_28359,N_28300);
and U29854 (N_29854,N_28383,N_27273);
and U29855 (N_29855,N_27675,N_27291);
or U29856 (N_29856,N_28187,N_27416);
xor U29857 (N_29857,N_27399,N_28251);
xor U29858 (N_29858,N_27372,N_27265);
xor U29859 (N_29859,N_28172,N_28378);
or U29860 (N_29860,N_27499,N_28351);
nor U29861 (N_29861,N_28270,N_27682);
or U29862 (N_29862,N_27373,N_27291);
nand U29863 (N_29863,N_27382,N_27837);
and U29864 (N_29864,N_28294,N_27320);
nor U29865 (N_29865,N_28008,N_27368);
nand U29866 (N_29866,N_28468,N_27074);
nand U29867 (N_29867,N_27200,N_27369);
xor U29868 (N_29868,N_27613,N_28173);
nand U29869 (N_29869,N_28034,N_28218);
or U29870 (N_29870,N_28434,N_27035);
or U29871 (N_29871,N_27679,N_28089);
nand U29872 (N_29872,N_27189,N_28326);
or U29873 (N_29873,N_27128,N_27900);
or U29874 (N_29874,N_27333,N_27579);
nor U29875 (N_29875,N_28259,N_27885);
or U29876 (N_29876,N_27759,N_27103);
nor U29877 (N_29877,N_28088,N_27469);
or U29878 (N_29878,N_27949,N_27699);
nand U29879 (N_29879,N_27478,N_27717);
or U29880 (N_29880,N_27330,N_28057);
xnor U29881 (N_29881,N_27795,N_27799);
or U29882 (N_29882,N_27520,N_28424);
xor U29883 (N_29883,N_27250,N_28247);
or U29884 (N_29884,N_27446,N_28322);
nand U29885 (N_29885,N_28275,N_28448);
nor U29886 (N_29886,N_27322,N_28324);
and U29887 (N_29887,N_27272,N_27129);
nand U29888 (N_29888,N_27219,N_27121);
nor U29889 (N_29889,N_27758,N_27002);
nand U29890 (N_29890,N_27311,N_28094);
or U29891 (N_29891,N_27114,N_28343);
xor U29892 (N_29892,N_27415,N_28352);
xor U29893 (N_29893,N_27859,N_27395);
or U29894 (N_29894,N_28350,N_27739);
nand U29895 (N_29895,N_27319,N_28467);
or U29896 (N_29896,N_28192,N_27911);
or U29897 (N_29897,N_27327,N_27386);
or U29898 (N_29898,N_27849,N_27087);
nand U29899 (N_29899,N_27195,N_28472);
and U29900 (N_29900,N_27557,N_28044);
nand U29901 (N_29901,N_28086,N_27347);
nand U29902 (N_29902,N_27072,N_27960);
nand U29903 (N_29903,N_27052,N_28440);
and U29904 (N_29904,N_27030,N_27674);
nand U29905 (N_29905,N_27390,N_27418);
or U29906 (N_29906,N_27954,N_27941);
xor U29907 (N_29907,N_28050,N_27670);
or U29908 (N_29908,N_27221,N_27044);
nand U29909 (N_29909,N_27367,N_27374);
xor U29910 (N_29910,N_28056,N_28426);
nor U29911 (N_29911,N_28095,N_28291);
and U29912 (N_29912,N_27170,N_27973);
nor U29913 (N_29913,N_27712,N_27029);
nand U29914 (N_29914,N_28076,N_28074);
nand U29915 (N_29915,N_27471,N_27329);
nor U29916 (N_29916,N_27113,N_27386);
and U29917 (N_29917,N_27937,N_27068);
xor U29918 (N_29918,N_27049,N_28499);
xnor U29919 (N_29919,N_28350,N_28494);
or U29920 (N_29920,N_27004,N_27910);
xnor U29921 (N_29921,N_27861,N_28343);
nor U29922 (N_29922,N_27647,N_27916);
and U29923 (N_29923,N_27957,N_27331);
or U29924 (N_29924,N_27726,N_28486);
xor U29925 (N_29925,N_28162,N_28100);
nor U29926 (N_29926,N_27732,N_27719);
or U29927 (N_29927,N_28122,N_27828);
xnor U29928 (N_29928,N_28423,N_27053);
or U29929 (N_29929,N_27645,N_27785);
nand U29930 (N_29930,N_27232,N_27354);
nor U29931 (N_29931,N_27468,N_27087);
nor U29932 (N_29932,N_28435,N_28136);
and U29933 (N_29933,N_28131,N_27976);
nor U29934 (N_29934,N_27778,N_28274);
or U29935 (N_29935,N_28091,N_27244);
nand U29936 (N_29936,N_27054,N_27487);
xnor U29937 (N_29937,N_27593,N_27509);
xnor U29938 (N_29938,N_27128,N_27743);
and U29939 (N_29939,N_27996,N_28174);
xor U29940 (N_29940,N_27029,N_28422);
and U29941 (N_29941,N_28074,N_27373);
xnor U29942 (N_29942,N_28337,N_27376);
xor U29943 (N_29943,N_28410,N_28489);
and U29944 (N_29944,N_28018,N_28440);
nor U29945 (N_29945,N_27774,N_27083);
nor U29946 (N_29946,N_28278,N_27267);
nor U29947 (N_29947,N_28487,N_28478);
nor U29948 (N_29948,N_28322,N_27787);
and U29949 (N_29949,N_27144,N_27878);
nor U29950 (N_29950,N_27327,N_27759);
or U29951 (N_29951,N_28028,N_27763);
or U29952 (N_29952,N_28489,N_27533);
xor U29953 (N_29953,N_27851,N_27674);
or U29954 (N_29954,N_27311,N_28156);
and U29955 (N_29955,N_28461,N_27457);
or U29956 (N_29956,N_27741,N_27222);
and U29957 (N_29957,N_27167,N_28170);
nand U29958 (N_29958,N_27684,N_28466);
and U29959 (N_29959,N_27096,N_27750);
or U29960 (N_29960,N_28185,N_27696);
and U29961 (N_29961,N_27137,N_27369);
nor U29962 (N_29962,N_27164,N_27378);
nand U29963 (N_29963,N_27290,N_28172);
nor U29964 (N_29964,N_27286,N_27897);
xor U29965 (N_29965,N_27368,N_28142);
or U29966 (N_29966,N_27405,N_28066);
or U29967 (N_29967,N_27759,N_27543);
nor U29968 (N_29968,N_27707,N_27706);
nor U29969 (N_29969,N_27087,N_27632);
xnor U29970 (N_29970,N_27456,N_27473);
xnor U29971 (N_29971,N_27246,N_27562);
nor U29972 (N_29972,N_28267,N_27279);
xnor U29973 (N_29973,N_27836,N_27788);
or U29974 (N_29974,N_28422,N_27209);
xor U29975 (N_29975,N_27521,N_28459);
and U29976 (N_29976,N_27374,N_27863);
nand U29977 (N_29977,N_27231,N_27919);
and U29978 (N_29978,N_27247,N_27498);
and U29979 (N_29979,N_27910,N_27557);
xnor U29980 (N_29980,N_27001,N_27171);
nor U29981 (N_29981,N_27112,N_27020);
nor U29982 (N_29982,N_28449,N_28040);
nor U29983 (N_29983,N_27484,N_27728);
or U29984 (N_29984,N_28393,N_27950);
and U29985 (N_29985,N_28102,N_27278);
nor U29986 (N_29986,N_27173,N_27292);
or U29987 (N_29987,N_27876,N_28474);
xnor U29988 (N_29988,N_28216,N_27112);
or U29989 (N_29989,N_27739,N_28268);
xnor U29990 (N_29990,N_28029,N_27463);
nand U29991 (N_29991,N_27902,N_27702);
nand U29992 (N_29992,N_27775,N_27257);
or U29993 (N_29993,N_27453,N_28497);
nor U29994 (N_29994,N_27637,N_27931);
nand U29995 (N_29995,N_28473,N_27309);
xor U29996 (N_29996,N_27653,N_27830);
nor U29997 (N_29997,N_27465,N_27091);
nand U29998 (N_29998,N_27864,N_28094);
and U29999 (N_29999,N_27917,N_27107);
and UO_0 (O_0,N_29054,N_28747);
or UO_1 (O_1,N_29508,N_28846);
and UO_2 (O_2,N_29643,N_29547);
nand UO_3 (O_3,N_29183,N_28556);
and UO_4 (O_4,N_28889,N_28604);
or UO_5 (O_5,N_29801,N_29088);
nand UO_6 (O_6,N_29991,N_29933);
xnor UO_7 (O_7,N_29463,N_29514);
xor UO_8 (O_8,N_29553,N_29256);
xnor UO_9 (O_9,N_29734,N_29525);
nand UO_10 (O_10,N_29151,N_28674);
xor UO_11 (O_11,N_29894,N_29860);
nor UO_12 (O_12,N_28797,N_28880);
xor UO_13 (O_13,N_29081,N_28829);
and UO_14 (O_14,N_29606,N_29021);
and UO_15 (O_15,N_29273,N_29826);
nand UO_16 (O_16,N_28985,N_29414);
xor UO_17 (O_17,N_28585,N_29371);
xor UO_18 (O_18,N_29281,N_29465);
nand UO_19 (O_19,N_29964,N_29951);
and UO_20 (O_20,N_29560,N_28969);
nand UO_21 (O_21,N_28714,N_29107);
or UO_22 (O_22,N_28896,N_28993);
and UO_23 (O_23,N_28529,N_29248);
nor UO_24 (O_24,N_29315,N_29191);
and UO_25 (O_25,N_29206,N_29272);
xor UO_26 (O_26,N_28678,N_29024);
xor UO_27 (O_27,N_28502,N_29989);
nor UO_28 (O_28,N_28720,N_29356);
nor UO_29 (O_29,N_29889,N_28620);
nor UO_30 (O_30,N_29457,N_29203);
nand UO_31 (O_31,N_29638,N_28961);
xor UO_32 (O_32,N_29723,N_29476);
xnor UO_33 (O_33,N_28559,N_28960);
or UO_34 (O_34,N_29498,N_28971);
nand UO_35 (O_35,N_28858,N_28723);
and UO_36 (O_36,N_29510,N_29393);
or UO_37 (O_37,N_29763,N_28929);
or UO_38 (O_38,N_29400,N_28534);
nor UO_39 (O_39,N_29780,N_28525);
xor UO_40 (O_40,N_28671,N_29350);
nand UO_41 (O_41,N_29701,N_29098);
nand UO_42 (O_42,N_29661,N_28700);
nand UO_43 (O_43,N_29781,N_29155);
xor UO_44 (O_44,N_29026,N_29806);
xor UO_45 (O_45,N_28857,N_29741);
xor UO_46 (O_46,N_28976,N_28801);
nor UO_47 (O_47,N_29527,N_29629);
or UO_48 (O_48,N_29852,N_29872);
nor UO_49 (O_49,N_29885,N_29966);
xor UO_50 (O_50,N_28580,N_29192);
nor UO_51 (O_51,N_29009,N_29022);
nor UO_52 (O_52,N_29302,N_28980);
xnor UO_53 (O_53,N_29607,N_29693);
nand UO_54 (O_54,N_29091,N_29044);
or UO_55 (O_55,N_28709,N_28788);
nand UO_56 (O_56,N_28560,N_28835);
and UO_57 (O_57,N_29522,N_29374);
or UO_58 (O_58,N_28901,N_29784);
nand UO_59 (O_59,N_29467,N_29268);
nor UO_60 (O_60,N_29765,N_29555);
and UO_61 (O_61,N_29039,N_29311);
nor UO_62 (O_62,N_29908,N_29848);
nand UO_63 (O_63,N_29533,N_28856);
or UO_64 (O_64,N_29717,N_28509);
xnor UO_65 (O_65,N_29450,N_29140);
nor UO_66 (O_66,N_29916,N_28806);
nand UO_67 (O_67,N_29484,N_29559);
nand UO_68 (O_68,N_29125,N_29278);
and UO_69 (O_69,N_28883,N_28643);
or UO_70 (O_70,N_29178,N_29149);
xnor UO_71 (O_71,N_29925,N_28787);
nor UO_72 (O_72,N_29391,N_29516);
nor UO_73 (O_73,N_29007,N_29558);
or UO_74 (O_74,N_29317,N_29095);
or UO_75 (O_75,N_29086,N_28996);
nor UO_76 (O_76,N_29697,N_29422);
or UO_77 (O_77,N_29029,N_29728);
nor UO_78 (O_78,N_28679,N_28545);
nor UO_79 (O_79,N_29347,N_28869);
nand UO_80 (O_80,N_29689,N_29677);
and UO_81 (O_81,N_28943,N_29799);
xor UO_82 (O_82,N_29865,N_28802);
xnor UO_83 (O_83,N_29645,N_29482);
xnor UO_84 (O_84,N_29575,N_29819);
nand UO_85 (O_85,N_28780,N_29491);
xor UO_86 (O_86,N_29232,N_29242);
and UO_87 (O_87,N_29705,N_28719);
and UO_88 (O_88,N_29968,N_29504);
nand UO_89 (O_89,N_29985,N_29500);
or UO_90 (O_90,N_28742,N_29461);
and UO_91 (O_91,N_29681,N_29941);
nor UO_92 (O_92,N_29818,N_28501);
xnor UO_93 (O_93,N_29675,N_28602);
xnor UO_94 (O_94,N_29950,N_29145);
and UO_95 (O_95,N_29593,N_28586);
xnor UO_96 (O_96,N_29032,N_29298);
xor UO_97 (O_97,N_29882,N_28812);
nor UO_98 (O_98,N_28956,N_28844);
and UO_99 (O_99,N_29481,N_29297);
and UO_100 (O_100,N_29313,N_29637);
and UO_101 (O_101,N_29582,N_29287);
or UO_102 (O_102,N_29770,N_29445);
nand UO_103 (O_103,N_28763,N_28800);
or UO_104 (O_104,N_29346,N_29518);
and UO_105 (O_105,N_29895,N_29390);
nand UO_106 (O_106,N_29167,N_28799);
xnor UO_107 (O_107,N_28725,N_28813);
or UO_108 (O_108,N_29613,N_29126);
nor UO_109 (O_109,N_29057,N_28745);
nand UO_110 (O_110,N_29303,N_29221);
or UO_111 (O_111,N_29674,N_29724);
or UO_112 (O_112,N_29364,N_29322);
xnor UO_113 (O_113,N_29434,N_29477);
nand UO_114 (O_114,N_29222,N_29657);
nand UO_115 (O_115,N_29425,N_28575);
or UO_116 (O_116,N_28652,N_29727);
nor UO_117 (O_117,N_28867,N_28931);
xnor UO_118 (O_118,N_29539,N_29932);
nor UO_119 (O_119,N_29887,N_28694);
nand UO_120 (O_120,N_29517,N_29744);
nor UO_121 (O_121,N_29199,N_28818);
xor UO_122 (O_122,N_28776,N_28657);
or UO_123 (O_123,N_29905,N_29284);
xor UO_124 (O_124,N_29580,N_29977);
and UO_125 (O_125,N_28614,N_29658);
and UO_126 (O_126,N_28630,N_28999);
nor UO_127 (O_127,N_29305,N_29684);
or UO_128 (O_128,N_29405,N_28702);
nand UO_129 (O_129,N_28979,N_28954);
nand UO_130 (O_130,N_28957,N_28850);
nor UO_131 (O_131,N_29033,N_29137);
nor UO_132 (O_132,N_29190,N_29802);
nor UO_133 (O_133,N_29402,N_29725);
and UO_134 (O_134,N_29992,N_29787);
or UO_135 (O_135,N_29075,N_29954);
xnor UO_136 (O_136,N_28705,N_28953);
xor UO_137 (O_137,N_29511,N_29479);
nor UO_138 (O_138,N_29016,N_28753);
and UO_139 (O_139,N_29939,N_29336);
and UO_140 (O_140,N_28734,N_29587);
nor UO_141 (O_141,N_28526,N_29691);
xnor UO_142 (O_142,N_28965,N_28613);
or UO_143 (O_143,N_29300,N_29170);
nor UO_144 (O_144,N_29421,N_28924);
nand UO_145 (O_145,N_28591,N_29225);
or UO_146 (O_146,N_28661,N_29620);
nor UO_147 (O_147,N_28918,N_29254);
nand UO_148 (O_148,N_29220,N_29460);
or UO_149 (O_149,N_28899,N_28992);
nor UO_150 (O_150,N_29357,N_29644);
nand UO_151 (O_151,N_28722,N_28530);
xor UO_152 (O_152,N_29093,N_28506);
and UO_153 (O_153,N_29902,N_29399);
or UO_154 (O_154,N_29233,N_29726);
nand UO_155 (O_155,N_29378,N_29280);
and UO_156 (O_156,N_28544,N_28547);
nor UO_157 (O_157,N_29212,N_29045);
or UO_158 (O_158,N_29528,N_28728);
nand UO_159 (O_159,N_28555,N_29569);
nand UO_160 (O_160,N_29270,N_29142);
or UO_161 (O_161,N_28771,N_29288);
xor UO_162 (O_162,N_29940,N_29229);
and UO_163 (O_163,N_29169,N_29005);
nand UO_164 (O_164,N_29634,N_29890);
or UO_165 (O_165,N_29217,N_29179);
nand UO_166 (O_166,N_28903,N_28936);
or UO_167 (O_167,N_28796,N_29490);
or UO_168 (O_168,N_28733,N_29168);
nand UO_169 (O_169,N_28981,N_28941);
xor UO_170 (O_170,N_29439,N_29963);
or UO_171 (O_171,N_29017,N_29130);
nand UO_172 (O_172,N_29538,N_29843);
xnor UO_173 (O_173,N_29507,N_29639);
and UO_174 (O_174,N_29811,N_28904);
nor UO_175 (O_175,N_29201,N_29863);
or UO_176 (O_176,N_29831,N_29108);
xor UO_177 (O_177,N_28807,N_29240);
and UO_178 (O_178,N_29856,N_29878);
or UO_179 (O_179,N_28647,N_29551);
and UO_180 (O_180,N_28637,N_29214);
xor UO_181 (O_181,N_29603,N_29982);
xor UO_182 (O_182,N_29216,N_29234);
nor UO_183 (O_183,N_29789,N_29330);
nor UO_184 (O_184,N_28754,N_29442);
and UO_185 (O_185,N_29830,N_29626);
and UO_186 (O_186,N_29002,N_29454);
nor UO_187 (O_187,N_29429,N_29565);
or UO_188 (O_188,N_29189,N_28540);
and UO_189 (O_189,N_29059,N_28810);
and UO_190 (O_190,N_29829,N_29880);
or UO_191 (O_191,N_28693,N_29523);
or UO_192 (O_192,N_29113,N_28503);
and UO_193 (O_193,N_29570,N_29124);
nand UO_194 (O_194,N_28589,N_29051);
and UO_195 (O_195,N_28911,N_29997);
nor UO_196 (O_196,N_28724,N_29325);
or UO_197 (O_197,N_28868,N_28762);
nand UO_198 (O_198,N_29572,N_29772);
nor UO_199 (O_199,N_28676,N_29680);
nor UO_200 (O_200,N_28665,N_29732);
and UO_201 (O_201,N_29420,N_29835);
and UO_202 (O_202,N_28794,N_28774);
nand UO_203 (O_203,N_29897,N_29244);
nand UO_204 (O_204,N_29839,N_29695);
and UO_205 (O_205,N_29837,N_29352);
nand UO_206 (O_206,N_29430,N_28877);
xnor UO_207 (O_207,N_29200,N_29064);
nand UO_208 (O_208,N_29825,N_29279);
xnor UO_209 (O_209,N_29836,N_28859);
nand UO_210 (O_210,N_28644,N_29253);
nand UO_211 (O_211,N_28949,N_29011);
nor UO_212 (O_212,N_29886,N_28793);
xnor UO_213 (O_213,N_28569,N_29102);
xor UO_214 (O_214,N_29785,N_29668);
xor UO_215 (O_215,N_29328,N_29573);
nand UO_216 (O_216,N_28595,N_29308);
nand UO_217 (O_217,N_29709,N_28898);
nor UO_218 (O_218,N_29803,N_29056);
nor UO_219 (O_219,N_28617,N_28703);
nand UO_220 (O_220,N_28914,N_29912);
nand UO_221 (O_221,N_29870,N_29990);
nor UO_222 (O_222,N_28521,N_28739);
nand UO_223 (O_223,N_28843,N_29683);
nand UO_224 (O_224,N_29584,N_28878);
or UO_225 (O_225,N_28716,N_28685);
and UO_226 (O_226,N_29568,N_29816);
xnor UO_227 (O_227,N_29259,N_29838);
nand UO_228 (O_228,N_28712,N_29773);
nand UO_229 (O_229,N_28891,N_29286);
nor UO_230 (O_230,N_29207,N_28633);
and UO_231 (O_231,N_29423,N_29814);
or UO_232 (O_232,N_28983,N_29269);
nor UO_233 (O_233,N_28950,N_29319);
or UO_234 (O_234,N_28792,N_28631);
or UO_235 (O_235,N_29704,N_28704);
nand UO_236 (O_236,N_29249,N_28650);
or UO_237 (O_237,N_29073,N_28554);
and UO_238 (O_238,N_29366,N_29502);
nor UO_239 (O_239,N_29735,N_28708);
nor UO_240 (O_240,N_28833,N_29060);
nor UO_241 (O_241,N_29031,N_29235);
nor UO_242 (O_242,N_29993,N_29731);
or UO_243 (O_243,N_29085,N_28565);
nand UO_244 (O_244,N_29118,N_28815);
and UO_245 (O_245,N_29129,N_29296);
nor UO_246 (O_246,N_29792,N_28582);
nand UO_247 (O_247,N_29141,N_29808);
and UO_248 (O_248,N_28975,N_28842);
and UO_249 (O_249,N_29299,N_28511);
nand UO_250 (O_250,N_29010,N_29664);
or UO_251 (O_251,N_28649,N_28594);
xor UO_252 (O_252,N_29715,N_29110);
and UO_253 (O_253,N_28860,N_29283);
nor UO_254 (O_254,N_29413,N_28915);
nand UO_255 (O_255,N_29426,N_29210);
or UO_256 (O_256,N_28849,N_29380);
nor UO_257 (O_257,N_28531,N_29497);
or UO_258 (O_258,N_29628,N_29080);
or UO_259 (O_259,N_29159,N_29219);
and UO_260 (O_260,N_29873,N_28938);
xor UO_261 (O_261,N_29550,N_28578);
xor UO_262 (O_262,N_29622,N_29228);
xor UO_263 (O_263,N_28504,N_29404);
xnor UO_264 (O_264,N_29632,N_28587);
or UO_265 (O_265,N_29227,N_28932);
nor UO_266 (O_266,N_29753,N_29903);
xnor UO_267 (O_267,N_29492,N_29275);
xor UO_268 (O_268,N_28851,N_28978);
and UO_269 (O_269,N_28951,N_29398);
and UO_270 (O_270,N_29358,N_29611);
xnor UO_271 (O_271,N_29961,N_29567);
and UO_272 (O_272,N_28513,N_29063);
nor UO_273 (O_273,N_29537,N_29354);
or UO_274 (O_274,N_29544,N_28832);
or UO_275 (O_275,N_29182,N_29708);
nor UO_276 (O_276,N_29237,N_29805);
xor UO_277 (O_277,N_29761,N_29438);
or UO_278 (O_278,N_29301,N_29769);
xor UO_279 (O_279,N_29771,N_29995);
nand UO_280 (O_280,N_29804,N_29304);
nand UO_281 (O_281,N_29659,N_29487);
xnor UO_282 (O_282,N_29410,N_28695);
and UO_283 (O_283,N_29911,N_29122);
nor UO_284 (O_284,N_29646,N_28872);
and UO_285 (O_285,N_29158,N_29036);
and UO_286 (O_286,N_29408,N_29791);
xnor UO_287 (O_287,N_29970,N_29417);
or UO_288 (O_288,N_29616,N_29764);
and UO_289 (O_289,N_28707,N_29180);
nor UO_290 (O_290,N_28748,N_29231);
nor UO_291 (O_291,N_28603,N_29174);
xnor UO_292 (O_292,N_29981,N_28579);
or UO_293 (O_293,N_28751,N_28567);
nor UO_294 (O_294,N_28536,N_28619);
or UO_295 (O_295,N_29250,N_29263);
and UO_296 (O_296,N_29447,N_29667);
and UO_297 (O_297,N_29333,N_28779);
and UO_298 (O_298,N_29337,N_29976);
or UO_299 (O_299,N_29810,N_29746);
nand UO_300 (O_300,N_28939,N_28744);
or UO_301 (O_301,N_29973,N_29071);
and UO_302 (O_302,N_29673,N_28824);
xnor UO_303 (O_303,N_29923,N_29419);
and UO_304 (O_304,N_29394,N_29261);
nand UO_305 (O_305,N_29412,N_29331);
nand UO_306 (O_306,N_28727,N_29285);
nand UO_307 (O_307,N_29758,N_29947);
and UO_308 (O_308,N_28928,N_29988);
nand UO_309 (O_309,N_28750,N_29849);
nor UO_310 (O_310,N_29891,N_28759);
nor UO_311 (O_311,N_29790,N_29562);
and UO_312 (O_312,N_29424,N_28615);
and UO_313 (O_313,N_29614,N_28863);
nand UO_314 (O_314,N_28618,N_29934);
and UO_315 (O_315,N_29531,N_29738);
and UO_316 (O_316,N_29332,N_29702);
nor UO_317 (O_317,N_29740,N_29166);
and UO_318 (O_318,N_29901,N_28923);
and UO_319 (O_319,N_28573,N_28522);
or UO_320 (O_320,N_29755,N_28684);
xor UO_321 (O_321,N_29822,N_28718);
and UO_322 (O_322,N_29640,N_29066);
or UO_323 (O_323,N_28523,N_28655);
and UO_324 (O_324,N_29707,N_29768);
xor UO_325 (O_325,N_28548,N_28596);
nand UO_326 (O_326,N_29416,N_29832);
nor UO_327 (O_327,N_29612,N_29660);
or UO_328 (O_328,N_29845,N_29339);
and UO_329 (O_329,N_29858,N_29062);
nand UO_330 (O_330,N_29750,N_29446);
nand UO_331 (O_331,N_28648,N_29716);
xnor UO_332 (O_332,N_29936,N_28970);
xnor UO_333 (O_333,N_29669,N_29209);
or UO_334 (O_334,N_28861,N_29969);
nor UO_335 (O_335,N_28786,N_29670);
or UO_336 (O_336,N_29957,N_29037);
or UO_337 (O_337,N_29195,N_29906);
nand UO_338 (O_338,N_29150,N_29376);
nor UO_339 (O_339,N_29453,N_29055);
xor UO_340 (O_340,N_28879,N_28730);
xor UO_341 (O_341,N_28895,N_29462);
nand UO_342 (O_342,N_29840,N_29774);
or UO_343 (O_343,N_29630,N_29899);
nand UO_344 (O_344,N_29942,N_29604);
and UO_345 (O_345,N_29441,N_28814);
nand UO_346 (O_346,N_28625,N_29312);
nand UO_347 (O_347,N_29069,N_29499);
or UO_348 (O_348,N_29967,N_28897);
nand UO_349 (O_349,N_29104,N_29058);
nor UO_350 (O_350,N_29318,N_29389);
nand UO_351 (O_351,N_29432,N_28775);
nand UO_352 (O_352,N_29271,N_29131);
xor UO_353 (O_353,N_29952,N_28638);
nor UO_354 (O_354,N_28549,N_29854);
nor UO_355 (O_355,N_29156,N_29900);
nor UO_356 (O_356,N_29935,N_29743);
xnor UO_357 (O_357,N_29241,N_28553);
or UO_358 (O_358,N_28538,N_28537);
and UO_359 (O_359,N_28566,N_29106);
nor UO_360 (O_360,N_29397,N_29184);
xor UO_361 (O_361,N_29139,N_29123);
nor UO_362 (O_362,N_28890,N_29003);
nor UO_363 (O_363,N_28873,N_29188);
xor UO_364 (O_364,N_29853,N_29436);
xnor UO_365 (O_365,N_29243,N_29898);
and UO_366 (O_366,N_29505,N_29605);
nand UO_367 (O_367,N_29842,N_28934);
or UO_368 (O_368,N_29996,N_29136);
nor UO_369 (O_369,N_28804,N_28917);
and UO_370 (O_370,N_29600,N_29914);
nand UO_371 (O_371,N_28527,N_28654);
nand UO_372 (O_372,N_28756,N_29355);
and UO_373 (O_373,N_29678,N_29049);
nor UO_374 (O_374,N_29395,N_29654);
nand UO_375 (O_375,N_29919,N_28701);
nand UO_376 (O_376,N_28601,N_29370);
nand UO_377 (O_377,N_29161,N_29160);
nor UO_378 (O_378,N_29172,N_28871);
nand UO_379 (O_379,N_29879,N_28838);
nor UO_380 (O_380,N_28598,N_29264);
xnor UO_381 (O_381,N_29987,N_29520);
or UO_382 (O_382,N_29909,N_29907);
nand UO_383 (O_383,N_29524,N_28822);
xor UO_384 (O_384,N_28721,N_28656);
or UO_385 (O_385,N_28584,N_29193);
nor UO_386 (O_386,N_29566,N_29546);
xor UO_387 (O_387,N_29353,N_28663);
and UO_388 (O_388,N_29928,N_29703);
xor UO_389 (O_389,N_28942,N_29592);
nor UO_390 (O_390,N_29515,N_29827);
nand UO_391 (O_391,N_29945,N_29962);
nand UO_392 (O_392,N_29030,N_29688);
and UO_393 (O_393,N_28680,N_28749);
or UO_394 (O_394,N_29470,N_29965);
nor UO_395 (O_395,N_29881,N_28827);
xnor UO_396 (O_396,N_29736,N_29023);
and UO_397 (O_397,N_29267,N_28768);
and UO_398 (O_398,N_29540,N_29314);
or UO_399 (O_399,N_29015,N_29164);
xor UO_400 (O_400,N_28855,N_29372);
xnor UO_401 (O_401,N_29089,N_29194);
and UO_402 (O_402,N_28532,N_28692);
xnor UO_403 (O_403,N_29653,N_29238);
or UO_404 (O_404,N_29449,N_29345);
and UO_405 (O_405,N_29767,N_28988);
xor UO_406 (O_406,N_29949,N_28533);
nand UO_407 (O_407,N_29588,N_28662);
and UO_408 (O_408,N_29642,N_28557);
nand UO_409 (O_409,N_29013,N_29114);
or UO_410 (O_410,N_28689,N_28885);
or UO_411 (O_411,N_29282,N_29722);
and UO_412 (O_412,N_28512,N_29795);
or UO_413 (O_413,N_29877,N_28845);
nand UO_414 (O_414,N_29586,N_28741);
and UO_415 (O_415,N_29087,N_28535);
and UO_416 (O_416,N_29888,N_28920);
nand UO_417 (O_417,N_29361,N_28852);
nand UO_418 (O_418,N_29589,N_29706);
or UO_419 (O_419,N_29101,N_28781);
xnor UO_420 (O_420,N_28516,N_28616);
nor UO_421 (O_421,N_28989,N_29921);
xnor UO_422 (O_422,N_29926,N_29742);
and UO_423 (O_423,N_29351,N_29014);
nand UO_424 (O_424,N_29618,N_29777);
and UO_425 (O_425,N_29134,N_28515);
and UO_426 (O_426,N_29163,N_29202);
or UO_427 (O_427,N_29809,N_28791);
or UO_428 (O_428,N_28974,N_29258);
xnor UO_429 (O_429,N_29309,N_29239);
or UO_430 (O_430,N_29197,N_28696);
xor UO_431 (O_431,N_29794,N_28933);
and UO_432 (O_432,N_28767,N_29496);
xor UO_433 (O_433,N_29262,N_29198);
and UO_434 (O_434,N_29624,N_29218);
nor UO_435 (O_435,N_29324,N_28621);
or UO_436 (O_436,N_28686,N_29748);
nand UO_437 (O_437,N_28823,N_28669);
or UO_438 (O_438,N_29652,N_29187);
or UO_439 (O_439,N_28769,N_29103);
or UO_440 (O_440,N_29096,N_28777);
and UO_441 (O_441,N_28706,N_29710);
nand UO_442 (O_442,N_29913,N_29672);
or UO_443 (O_443,N_29375,N_29291);
nand UO_444 (O_444,N_29247,N_28715);
nor UO_445 (O_445,N_28607,N_29224);
nand UO_446 (O_446,N_29685,N_29548);
and UO_447 (O_447,N_29115,N_29834);
nor UO_448 (O_448,N_29396,N_29974);
and UO_449 (O_449,N_28510,N_29177);
and UO_450 (O_450,N_28927,N_28610);
nor UO_451 (O_451,N_28605,N_29501);
nand UO_452 (O_452,N_28600,N_28760);
xor UO_453 (O_453,N_28524,N_29427);
nor UO_454 (O_454,N_28935,N_28593);
nor UO_455 (O_455,N_29367,N_28991);
and UO_456 (O_456,N_29876,N_29542);
nor UO_457 (O_457,N_28713,N_29931);
nand UO_458 (O_458,N_29448,N_28546);
xor UO_459 (O_459,N_29513,N_29257);
xor UO_460 (O_460,N_29100,N_29175);
xnor UO_461 (O_461,N_29379,N_29984);
nand UO_462 (O_462,N_28825,N_29557);
or UO_463 (O_463,N_28597,N_29117);
nand UO_464 (O_464,N_29671,N_29821);
nand UO_465 (O_465,N_28570,N_28562);
or UO_466 (O_466,N_28925,N_28726);
xnor UO_467 (O_467,N_29488,N_29363);
nand UO_468 (O_468,N_28922,N_29956);
nor UO_469 (O_469,N_28641,N_29368);
xor UO_470 (O_470,N_29998,N_29920);
nand UO_471 (O_471,N_29532,N_29290);
or UO_472 (O_472,N_28886,N_28893);
or UO_473 (O_473,N_28913,N_29910);
xor UO_474 (O_474,N_28977,N_28926);
nand UO_475 (O_475,N_29721,N_28987);
nand UO_476 (O_476,N_29937,N_29623);
nor UO_477 (O_477,N_29121,N_29428);
and UO_478 (O_478,N_28995,N_28561);
and UO_479 (O_479,N_29148,N_29892);
nand UO_480 (O_480,N_29800,N_28563);
xor UO_481 (O_481,N_29068,N_29274);
or UO_482 (O_482,N_29844,N_28778);
nor UO_483 (O_483,N_29329,N_29700);
nand UO_484 (O_484,N_29266,N_29841);
nor UO_485 (O_485,N_29340,N_29381);
nand UO_486 (O_486,N_29452,N_29050);
and UO_487 (O_487,N_29230,N_29884);
nand UO_488 (O_488,N_28930,N_29493);
xnor UO_489 (O_489,N_28690,N_28606);
nor UO_490 (O_490,N_29483,N_29000);
or UO_491 (O_491,N_29245,N_29615);
nand UO_492 (O_492,N_29369,N_29651);
xnor UO_493 (O_493,N_29655,N_29338);
or UO_494 (O_494,N_29946,N_28518);
or UO_495 (O_495,N_29144,N_29128);
and UO_496 (O_496,N_28803,N_28811);
nor UO_497 (O_497,N_29074,N_28550);
or UO_498 (O_498,N_29489,N_29083);
and UO_499 (O_499,N_29676,N_28820);
xor UO_500 (O_500,N_29759,N_29687);
xnor UO_501 (O_501,N_28821,N_29306);
nand UO_502 (O_502,N_29571,N_28539);
nand UO_503 (O_503,N_28944,N_28636);
and UO_504 (O_504,N_29327,N_29383);
nand UO_505 (O_505,N_28507,N_29132);
xnor UO_506 (O_506,N_28964,N_29040);
xor UO_507 (O_507,N_29756,N_29929);
nand UO_508 (O_508,N_28919,N_28738);
nand UO_509 (O_509,N_29173,N_29798);
or UO_510 (O_510,N_29409,N_29627);
and UO_511 (O_511,N_29116,N_28809);
nor UO_512 (O_512,N_29574,N_29323);
and UO_513 (O_513,N_28909,N_29578);
nand UO_514 (O_514,N_28910,N_29666);
nor UO_515 (O_515,N_29035,N_29475);
nand UO_516 (O_516,N_29472,N_28746);
xor UO_517 (O_517,N_28841,N_29869);
or UO_518 (O_518,N_29601,N_29435);
nor UO_519 (O_519,N_29406,N_28672);
and UO_520 (O_520,N_28805,N_29146);
nor UO_521 (O_521,N_29260,N_29464);
nor UO_522 (O_522,N_29373,N_28862);
xnor UO_523 (O_523,N_29480,N_28959);
xor UO_524 (O_524,N_29001,N_29679);
or UO_525 (O_525,N_29341,N_28998);
or UO_526 (O_526,N_28834,N_29165);
nor UO_527 (O_527,N_28752,N_29552);
nand UO_528 (O_528,N_29563,N_29152);
nand UO_529 (O_529,N_28984,N_28732);
and UO_530 (O_530,N_29181,N_29788);
and UO_531 (O_531,N_28795,N_28731);
nand UO_532 (O_532,N_29008,N_29943);
nand UO_533 (O_533,N_28590,N_29815);
xor UO_534 (O_534,N_29545,N_29521);
and UO_535 (O_535,N_29478,N_29042);
nand UO_536 (O_536,N_28666,N_29757);
xor UO_537 (O_537,N_28937,N_28798);
or UO_538 (O_538,N_28711,N_28514);
nor UO_539 (O_539,N_29893,N_29255);
nor UO_540 (O_540,N_28836,N_28612);
xor UO_541 (O_541,N_29762,N_29211);
nand UO_542 (O_542,N_28541,N_29813);
xor UO_543 (O_543,N_29485,N_29930);
nand UO_544 (O_544,N_29823,N_29147);
or UO_545 (O_545,N_29745,N_28888);
nor UO_546 (O_546,N_29599,N_28639);
or UO_547 (O_547,N_29120,N_28972);
or UO_548 (O_548,N_29292,N_28627);
xnor UO_549 (O_549,N_28945,N_29783);
or UO_550 (O_550,N_28765,N_28740);
or UO_551 (O_551,N_29904,N_29851);
nor UO_552 (O_552,N_29749,N_29316);
nand UO_553 (O_553,N_29223,N_29739);
nand UO_554 (O_554,N_29365,N_28645);
nand UO_555 (O_555,N_28766,N_29204);
and UO_556 (O_556,N_29647,N_28543);
and UO_557 (O_557,N_29536,N_29663);
and UO_558 (O_558,N_28789,N_29766);
or UO_559 (O_559,N_29980,N_28628);
nor UO_560 (O_560,N_28592,N_28629);
nand UO_561 (O_561,N_28884,N_29162);
and UO_562 (O_562,N_28837,N_28508);
or UO_563 (O_563,N_29859,N_29662);
or UO_564 (O_564,N_28572,N_29526);
nand UO_565 (O_565,N_29621,N_28736);
nand UO_566 (O_566,N_29978,N_29577);
nand UO_567 (O_567,N_29924,N_29874);
nor UO_568 (O_568,N_29486,N_29135);
or UO_569 (O_569,N_28743,N_29138);
and UO_570 (O_570,N_29041,N_29712);
nand UO_571 (O_571,N_29360,N_29714);
or UO_572 (O_572,N_29437,N_28952);
or UO_573 (O_573,N_29444,N_29385);
or UO_574 (O_574,N_28864,N_29529);
nor UO_575 (O_575,N_29752,N_29648);
nand UO_576 (O_576,N_29796,N_29718);
xor UO_577 (O_577,N_29959,N_29633);
xor UO_578 (O_578,N_29953,N_29387);
nor UO_579 (O_579,N_28881,N_29466);
nand UO_580 (O_580,N_29564,N_29061);
or UO_581 (O_581,N_29154,N_29344);
xor UO_582 (O_582,N_29699,N_28902);
and UO_583 (O_583,N_29733,N_29585);
nand UO_584 (O_584,N_29864,N_28576);
nor UO_585 (O_585,N_29293,N_29276);
and UO_586 (O_586,N_29006,N_28697);
or UO_587 (O_587,N_29994,N_29922);
nand UO_588 (O_588,N_28848,N_29534);
xnor UO_589 (O_589,N_29343,N_29215);
or UO_590 (O_590,N_28632,N_29236);
nor UO_591 (O_591,N_29451,N_29143);
xor UO_592 (O_592,N_29594,N_29983);
or UO_593 (O_593,N_29690,N_28729);
or UO_594 (O_594,N_29649,N_29631);
nand UO_595 (O_595,N_28640,N_28611);
nand UO_596 (O_596,N_29561,N_29938);
and UO_597 (O_597,N_29775,N_29760);
nand UO_598 (O_598,N_29597,N_29595);
xor UO_599 (O_599,N_29349,N_28528);
and UO_600 (O_600,N_29915,N_28817);
nand UO_601 (O_601,N_29295,N_28816);
xnor UO_602 (O_602,N_29157,N_29456);
xnor UO_603 (O_603,N_29857,N_29046);
or UO_604 (O_604,N_29289,N_29871);
nor UO_605 (O_605,N_28962,N_29541);
nand UO_606 (O_606,N_29535,N_28735);
nand UO_607 (O_607,N_29641,N_29020);
nor UO_608 (O_608,N_29433,N_29186);
nand UO_609 (O_609,N_28737,N_29065);
and UO_610 (O_610,N_29543,N_28688);
nor UO_611 (O_611,N_29944,N_28658);
nand UO_612 (O_612,N_28757,N_28947);
or UO_613 (O_613,N_29119,N_29208);
nor UO_614 (O_614,N_29636,N_28773);
nor UO_615 (O_615,N_29948,N_29321);
xor UO_616 (O_616,N_29384,N_29474);
xor UO_617 (O_617,N_28588,N_29415);
nand UO_618 (O_618,N_29955,N_28758);
xor UO_619 (O_619,N_29617,N_28882);
xnor UO_620 (O_620,N_29509,N_29530);
or UO_621 (O_621,N_29326,N_29918);
nor UO_622 (O_622,N_29418,N_28830);
nor UO_623 (O_623,N_29554,N_29112);
or UO_624 (O_624,N_28624,N_28790);
xor UO_625 (O_625,N_28785,N_28865);
or UO_626 (O_626,N_29028,N_29094);
or UO_627 (O_627,N_29078,N_29111);
or UO_628 (O_628,N_29440,N_28784);
xor UO_629 (O_629,N_28900,N_29053);
xor UO_630 (O_630,N_29751,N_28772);
nand UO_631 (O_631,N_29067,N_29596);
nand UO_632 (O_632,N_29294,N_29576);
xor UO_633 (O_633,N_29506,N_29720);
nand UO_634 (O_634,N_29875,N_29719);
xnor UO_635 (O_635,N_29105,N_29556);
nand UO_636 (O_636,N_29251,N_29459);
or UO_637 (O_637,N_29153,N_29867);
nor UO_638 (O_638,N_29411,N_29579);
or UO_639 (O_639,N_28905,N_29277);
and UO_640 (O_640,N_29682,N_29362);
xor UO_641 (O_641,N_28912,N_28839);
or UO_642 (O_642,N_29386,N_28854);
xor UO_643 (O_643,N_29004,N_28874);
or UO_644 (O_644,N_29999,N_29782);
xor UO_645 (O_645,N_28667,N_29591);
or UO_646 (O_646,N_29824,N_29034);
nor UO_647 (O_647,N_29598,N_29917);
nand UO_648 (O_648,N_29686,N_28574);
nor UO_649 (O_649,N_29833,N_29807);
nand UO_650 (O_650,N_29986,N_29213);
nor UO_651 (O_651,N_28571,N_28599);
nor UO_652 (O_652,N_29590,N_28958);
nand UO_653 (O_653,N_28564,N_29401);
and UO_654 (O_654,N_29495,N_29503);
nor UO_655 (O_655,N_29820,N_29443);
nand UO_656 (O_656,N_28660,N_29855);
xnor UO_657 (O_657,N_28577,N_29812);
and UO_658 (O_658,N_29583,N_29072);
nand UO_659 (O_659,N_29958,N_29581);
xnor UO_660 (O_660,N_29388,N_28646);
nor UO_661 (O_661,N_29127,N_28916);
xor UO_662 (O_662,N_28609,N_29310);
or UO_663 (O_663,N_29458,N_29625);
nor UO_664 (O_664,N_28770,N_28948);
and UO_665 (O_665,N_28675,N_29828);
nand UO_666 (O_666,N_28826,N_28622);
nand UO_667 (O_667,N_28876,N_29047);
nor UO_668 (O_668,N_29776,N_28828);
and UO_669 (O_669,N_29043,N_29711);
or UO_670 (O_670,N_29866,N_28651);
and UO_671 (O_671,N_28668,N_29052);
xnor UO_672 (O_672,N_29252,N_29896);
xnor UO_673 (O_673,N_28659,N_28664);
nor UO_674 (O_674,N_29469,N_28699);
or UO_675 (O_675,N_29092,N_28623);
and UO_676 (O_676,N_29747,N_29754);
xnor UO_677 (O_677,N_28520,N_29862);
nand UO_678 (O_678,N_29609,N_29737);
or UO_679 (O_679,N_28840,N_29975);
and UO_680 (O_680,N_29307,N_29665);
nand UO_681 (O_681,N_28847,N_29082);
nand UO_682 (O_682,N_28500,N_29519);
nor UO_683 (O_683,N_29079,N_29471);
or UO_684 (O_684,N_28997,N_29713);
xor UO_685 (O_685,N_29850,N_29019);
or UO_686 (O_686,N_29696,N_29018);
xnor UO_687 (O_687,N_28819,N_28906);
and UO_688 (O_688,N_29226,N_28955);
nand UO_689 (O_689,N_29171,N_28940);
nor UO_690 (O_690,N_28982,N_28717);
nor UO_691 (O_691,N_29133,N_28782);
xor UO_692 (O_692,N_29246,N_28635);
or UO_693 (O_693,N_28908,N_28783);
xor UO_694 (O_694,N_28966,N_28682);
nand UO_695 (O_695,N_29797,N_29176);
nand UO_696 (O_696,N_29927,N_29084);
nor UO_697 (O_697,N_29359,N_29650);
or UO_698 (O_698,N_29334,N_29109);
or UO_699 (O_699,N_28892,N_28519);
or UO_700 (O_700,N_28990,N_28710);
nor UO_701 (O_701,N_28907,N_29656);
nand UO_702 (O_702,N_29205,N_29090);
nor UO_703 (O_703,N_28875,N_29455);
and UO_704 (O_704,N_28894,N_29694);
nor UO_705 (O_705,N_28761,N_28866);
nand UO_706 (O_706,N_29382,N_28764);
and UO_707 (O_707,N_28642,N_29342);
nand UO_708 (O_708,N_28542,N_28551);
and UO_709 (O_709,N_29012,N_28698);
xnor UO_710 (O_710,N_29779,N_29099);
or UO_711 (O_711,N_28653,N_28626);
or UO_712 (O_712,N_29320,N_28808);
and UO_713 (O_713,N_28687,N_29971);
and UO_714 (O_714,N_29861,N_29077);
nand UO_715 (O_715,N_29549,N_28683);
nor UO_716 (O_716,N_28963,N_28973);
nand UO_717 (O_717,N_29960,N_29038);
xor UO_718 (O_718,N_28968,N_28853);
or UO_719 (O_719,N_29610,N_29097);
and UO_720 (O_720,N_28755,N_29070);
and UO_721 (O_721,N_29635,N_28517);
nor UO_722 (O_722,N_28634,N_28870);
nand UO_723 (O_723,N_29786,N_29335);
or UO_724 (O_724,N_29793,N_29473);
and UO_725 (O_725,N_28581,N_28921);
nand UO_726 (O_726,N_28505,N_29407);
nor UO_727 (O_727,N_29817,N_29883);
xor UO_728 (O_728,N_29730,N_29265);
and UO_729 (O_729,N_29025,N_28946);
xor UO_730 (O_730,N_28986,N_28994);
or UO_731 (O_731,N_29608,N_28583);
xnor UO_732 (O_732,N_28677,N_29972);
nor UO_733 (O_733,N_29377,N_29778);
nand UO_734 (O_734,N_28673,N_28558);
nor UO_735 (O_735,N_29619,N_28670);
xnor UO_736 (O_736,N_28691,N_29431);
nand UO_737 (O_737,N_29846,N_29692);
and UO_738 (O_738,N_29048,N_29468);
xnor UO_739 (O_739,N_29348,N_29196);
nand UO_740 (O_740,N_28568,N_29847);
xor UO_741 (O_741,N_29602,N_28887);
nand UO_742 (O_742,N_29729,N_29698);
xnor UO_743 (O_743,N_29979,N_29512);
nand UO_744 (O_744,N_29076,N_28608);
xor UO_745 (O_745,N_28552,N_29403);
or UO_746 (O_746,N_29027,N_28967);
and UO_747 (O_747,N_29494,N_29185);
nor UO_748 (O_748,N_29868,N_28681);
or UO_749 (O_749,N_28831,N_29392);
and UO_750 (O_750,N_28809,N_28835);
nor UO_751 (O_751,N_29304,N_28512);
or UO_752 (O_752,N_28728,N_29591);
xnor UO_753 (O_753,N_29674,N_28872);
nand UO_754 (O_754,N_28684,N_28580);
and UO_755 (O_755,N_28645,N_29014);
nand UO_756 (O_756,N_29088,N_29825);
or UO_757 (O_757,N_28933,N_28574);
or UO_758 (O_758,N_29887,N_29672);
and UO_759 (O_759,N_29008,N_28531);
or UO_760 (O_760,N_28582,N_28651);
xnor UO_761 (O_761,N_29575,N_29227);
nor UO_762 (O_762,N_29023,N_29737);
nor UO_763 (O_763,N_29777,N_28509);
nand UO_764 (O_764,N_29344,N_28931);
nand UO_765 (O_765,N_29782,N_29812);
and UO_766 (O_766,N_29663,N_28985);
nor UO_767 (O_767,N_29457,N_29456);
nand UO_768 (O_768,N_29792,N_28948);
or UO_769 (O_769,N_29997,N_29025);
nand UO_770 (O_770,N_29667,N_28557);
or UO_771 (O_771,N_29749,N_29149);
xnor UO_772 (O_772,N_29426,N_29561);
or UO_773 (O_773,N_28928,N_29319);
or UO_774 (O_774,N_29073,N_29880);
nand UO_775 (O_775,N_28883,N_28771);
nor UO_776 (O_776,N_29338,N_28907);
or UO_777 (O_777,N_29244,N_29549);
nand UO_778 (O_778,N_29364,N_28637);
xnor UO_779 (O_779,N_29096,N_28887);
xor UO_780 (O_780,N_29722,N_28917);
nand UO_781 (O_781,N_29017,N_29745);
or UO_782 (O_782,N_28897,N_28659);
and UO_783 (O_783,N_29640,N_29883);
nand UO_784 (O_784,N_29777,N_28625);
xor UO_785 (O_785,N_29516,N_29030);
and UO_786 (O_786,N_29453,N_29633);
nand UO_787 (O_787,N_28575,N_28923);
and UO_788 (O_788,N_29081,N_29712);
nand UO_789 (O_789,N_29657,N_29865);
or UO_790 (O_790,N_29361,N_29298);
xnor UO_791 (O_791,N_28511,N_28780);
xor UO_792 (O_792,N_28925,N_29959);
nand UO_793 (O_793,N_28920,N_28959);
and UO_794 (O_794,N_29020,N_28602);
or UO_795 (O_795,N_28646,N_28954);
nand UO_796 (O_796,N_29347,N_29550);
and UO_797 (O_797,N_28720,N_29057);
or UO_798 (O_798,N_29752,N_29944);
nor UO_799 (O_799,N_28931,N_28556);
nor UO_800 (O_800,N_29763,N_29195);
nand UO_801 (O_801,N_28939,N_29166);
or UO_802 (O_802,N_29434,N_29773);
xor UO_803 (O_803,N_29234,N_29928);
or UO_804 (O_804,N_29117,N_28789);
and UO_805 (O_805,N_28696,N_28689);
nor UO_806 (O_806,N_28696,N_28682);
nand UO_807 (O_807,N_28565,N_29289);
nand UO_808 (O_808,N_29153,N_29311);
or UO_809 (O_809,N_29331,N_28507);
and UO_810 (O_810,N_29190,N_29638);
or UO_811 (O_811,N_29892,N_29618);
and UO_812 (O_812,N_29298,N_28819);
and UO_813 (O_813,N_28739,N_28727);
or UO_814 (O_814,N_29115,N_28640);
nand UO_815 (O_815,N_29929,N_28522);
xnor UO_816 (O_816,N_29894,N_28714);
or UO_817 (O_817,N_29496,N_29383);
and UO_818 (O_818,N_29894,N_29332);
and UO_819 (O_819,N_29705,N_29497);
nor UO_820 (O_820,N_29745,N_29630);
xor UO_821 (O_821,N_29001,N_29476);
or UO_822 (O_822,N_29305,N_29278);
nand UO_823 (O_823,N_29260,N_29291);
nand UO_824 (O_824,N_29167,N_29211);
and UO_825 (O_825,N_29579,N_29099);
and UO_826 (O_826,N_28753,N_29408);
or UO_827 (O_827,N_29313,N_29216);
and UO_828 (O_828,N_28639,N_29444);
and UO_829 (O_829,N_28598,N_28615);
xnor UO_830 (O_830,N_28658,N_29847);
xor UO_831 (O_831,N_29964,N_29008);
nor UO_832 (O_832,N_29651,N_28827);
or UO_833 (O_833,N_29995,N_29892);
nor UO_834 (O_834,N_29595,N_28867);
nand UO_835 (O_835,N_29902,N_28632);
nor UO_836 (O_836,N_29228,N_29473);
or UO_837 (O_837,N_29075,N_29508);
or UO_838 (O_838,N_29611,N_28898);
xnor UO_839 (O_839,N_29786,N_28805);
and UO_840 (O_840,N_29382,N_29317);
xor UO_841 (O_841,N_29064,N_29964);
and UO_842 (O_842,N_28540,N_29980);
nand UO_843 (O_843,N_28555,N_29131);
nor UO_844 (O_844,N_29846,N_28584);
nor UO_845 (O_845,N_29377,N_29949);
xnor UO_846 (O_846,N_29974,N_29936);
xor UO_847 (O_847,N_28681,N_29503);
nand UO_848 (O_848,N_29766,N_29525);
or UO_849 (O_849,N_28867,N_29908);
and UO_850 (O_850,N_29391,N_29771);
nand UO_851 (O_851,N_29367,N_28642);
xnor UO_852 (O_852,N_29335,N_29337);
xnor UO_853 (O_853,N_28952,N_29984);
nand UO_854 (O_854,N_28649,N_29934);
nand UO_855 (O_855,N_29034,N_29569);
xnor UO_856 (O_856,N_29276,N_29911);
xor UO_857 (O_857,N_28907,N_28642);
or UO_858 (O_858,N_29993,N_28817);
nand UO_859 (O_859,N_28961,N_29623);
or UO_860 (O_860,N_29366,N_29929);
nor UO_861 (O_861,N_28616,N_28631);
and UO_862 (O_862,N_29993,N_29754);
and UO_863 (O_863,N_29827,N_29482);
and UO_864 (O_864,N_28518,N_29318);
and UO_865 (O_865,N_28506,N_28720);
xor UO_866 (O_866,N_29007,N_29718);
nand UO_867 (O_867,N_28955,N_28985);
nor UO_868 (O_868,N_28878,N_28720);
nor UO_869 (O_869,N_29103,N_29053);
xnor UO_870 (O_870,N_29613,N_29851);
nand UO_871 (O_871,N_28631,N_28847);
xor UO_872 (O_872,N_29146,N_29078);
nor UO_873 (O_873,N_29938,N_29121);
and UO_874 (O_874,N_29050,N_28860);
xor UO_875 (O_875,N_29103,N_29855);
and UO_876 (O_876,N_28825,N_28693);
or UO_877 (O_877,N_29091,N_29548);
or UO_878 (O_878,N_29949,N_28565);
xor UO_879 (O_879,N_29304,N_29437);
nand UO_880 (O_880,N_29961,N_29936);
xor UO_881 (O_881,N_29016,N_29870);
xnor UO_882 (O_882,N_29278,N_28754);
or UO_883 (O_883,N_29231,N_28984);
or UO_884 (O_884,N_29027,N_28858);
xor UO_885 (O_885,N_29087,N_29329);
or UO_886 (O_886,N_29216,N_29809);
or UO_887 (O_887,N_28788,N_29230);
nand UO_888 (O_888,N_28932,N_29682);
or UO_889 (O_889,N_29267,N_28731);
nand UO_890 (O_890,N_28687,N_29154);
xor UO_891 (O_891,N_28969,N_29999);
and UO_892 (O_892,N_28724,N_29630);
or UO_893 (O_893,N_29937,N_28808);
nand UO_894 (O_894,N_29005,N_29123);
and UO_895 (O_895,N_29479,N_29339);
xnor UO_896 (O_896,N_29549,N_28610);
and UO_897 (O_897,N_28874,N_29964);
nand UO_898 (O_898,N_28616,N_29625);
nand UO_899 (O_899,N_29136,N_28626);
nor UO_900 (O_900,N_29856,N_29673);
nor UO_901 (O_901,N_28677,N_29637);
nand UO_902 (O_902,N_28968,N_29019);
nor UO_903 (O_903,N_29142,N_29780);
and UO_904 (O_904,N_29770,N_29211);
or UO_905 (O_905,N_29257,N_29391);
and UO_906 (O_906,N_28832,N_29331);
nand UO_907 (O_907,N_29829,N_29473);
nor UO_908 (O_908,N_29987,N_28641);
or UO_909 (O_909,N_28841,N_29822);
xor UO_910 (O_910,N_28535,N_29851);
or UO_911 (O_911,N_29076,N_29195);
nor UO_912 (O_912,N_29345,N_29726);
or UO_913 (O_913,N_29589,N_28738);
or UO_914 (O_914,N_29867,N_28766);
xnor UO_915 (O_915,N_28799,N_29288);
nand UO_916 (O_916,N_29358,N_28734);
or UO_917 (O_917,N_29122,N_29962);
and UO_918 (O_918,N_28826,N_28901);
and UO_919 (O_919,N_28865,N_29497);
xor UO_920 (O_920,N_28688,N_29207);
nor UO_921 (O_921,N_29616,N_28583);
or UO_922 (O_922,N_28687,N_29457);
and UO_923 (O_923,N_28869,N_29133);
or UO_924 (O_924,N_28905,N_29616);
nor UO_925 (O_925,N_28953,N_28680);
nor UO_926 (O_926,N_28582,N_29983);
nor UO_927 (O_927,N_29708,N_29495);
nand UO_928 (O_928,N_29914,N_28866);
nor UO_929 (O_929,N_29739,N_29838);
and UO_930 (O_930,N_29322,N_28790);
xor UO_931 (O_931,N_29760,N_28770);
or UO_932 (O_932,N_29182,N_29098);
or UO_933 (O_933,N_28992,N_29410);
nor UO_934 (O_934,N_28605,N_29924);
nand UO_935 (O_935,N_28779,N_29919);
or UO_936 (O_936,N_28543,N_29189);
and UO_937 (O_937,N_28730,N_28943);
nand UO_938 (O_938,N_29104,N_28796);
or UO_939 (O_939,N_28705,N_29318);
xor UO_940 (O_940,N_29493,N_28795);
nor UO_941 (O_941,N_28615,N_28681);
and UO_942 (O_942,N_28794,N_28942);
and UO_943 (O_943,N_29870,N_29596);
nand UO_944 (O_944,N_28703,N_28754);
and UO_945 (O_945,N_28954,N_29096);
xnor UO_946 (O_946,N_29914,N_28965);
nand UO_947 (O_947,N_28699,N_29716);
nor UO_948 (O_948,N_29704,N_28829);
and UO_949 (O_949,N_29401,N_29954);
nor UO_950 (O_950,N_29978,N_29293);
or UO_951 (O_951,N_29296,N_29846);
nand UO_952 (O_952,N_29040,N_29302);
nor UO_953 (O_953,N_29877,N_29688);
nand UO_954 (O_954,N_28518,N_28893);
nand UO_955 (O_955,N_28984,N_28760);
xnor UO_956 (O_956,N_29559,N_28579);
and UO_957 (O_957,N_28689,N_29677);
nor UO_958 (O_958,N_29914,N_29100);
xnor UO_959 (O_959,N_29375,N_28723);
and UO_960 (O_960,N_29366,N_28919);
and UO_961 (O_961,N_29964,N_29053);
or UO_962 (O_962,N_28544,N_29468);
nand UO_963 (O_963,N_29647,N_29390);
nor UO_964 (O_964,N_28830,N_29782);
xor UO_965 (O_965,N_29156,N_29055);
nand UO_966 (O_966,N_28510,N_29407);
xnor UO_967 (O_967,N_29524,N_29471);
nor UO_968 (O_968,N_29845,N_29919);
and UO_969 (O_969,N_28971,N_29048);
nand UO_970 (O_970,N_29525,N_29826);
nor UO_971 (O_971,N_29472,N_28503);
nand UO_972 (O_972,N_28661,N_28765);
xnor UO_973 (O_973,N_28738,N_28928);
nor UO_974 (O_974,N_29572,N_29586);
nand UO_975 (O_975,N_28645,N_29358);
nand UO_976 (O_976,N_29824,N_29784);
nand UO_977 (O_977,N_29903,N_29342);
and UO_978 (O_978,N_29999,N_29589);
xor UO_979 (O_979,N_28749,N_28567);
and UO_980 (O_980,N_29037,N_28725);
and UO_981 (O_981,N_29051,N_29110);
and UO_982 (O_982,N_29809,N_28978);
xnor UO_983 (O_983,N_29663,N_29669);
nand UO_984 (O_984,N_29439,N_29097);
nand UO_985 (O_985,N_29781,N_28906);
xnor UO_986 (O_986,N_28780,N_29639);
nor UO_987 (O_987,N_29832,N_29856);
nand UO_988 (O_988,N_28506,N_29380);
and UO_989 (O_989,N_28644,N_29949);
or UO_990 (O_990,N_29635,N_29598);
nand UO_991 (O_991,N_29876,N_28767);
nor UO_992 (O_992,N_29239,N_28790);
and UO_993 (O_993,N_29773,N_29827);
and UO_994 (O_994,N_29943,N_29513);
xor UO_995 (O_995,N_29966,N_29676);
and UO_996 (O_996,N_29142,N_29363);
nor UO_997 (O_997,N_28776,N_29576);
or UO_998 (O_998,N_29070,N_28626);
and UO_999 (O_999,N_29534,N_29195);
xnor UO_1000 (O_1000,N_29230,N_29265);
nor UO_1001 (O_1001,N_29437,N_29620);
or UO_1002 (O_1002,N_28729,N_29532);
nor UO_1003 (O_1003,N_29436,N_29723);
xnor UO_1004 (O_1004,N_28792,N_29815);
and UO_1005 (O_1005,N_29296,N_28800);
or UO_1006 (O_1006,N_28936,N_28994);
nor UO_1007 (O_1007,N_28746,N_28839);
nand UO_1008 (O_1008,N_29637,N_29029);
and UO_1009 (O_1009,N_29720,N_29696);
or UO_1010 (O_1010,N_29413,N_29707);
xor UO_1011 (O_1011,N_29180,N_28531);
xnor UO_1012 (O_1012,N_29074,N_28894);
nor UO_1013 (O_1013,N_28845,N_29839);
and UO_1014 (O_1014,N_29059,N_28603);
nand UO_1015 (O_1015,N_28695,N_29345);
nor UO_1016 (O_1016,N_29412,N_29303);
nand UO_1017 (O_1017,N_29557,N_29738);
nor UO_1018 (O_1018,N_29253,N_28737);
xor UO_1019 (O_1019,N_28940,N_28654);
nor UO_1020 (O_1020,N_29257,N_28522);
xor UO_1021 (O_1021,N_28721,N_29973);
xnor UO_1022 (O_1022,N_28781,N_29181);
or UO_1023 (O_1023,N_28680,N_29877);
or UO_1024 (O_1024,N_29417,N_28771);
nand UO_1025 (O_1025,N_28765,N_29369);
nor UO_1026 (O_1026,N_29242,N_29504);
or UO_1027 (O_1027,N_29519,N_28924);
or UO_1028 (O_1028,N_29698,N_29645);
nand UO_1029 (O_1029,N_29657,N_28879);
or UO_1030 (O_1030,N_28616,N_29849);
and UO_1031 (O_1031,N_29102,N_28853);
nand UO_1032 (O_1032,N_29316,N_28958);
xnor UO_1033 (O_1033,N_28790,N_29069);
nor UO_1034 (O_1034,N_29949,N_29533);
xnor UO_1035 (O_1035,N_28984,N_29578);
or UO_1036 (O_1036,N_28568,N_29725);
or UO_1037 (O_1037,N_29908,N_29337);
nor UO_1038 (O_1038,N_28653,N_29011);
and UO_1039 (O_1039,N_28978,N_28613);
xnor UO_1040 (O_1040,N_29542,N_29546);
nand UO_1041 (O_1041,N_28550,N_29646);
or UO_1042 (O_1042,N_28662,N_29508);
and UO_1043 (O_1043,N_28771,N_29244);
xor UO_1044 (O_1044,N_29556,N_29733);
xnor UO_1045 (O_1045,N_28790,N_29475);
and UO_1046 (O_1046,N_28999,N_29608);
xor UO_1047 (O_1047,N_28581,N_28687);
or UO_1048 (O_1048,N_28743,N_29724);
or UO_1049 (O_1049,N_28628,N_28880);
nand UO_1050 (O_1050,N_29351,N_29476);
xnor UO_1051 (O_1051,N_28755,N_29974);
or UO_1052 (O_1052,N_28882,N_29178);
or UO_1053 (O_1053,N_28715,N_29141);
and UO_1054 (O_1054,N_29176,N_28577);
nor UO_1055 (O_1055,N_29228,N_29538);
and UO_1056 (O_1056,N_29042,N_29455);
xor UO_1057 (O_1057,N_28773,N_29994);
nor UO_1058 (O_1058,N_29162,N_29166);
nor UO_1059 (O_1059,N_28717,N_28797);
xor UO_1060 (O_1060,N_29042,N_29972);
nor UO_1061 (O_1061,N_29535,N_29372);
nor UO_1062 (O_1062,N_29195,N_28907);
or UO_1063 (O_1063,N_28623,N_28607);
or UO_1064 (O_1064,N_28736,N_28854);
xnor UO_1065 (O_1065,N_28923,N_28549);
nor UO_1066 (O_1066,N_28935,N_29310);
and UO_1067 (O_1067,N_29284,N_28862);
and UO_1068 (O_1068,N_28665,N_28686);
or UO_1069 (O_1069,N_29290,N_29252);
and UO_1070 (O_1070,N_29149,N_29028);
nor UO_1071 (O_1071,N_28806,N_29754);
or UO_1072 (O_1072,N_29952,N_29644);
xor UO_1073 (O_1073,N_29506,N_28674);
and UO_1074 (O_1074,N_28772,N_29373);
xor UO_1075 (O_1075,N_29917,N_28687);
nand UO_1076 (O_1076,N_29286,N_29544);
and UO_1077 (O_1077,N_29713,N_29047);
nor UO_1078 (O_1078,N_28643,N_29215);
xor UO_1079 (O_1079,N_29866,N_28606);
xor UO_1080 (O_1080,N_29611,N_29990);
xor UO_1081 (O_1081,N_28666,N_28853);
xor UO_1082 (O_1082,N_29353,N_28818);
or UO_1083 (O_1083,N_28780,N_29536);
nand UO_1084 (O_1084,N_28614,N_28932);
nor UO_1085 (O_1085,N_29028,N_28675);
and UO_1086 (O_1086,N_29636,N_29318);
nor UO_1087 (O_1087,N_28999,N_29705);
nor UO_1088 (O_1088,N_29439,N_28565);
nor UO_1089 (O_1089,N_29044,N_29252);
nor UO_1090 (O_1090,N_28711,N_29080);
and UO_1091 (O_1091,N_29165,N_28782);
nand UO_1092 (O_1092,N_29121,N_29876);
nor UO_1093 (O_1093,N_29715,N_29850);
or UO_1094 (O_1094,N_29936,N_28667);
nor UO_1095 (O_1095,N_28527,N_29838);
xor UO_1096 (O_1096,N_29768,N_29763);
nor UO_1097 (O_1097,N_28735,N_29816);
nand UO_1098 (O_1098,N_29378,N_29395);
and UO_1099 (O_1099,N_28848,N_29801);
nand UO_1100 (O_1100,N_29985,N_28547);
nand UO_1101 (O_1101,N_29391,N_29304);
and UO_1102 (O_1102,N_29446,N_28908);
nand UO_1103 (O_1103,N_29154,N_29538);
xnor UO_1104 (O_1104,N_29787,N_29130);
or UO_1105 (O_1105,N_29721,N_29893);
nand UO_1106 (O_1106,N_28878,N_29727);
or UO_1107 (O_1107,N_29955,N_29764);
and UO_1108 (O_1108,N_29404,N_28607);
xnor UO_1109 (O_1109,N_29228,N_29210);
or UO_1110 (O_1110,N_29561,N_29308);
and UO_1111 (O_1111,N_29036,N_29854);
xor UO_1112 (O_1112,N_29628,N_29655);
or UO_1113 (O_1113,N_29045,N_28698);
or UO_1114 (O_1114,N_28978,N_29419);
and UO_1115 (O_1115,N_29579,N_29927);
nand UO_1116 (O_1116,N_29386,N_29437);
xor UO_1117 (O_1117,N_28619,N_29057);
nand UO_1118 (O_1118,N_29376,N_28781);
and UO_1119 (O_1119,N_28507,N_29976);
or UO_1120 (O_1120,N_29015,N_28955);
and UO_1121 (O_1121,N_29764,N_28761);
xor UO_1122 (O_1122,N_29362,N_29687);
nand UO_1123 (O_1123,N_28703,N_28925);
xor UO_1124 (O_1124,N_29202,N_28930);
or UO_1125 (O_1125,N_29543,N_29241);
nor UO_1126 (O_1126,N_28617,N_28975);
nand UO_1127 (O_1127,N_29258,N_28763);
and UO_1128 (O_1128,N_28539,N_28639);
and UO_1129 (O_1129,N_28664,N_29118);
and UO_1130 (O_1130,N_28692,N_28881);
nand UO_1131 (O_1131,N_29263,N_29189);
nor UO_1132 (O_1132,N_28963,N_29946);
or UO_1133 (O_1133,N_29223,N_29874);
nand UO_1134 (O_1134,N_29697,N_28762);
nand UO_1135 (O_1135,N_29561,N_29289);
xnor UO_1136 (O_1136,N_29605,N_29565);
nand UO_1137 (O_1137,N_29760,N_29747);
and UO_1138 (O_1138,N_29195,N_29034);
nand UO_1139 (O_1139,N_29967,N_29771);
nor UO_1140 (O_1140,N_29735,N_29908);
and UO_1141 (O_1141,N_29440,N_28968);
nand UO_1142 (O_1142,N_29361,N_29141);
and UO_1143 (O_1143,N_29907,N_29226);
nand UO_1144 (O_1144,N_29697,N_29315);
nor UO_1145 (O_1145,N_28937,N_28721);
nand UO_1146 (O_1146,N_29781,N_29368);
xor UO_1147 (O_1147,N_29069,N_28793);
nor UO_1148 (O_1148,N_29510,N_29877);
xnor UO_1149 (O_1149,N_28636,N_29559);
xnor UO_1150 (O_1150,N_29789,N_29139);
or UO_1151 (O_1151,N_29036,N_29263);
or UO_1152 (O_1152,N_29348,N_29801);
nor UO_1153 (O_1153,N_29921,N_29048);
or UO_1154 (O_1154,N_28518,N_29324);
nand UO_1155 (O_1155,N_29675,N_29574);
and UO_1156 (O_1156,N_28501,N_29275);
and UO_1157 (O_1157,N_29872,N_29922);
and UO_1158 (O_1158,N_29319,N_28640);
and UO_1159 (O_1159,N_29545,N_29322);
and UO_1160 (O_1160,N_28560,N_29787);
or UO_1161 (O_1161,N_29739,N_28756);
or UO_1162 (O_1162,N_28552,N_29888);
and UO_1163 (O_1163,N_29248,N_28638);
or UO_1164 (O_1164,N_29714,N_29412);
and UO_1165 (O_1165,N_28751,N_29132);
nand UO_1166 (O_1166,N_29686,N_28708);
and UO_1167 (O_1167,N_29625,N_29369);
xnor UO_1168 (O_1168,N_29158,N_29607);
nor UO_1169 (O_1169,N_29192,N_29669);
nand UO_1170 (O_1170,N_29348,N_29838);
nor UO_1171 (O_1171,N_29435,N_29923);
and UO_1172 (O_1172,N_29865,N_28822);
and UO_1173 (O_1173,N_28964,N_29378);
and UO_1174 (O_1174,N_28535,N_29068);
nor UO_1175 (O_1175,N_29283,N_29356);
nor UO_1176 (O_1176,N_29515,N_28948);
nand UO_1177 (O_1177,N_29436,N_28822);
or UO_1178 (O_1178,N_29712,N_29389);
and UO_1179 (O_1179,N_29310,N_28733);
or UO_1180 (O_1180,N_29567,N_29122);
nand UO_1181 (O_1181,N_28976,N_28742);
or UO_1182 (O_1182,N_29321,N_29736);
nand UO_1183 (O_1183,N_28804,N_29094);
xnor UO_1184 (O_1184,N_29898,N_29911);
or UO_1185 (O_1185,N_29679,N_29669);
nor UO_1186 (O_1186,N_29411,N_29873);
nand UO_1187 (O_1187,N_28995,N_29196);
or UO_1188 (O_1188,N_29474,N_28573);
xnor UO_1189 (O_1189,N_29743,N_29549);
nand UO_1190 (O_1190,N_29599,N_29819);
nor UO_1191 (O_1191,N_29902,N_29235);
nand UO_1192 (O_1192,N_29842,N_29297);
nor UO_1193 (O_1193,N_28814,N_29407);
or UO_1194 (O_1194,N_28691,N_29451);
nand UO_1195 (O_1195,N_29784,N_28879);
nand UO_1196 (O_1196,N_29279,N_29297);
nor UO_1197 (O_1197,N_28969,N_29954);
xnor UO_1198 (O_1198,N_28891,N_29962);
and UO_1199 (O_1199,N_28719,N_29641);
nor UO_1200 (O_1200,N_28696,N_29947);
xnor UO_1201 (O_1201,N_29584,N_29212);
nor UO_1202 (O_1202,N_29604,N_29764);
xor UO_1203 (O_1203,N_28613,N_28855);
nand UO_1204 (O_1204,N_29760,N_29039);
xor UO_1205 (O_1205,N_29468,N_29467);
nor UO_1206 (O_1206,N_28955,N_29363);
nand UO_1207 (O_1207,N_29976,N_28721);
or UO_1208 (O_1208,N_29282,N_29742);
xnor UO_1209 (O_1209,N_29609,N_29017);
or UO_1210 (O_1210,N_29041,N_29252);
xor UO_1211 (O_1211,N_28605,N_29832);
xnor UO_1212 (O_1212,N_29928,N_29902);
nand UO_1213 (O_1213,N_29079,N_28557);
nand UO_1214 (O_1214,N_28667,N_29754);
and UO_1215 (O_1215,N_28859,N_29419);
nand UO_1216 (O_1216,N_29997,N_29160);
and UO_1217 (O_1217,N_28512,N_29193);
or UO_1218 (O_1218,N_29947,N_28774);
or UO_1219 (O_1219,N_29431,N_29091);
nor UO_1220 (O_1220,N_29866,N_29568);
nor UO_1221 (O_1221,N_29637,N_28976);
nand UO_1222 (O_1222,N_28543,N_29421);
nand UO_1223 (O_1223,N_29869,N_29298);
or UO_1224 (O_1224,N_28972,N_29035);
and UO_1225 (O_1225,N_29718,N_28922);
and UO_1226 (O_1226,N_29808,N_28836);
and UO_1227 (O_1227,N_29072,N_29454);
nor UO_1228 (O_1228,N_29100,N_29541);
xnor UO_1229 (O_1229,N_29130,N_28582);
nand UO_1230 (O_1230,N_28527,N_28513);
xor UO_1231 (O_1231,N_28523,N_29567);
nor UO_1232 (O_1232,N_29798,N_29223);
and UO_1233 (O_1233,N_29323,N_28992);
and UO_1234 (O_1234,N_29243,N_29052);
nand UO_1235 (O_1235,N_29759,N_29160);
nor UO_1236 (O_1236,N_29587,N_29772);
or UO_1237 (O_1237,N_29934,N_28842);
and UO_1238 (O_1238,N_29759,N_29964);
xor UO_1239 (O_1239,N_28674,N_29910);
or UO_1240 (O_1240,N_29145,N_28578);
xnor UO_1241 (O_1241,N_29115,N_29264);
or UO_1242 (O_1242,N_28805,N_29060);
nor UO_1243 (O_1243,N_29044,N_29188);
xor UO_1244 (O_1244,N_28844,N_29840);
or UO_1245 (O_1245,N_29129,N_29439);
nor UO_1246 (O_1246,N_29748,N_28765);
and UO_1247 (O_1247,N_28532,N_29619);
nand UO_1248 (O_1248,N_29442,N_29766);
nand UO_1249 (O_1249,N_29109,N_28752);
or UO_1250 (O_1250,N_28776,N_29628);
and UO_1251 (O_1251,N_28550,N_29107);
nor UO_1252 (O_1252,N_29603,N_29590);
xnor UO_1253 (O_1253,N_28749,N_28646);
nand UO_1254 (O_1254,N_29056,N_29337);
or UO_1255 (O_1255,N_29306,N_28994);
nor UO_1256 (O_1256,N_29461,N_29177);
nand UO_1257 (O_1257,N_28858,N_29306);
nor UO_1258 (O_1258,N_29601,N_28596);
xnor UO_1259 (O_1259,N_29041,N_29580);
xnor UO_1260 (O_1260,N_29596,N_29748);
or UO_1261 (O_1261,N_28631,N_28638);
nor UO_1262 (O_1262,N_29936,N_29198);
or UO_1263 (O_1263,N_29858,N_29865);
nand UO_1264 (O_1264,N_29453,N_29410);
and UO_1265 (O_1265,N_29280,N_29897);
and UO_1266 (O_1266,N_28540,N_28662);
nand UO_1267 (O_1267,N_29540,N_29668);
nand UO_1268 (O_1268,N_29193,N_28783);
and UO_1269 (O_1269,N_29844,N_28522);
xor UO_1270 (O_1270,N_28975,N_29864);
nand UO_1271 (O_1271,N_29491,N_29962);
nand UO_1272 (O_1272,N_28748,N_29817);
nor UO_1273 (O_1273,N_29405,N_28691);
nor UO_1274 (O_1274,N_28962,N_28717);
or UO_1275 (O_1275,N_29097,N_29111);
nand UO_1276 (O_1276,N_28965,N_29014);
and UO_1277 (O_1277,N_29414,N_29232);
xnor UO_1278 (O_1278,N_28658,N_29111);
and UO_1279 (O_1279,N_29946,N_28896);
nor UO_1280 (O_1280,N_29047,N_29768);
nor UO_1281 (O_1281,N_29586,N_29905);
or UO_1282 (O_1282,N_28611,N_29318);
nand UO_1283 (O_1283,N_29645,N_28523);
and UO_1284 (O_1284,N_28674,N_29803);
xnor UO_1285 (O_1285,N_29332,N_28674);
xnor UO_1286 (O_1286,N_29491,N_29242);
xor UO_1287 (O_1287,N_28608,N_29235);
or UO_1288 (O_1288,N_28532,N_29806);
nor UO_1289 (O_1289,N_28866,N_29134);
xor UO_1290 (O_1290,N_29899,N_29382);
nand UO_1291 (O_1291,N_29457,N_29886);
or UO_1292 (O_1292,N_29255,N_29154);
xor UO_1293 (O_1293,N_28793,N_28978);
nor UO_1294 (O_1294,N_28637,N_28618);
nand UO_1295 (O_1295,N_28798,N_29806);
nand UO_1296 (O_1296,N_29193,N_29318);
or UO_1297 (O_1297,N_29250,N_28945);
or UO_1298 (O_1298,N_29309,N_29804);
nor UO_1299 (O_1299,N_29866,N_28785);
or UO_1300 (O_1300,N_29355,N_29930);
nand UO_1301 (O_1301,N_29262,N_29650);
nor UO_1302 (O_1302,N_28594,N_29416);
and UO_1303 (O_1303,N_28834,N_28802);
and UO_1304 (O_1304,N_28838,N_28721);
xor UO_1305 (O_1305,N_28917,N_29474);
xnor UO_1306 (O_1306,N_28831,N_28772);
and UO_1307 (O_1307,N_29509,N_28965);
nor UO_1308 (O_1308,N_28718,N_28821);
xor UO_1309 (O_1309,N_29710,N_28534);
nand UO_1310 (O_1310,N_29611,N_29663);
and UO_1311 (O_1311,N_29142,N_29913);
xor UO_1312 (O_1312,N_29244,N_28922);
nand UO_1313 (O_1313,N_29312,N_28533);
and UO_1314 (O_1314,N_29526,N_29545);
nor UO_1315 (O_1315,N_29871,N_28703);
xnor UO_1316 (O_1316,N_29283,N_28640);
nor UO_1317 (O_1317,N_29736,N_29770);
or UO_1318 (O_1318,N_29848,N_29088);
and UO_1319 (O_1319,N_28784,N_28615);
nand UO_1320 (O_1320,N_29647,N_29696);
or UO_1321 (O_1321,N_29107,N_29387);
nor UO_1322 (O_1322,N_28857,N_29955);
xnor UO_1323 (O_1323,N_28681,N_28900);
or UO_1324 (O_1324,N_28770,N_29364);
or UO_1325 (O_1325,N_29262,N_29969);
nand UO_1326 (O_1326,N_29096,N_29375);
and UO_1327 (O_1327,N_29628,N_29645);
xnor UO_1328 (O_1328,N_29085,N_29418);
nand UO_1329 (O_1329,N_29132,N_29738);
nand UO_1330 (O_1330,N_28800,N_29174);
xnor UO_1331 (O_1331,N_29801,N_29332);
xnor UO_1332 (O_1332,N_28962,N_28827);
xor UO_1333 (O_1333,N_29550,N_29559);
xor UO_1334 (O_1334,N_29249,N_28668);
or UO_1335 (O_1335,N_29755,N_28604);
xnor UO_1336 (O_1336,N_29587,N_29751);
nor UO_1337 (O_1337,N_29576,N_29316);
nand UO_1338 (O_1338,N_29331,N_28665);
and UO_1339 (O_1339,N_28649,N_29984);
or UO_1340 (O_1340,N_29514,N_29255);
or UO_1341 (O_1341,N_28925,N_29279);
and UO_1342 (O_1342,N_29361,N_29876);
or UO_1343 (O_1343,N_28686,N_29448);
or UO_1344 (O_1344,N_29331,N_28672);
and UO_1345 (O_1345,N_29661,N_29696);
xnor UO_1346 (O_1346,N_28615,N_29115);
or UO_1347 (O_1347,N_29994,N_29796);
nor UO_1348 (O_1348,N_29361,N_28907);
xor UO_1349 (O_1349,N_29385,N_29686);
and UO_1350 (O_1350,N_28927,N_29034);
nor UO_1351 (O_1351,N_29846,N_29606);
and UO_1352 (O_1352,N_28513,N_28602);
or UO_1353 (O_1353,N_29700,N_29090);
or UO_1354 (O_1354,N_28700,N_29912);
or UO_1355 (O_1355,N_28916,N_29943);
nand UO_1356 (O_1356,N_29483,N_28765);
or UO_1357 (O_1357,N_29168,N_28568);
or UO_1358 (O_1358,N_29766,N_29003);
and UO_1359 (O_1359,N_29985,N_29851);
and UO_1360 (O_1360,N_29389,N_28607);
nand UO_1361 (O_1361,N_29589,N_29569);
nand UO_1362 (O_1362,N_28665,N_29725);
or UO_1363 (O_1363,N_29603,N_28769);
xor UO_1364 (O_1364,N_29325,N_29948);
xor UO_1365 (O_1365,N_28628,N_29665);
nand UO_1366 (O_1366,N_28834,N_28993);
and UO_1367 (O_1367,N_29062,N_28687);
and UO_1368 (O_1368,N_29042,N_28725);
xnor UO_1369 (O_1369,N_29501,N_29906);
xor UO_1370 (O_1370,N_29382,N_29310);
nand UO_1371 (O_1371,N_28634,N_29871);
nand UO_1372 (O_1372,N_29157,N_28763);
nor UO_1373 (O_1373,N_29569,N_28906);
nor UO_1374 (O_1374,N_29520,N_29436);
nand UO_1375 (O_1375,N_29584,N_29717);
and UO_1376 (O_1376,N_29608,N_29296);
and UO_1377 (O_1377,N_29965,N_29687);
or UO_1378 (O_1378,N_29588,N_28710);
nand UO_1379 (O_1379,N_29921,N_28897);
or UO_1380 (O_1380,N_29173,N_29622);
and UO_1381 (O_1381,N_29926,N_29853);
nor UO_1382 (O_1382,N_28598,N_29831);
xor UO_1383 (O_1383,N_29021,N_28999);
nand UO_1384 (O_1384,N_29639,N_29251);
or UO_1385 (O_1385,N_28826,N_29422);
nor UO_1386 (O_1386,N_28929,N_28782);
nand UO_1387 (O_1387,N_29330,N_28519);
xor UO_1388 (O_1388,N_28878,N_29401);
nand UO_1389 (O_1389,N_29095,N_29671);
and UO_1390 (O_1390,N_29240,N_29396);
nor UO_1391 (O_1391,N_29452,N_28820);
xnor UO_1392 (O_1392,N_28998,N_28729);
and UO_1393 (O_1393,N_29529,N_29565);
nor UO_1394 (O_1394,N_29089,N_29356);
xor UO_1395 (O_1395,N_28517,N_28592);
nor UO_1396 (O_1396,N_29156,N_29816);
or UO_1397 (O_1397,N_28676,N_28529);
nor UO_1398 (O_1398,N_29802,N_28773);
nor UO_1399 (O_1399,N_28576,N_29729);
nand UO_1400 (O_1400,N_29994,N_28793);
nor UO_1401 (O_1401,N_29367,N_28744);
xnor UO_1402 (O_1402,N_29532,N_28857);
nand UO_1403 (O_1403,N_28773,N_29187);
or UO_1404 (O_1404,N_29957,N_29371);
nor UO_1405 (O_1405,N_29032,N_28686);
nand UO_1406 (O_1406,N_29480,N_29729);
or UO_1407 (O_1407,N_29307,N_29968);
nand UO_1408 (O_1408,N_28899,N_28901);
nand UO_1409 (O_1409,N_28510,N_28956);
nand UO_1410 (O_1410,N_28692,N_29919);
nor UO_1411 (O_1411,N_28875,N_29259);
or UO_1412 (O_1412,N_29517,N_29748);
or UO_1413 (O_1413,N_28813,N_28870);
nand UO_1414 (O_1414,N_28940,N_29766);
nand UO_1415 (O_1415,N_28678,N_29017);
or UO_1416 (O_1416,N_29526,N_29511);
or UO_1417 (O_1417,N_29054,N_28910);
nand UO_1418 (O_1418,N_28927,N_29901);
nor UO_1419 (O_1419,N_29094,N_28821);
xnor UO_1420 (O_1420,N_28564,N_29823);
xor UO_1421 (O_1421,N_29693,N_29420);
xnor UO_1422 (O_1422,N_28503,N_29836);
xor UO_1423 (O_1423,N_28802,N_29561);
or UO_1424 (O_1424,N_29091,N_29866);
and UO_1425 (O_1425,N_29420,N_28589);
nand UO_1426 (O_1426,N_29610,N_29159);
nor UO_1427 (O_1427,N_29080,N_29543);
xor UO_1428 (O_1428,N_29230,N_29269);
xor UO_1429 (O_1429,N_29149,N_29941);
or UO_1430 (O_1430,N_29882,N_29496);
or UO_1431 (O_1431,N_28847,N_28663);
nor UO_1432 (O_1432,N_29865,N_28717);
xor UO_1433 (O_1433,N_29642,N_29605);
and UO_1434 (O_1434,N_29956,N_29318);
and UO_1435 (O_1435,N_28583,N_29035);
nor UO_1436 (O_1436,N_29944,N_29789);
nand UO_1437 (O_1437,N_29579,N_28694);
or UO_1438 (O_1438,N_29076,N_28912);
nor UO_1439 (O_1439,N_29550,N_29875);
nand UO_1440 (O_1440,N_29694,N_28764);
xor UO_1441 (O_1441,N_29467,N_29210);
nor UO_1442 (O_1442,N_29168,N_29899);
nand UO_1443 (O_1443,N_29695,N_28811);
and UO_1444 (O_1444,N_29996,N_29063);
nor UO_1445 (O_1445,N_29173,N_28684);
xnor UO_1446 (O_1446,N_28997,N_29893);
nor UO_1447 (O_1447,N_28862,N_28657);
nand UO_1448 (O_1448,N_29536,N_29417);
nor UO_1449 (O_1449,N_29079,N_29825);
or UO_1450 (O_1450,N_29376,N_28542);
nand UO_1451 (O_1451,N_29146,N_29463);
nor UO_1452 (O_1452,N_28903,N_29289);
and UO_1453 (O_1453,N_28857,N_29244);
or UO_1454 (O_1454,N_29157,N_29782);
xnor UO_1455 (O_1455,N_29338,N_29099);
nor UO_1456 (O_1456,N_29720,N_29020);
xnor UO_1457 (O_1457,N_29020,N_28864);
nor UO_1458 (O_1458,N_28610,N_29510);
and UO_1459 (O_1459,N_29446,N_29906);
or UO_1460 (O_1460,N_29637,N_28592);
and UO_1461 (O_1461,N_29689,N_29093);
nand UO_1462 (O_1462,N_29036,N_28856);
nor UO_1463 (O_1463,N_29585,N_29239);
nor UO_1464 (O_1464,N_29685,N_29118);
or UO_1465 (O_1465,N_28898,N_29747);
or UO_1466 (O_1466,N_28820,N_29605);
and UO_1467 (O_1467,N_28782,N_28538);
nor UO_1468 (O_1468,N_29880,N_29242);
xor UO_1469 (O_1469,N_29723,N_29996);
nor UO_1470 (O_1470,N_28714,N_29619);
nand UO_1471 (O_1471,N_29411,N_28545);
and UO_1472 (O_1472,N_28834,N_29161);
nor UO_1473 (O_1473,N_28852,N_29881);
nor UO_1474 (O_1474,N_29497,N_29789);
xnor UO_1475 (O_1475,N_29154,N_29127);
or UO_1476 (O_1476,N_29316,N_29138);
or UO_1477 (O_1477,N_28544,N_28993);
or UO_1478 (O_1478,N_29192,N_29291);
and UO_1479 (O_1479,N_28897,N_29005);
xnor UO_1480 (O_1480,N_29368,N_29227);
xor UO_1481 (O_1481,N_29004,N_29769);
and UO_1482 (O_1482,N_28981,N_29328);
and UO_1483 (O_1483,N_29388,N_28757);
nor UO_1484 (O_1484,N_29710,N_28563);
xnor UO_1485 (O_1485,N_29730,N_29068);
xnor UO_1486 (O_1486,N_29312,N_28676);
or UO_1487 (O_1487,N_29429,N_29984);
xor UO_1488 (O_1488,N_28618,N_29317);
xor UO_1489 (O_1489,N_28583,N_28655);
nor UO_1490 (O_1490,N_28643,N_28525);
nor UO_1491 (O_1491,N_28967,N_28643);
and UO_1492 (O_1492,N_28607,N_28655);
or UO_1493 (O_1493,N_28805,N_28851);
and UO_1494 (O_1494,N_29609,N_29338);
or UO_1495 (O_1495,N_29402,N_29233);
xnor UO_1496 (O_1496,N_29078,N_28638);
or UO_1497 (O_1497,N_28500,N_28661);
nand UO_1498 (O_1498,N_28527,N_28645);
xnor UO_1499 (O_1499,N_29662,N_29434);
nor UO_1500 (O_1500,N_29311,N_29848);
nand UO_1501 (O_1501,N_28569,N_29131);
nand UO_1502 (O_1502,N_29910,N_28854);
xor UO_1503 (O_1503,N_29784,N_29523);
nand UO_1504 (O_1504,N_29038,N_29459);
and UO_1505 (O_1505,N_29799,N_28522);
or UO_1506 (O_1506,N_29238,N_29413);
xnor UO_1507 (O_1507,N_29396,N_29100);
or UO_1508 (O_1508,N_29619,N_28671);
nor UO_1509 (O_1509,N_29354,N_29697);
nand UO_1510 (O_1510,N_29104,N_29120);
and UO_1511 (O_1511,N_28994,N_29322);
or UO_1512 (O_1512,N_29886,N_28556);
or UO_1513 (O_1513,N_29805,N_28976);
nand UO_1514 (O_1514,N_28667,N_28770);
nor UO_1515 (O_1515,N_29146,N_28878);
nand UO_1516 (O_1516,N_29213,N_29373);
nor UO_1517 (O_1517,N_29837,N_28729);
nor UO_1518 (O_1518,N_28798,N_29918);
nand UO_1519 (O_1519,N_29557,N_29042);
and UO_1520 (O_1520,N_29466,N_29063);
xor UO_1521 (O_1521,N_28931,N_28836);
and UO_1522 (O_1522,N_29614,N_28590);
and UO_1523 (O_1523,N_29156,N_28969);
xnor UO_1524 (O_1524,N_29575,N_29501);
or UO_1525 (O_1525,N_29567,N_29566);
and UO_1526 (O_1526,N_29034,N_29891);
xor UO_1527 (O_1527,N_29928,N_28907);
nand UO_1528 (O_1528,N_29442,N_29794);
nand UO_1529 (O_1529,N_29123,N_29842);
nand UO_1530 (O_1530,N_28527,N_29685);
and UO_1531 (O_1531,N_28525,N_28601);
and UO_1532 (O_1532,N_29545,N_28511);
or UO_1533 (O_1533,N_29570,N_29144);
nand UO_1534 (O_1534,N_28903,N_29395);
or UO_1535 (O_1535,N_29728,N_29136);
nand UO_1536 (O_1536,N_28837,N_28733);
nor UO_1537 (O_1537,N_28975,N_29796);
nand UO_1538 (O_1538,N_28654,N_28800);
and UO_1539 (O_1539,N_29800,N_29856);
nor UO_1540 (O_1540,N_28958,N_28517);
nor UO_1541 (O_1541,N_28996,N_28723);
nand UO_1542 (O_1542,N_28552,N_28788);
nand UO_1543 (O_1543,N_28925,N_29740);
or UO_1544 (O_1544,N_29799,N_29045);
nand UO_1545 (O_1545,N_28807,N_29351);
and UO_1546 (O_1546,N_28790,N_29366);
nand UO_1547 (O_1547,N_29464,N_28990);
nand UO_1548 (O_1548,N_29347,N_28787);
and UO_1549 (O_1549,N_29715,N_29385);
xnor UO_1550 (O_1550,N_29050,N_29164);
nor UO_1551 (O_1551,N_28619,N_29322);
nor UO_1552 (O_1552,N_29558,N_29937);
nor UO_1553 (O_1553,N_29339,N_29865);
or UO_1554 (O_1554,N_28672,N_29433);
and UO_1555 (O_1555,N_29531,N_29054);
nand UO_1556 (O_1556,N_29862,N_28883);
or UO_1557 (O_1557,N_29082,N_29434);
xor UO_1558 (O_1558,N_29234,N_28887);
or UO_1559 (O_1559,N_28500,N_28788);
nand UO_1560 (O_1560,N_29691,N_29205);
nand UO_1561 (O_1561,N_29043,N_29533);
and UO_1562 (O_1562,N_28532,N_29111);
or UO_1563 (O_1563,N_29604,N_29233);
and UO_1564 (O_1564,N_29956,N_28579);
nor UO_1565 (O_1565,N_29157,N_28781);
nor UO_1566 (O_1566,N_28651,N_29583);
or UO_1567 (O_1567,N_29857,N_29548);
xor UO_1568 (O_1568,N_28690,N_28947);
or UO_1569 (O_1569,N_29747,N_29716);
nor UO_1570 (O_1570,N_28688,N_29009);
nand UO_1571 (O_1571,N_29417,N_28659);
and UO_1572 (O_1572,N_28864,N_28567);
and UO_1573 (O_1573,N_29404,N_28636);
or UO_1574 (O_1574,N_29451,N_28644);
nand UO_1575 (O_1575,N_28642,N_28551);
nand UO_1576 (O_1576,N_29778,N_28615);
and UO_1577 (O_1577,N_28555,N_28791);
or UO_1578 (O_1578,N_29542,N_29476);
xnor UO_1579 (O_1579,N_29596,N_29914);
or UO_1580 (O_1580,N_28598,N_29302);
xor UO_1581 (O_1581,N_29636,N_29537);
nor UO_1582 (O_1582,N_29915,N_28845);
or UO_1583 (O_1583,N_28913,N_29765);
or UO_1584 (O_1584,N_28579,N_29693);
nand UO_1585 (O_1585,N_28878,N_29829);
or UO_1586 (O_1586,N_28865,N_29125);
or UO_1587 (O_1587,N_29079,N_29775);
xnor UO_1588 (O_1588,N_29773,N_28880);
or UO_1589 (O_1589,N_29485,N_28695);
nor UO_1590 (O_1590,N_29839,N_29880);
and UO_1591 (O_1591,N_28628,N_29147);
xor UO_1592 (O_1592,N_29373,N_29796);
nand UO_1593 (O_1593,N_28631,N_29426);
and UO_1594 (O_1594,N_28928,N_29512);
nand UO_1595 (O_1595,N_29840,N_29130);
or UO_1596 (O_1596,N_28658,N_29493);
nor UO_1597 (O_1597,N_29702,N_29882);
and UO_1598 (O_1598,N_29469,N_28859);
nand UO_1599 (O_1599,N_29800,N_29882);
nor UO_1600 (O_1600,N_28746,N_29746);
nor UO_1601 (O_1601,N_28818,N_28665);
xnor UO_1602 (O_1602,N_29322,N_29963);
nor UO_1603 (O_1603,N_29258,N_29733);
and UO_1604 (O_1604,N_29273,N_29270);
xnor UO_1605 (O_1605,N_28884,N_29758);
nand UO_1606 (O_1606,N_29952,N_29463);
nor UO_1607 (O_1607,N_29481,N_29224);
and UO_1608 (O_1608,N_29552,N_28861);
or UO_1609 (O_1609,N_28703,N_28759);
and UO_1610 (O_1610,N_29475,N_29717);
and UO_1611 (O_1611,N_29748,N_29256);
or UO_1612 (O_1612,N_29356,N_29907);
xnor UO_1613 (O_1613,N_28511,N_28908);
nor UO_1614 (O_1614,N_29525,N_28947);
nor UO_1615 (O_1615,N_28653,N_28850);
or UO_1616 (O_1616,N_29962,N_28996);
nand UO_1617 (O_1617,N_28883,N_29207);
or UO_1618 (O_1618,N_29015,N_29360);
xor UO_1619 (O_1619,N_29704,N_28871);
nor UO_1620 (O_1620,N_29271,N_29762);
nand UO_1621 (O_1621,N_29669,N_28915);
nand UO_1622 (O_1622,N_29202,N_29285);
xor UO_1623 (O_1623,N_29099,N_29494);
nand UO_1624 (O_1624,N_28977,N_29264);
nand UO_1625 (O_1625,N_29357,N_29991);
and UO_1626 (O_1626,N_29378,N_29230);
nor UO_1627 (O_1627,N_29648,N_29330);
and UO_1628 (O_1628,N_29559,N_29979);
nor UO_1629 (O_1629,N_29653,N_29990);
xnor UO_1630 (O_1630,N_28687,N_29299);
nor UO_1631 (O_1631,N_28710,N_28838);
and UO_1632 (O_1632,N_29816,N_28566);
or UO_1633 (O_1633,N_29614,N_29442);
nor UO_1634 (O_1634,N_29748,N_29981);
nor UO_1635 (O_1635,N_28641,N_29429);
and UO_1636 (O_1636,N_29722,N_29171);
xor UO_1637 (O_1637,N_29653,N_29813);
xnor UO_1638 (O_1638,N_29560,N_29828);
nor UO_1639 (O_1639,N_28985,N_29605);
nor UO_1640 (O_1640,N_29792,N_28802);
nor UO_1641 (O_1641,N_29195,N_29733);
xor UO_1642 (O_1642,N_29251,N_29662);
xor UO_1643 (O_1643,N_29287,N_29378);
nor UO_1644 (O_1644,N_29744,N_29887);
nand UO_1645 (O_1645,N_29829,N_28511);
and UO_1646 (O_1646,N_29937,N_29586);
and UO_1647 (O_1647,N_28572,N_28718);
nor UO_1648 (O_1648,N_29750,N_29052);
and UO_1649 (O_1649,N_29698,N_29067);
nor UO_1650 (O_1650,N_29366,N_29025);
nor UO_1651 (O_1651,N_29942,N_28703);
nor UO_1652 (O_1652,N_29931,N_29021);
nor UO_1653 (O_1653,N_28552,N_29593);
nand UO_1654 (O_1654,N_28616,N_29292);
and UO_1655 (O_1655,N_28797,N_29948);
nor UO_1656 (O_1656,N_28627,N_28955);
xor UO_1657 (O_1657,N_28829,N_29620);
nor UO_1658 (O_1658,N_29253,N_29810);
and UO_1659 (O_1659,N_28993,N_28829);
xor UO_1660 (O_1660,N_29294,N_29225);
and UO_1661 (O_1661,N_28692,N_28667);
nand UO_1662 (O_1662,N_29702,N_29402);
nor UO_1663 (O_1663,N_28892,N_29652);
nor UO_1664 (O_1664,N_28848,N_29965);
nand UO_1665 (O_1665,N_29365,N_28531);
or UO_1666 (O_1666,N_29877,N_29126);
and UO_1667 (O_1667,N_28624,N_28919);
nand UO_1668 (O_1668,N_29392,N_28670);
or UO_1669 (O_1669,N_29290,N_29076);
and UO_1670 (O_1670,N_29530,N_29348);
or UO_1671 (O_1671,N_28956,N_29730);
nor UO_1672 (O_1672,N_29621,N_29836);
nor UO_1673 (O_1673,N_29637,N_29880);
nand UO_1674 (O_1674,N_29222,N_29597);
or UO_1675 (O_1675,N_29566,N_29187);
and UO_1676 (O_1676,N_29205,N_29498);
nand UO_1677 (O_1677,N_28762,N_28551);
or UO_1678 (O_1678,N_29069,N_29950);
or UO_1679 (O_1679,N_29494,N_28921);
nor UO_1680 (O_1680,N_29376,N_29897);
or UO_1681 (O_1681,N_28679,N_29861);
nand UO_1682 (O_1682,N_29920,N_28873);
nand UO_1683 (O_1683,N_29043,N_29336);
nand UO_1684 (O_1684,N_28697,N_28663);
xor UO_1685 (O_1685,N_29435,N_29072);
or UO_1686 (O_1686,N_29137,N_28860);
nand UO_1687 (O_1687,N_29201,N_28918);
xor UO_1688 (O_1688,N_28994,N_28908);
nor UO_1689 (O_1689,N_29631,N_28934);
or UO_1690 (O_1690,N_29189,N_28804);
and UO_1691 (O_1691,N_29562,N_29585);
or UO_1692 (O_1692,N_29624,N_28804);
nand UO_1693 (O_1693,N_29303,N_28908);
or UO_1694 (O_1694,N_28635,N_29638);
nand UO_1695 (O_1695,N_28820,N_29880);
or UO_1696 (O_1696,N_29056,N_29840);
nor UO_1697 (O_1697,N_28993,N_29279);
or UO_1698 (O_1698,N_28649,N_29164);
and UO_1699 (O_1699,N_29524,N_28648);
nor UO_1700 (O_1700,N_29539,N_28801);
nor UO_1701 (O_1701,N_29202,N_28919);
xnor UO_1702 (O_1702,N_28943,N_29681);
and UO_1703 (O_1703,N_29131,N_29852);
or UO_1704 (O_1704,N_29644,N_29316);
nand UO_1705 (O_1705,N_29004,N_29604);
or UO_1706 (O_1706,N_28678,N_28681);
nand UO_1707 (O_1707,N_28861,N_29751);
or UO_1708 (O_1708,N_28592,N_29548);
nand UO_1709 (O_1709,N_29850,N_28565);
nor UO_1710 (O_1710,N_29193,N_29771);
nor UO_1711 (O_1711,N_29598,N_28680);
nand UO_1712 (O_1712,N_28755,N_29625);
nor UO_1713 (O_1713,N_29492,N_28659);
and UO_1714 (O_1714,N_28683,N_29126);
and UO_1715 (O_1715,N_28666,N_29941);
xnor UO_1716 (O_1716,N_29119,N_29088);
and UO_1717 (O_1717,N_29866,N_28671);
and UO_1718 (O_1718,N_29555,N_29961);
xnor UO_1719 (O_1719,N_29897,N_28665);
and UO_1720 (O_1720,N_29724,N_28902);
nor UO_1721 (O_1721,N_29824,N_28962);
nor UO_1722 (O_1722,N_28987,N_28585);
or UO_1723 (O_1723,N_29342,N_29640);
nand UO_1724 (O_1724,N_29412,N_28598);
nor UO_1725 (O_1725,N_28927,N_28534);
nor UO_1726 (O_1726,N_28896,N_29692);
nor UO_1727 (O_1727,N_29619,N_29847);
xnor UO_1728 (O_1728,N_29975,N_28820);
xnor UO_1729 (O_1729,N_29515,N_29748);
nor UO_1730 (O_1730,N_29120,N_28804);
or UO_1731 (O_1731,N_29333,N_28847);
or UO_1732 (O_1732,N_29328,N_29235);
and UO_1733 (O_1733,N_28913,N_29794);
xnor UO_1734 (O_1734,N_28544,N_28689);
or UO_1735 (O_1735,N_29521,N_29978);
xor UO_1736 (O_1736,N_29460,N_29523);
and UO_1737 (O_1737,N_29017,N_29885);
xor UO_1738 (O_1738,N_28605,N_29440);
xnor UO_1739 (O_1739,N_29704,N_29467);
nand UO_1740 (O_1740,N_29428,N_29096);
nor UO_1741 (O_1741,N_29447,N_29180);
nor UO_1742 (O_1742,N_29028,N_29937);
nand UO_1743 (O_1743,N_28871,N_29636);
and UO_1744 (O_1744,N_28710,N_29935);
xor UO_1745 (O_1745,N_28745,N_28978);
nor UO_1746 (O_1746,N_28675,N_29495);
and UO_1747 (O_1747,N_28944,N_28691);
nor UO_1748 (O_1748,N_29232,N_29972);
nor UO_1749 (O_1749,N_29445,N_29868);
xor UO_1750 (O_1750,N_29130,N_29186);
nor UO_1751 (O_1751,N_29529,N_29967);
nand UO_1752 (O_1752,N_28738,N_28612);
or UO_1753 (O_1753,N_28611,N_29133);
or UO_1754 (O_1754,N_29617,N_28621);
nand UO_1755 (O_1755,N_28844,N_28528);
and UO_1756 (O_1756,N_28757,N_29809);
or UO_1757 (O_1757,N_29457,N_28721);
nand UO_1758 (O_1758,N_29614,N_29123);
xor UO_1759 (O_1759,N_28574,N_29119);
and UO_1760 (O_1760,N_29790,N_28813);
nor UO_1761 (O_1761,N_29963,N_29711);
and UO_1762 (O_1762,N_29750,N_29873);
xor UO_1763 (O_1763,N_29482,N_29225);
nand UO_1764 (O_1764,N_29694,N_28984);
xor UO_1765 (O_1765,N_29841,N_29676);
and UO_1766 (O_1766,N_29728,N_28890);
nor UO_1767 (O_1767,N_29868,N_28505);
xnor UO_1768 (O_1768,N_29605,N_28943);
or UO_1769 (O_1769,N_29346,N_29791);
nor UO_1770 (O_1770,N_28628,N_29326);
or UO_1771 (O_1771,N_28842,N_29788);
xnor UO_1772 (O_1772,N_28798,N_28513);
nor UO_1773 (O_1773,N_29703,N_28525);
nand UO_1774 (O_1774,N_29931,N_29682);
nand UO_1775 (O_1775,N_29775,N_28647);
nor UO_1776 (O_1776,N_29767,N_29447);
nand UO_1777 (O_1777,N_29337,N_29713);
and UO_1778 (O_1778,N_28846,N_28890);
nand UO_1779 (O_1779,N_28918,N_29379);
nand UO_1780 (O_1780,N_29727,N_29781);
nand UO_1781 (O_1781,N_29592,N_28709);
nand UO_1782 (O_1782,N_29890,N_29552);
and UO_1783 (O_1783,N_29620,N_29006);
nand UO_1784 (O_1784,N_29088,N_28808);
and UO_1785 (O_1785,N_28996,N_29464);
or UO_1786 (O_1786,N_29192,N_29336);
nor UO_1787 (O_1787,N_29727,N_28952);
and UO_1788 (O_1788,N_29071,N_28565);
and UO_1789 (O_1789,N_28654,N_28699);
nor UO_1790 (O_1790,N_29679,N_29798);
and UO_1791 (O_1791,N_29297,N_28847);
or UO_1792 (O_1792,N_28995,N_29065);
nand UO_1793 (O_1793,N_28631,N_28644);
nor UO_1794 (O_1794,N_28571,N_29502);
xnor UO_1795 (O_1795,N_29476,N_28848);
and UO_1796 (O_1796,N_28948,N_29700);
or UO_1797 (O_1797,N_28807,N_28508);
and UO_1798 (O_1798,N_29861,N_29405);
xor UO_1799 (O_1799,N_29159,N_28726);
nand UO_1800 (O_1800,N_29129,N_29533);
nand UO_1801 (O_1801,N_29125,N_29859);
xnor UO_1802 (O_1802,N_29137,N_29756);
nand UO_1803 (O_1803,N_29578,N_29223);
or UO_1804 (O_1804,N_29122,N_28545);
nand UO_1805 (O_1805,N_29802,N_28564);
and UO_1806 (O_1806,N_29828,N_29831);
and UO_1807 (O_1807,N_29940,N_29416);
xor UO_1808 (O_1808,N_28919,N_28730);
xor UO_1809 (O_1809,N_29093,N_28584);
nor UO_1810 (O_1810,N_29588,N_28848);
nand UO_1811 (O_1811,N_28879,N_29115);
nand UO_1812 (O_1812,N_29278,N_29114);
and UO_1813 (O_1813,N_29735,N_29467);
xor UO_1814 (O_1814,N_29512,N_28787);
and UO_1815 (O_1815,N_29011,N_28538);
nand UO_1816 (O_1816,N_29182,N_29271);
nand UO_1817 (O_1817,N_29936,N_29555);
nand UO_1818 (O_1818,N_29204,N_28742);
or UO_1819 (O_1819,N_29381,N_28906);
and UO_1820 (O_1820,N_28846,N_28853);
and UO_1821 (O_1821,N_28763,N_28803);
nor UO_1822 (O_1822,N_29273,N_28738);
nand UO_1823 (O_1823,N_28615,N_29397);
or UO_1824 (O_1824,N_28880,N_28776);
nor UO_1825 (O_1825,N_29692,N_29517);
nor UO_1826 (O_1826,N_29054,N_28702);
or UO_1827 (O_1827,N_28811,N_28907);
nor UO_1828 (O_1828,N_28879,N_29669);
nand UO_1829 (O_1829,N_29714,N_29615);
and UO_1830 (O_1830,N_28604,N_29360);
or UO_1831 (O_1831,N_28742,N_28974);
nand UO_1832 (O_1832,N_29737,N_29983);
or UO_1833 (O_1833,N_29808,N_29533);
or UO_1834 (O_1834,N_28767,N_28997);
and UO_1835 (O_1835,N_29864,N_29719);
nor UO_1836 (O_1836,N_29924,N_28776);
nor UO_1837 (O_1837,N_29005,N_29077);
nand UO_1838 (O_1838,N_29243,N_29289);
or UO_1839 (O_1839,N_28611,N_29475);
xnor UO_1840 (O_1840,N_28848,N_29677);
or UO_1841 (O_1841,N_28848,N_29223);
xnor UO_1842 (O_1842,N_29601,N_28503);
nand UO_1843 (O_1843,N_28815,N_29369);
nand UO_1844 (O_1844,N_28987,N_29163);
nor UO_1845 (O_1845,N_28777,N_29203);
or UO_1846 (O_1846,N_29723,N_29713);
xor UO_1847 (O_1847,N_29650,N_29693);
or UO_1848 (O_1848,N_29182,N_28788);
xor UO_1849 (O_1849,N_29717,N_29183);
and UO_1850 (O_1850,N_29620,N_28890);
or UO_1851 (O_1851,N_29732,N_29103);
nand UO_1852 (O_1852,N_28709,N_29085);
or UO_1853 (O_1853,N_28782,N_29108);
or UO_1854 (O_1854,N_29896,N_28791);
and UO_1855 (O_1855,N_28757,N_29335);
nand UO_1856 (O_1856,N_29010,N_29082);
nand UO_1857 (O_1857,N_29342,N_29840);
or UO_1858 (O_1858,N_28621,N_28509);
nor UO_1859 (O_1859,N_29118,N_29023);
xnor UO_1860 (O_1860,N_29581,N_28937);
xnor UO_1861 (O_1861,N_29558,N_29932);
or UO_1862 (O_1862,N_29753,N_29115);
and UO_1863 (O_1863,N_29822,N_28838);
xor UO_1864 (O_1864,N_28592,N_28695);
nand UO_1865 (O_1865,N_29935,N_28581);
nor UO_1866 (O_1866,N_29300,N_29962);
or UO_1867 (O_1867,N_29252,N_29079);
xnor UO_1868 (O_1868,N_29006,N_29884);
nor UO_1869 (O_1869,N_28530,N_29713);
nor UO_1870 (O_1870,N_29060,N_29720);
and UO_1871 (O_1871,N_29085,N_28636);
and UO_1872 (O_1872,N_29603,N_29806);
xnor UO_1873 (O_1873,N_29515,N_29736);
nand UO_1874 (O_1874,N_29635,N_28524);
xor UO_1875 (O_1875,N_29545,N_29800);
and UO_1876 (O_1876,N_28568,N_29058);
and UO_1877 (O_1877,N_28908,N_29775);
and UO_1878 (O_1878,N_28578,N_29860);
xnor UO_1879 (O_1879,N_28600,N_29843);
nand UO_1880 (O_1880,N_28904,N_29853);
nand UO_1881 (O_1881,N_28934,N_29130);
or UO_1882 (O_1882,N_29238,N_29706);
nor UO_1883 (O_1883,N_28803,N_28782);
and UO_1884 (O_1884,N_28560,N_29372);
and UO_1885 (O_1885,N_29454,N_28795);
nand UO_1886 (O_1886,N_29708,N_29143);
nor UO_1887 (O_1887,N_29176,N_28758);
nand UO_1888 (O_1888,N_28581,N_28834);
and UO_1889 (O_1889,N_29092,N_29548);
nor UO_1890 (O_1890,N_29589,N_29719);
nand UO_1891 (O_1891,N_29318,N_29346);
nor UO_1892 (O_1892,N_29019,N_28697);
xnor UO_1893 (O_1893,N_29362,N_29596);
or UO_1894 (O_1894,N_29818,N_28722);
xor UO_1895 (O_1895,N_29292,N_29228);
or UO_1896 (O_1896,N_29781,N_28769);
xnor UO_1897 (O_1897,N_29725,N_29063);
and UO_1898 (O_1898,N_29303,N_29992);
xor UO_1899 (O_1899,N_29811,N_28686);
and UO_1900 (O_1900,N_29532,N_29849);
nand UO_1901 (O_1901,N_28774,N_28930);
and UO_1902 (O_1902,N_28677,N_28735);
nor UO_1903 (O_1903,N_28876,N_28962);
nor UO_1904 (O_1904,N_29104,N_28555);
nor UO_1905 (O_1905,N_29565,N_29935);
xor UO_1906 (O_1906,N_29762,N_28778);
xor UO_1907 (O_1907,N_29859,N_29225);
xor UO_1908 (O_1908,N_28798,N_28707);
nand UO_1909 (O_1909,N_29685,N_29489);
nand UO_1910 (O_1910,N_29981,N_29983);
nand UO_1911 (O_1911,N_28813,N_28574);
xor UO_1912 (O_1912,N_28708,N_29565);
or UO_1913 (O_1913,N_29793,N_29000);
or UO_1914 (O_1914,N_29173,N_28783);
nand UO_1915 (O_1915,N_28959,N_29676);
and UO_1916 (O_1916,N_29778,N_29324);
nor UO_1917 (O_1917,N_29246,N_28728);
xnor UO_1918 (O_1918,N_29751,N_29585);
and UO_1919 (O_1919,N_29729,N_29308);
or UO_1920 (O_1920,N_29001,N_28607);
or UO_1921 (O_1921,N_29018,N_28984);
nor UO_1922 (O_1922,N_29992,N_29098);
nor UO_1923 (O_1923,N_29878,N_29716);
nor UO_1924 (O_1924,N_29079,N_29208);
or UO_1925 (O_1925,N_29463,N_28501);
xor UO_1926 (O_1926,N_29942,N_29587);
or UO_1927 (O_1927,N_28856,N_29872);
and UO_1928 (O_1928,N_29654,N_29683);
and UO_1929 (O_1929,N_29230,N_29820);
xor UO_1930 (O_1930,N_28822,N_28515);
nand UO_1931 (O_1931,N_28853,N_29592);
nor UO_1932 (O_1932,N_29103,N_29496);
nor UO_1933 (O_1933,N_29994,N_29932);
nor UO_1934 (O_1934,N_29141,N_29605);
xor UO_1935 (O_1935,N_28673,N_29118);
xor UO_1936 (O_1936,N_29661,N_29908);
or UO_1937 (O_1937,N_29190,N_28826);
and UO_1938 (O_1938,N_29478,N_29293);
nor UO_1939 (O_1939,N_29302,N_29942);
nand UO_1940 (O_1940,N_29396,N_28958);
and UO_1941 (O_1941,N_29246,N_29358);
nor UO_1942 (O_1942,N_29961,N_29812);
nor UO_1943 (O_1943,N_29774,N_29947);
nor UO_1944 (O_1944,N_29085,N_29395);
and UO_1945 (O_1945,N_28849,N_29247);
nand UO_1946 (O_1946,N_29257,N_29171);
nor UO_1947 (O_1947,N_29510,N_29064);
or UO_1948 (O_1948,N_29937,N_28727);
or UO_1949 (O_1949,N_29061,N_29485);
xnor UO_1950 (O_1950,N_29511,N_29840);
or UO_1951 (O_1951,N_29392,N_29386);
nor UO_1952 (O_1952,N_29172,N_28886);
nor UO_1953 (O_1953,N_29023,N_29543);
nor UO_1954 (O_1954,N_28609,N_28948);
and UO_1955 (O_1955,N_29836,N_28825);
xnor UO_1956 (O_1956,N_28860,N_29768);
or UO_1957 (O_1957,N_28921,N_28898);
nand UO_1958 (O_1958,N_29915,N_29276);
or UO_1959 (O_1959,N_28947,N_29625);
nor UO_1960 (O_1960,N_28535,N_29628);
nor UO_1961 (O_1961,N_29917,N_29366);
nor UO_1962 (O_1962,N_28557,N_29671);
nor UO_1963 (O_1963,N_28901,N_29545);
or UO_1964 (O_1964,N_29071,N_28923);
nor UO_1965 (O_1965,N_29664,N_29847);
nand UO_1966 (O_1966,N_29232,N_29746);
xor UO_1967 (O_1967,N_29205,N_29051);
and UO_1968 (O_1968,N_29127,N_29718);
or UO_1969 (O_1969,N_28988,N_29078);
nand UO_1970 (O_1970,N_29473,N_29801);
and UO_1971 (O_1971,N_29511,N_29079);
xor UO_1972 (O_1972,N_28888,N_29951);
nand UO_1973 (O_1973,N_29666,N_28869);
xor UO_1974 (O_1974,N_29223,N_28643);
or UO_1975 (O_1975,N_29724,N_29141);
nand UO_1976 (O_1976,N_29798,N_28561);
nor UO_1977 (O_1977,N_28997,N_29545);
nand UO_1978 (O_1978,N_29055,N_28574);
and UO_1979 (O_1979,N_29775,N_29922);
nand UO_1980 (O_1980,N_29285,N_29990);
nor UO_1981 (O_1981,N_28717,N_29112);
nor UO_1982 (O_1982,N_29787,N_29797);
nor UO_1983 (O_1983,N_28506,N_29052);
xnor UO_1984 (O_1984,N_28975,N_28788);
or UO_1985 (O_1985,N_29075,N_29341);
nor UO_1986 (O_1986,N_29060,N_29682);
and UO_1987 (O_1987,N_28692,N_28661);
and UO_1988 (O_1988,N_29872,N_29549);
nor UO_1989 (O_1989,N_28774,N_29135);
and UO_1990 (O_1990,N_29388,N_29218);
nand UO_1991 (O_1991,N_29437,N_29273);
nand UO_1992 (O_1992,N_29032,N_28562);
or UO_1993 (O_1993,N_29338,N_29464);
xnor UO_1994 (O_1994,N_28884,N_29813);
xor UO_1995 (O_1995,N_29908,N_28599);
nand UO_1996 (O_1996,N_29875,N_29330);
xor UO_1997 (O_1997,N_29073,N_29401);
and UO_1998 (O_1998,N_29700,N_29965);
or UO_1999 (O_1999,N_28815,N_29850);
and UO_2000 (O_2000,N_29273,N_29958);
or UO_2001 (O_2001,N_29192,N_29238);
nand UO_2002 (O_2002,N_29484,N_29618);
or UO_2003 (O_2003,N_29268,N_28518);
nand UO_2004 (O_2004,N_29273,N_29868);
nand UO_2005 (O_2005,N_29782,N_28863);
nand UO_2006 (O_2006,N_29844,N_28561);
nand UO_2007 (O_2007,N_29093,N_28848);
xor UO_2008 (O_2008,N_28675,N_29115);
or UO_2009 (O_2009,N_29238,N_29746);
nand UO_2010 (O_2010,N_29889,N_29565);
nand UO_2011 (O_2011,N_28757,N_29516);
xor UO_2012 (O_2012,N_28508,N_28643);
nor UO_2013 (O_2013,N_29286,N_28751);
or UO_2014 (O_2014,N_29305,N_29639);
and UO_2015 (O_2015,N_29219,N_28773);
xnor UO_2016 (O_2016,N_28980,N_29577);
xor UO_2017 (O_2017,N_28869,N_28541);
xnor UO_2018 (O_2018,N_28501,N_29084);
and UO_2019 (O_2019,N_28602,N_29739);
nor UO_2020 (O_2020,N_28801,N_29536);
or UO_2021 (O_2021,N_28533,N_28938);
or UO_2022 (O_2022,N_29238,N_29171);
nor UO_2023 (O_2023,N_29820,N_29607);
xnor UO_2024 (O_2024,N_29314,N_29381);
xor UO_2025 (O_2025,N_28564,N_29115);
xnor UO_2026 (O_2026,N_28982,N_28981);
or UO_2027 (O_2027,N_29744,N_29335);
nor UO_2028 (O_2028,N_29517,N_29662);
xor UO_2029 (O_2029,N_29077,N_29844);
nand UO_2030 (O_2030,N_29578,N_29724);
xor UO_2031 (O_2031,N_29927,N_29158);
nand UO_2032 (O_2032,N_28568,N_29730);
nand UO_2033 (O_2033,N_29560,N_29460);
or UO_2034 (O_2034,N_28880,N_28514);
nor UO_2035 (O_2035,N_29184,N_29676);
nand UO_2036 (O_2036,N_28646,N_29804);
and UO_2037 (O_2037,N_29134,N_29698);
nand UO_2038 (O_2038,N_28790,N_29391);
or UO_2039 (O_2039,N_28718,N_28897);
xnor UO_2040 (O_2040,N_28824,N_29270);
and UO_2041 (O_2041,N_29040,N_29819);
nor UO_2042 (O_2042,N_29348,N_29978);
nand UO_2043 (O_2043,N_28827,N_29411);
nor UO_2044 (O_2044,N_29464,N_28756);
and UO_2045 (O_2045,N_28510,N_28681);
and UO_2046 (O_2046,N_29236,N_29353);
xnor UO_2047 (O_2047,N_28633,N_29951);
xor UO_2048 (O_2048,N_29543,N_29991);
nor UO_2049 (O_2049,N_28878,N_28520);
xor UO_2050 (O_2050,N_28868,N_29026);
nand UO_2051 (O_2051,N_29422,N_29291);
nor UO_2052 (O_2052,N_29190,N_29641);
and UO_2053 (O_2053,N_28786,N_28827);
nand UO_2054 (O_2054,N_29207,N_28653);
nor UO_2055 (O_2055,N_29075,N_29974);
xnor UO_2056 (O_2056,N_28596,N_29419);
or UO_2057 (O_2057,N_29645,N_29134);
and UO_2058 (O_2058,N_29721,N_29886);
and UO_2059 (O_2059,N_29271,N_28746);
nand UO_2060 (O_2060,N_29671,N_29254);
nand UO_2061 (O_2061,N_28597,N_28625);
and UO_2062 (O_2062,N_28828,N_29821);
nand UO_2063 (O_2063,N_29625,N_29181);
nand UO_2064 (O_2064,N_29596,N_28621);
nand UO_2065 (O_2065,N_29813,N_29530);
xnor UO_2066 (O_2066,N_28500,N_29841);
nor UO_2067 (O_2067,N_28951,N_29411);
and UO_2068 (O_2068,N_28511,N_29577);
nand UO_2069 (O_2069,N_29851,N_29629);
nand UO_2070 (O_2070,N_29250,N_29582);
nand UO_2071 (O_2071,N_28557,N_28758);
or UO_2072 (O_2072,N_29167,N_29034);
nor UO_2073 (O_2073,N_29546,N_29007);
xor UO_2074 (O_2074,N_29592,N_29195);
nand UO_2075 (O_2075,N_29343,N_28853);
xor UO_2076 (O_2076,N_29992,N_28874);
or UO_2077 (O_2077,N_29591,N_28602);
and UO_2078 (O_2078,N_29647,N_29946);
or UO_2079 (O_2079,N_28894,N_29503);
and UO_2080 (O_2080,N_29641,N_29864);
nor UO_2081 (O_2081,N_29498,N_29387);
xor UO_2082 (O_2082,N_29808,N_29124);
xor UO_2083 (O_2083,N_28545,N_28790);
xnor UO_2084 (O_2084,N_29510,N_28514);
nand UO_2085 (O_2085,N_29604,N_29911);
or UO_2086 (O_2086,N_29793,N_28776);
xor UO_2087 (O_2087,N_29148,N_28539);
nor UO_2088 (O_2088,N_28536,N_29479);
nand UO_2089 (O_2089,N_29791,N_28767);
nand UO_2090 (O_2090,N_28595,N_29325);
or UO_2091 (O_2091,N_28952,N_29244);
nor UO_2092 (O_2092,N_29798,N_29353);
nor UO_2093 (O_2093,N_29004,N_28524);
nand UO_2094 (O_2094,N_29811,N_29156);
nor UO_2095 (O_2095,N_29187,N_29692);
xnor UO_2096 (O_2096,N_29457,N_28940);
nand UO_2097 (O_2097,N_29123,N_29013);
and UO_2098 (O_2098,N_28794,N_29143);
xor UO_2099 (O_2099,N_28733,N_28738);
nor UO_2100 (O_2100,N_29217,N_29658);
and UO_2101 (O_2101,N_29161,N_29143);
nand UO_2102 (O_2102,N_28829,N_28803);
nand UO_2103 (O_2103,N_29506,N_28806);
nor UO_2104 (O_2104,N_29290,N_29261);
nand UO_2105 (O_2105,N_29568,N_28597);
nor UO_2106 (O_2106,N_29964,N_29646);
nor UO_2107 (O_2107,N_29716,N_28535);
nor UO_2108 (O_2108,N_28581,N_29265);
and UO_2109 (O_2109,N_28843,N_29561);
and UO_2110 (O_2110,N_28960,N_29326);
or UO_2111 (O_2111,N_29113,N_29689);
and UO_2112 (O_2112,N_29909,N_28652);
nand UO_2113 (O_2113,N_29305,N_29319);
nand UO_2114 (O_2114,N_28529,N_29136);
nand UO_2115 (O_2115,N_28584,N_28512);
nand UO_2116 (O_2116,N_29451,N_29329);
xnor UO_2117 (O_2117,N_28689,N_29495);
nor UO_2118 (O_2118,N_28978,N_29131);
and UO_2119 (O_2119,N_29439,N_29574);
xnor UO_2120 (O_2120,N_29057,N_29097);
nor UO_2121 (O_2121,N_29505,N_29383);
or UO_2122 (O_2122,N_29083,N_28529);
nand UO_2123 (O_2123,N_29981,N_29887);
xnor UO_2124 (O_2124,N_29179,N_29817);
nand UO_2125 (O_2125,N_29752,N_28682);
nand UO_2126 (O_2126,N_28710,N_29576);
nor UO_2127 (O_2127,N_29337,N_29424);
nor UO_2128 (O_2128,N_28728,N_29613);
nor UO_2129 (O_2129,N_29780,N_28721);
nor UO_2130 (O_2130,N_29502,N_29324);
nor UO_2131 (O_2131,N_28726,N_29718);
nand UO_2132 (O_2132,N_29555,N_29922);
xnor UO_2133 (O_2133,N_28671,N_28776);
and UO_2134 (O_2134,N_29100,N_29392);
xnor UO_2135 (O_2135,N_29933,N_29254);
nand UO_2136 (O_2136,N_29671,N_28872);
nor UO_2137 (O_2137,N_29835,N_29177);
and UO_2138 (O_2138,N_29734,N_29505);
xor UO_2139 (O_2139,N_29317,N_29330);
nand UO_2140 (O_2140,N_28534,N_29959);
nand UO_2141 (O_2141,N_29819,N_29940);
xnor UO_2142 (O_2142,N_28848,N_29290);
nand UO_2143 (O_2143,N_28972,N_28901);
xor UO_2144 (O_2144,N_29779,N_29344);
and UO_2145 (O_2145,N_28921,N_28959);
xnor UO_2146 (O_2146,N_28657,N_28539);
and UO_2147 (O_2147,N_28888,N_29188);
xnor UO_2148 (O_2148,N_28750,N_29989);
and UO_2149 (O_2149,N_28823,N_29941);
or UO_2150 (O_2150,N_29795,N_29659);
nand UO_2151 (O_2151,N_28526,N_28746);
and UO_2152 (O_2152,N_29141,N_28512);
nor UO_2153 (O_2153,N_28775,N_29024);
and UO_2154 (O_2154,N_28689,N_28758);
and UO_2155 (O_2155,N_28849,N_29221);
xnor UO_2156 (O_2156,N_28615,N_29039);
or UO_2157 (O_2157,N_28826,N_28974);
xor UO_2158 (O_2158,N_29471,N_29815);
or UO_2159 (O_2159,N_29125,N_28968);
nand UO_2160 (O_2160,N_28786,N_29452);
and UO_2161 (O_2161,N_29768,N_28665);
nand UO_2162 (O_2162,N_28881,N_29417);
xnor UO_2163 (O_2163,N_29017,N_29786);
xor UO_2164 (O_2164,N_29341,N_29058);
and UO_2165 (O_2165,N_29950,N_29829);
nor UO_2166 (O_2166,N_29403,N_29001);
xnor UO_2167 (O_2167,N_29557,N_29162);
nand UO_2168 (O_2168,N_28817,N_28794);
xor UO_2169 (O_2169,N_29010,N_29830);
nor UO_2170 (O_2170,N_29403,N_29204);
or UO_2171 (O_2171,N_28562,N_29290);
nor UO_2172 (O_2172,N_28601,N_29249);
nand UO_2173 (O_2173,N_29904,N_29840);
nor UO_2174 (O_2174,N_28704,N_28604);
nor UO_2175 (O_2175,N_29333,N_29019);
and UO_2176 (O_2176,N_29949,N_29620);
and UO_2177 (O_2177,N_29270,N_28766);
xor UO_2178 (O_2178,N_29221,N_29409);
and UO_2179 (O_2179,N_29663,N_28621);
nand UO_2180 (O_2180,N_28765,N_28992);
or UO_2181 (O_2181,N_29923,N_29442);
nand UO_2182 (O_2182,N_29683,N_28991);
nor UO_2183 (O_2183,N_29465,N_29818);
and UO_2184 (O_2184,N_28825,N_28971);
or UO_2185 (O_2185,N_28921,N_28656);
nand UO_2186 (O_2186,N_29006,N_29222);
and UO_2187 (O_2187,N_29379,N_29786);
xnor UO_2188 (O_2188,N_29563,N_28775);
or UO_2189 (O_2189,N_28772,N_29781);
or UO_2190 (O_2190,N_29065,N_29655);
nor UO_2191 (O_2191,N_29052,N_29849);
nor UO_2192 (O_2192,N_28820,N_29536);
nor UO_2193 (O_2193,N_29341,N_29544);
xor UO_2194 (O_2194,N_29346,N_28855);
and UO_2195 (O_2195,N_29297,N_29021);
xor UO_2196 (O_2196,N_29394,N_29077);
nor UO_2197 (O_2197,N_29782,N_29177);
or UO_2198 (O_2198,N_29432,N_29445);
nand UO_2199 (O_2199,N_29014,N_29282);
nand UO_2200 (O_2200,N_29042,N_29934);
nor UO_2201 (O_2201,N_29569,N_29993);
nand UO_2202 (O_2202,N_28563,N_29380);
nand UO_2203 (O_2203,N_29937,N_29569);
nor UO_2204 (O_2204,N_29143,N_29886);
nor UO_2205 (O_2205,N_28786,N_29252);
xor UO_2206 (O_2206,N_29716,N_29254);
nand UO_2207 (O_2207,N_29197,N_28718);
and UO_2208 (O_2208,N_29931,N_28989);
and UO_2209 (O_2209,N_29554,N_29333);
nand UO_2210 (O_2210,N_29687,N_29173);
or UO_2211 (O_2211,N_28857,N_29922);
nand UO_2212 (O_2212,N_29361,N_29129);
or UO_2213 (O_2213,N_28996,N_28626);
or UO_2214 (O_2214,N_28586,N_29158);
nand UO_2215 (O_2215,N_29445,N_29754);
xnor UO_2216 (O_2216,N_29970,N_29836);
nor UO_2217 (O_2217,N_29256,N_29805);
nand UO_2218 (O_2218,N_28562,N_28813);
nor UO_2219 (O_2219,N_29815,N_29419);
or UO_2220 (O_2220,N_29828,N_29687);
nand UO_2221 (O_2221,N_28879,N_29682);
nand UO_2222 (O_2222,N_29908,N_29391);
xnor UO_2223 (O_2223,N_28589,N_28916);
nand UO_2224 (O_2224,N_29505,N_29237);
nor UO_2225 (O_2225,N_28750,N_28574);
or UO_2226 (O_2226,N_28935,N_29010);
nor UO_2227 (O_2227,N_29572,N_29281);
or UO_2228 (O_2228,N_29864,N_29941);
nand UO_2229 (O_2229,N_29171,N_29665);
nand UO_2230 (O_2230,N_29880,N_29492);
nand UO_2231 (O_2231,N_28835,N_29378);
and UO_2232 (O_2232,N_28904,N_28578);
xnor UO_2233 (O_2233,N_29218,N_28623);
or UO_2234 (O_2234,N_28663,N_29318);
xor UO_2235 (O_2235,N_28817,N_28819);
or UO_2236 (O_2236,N_28668,N_29948);
and UO_2237 (O_2237,N_28696,N_29483);
and UO_2238 (O_2238,N_29509,N_28609);
and UO_2239 (O_2239,N_29148,N_29928);
or UO_2240 (O_2240,N_29561,N_29095);
or UO_2241 (O_2241,N_29046,N_29709);
nor UO_2242 (O_2242,N_29477,N_29245);
nor UO_2243 (O_2243,N_29750,N_29186);
nor UO_2244 (O_2244,N_28670,N_28946);
or UO_2245 (O_2245,N_28539,N_29773);
or UO_2246 (O_2246,N_29175,N_29533);
or UO_2247 (O_2247,N_29872,N_28841);
nand UO_2248 (O_2248,N_29167,N_29860);
or UO_2249 (O_2249,N_29540,N_29357);
and UO_2250 (O_2250,N_28959,N_29477);
and UO_2251 (O_2251,N_29813,N_28810);
or UO_2252 (O_2252,N_29343,N_28917);
or UO_2253 (O_2253,N_28885,N_28977);
nor UO_2254 (O_2254,N_29879,N_29031);
xor UO_2255 (O_2255,N_29362,N_28694);
nor UO_2256 (O_2256,N_29043,N_28765);
or UO_2257 (O_2257,N_28721,N_29607);
nand UO_2258 (O_2258,N_29371,N_29479);
xnor UO_2259 (O_2259,N_28857,N_29100);
or UO_2260 (O_2260,N_29855,N_29818);
and UO_2261 (O_2261,N_29907,N_28959);
and UO_2262 (O_2262,N_28999,N_29614);
and UO_2263 (O_2263,N_28576,N_29873);
and UO_2264 (O_2264,N_29140,N_28596);
nand UO_2265 (O_2265,N_29953,N_29383);
and UO_2266 (O_2266,N_29003,N_28589);
xnor UO_2267 (O_2267,N_28991,N_29870);
and UO_2268 (O_2268,N_29363,N_28959);
or UO_2269 (O_2269,N_28934,N_29688);
nand UO_2270 (O_2270,N_29684,N_29125);
nor UO_2271 (O_2271,N_29453,N_29814);
nor UO_2272 (O_2272,N_28995,N_29000);
or UO_2273 (O_2273,N_29571,N_29265);
or UO_2274 (O_2274,N_28652,N_28909);
xnor UO_2275 (O_2275,N_29290,N_29026);
xor UO_2276 (O_2276,N_29404,N_28513);
or UO_2277 (O_2277,N_29134,N_29817);
and UO_2278 (O_2278,N_29744,N_28878);
nand UO_2279 (O_2279,N_29706,N_29268);
and UO_2280 (O_2280,N_28525,N_29484);
nand UO_2281 (O_2281,N_29468,N_28689);
xor UO_2282 (O_2282,N_28819,N_29050);
or UO_2283 (O_2283,N_28511,N_29773);
xnor UO_2284 (O_2284,N_28780,N_29783);
nor UO_2285 (O_2285,N_28860,N_29978);
or UO_2286 (O_2286,N_28967,N_29655);
xnor UO_2287 (O_2287,N_28834,N_29745);
or UO_2288 (O_2288,N_29871,N_28555);
xnor UO_2289 (O_2289,N_29815,N_29404);
or UO_2290 (O_2290,N_29151,N_29105);
nand UO_2291 (O_2291,N_28800,N_28885);
or UO_2292 (O_2292,N_28545,N_28586);
xnor UO_2293 (O_2293,N_29409,N_29142);
nand UO_2294 (O_2294,N_29765,N_28551);
xor UO_2295 (O_2295,N_29384,N_29876);
and UO_2296 (O_2296,N_29074,N_29817);
nand UO_2297 (O_2297,N_29660,N_29853);
and UO_2298 (O_2298,N_29369,N_28936);
or UO_2299 (O_2299,N_28956,N_28812);
or UO_2300 (O_2300,N_28974,N_28702);
and UO_2301 (O_2301,N_29089,N_29854);
nand UO_2302 (O_2302,N_29158,N_29555);
nor UO_2303 (O_2303,N_29841,N_29949);
and UO_2304 (O_2304,N_28841,N_29422);
nor UO_2305 (O_2305,N_29827,N_29686);
xor UO_2306 (O_2306,N_28879,N_28770);
or UO_2307 (O_2307,N_29875,N_29874);
nand UO_2308 (O_2308,N_28630,N_29013);
nor UO_2309 (O_2309,N_29577,N_29990);
nor UO_2310 (O_2310,N_29444,N_28860);
or UO_2311 (O_2311,N_29316,N_29242);
nor UO_2312 (O_2312,N_29909,N_29377);
nand UO_2313 (O_2313,N_29722,N_29291);
xor UO_2314 (O_2314,N_29203,N_29982);
nor UO_2315 (O_2315,N_29720,N_29898);
or UO_2316 (O_2316,N_28657,N_29075);
nor UO_2317 (O_2317,N_29595,N_29441);
nor UO_2318 (O_2318,N_29523,N_29102);
nor UO_2319 (O_2319,N_29304,N_29050);
nor UO_2320 (O_2320,N_28681,N_28650);
nand UO_2321 (O_2321,N_28658,N_29203);
or UO_2322 (O_2322,N_29604,N_28648);
xnor UO_2323 (O_2323,N_28796,N_29587);
nand UO_2324 (O_2324,N_28953,N_28750);
or UO_2325 (O_2325,N_29805,N_28884);
or UO_2326 (O_2326,N_29349,N_28557);
and UO_2327 (O_2327,N_29576,N_29160);
and UO_2328 (O_2328,N_29989,N_29174);
xnor UO_2329 (O_2329,N_29514,N_28898);
nand UO_2330 (O_2330,N_29458,N_29687);
and UO_2331 (O_2331,N_28972,N_28920);
and UO_2332 (O_2332,N_29830,N_29755);
xor UO_2333 (O_2333,N_29678,N_29737);
nor UO_2334 (O_2334,N_29029,N_28974);
or UO_2335 (O_2335,N_29341,N_29215);
nand UO_2336 (O_2336,N_29245,N_29593);
and UO_2337 (O_2337,N_29592,N_29649);
xor UO_2338 (O_2338,N_29516,N_29962);
nor UO_2339 (O_2339,N_29864,N_29792);
nor UO_2340 (O_2340,N_29552,N_28627);
nor UO_2341 (O_2341,N_29106,N_28506);
or UO_2342 (O_2342,N_28517,N_28579);
xnor UO_2343 (O_2343,N_29951,N_28779);
nand UO_2344 (O_2344,N_29488,N_28668);
or UO_2345 (O_2345,N_28548,N_28800);
or UO_2346 (O_2346,N_29142,N_28733);
nor UO_2347 (O_2347,N_29268,N_29965);
nand UO_2348 (O_2348,N_29715,N_28958);
nor UO_2349 (O_2349,N_29372,N_29600);
and UO_2350 (O_2350,N_29423,N_28966);
nor UO_2351 (O_2351,N_29240,N_29303);
nand UO_2352 (O_2352,N_29464,N_29574);
nand UO_2353 (O_2353,N_28625,N_28661);
and UO_2354 (O_2354,N_29882,N_29575);
nand UO_2355 (O_2355,N_29448,N_28865);
xor UO_2356 (O_2356,N_28769,N_28774);
xor UO_2357 (O_2357,N_29497,N_29278);
nand UO_2358 (O_2358,N_28612,N_29957);
nor UO_2359 (O_2359,N_28825,N_29683);
and UO_2360 (O_2360,N_29735,N_29748);
nor UO_2361 (O_2361,N_28830,N_29790);
xor UO_2362 (O_2362,N_28962,N_29777);
or UO_2363 (O_2363,N_29715,N_29466);
nand UO_2364 (O_2364,N_29212,N_29979);
xor UO_2365 (O_2365,N_29968,N_29698);
or UO_2366 (O_2366,N_28847,N_29661);
nor UO_2367 (O_2367,N_29725,N_29846);
or UO_2368 (O_2368,N_28952,N_29797);
nor UO_2369 (O_2369,N_29915,N_29265);
nand UO_2370 (O_2370,N_29046,N_28872);
or UO_2371 (O_2371,N_28536,N_29316);
or UO_2372 (O_2372,N_29432,N_28904);
nand UO_2373 (O_2373,N_29407,N_29696);
and UO_2374 (O_2374,N_29492,N_29751);
and UO_2375 (O_2375,N_29767,N_28897);
xor UO_2376 (O_2376,N_29430,N_28637);
nor UO_2377 (O_2377,N_29505,N_29653);
or UO_2378 (O_2378,N_29417,N_29633);
and UO_2379 (O_2379,N_28857,N_28950);
and UO_2380 (O_2380,N_29018,N_28577);
or UO_2381 (O_2381,N_28957,N_29464);
nand UO_2382 (O_2382,N_29639,N_28540);
xnor UO_2383 (O_2383,N_28910,N_29178);
and UO_2384 (O_2384,N_29209,N_28813);
xor UO_2385 (O_2385,N_29791,N_29049);
or UO_2386 (O_2386,N_28759,N_28921);
nor UO_2387 (O_2387,N_29540,N_28637);
and UO_2388 (O_2388,N_28719,N_28507);
nor UO_2389 (O_2389,N_29265,N_28964);
and UO_2390 (O_2390,N_29763,N_29453);
or UO_2391 (O_2391,N_29385,N_29473);
or UO_2392 (O_2392,N_28628,N_29154);
or UO_2393 (O_2393,N_29109,N_28727);
or UO_2394 (O_2394,N_29692,N_29565);
nor UO_2395 (O_2395,N_28726,N_29317);
nor UO_2396 (O_2396,N_29544,N_29676);
xnor UO_2397 (O_2397,N_29085,N_28885);
or UO_2398 (O_2398,N_29220,N_29938);
nor UO_2399 (O_2399,N_29528,N_29846);
nor UO_2400 (O_2400,N_28585,N_29079);
xor UO_2401 (O_2401,N_29784,N_29207);
nand UO_2402 (O_2402,N_29237,N_28665);
or UO_2403 (O_2403,N_29900,N_28968);
nor UO_2404 (O_2404,N_29987,N_29931);
nand UO_2405 (O_2405,N_29769,N_29765);
xor UO_2406 (O_2406,N_29754,N_29241);
xnor UO_2407 (O_2407,N_29399,N_29782);
nor UO_2408 (O_2408,N_29498,N_28592);
xor UO_2409 (O_2409,N_28949,N_29116);
xor UO_2410 (O_2410,N_28994,N_28534);
and UO_2411 (O_2411,N_29087,N_29624);
and UO_2412 (O_2412,N_29060,N_28582);
or UO_2413 (O_2413,N_28835,N_29280);
nor UO_2414 (O_2414,N_29689,N_28509);
xnor UO_2415 (O_2415,N_29048,N_28757);
and UO_2416 (O_2416,N_29314,N_28840);
xor UO_2417 (O_2417,N_29069,N_29927);
xor UO_2418 (O_2418,N_29941,N_28520);
and UO_2419 (O_2419,N_29403,N_29702);
xnor UO_2420 (O_2420,N_28549,N_29189);
or UO_2421 (O_2421,N_29667,N_28840);
or UO_2422 (O_2422,N_28935,N_28819);
nand UO_2423 (O_2423,N_29888,N_29459);
or UO_2424 (O_2424,N_29649,N_28689);
nand UO_2425 (O_2425,N_29292,N_28701);
nand UO_2426 (O_2426,N_28583,N_28828);
nand UO_2427 (O_2427,N_28624,N_29809);
or UO_2428 (O_2428,N_29273,N_29516);
xor UO_2429 (O_2429,N_29423,N_29792);
or UO_2430 (O_2430,N_28566,N_28699);
xor UO_2431 (O_2431,N_29395,N_29750);
and UO_2432 (O_2432,N_29903,N_29867);
and UO_2433 (O_2433,N_29680,N_29783);
or UO_2434 (O_2434,N_29878,N_29596);
nand UO_2435 (O_2435,N_28658,N_29523);
and UO_2436 (O_2436,N_29943,N_29947);
nor UO_2437 (O_2437,N_28644,N_29840);
or UO_2438 (O_2438,N_28735,N_29696);
or UO_2439 (O_2439,N_28883,N_29267);
xnor UO_2440 (O_2440,N_29623,N_29283);
nand UO_2441 (O_2441,N_29400,N_28575);
nand UO_2442 (O_2442,N_29040,N_28544);
nor UO_2443 (O_2443,N_28697,N_29175);
nor UO_2444 (O_2444,N_29164,N_29347);
xor UO_2445 (O_2445,N_29068,N_29692);
xor UO_2446 (O_2446,N_29701,N_29571);
or UO_2447 (O_2447,N_29436,N_29884);
nor UO_2448 (O_2448,N_28595,N_29684);
and UO_2449 (O_2449,N_29055,N_28941);
xor UO_2450 (O_2450,N_28656,N_29999);
and UO_2451 (O_2451,N_29774,N_29228);
nand UO_2452 (O_2452,N_28786,N_29521);
and UO_2453 (O_2453,N_28616,N_28524);
xor UO_2454 (O_2454,N_29045,N_29608);
nor UO_2455 (O_2455,N_29865,N_29022);
and UO_2456 (O_2456,N_28982,N_28893);
xor UO_2457 (O_2457,N_28941,N_28596);
xor UO_2458 (O_2458,N_29753,N_29380);
or UO_2459 (O_2459,N_29612,N_29067);
xnor UO_2460 (O_2460,N_28564,N_29932);
nor UO_2461 (O_2461,N_29551,N_29501);
nand UO_2462 (O_2462,N_29305,N_29682);
nand UO_2463 (O_2463,N_29730,N_28897);
nand UO_2464 (O_2464,N_29269,N_29685);
nor UO_2465 (O_2465,N_29420,N_29337);
nand UO_2466 (O_2466,N_28755,N_28811);
and UO_2467 (O_2467,N_29708,N_29810);
nor UO_2468 (O_2468,N_29829,N_28894);
or UO_2469 (O_2469,N_29270,N_29488);
or UO_2470 (O_2470,N_29767,N_28857);
nor UO_2471 (O_2471,N_29060,N_29893);
nor UO_2472 (O_2472,N_29824,N_29807);
nor UO_2473 (O_2473,N_28699,N_29154);
nand UO_2474 (O_2474,N_29556,N_29150);
nand UO_2475 (O_2475,N_29593,N_29380);
nor UO_2476 (O_2476,N_28706,N_28800);
or UO_2477 (O_2477,N_29124,N_28964);
xor UO_2478 (O_2478,N_28781,N_28691);
nor UO_2479 (O_2479,N_29323,N_29347);
nand UO_2480 (O_2480,N_29474,N_28890);
nand UO_2481 (O_2481,N_29343,N_28535);
nand UO_2482 (O_2482,N_29920,N_29566);
or UO_2483 (O_2483,N_28750,N_29543);
or UO_2484 (O_2484,N_28624,N_29375);
and UO_2485 (O_2485,N_29308,N_29333);
nand UO_2486 (O_2486,N_28723,N_29383);
nor UO_2487 (O_2487,N_29434,N_28950);
nand UO_2488 (O_2488,N_28979,N_29754);
xnor UO_2489 (O_2489,N_29535,N_29039);
and UO_2490 (O_2490,N_28670,N_28948);
nand UO_2491 (O_2491,N_29562,N_29639);
or UO_2492 (O_2492,N_29017,N_28533);
and UO_2493 (O_2493,N_28935,N_28767);
and UO_2494 (O_2494,N_28582,N_28906);
xnor UO_2495 (O_2495,N_29407,N_29561);
xor UO_2496 (O_2496,N_28879,N_29750);
xor UO_2497 (O_2497,N_29453,N_29137);
xor UO_2498 (O_2498,N_29715,N_28757);
or UO_2499 (O_2499,N_29172,N_29973);
nand UO_2500 (O_2500,N_28705,N_29600);
nor UO_2501 (O_2501,N_28950,N_29945);
and UO_2502 (O_2502,N_29866,N_29794);
nor UO_2503 (O_2503,N_28939,N_28687);
nor UO_2504 (O_2504,N_28950,N_29757);
nand UO_2505 (O_2505,N_28788,N_28973);
nand UO_2506 (O_2506,N_29753,N_29554);
and UO_2507 (O_2507,N_28789,N_28538);
and UO_2508 (O_2508,N_29110,N_28942);
nand UO_2509 (O_2509,N_28574,N_28935);
or UO_2510 (O_2510,N_29267,N_29690);
or UO_2511 (O_2511,N_28604,N_29731);
nand UO_2512 (O_2512,N_29000,N_29577);
and UO_2513 (O_2513,N_28691,N_29177);
nor UO_2514 (O_2514,N_29828,N_28791);
xnor UO_2515 (O_2515,N_29616,N_29437);
nand UO_2516 (O_2516,N_29006,N_29187);
and UO_2517 (O_2517,N_29559,N_29499);
and UO_2518 (O_2518,N_29587,N_28748);
nor UO_2519 (O_2519,N_29527,N_29491);
nand UO_2520 (O_2520,N_29572,N_28960);
nor UO_2521 (O_2521,N_29181,N_29226);
nand UO_2522 (O_2522,N_29701,N_29177);
nor UO_2523 (O_2523,N_28918,N_28866);
nand UO_2524 (O_2524,N_29113,N_29950);
nor UO_2525 (O_2525,N_28883,N_28888);
or UO_2526 (O_2526,N_29106,N_29305);
nand UO_2527 (O_2527,N_29962,N_28905);
and UO_2528 (O_2528,N_29243,N_28553);
nor UO_2529 (O_2529,N_28820,N_29159);
nand UO_2530 (O_2530,N_29116,N_29205);
nand UO_2531 (O_2531,N_29702,N_29613);
and UO_2532 (O_2532,N_28737,N_28942);
nand UO_2533 (O_2533,N_29100,N_29803);
nor UO_2534 (O_2534,N_29366,N_29220);
and UO_2535 (O_2535,N_28816,N_29149);
nor UO_2536 (O_2536,N_29817,N_28648);
and UO_2537 (O_2537,N_28906,N_29038);
nand UO_2538 (O_2538,N_29346,N_28888);
or UO_2539 (O_2539,N_29157,N_28893);
xor UO_2540 (O_2540,N_29068,N_29480);
xnor UO_2541 (O_2541,N_28942,N_28816);
nand UO_2542 (O_2542,N_29216,N_29952);
xor UO_2543 (O_2543,N_28797,N_29341);
nor UO_2544 (O_2544,N_29104,N_29176);
xor UO_2545 (O_2545,N_28586,N_28849);
or UO_2546 (O_2546,N_28551,N_29489);
and UO_2547 (O_2547,N_28976,N_29005);
nand UO_2548 (O_2548,N_28752,N_29397);
or UO_2549 (O_2549,N_28880,N_29487);
nor UO_2550 (O_2550,N_28920,N_29402);
xor UO_2551 (O_2551,N_29623,N_29998);
nor UO_2552 (O_2552,N_29557,N_28694);
nor UO_2553 (O_2553,N_28745,N_29215);
or UO_2554 (O_2554,N_28665,N_28737);
xnor UO_2555 (O_2555,N_29574,N_29495);
xor UO_2556 (O_2556,N_29911,N_29472);
nand UO_2557 (O_2557,N_29336,N_29082);
nor UO_2558 (O_2558,N_28593,N_28587);
nand UO_2559 (O_2559,N_29981,N_29437);
and UO_2560 (O_2560,N_28627,N_29049);
or UO_2561 (O_2561,N_28583,N_28751);
and UO_2562 (O_2562,N_29766,N_28621);
nand UO_2563 (O_2563,N_28809,N_28602);
xnor UO_2564 (O_2564,N_28911,N_29897);
nor UO_2565 (O_2565,N_29689,N_28581);
or UO_2566 (O_2566,N_29724,N_29319);
or UO_2567 (O_2567,N_28981,N_29139);
or UO_2568 (O_2568,N_29710,N_28835);
xor UO_2569 (O_2569,N_29787,N_28677);
or UO_2570 (O_2570,N_29451,N_29270);
nand UO_2571 (O_2571,N_29245,N_28978);
or UO_2572 (O_2572,N_28758,N_29964);
and UO_2573 (O_2573,N_29569,N_29083);
or UO_2574 (O_2574,N_29201,N_29323);
or UO_2575 (O_2575,N_29897,N_29693);
nor UO_2576 (O_2576,N_29858,N_28703);
or UO_2577 (O_2577,N_29283,N_29559);
nor UO_2578 (O_2578,N_29210,N_29802);
nor UO_2579 (O_2579,N_29392,N_29793);
xor UO_2580 (O_2580,N_29523,N_28605);
nor UO_2581 (O_2581,N_29160,N_29560);
and UO_2582 (O_2582,N_29797,N_29100);
nor UO_2583 (O_2583,N_29243,N_29311);
and UO_2584 (O_2584,N_29007,N_28796);
or UO_2585 (O_2585,N_29051,N_28743);
nand UO_2586 (O_2586,N_29787,N_29041);
nand UO_2587 (O_2587,N_29591,N_28693);
nand UO_2588 (O_2588,N_28951,N_29960);
xnor UO_2589 (O_2589,N_28847,N_28658);
and UO_2590 (O_2590,N_29217,N_29580);
xnor UO_2591 (O_2591,N_29627,N_28773);
nand UO_2592 (O_2592,N_29775,N_28793);
xor UO_2593 (O_2593,N_29316,N_29063);
or UO_2594 (O_2594,N_29951,N_28539);
xor UO_2595 (O_2595,N_29731,N_28725);
nor UO_2596 (O_2596,N_29494,N_28948);
or UO_2597 (O_2597,N_29349,N_29714);
or UO_2598 (O_2598,N_29457,N_28635);
or UO_2599 (O_2599,N_29223,N_29381);
xnor UO_2600 (O_2600,N_29700,N_29766);
or UO_2601 (O_2601,N_28667,N_29947);
or UO_2602 (O_2602,N_29744,N_29390);
nand UO_2603 (O_2603,N_28773,N_29061);
nand UO_2604 (O_2604,N_29740,N_28812);
or UO_2605 (O_2605,N_28660,N_29928);
and UO_2606 (O_2606,N_29134,N_29838);
nor UO_2607 (O_2607,N_28771,N_29203);
or UO_2608 (O_2608,N_29546,N_28580);
nor UO_2609 (O_2609,N_28501,N_29683);
xor UO_2610 (O_2610,N_29525,N_29117);
nand UO_2611 (O_2611,N_29692,N_29798);
nand UO_2612 (O_2612,N_29409,N_29608);
and UO_2613 (O_2613,N_28603,N_29808);
or UO_2614 (O_2614,N_28943,N_28795);
nand UO_2615 (O_2615,N_29418,N_29507);
nor UO_2616 (O_2616,N_29829,N_28518);
and UO_2617 (O_2617,N_29428,N_28961);
or UO_2618 (O_2618,N_28954,N_28765);
xnor UO_2619 (O_2619,N_28974,N_29820);
or UO_2620 (O_2620,N_29567,N_29236);
xnor UO_2621 (O_2621,N_29545,N_29803);
nor UO_2622 (O_2622,N_29907,N_29725);
nor UO_2623 (O_2623,N_29757,N_28554);
or UO_2624 (O_2624,N_29901,N_28688);
nand UO_2625 (O_2625,N_29227,N_28549);
and UO_2626 (O_2626,N_29837,N_28991);
and UO_2627 (O_2627,N_29821,N_29856);
and UO_2628 (O_2628,N_28655,N_28661);
xnor UO_2629 (O_2629,N_29749,N_29840);
nor UO_2630 (O_2630,N_29821,N_29289);
nor UO_2631 (O_2631,N_29179,N_29941);
nand UO_2632 (O_2632,N_29095,N_29829);
xnor UO_2633 (O_2633,N_28511,N_29061);
or UO_2634 (O_2634,N_29108,N_28591);
and UO_2635 (O_2635,N_29125,N_29142);
nand UO_2636 (O_2636,N_29869,N_28575);
or UO_2637 (O_2637,N_29315,N_28739);
or UO_2638 (O_2638,N_29598,N_28835);
or UO_2639 (O_2639,N_28866,N_28544);
and UO_2640 (O_2640,N_29146,N_28594);
or UO_2641 (O_2641,N_29946,N_29640);
nand UO_2642 (O_2642,N_29510,N_28888);
nand UO_2643 (O_2643,N_28766,N_28534);
nor UO_2644 (O_2644,N_29645,N_28880);
nor UO_2645 (O_2645,N_29519,N_29594);
xor UO_2646 (O_2646,N_29458,N_28544);
or UO_2647 (O_2647,N_29903,N_28984);
xnor UO_2648 (O_2648,N_29841,N_28987);
and UO_2649 (O_2649,N_29170,N_29533);
or UO_2650 (O_2650,N_29673,N_28586);
xor UO_2651 (O_2651,N_29802,N_29207);
xor UO_2652 (O_2652,N_28765,N_28628);
xor UO_2653 (O_2653,N_29284,N_29987);
and UO_2654 (O_2654,N_28777,N_29924);
or UO_2655 (O_2655,N_29753,N_29704);
nor UO_2656 (O_2656,N_29239,N_28716);
xnor UO_2657 (O_2657,N_28761,N_28725);
nand UO_2658 (O_2658,N_28659,N_28658);
or UO_2659 (O_2659,N_28748,N_28583);
nand UO_2660 (O_2660,N_28952,N_29077);
nor UO_2661 (O_2661,N_28608,N_29588);
or UO_2662 (O_2662,N_29067,N_29322);
or UO_2663 (O_2663,N_29762,N_29992);
xor UO_2664 (O_2664,N_29649,N_29832);
nor UO_2665 (O_2665,N_28949,N_28851);
or UO_2666 (O_2666,N_28622,N_28627);
or UO_2667 (O_2667,N_28932,N_29297);
nor UO_2668 (O_2668,N_28591,N_29659);
nand UO_2669 (O_2669,N_29259,N_29078);
nand UO_2670 (O_2670,N_29688,N_29724);
and UO_2671 (O_2671,N_29061,N_29681);
or UO_2672 (O_2672,N_29392,N_29010);
nor UO_2673 (O_2673,N_28649,N_29784);
nor UO_2674 (O_2674,N_29757,N_28760);
or UO_2675 (O_2675,N_29194,N_29842);
and UO_2676 (O_2676,N_29811,N_29066);
nand UO_2677 (O_2677,N_29233,N_28974);
nand UO_2678 (O_2678,N_29133,N_28754);
xnor UO_2679 (O_2679,N_28519,N_29157);
or UO_2680 (O_2680,N_28836,N_29578);
xor UO_2681 (O_2681,N_28768,N_29268);
xor UO_2682 (O_2682,N_28576,N_29454);
nor UO_2683 (O_2683,N_29806,N_29509);
xnor UO_2684 (O_2684,N_29912,N_28847);
and UO_2685 (O_2685,N_29263,N_28696);
xnor UO_2686 (O_2686,N_29567,N_28573);
and UO_2687 (O_2687,N_29531,N_29841);
nor UO_2688 (O_2688,N_28792,N_29941);
and UO_2689 (O_2689,N_29743,N_29180);
and UO_2690 (O_2690,N_29436,N_29531);
xnor UO_2691 (O_2691,N_28640,N_28815);
and UO_2692 (O_2692,N_29868,N_29027);
nor UO_2693 (O_2693,N_29911,N_29696);
nor UO_2694 (O_2694,N_28578,N_29763);
xor UO_2695 (O_2695,N_28596,N_29491);
or UO_2696 (O_2696,N_29038,N_29021);
nand UO_2697 (O_2697,N_29335,N_28925);
nor UO_2698 (O_2698,N_29423,N_29640);
nor UO_2699 (O_2699,N_28655,N_28847);
and UO_2700 (O_2700,N_29807,N_29380);
xor UO_2701 (O_2701,N_29092,N_28937);
and UO_2702 (O_2702,N_29232,N_29362);
nand UO_2703 (O_2703,N_29038,N_29774);
xnor UO_2704 (O_2704,N_29997,N_29806);
xor UO_2705 (O_2705,N_29955,N_29495);
or UO_2706 (O_2706,N_29140,N_28701);
nor UO_2707 (O_2707,N_28561,N_29514);
nor UO_2708 (O_2708,N_28846,N_29780);
or UO_2709 (O_2709,N_28597,N_29471);
nand UO_2710 (O_2710,N_29966,N_28676);
xnor UO_2711 (O_2711,N_29109,N_29252);
nand UO_2712 (O_2712,N_29498,N_29052);
nor UO_2713 (O_2713,N_29555,N_29471);
nor UO_2714 (O_2714,N_28535,N_29934);
xnor UO_2715 (O_2715,N_28689,N_29239);
or UO_2716 (O_2716,N_29917,N_28606);
nor UO_2717 (O_2717,N_29297,N_29916);
nand UO_2718 (O_2718,N_28947,N_29481);
and UO_2719 (O_2719,N_29753,N_28811);
xnor UO_2720 (O_2720,N_29737,N_29347);
nor UO_2721 (O_2721,N_29786,N_28907);
nor UO_2722 (O_2722,N_29338,N_29549);
xnor UO_2723 (O_2723,N_28783,N_29221);
or UO_2724 (O_2724,N_28514,N_29854);
nor UO_2725 (O_2725,N_28580,N_29463);
nor UO_2726 (O_2726,N_28853,N_28646);
nand UO_2727 (O_2727,N_29219,N_28700);
nand UO_2728 (O_2728,N_28791,N_29283);
or UO_2729 (O_2729,N_28749,N_28745);
nand UO_2730 (O_2730,N_29843,N_28626);
xnor UO_2731 (O_2731,N_29801,N_28734);
or UO_2732 (O_2732,N_28975,N_28864);
and UO_2733 (O_2733,N_29823,N_28845);
nand UO_2734 (O_2734,N_28864,N_29486);
nor UO_2735 (O_2735,N_29711,N_29879);
nand UO_2736 (O_2736,N_29993,N_29075);
xnor UO_2737 (O_2737,N_29269,N_29766);
nand UO_2738 (O_2738,N_29607,N_29108);
and UO_2739 (O_2739,N_29273,N_29965);
xor UO_2740 (O_2740,N_29943,N_29033);
or UO_2741 (O_2741,N_28866,N_29195);
or UO_2742 (O_2742,N_29603,N_28744);
or UO_2743 (O_2743,N_29727,N_28775);
xor UO_2744 (O_2744,N_28784,N_29897);
nor UO_2745 (O_2745,N_29995,N_29901);
nor UO_2746 (O_2746,N_29801,N_29695);
xnor UO_2747 (O_2747,N_28570,N_29203);
nand UO_2748 (O_2748,N_28559,N_28593);
xor UO_2749 (O_2749,N_28747,N_29362);
nor UO_2750 (O_2750,N_28573,N_28996);
xor UO_2751 (O_2751,N_29450,N_28836);
and UO_2752 (O_2752,N_28563,N_29482);
nor UO_2753 (O_2753,N_29237,N_29995);
or UO_2754 (O_2754,N_29238,N_29142);
nand UO_2755 (O_2755,N_29072,N_28935);
xnor UO_2756 (O_2756,N_28567,N_28615);
nand UO_2757 (O_2757,N_28586,N_28658);
nor UO_2758 (O_2758,N_28920,N_29630);
nor UO_2759 (O_2759,N_28564,N_29541);
xor UO_2760 (O_2760,N_29777,N_28647);
or UO_2761 (O_2761,N_28533,N_29502);
nor UO_2762 (O_2762,N_29061,N_28920);
and UO_2763 (O_2763,N_29026,N_29456);
nand UO_2764 (O_2764,N_29663,N_28574);
xnor UO_2765 (O_2765,N_29675,N_29678);
nand UO_2766 (O_2766,N_28618,N_29478);
nor UO_2767 (O_2767,N_28708,N_29085);
or UO_2768 (O_2768,N_29404,N_29418);
or UO_2769 (O_2769,N_29230,N_29695);
and UO_2770 (O_2770,N_29052,N_29467);
and UO_2771 (O_2771,N_29788,N_29790);
xnor UO_2772 (O_2772,N_29591,N_29315);
and UO_2773 (O_2773,N_29544,N_29011);
xor UO_2774 (O_2774,N_29059,N_29349);
nand UO_2775 (O_2775,N_29546,N_28845);
nor UO_2776 (O_2776,N_28629,N_28659);
or UO_2777 (O_2777,N_29957,N_29119);
xnor UO_2778 (O_2778,N_29335,N_29153);
nand UO_2779 (O_2779,N_29472,N_29817);
xor UO_2780 (O_2780,N_29263,N_29182);
and UO_2781 (O_2781,N_28752,N_29402);
and UO_2782 (O_2782,N_29597,N_28565);
xnor UO_2783 (O_2783,N_29314,N_29894);
nand UO_2784 (O_2784,N_29513,N_28996);
or UO_2785 (O_2785,N_29484,N_28911);
xor UO_2786 (O_2786,N_29485,N_29218);
nand UO_2787 (O_2787,N_29850,N_29855);
xnor UO_2788 (O_2788,N_29870,N_29341);
and UO_2789 (O_2789,N_29959,N_28780);
or UO_2790 (O_2790,N_29738,N_28677);
nand UO_2791 (O_2791,N_29757,N_29438);
xnor UO_2792 (O_2792,N_29522,N_28752);
and UO_2793 (O_2793,N_29522,N_29157);
xor UO_2794 (O_2794,N_29621,N_29239);
and UO_2795 (O_2795,N_29559,N_29517);
nand UO_2796 (O_2796,N_28511,N_29338);
nand UO_2797 (O_2797,N_29893,N_29960);
or UO_2798 (O_2798,N_28805,N_28975);
or UO_2799 (O_2799,N_29060,N_29566);
or UO_2800 (O_2800,N_28596,N_29051);
nand UO_2801 (O_2801,N_29202,N_29987);
and UO_2802 (O_2802,N_29808,N_29801);
and UO_2803 (O_2803,N_29657,N_29495);
and UO_2804 (O_2804,N_29102,N_29725);
and UO_2805 (O_2805,N_28803,N_29901);
and UO_2806 (O_2806,N_29025,N_29023);
or UO_2807 (O_2807,N_28607,N_29604);
nand UO_2808 (O_2808,N_29676,N_29812);
nor UO_2809 (O_2809,N_28690,N_29436);
nor UO_2810 (O_2810,N_29376,N_29061);
nand UO_2811 (O_2811,N_28802,N_29725);
or UO_2812 (O_2812,N_29260,N_28583);
xnor UO_2813 (O_2813,N_29535,N_28715);
or UO_2814 (O_2814,N_28604,N_29278);
nor UO_2815 (O_2815,N_28860,N_28571);
xor UO_2816 (O_2816,N_28598,N_29374);
or UO_2817 (O_2817,N_29218,N_29939);
and UO_2818 (O_2818,N_28853,N_28881);
or UO_2819 (O_2819,N_29681,N_29207);
nand UO_2820 (O_2820,N_28554,N_29560);
nor UO_2821 (O_2821,N_29509,N_29869);
and UO_2822 (O_2822,N_28512,N_29613);
nand UO_2823 (O_2823,N_29316,N_28786);
nor UO_2824 (O_2824,N_28916,N_28964);
xor UO_2825 (O_2825,N_29831,N_28968);
or UO_2826 (O_2826,N_28648,N_28776);
or UO_2827 (O_2827,N_28730,N_28543);
and UO_2828 (O_2828,N_29551,N_29018);
nor UO_2829 (O_2829,N_28548,N_29494);
and UO_2830 (O_2830,N_29640,N_29031);
xnor UO_2831 (O_2831,N_28597,N_29320);
or UO_2832 (O_2832,N_28843,N_29846);
xor UO_2833 (O_2833,N_29605,N_29259);
nor UO_2834 (O_2834,N_29518,N_29130);
nor UO_2835 (O_2835,N_28807,N_29885);
and UO_2836 (O_2836,N_29848,N_29236);
nand UO_2837 (O_2837,N_28940,N_29310);
nand UO_2838 (O_2838,N_29695,N_28872);
nand UO_2839 (O_2839,N_29970,N_29659);
nand UO_2840 (O_2840,N_28595,N_29950);
or UO_2841 (O_2841,N_29461,N_29045);
xnor UO_2842 (O_2842,N_29741,N_29890);
nor UO_2843 (O_2843,N_28910,N_29659);
nand UO_2844 (O_2844,N_28997,N_29825);
nor UO_2845 (O_2845,N_29481,N_29165);
nor UO_2846 (O_2846,N_29572,N_29372);
nor UO_2847 (O_2847,N_29432,N_29142);
xor UO_2848 (O_2848,N_29478,N_29467);
nor UO_2849 (O_2849,N_28788,N_29986);
and UO_2850 (O_2850,N_28501,N_29446);
or UO_2851 (O_2851,N_29928,N_29796);
nand UO_2852 (O_2852,N_28698,N_28627);
and UO_2853 (O_2853,N_29335,N_29271);
nor UO_2854 (O_2854,N_29598,N_29014);
and UO_2855 (O_2855,N_29593,N_29870);
nand UO_2856 (O_2856,N_29487,N_29615);
xor UO_2857 (O_2857,N_28792,N_29066);
nand UO_2858 (O_2858,N_28688,N_29544);
nand UO_2859 (O_2859,N_29976,N_29811);
nor UO_2860 (O_2860,N_29311,N_29423);
xor UO_2861 (O_2861,N_28587,N_28510);
nor UO_2862 (O_2862,N_29395,N_28705);
nand UO_2863 (O_2863,N_29119,N_29224);
and UO_2864 (O_2864,N_29324,N_29960);
nand UO_2865 (O_2865,N_28532,N_29528);
nor UO_2866 (O_2866,N_29607,N_28984);
xnor UO_2867 (O_2867,N_29786,N_29012);
xnor UO_2868 (O_2868,N_29934,N_29817);
nor UO_2869 (O_2869,N_28604,N_29615);
xnor UO_2870 (O_2870,N_29427,N_29798);
or UO_2871 (O_2871,N_29541,N_29989);
xnor UO_2872 (O_2872,N_29316,N_29655);
and UO_2873 (O_2873,N_29675,N_28913);
nor UO_2874 (O_2874,N_29034,N_29624);
xnor UO_2875 (O_2875,N_29154,N_28884);
nand UO_2876 (O_2876,N_28804,N_29687);
and UO_2877 (O_2877,N_28890,N_29691);
nand UO_2878 (O_2878,N_29383,N_29261);
or UO_2879 (O_2879,N_29749,N_29538);
xnor UO_2880 (O_2880,N_28625,N_29366);
xnor UO_2881 (O_2881,N_28522,N_29828);
nor UO_2882 (O_2882,N_28846,N_29712);
or UO_2883 (O_2883,N_28929,N_28952);
nor UO_2884 (O_2884,N_28748,N_28658);
and UO_2885 (O_2885,N_28846,N_29533);
or UO_2886 (O_2886,N_29340,N_29024);
xnor UO_2887 (O_2887,N_29520,N_28633);
and UO_2888 (O_2888,N_29575,N_29816);
or UO_2889 (O_2889,N_28611,N_29107);
nand UO_2890 (O_2890,N_29927,N_29047);
xor UO_2891 (O_2891,N_29388,N_28912);
or UO_2892 (O_2892,N_29262,N_29873);
and UO_2893 (O_2893,N_29902,N_29547);
or UO_2894 (O_2894,N_28759,N_28629);
or UO_2895 (O_2895,N_29124,N_29225);
nand UO_2896 (O_2896,N_28563,N_28675);
nand UO_2897 (O_2897,N_29601,N_29619);
or UO_2898 (O_2898,N_29073,N_29395);
nand UO_2899 (O_2899,N_28761,N_29517);
and UO_2900 (O_2900,N_28502,N_29206);
or UO_2901 (O_2901,N_29795,N_29054);
nand UO_2902 (O_2902,N_28874,N_28698);
nand UO_2903 (O_2903,N_29520,N_29357);
xor UO_2904 (O_2904,N_28966,N_29855);
xnor UO_2905 (O_2905,N_29725,N_29072);
xnor UO_2906 (O_2906,N_29113,N_29876);
xnor UO_2907 (O_2907,N_28926,N_29906);
nand UO_2908 (O_2908,N_28837,N_29900);
nor UO_2909 (O_2909,N_29539,N_29610);
nor UO_2910 (O_2910,N_29557,N_29802);
nand UO_2911 (O_2911,N_29829,N_28564);
or UO_2912 (O_2912,N_29535,N_29516);
or UO_2913 (O_2913,N_29055,N_29889);
and UO_2914 (O_2914,N_28697,N_28527);
or UO_2915 (O_2915,N_29535,N_29188);
nor UO_2916 (O_2916,N_29449,N_29081);
and UO_2917 (O_2917,N_29079,N_29551);
xor UO_2918 (O_2918,N_29622,N_28968);
or UO_2919 (O_2919,N_28755,N_29927);
nor UO_2920 (O_2920,N_29761,N_29376);
xnor UO_2921 (O_2921,N_29130,N_29610);
or UO_2922 (O_2922,N_28636,N_29002);
or UO_2923 (O_2923,N_28819,N_29957);
or UO_2924 (O_2924,N_28952,N_28685);
and UO_2925 (O_2925,N_29729,N_29179);
or UO_2926 (O_2926,N_29296,N_29399);
nor UO_2927 (O_2927,N_29556,N_29781);
nand UO_2928 (O_2928,N_28773,N_29445);
xnor UO_2929 (O_2929,N_29084,N_29523);
nand UO_2930 (O_2930,N_29091,N_28658);
xor UO_2931 (O_2931,N_29110,N_28839);
nand UO_2932 (O_2932,N_29000,N_29163);
xor UO_2933 (O_2933,N_29146,N_29025);
nand UO_2934 (O_2934,N_28543,N_28659);
and UO_2935 (O_2935,N_29052,N_28989);
xor UO_2936 (O_2936,N_28891,N_29672);
nand UO_2937 (O_2937,N_28502,N_29149);
nand UO_2938 (O_2938,N_29643,N_29395);
xnor UO_2939 (O_2939,N_28525,N_28826);
nand UO_2940 (O_2940,N_29638,N_28923);
or UO_2941 (O_2941,N_29283,N_28529);
xor UO_2942 (O_2942,N_29763,N_28623);
and UO_2943 (O_2943,N_29536,N_28545);
or UO_2944 (O_2944,N_28555,N_28601);
and UO_2945 (O_2945,N_28933,N_29191);
nor UO_2946 (O_2946,N_29856,N_29658);
and UO_2947 (O_2947,N_29604,N_28940);
and UO_2948 (O_2948,N_29877,N_29286);
xnor UO_2949 (O_2949,N_29814,N_28959);
xnor UO_2950 (O_2950,N_28967,N_28952);
nand UO_2951 (O_2951,N_29330,N_29838);
or UO_2952 (O_2952,N_29431,N_29617);
xnor UO_2953 (O_2953,N_29182,N_29383);
or UO_2954 (O_2954,N_28741,N_29962);
xnor UO_2955 (O_2955,N_29077,N_29057);
or UO_2956 (O_2956,N_28617,N_28754);
xor UO_2957 (O_2957,N_28533,N_29948);
nor UO_2958 (O_2958,N_29247,N_29552);
xnor UO_2959 (O_2959,N_28747,N_29448);
xnor UO_2960 (O_2960,N_29895,N_29211);
or UO_2961 (O_2961,N_28727,N_29004);
or UO_2962 (O_2962,N_28982,N_29100);
nor UO_2963 (O_2963,N_29837,N_29548);
nor UO_2964 (O_2964,N_29798,N_29669);
or UO_2965 (O_2965,N_28853,N_29770);
and UO_2966 (O_2966,N_28880,N_29985);
nand UO_2967 (O_2967,N_29480,N_28655);
nor UO_2968 (O_2968,N_28628,N_28738);
nor UO_2969 (O_2969,N_28573,N_29221);
xor UO_2970 (O_2970,N_29222,N_29312);
or UO_2971 (O_2971,N_29378,N_29909);
xor UO_2972 (O_2972,N_29384,N_29579);
xor UO_2973 (O_2973,N_28961,N_29096);
or UO_2974 (O_2974,N_29760,N_29004);
nor UO_2975 (O_2975,N_29751,N_28980);
nand UO_2976 (O_2976,N_29249,N_29979);
or UO_2977 (O_2977,N_28751,N_29930);
and UO_2978 (O_2978,N_29383,N_28973);
nand UO_2979 (O_2979,N_29346,N_28556);
or UO_2980 (O_2980,N_29274,N_28880);
nor UO_2981 (O_2981,N_29090,N_29853);
xnor UO_2982 (O_2982,N_28955,N_29693);
and UO_2983 (O_2983,N_29078,N_29784);
nand UO_2984 (O_2984,N_29224,N_28785);
and UO_2985 (O_2985,N_28977,N_28781);
nand UO_2986 (O_2986,N_29800,N_29767);
nand UO_2987 (O_2987,N_29115,N_28806);
nor UO_2988 (O_2988,N_29889,N_28686);
and UO_2989 (O_2989,N_29380,N_29632);
xnor UO_2990 (O_2990,N_28849,N_28598);
and UO_2991 (O_2991,N_29466,N_29953);
and UO_2992 (O_2992,N_29330,N_29944);
nor UO_2993 (O_2993,N_29840,N_28714);
xnor UO_2994 (O_2994,N_29871,N_28600);
or UO_2995 (O_2995,N_28766,N_28883);
nor UO_2996 (O_2996,N_29206,N_29624);
or UO_2997 (O_2997,N_29607,N_28800);
and UO_2998 (O_2998,N_28935,N_29736);
or UO_2999 (O_2999,N_29674,N_28505);
xnor UO_3000 (O_3000,N_28606,N_29001);
nor UO_3001 (O_3001,N_29533,N_28805);
or UO_3002 (O_3002,N_29756,N_28651);
or UO_3003 (O_3003,N_28871,N_29765);
nor UO_3004 (O_3004,N_28511,N_29029);
and UO_3005 (O_3005,N_29576,N_28584);
and UO_3006 (O_3006,N_28586,N_29364);
and UO_3007 (O_3007,N_28738,N_29934);
xnor UO_3008 (O_3008,N_29755,N_29301);
xnor UO_3009 (O_3009,N_28553,N_28917);
and UO_3010 (O_3010,N_28745,N_29983);
and UO_3011 (O_3011,N_29665,N_29602);
or UO_3012 (O_3012,N_29830,N_28840);
xor UO_3013 (O_3013,N_29806,N_28931);
or UO_3014 (O_3014,N_29238,N_28674);
nand UO_3015 (O_3015,N_29705,N_29409);
nor UO_3016 (O_3016,N_29311,N_29046);
or UO_3017 (O_3017,N_29991,N_28817);
and UO_3018 (O_3018,N_29948,N_29755);
or UO_3019 (O_3019,N_29946,N_29323);
or UO_3020 (O_3020,N_29285,N_28633);
and UO_3021 (O_3021,N_28843,N_29886);
or UO_3022 (O_3022,N_29074,N_29962);
nor UO_3023 (O_3023,N_29083,N_29948);
and UO_3024 (O_3024,N_29475,N_29003);
nand UO_3025 (O_3025,N_29058,N_29250);
nand UO_3026 (O_3026,N_29729,N_29114);
and UO_3027 (O_3027,N_28652,N_29135);
xnor UO_3028 (O_3028,N_28611,N_28625);
and UO_3029 (O_3029,N_29199,N_29341);
and UO_3030 (O_3030,N_29154,N_29999);
xnor UO_3031 (O_3031,N_29971,N_29450);
xnor UO_3032 (O_3032,N_29696,N_29445);
nand UO_3033 (O_3033,N_29401,N_28552);
nor UO_3034 (O_3034,N_29351,N_28968);
and UO_3035 (O_3035,N_29749,N_28540);
xor UO_3036 (O_3036,N_28816,N_28621);
xor UO_3037 (O_3037,N_28899,N_29488);
and UO_3038 (O_3038,N_29511,N_29405);
xor UO_3039 (O_3039,N_29571,N_29445);
and UO_3040 (O_3040,N_29513,N_29240);
xor UO_3041 (O_3041,N_29542,N_29012);
nand UO_3042 (O_3042,N_28707,N_29105);
nor UO_3043 (O_3043,N_29365,N_28971);
or UO_3044 (O_3044,N_29179,N_28870);
xnor UO_3045 (O_3045,N_29624,N_28949);
or UO_3046 (O_3046,N_29579,N_28657);
and UO_3047 (O_3047,N_28862,N_29795);
nand UO_3048 (O_3048,N_29352,N_29699);
and UO_3049 (O_3049,N_28790,N_28748);
nand UO_3050 (O_3050,N_28565,N_29375);
or UO_3051 (O_3051,N_29738,N_29176);
nor UO_3052 (O_3052,N_28847,N_29886);
nand UO_3053 (O_3053,N_29593,N_29227);
xnor UO_3054 (O_3054,N_29057,N_29716);
nand UO_3055 (O_3055,N_29762,N_29173);
xnor UO_3056 (O_3056,N_28529,N_29540);
and UO_3057 (O_3057,N_28670,N_28613);
nand UO_3058 (O_3058,N_29244,N_29394);
xor UO_3059 (O_3059,N_28958,N_28856);
xnor UO_3060 (O_3060,N_28701,N_29953);
nor UO_3061 (O_3061,N_28769,N_29870);
or UO_3062 (O_3062,N_29993,N_29359);
or UO_3063 (O_3063,N_28945,N_29796);
and UO_3064 (O_3064,N_29897,N_28834);
nand UO_3065 (O_3065,N_28760,N_29109);
or UO_3066 (O_3066,N_29748,N_28903);
and UO_3067 (O_3067,N_29621,N_28616);
nand UO_3068 (O_3068,N_29344,N_28521);
nand UO_3069 (O_3069,N_28550,N_29950);
xor UO_3070 (O_3070,N_29841,N_29857);
nor UO_3071 (O_3071,N_29991,N_29443);
or UO_3072 (O_3072,N_29871,N_29364);
xnor UO_3073 (O_3073,N_29790,N_29750);
nand UO_3074 (O_3074,N_29901,N_28948);
nor UO_3075 (O_3075,N_29485,N_28754);
and UO_3076 (O_3076,N_29409,N_28868);
and UO_3077 (O_3077,N_29729,N_28828);
nand UO_3078 (O_3078,N_28598,N_28603);
or UO_3079 (O_3079,N_29148,N_28793);
nor UO_3080 (O_3080,N_29671,N_29950);
and UO_3081 (O_3081,N_29495,N_28545);
xnor UO_3082 (O_3082,N_29018,N_29452);
and UO_3083 (O_3083,N_28952,N_29410);
xor UO_3084 (O_3084,N_28729,N_29373);
and UO_3085 (O_3085,N_29947,N_29310);
nand UO_3086 (O_3086,N_29689,N_28909);
nor UO_3087 (O_3087,N_29215,N_29723);
and UO_3088 (O_3088,N_29788,N_29845);
nor UO_3089 (O_3089,N_29395,N_28582);
nand UO_3090 (O_3090,N_29260,N_29529);
and UO_3091 (O_3091,N_29464,N_28610);
nand UO_3092 (O_3092,N_28583,N_29122);
nand UO_3093 (O_3093,N_29261,N_28902);
or UO_3094 (O_3094,N_29468,N_29369);
and UO_3095 (O_3095,N_29334,N_29222);
nor UO_3096 (O_3096,N_28620,N_28931);
nand UO_3097 (O_3097,N_29748,N_28741);
nor UO_3098 (O_3098,N_29271,N_28870);
xor UO_3099 (O_3099,N_29812,N_28755);
nor UO_3100 (O_3100,N_28923,N_29599);
and UO_3101 (O_3101,N_28767,N_29953);
nor UO_3102 (O_3102,N_29383,N_28849);
xor UO_3103 (O_3103,N_29729,N_28739);
and UO_3104 (O_3104,N_29140,N_28996);
nand UO_3105 (O_3105,N_28511,N_29653);
nand UO_3106 (O_3106,N_29332,N_29317);
xnor UO_3107 (O_3107,N_28853,N_28868);
nor UO_3108 (O_3108,N_28745,N_29438);
and UO_3109 (O_3109,N_28895,N_28828);
and UO_3110 (O_3110,N_29862,N_29207);
or UO_3111 (O_3111,N_29517,N_29297);
nor UO_3112 (O_3112,N_29350,N_28751);
xnor UO_3113 (O_3113,N_29821,N_29941);
xnor UO_3114 (O_3114,N_29149,N_28505);
nand UO_3115 (O_3115,N_29373,N_29506);
nor UO_3116 (O_3116,N_29313,N_29570);
or UO_3117 (O_3117,N_28817,N_29701);
nor UO_3118 (O_3118,N_29879,N_29166);
xor UO_3119 (O_3119,N_29406,N_29715);
xnor UO_3120 (O_3120,N_29597,N_29843);
nor UO_3121 (O_3121,N_29883,N_28857);
nand UO_3122 (O_3122,N_29391,N_29972);
xnor UO_3123 (O_3123,N_28891,N_29852);
and UO_3124 (O_3124,N_28798,N_29576);
nor UO_3125 (O_3125,N_28659,N_29302);
nor UO_3126 (O_3126,N_29790,N_29696);
xor UO_3127 (O_3127,N_28684,N_28979);
nor UO_3128 (O_3128,N_28916,N_29950);
nor UO_3129 (O_3129,N_29055,N_29945);
xnor UO_3130 (O_3130,N_29483,N_29358);
xnor UO_3131 (O_3131,N_29263,N_29633);
or UO_3132 (O_3132,N_29538,N_28665);
xnor UO_3133 (O_3133,N_29348,N_29043);
and UO_3134 (O_3134,N_29878,N_29374);
nor UO_3135 (O_3135,N_29633,N_29748);
nand UO_3136 (O_3136,N_29582,N_29897);
xor UO_3137 (O_3137,N_29447,N_28543);
or UO_3138 (O_3138,N_29421,N_29668);
or UO_3139 (O_3139,N_29516,N_28774);
xnor UO_3140 (O_3140,N_29989,N_29166);
nor UO_3141 (O_3141,N_29554,N_28623);
or UO_3142 (O_3142,N_28918,N_28522);
and UO_3143 (O_3143,N_29732,N_28923);
nor UO_3144 (O_3144,N_29805,N_29485);
or UO_3145 (O_3145,N_28629,N_29038);
nand UO_3146 (O_3146,N_28891,N_28830);
nand UO_3147 (O_3147,N_29299,N_29261);
or UO_3148 (O_3148,N_28875,N_29499);
xnor UO_3149 (O_3149,N_29702,N_28704);
nand UO_3150 (O_3150,N_29472,N_28694);
or UO_3151 (O_3151,N_28694,N_29933);
xor UO_3152 (O_3152,N_29490,N_29770);
xor UO_3153 (O_3153,N_29827,N_29828);
or UO_3154 (O_3154,N_29360,N_29119);
nor UO_3155 (O_3155,N_29216,N_29894);
nand UO_3156 (O_3156,N_28981,N_28861);
nand UO_3157 (O_3157,N_29744,N_29459);
xor UO_3158 (O_3158,N_29515,N_28531);
xnor UO_3159 (O_3159,N_29040,N_29132);
nand UO_3160 (O_3160,N_28784,N_29350);
nand UO_3161 (O_3161,N_29272,N_29072);
and UO_3162 (O_3162,N_29689,N_28972);
or UO_3163 (O_3163,N_28773,N_28802);
or UO_3164 (O_3164,N_28642,N_29308);
and UO_3165 (O_3165,N_28820,N_29400);
or UO_3166 (O_3166,N_29971,N_29592);
nand UO_3167 (O_3167,N_29303,N_29305);
nor UO_3168 (O_3168,N_28983,N_28540);
and UO_3169 (O_3169,N_28878,N_29018);
xor UO_3170 (O_3170,N_28779,N_29155);
and UO_3171 (O_3171,N_28733,N_28746);
nor UO_3172 (O_3172,N_29453,N_29932);
xor UO_3173 (O_3173,N_28568,N_29760);
or UO_3174 (O_3174,N_29528,N_29810);
or UO_3175 (O_3175,N_29305,N_29670);
nand UO_3176 (O_3176,N_29616,N_28715);
nand UO_3177 (O_3177,N_28960,N_29692);
xor UO_3178 (O_3178,N_29401,N_28579);
or UO_3179 (O_3179,N_29152,N_29773);
and UO_3180 (O_3180,N_28528,N_29874);
nor UO_3181 (O_3181,N_29812,N_29919);
nand UO_3182 (O_3182,N_29333,N_29189);
nand UO_3183 (O_3183,N_29438,N_29779);
nor UO_3184 (O_3184,N_29402,N_28850);
and UO_3185 (O_3185,N_29419,N_29354);
nor UO_3186 (O_3186,N_29099,N_29703);
and UO_3187 (O_3187,N_29355,N_29664);
or UO_3188 (O_3188,N_29877,N_28661);
or UO_3189 (O_3189,N_29694,N_28565);
xnor UO_3190 (O_3190,N_28921,N_29351);
and UO_3191 (O_3191,N_29077,N_28970);
and UO_3192 (O_3192,N_29278,N_29521);
or UO_3193 (O_3193,N_29643,N_28737);
xnor UO_3194 (O_3194,N_28919,N_28678);
nor UO_3195 (O_3195,N_29564,N_29605);
xor UO_3196 (O_3196,N_28592,N_28808);
and UO_3197 (O_3197,N_29505,N_29945);
nor UO_3198 (O_3198,N_29258,N_29573);
xor UO_3199 (O_3199,N_28697,N_29524);
nand UO_3200 (O_3200,N_29354,N_28871);
xor UO_3201 (O_3201,N_29885,N_28566);
xor UO_3202 (O_3202,N_29305,N_29012);
xor UO_3203 (O_3203,N_29312,N_28751);
or UO_3204 (O_3204,N_29832,N_29834);
nand UO_3205 (O_3205,N_29253,N_29382);
xor UO_3206 (O_3206,N_29309,N_29374);
xnor UO_3207 (O_3207,N_29515,N_29506);
nand UO_3208 (O_3208,N_28705,N_28877);
xnor UO_3209 (O_3209,N_28771,N_28544);
nand UO_3210 (O_3210,N_29480,N_29335);
and UO_3211 (O_3211,N_29451,N_29209);
nand UO_3212 (O_3212,N_28603,N_29529);
xor UO_3213 (O_3213,N_28923,N_29182);
or UO_3214 (O_3214,N_28839,N_29211);
xnor UO_3215 (O_3215,N_28686,N_29126);
xor UO_3216 (O_3216,N_29473,N_29606);
nor UO_3217 (O_3217,N_29356,N_28614);
nor UO_3218 (O_3218,N_28948,N_29777);
or UO_3219 (O_3219,N_29634,N_28601);
nand UO_3220 (O_3220,N_28518,N_28616);
or UO_3221 (O_3221,N_29020,N_29506);
xnor UO_3222 (O_3222,N_29525,N_29722);
nand UO_3223 (O_3223,N_29014,N_28719);
or UO_3224 (O_3224,N_29380,N_29808);
or UO_3225 (O_3225,N_29794,N_29768);
nand UO_3226 (O_3226,N_28713,N_29065);
or UO_3227 (O_3227,N_29401,N_29970);
nand UO_3228 (O_3228,N_28985,N_28826);
xnor UO_3229 (O_3229,N_29989,N_28694);
or UO_3230 (O_3230,N_29313,N_29277);
and UO_3231 (O_3231,N_29229,N_28873);
nand UO_3232 (O_3232,N_29893,N_29565);
or UO_3233 (O_3233,N_28616,N_28679);
xnor UO_3234 (O_3234,N_29029,N_29753);
or UO_3235 (O_3235,N_29511,N_29077);
or UO_3236 (O_3236,N_29089,N_28672);
and UO_3237 (O_3237,N_29313,N_29987);
or UO_3238 (O_3238,N_28612,N_29250);
or UO_3239 (O_3239,N_29536,N_29807);
nor UO_3240 (O_3240,N_29299,N_29367);
or UO_3241 (O_3241,N_29842,N_29627);
and UO_3242 (O_3242,N_29268,N_28752);
and UO_3243 (O_3243,N_29436,N_29070);
xnor UO_3244 (O_3244,N_29280,N_28936);
xor UO_3245 (O_3245,N_29413,N_29561);
nor UO_3246 (O_3246,N_28753,N_28957);
and UO_3247 (O_3247,N_28543,N_29973);
xnor UO_3248 (O_3248,N_29259,N_29621);
nand UO_3249 (O_3249,N_29285,N_29081);
nor UO_3250 (O_3250,N_29076,N_29977);
nand UO_3251 (O_3251,N_29449,N_29403);
nand UO_3252 (O_3252,N_29493,N_29325);
or UO_3253 (O_3253,N_29077,N_29937);
or UO_3254 (O_3254,N_29083,N_29233);
nor UO_3255 (O_3255,N_28737,N_29347);
nor UO_3256 (O_3256,N_29330,N_28766);
nand UO_3257 (O_3257,N_28876,N_29353);
or UO_3258 (O_3258,N_28817,N_28867);
nand UO_3259 (O_3259,N_28654,N_28662);
nand UO_3260 (O_3260,N_28505,N_29946);
and UO_3261 (O_3261,N_28960,N_29915);
nand UO_3262 (O_3262,N_29331,N_28807);
or UO_3263 (O_3263,N_29193,N_28639);
nor UO_3264 (O_3264,N_28759,N_29237);
or UO_3265 (O_3265,N_28577,N_29294);
and UO_3266 (O_3266,N_29836,N_29819);
and UO_3267 (O_3267,N_29814,N_29001);
xor UO_3268 (O_3268,N_29922,N_29007);
nor UO_3269 (O_3269,N_28607,N_29084);
or UO_3270 (O_3270,N_29631,N_28807);
and UO_3271 (O_3271,N_29748,N_29458);
and UO_3272 (O_3272,N_28513,N_29913);
and UO_3273 (O_3273,N_29478,N_28911);
nor UO_3274 (O_3274,N_29179,N_29580);
or UO_3275 (O_3275,N_29068,N_29591);
xnor UO_3276 (O_3276,N_28931,N_29020);
nand UO_3277 (O_3277,N_29851,N_29126);
nor UO_3278 (O_3278,N_28634,N_28599);
or UO_3279 (O_3279,N_29591,N_28615);
xnor UO_3280 (O_3280,N_28746,N_29064);
nand UO_3281 (O_3281,N_29214,N_28828);
nand UO_3282 (O_3282,N_29325,N_28509);
xor UO_3283 (O_3283,N_29314,N_28599);
nor UO_3284 (O_3284,N_29006,N_29632);
or UO_3285 (O_3285,N_28891,N_28955);
xnor UO_3286 (O_3286,N_29795,N_28979);
or UO_3287 (O_3287,N_29409,N_28612);
xor UO_3288 (O_3288,N_29327,N_29740);
or UO_3289 (O_3289,N_29662,N_28648);
or UO_3290 (O_3290,N_29333,N_29859);
nand UO_3291 (O_3291,N_29723,N_29639);
xnor UO_3292 (O_3292,N_28502,N_29003);
nand UO_3293 (O_3293,N_29774,N_29083);
nand UO_3294 (O_3294,N_29532,N_29851);
nand UO_3295 (O_3295,N_29042,N_29201);
or UO_3296 (O_3296,N_28980,N_29371);
nand UO_3297 (O_3297,N_28798,N_29240);
xor UO_3298 (O_3298,N_29500,N_28686);
xor UO_3299 (O_3299,N_29234,N_29070);
or UO_3300 (O_3300,N_28846,N_29454);
or UO_3301 (O_3301,N_29457,N_28629);
nor UO_3302 (O_3302,N_29430,N_29420);
nor UO_3303 (O_3303,N_28596,N_29621);
or UO_3304 (O_3304,N_28548,N_28654);
and UO_3305 (O_3305,N_29444,N_28638);
xor UO_3306 (O_3306,N_29145,N_29074);
nor UO_3307 (O_3307,N_29362,N_29179);
xnor UO_3308 (O_3308,N_29999,N_28773);
nor UO_3309 (O_3309,N_28682,N_29751);
nand UO_3310 (O_3310,N_29804,N_28755);
and UO_3311 (O_3311,N_29451,N_29485);
or UO_3312 (O_3312,N_29851,N_29378);
and UO_3313 (O_3313,N_28902,N_29485);
xor UO_3314 (O_3314,N_29036,N_29171);
or UO_3315 (O_3315,N_28516,N_29460);
and UO_3316 (O_3316,N_28662,N_29776);
nor UO_3317 (O_3317,N_29444,N_29171);
nand UO_3318 (O_3318,N_29626,N_29985);
nand UO_3319 (O_3319,N_29600,N_29135);
nor UO_3320 (O_3320,N_29589,N_28686);
nor UO_3321 (O_3321,N_29347,N_29657);
and UO_3322 (O_3322,N_29391,N_29158);
xnor UO_3323 (O_3323,N_29694,N_29674);
nand UO_3324 (O_3324,N_28640,N_29775);
and UO_3325 (O_3325,N_28657,N_28685);
nor UO_3326 (O_3326,N_28785,N_28618);
nand UO_3327 (O_3327,N_29236,N_29216);
nand UO_3328 (O_3328,N_28848,N_28637);
nor UO_3329 (O_3329,N_29884,N_29424);
and UO_3330 (O_3330,N_28839,N_28717);
xnor UO_3331 (O_3331,N_29451,N_29933);
nor UO_3332 (O_3332,N_29439,N_28683);
or UO_3333 (O_3333,N_29945,N_29229);
xnor UO_3334 (O_3334,N_28899,N_29051);
xnor UO_3335 (O_3335,N_29171,N_29608);
nand UO_3336 (O_3336,N_29475,N_29243);
nand UO_3337 (O_3337,N_29172,N_29272);
and UO_3338 (O_3338,N_29819,N_29132);
and UO_3339 (O_3339,N_28904,N_29909);
and UO_3340 (O_3340,N_29287,N_29992);
or UO_3341 (O_3341,N_29670,N_29599);
and UO_3342 (O_3342,N_29395,N_29341);
nor UO_3343 (O_3343,N_28624,N_28963);
and UO_3344 (O_3344,N_29388,N_28519);
nor UO_3345 (O_3345,N_28935,N_29332);
or UO_3346 (O_3346,N_29308,N_29903);
nand UO_3347 (O_3347,N_28567,N_29000);
and UO_3348 (O_3348,N_29950,N_29467);
and UO_3349 (O_3349,N_28505,N_29458);
or UO_3350 (O_3350,N_29964,N_28624);
or UO_3351 (O_3351,N_29637,N_28673);
or UO_3352 (O_3352,N_28930,N_28779);
nor UO_3353 (O_3353,N_28711,N_29840);
or UO_3354 (O_3354,N_29117,N_29949);
and UO_3355 (O_3355,N_29844,N_28730);
or UO_3356 (O_3356,N_29780,N_29771);
nor UO_3357 (O_3357,N_29571,N_28976);
nor UO_3358 (O_3358,N_29465,N_28570);
nor UO_3359 (O_3359,N_28937,N_29748);
nand UO_3360 (O_3360,N_29108,N_29530);
nor UO_3361 (O_3361,N_29034,N_29963);
nor UO_3362 (O_3362,N_28747,N_28610);
nand UO_3363 (O_3363,N_28728,N_28819);
or UO_3364 (O_3364,N_28977,N_29313);
nor UO_3365 (O_3365,N_29236,N_29075);
nor UO_3366 (O_3366,N_29908,N_29999);
and UO_3367 (O_3367,N_29388,N_28599);
nand UO_3368 (O_3368,N_28828,N_29424);
nand UO_3369 (O_3369,N_29216,N_29126);
nand UO_3370 (O_3370,N_28673,N_29091);
or UO_3371 (O_3371,N_29228,N_29080);
nor UO_3372 (O_3372,N_28784,N_28860);
xnor UO_3373 (O_3373,N_29485,N_29132);
nor UO_3374 (O_3374,N_29713,N_28673);
or UO_3375 (O_3375,N_29729,N_28773);
or UO_3376 (O_3376,N_29672,N_28739);
or UO_3377 (O_3377,N_28741,N_29092);
and UO_3378 (O_3378,N_29061,N_28641);
nand UO_3379 (O_3379,N_28672,N_29461);
xnor UO_3380 (O_3380,N_28815,N_29138);
nor UO_3381 (O_3381,N_29254,N_29210);
xor UO_3382 (O_3382,N_28553,N_29288);
or UO_3383 (O_3383,N_29736,N_29431);
nor UO_3384 (O_3384,N_29974,N_29549);
nand UO_3385 (O_3385,N_29092,N_29858);
nor UO_3386 (O_3386,N_28600,N_29167);
and UO_3387 (O_3387,N_29572,N_29354);
nor UO_3388 (O_3388,N_29572,N_29730);
nor UO_3389 (O_3389,N_29418,N_28958);
nand UO_3390 (O_3390,N_28889,N_29036);
and UO_3391 (O_3391,N_29679,N_29771);
nor UO_3392 (O_3392,N_29866,N_29347);
and UO_3393 (O_3393,N_29559,N_29531);
and UO_3394 (O_3394,N_29460,N_29704);
or UO_3395 (O_3395,N_28856,N_29524);
nand UO_3396 (O_3396,N_29468,N_28524);
and UO_3397 (O_3397,N_28769,N_29161);
nor UO_3398 (O_3398,N_28554,N_28713);
and UO_3399 (O_3399,N_29231,N_28523);
and UO_3400 (O_3400,N_28630,N_28970);
nand UO_3401 (O_3401,N_29805,N_28594);
nand UO_3402 (O_3402,N_29836,N_29174);
or UO_3403 (O_3403,N_29217,N_29492);
and UO_3404 (O_3404,N_29621,N_28940);
xor UO_3405 (O_3405,N_28788,N_28863);
or UO_3406 (O_3406,N_29843,N_29221);
or UO_3407 (O_3407,N_28528,N_29437);
nand UO_3408 (O_3408,N_28669,N_28722);
or UO_3409 (O_3409,N_29099,N_28981);
or UO_3410 (O_3410,N_29128,N_29509);
nand UO_3411 (O_3411,N_29748,N_28848);
xnor UO_3412 (O_3412,N_29331,N_28743);
nor UO_3413 (O_3413,N_29997,N_29127);
or UO_3414 (O_3414,N_29047,N_29285);
or UO_3415 (O_3415,N_29770,N_29631);
or UO_3416 (O_3416,N_29829,N_29434);
and UO_3417 (O_3417,N_29206,N_29679);
nor UO_3418 (O_3418,N_28654,N_29259);
nand UO_3419 (O_3419,N_29077,N_28596);
nor UO_3420 (O_3420,N_29948,N_28800);
nor UO_3421 (O_3421,N_29483,N_29849);
nand UO_3422 (O_3422,N_28771,N_29155);
nand UO_3423 (O_3423,N_29734,N_29674);
or UO_3424 (O_3424,N_29533,N_28972);
or UO_3425 (O_3425,N_29363,N_29933);
nand UO_3426 (O_3426,N_28610,N_29951);
xor UO_3427 (O_3427,N_29246,N_28608);
xor UO_3428 (O_3428,N_29120,N_28698);
and UO_3429 (O_3429,N_28821,N_29860);
nand UO_3430 (O_3430,N_28875,N_29338);
nand UO_3431 (O_3431,N_28644,N_28986);
or UO_3432 (O_3432,N_28675,N_29730);
and UO_3433 (O_3433,N_28752,N_28557);
nor UO_3434 (O_3434,N_28669,N_28984);
and UO_3435 (O_3435,N_29782,N_29415);
nor UO_3436 (O_3436,N_29626,N_29400);
xnor UO_3437 (O_3437,N_28515,N_29118);
nand UO_3438 (O_3438,N_29097,N_29223);
and UO_3439 (O_3439,N_28937,N_29336);
nand UO_3440 (O_3440,N_29802,N_29204);
nor UO_3441 (O_3441,N_28804,N_29150);
and UO_3442 (O_3442,N_29409,N_29060);
xor UO_3443 (O_3443,N_28774,N_29538);
nor UO_3444 (O_3444,N_29545,N_29073);
xnor UO_3445 (O_3445,N_29511,N_28730);
and UO_3446 (O_3446,N_29931,N_29655);
or UO_3447 (O_3447,N_29086,N_28686);
nor UO_3448 (O_3448,N_28840,N_28609);
xnor UO_3449 (O_3449,N_29536,N_28786);
nand UO_3450 (O_3450,N_28637,N_28972);
or UO_3451 (O_3451,N_29139,N_29735);
xnor UO_3452 (O_3452,N_29063,N_29675);
nor UO_3453 (O_3453,N_29401,N_28699);
nor UO_3454 (O_3454,N_28646,N_29242);
nand UO_3455 (O_3455,N_28783,N_29201);
or UO_3456 (O_3456,N_29057,N_28681);
or UO_3457 (O_3457,N_28923,N_29559);
and UO_3458 (O_3458,N_29146,N_29730);
xor UO_3459 (O_3459,N_29840,N_28843);
and UO_3460 (O_3460,N_28595,N_29962);
nor UO_3461 (O_3461,N_29064,N_29229);
or UO_3462 (O_3462,N_28631,N_29888);
xnor UO_3463 (O_3463,N_29175,N_29178);
xor UO_3464 (O_3464,N_29717,N_29153);
or UO_3465 (O_3465,N_29784,N_29140);
and UO_3466 (O_3466,N_29989,N_29191);
nand UO_3467 (O_3467,N_29435,N_28709);
or UO_3468 (O_3468,N_29214,N_29810);
xor UO_3469 (O_3469,N_29043,N_28744);
xor UO_3470 (O_3470,N_29952,N_29595);
nor UO_3471 (O_3471,N_29927,N_28994);
nand UO_3472 (O_3472,N_29603,N_28947);
nor UO_3473 (O_3473,N_28828,N_29639);
and UO_3474 (O_3474,N_29360,N_29669);
and UO_3475 (O_3475,N_29610,N_29136);
nand UO_3476 (O_3476,N_29295,N_28614);
or UO_3477 (O_3477,N_29930,N_29070);
and UO_3478 (O_3478,N_29831,N_29148);
nand UO_3479 (O_3479,N_29704,N_28565);
or UO_3480 (O_3480,N_29813,N_29323);
nand UO_3481 (O_3481,N_28917,N_29919);
and UO_3482 (O_3482,N_29622,N_28803);
and UO_3483 (O_3483,N_29644,N_29830);
xnor UO_3484 (O_3484,N_29787,N_29934);
nand UO_3485 (O_3485,N_29345,N_28520);
nor UO_3486 (O_3486,N_28520,N_29258);
xnor UO_3487 (O_3487,N_28602,N_29293);
nand UO_3488 (O_3488,N_29409,N_28539);
nor UO_3489 (O_3489,N_28505,N_29490);
nand UO_3490 (O_3490,N_28640,N_29193);
nand UO_3491 (O_3491,N_29719,N_28846);
xnor UO_3492 (O_3492,N_29123,N_29181);
xor UO_3493 (O_3493,N_28759,N_29878);
or UO_3494 (O_3494,N_29355,N_28860);
nand UO_3495 (O_3495,N_29380,N_28503);
xor UO_3496 (O_3496,N_28891,N_29733);
or UO_3497 (O_3497,N_29784,N_29994);
nand UO_3498 (O_3498,N_29045,N_28543);
and UO_3499 (O_3499,N_29414,N_28626);
endmodule