module basic_2000_20000_2500_5_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_593,In_1896);
xor U1 (N_1,In_290,In_1124);
or U2 (N_2,In_1965,In_1482);
nor U3 (N_3,In_1433,In_928);
or U4 (N_4,In_1539,In_1932);
xor U5 (N_5,In_1629,In_1074);
nand U6 (N_6,In_1224,In_1912);
nor U7 (N_7,In_1516,In_1577);
nand U8 (N_8,In_994,In_655);
xor U9 (N_9,In_199,In_883);
nor U10 (N_10,In_367,In_658);
or U11 (N_11,In_87,In_1385);
nor U12 (N_12,In_279,In_1678);
and U13 (N_13,In_784,In_891);
and U14 (N_14,In_445,In_996);
nor U15 (N_15,In_912,In_634);
nand U16 (N_16,In_532,In_1378);
or U17 (N_17,In_288,In_1758);
nor U18 (N_18,In_638,In_519);
and U19 (N_19,In_1493,In_326);
and U20 (N_20,In_599,In_921);
and U21 (N_21,In_1698,In_779);
or U22 (N_22,In_647,In_1807);
nand U23 (N_23,In_1504,In_1809);
nand U24 (N_24,In_535,In_556);
xor U25 (N_25,In_1012,In_464);
nand U26 (N_26,In_569,In_622);
nand U27 (N_27,In_1197,In_366);
xor U28 (N_28,In_1257,In_235);
or U29 (N_29,In_1788,In_160);
nand U30 (N_30,In_1680,In_866);
xor U31 (N_31,In_75,In_377);
nor U32 (N_32,In_1514,In_1507);
xnor U33 (N_33,In_1239,In_678);
nor U34 (N_34,In_713,In_1953);
or U35 (N_35,In_1963,In_938);
and U36 (N_36,In_566,In_1242);
xnor U37 (N_37,In_1112,In_188);
and U38 (N_38,In_1931,In_1861);
nor U39 (N_39,In_1848,In_208);
nand U40 (N_40,In_1043,In_1558);
nand U41 (N_41,In_1110,In_1187);
nor U42 (N_42,In_819,In_1238);
nor U43 (N_43,In_1707,In_1595);
nor U44 (N_44,In_325,In_1997);
or U45 (N_45,In_1284,In_958);
nand U46 (N_46,In_1644,In_1713);
and U47 (N_47,In_344,In_1761);
xnor U48 (N_48,In_1938,In_1515);
nor U49 (N_49,In_969,In_776);
nor U50 (N_50,In_1007,In_1361);
nor U51 (N_51,In_523,In_567);
and U52 (N_52,In_1729,In_1479);
and U53 (N_53,In_1762,In_162);
xor U54 (N_54,In_336,In_9);
nand U55 (N_55,In_330,In_1078);
xor U56 (N_56,In_312,In_861);
or U57 (N_57,In_868,In_792);
nand U58 (N_58,In_474,In_213);
nand U59 (N_59,In_459,In_31);
nor U60 (N_60,In_973,In_251);
nor U61 (N_61,In_1768,In_1153);
xnor U62 (N_62,In_1203,In_796);
xnor U63 (N_63,In_1205,In_1233);
and U64 (N_64,In_21,In_739);
nand U65 (N_65,In_151,In_541);
and U66 (N_66,In_1796,In_942);
xnor U67 (N_67,In_1247,In_730);
and U68 (N_68,In_1827,In_483);
and U69 (N_69,In_1062,In_867);
nor U70 (N_70,In_1534,In_1279);
xnor U71 (N_71,In_129,In_1955);
or U72 (N_72,In_1977,In_153);
nand U73 (N_73,In_1744,In_350);
nor U74 (N_74,In_1402,In_285);
nor U75 (N_75,In_1817,In_494);
and U76 (N_76,In_505,In_1556);
xor U77 (N_77,In_990,In_1119);
or U78 (N_78,In_1494,In_1355);
or U79 (N_79,In_114,In_1142);
nand U80 (N_80,In_1430,In_1008);
nor U81 (N_81,In_1170,In_962);
nand U82 (N_82,In_14,In_1816);
and U83 (N_83,In_1206,In_863);
or U84 (N_84,In_424,In_1683);
and U85 (N_85,In_738,In_1488);
or U86 (N_86,In_1669,In_1199);
and U87 (N_87,In_747,In_578);
xnor U88 (N_88,In_1580,In_499);
or U89 (N_89,In_1612,In_1551);
nor U90 (N_90,In_502,In_1892);
or U91 (N_91,In_1332,In_1312);
xor U92 (N_92,In_1180,In_995);
and U93 (N_93,In_431,In_628);
nor U94 (N_94,In_262,In_1389);
and U95 (N_95,In_753,In_309);
and U96 (N_96,In_763,In_98);
nand U97 (N_97,In_1511,In_138);
or U98 (N_98,In_191,In_358);
xnor U99 (N_99,In_1626,In_1292);
xnor U100 (N_100,In_101,In_793);
nor U101 (N_101,In_1418,In_444);
nand U102 (N_102,In_758,In_313);
or U103 (N_103,In_531,In_1065);
nand U104 (N_104,In_1502,In_1081);
xnor U105 (N_105,In_572,In_1091);
or U106 (N_106,In_1130,In_843);
and U107 (N_107,In_676,In_911);
and U108 (N_108,In_882,In_1277);
nor U109 (N_109,In_828,In_55);
or U110 (N_110,In_415,In_1679);
and U111 (N_111,In_489,In_948);
nor U112 (N_112,In_1020,In_675);
nor U113 (N_113,In_1567,In_1191);
or U114 (N_114,In_605,In_1623);
or U115 (N_115,In_36,In_1675);
xnor U116 (N_116,In_1976,In_1655);
nand U117 (N_117,In_210,In_732);
xnor U118 (N_118,In_301,In_1275);
xnor U119 (N_119,In_60,In_1473);
nor U120 (N_120,In_1631,In_805);
nor U121 (N_121,In_315,In_1523);
nand U122 (N_122,In_546,In_1789);
or U123 (N_123,In_1957,In_1146);
nand U124 (N_124,In_1314,In_910);
or U125 (N_125,In_1177,In_1392);
or U126 (N_126,In_1806,In_1252);
or U127 (N_127,In_660,In_583);
or U128 (N_128,In_1717,In_621);
nor U129 (N_129,In_34,In_1791);
xor U130 (N_130,In_1475,In_937);
nor U131 (N_131,In_1060,In_652);
and U132 (N_132,In_146,In_1540);
nand U133 (N_133,In_29,In_1337);
xnor U134 (N_134,In_349,In_799);
and U135 (N_135,In_1016,In_554);
and U136 (N_136,In_156,In_81);
and U137 (N_137,In_1310,In_832);
nand U138 (N_138,In_611,In_1071);
or U139 (N_139,In_186,In_137);
nor U140 (N_140,In_1015,In_1363);
and U141 (N_141,In_511,In_764);
xnor U142 (N_142,In_694,In_951);
or U143 (N_143,In_1001,In_1244);
nand U144 (N_144,In_1321,In_394);
or U145 (N_145,In_51,In_218);
nand U146 (N_146,In_1625,In_1716);
or U147 (N_147,In_930,In_277);
xor U148 (N_148,In_52,In_573);
xor U149 (N_149,In_1155,In_1921);
xor U150 (N_150,In_1906,In_1525);
and U151 (N_151,In_976,In_47);
and U152 (N_152,In_95,In_968);
nand U153 (N_153,In_723,In_1601);
and U154 (N_154,In_1113,In_636);
and U155 (N_155,In_1111,In_1743);
or U156 (N_156,In_524,In_440);
nand U157 (N_157,In_812,In_897);
nand U158 (N_158,In_1777,In_1077);
or U159 (N_159,In_1779,In_376);
nand U160 (N_160,In_69,In_192);
and U161 (N_161,In_159,In_515);
or U162 (N_162,In_771,In_1182);
and U163 (N_163,In_952,In_507);
nand U164 (N_164,In_368,In_437);
xnor U165 (N_165,In_731,In_632);
or U166 (N_166,In_372,In_347);
nand U167 (N_167,In_865,In_1227);
nor U168 (N_168,In_182,In_801);
xor U169 (N_169,In_365,In_261);
or U170 (N_170,In_1573,In_979);
and U171 (N_171,In_878,In_1653);
or U172 (N_172,In_1045,In_205);
or U173 (N_173,In_77,In_1395);
nand U174 (N_174,In_896,In_1588);
or U175 (N_175,In_1042,In_206);
nor U176 (N_176,In_1018,In_913);
nor U177 (N_177,In_209,In_999);
xor U178 (N_178,In_1368,In_1465);
xor U179 (N_179,In_224,In_787);
or U180 (N_180,In_710,In_1838);
or U181 (N_181,In_1952,In_1569);
nor U182 (N_182,In_462,In_1427);
xor U183 (N_183,In_1181,In_1178);
xor U184 (N_184,In_1087,In_927);
nor U185 (N_185,In_1386,In_693);
xnor U186 (N_186,In_613,In_1832);
nand U187 (N_187,In_1200,In_324);
nor U188 (N_188,In_1903,In_1428);
and U189 (N_189,In_1581,In_306);
nand U190 (N_190,In_791,In_1797);
xor U191 (N_191,In_830,In_1608);
nand U192 (N_192,In_1725,In_1021);
nand U193 (N_193,In_899,In_419);
nor U194 (N_194,In_1373,In_1715);
and U195 (N_195,In_1223,In_598);
and U196 (N_196,In_1167,In_308);
nor U197 (N_197,In_201,In_550);
and U198 (N_198,In_269,In_722);
nor U199 (N_199,In_1867,In_1923);
and U200 (N_200,In_1876,In_1519);
or U201 (N_201,In_1936,In_1943);
nand U202 (N_202,In_687,In_1900);
nand U203 (N_203,In_1415,In_1097);
nand U204 (N_204,In_1571,In_557);
and U205 (N_205,In_1591,In_981);
nand U206 (N_206,In_603,In_945);
xor U207 (N_207,In_536,In_1336);
or U208 (N_208,In_1741,In_625);
and U209 (N_209,In_490,In_1347);
nor U210 (N_210,In_860,In_1868);
xor U211 (N_211,In_1422,In_1413);
nor U212 (N_212,In_955,In_534);
nand U213 (N_213,In_1432,In_418);
nor U214 (N_214,In_1627,In_1033);
or U215 (N_215,In_1787,In_400);
xor U216 (N_216,In_1663,In_941);
or U217 (N_217,In_1228,In_1617);
xnor U218 (N_218,In_1559,In_1100);
nor U219 (N_219,In_1891,In_271);
and U220 (N_220,In_525,In_10);
nand U221 (N_221,In_715,In_1179);
and U222 (N_222,In_1492,In_905);
nor U223 (N_223,In_1118,In_1184);
xnor U224 (N_224,In_1527,In_439);
or U225 (N_225,In_749,In_1150);
and U226 (N_226,In_466,In_155);
nand U227 (N_227,In_1901,In_1348);
or U228 (N_228,In_266,In_944);
nor U229 (N_229,In_1701,In_1498);
xnor U230 (N_230,In_1276,In_983);
nor U231 (N_231,In_1889,In_846);
and U232 (N_232,In_193,In_1798);
and U233 (N_233,In_518,In_1562);
or U234 (N_234,In_811,In_311);
xor U235 (N_235,In_1460,In_1667);
nand U236 (N_236,In_870,In_641);
nor U237 (N_237,In_1391,In_456);
nor U238 (N_238,In_1870,In_480);
nor U239 (N_239,In_920,In_873);
nand U240 (N_240,In_1824,In_391);
and U241 (N_241,In_496,In_178);
nand U242 (N_242,In_1795,In_1894);
and U243 (N_243,In_45,In_1711);
xnor U244 (N_244,In_1121,In_1481);
nor U245 (N_245,In_1751,In_1513);
xor U246 (N_246,In_327,In_12);
xnor U247 (N_247,In_1420,In_1727);
and U248 (N_248,In_1149,In_1114);
and U249 (N_249,In_664,In_551);
or U250 (N_250,In_173,In_1636);
xor U251 (N_251,In_665,In_1546);
or U252 (N_252,In_1596,In_752);
nor U253 (N_253,In_931,In_702);
and U254 (N_254,In_19,In_380);
nand U255 (N_255,In_1173,In_1555);
nand U256 (N_256,In_161,In_893);
xnor U257 (N_257,In_650,In_409);
xnor U258 (N_258,In_390,In_1140);
nor U259 (N_259,In_1353,In_708);
nand U260 (N_260,In_1878,In_1472);
and U261 (N_261,In_925,In_94);
or U262 (N_262,In_1995,In_840);
nand U263 (N_263,In_1226,In_392);
xor U264 (N_264,In_1994,In_1086);
xnor U265 (N_265,In_1750,In_1532);
nor U266 (N_266,In_1444,In_959);
nor U267 (N_267,In_552,In_1726);
nor U268 (N_268,In_130,In_1917);
nor U269 (N_269,In_128,In_1435);
nand U270 (N_270,In_1721,In_1880);
nand U271 (N_271,In_1800,In_1530);
nand U272 (N_272,In_1377,In_1677);
xor U273 (N_273,In_1874,In_1927);
and U274 (N_274,In_273,In_1640);
xnor U275 (N_275,In_280,In_1773);
xor U276 (N_276,In_1454,In_736);
nand U277 (N_277,In_355,In_1553);
xor U278 (N_278,In_106,In_644);
nor U279 (N_279,In_3,In_1783);
nor U280 (N_280,In_718,In_895);
xor U281 (N_281,In_124,In_303);
and U282 (N_282,In_1786,In_16);
nor U283 (N_283,In_1875,In_341);
nor U284 (N_284,In_1297,In_1823);
or U285 (N_285,In_84,In_877);
nand U286 (N_286,In_1175,In_508);
or U287 (N_287,In_1372,In_1584);
xor U288 (N_288,In_282,In_671);
or U289 (N_289,In_1857,In_339);
xnor U290 (N_290,In_699,In_1524);
and U291 (N_291,In_1854,In_481);
nor U292 (N_292,In_1911,In_381);
or U293 (N_293,In_510,In_397);
or U294 (N_294,In_1080,In_1067);
or U295 (N_295,In_681,In_453);
nand U296 (N_296,In_645,In_1886);
and U297 (N_297,In_1287,In_818);
nand U298 (N_298,In_744,In_705);
or U299 (N_299,In_475,In_62);
xnor U300 (N_300,In_1548,In_755);
nand U301 (N_301,In_86,In_420);
and U302 (N_302,In_1172,In_610);
or U303 (N_303,In_1772,In_1426);
and U304 (N_304,In_232,In_1594);
and U305 (N_305,In_961,In_144);
and U306 (N_306,In_1141,In_822);
xor U307 (N_307,In_1710,In_964);
or U308 (N_308,In_1941,In_184);
or U309 (N_309,In_1869,In_152);
xnor U310 (N_310,In_1478,In_1736);
nand U311 (N_311,In_348,In_1985);
nor U312 (N_312,In_165,In_56);
and U313 (N_313,In_1542,In_382);
or U314 (N_314,In_1737,In_24);
xor U315 (N_315,In_781,In_195);
and U316 (N_316,In_1014,In_1775);
nand U317 (N_317,In_1714,In_1047);
or U318 (N_318,In_1811,In_890);
nor U319 (N_319,In_1437,In_1381);
nand U320 (N_320,In_1293,In_806);
xnor U321 (N_321,In_614,In_1245);
or U322 (N_322,In_1039,In_587);
nor U323 (N_323,In_207,In_1449);
and U324 (N_324,In_751,In_1933);
nor U325 (N_325,In_1445,In_371);
nor U326 (N_326,In_1946,In_1157);
nand U327 (N_327,In_1024,In_40);
nand U328 (N_328,In_287,In_1535);
or U329 (N_329,In_136,In_472);
xnor U330 (N_330,In_698,In_1213);
and U331 (N_331,In_922,In_417);
nor U332 (N_332,In_986,In_559);
and U333 (N_333,In_1417,In_1628);
nand U334 (N_334,In_737,In_85);
and U335 (N_335,In_1910,In_839);
xnor U336 (N_336,In_1704,In_1412);
nand U337 (N_337,In_221,In_1464);
and U338 (N_338,In_875,In_297);
xor U339 (N_339,In_1019,In_1723);
xor U340 (N_340,In_1258,In_64);
nand U341 (N_341,In_38,In_1063);
and U342 (N_342,In_858,In_1508);
and U343 (N_343,In_204,In_461);
nor U344 (N_344,In_856,In_1068);
or U345 (N_345,In_909,In_1645);
or U346 (N_346,In_321,In_667);
nand U347 (N_347,In_734,In_1485);
and U348 (N_348,In_824,In_1316);
nor U349 (N_349,In_216,In_1984);
and U350 (N_350,In_406,In_1810);
nand U351 (N_351,In_960,In_452);
nor U352 (N_352,In_1283,In_322);
and U353 (N_353,In_1954,In_545);
xor U354 (N_354,In_1154,In_924);
xor U355 (N_355,In_1414,In_504);
nand U356 (N_356,In_447,In_1632);
xnor U357 (N_357,In_590,In_1094);
or U358 (N_358,In_1541,In_42);
nand U359 (N_359,In_435,In_226);
and U360 (N_360,In_783,In_170);
nor U361 (N_361,In_278,In_1755);
nand U362 (N_362,In_1937,In_1248);
nand U363 (N_363,In_393,In_1904);
nor U364 (N_364,In_1766,In_1820);
xor U365 (N_365,In_529,In_479);
and U366 (N_366,In_1700,In_1318);
nand U367 (N_367,In_468,In_1990);
xnor U368 (N_368,In_18,In_1421);
and U369 (N_369,In_1855,In_797);
xnor U370 (N_370,In_1302,In_39);
nand U371 (N_371,In_107,In_1674);
nand U372 (N_372,In_754,In_851);
nand U373 (N_373,In_1225,In_1123);
nand U374 (N_374,In_1176,In_1185);
nand U375 (N_375,In_1607,In_310);
nand U376 (N_376,In_258,In_1948);
and U377 (N_377,In_773,In_169);
nand U378 (N_378,In_149,In_1748);
xor U379 (N_379,In_1572,In_778);
nor U380 (N_380,In_1400,In_1659);
and U381 (N_381,In_427,In_1740);
or U382 (N_382,In_1489,In_1974);
xor U383 (N_383,In_300,In_1784);
and U384 (N_384,In_886,In_820);
or U385 (N_385,In_386,In_500);
xor U386 (N_386,In_436,In_1693);
nand U387 (N_387,In_111,In_401);
xnor U388 (N_388,In_148,In_788);
nand U389 (N_389,In_1968,In_1339);
nor U390 (N_390,In_289,In_618);
and U391 (N_391,In_1064,In_543);
or U392 (N_392,In_477,In_1805);
nand U393 (N_393,In_757,In_1458);
or U394 (N_394,In_1059,In_395);
xor U395 (N_395,In_821,In_1329);
xnor U396 (N_396,In_384,In_790);
xor U397 (N_397,In_426,In_1672);
nand U398 (N_398,In_1186,In_1637);
nor U399 (N_399,In_700,In_596);
nor U400 (N_400,In_1333,In_1046);
xor U401 (N_401,In_1560,In_172);
nand U402 (N_402,In_1126,In_1533);
and U403 (N_403,In_412,In_714);
nand U404 (N_404,In_1349,In_1920);
or U405 (N_405,In_1267,In_1424);
or U406 (N_406,In_441,In_1735);
or U407 (N_407,In_1011,In_1406);
and U408 (N_408,In_1394,In_786);
nand U409 (N_409,In_359,In_212);
xnor U410 (N_410,In_1928,In_1918);
and U411 (N_411,In_759,In_1243);
and U412 (N_412,In_143,In_150);
and U413 (N_413,In_1327,In_413);
nand U414 (N_414,In_654,In_8);
xnor U415 (N_415,In_795,In_985);
and U416 (N_416,In_1668,In_582);
nor U417 (N_417,In_906,In_1448);
nor U418 (N_418,In_637,In_1752);
nor U419 (N_419,In_132,In_853);
or U420 (N_420,In_74,In_1908);
or U421 (N_421,In_1696,In_404);
and U422 (N_422,In_211,In_847);
or U423 (N_423,In_1005,In_1660);
xor U424 (N_424,In_1354,In_1027);
nor U425 (N_425,In_110,In_862);
xnor U426 (N_426,In_1265,In_48);
and U427 (N_427,In_1281,In_168);
xnor U428 (N_428,In_1501,In_850);
xnor U429 (N_429,In_263,In_544);
and U430 (N_430,In_1983,In_568);
xnor U431 (N_431,In_1552,In_549);
xnor U432 (N_432,In_1801,In_72);
nand U433 (N_433,In_537,In_1143);
nor U434 (N_434,In_1076,In_635);
nand U435 (N_435,In_1235,In_50);
nand U436 (N_436,In_1108,In_1044);
nand U437 (N_437,In_1096,In_735);
nor U438 (N_438,In_363,In_876);
and U439 (N_439,In_1366,In_1375);
and U440 (N_440,In_1847,In_323);
nand U441 (N_441,In_131,In_345);
nor U442 (N_442,In_1006,In_814);
or U443 (N_443,In_974,In_1307);
nand U444 (N_444,In_1671,In_1313);
nor U445 (N_445,In_399,In_1338);
or U446 (N_446,In_1959,In_1898);
nand U447 (N_447,In_980,In_1497);
or U448 (N_448,In_1945,In_826);
nor U449 (N_449,In_1536,In_1545);
xor U450 (N_450,In_1563,In_743);
or U451 (N_451,In_1220,In_1961);
or U452 (N_452,In_1122,In_457);
nor U453 (N_453,In_1575,In_885);
and U454 (N_454,In_662,In_646);
and U455 (N_455,In_1641,In_17);
or U456 (N_456,In_1237,In_433);
or U457 (N_457,In_1212,In_1330);
and U458 (N_458,In_1621,In_1966);
or U459 (N_459,In_70,In_1753);
nand U460 (N_460,In_1057,In_668);
nand U461 (N_461,In_988,In_120);
or U462 (N_462,In_695,In_1317);
nor U463 (N_463,In_1526,In_1259);
nand U464 (N_464,In_133,In_1382);
or U465 (N_465,In_1881,In_1897);
or U466 (N_466,In_777,In_43);
and U467 (N_467,In_1684,In_1708);
and U468 (N_468,In_1164,In_1825);
xor U469 (N_469,In_1278,In_520);
nor U470 (N_470,In_91,In_1134);
xor U471 (N_471,In_304,In_1319);
or U472 (N_472,In_1129,In_166);
xnor U473 (N_473,In_1962,In_601);
nand U474 (N_474,In_1250,In_1371);
nor U475 (N_475,In_1072,In_802);
xor U476 (N_476,In_1073,In_1503);
and U477 (N_477,In_594,In_118);
nand U478 (N_478,In_1598,In_293);
or U479 (N_479,In_57,In_689);
nand U480 (N_480,In_581,In_1763);
and U481 (N_481,In_1152,In_1358);
nor U482 (N_482,In_794,In_1720);
and U483 (N_483,In_880,In_857);
nor U484 (N_484,In_1688,In_1095);
nand U485 (N_485,In_1812,In_242);
nor U486 (N_486,In_1219,In_252);
nor U487 (N_487,In_1230,In_1712);
or U488 (N_488,In_827,In_720);
nor U489 (N_489,In_93,In_1010);
nand U490 (N_490,In_1168,In_7);
nand U491 (N_491,In_1169,In_1116);
nor U492 (N_492,In_1370,In_421);
xnor U493 (N_493,In_1408,In_498);
or U494 (N_494,In_1656,In_712);
and U495 (N_495,In_1872,In_1829);
or U496 (N_496,In_163,In_1231);
xnor U497 (N_497,In_1144,In_721);
nand U498 (N_498,In_82,In_214);
nor U499 (N_499,In_248,In_181);
or U500 (N_500,In_378,In_1620);
nand U501 (N_501,In_102,In_387);
nand U502 (N_502,In_1051,In_1731);
nor U503 (N_503,In_22,In_227);
and U504 (N_504,In_809,In_816);
or U505 (N_505,In_501,In_1537);
nor U506 (N_506,In_1564,In_1171);
xor U507 (N_507,In_1038,In_604);
nor U508 (N_508,In_100,In_1879);
xor U509 (N_509,In_672,In_1017);
nand U510 (N_510,In_918,In_1052);
nor U511 (N_511,In_49,In_465);
nand U512 (N_512,In_1282,In_1981);
xnor U513 (N_513,In_626,In_746);
nand U514 (N_514,In_589,In_1029);
nor U515 (N_515,In_1442,In_1888);
xnor U516 (N_516,In_495,In_666);
nand U517 (N_517,In_1967,In_1619);
xor U518 (N_518,In_405,In_528);
or U519 (N_519,In_1603,In_329);
nor U520 (N_520,In_1858,In_1939);
xor U521 (N_521,In_316,In_233);
xnor U522 (N_522,In_1771,In_1273);
nand U523 (N_523,In_1022,In_487);
or U524 (N_524,In_1808,In_1298);
or U525 (N_525,In_116,In_281);
or U526 (N_526,In_1837,In_147);
nand U527 (N_527,In_1241,In_183);
xnor U528 (N_528,In_292,In_934);
and U529 (N_529,In_1924,In_1461);
or U530 (N_530,In_1264,In_1369);
or U531 (N_531,In_1376,In_711);
xor U532 (N_532,In_286,In_997);
xor U533 (N_533,In_1379,In_1860);
or U534 (N_534,In_1125,In_894);
and U535 (N_535,In_240,In_879);
xnor U536 (N_536,In_1434,In_1411);
or U537 (N_537,In_291,In_1942);
and U538 (N_538,In_527,In_274);
and U539 (N_539,In_1885,In_834);
xnor U540 (N_540,In_187,In_1346);
xor U541 (N_541,In_765,In_236);
nand U542 (N_542,In_1500,In_1951);
or U543 (N_543,In_936,In_140);
nand U544 (N_544,In_108,In_852);
or U545 (N_545,In_264,In_874);
nand U546 (N_546,In_334,In_935);
nand U547 (N_547,In_674,In_888);
and U548 (N_548,In_1873,In_591);
nand U549 (N_549,In_352,In_123);
and U550 (N_550,In_0,In_1998);
and U551 (N_551,In_180,In_1510);
and U552 (N_552,In_239,In_683);
and U553 (N_553,In_1048,In_1356);
and U554 (N_554,In_745,In_442);
xnor U555 (N_555,In_105,In_1505);
or U556 (N_556,In_1383,In_1635);
xnor U557 (N_557,In_539,In_1697);
nor U558 (N_558,In_588,In_99);
nor U559 (N_559,In_949,In_975);
nand U560 (N_560,In_374,In_1614);
nor U561 (N_561,In_276,In_1831);
and U562 (N_562,In_1597,In_32);
xor U563 (N_563,In_328,In_1301);
nor U564 (N_564,In_1681,In_648);
nand U565 (N_565,In_254,In_492);
or U566 (N_566,In_37,In_1296);
nor U567 (N_567,In_1031,In_701);
nand U568 (N_568,In_1082,In_307);
or U569 (N_569,In_1261,In_228);
nor U570 (N_570,In_1089,In_1192);
xor U571 (N_571,In_1993,In_1331);
and U572 (N_572,In_243,In_926);
nand U573 (N_573,In_1686,In_449);
and U574 (N_574,In_175,In_1522);
and U575 (N_575,In_1162,In_685);
nand U576 (N_576,In_1470,In_225);
xnor U577 (N_577,In_798,In_620);
xnor U578 (N_578,In_154,In_1439);
nor U579 (N_579,In_1618,In_1565);
or U580 (N_580,In_993,In_522);
and U581 (N_581,In_831,In_179);
nand U582 (N_582,In_298,In_1724);
or U583 (N_583,In_317,In_933);
xor U584 (N_584,In_898,In_1028);
xnor U585 (N_585,In_1842,In_30);
or U586 (N_586,In_396,In_272);
xor U587 (N_587,In_750,In_1050);
or U588 (N_588,In_1739,In_517);
nor U589 (N_589,In_1308,In_627);
nor U590 (N_590,In_194,In_1013);
nor U591 (N_591,In_904,In_488);
or U592 (N_592,In_398,In_884);
nand U593 (N_593,In_1055,In_1651);
and U594 (N_594,In_1856,In_584);
or U595 (N_595,In_1483,In_234);
nand U596 (N_596,In_6,In_11);
nor U597 (N_597,In_514,In_977);
and U598 (N_598,In_923,In_202);
or U599 (N_599,In_467,In_810);
and U600 (N_600,In_1647,In_521);
nand U601 (N_601,In_185,In_458);
and U602 (N_602,In_919,In_503);
xnor U603 (N_603,In_1665,In_767);
or U604 (N_604,In_1925,In_389);
nor U605 (N_605,In_1106,In_1328);
nand U606 (N_606,In_1978,In_364);
nand U607 (N_607,In_1127,In_1996);
or U608 (N_608,In_65,In_255);
or U609 (N_609,In_1266,In_259);
nor U610 (N_610,In_1790,In_1913);
and U611 (N_611,In_1661,In_903);
and U612 (N_612,In_237,In_353);
or U613 (N_613,In_1133,In_422);
xnor U614 (N_614,In_23,In_1204);
nand U615 (N_615,In_1570,In_158);
or U616 (N_616,In_615,In_770);
nor U617 (N_617,In_1166,In_570);
nand U618 (N_618,In_1722,In_1484);
nor U619 (N_619,In_1852,In_1341);
or U620 (N_620,In_1294,In_1834);
or U621 (N_621,In_842,In_1528);
or U622 (N_622,In_1299,In_555);
or U623 (N_623,In_1407,In_103);
or U624 (N_624,In_1746,In_1670);
nor U625 (N_625,In_369,In_1260);
and U626 (N_626,In_383,In_967);
nand U627 (N_627,In_1760,In_1944);
nor U628 (N_628,In_1357,In_1517);
nand U629 (N_629,In_633,In_1253);
or U630 (N_630,In_2,In_696);
or U631 (N_631,In_25,In_1576);
nand U632 (N_632,In_1305,In_1456);
or U633 (N_633,In_1989,In_725);
or U634 (N_634,In_497,In_709);
and U635 (N_635,In_728,In_844);
or U636 (N_636,In_1590,In_780);
nand U637 (N_637,In_769,In_58);
and U638 (N_638,In_1747,In_916);
xor U639 (N_639,In_1304,In_1616);
or U640 (N_640,In_1592,In_690);
nand U641 (N_641,In_1685,In_1486);
nor U642 (N_642,In_73,In_1915);
xnor U643 (N_643,In_1438,In_379);
nand U644 (N_644,In_63,In_1843);
or U645 (N_645,In_971,In_1269);
xor U646 (N_646,In_59,In_617);
xnor U647 (N_647,In_1208,In_561);
or U648 (N_648,In_1107,In_260);
or U649 (N_649,In_1813,In_1104);
nor U650 (N_650,In_1088,In_1890);
and U651 (N_651,In_1781,In_686);
and U652 (N_652,In_113,In_78);
and U653 (N_653,In_688,In_1871);
nand U654 (N_654,In_1907,In_1272);
nand U655 (N_655,In_1703,In_1249);
or U656 (N_656,In_1605,In_1971);
xnor U657 (N_657,In_229,In_1075);
nor U658 (N_658,In_1664,In_1070);
nand U659 (N_659,In_1499,In_1922);
xnor U660 (N_660,In_657,In_1506);
nor U661 (N_661,In_346,In_609);
or U662 (N_662,In_1101,In_1919);
xor U663 (N_663,In_1574,In_139);
or U664 (N_664,In_1599,In_1251);
xnor U665 (N_665,In_1324,In_800);
nor U666 (N_666,In_342,In_1844);
xor U667 (N_667,In_1794,In_1730);
or U668 (N_668,In_249,In_1135);
xnor U669 (N_669,In_987,In_1455);
nor U670 (N_670,In_595,In_600);
and U671 (N_671,In_104,In_756);
nand U672 (N_672,In_343,In_1344);
nor U673 (N_673,In_864,In_1793);
and U674 (N_674,In_607,In_577);
nand U675 (N_675,In_403,In_1462);
nor U676 (N_676,In_1409,In_112);
and U677 (N_677,In_189,In_1345);
or U678 (N_678,In_1419,In_630);
nand U679 (N_679,In_1090,In_1905);
xor U680 (N_680,In_1222,In_565);
and U681 (N_681,In_574,In_1694);
xnor U682 (N_682,In_28,In_177);
and U683 (N_683,In_1084,In_471);
xnor U684 (N_684,In_1764,In_1466);
xor U685 (N_685,In_616,In_1495);
xnor U686 (N_686,In_428,In_314);
and U687 (N_687,In_560,In_1549);
nand U688 (N_688,In_716,In_663);
nand U689 (N_689,In_1457,In_1830);
and U690 (N_690,In_302,In_469);
nor U691 (N_691,In_265,In_592);
or U692 (N_692,In_1652,In_1139);
and U693 (N_693,In_585,In_513);
xnor U694 (N_694,In_1158,In_1899);
xor U695 (N_695,In_1639,In_1676);
nor U696 (N_696,In_331,In_1374);
nand U697 (N_697,In_1648,In_1866);
or U698 (N_698,In_121,In_1705);
or U699 (N_699,In_1053,In_1023);
nand U700 (N_700,In_1579,In_1819);
nor U701 (N_701,In_932,In_1557);
nand U702 (N_702,In_606,In_167);
xnor U703 (N_703,In_1365,In_1161);
and U704 (N_704,In_1380,In_533);
or U705 (N_705,In_1964,In_268);
nand U706 (N_706,In_1000,In_247);
or U707 (N_707,In_80,In_267);
nand U708 (N_708,In_1004,In_1582);
xor U709 (N_709,In_1194,In_1359);
xor U710 (N_710,In_174,In_354);
or U711 (N_711,In_1255,In_463);
or U712 (N_712,In_1759,In_669);
nand U713 (N_713,In_250,In_126);
nand U714 (N_714,In_1709,In_953);
xor U715 (N_715,In_1836,In_1649);
xnor U716 (N_716,In_1972,In_1263);
nand U717 (N_717,In_1190,In_1529);
xnor U718 (N_718,In_1032,In_1692);
and U719 (N_719,In_1303,In_972);
nand U720 (N_720,In_1286,In_1699);
nor U721 (N_721,In_454,In_1401);
and U722 (N_722,In_915,In_1926);
nand U723 (N_723,In_370,In_1446);
xnor U724 (N_724,In_717,In_270);
xnor U725 (N_725,In_1474,In_1209);
nor U726 (N_726,In_1362,In_1036);
nor U727 (N_727,In_1988,In_1221);
nor U728 (N_728,In_859,In_294);
and U729 (N_729,In_1102,In_434);
xor U730 (N_730,In_1992,In_1568);
and U731 (N_731,In_245,In_1002);
nor U732 (N_732,In_1865,In_1826);
or U733 (N_733,In_1295,In_1949);
and U734 (N_734,In_1211,In_13);
or U735 (N_735,In_1289,In_1554);
nand U736 (N_736,In_692,In_1509);
nand U737 (N_737,In_425,In_1058);
nor U738 (N_738,In_1256,In_1650);
or U739 (N_739,In_486,In_1128);
xnor U740 (N_740,In_1950,In_1441);
nand U741 (N_741,In_44,In_66);
xnor U742 (N_742,In_506,In_1138);
nand U743 (N_743,In_1657,In_639);
and U744 (N_744,In_772,In_1459);
and U745 (N_745,In_1561,In_4);
nor U746 (N_746,In_1151,In_1882);
nor U747 (N_747,In_1034,In_1300);
or U748 (N_748,In_1160,In_176);
and U749 (N_749,In_231,In_1638);
nor U750 (N_750,In_1280,In_1056);
nand U751 (N_751,In_1833,In_917);
and U752 (N_752,In_946,In_530);
nand U753 (N_753,In_299,In_318);
nand U754 (N_754,In_1098,In_135);
or U755 (N_755,In_351,In_117);
xnor U756 (N_756,In_1666,In_998);
nor U757 (N_757,In_1403,In_109);
nand U758 (N_758,In_516,In_1585);
nor U759 (N_759,In_727,In_1291);
xnor U760 (N_760,In_1246,In_1543);
nor U761 (N_761,In_1274,In_869);
or U762 (N_762,In_789,In_564);
and U763 (N_763,In_1658,In_1447);
xor U764 (N_764,In_1884,In_813);
and U765 (N_765,In_1183,In_1774);
and U766 (N_766,In_1054,In_1351);
and U767 (N_767,In_335,In_1285);
or U768 (N_768,In_670,In_845);
or U769 (N_769,In_1451,In_1969);
and U770 (N_770,In_579,In_141);
and U771 (N_771,In_651,In_1360);
nand U772 (N_772,In_704,In_1643);
nand U773 (N_773,In_950,In_1799);
and U774 (N_774,In_1342,In_729);
xnor U775 (N_775,In_197,In_448);
nor U776 (N_776,In_540,In_432);
xor U777 (N_777,In_1240,In_246);
nor U778 (N_778,In_1,In_892);
nand U779 (N_779,In_1136,In_629);
or U780 (N_780,In_1782,In_1218);
nand U781 (N_781,In_1234,In_748);
xor U782 (N_782,In_455,In_1960);
or U783 (N_783,In_1431,In_1037);
nor U784 (N_784,In_438,In_1728);
and U785 (N_785,In_1387,In_608);
xnor U786 (N_786,In_90,In_46);
nor U787 (N_787,In_1803,In_742);
nand U788 (N_788,In_1613,In_1270);
and U789 (N_789,In_1120,In_1117);
and U790 (N_790,In_1550,In_766);
and U791 (N_791,In_223,In_1322);
nand U792 (N_792,In_978,In_68);
nand U793 (N_793,In_157,In_97);
xnor U794 (N_794,In_836,In_1290);
or U795 (N_795,In_597,In_1079);
nand U796 (N_796,In_833,In_1864);
nor U797 (N_797,In_337,In_558);
xor U798 (N_798,In_1689,In_697);
or U799 (N_799,In_360,In_943);
or U800 (N_800,In_1352,In_1770);
nand U801 (N_801,In_643,In_1818);
or U802 (N_802,In_1188,In_726);
xnor U803 (N_803,In_1163,In_1217);
nor U804 (N_804,In_1207,In_88);
nor U805 (N_805,In_83,In_416);
xnor U806 (N_806,In_782,In_1520);
or U807 (N_807,In_92,In_1769);
or U808 (N_808,In_1850,In_1436);
xor U809 (N_809,In_1745,In_1934);
xor U810 (N_810,In_1975,In_1956);
nand U811 (N_811,In_733,In_423);
xor U812 (N_812,In_1092,In_1624);
xnor U813 (N_813,In_119,In_1350);
nor U814 (N_814,In_1364,In_649);
nor U815 (N_815,In_1061,In_835);
and U816 (N_816,In_900,In_1973);
nor U817 (N_817,In_76,In_642);
nand U818 (N_818,In_1785,In_241);
xnor U819 (N_819,In_1815,In_1757);
nor U820 (N_820,In_1853,In_602);
or U821 (N_821,In_1463,In_283);
and U822 (N_822,In_373,In_965);
nand U823 (N_823,In_142,In_1883);
and U824 (N_824,In_1691,In_1991);
nor U825 (N_825,In_1544,In_775);
nand U826 (N_826,In_1778,In_656);
nor U827 (N_827,In_1398,In_71);
xor U828 (N_828,In_881,In_740);
nand U829 (N_829,In_402,In_473);
and U830 (N_830,In_215,In_807);
xor U831 (N_831,In_5,In_1622);
nand U832 (N_832,In_244,In_680);
xor U833 (N_833,In_719,In_375);
nand U834 (N_834,In_1202,In_774);
xor U835 (N_835,In_1851,In_1109);
nor U836 (N_836,In_1399,In_1914);
xor U837 (N_837,In_768,In_804);
and U838 (N_838,In_553,In_1216);
nor U839 (N_839,In_838,In_1210);
and U840 (N_840,In_493,In_1862);
and U841 (N_841,In_1132,In_15);
or U842 (N_842,In_823,In_451);
and U843 (N_843,In_837,In_1958);
nand U844 (N_844,In_1610,In_333);
nor U845 (N_845,In_1615,In_122);
nor U846 (N_846,In_509,In_361);
nor U847 (N_847,In_939,In_526);
nand U848 (N_848,In_1423,In_803);
xnor U849 (N_849,In_1767,In_512);
or U850 (N_850,In_1309,In_1452);
nor U851 (N_851,In_1583,In_1987);
and U852 (N_852,In_1756,In_450);
and U853 (N_853,In_1863,In_1069);
nor U854 (N_854,In_1103,In_411);
and U855 (N_855,In_1646,In_1999);
or U856 (N_856,In_476,In_762);
and U857 (N_857,In_1137,In_1673);
nand U858 (N_858,In_1334,In_296);
xor U859 (N_859,In_872,In_1593);
nand U860 (N_860,In_485,In_954);
nand U861 (N_861,In_1468,In_956);
and U862 (N_862,In_1405,In_907);
or U863 (N_863,In_1093,In_1634);
nand U864 (N_864,In_134,In_1026);
or U865 (N_865,In_1887,In_1578);
and U866 (N_866,In_1035,In_929);
nor U867 (N_867,In_460,In_580);
nor U868 (N_868,In_682,In_575);
nand U869 (N_869,In_571,In_1547);
nor U870 (N_870,In_1443,In_1174);
nor U871 (N_871,In_1706,In_491);
xnor U872 (N_872,In_889,In_1198);
xnor U873 (N_873,In_1849,In_478);
nor U874 (N_874,In_901,In_1749);
nand U875 (N_875,In_1105,In_1841);
xnor U876 (N_876,In_1835,In_1214);
nor U877 (N_877,In_1609,In_849);
or U878 (N_878,In_1390,In_984);
xor U879 (N_879,In_20,In_1429);
nand U880 (N_880,In_305,In_79);
nor U881 (N_881,In_1320,In_429);
xor U882 (N_882,In_230,In_661);
and U883 (N_883,In_96,In_623);
xor U884 (N_884,In_659,In_992);
and U885 (N_885,In_200,In_1980);
xnor U886 (N_886,In_825,In_808);
nor U887 (N_887,In_1940,In_1893);
and U888 (N_888,In_871,In_1476);
and U889 (N_889,In_1315,In_1325);
nand U890 (N_890,In_576,In_1930);
nor U891 (N_891,In_1611,In_1538);
and U892 (N_892,In_1232,In_1780);
nand U893 (N_893,In_1822,In_1326);
or U894 (N_894,In_1083,In_443);
nor U895 (N_895,In_1916,In_1765);
nor U896 (N_896,In_67,In_1738);
and U897 (N_897,In_1388,In_1754);
or U898 (N_898,In_854,In_89);
xor U899 (N_899,In_1695,In_127);
and U900 (N_900,In_631,In_125);
nor U901 (N_901,In_196,In_1254);
nor U902 (N_902,In_1416,In_356);
nand U903 (N_903,In_1490,In_855);
xor U904 (N_904,In_362,In_991);
or U905 (N_905,In_1440,In_619);
xnor U906 (N_906,In_1201,In_408);
nor U907 (N_907,In_484,In_1471);
and U908 (N_908,In_198,In_1397);
xnor U909 (N_909,In_586,In_785);
or U910 (N_910,In_1145,In_1323);
nand U911 (N_911,In_253,In_1236);
nor U912 (N_912,In_1009,In_547);
xor U913 (N_913,In_1970,In_970);
or U914 (N_914,In_1410,In_1195);
and U915 (N_915,In_914,In_1311);
and U916 (N_916,In_54,In_1909);
nor U917 (N_917,In_1902,In_410);
nand U918 (N_918,In_1895,In_966);
nor U919 (N_919,In_1193,In_1845);
xor U920 (N_920,In_1566,In_908);
nor U921 (N_921,In_1189,In_1821);
nand U922 (N_922,In_1690,In_1367);
nand U923 (N_923,In_982,In_1877);
xnor U924 (N_924,In_1802,In_1982);
or U925 (N_925,In_1512,In_679);
xor U926 (N_926,In_673,In_1165);
nand U927 (N_927,In_724,In_1040);
nand U928 (N_928,In_284,In_848);
or U929 (N_929,In_1085,In_61);
xor U930 (N_930,In_1131,In_1099);
or U931 (N_931,In_1288,In_1335);
nand U932 (N_932,In_1742,In_1531);
nor U933 (N_933,In_1814,In_1947);
and U934 (N_934,In_1586,In_145);
nand U935 (N_935,In_989,In_1343);
nand U936 (N_936,In_257,In_760);
or U937 (N_937,In_295,In_684);
and U938 (N_938,In_741,In_1156);
and U939 (N_939,In_320,In_407);
xnor U940 (N_940,In_957,In_815);
and U941 (N_941,In_1718,In_164);
nor U942 (N_942,In_1450,In_1846);
or U943 (N_943,In_612,In_1630);
or U944 (N_944,In_841,In_1840);
and U945 (N_945,In_947,In_190);
nand U946 (N_946,In_691,In_1030);
nor U947 (N_947,In_677,In_1404);
and U948 (N_948,In_940,In_1159);
nor U949 (N_949,In_332,In_482);
and U950 (N_950,In_1262,In_1340);
and U951 (N_951,In_887,In_219);
nand U952 (N_952,In_1828,In_1979);
and U953 (N_953,In_1734,In_1453);
and U954 (N_954,In_222,In_542);
or U955 (N_955,In_1467,In_1025);
or U956 (N_956,In_35,In_562);
nor U957 (N_957,In_703,In_340);
nand U958 (N_958,In_430,In_963);
and U959 (N_959,In_1859,In_707);
or U960 (N_960,In_470,In_1719);
xnor U961 (N_961,In_217,In_653);
xor U962 (N_962,In_1662,In_41);
or U963 (N_963,In_1229,In_624);
nand U964 (N_964,In_1935,In_1687);
or U965 (N_965,In_1839,In_1306);
or U966 (N_966,In_902,In_1425);
nand U967 (N_967,In_1496,In_1654);
and U968 (N_968,In_1600,In_1215);
nor U969 (N_969,In_1477,In_1602);
and U970 (N_970,In_548,In_1148);
nand U971 (N_971,In_1604,In_357);
or U972 (N_972,In_1384,In_1633);
and U973 (N_973,In_1041,In_1491);
nand U974 (N_974,In_1049,In_1396);
and U975 (N_975,In_706,In_538);
or U976 (N_976,In_115,In_1115);
and U977 (N_977,In_761,In_1587);
and U978 (N_978,In_1271,In_27);
nand U979 (N_979,In_1393,In_1196);
and U980 (N_980,In_1776,In_1804);
and U981 (N_981,In_53,In_1518);
nor U982 (N_982,In_414,In_275);
xnor U983 (N_983,In_1469,In_203);
or U984 (N_984,In_1066,In_1487);
or U985 (N_985,In_1929,In_829);
or U986 (N_986,In_26,In_1732);
nor U987 (N_987,In_256,In_388);
nand U988 (N_988,In_1589,In_1986);
nand U989 (N_989,In_1521,In_1606);
or U990 (N_990,In_817,In_1733);
and U991 (N_991,In_338,In_1268);
or U992 (N_992,In_1682,In_171);
nor U993 (N_993,In_1480,In_640);
or U994 (N_994,In_220,In_238);
nand U995 (N_995,In_1642,In_563);
nor U996 (N_996,In_385,In_319);
xor U997 (N_997,In_1003,In_1792);
nor U998 (N_998,In_1147,In_446);
nor U999 (N_999,In_33,In_1702);
nor U1000 (N_1000,In_215,In_160);
nor U1001 (N_1001,In_685,In_84);
nor U1002 (N_1002,In_1471,In_842);
xor U1003 (N_1003,In_1318,In_412);
nor U1004 (N_1004,In_131,In_457);
nand U1005 (N_1005,In_1378,In_1395);
or U1006 (N_1006,In_1535,In_1631);
xor U1007 (N_1007,In_1633,In_1929);
nand U1008 (N_1008,In_954,In_583);
or U1009 (N_1009,In_1953,In_1839);
and U1010 (N_1010,In_1145,In_1692);
xor U1011 (N_1011,In_837,In_1651);
nand U1012 (N_1012,In_1012,In_1989);
and U1013 (N_1013,In_1400,In_407);
or U1014 (N_1014,In_788,In_769);
and U1015 (N_1015,In_58,In_987);
nor U1016 (N_1016,In_1999,In_147);
nor U1017 (N_1017,In_1779,In_924);
xor U1018 (N_1018,In_619,In_1161);
nand U1019 (N_1019,In_155,In_732);
and U1020 (N_1020,In_1906,In_126);
nand U1021 (N_1021,In_1508,In_1993);
nor U1022 (N_1022,In_1100,In_1970);
or U1023 (N_1023,In_1642,In_1868);
xnor U1024 (N_1024,In_22,In_100);
nor U1025 (N_1025,In_1646,In_757);
nor U1026 (N_1026,In_398,In_486);
nor U1027 (N_1027,In_53,In_1781);
or U1028 (N_1028,In_1319,In_709);
and U1029 (N_1029,In_1260,In_686);
and U1030 (N_1030,In_48,In_323);
nor U1031 (N_1031,In_1009,In_1973);
nor U1032 (N_1032,In_1902,In_1945);
and U1033 (N_1033,In_1740,In_537);
and U1034 (N_1034,In_235,In_1921);
xnor U1035 (N_1035,In_832,In_1230);
nand U1036 (N_1036,In_1699,In_1740);
xnor U1037 (N_1037,In_551,In_787);
and U1038 (N_1038,In_811,In_1896);
and U1039 (N_1039,In_917,In_1348);
or U1040 (N_1040,In_1091,In_963);
nand U1041 (N_1041,In_1477,In_1677);
xor U1042 (N_1042,In_1758,In_1133);
nand U1043 (N_1043,In_1754,In_1180);
xnor U1044 (N_1044,In_873,In_1377);
nand U1045 (N_1045,In_18,In_847);
or U1046 (N_1046,In_631,In_468);
or U1047 (N_1047,In_35,In_24);
nand U1048 (N_1048,In_684,In_453);
and U1049 (N_1049,In_1211,In_1483);
nand U1050 (N_1050,In_385,In_1310);
and U1051 (N_1051,In_1481,In_191);
and U1052 (N_1052,In_1353,In_459);
nor U1053 (N_1053,In_32,In_292);
nor U1054 (N_1054,In_1457,In_156);
or U1055 (N_1055,In_76,In_1535);
or U1056 (N_1056,In_836,In_1034);
nor U1057 (N_1057,In_903,In_1776);
nand U1058 (N_1058,In_282,In_1024);
or U1059 (N_1059,In_1118,In_1855);
nand U1060 (N_1060,In_843,In_1020);
xor U1061 (N_1061,In_884,In_1326);
nor U1062 (N_1062,In_1131,In_1454);
nand U1063 (N_1063,In_124,In_948);
or U1064 (N_1064,In_437,In_1766);
xnor U1065 (N_1065,In_1383,In_31);
nand U1066 (N_1066,In_1016,In_1465);
xnor U1067 (N_1067,In_760,In_1187);
nand U1068 (N_1068,In_1518,In_1626);
nand U1069 (N_1069,In_1827,In_730);
nand U1070 (N_1070,In_1503,In_87);
or U1071 (N_1071,In_14,In_906);
nor U1072 (N_1072,In_263,In_1811);
nand U1073 (N_1073,In_1005,In_1976);
nand U1074 (N_1074,In_1499,In_1421);
and U1075 (N_1075,In_641,In_553);
nor U1076 (N_1076,In_1394,In_1634);
or U1077 (N_1077,In_768,In_1753);
nand U1078 (N_1078,In_1828,In_1035);
or U1079 (N_1079,In_1847,In_758);
nand U1080 (N_1080,In_230,In_1119);
xor U1081 (N_1081,In_85,In_817);
nor U1082 (N_1082,In_660,In_1969);
nor U1083 (N_1083,In_813,In_1635);
xnor U1084 (N_1084,In_1359,In_1410);
xnor U1085 (N_1085,In_1976,In_837);
and U1086 (N_1086,In_320,In_1983);
or U1087 (N_1087,In_200,In_1845);
nor U1088 (N_1088,In_1415,In_558);
nand U1089 (N_1089,In_1439,In_178);
or U1090 (N_1090,In_776,In_1304);
nand U1091 (N_1091,In_624,In_1127);
nand U1092 (N_1092,In_376,In_878);
nor U1093 (N_1093,In_1087,In_932);
xnor U1094 (N_1094,In_284,In_270);
nor U1095 (N_1095,In_1542,In_373);
nor U1096 (N_1096,In_896,In_626);
nand U1097 (N_1097,In_424,In_1739);
nor U1098 (N_1098,In_1838,In_1005);
and U1099 (N_1099,In_839,In_275);
nor U1100 (N_1100,In_844,In_1126);
nand U1101 (N_1101,In_756,In_649);
and U1102 (N_1102,In_178,In_316);
or U1103 (N_1103,In_1995,In_367);
nand U1104 (N_1104,In_703,In_827);
and U1105 (N_1105,In_1620,In_797);
nor U1106 (N_1106,In_1905,In_769);
xnor U1107 (N_1107,In_19,In_850);
or U1108 (N_1108,In_511,In_396);
xor U1109 (N_1109,In_833,In_1877);
xor U1110 (N_1110,In_1140,In_608);
and U1111 (N_1111,In_1709,In_1540);
and U1112 (N_1112,In_164,In_1959);
or U1113 (N_1113,In_1704,In_869);
nor U1114 (N_1114,In_25,In_763);
nand U1115 (N_1115,In_1059,In_1868);
nor U1116 (N_1116,In_1632,In_1536);
and U1117 (N_1117,In_8,In_131);
nor U1118 (N_1118,In_503,In_1495);
nand U1119 (N_1119,In_456,In_1854);
nor U1120 (N_1120,In_1323,In_61);
nand U1121 (N_1121,In_1299,In_508);
or U1122 (N_1122,In_1801,In_716);
xor U1123 (N_1123,In_1161,In_1580);
nor U1124 (N_1124,In_1111,In_1390);
nand U1125 (N_1125,In_895,In_1247);
and U1126 (N_1126,In_1552,In_266);
or U1127 (N_1127,In_741,In_378);
and U1128 (N_1128,In_817,In_241);
nand U1129 (N_1129,In_1208,In_522);
nand U1130 (N_1130,In_1779,In_1701);
nor U1131 (N_1131,In_913,In_585);
and U1132 (N_1132,In_1517,In_1461);
xnor U1133 (N_1133,In_946,In_326);
nand U1134 (N_1134,In_518,In_732);
nand U1135 (N_1135,In_1551,In_1735);
and U1136 (N_1136,In_1689,In_167);
xor U1137 (N_1137,In_1637,In_365);
and U1138 (N_1138,In_708,In_1738);
and U1139 (N_1139,In_993,In_1203);
and U1140 (N_1140,In_1632,In_981);
nand U1141 (N_1141,In_731,In_1247);
or U1142 (N_1142,In_32,In_751);
and U1143 (N_1143,In_331,In_1415);
and U1144 (N_1144,In_1813,In_718);
nor U1145 (N_1145,In_630,In_1260);
xnor U1146 (N_1146,In_1918,In_227);
and U1147 (N_1147,In_1499,In_866);
or U1148 (N_1148,In_447,In_401);
and U1149 (N_1149,In_1743,In_506);
nand U1150 (N_1150,In_142,In_698);
nor U1151 (N_1151,In_364,In_727);
and U1152 (N_1152,In_932,In_1352);
and U1153 (N_1153,In_523,In_1087);
nor U1154 (N_1154,In_144,In_205);
xnor U1155 (N_1155,In_677,In_1973);
nor U1156 (N_1156,In_1912,In_555);
or U1157 (N_1157,In_797,In_487);
nand U1158 (N_1158,In_231,In_500);
nand U1159 (N_1159,In_625,In_685);
and U1160 (N_1160,In_1775,In_1125);
nor U1161 (N_1161,In_1027,In_1480);
nor U1162 (N_1162,In_926,In_1523);
nand U1163 (N_1163,In_1046,In_1591);
nand U1164 (N_1164,In_1190,In_1136);
or U1165 (N_1165,In_1660,In_314);
xnor U1166 (N_1166,In_1346,In_1671);
xor U1167 (N_1167,In_655,In_836);
and U1168 (N_1168,In_1866,In_558);
or U1169 (N_1169,In_1247,In_1993);
xor U1170 (N_1170,In_1805,In_878);
nand U1171 (N_1171,In_1973,In_415);
xnor U1172 (N_1172,In_1460,In_148);
xnor U1173 (N_1173,In_1269,In_1017);
or U1174 (N_1174,In_460,In_940);
or U1175 (N_1175,In_47,In_462);
or U1176 (N_1176,In_1518,In_1219);
and U1177 (N_1177,In_1803,In_1363);
xnor U1178 (N_1178,In_425,In_77);
nor U1179 (N_1179,In_119,In_812);
xnor U1180 (N_1180,In_1182,In_1238);
xor U1181 (N_1181,In_1153,In_1028);
or U1182 (N_1182,In_1108,In_293);
nor U1183 (N_1183,In_622,In_1916);
nor U1184 (N_1184,In_1471,In_1118);
or U1185 (N_1185,In_369,In_1925);
nand U1186 (N_1186,In_1566,In_81);
nand U1187 (N_1187,In_405,In_388);
and U1188 (N_1188,In_315,In_788);
nor U1189 (N_1189,In_931,In_61);
or U1190 (N_1190,In_108,In_1966);
or U1191 (N_1191,In_1674,In_1676);
xor U1192 (N_1192,In_7,In_1076);
or U1193 (N_1193,In_665,In_312);
xor U1194 (N_1194,In_285,In_1397);
nand U1195 (N_1195,In_1862,In_549);
and U1196 (N_1196,In_1284,In_1763);
or U1197 (N_1197,In_874,In_1610);
or U1198 (N_1198,In_1433,In_1800);
nand U1199 (N_1199,In_1778,In_1650);
or U1200 (N_1200,In_1246,In_213);
nand U1201 (N_1201,In_1171,In_84);
and U1202 (N_1202,In_1244,In_414);
or U1203 (N_1203,In_1234,In_1962);
xor U1204 (N_1204,In_1505,In_833);
nand U1205 (N_1205,In_881,In_259);
xnor U1206 (N_1206,In_1522,In_1616);
or U1207 (N_1207,In_222,In_1763);
nand U1208 (N_1208,In_1511,In_1057);
and U1209 (N_1209,In_439,In_1569);
and U1210 (N_1210,In_398,In_1170);
and U1211 (N_1211,In_332,In_1733);
and U1212 (N_1212,In_258,In_910);
or U1213 (N_1213,In_1891,In_653);
nand U1214 (N_1214,In_1291,In_518);
and U1215 (N_1215,In_35,In_1507);
or U1216 (N_1216,In_1288,In_384);
and U1217 (N_1217,In_1863,In_637);
xor U1218 (N_1218,In_608,In_215);
xor U1219 (N_1219,In_145,In_912);
or U1220 (N_1220,In_392,In_1178);
nor U1221 (N_1221,In_505,In_6);
xnor U1222 (N_1222,In_602,In_1121);
nand U1223 (N_1223,In_1427,In_939);
or U1224 (N_1224,In_966,In_1693);
or U1225 (N_1225,In_26,In_254);
nor U1226 (N_1226,In_529,In_30);
nand U1227 (N_1227,In_566,In_675);
and U1228 (N_1228,In_974,In_421);
xor U1229 (N_1229,In_132,In_1336);
nor U1230 (N_1230,In_286,In_1585);
nand U1231 (N_1231,In_1115,In_1754);
and U1232 (N_1232,In_1229,In_1677);
and U1233 (N_1233,In_781,In_447);
nand U1234 (N_1234,In_1696,In_650);
nand U1235 (N_1235,In_791,In_1078);
nor U1236 (N_1236,In_881,In_460);
nand U1237 (N_1237,In_1953,In_128);
nor U1238 (N_1238,In_344,In_1330);
nand U1239 (N_1239,In_699,In_1789);
nor U1240 (N_1240,In_182,In_1491);
or U1241 (N_1241,In_1589,In_981);
xor U1242 (N_1242,In_276,In_1666);
and U1243 (N_1243,In_599,In_1167);
xnor U1244 (N_1244,In_418,In_423);
nand U1245 (N_1245,In_35,In_576);
and U1246 (N_1246,In_1859,In_121);
nand U1247 (N_1247,In_54,In_214);
or U1248 (N_1248,In_1022,In_1072);
or U1249 (N_1249,In_265,In_449);
nor U1250 (N_1250,In_1256,In_639);
and U1251 (N_1251,In_1680,In_1604);
xnor U1252 (N_1252,In_904,In_1336);
nor U1253 (N_1253,In_66,In_1604);
nor U1254 (N_1254,In_1068,In_980);
and U1255 (N_1255,In_1481,In_819);
or U1256 (N_1256,In_1918,In_621);
or U1257 (N_1257,In_252,In_555);
xor U1258 (N_1258,In_1,In_1990);
or U1259 (N_1259,In_1157,In_383);
and U1260 (N_1260,In_1280,In_1254);
and U1261 (N_1261,In_1173,In_1388);
or U1262 (N_1262,In_647,In_1533);
nand U1263 (N_1263,In_1524,In_69);
nor U1264 (N_1264,In_131,In_1656);
nand U1265 (N_1265,In_1650,In_1730);
nand U1266 (N_1266,In_1842,In_430);
xor U1267 (N_1267,In_1033,In_290);
and U1268 (N_1268,In_908,In_1525);
and U1269 (N_1269,In_1935,In_753);
and U1270 (N_1270,In_656,In_48);
xnor U1271 (N_1271,In_1386,In_377);
or U1272 (N_1272,In_518,In_432);
nor U1273 (N_1273,In_869,In_303);
nand U1274 (N_1274,In_449,In_1856);
nand U1275 (N_1275,In_721,In_936);
xor U1276 (N_1276,In_862,In_1707);
nor U1277 (N_1277,In_758,In_1848);
xor U1278 (N_1278,In_329,In_1079);
or U1279 (N_1279,In_1932,In_1907);
and U1280 (N_1280,In_670,In_1570);
or U1281 (N_1281,In_1322,In_918);
nand U1282 (N_1282,In_179,In_1309);
xor U1283 (N_1283,In_334,In_1055);
xnor U1284 (N_1284,In_122,In_94);
xor U1285 (N_1285,In_1598,In_450);
nor U1286 (N_1286,In_1173,In_1259);
xnor U1287 (N_1287,In_1433,In_1172);
and U1288 (N_1288,In_1560,In_1962);
nand U1289 (N_1289,In_1403,In_1320);
or U1290 (N_1290,In_630,In_378);
and U1291 (N_1291,In_279,In_560);
and U1292 (N_1292,In_1304,In_778);
nor U1293 (N_1293,In_1824,In_455);
or U1294 (N_1294,In_324,In_1913);
or U1295 (N_1295,In_683,In_1153);
and U1296 (N_1296,In_1624,In_1329);
nand U1297 (N_1297,In_726,In_245);
and U1298 (N_1298,In_1229,In_1468);
nand U1299 (N_1299,In_789,In_871);
nor U1300 (N_1300,In_1577,In_697);
nor U1301 (N_1301,In_9,In_1370);
xnor U1302 (N_1302,In_843,In_796);
or U1303 (N_1303,In_95,In_1465);
xnor U1304 (N_1304,In_1702,In_367);
nand U1305 (N_1305,In_248,In_1531);
and U1306 (N_1306,In_1336,In_38);
and U1307 (N_1307,In_1108,In_849);
and U1308 (N_1308,In_208,In_420);
or U1309 (N_1309,In_1942,In_662);
xnor U1310 (N_1310,In_1312,In_50);
or U1311 (N_1311,In_1046,In_1455);
xor U1312 (N_1312,In_84,In_1994);
nor U1313 (N_1313,In_660,In_615);
and U1314 (N_1314,In_1721,In_1240);
nand U1315 (N_1315,In_1659,In_1859);
nand U1316 (N_1316,In_1843,In_377);
or U1317 (N_1317,In_1078,In_591);
or U1318 (N_1318,In_1850,In_1994);
or U1319 (N_1319,In_1084,In_994);
or U1320 (N_1320,In_766,In_1669);
nor U1321 (N_1321,In_992,In_1581);
nand U1322 (N_1322,In_318,In_530);
and U1323 (N_1323,In_826,In_614);
nand U1324 (N_1324,In_1721,In_775);
nor U1325 (N_1325,In_949,In_466);
or U1326 (N_1326,In_1340,In_50);
xnor U1327 (N_1327,In_1345,In_769);
nand U1328 (N_1328,In_1364,In_1777);
xnor U1329 (N_1329,In_1580,In_572);
or U1330 (N_1330,In_1769,In_1608);
or U1331 (N_1331,In_691,In_900);
or U1332 (N_1332,In_1795,In_1645);
xnor U1333 (N_1333,In_1501,In_991);
and U1334 (N_1334,In_492,In_1797);
nor U1335 (N_1335,In_705,In_403);
or U1336 (N_1336,In_1879,In_284);
and U1337 (N_1337,In_578,In_285);
nor U1338 (N_1338,In_991,In_328);
nor U1339 (N_1339,In_980,In_1958);
nand U1340 (N_1340,In_126,In_1453);
and U1341 (N_1341,In_1898,In_1571);
or U1342 (N_1342,In_844,In_1490);
nor U1343 (N_1343,In_1082,In_760);
and U1344 (N_1344,In_507,In_1282);
xnor U1345 (N_1345,In_808,In_1460);
or U1346 (N_1346,In_463,In_50);
or U1347 (N_1347,In_706,In_1018);
or U1348 (N_1348,In_664,In_754);
xnor U1349 (N_1349,In_147,In_1113);
xnor U1350 (N_1350,In_98,In_1395);
nand U1351 (N_1351,In_1927,In_1380);
or U1352 (N_1352,In_19,In_1689);
xnor U1353 (N_1353,In_1550,In_292);
and U1354 (N_1354,In_1112,In_1019);
or U1355 (N_1355,In_806,In_1218);
xor U1356 (N_1356,In_351,In_1259);
nand U1357 (N_1357,In_808,In_1658);
nand U1358 (N_1358,In_79,In_1735);
or U1359 (N_1359,In_841,In_1323);
and U1360 (N_1360,In_1403,In_175);
xnor U1361 (N_1361,In_1971,In_38);
or U1362 (N_1362,In_1700,In_1405);
nor U1363 (N_1363,In_1185,In_1764);
and U1364 (N_1364,In_97,In_957);
nand U1365 (N_1365,In_889,In_1997);
xnor U1366 (N_1366,In_1437,In_515);
xor U1367 (N_1367,In_24,In_1619);
and U1368 (N_1368,In_1845,In_1275);
nand U1369 (N_1369,In_1763,In_1616);
nor U1370 (N_1370,In_331,In_1723);
nand U1371 (N_1371,In_1069,In_638);
xnor U1372 (N_1372,In_1174,In_645);
nor U1373 (N_1373,In_174,In_1834);
and U1374 (N_1374,In_649,In_759);
xor U1375 (N_1375,In_650,In_474);
nand U1376 (N_1376,In_367,In_1854);
and U1377 (N_1377,In_1862,In_1853);
nand U1378 (N_1378,In_1098,In_1467);
xnor U1379 (N_1379,In_1885,In_1377);
and U1380 (N_1380,In_124,In_1079);
and U1381 (N_1381,In_363,In_249);
or U1382 (N_1382,In_1609,In_1473);
nor U1383 (N_1383,In_1300,In_773);
and U1384 (N_1384,In_916,In_1562);
or U1385 (N_1385,In_349,In_1967);
and U1386 (N_1386,In_1477,In_689);
xor U1387 (N_1387,In_733,In_1564);
and U1388 (N_1388,In_332,In_275);
and U1389 (N_1389,In_558,In_1539);
xor U1390 (N_1390,In_541,In_1869);
and U1391 (N_1391,In_1273,In_1948);
nor U1392 (N_1392,In_1996,In_1946);
nor U1393 (N_1393,In_1330,In_1587);
nor U1394 (N_1394,In_1283,In_634);
xor U1395 (N_1395,In_135,In_782);
nand U1396 (N_1396,In_1227,In_842);
or U1397 (N_1397,In_886,In_1043);
nand U1398 (N_1398,In_1915,In_1277);
nand U1399 (N_1399,In_725,In_826);
or U1400 (N_1400,In_169,In_534);
nand U1401 (N_1401,In_1378,In_871);
and U1402 (N_1402,In_793,In_1709);
nand U1403 (N_1403,In_998,In_1810);
or U1404 (N_1404,In_675,In_1);
nand U1405 (N_1405,In_1992,In_1662);
or U1406 (N_1406,In_1130,In_976);
and U1407 (N_1407,In_591,In_1785);
xnor U1408 (N_1408,In_1690,In_638);
or U1409 (N_1409,In_1639,In_1007);
xnor U1410 (N_1410,In_590,In_680);
nand U1411 (N_1411,In_862,In_846);
or U1412 (N_1412,In_108,In_1267);
nand U1413 (N_1413,In_88,In_388);
and U1414 (N_1414,In_1867,In_1870);
and U1415 (N_1415,In_1154,In_583);
nand U1416 (N_1416,In_318,In_665);
nand U1417 (N_1417,In_982,In_383);
nand U1418 (N_1418,In_741,In_167);
nor U1419 (N_1419,In_690,In_371);
xor U1420 (N_1420,In_1069,In_153);
xnor U1421 (N_1421,In_1078,In_643);
xor U1422 (N_1422,In_1323,In_1848);
nand U1423 (N_1423,In_1242,In_98);
nor U1424 (N_1424,In_376,In_266);
or U1425 (N_1425,In_309,In_1265);
nor U1426 (N_1426,In_59,In_1937);
nor U1427 (N_1427,In_1035,In_804);
or U1428 (N_1428,In_1859,In_1105);
xnor U1429 (N_1429,In_1196,In_1916);
nand U1430 (N_1430,In_257,In_1968);
nand U1431 (N_1431,In_355,In_1367);
nand U1432 (N_1432,In_1336,In_1802);
nand U1433 (N_1433,In_1873,In_773);
nand U1434 (N_1434,In_1615,In_272);
xor U1435 (N_1435,In_498,In_1541);
xor U1436 (N_1436,In_1314,In_743);
and U1437 (N_1437,In_1944,In_423);
or U1438 (N_1438,In_451,In_1596);
xnor U1439 (N_1439,In_2,In_1351);
nand U1440 (N_1440,In_134,In_488);
xnor U1441 (N_1441,In_224,In_1932);
nor U1442 (N_1442,In_1690,In_1903);
or U1443 (N_1443,In_1351,In_541);
or U1444 (N_1444,In_442,In_732);
nand U1445 (N_1445,In_111,In_1744);
or U1446 (N_1446,In_1405,In_546);
and U1447 (N_1447,In_16,In_1766);
nand U1448 (N_1448,In_1043,In_1851);
nand U1449 (N_1449,In_1877,In_1086);
nand U1450 (N_1450,In_831,In_564);
and U1451 (N_1451,In_506,In_1338);
or U1452 (N_1452,In_1730,In_1156);
nand U1453 (N_1453,In_1174,In_1187);
and U1454 (N_1454,In_834,In_1072);
xor U1455 (N_1455,In_1304,In_802);
and U1456 (N_1456,In_1720,In_47);
or U1457 (N_1457,In_1611,In_1206);
or U1458 (N_1458,In_1750,In_188);
xnor U1459 (N_1459,In_647,In_850);
nor U1460 (N_1460,In_800,In_60);
or U1461 (N_1461,In_960,In_1993);
nor U1462 (N_1462,In_437,In_424);
and U1463 (N_1463,In_426,In_919);
xor U1464 (N_1464,In_1300,In_272);
and U1465 (N_1465,In_1884,In_797);
and U1466 (N_1466,In_1902,In_371);
or U1467 (N_1467,In_523,In_736);
xor U1468 (N_1468,In_1477,In_1522);
and U1469 (N_1469,In_252,In_1135);
xor U1470 (N_1470,In_776,In_564);
nand U1471 (N_1471,In_862,In_1166);
xor U1472 (N_1472,In_960,In_495);
or U1473 (N_1473,In_46,In_127);
or U1474 (N_1474,In_1069,In_474);
and U1475 (N_1475,In_381,In_794);
nor U1476 (N_1476,In_1168,In_363);
nor U1477 (N_1477,In_1769,In_1236);
nand U1478 (N_1478,In_680,In_1332);
nand U1479 (N_1479,In_1825,In_1850);
nand U1480 (N_1480,In_188,In_1937);
and U1481 (N_1481,In_1795,In_1165);
and U1482 (N_1482,In_1856,In_1936);
and U1483 (N_1483,In_1825,In_1578);
and U1484 (N_1484,In_1775,In_191);
xor U1485 (N_1485,In_435,In_423);
xnor U1486 (N_1486,In_1569,In_449);
or U1487 (N_1487,In_222,In_627);
nand U1488 (N_1488,In_798,In_1811);
nand U1489 (N_1489,In_1420,In_1912);
xnor U1490 (N_1490,In_1226,In_973);
or U1491 (N_1491,In_1047,In_1819);
nor U1492 (N_1492,In_1360,In_911);
or U1493 (N_1493,In_1819,In_1524);
nand U1494 (N_1494,In_631,In_348);
and U1495 (N_1495,In_1844,In_1719);
nand U1496 (N_1496,In_423,In_1198);
nor U1497 (N_1497,In_324,In_1267);
or U1498 (N_1498,In_621,In_617);
or U1499 (N_1499,In_1495,In_1919);
or U1500 (N_1500,In_1793,In_948);
nor U1501 (N_1501,In_557,In_320);
xor U1502 (N_1502,In_270,In_1078);
and U1503 (N_1503,In_816,In_229);
or U1504 (N_1504,In_115,In_782);
xnor U1505 (N_1505,In_1689,In_1607);
nand U1506 (N_1506,In_889,In_1496);
xnor U1507 (N_1507,In_617,In_62);
xor U1508 (N_1508,In_929,In_198);
nor U1509 (N_1509,In_1494,In_1548);
nor U1510 (N_1510,In_1932,In_513);
xor U1511 (N_1511,In_752,In_1078);
or U1512 (N_1512,In_148,In_1407);
xor U1513 (N_1513,In_1441,In_1462);
and U1514 (N_1514,In_1330,In_506);
or U1515 (N_1515,In_1342,In_1928);
nor U1516 (N_1516,In_1575,In_1435);
nand U1517 (N_1517,In_1562,In_1756);
xnor U1518 (N_1518,In_289,In_252);
or U1519 (N_1519,In_1532,In_787);
nand U1520 (N_1520,In_1604,In_355);
nor U1521 (N_1521,In_585,In_1018);
nand U1522 (N_1522,In_1153,In_492);
nand U1523 (N_1523,In_30,In_598);
nand U1524 (N_1524,In_1848,In_51);
nand U1525 (N_1525,In_1966,In_145);
or U1526 (N_1526,In_566,In_7);
and U1527 (N_1527,In_1069,In_1478);
xnor U1528 (N_1528,In_1954,In_1210);
nand U1529 (N_1529,In_920,In_610);
or U1530 (N_1530,In_859,In_228);
nand U1531 (N_1531,In_947,In_1956);
and U1532 (N_1532,In_1303,In_252);
nand U1533 (N_1533,In_1752,In_842);
nand U1534 (N_1534,In_1731,In_1746);
nor U1535 (N_1535,In_755,In_1435);
nand U1536 (N_1536,In_1795,In_1063);
xor U1537 (N_1537,In_1254,In_1878);
nor U1538 (N_1538,In_52,In_460);
or U1539 (N_1539,In_219,In_1299);
or U1540 (N_1540,In_1200,In_1209);
xnor U1541 (N_1541,In_1276,In_1128);
nand U1542 (N_1542,In_1264,In_931);
nor U1543 (N_1543,In_1524,In_1488);
xor U1544 (N_1544,In_745,In_941);
nor U1545 (N_1545,In_637,In_1472);
nand U1546 (N_1546,In_93,In_1924);
nand U1547 (N_1547,In_1127,In_1960);
or U1548 (N_1548,In_1333,In_999);
xnor U1549 (N_1549,In_1168,In_365);
and U1550 (N_1550,In_1868,In_1299);
nor U1551 (N_1551,In_280,In_1361);
xor U1552 (N_1552,In_847,In_991);
nand U1553 (N_1553,In_847,In_434);
and U1554 (N_1554,In_1013,In_192);
or U1555 (N_1555,In_1875,In_401);
and U1556 (N_1556,In_462,In_350);
or U1557 (N_1557,In_732,In_1220);
or U1558 (N_1558,In_1655,In_219);
nand U1559 (N_1559,In_509,In_503);
xnor U1560 (N_1560,In_1028,In_1949);
or U1561 (N_1561,In_616,In_1665);
xnor U1562 (N_1562,In_1351,In_655);
nand U1563 (N_1563,In_1912,In_1899);
or U1564 (N_1564,In_1148,In_541);
nand U1565 (N_1565,In_330,In_849);
nor U1566 (N_1566,In_250,In_1142);
nand U1567 (N_1567,In_1836,In_1535);
and U1568 (N_1568,In_846,In_1893);
nand U1569 (N_1569,In_69,In_1047);
and U1570 (N_1570,In_821,In_1872);
or U1571 (N_1571,In_814,In_599);
or U1572 (N_1572,In_959,In_1889);
or U1573 (N_1573,In_604,In_250);
xnor U1574 (N_1574,In_1205,In_216);
or U1575 (N_1575,In_1251,In_1727);
or U1576 (N_1576,In_676,In_1656);
nor U1577 (N_1577,In_1341,In_576);
xnor U1578 (N_1578,In_715,In_606);
and U1579 (N_1579,In_457,In_1953);
and U1580 (N_1580,In_1951,In_1520);
and U1581 (N_1581,In_1755,In_952);
nand U1582 (N_1582,In_1485,In_38);
nand U1583 (N_1583,In_631,In_1967);
or U1584 (N_1584,In_623,In_767);
nor U1585 (N_1585,In_1253,In_600);
and U1586 (N_1586,In_1223,In_759);
xnor U1587 (N_1587,In_588,In_1194);
nand U1588 (N_1588,In_707,In_910);
xor U1589 (N_1589,In_924,In_524);
or U1590 (N_1590,In_1375,In_1612);
nand U1591 (N_1591,In_1865,In_1720);
and U1592 (N_1592,In_986,In_1537);
nand U1593 (N_1593,In_225,In_1076);
xor U1594 (N_1594,In_938,In_1620);
or U1595 (N_1595,In_129,In_99);
and U1596 (N_1596,In_49,In_796);
and U1597 (N_1597,In_1361,In_505);
nor U1598 (N_1598,In_1425,In_1417);
nand U1599 (N_1599,In_165,In_611);
and U1600 (N_1600,In_1012,In_902);
nand U1601 (N_1601,In_1705,In_585);
and U1602 (N_1602,In_1469,In_1716);
xnor U1603 (N_1603,In_646,In_678);
xor U1604 (N_1604,In_1167,In_474);
or U1605 (N_1605,In_1007,In_376);
xnor U1606 (N_1606,In_1864,In_209);
nand U1607 (N_1607,In_1761,In_27);
nand U1608 (N_1608,In_894,In_1925);
and U1609 (N_1609,In_722,In_1127);
nand U1610 (N_1610,In_1112,In_1677);
xor U1611 (N_1611,In_537,In_1782);
xnor U1612 (N_1612,In_1610,In_1643);
xor U1613 (N_1613,In_828,In_382);
nand U1614 (N_1614,In_135,In_36);
and U1615 (N_1615,In_47,In_577);
xnor U1616 (N_1616,In_593,In_1530);
or U1617 (N_1617,In_1143,In_627);
xnor U1618 (N_1618,In_312,In_458);
and U1619 (N_1619,In_497,In_513);
and U1620 (N_1620,In_751,In_1308);
and U1621 (N_1621,In_395,In_1413);
nand U1622 (N_1622,In_1425,In_654);
nand U1623 (N_1623,In_1728,In_1474);
or U1624 (N_1624,In_951,In_1344);
and U1625 (N_1625,In_192,In_35);
or U1626 (N_1626,In_1499,In_86);
nor U1627 (N_1627,In_150,In_156);
nor U1628 (N_1628,In_513,In_1611);
nand U1629 (N_1629,In_1219,In_115);
xnor U1630 (N_1630,In_1066,In_1722);
nor U1631 (N_1631,In_792,In_1540);
xnor U1632 (N_1632,In_1315,In_1168);
xnor U1633 (N_1633,In_1008,In_933);
xor U1634 (N_1634,In_151,In_1599);
xnor U1635 (N_1635,In_1935,In_883);
or U1636 (N_1636,In_874,In_1325);
xor U1637 (N_1637,In_46,In_471);
nor U1638 (N_1638,In_253,In_185);
nor U1639 (N_1639,In_1148,In_61);
or U1640 (N_1640,In_1918,In_1398);
xor U1641 (N_1641,In_1750,In_274);
or U1642 (N_1642,In_838,In_941);
nor U1643 (N_1643,In_609,In_557);
nor U1644 (N_1644,In_576,In_1779);
nand U1645 (N_1645,In_1029,In_1960);
nand U1646 (N_1646,In_345,In_833);
and U1647 (N_1647,In_1229,In_1662);
or U1648 (N_1648,In_608,In_68);
or U1649 (N_1649,In_1855,In_421);
nand U1650 (N_1650,In_865,In_805);
and U1651 (N_1651,In_385,In_906);
nand U1652 (N_1652,In_948,In_513);
xor U1653 (N_1653,In_306,In_205);
and U1654 (N_1654,In_875,In_1113);
nand U1655 (N_1655,In_1580,In_875);
and U1656 (N_1656,In_1056,In_16);
xnor U1657 (N_1657,In_1154,In_262);
xor U1658 (N_1658,In_1985,In_318);
or U1659 (N_1659,In_1802,In_1902);
xor U1660 (N_1660,In_899,In_487);
nand U1661 (N_1661,In_1650,In_1836);
or U1662 (N_1662,In_1615,In_362);
nand U1663 (N_1663,In_1177,In_1980);
or U1664 (N_1664,In_365,In_1855);
xnor U1665 (N_1665,In_88,In_950);
nand U1666 (N_1666,In_1456,In_487);
or U1667 (N_1667,In_891,In_389);
xor U1668 (N_1668,In_12,In_264);
and U1669 (N_1669,In_655,In_488);
or U1670 (N_1670,In_234,In_795);
nand U1671 (N_1671,In_837,In_1667);
nor U1672 (N_1672,In_239,In_206);
nor U1673 (N_1673,In_967,In_1952);
or U1674 (N_1674,In_381,In_1421);
or U1675 (N_1675,In_95,In_1929);
or U1676 (N_1676,In_310,In_1656);
nor U1677 (N_1677,In_924,In_1946);
xnor U1678 (N_1678,In_1114,In_645);
nor U1679 (N_1679,In_168,In_874);
nor U1680 (N_1680,In_1457,In_387);
xnor U1681 (N_1681,In_1723,In_1496);
nand U1682 (N_1682,In_1054,In_1119);
and U1683 (N_1683,In_1458,In_1162);
nand U1684 (N_1684,In_1720,In_5);
xor U1685 (N_1685,In_1338,In_132);
nand U1686 (N_1686,In_616,In_1188);
xnor U1687 (N_1687,In_761,In_1742);
and U1688 (N_1688,In_1509,In_851);
or U1689 (N_1689,In_259,In_1217);
nor U1690 (N_1690,In_1558,In_1229);
or U1691 (N_1691,In_962,In_1467);
nor U1692 (N_1692,In_140,In_1122);
nor U1693 (N_1693,In_1038,In_1678);
nand U1694 (N_1694,In_756,In_1355);
xnor U1695 (N_1695,In_1413,In_906);
nand U1696 (N_1696,In_154,In_1128);
nand U1697 (N_1697,In_827,In_1401);
or U1698 (N_1698,In_1627,In_549);
and U1699 (N_1699,In_467,In_1193);
nor U1700 (N_1700,In_1058,In_1780);
nor U1701 (N_1701,In_1595,In_374);
and U1702 (N_1702,In_646,In_341);
nor U1703 (N_1703,In_1382,In_261);
xor U1704 (N_1704,In_1157,In_1744);
or U1705 (N_1705,In_949,In_1582);
and U1706 (N_1706,In_776,In_1531);
nand U1707 (N_1707,In_901,In_909);
nor U1708 (N_1708,In_1598,In_857);
nand U1709 (N_1709,In_1784,In_625);
nor U1710 (N_1710,In_226,In_1287);
xor U1711 (N_1711,In_674,In_658);
nand U1712 (N_1712,In_1585,In_1559);
or U1713 (N_1713,In_161,In_1223);
xor U1714 (N_1714,In_1161,In_480);
nor U1715 (N_1715,In_1501,In_1595);
or U1716 (N_1716,In_1668,In_1764);
or U1717 (N_1717,In_1073,In_1838);
and U1718 (N_1718,In_1942,In_475);
and U1719 (N_1719,In_1972,In_1132);
nor U1720 (N_1720,In_723,In_594);
xnor U1721 (N_1721,In_1610,In_1413);
and U1722 (N_1722,In_1314,In_43);
and U1723 (N_1723,In_282,In_539);
nor U1724 (N_1724,In_94,In_791);
nand U1725 (N_1725,In_892,In_1917);
nand U1726 (N_1726,In_1137,In_1431);
nand U1727 (N_1727,In_1083,In_1438);
and U1728 (N_1728,In_1689,In_1185);
or U1729 (N_1729,In_1605,In_527);
nand U1730 (N_1730,In_1440,In_772);
xnor U1731 (N_1731,In_1856,In_1423);
nand U1732 (N_1732,In_1721,In_748);
nor U1733 (N_1733,In_1326,In_746);
and U1734 (N_1734,In_1014,In_1257);
and U1735 (N_1735,In_658,In_1909);
nand U1736 (N_1736,In_1747,In_63);
nor U1737 (N_1737,In_1314,In_515);
nand U1738 (N_1738,In_785,In_429);
nand U1739 (N_1739,In_1344,In_1159);
nand U1740 (N_1740,In_1776,In_1289);
xor U1741 (N_1741,In_887,In_1597);
or U1742 (N_1742,In_495,In_1209);
xnor U1743 (N_1743,In_1115,In_855);
nand U1744 (N_1744,In_320,In_1218);
xor U1745 (N_1745,In_928,In_1095);
and U1746 (N_1746,In_1106,In_212);
nand U1747 (N_1747,In_411,In_358);
nor U1748 (N_1748,In_94,In_1983);
nor U1749 (N_1749,In_1883,In_864);
nand U1750 (N_1750,In_1973,In_1264);
nor U1751 (N_1751,In_1104,In_186);
and U1752 (N_1752,In_838,In_701);
nor U1753 (N_1753,In_389,In_1100);
or U1754 (N_1754,In_1038,In_245);
nand U1755 (N_1755,In_1965,In_1316);
and U1756 (N_1756,In_776,In_198);
nor U1757 (N_1757,In_1945,In_40);
nand U1758 (N_1758,In_1721,In_346);
xor U1759 (N_1759,In_1647,In_59);
or U1760 (N_1760,In_1164,In_1266);
nand U1761 (N_1761,In_1693,In_1347);
or U1762 (N_1762,In_173,In_841);
xor U1763 (N_1763,In_1556,In_1800);
and U1764 (N_1764,In_108,In_267);
nor U1765 (N_1765,In_1696,In_506);
or U1766 (N_1766,In_1623,In_655);
nand U1767 (N_1767,In_278,In_728);
and U1768 (N_1768,In_131,In_167);
nor U1769 (N_1769,In_226,In_1805);
xnor U1770 (N_1770,In_1676,In_1013);
or U1771 (N_1771,In_1959,In_246);
and U1772 (N_1772,In_1149,In_1733);
or U1773 (N_1773,In_34,In_1345);
nor U1774 (N_1774,In_806,In_392);
nor U1775 (N_1775,In_668,In_1659);
and U1776 (N_1776,In_1674,In_362);
nor U1777 (N_1777,In_1014,In_1213);
or U1778 (N_1778,In_1591,In_1394);
or U1779 (N_1779,In_1625,In_1082);
xnor U1780 (N_1780,In_1591,In_646);
or U1781 (N_1781,In_1312,In_296);
xnor U1782 (N_1782,In_1115,In_1414);
or U1783 (N_1783,In_1997,In_12);
nand U1784 (N_1784,In_1741,In_1958);
and U1785 (N_1785,In_595,In_100);
nand U1786 (N_1786,In_53,In_550);
or U1787 (N_1787,In_780,In_1928);
xor U1788 (N_1788,In_1410,In_1623);
nor U1789 (N_1789,In_1573,In_315);
xor U1790 (N_1790,In_172,In_323);
xnor U1791 (N_1791,In_1403,In_1557);
nand U1792 (N_1792,In_176,In_1304);
nand U1793 (N_1793,In_1849,In_909);
nand U1794 (N_1794,In_236,In_1688);
nand U1795 (N_1795,In_364,In_1309);
and U1796 (N_1796,In_1489,In_403);
or U1797 (N_1797,In_12,In_1878);
nor U1798 (N_1798,In_376,In_748);
xor U1799 (N_1799,In_1589,In_1280);
nand U1800 (N_1800,In_1269,In_1129);
nor U1801 (N_1801,In_820,In_1569);
and U1802 (N_1802,In_855,In_512);
nor U1803 (N_1803,In_441,In_756);
nand U1804 (N_1804,In_13,In_1979);
xor U1805 (N_1805,In_180,In_185);
nor U1806 (N_1806,In_11,In_682);
nor U1807 (N_1807,In_920,In_97);
xor U1808 (N_1808,In_1192,In_1071);
xnor U1809 (N_1809,In_81,In_1020);
and U1810 (N_1810,In_1363,In_1169);
nand U1811 (N_1811,In_1597,In_1760);
xnor U1812 (N_1812,In_13,In_1995);
or U1813 (N_1813,In_967,In_152);
nand U1814 (N_1814,In_1809,In_889);
nor U1815 (N_1815,In_402,In_537);
or U1816 (N_1816,In_1623,In_734);
and U1817 (N_1817,In_332,In_1357);
xor U1818 (N_1818,In_400,In_1383);
xor U1819 (N_1819,In_708,In_1798);
or U1820 (N_1820,In_536,In_715);
nand U1821 (N_1821,In_1879,In_1062);
and U1822 (N_1822,In_1488,In_348);
xor U1823 (N_1823,In_419,In_1567);
nor U1824 (N_1824,In_1626,In_1251);
nor U1825 (N_1825,In_739,In_1105);
and U1826 (N_1826,In_487,In_279);
xnor U1827 (N_1827,In_1942,In_672);
and U1828 (N_1828,In_1243,In_375);
nand U1829 (N_1829,In_1531,In_1440);
nor U1830 (N_1830,In_664,In_330);
and U1831 (N_1831,In_1716,In_182);
xor U1832 (N_1832,In_1853,In_1270);
nand U1833 (N_1833,In_667,In_261);
nor U1834 (N_1834,In_103,In_985);
xor U1835 (N_1835,In_1385,In_395);
and U1836 (N_1836,In_1264,In_954);
or U1837 (N_1837,In_178,In_1590);
nor U1838 (N_1838,In_655,In_817);
nand U1839 (N_1839,In_1961,In_180);
xor U1840 (N_1840,In_282,In_747);
nor U1841 (N_1841,In_758,In_472);
or U1842 (N_1842,In_949,In_837);
or U1843 (N_1843,In_1463,In_995);
or U1844 (N_1844,In_685,In_1769);
nor U1845 (N_1845,In_1058,In_1610);
and U1846 (N_1846,In_364,In_60);
xor U1847 (N_1847,In_1802,In_1501);
and U1848 (N_1848,In_1799,In_1914);
or U1849 (N_1849,In_1293,In_1968);
nand U1850 (N_1850,In_683,In_579);
and U1851 (N_1851,In_1146,In_1505);
nor U1852 (N_1852,In_1521,In_216);
xnor U1853 (N_1853,In_213,In_569);
nor U1854 (N_1854,In_1466,In_341);
xor U1855 (N_1855,In_1295,In_682);
nor U1856 (N_1856,In_769,In_1941);
nand U1857 (N_1857,In_304,In_350);
and U1858 (N_1858,In_922,In_870);
nand U1859 (N_1859,In_1842,In_457);
nor U1860 (N_1860,In_1990,In_753);
xor U1861 (N_1861,In_1452,In_1974);
xnor U1862 (N_1862,In_538,In_308);
and U1863 (N_1863,In_193,In_923);
nand U1864 (N_1864,In_1295,In_26);
xnor U1865 (N_1865,In_1534,In_1558);
and U1866 (N_1866,In_1113,In_1793);
nor U1867 (N_1867,In_185,In_1360);
or U1868 (N_1868,In_1944,In_1082);
or U1869 (N_1869,In_1069,In_424);
nor U1870 (N_1870,In_1166,In_507);
or U1871 (N_1871,In_1783,In_1627);
nor U1872 (N_1872,In_1184,In_1304);
xnor U1873 (N_1873,In_1805,In_1104);
xnor U1874 (N_1874,In_897,In_974);
or U1875 (N_1875,In_1402,In_1619);
nor U1876 (N_1876,In_974,In_1267);
nor U1877 (N_1877,In_1979,In_1331);
or U1878 (N_1878,In_1195,In_166);
nor U1879 (N_1879,In_71,In_491);
and U1880 (N_1880,In_1486,In_1508);
xnor U1881 (N_1881,In_1484,In_838);
and U1882 (N_1882,In_631,In_1762);
or U1883 (N_1883,In_931,In_1549);
and U1884 (N_1884,In_83,In_1292);
nand U1885 (N_1885,In_1826,In_1124);
nor U1886 (N_1886,In_591,In_1130);
or U1887 (N_1887,In_381,In_1035);
or U1888 (N_1888,In_1976,In_566);
and U1889 (N_1889,In_347,In_689);
nor U1890 (N_1890,In_1088,In_448);
nand U1891 (N_1891,In_647,In_1375);
nand U1892 (N_1892,In_485,In_621);
nor U1893 (N_1893,In_699,In_1597);
nand U1894 (N_1894,In_1403,In_184);
nand U1895 (N_1895,In_280,In_1038);
nand U1896 (N_1896,In_1712,In_313);
or U1897 (N_1897,In_95,In_1605);
nor U1898 (N_1898,In_1755,In_229);
or U1899 (N_1899,In_1008,In_1781);
nand U1900 (N_1900,In_935,In_316);
and U1901 (N_1901,In_1103,In_906);
nor U1902 (N_1902,In_1427,In_1919);
or U1903 (N_1903,In_851,In_1827);
or U1904 (N_1904,In_990,In_56);
xnor U1905 (N_1905,In_975,In_1915);
or U1906 (N_1906,In_73,In_226);
and U1907 (N_1907,In_881,In_479);
xor U1908 (N_1908,In_1675,In_1622);
and U1909 (N_1909,In_1819,In_147);
nor U1910 (N_1910,In_1319,In_1011);
and U1911 (N_1911,In_1981,In_824);
nand U1912 (N_1912,In_390,In_241);
nor U1913 (N_1913,In_829,In_1435);
and U1914 (N_1914,In_1478,In_32);
nand U1915 (N_1915,In_1114,In_1580);
nand U1916 (N_1916,In_1275,In_1976);
and U1917 (N_1917,In_62,In_35);
and U1918 (N_1918,In_1157,In_314);
xor U1919 (N_1919,In_1192,In_286);
nor U1920 (N_1920,In_794,In_1719);
xor U1921 (N_1921,In_1645,In_1397);
nor U1922 (N_1922,In_526,In_196);
and U1923 (N_1923,In_828,In_172);
nand U1924 (N_1924,In_460,In_360);
nand U1925 (N_1925,In_5,In_166);
nand U1926 (N_1926,In_816,In_285);
nand U1927 (N_1927,In_1439,In_480);
nor U1928 (N_1928,In_364,In_652);
nand U1929 (N_1929,In_1982,In_76);
or U1930 (N_1930,In_40,In_419);
or U1931 (N_1931,In_226,In_270);
nor U1932 (N_1932,In_70,In_126);
nand U1933 (N_1933,In_400,In_1732);
xor U1934 (N_1934,In_217,In_124);
nand U1935 (N_1935,In_595,In_1588);
and U1936 (N_1936,In_125,In_653);
and U1937 (N_1937,In_819,In_664);
xor U1938 (N_1938,In_1276,In_10);
nand U1939 (N_1939,In_747,In_948);
nand U1940 (N_1940,In_1621,In_776);
nor U1941 (N_1941,In_741,In_1177);
nor U1942 (N_1942,In_1233,In_1091);
nor U1943 (N_1943,In_1126,In_778);
xnor U1944 (N_1944,In_930,In_1583);
nor U1945 (N_1945,In_1087,In_360);
xor U1946 (N_1946,In_1672,In_132);
xnor U1947 (N_1947,In_824,In_1598);
or U1948 (N_1948,In_1612,In_502);
xor U1949 (N_1949,In_1814,In_1328);
xor U1950 (N_1950,In_1313,In_1822);
nand U1951 (N_1951,In_1070,In_1572);
and U1952 (N_1952,In_204,In_1834);
nand U1953 (N_1953,In_1025,In_914);
nor U1954 (N_1954,In_346,In_560);
nand U1955 (N_1955,In_637,In_1934);
nor U1956 (N_1956,In_1479,In_1915);
or U1957 (N_1957,In_94,In_1000);
nand U1958 (N_1958,In_772,In_354);
or U1959 (N_1959,In_160,In_980);
and U1960 (N_1960,In_324,In_769);
or U1961 (N_1961,In_22,In_1884);
xnor U1962 (N_1962,In_1648,In_222);
or U1963 (N_1963,In_37,In_405);
or U1964 (N_1964,In_1308,In_552);
or U1965 (N_1965,In_1751,In_1989);
and U1966 (N_1966,In_191,In_1865);
nor U1967 (N_1967,In_327,In_1344);
nand U1968 (N_1968,In_339,In_1906);
nand U1969 (N_1969,In_493,In_1500);
or U1970 (N_1970,In_461,In_1741);
nand U1971 (N_1971,In_1123,In_786);
nand U1972 (N_1972,In_1592,In_167);
or U1973 (N_1973,In_1811,In_1223);
or U1974 (N_1974,In_420,In_1417);
or U1975 (N_1975,In_1421,In_650);
nand U1976 (N_1976,In_23,In_283);
xnor U1977 (N_1977,In_102,In_1714);
nor U1978 (N_1978,In_744,In_1329);
and U1979 (N_1979,In_1190,In_851);
or U1980 (N_1980,In_1371,In_1247);
or U1981 (N_1981,In_427,In_1225);
nand U1982 (N_1982,In_1606,In_1118);
xnor U1983 (N_1983,In_1019,In_360);
nor U1984 (N_1984,In_1845,In_1361);
xor U1985 (N_1985,In_334,In_1705);
xnor U1986 (N_1986,In_1498,In_1185);
xor U1987 (N_1987,In_1773,In_1162);
and U1988 (N_1988,In_34,In_1058);
or U1989 (N_1989,In_1159,In_1112);
and U1990 (N_1990,In_247,In_1361);
or U1991 (N_1991,In_834,In_1123);
or U1992 (N_1992,In_80,In_217);
or U1993 (N_1993,In_886,In_1895);
and U1994 (N_1994,In_1149,In_1496);
nand U1995 (N_1995,In_1018,In_661);
nor U1996 (N_1996,In_858,In_275);
and U1997 (N_1997,In_529,In_43);
or U1998 (N_1998,In_66,In_293);
nand U1999 (N_1999,In_343,In_746);
xnor U2000 (N_2000,In_1676,In_1905);
xnor U2001 (N_2001,In_1813,In_1498);
or U2002 (N_2002,In_243,In_1863);
or U2003 (N_2003,In_1367,In_1063);
or U2004 (N_2004,In_372,In_1413);
nand U2005 (N_2005,In_1079,In_1870);
xnor U2006 (N_2006,In_60,In_1007);
xor U2007 (N_2007,In_1028,In_436);
nand U2008 (N_2008,In_1012,In_41);
or U2009 (N_2009,In_513,In_1215);
xor U2010 (N_2010,In_1983,In_1333);
nand U2011 (N_2011,In_1879,In_161);
nand U2012 (N_2012,In_623,In_1211);
nand U2013 (N_2013,In_1954,In_1464);
nand U2014 (N_2014,In_73,In_799);
xor U2015 (N_2015,In_1107,In_1741);
or U2016 (N_2016,In_1048,In_1140);
xnor U2017 (N_2017,In_1062,In_877);
or U2018 (N_2018,In_853,In_1284);
or U2019 (N_2019,In_351,In_388);
and U2020 (N_2020,In_312,In_151);
xor U2021 (N_2021,In_982,In_282);
and U2022 (N_2022,In_343,In_437);
nand U2023 (N_2023,In_1811,In_1832);
and U2024 (N_2024,In_1691,In_1687);
or U2025 (N_2025,In_345,In_1767);
and U2026 (N_2026,In_973,In_1109);
nand U2027 (N_2027,In_234,In_1218);
nor U2028 (N_2028,In_1278,In_1036);
and U2029 (N_2029,In_154,In_339);
or U2030 (N_2030,In_101,In_1306);
nor U2031 (N_2031,In_583,In_1678);
nor U2032 (N_2032,In_52,In_1928);
or U2033 (N_2033,In_1682,In_1221);
and U2034 (N_2034,In_999,In_1968);
and U2035 (N_2035,In_1491,In_255);
xor U2036 (N_2036,In_148,In_1944);
or U2037 (N_2037,In_22,In_1905);
nor U2038 (N_2038,In_24,In_1779);
and U2039 (N_2039,In_1966,In_719);
and U2040 (N_2040,In_1227,In_1244);
or U2041 (N_2041,In_13,In_1890);
or U2042 (N_2042,In_656,In_1251);
nand U2043 (N_2043,In_687,In_1762);
nand U2044 (N_2044,In_1950,In_397);
xnor U2045 (N_2045,In_1938,In_1842);
nor U2046 (N_2046,In_640,In_1481);
and U2047 (N_2047,In_872,In_1484);
xnor U2048 (N_2048,In_1185,In_392);
and U2049 (N_2049,In_154,In_1156);
nand U2050 (N_2050,In_1,In_1522);
and U2051 (N_2051,In_1794,In_1275);
nor U2052 (N_2052,In_1228,In_1198);
nor U2053 (N_2053,In_501,In_812);
nand U2054 (N_2054,In_472,In_848);
nor U2055 (N_2055,In_1627,In_1740);
or U2056 (N_2056,In_1452,In_301);
or U2057 (N_2057,In_283,In_1698);
and U2058 (N_2058,In_230,In_559);
and U2059 (N_2059,In_927,In_1551);
nand U2060 (N_2060,In_577,In_994);
xor U2061 (N_2061,In_990,In_1282);
or U2062 (N_2062,In_216,In_553);
or U2063 (N_2063,In_1081,In_1432);
nand U2064 (N_2064,In_1983,In_1729);
or U2065 (N_2065,In_402,In_1956);
xnor U2066 (N_2066,In_661,In_1447);
nor U2067 (N_2067,In_465,In_957);
nor U2068 (N_2068,In_1034,In_1594);
xnor U2069 (N_2069,In_1645,In_466);
and U2070 (N_2070,In_1933,In_1774);
or U2071 (N_2071,In_1096,In_644);
nor U2072 (N_2072,In_444,In_33);
nor U2073 (N_2073,In_283,In_1525);
and U2074 (N_2074,In_1482,In_1194);
or U2075 (N_2075,In_518,In_1951);
or U2076 (N_2076,In_1363,In_1245);
nor U2077 (N_2077,In_171,In_71);
nand U2078 (N_2078,In_1834,In_28);
nor U2079 (N_2079,In_1549,In_111);
nor U2080 (N_2080,In_986,In_749);
xnor U2081 (N_2081,In_1838,In_1827);
and U2082 (N_2082,In_1846,In_969);
nor U2083 (N_2083,In_1422,In_1971);
nor U2084 (N_2084,In_1130,In_770);
nand U2085 (N_2085,In_1388,In_1237);
or U2086 (N_2086,In_1617,In_1731);
and U2087 (N_2087,In_293,In_1969);
nor U2088 (N_2088,In_356,In_514);
nor U2089 (N_2089,In_1500,In_82);
and U2090 (N_2090,In_1363,In_956);
nand U2091 (N_2091,In_1366,In_1766);
nand U2092 (N_2092,In_806,In_912);
and U2093 (N_2093,In_349,In_70);
or U2094 (N_2094,In_196,In_784);
or U2095 (N_2095,In_1267,In_1164);
or U2096 (N_2096,In_756,In_1269);
nor U2097 (N_2097,In_872,In_1816);
nand U2098 (N_2098,In_844,In_1445);
xnor U2099 (N_2099,In_1766,In_1466);
xor U2100 (N_2100,In_1675,In_831);
and U2101 (N_2101,In_496,In_1994);
nand U2102 (N_2102,In_281,In_1000);
and U2103 (N_2103,In_833,In_1231);
xor U2104 (N_2104,In_226,In_512);
or U2105 (N_2105,In_1348,In_322);
or U2106 (N_2106,In_896,In_389);
or U2107 (N_2107,In_1825,In_334);
nor U2108 (N_2108,In_1848,In_1710);
nand U2109 (N_2109,In_462,In_1914);
and U2110 (N_2110,In_570,In_940);
nor U2111 (N_2111,In_1559,In_444);
or U2112 (N_2112,In_647,In_896);
nor U2113 (N_2113,In_1738,In_1197);
xor U2114 (N_2114,In_364,In_960);
or U2115 (N_2115,In_889,In_834);
nand U2116 (N_2116,In_387,In_1589);
xor U2117 (N_2117,In_1445,In_179);
xor U2118 (N_2118,In_1162,In_427);
xnor U2119 (N_2119,In_641,In_1757);
nand U2120 (N_2120,In_1772,In_802);
and U2121 (N_2121,In_1245,In_1213);
or U2122 (N_2122,In_197,In_1757);
and U2123 (N_2123,In_1664,In_945);
and U2124 (N_2124,In_627,In_642);
nor U2125 (N_2125,In_1773,In_1980);
and U2126 (N_2126,In_707,In_587);
nor U2127 (N_2127,In_1042,In_169);
nor U2128 (N_2128,In_362,In_1841);
or U2129 (N_2129,In_1062,In_302);
and U2130 (N_2130,In_1952,In_21);
xnor U2131 (N_2131,In_1048,In_1625);
xor U2132 (N_2132,In_762,In_341);
nor U2133 (N_2133,In_28,In_1694);
nand U2134 (N_2134,In_1908,In_547);
xnor U2135 (N_2135,In_1354,In_224);
xor U2136 (N_2136,In_1629,In_143);
nor U2137 (N_2137,In_1724,In_1065);
xor U2138 (N_2138,In_697,In_1044);
or U2139 (N_2139,In_758,In_1256);
and U2140 (N_2140,In_1294,In_1719);
nor U2141 (N_2141,In_1175,In_1067);
or U2142 (N_2142,In_4,In_1783);
and U2143 (N_2143,In_1514,In_755);
xor U2144 (N_2144,In_1109,In_1960);
and U2145 (N_2145,In_568,In_261);
and U2146 (N_2146,In_246,In_670);
and U2147 (N_2147,In_1192,In_814);
nand U2148 (N_2148,In_473,In_1499);
or U2149 (N_2149,In_1771,In_719);
nand U2150 (N_2150,In_1713,In_627);
xor U2151 (N_2151,In_1307,In_1744);
nand U2152 (N_2152,In_730,In_1507);
nor U2153 (N_2153,In_1168,In_164);
nor U2154 (N_2154,In_235,In_640);
nor U2155 (N_2155,In_1010,In_1243);
xor U2156 (N_2156,In_1054,In_1599);
xor U2157 (N_2157,In_478,In_190);
xor U2158 (N_2158,In_1835,In_749);
or U2159 (N_2159,In_891,In_525);
or U2160 (N_2160,In_1242,In_1178);
nor U2161 (N_2161,In_1831,In_1673);
and U2162 (N_2162,In_1924,In_976);
xnor U2163 (N_2163,In_711,In_1949);
and U2164 (N_2164,In_926,In_1753);
or U2165 (N_2165,In_1780,In_1999);
nor U2166 (N_2166,In_1745,In_1817);
xnor U2167 (N_2167,In_960,In_33);
or U2168 (N_2168,In_540,In_1914);
or U2169 (N_2169,In_991,In_105);
and U2170 (N_2170,In_1420,In_872);
xor U2171 (N_2171,In_1822,In_521);
or U2172 (N_2172,In_1749,In_1897);
and U2173 (N_2173,In_1927,In_551);
and U2174 (N_2174,In_1983,In_788);
xor U2175 (N_2175,In_1135,In_951);
and U2176 (N_2176,In_1919,In_1657);
and U2177 (N_2177,In_617,In_794);
nand U2178 (N_2178,In_1775,In_416);
xor U2179 (N_2179,In_872,In_74);
and U2180 (N_2180,In_822,In_91);
nor U2181 (N_2181,In_1317,In_1958);
nor U2182 (N_2182,In_320,In_1011);
xnor U2183 (N_2183,In_1381,In_1326);
xnor U2184 (N_2184,In_1005,In_717);
or U2185 (N_2185,In_186,In_1259);
or U2186 (N_2186,In_391,In_1622);
or U2187 (N_2187,In_1633,In_1622);
or U2188 (N_2188,In_1915,In_604);
xnor U2189 (N_2189,In_1719,In_763);
or U2190 (N_2190,In_375,In_793);
nand U2191 (N_2191,In_1941,In_1998);
nor U2192 (N_2192,In_982,In_1305);
and U2193 (N_2193,In_127,In_1700);
nor U2194 (N_2194,In_1108,In_767);
and U2195 (N_2195,In_1084,In_102);
nand U2196 (N_2196,In_1136,In_654);
nor U2197 (N_2197,In_698,In_1863);
xnor U2198 (N_2198,In_1233,In_43);
xnor U2199 (N_2199,In_1865,In_1831);
xnor U2200 (N_2200,In_578,In_11);
xnor U2201 (N_2201,In_1339,In_1476);
and U2202 (N_2202,In_1919,In_1451);
xor U2203 (N_2203,In_1530,In_1152);
nor U2204 (N_2204,In_1671,In_1925);
xnor U2205 (N_2205,In_913,In_860);
nand U2206 (N_2206,In_1709,In_910);
and U2207 (N_2207,In_1541,In_800);
and U2208 (N_2208,In_1369,In_1665);
and U2209 (N_2209,In_709,In_1146);
and U2210 (N_2210,In_1947,In_1637);
nand U2211 (N_2211,In_1941,In_1243);
xor U2212 (N_2212,In_945,In_1977);
nor U2213 (N_2213,In_1964,In_1102);
nor U2214 (N_2214,In_953,In_1195);
and U2215 (N_2215,In_790,In_345);
and U2216 (N_2216,In_94,In_1858);
nor U2217 (N_2217,In_1874,In_717);
nand U2218 (N_2218,In_1185,In_1968);
or U2219 (N_2219,In_584,In_1598);
and U2220 (N_2220,In_1400,In_873);
xnor U2221 (N_2221,In_1593,In_1063);
nand U2222 (N_2222,In_871,In_144);
and U2223 (N_2223,In_1757,In_1591);
nand U2224 (N_2224,In_1445,In_250);
or U2225 (N_2225,In_1350,In_1360);
and U2226 (N_2226,In_491,In_275);
and U2227 (N_2227,In_1422,In_1130);
and U2228 (N_2228,In_1752,In_419);
or U2229 (N_2229,In_607,In_649);
and U2230 (N_2230,In_1908,In_721);
nand U2231 (N_2231,In_1059,In_213);
and U2232 (N_2232,In_1817,In_1356);
and U2233 (N_2233,In_261,In_841);
xnor U2234 (N_2234,In_15,In_352);
xor U2235 (N_2235,In_863,In_771);
or U2236 (N_2236,In_749,In_556);
nand U2237 (N_2237,In_381,In_201);
or U2238 (N_2238,In_1022,In_1480);
and U2239 (N_2239,In_1980,In_1353);
xor U2240 (N_2240,In_86,In_1349);
nor U2241 (N_2241,In_908,In_326);
nor U2242 (N_2242,In_768,In_1859);
and U2243 (N_2243,In_137,In_1853);
or U2244 (N_2244,In_772,In_1304);
xor U2245 (N_2245,In_1773,In_1943);
nor U2246 (N_2246,In_820,In_694);
nand U2247 (N_2247,In_235,In_1722);
and U2248 (N_2248,In_1889,In_1512);
xnor U2249 (N_2249,In_1607,In_1044);
nor U2250 (N_2250,In_338,In_1069);
or U2251 (N_2251,In_13,In_238);
nand U2252 (N_2252,In_659,In_1648);
nand U2253 (N_2253,In_1142,In_1341);
nand U2254 (N_2254,In_532,In_10);
nor U2255 (N_2255,In_224,In_1125);
xor U2256 (N_2256,In_1041,In_957);
nor U2257 (N_2257,In_1954,In_1109);
or U2258 (N_2258,In_1673,In_574);
or U2259 (N_2259,In_1926,In_679);
nand U2260 (N_2260,In_919,In_968);
and U2261 (N_2261,In_484,In_1867);
nor U2262 (N_2262,In_875,In_473);
xor U2263 (N_2263,In_909,In_1143);
xor U2264 (N_2264,In_1556,In_519);
nand U2265 (N_2265,In_1071,In_1028);
or U2266 (N_2266,In_867,In_242);
xnor U2267 (N_2267,In_667,In_1320);
and U2268 (N_2268,In_286,In_1306);
nor U2269 (N_2269,In_798,In_1912);
and U2270 (N_2270,In_329,In_755);
nor U2271 (N_2271,In_1257,In_1728);
nor U2272 (N_2272,In_1622,In_173);
and U2273 (N_2273,In_489,In_324);
or U2274 (N_2274,In_254,In_1637);
or U2275 (N_2275,In_547,In_1670);
nand U2276 (N_2276,In_1319,In_488);
and U2277 (N_2277,In_1636,In_328);
xnor U2278 (N_2278,In_629,In_512);
xnor U2279 (N_2279,In_668,In_1935);
and U2280 (N_2280,In_459,In_528);
or U2281 (N_2281,In_1850,In_1122);
nand U2282 (N_2282,In_1208,In_194);
nand U2283 (N_2283,In_461,In_705);
nor U2284 (N_2284,In_223,In_1480);
nor U2285 (N_2285,In_1703,In_1941);
xnor U2286 (N_2286,In_914,In_1132);
nor U2287 (N_2287,In_454,In_705);
nand U2288 (N_2288,In_852,In_1567);
xor U2289 (N_2289,In_15,In_960);
xor U2290 (N_2290,In_522,In_1851);
and U2291 (N_2291,In_1620,In_366);
and U2292 (N_2292,In_108,In_363);
nand U2293 (N_2293,In_1599,In_1580);
nand U2294 (N_2294,In_1516,In_662);
nand U2295 (N_2295,In_1289,In_1503);
and U2296 (N_2296,In_179,In_251);
xor U2297 (N_2297,In_1459,In_82);
nand U2298 (N_2298,In_814,In_1840);
nand U2299 (N_2299,In_1894,In_1316);
nand U2300 (N_2300,In_487,In_1834);
nor U2301 (N_2301,In_1456,In_1527);
nor U2302 (N_2302,In_446,In_973);
xnor U2303 (N_2303,In_1976,In_600);
and U2304 (N_2304,In_422,In_1085);
or U2305 (N_2305,In_1253,In_504);
xnor U2306 (N_2306,In_348,In_1473);
and U2307 (N_2307,In_169,In_1655);
nor U2308 (N_2308,In_62,In_598);
or U2309 (N_2309,In_1288,In_1702);
and U2310 (N_2310,In_826,In_1392);
nor U2311 (N_2311,In_1176,In_1289);
nand U2312 (N_2312,In_1834,In_18);
nand U2313 (N_2313,In_1366,In_177);
xnor U2314 (N_2314,In_1100,In_1201);
xnor U2315 (N_2315,In_739,In_1772);
or U2316 (N_2316,In_240,In_1159);
xor U2317 (N_2317,In_74,In_385);
and U2318 (N_2318,In_1516,In_1611);
nor U2319 (N_2319,In_1389,In_153);
or U2320 (N_2320,In_1409,In_1851);
and U2321 (N_2321,In_1477,In_844);
nor U2322 (N_2322,In_268,In_337);
xnor U2323 (N_2323,In_1837,In_1741);
or U2324 (N_2324,In_1067,In_71);
or U2325 (N_2325,In_1753,In_202);
xnor U2326 (N_2326,In_464,In_326);
nor U2327 (N_2327,In_205,In_1517);
and U2328 (N_2328,In_1753,In_1575);
nand U2329 (N_2329,In_1950,In_342);
nor U2330 (N_2330,In_507,In_983);
xor U2331 (N_2331,In_1359,In_1292);
and U2332 (N_2332,In_640,In_21);
nor U2333 (N_2333,In_1197,In_1500);
nor U2334 (N_2334,In_1346,In_1645);
nor U2335 (N_2335,In_1215,In_458);
and U2336 (N_2336,In_1936,In_1878);
xor U2337 (N_2337,In_1748,In_1173);
nor U2338 (N_2338,In_598,In_1207);
and U2339 (N_2339,In_1123,In_435);
and U2340 (N_2340,In_475,In_234);
nor U2341 (N_2341,In_1965,In_1613);
or U2342 (N_2342,In_666,In_366);
or U2343 (N_2343,In_1429,In_1025);
nand U2344 (N_2344,In_1659,In_725);
nand U2345 (N_2345,In_453,In_442);
or U2346 (N_2346,In_255,In_683);
nor U2347 (N_2347,In_1578,In_411);
and U2348 (N_2348,In_767,In_1098);
xnor U2349 (N_2349,In_1989,In_1926);
nor U2350 (N_2350,In_1926,In_1368);
nor U2351 (N_2351,In_1608,In_1388);
nand U2352 (N_2352,In_141,In_402);
and U2353 (N_2353,In_1343,In_1701);
nor U2354 (N_2354,In_193,In_1144);
xnor U2355 (N_2355,In_1486,In_496);
nor U2356 (N_2356,In_203,In_469);
xnor U2357 (N_2357,In_530,In_764);
and U2358 (N_2358,In_1260,In_1461);
xnor U2359 (N_2359,In_212,In_241);
nor U2360 (N_2360,In_701,In_1306);
nor U2361 (N_2361,In_597,In_1165);
nand U2362 (N_2362,In_575,In_1105);
nand U2363 (N_2363,In_349,In_131);
or U2364 (N_2364,In_1195,In_187);
xnor U2365 (N_2365,In_946,In_1855);
and U2366 (N_2366,In_344,In_1526);
nand U2367 (N_2367,In_1586,In_1048);
nor U2368 (N_2368,In_1536,In_1458);
xor U2369 (N_2369,In_304,In_1866);
xor U2370 (N_2370,In_1323,In_895);
nor U2371 (N_2371,In_326,In_334);
nor U2372 (N_2372,In_887,In_1069);
and U2373 (N_2373,In_1378,In_625);
or U2374 (N_2374,In_722,In_1385);
nand U2375 (N_2375,In_1502,In_444);
or U2376 (N_2376,In_1027,In_38);
or U2377 (N_2377,In_1103,In_1087);
or U2378 (N_2378,In_1049,In_1184);
xnor U2379 (N_2379,In_292,In_1831);
xnor U2380 (N_2380,In_710,In_505);
and U2381 (N_2381,In_1630,In_178);
nand U2382 (N_2382,In_976,In_670);
nor U2383 (N_2383,In_1255,In_1928);
and U2384 (N_2384,In_702,In_1955);
nand U2385 (N_2385,In_1787,In_289);
nor U2386 (N_2386,In_858,In_1766);
or U2387 (N_2387,In_587,In_799);
nor U2388 (N_2388,In_1662,In_1311);
and U2389 (N_2389,In_1930,In_1293);
or U2390 (N_2390,In_1747,In_265);
xor U2391 (N_2391,In_1251,In_745);
and U2392 (N_2392,In_87,In_1248);
and U2393 (N_2393,In_544,In_1357);
nor U2394 (N_2394,In_1921,In_1172);
xnor U2395 (N_2395,In_56,In_1152);
nor U2396 (N_2396,In_893,In_1456);
and U2397 (N_2397,In_1160,In_499);
or U2398 (N_2398,In_1168,In_1278);
or U2399 (N_2399,In_1602,In_1950);
and U2400 (N_2400,In_1109,In_1641);
xor U2401 (N_2401,In_1895,In_1584);
and U2402 (N_2402,In_1733,In_1825);
and U2403 (N_2403,In_1982,In_916);
nor U2404 (N_2404,In_95,In_272);
or U2405 (N_2405,In_1110,In_205);
nor U2406 (N_2406,In_265,In_1221);
and U2407 (N_2407,In_1168,In_1740);
or U2408 (N_2408,In_212,In_1473);
or U2409 (N_2409,In_190,In_1773);
xnor U2410 (N_2410,In_416,In_859);
xnor U2411 (N_2411,In_309,In_707);
and U2412 (N_2412,In_1078,In_74);
nor U2413 (N_2413,In_1152,In_1970);
and U2414 (N_2414,In_1501,In_1144);
nor U2415 (N_2415,In_1564,In_1542);
and U2416 (N_2416,In_814,In_1679);
xor U2417 (N_2417,In_1794,In_572);
xnor U2418 (N_2418,In_1068,In_126);
or U2419 (N_2419,In_1151,In_709);
nand U2420 (N_2420,In_166,In_45);
or U2421 (N_2421,In_1343,In_1950);
xor U2422 (N_2422,In_277,In_1084);
or U2423 (N_2423,In_1054,In_1472);
and U2424 (N_2424,In_363,In_1639);
nor U2425 (N_2425,In_1406,In_968);
nand U2426 (N_2426,In_1918,In_824);
xor U2427 (N_2427,In_329,In_561);
xor U2428 (N_2428,In_826,In_1931);
and U2429 (N_2429,In_558,In_1642);
xor U2430 (N_2430,In_1664,In_47);
xnor U2431 (N_2431,In_314,In_139);
or U2432 (N_2432,In_319,In_1445);
xor U2433 (N_2433,In_384,In_284);
nand U2434 (N_2434,In_246,In_672);
nor U2435 (N_2435,In_1678,In_1098);
and U2436 (N_2436,In_1888,In_1846);
xor U2437 (N_2437,In_1189,In_100);
nand U2438 (N_2438,In_632,In_1378);
xor U2439 (N_2439,In_763,In_828);
nor U2440 (N_2440,In_1240,In_1590);
and U2441 (N_2441,In_1625,In_214);
or U2442 (N_2442,In_1916,In_1638);
nor U2443 (N_2443,In_968,In_1585);
nand U2444 (N_2444,In_1061,In_1974);
nand U2445 (N_2445,In_1229,In_649);
and U2446 (N_2446,In_1917,In_1835);
xor U2447 (N_2447,In_401,In_1214);
nand U2448 (N_2448,In_164,In_342);
nand U2449 (N_2449,In_770,In_67);
or U2450 (N_2450,In_409,In_1850);
and U2451 (N_2451,In_843,In_1857);
and U2452 (N_2452,In_1508,In_1997);
xnor U2453 (N_2453,In_1672,In_1581);
xnor U2454 (N_2454,In_1607,In_1224);
or U2455 (N_2455,In_1442,In_883);
and U2456 (N_2456,In_759,In_1912);
nor U2457 (N_2457,In_117,In_1798);
and U2458 (N_2458,In_709,In_626);
or U2459 (N_2459,In_1938,In_1293);
and U2460 (N_2460,In_856,In_1338);
and U2461 (N_2461,In_724,In_569);
xnor U2462 (N_2462,In_1734,In_506);
or U2463 (N_2463,In_14,In_1140);
nor U2464 (N_2464,In_969,In_1858);
and U2465 (N_2465,In_1263,In_200);
nor U2466 (N_2466,In_662,In_1697);
and U2467 (N_2467,In_1663,In_400);
and U2468 (N_2468,In_524,In_1390);
or U2469 (N_2469,In_1104,In_1730);
or U2470 (N_2470,In_581,In_344);
and U2471 (N_2471,In_621,In_344);
nor U2472 (N_2472,In_1557,In_1626);
xnor U2473 (N_2473,In_1828,In_602);
or U2474 (N_2474,In_1389,In_1505);
nor U2475 (N_2475,In_1183,In_1397);
nand U2476 (N_2476,In_274,In_972);
or U2477 (N_2477,In_1758,In_1042);
or U2478 (N_2478,In_493,In_1104);
nor U2479 (N_2479,In_1088,In_1778);
nand U2480 (N_2480,In_1029,In_1834);
nand U2481 (N_2481,In_983,In_262);
xnor U2482 (N_2482,In_1919,In_1256);
nor U2483 (N_2483,In_533,In_798);
or U2484 (N_2484,In_1965,In_1339);
nand U2485 (N_2485,In_746,In_1626);
and U2486 (N_2486,In_919,In_1);
nand U2487 (N_2487,In_281,In_279);
nor U2488 (N_2488,In_1259,In_1144);
xor U2489 (N_2489,In_176,In_1043);
xnor U2490 (N_2490,In_1875,In_447);
xnor U2491 (N_2491,In_66,In_501);
xnor U2492 (N_2492,In_1510,In_60);
nor U2493 (N_2493,In_436,In_13);
nor U2494 (N_2494,In_1322,In_1515);
nand U2495 (N_2495,In_1084,In_192);
xor U2496 (N_2496,In_526,In_377);
nand U2497 (N_2497,In_261,In_951);
nand U2498 (N_2498,In_1297,In_1655);
xor U2499 (N_2499,In_1067,In_401);
xor U2500 (N_2500,In_953,In_1192);
or U2501 (N_2501,In_1404,In_1874);
and U2502 (N_2502,In_473,In_867);
xor U2503 (N_2503,In_359,In_1434);
nor U2504 (N_2504,In_403,In_799);
xor U2505 (N_2505,In_1223,In_332);
or U2506 (N_2506,In_1512,In_479);
or U2507 (N_2507,In_1211,In_311);
nand U2508 (N_2508,In_1947,In_552);
nand U2509 (N_2509,In_1723,In_1811);
nor U2510 (N_2510,In_1384,In_341);
nand U2511 (N_2511,In_808,In_1100);
and U2512 (N_2512,In_646,In_531);
nor U2513 (N_2513,In_1400,In_201);
nand U2514 (N_2514,In_1286,In_1157);
nor U2515 (N_2515,In_1308,In_586);
nor U2516 (N_2516,In_32,In_843);
and U2517 (N_2517,In_1263,In_2);
or U2518 (N_2518,In_1815,In_193);
nand U2519 (N_2519,In_351,In_1204);
nor U2520 (N_2520,In_977,In_1681);
xor U2521 (N_2521,In_195,In_1876);
nand U2522 (N_2522,In_1304,In_1030);
nand U2523 (N_2523,In_690,In_573);
nor U2524 (N_2524,In_1956,In_1015);
nor U2525 (N_2525,In_995,In_818);
and U2526 (N_2526,In_1835,In_1336);
or U2527 (N_2527,In_993,In_725);
nand U2528 (N_2528,In_807,In_829);
and U2529 (N_2529,In_159,In_1055);
and U2530 (N_2530,In_1728,In_1867);
nand U2531 (N_2531,In_278,In_408);
nand U2532 (N_2532,In_1993,In_407);
or U2533 (N_2533,In_145,In_1783);
nor U2534 (N_2534,In_1935,In_841);
nand U2535 (N_2535,In_612,In_774);
or U2536 (N_2536,In_224,In_1529);
nand U2537 (N_2537,In_1242,In_466);
nor U2538 (N_2538,In_1224,In_678);
or U2539 (N_2539,In_1067,In_453);
or U2540 (N_2540,In_190,In_753);
or U2541 (N_2541,In_1494,In_90);
nand U2542 (N_2542,In_463,In_885);
nand U2543 (N_2543,In_385,In_119);
nor U2544 (N_2544,In_875,In_1687);
nor U2545 (N_2545,In_1436,In_192);
nand U2546 (N_2546,In_983,In_846);
nor U2547 (N_2547,In_1228,In_736);
xor U2548 (N_2548,In_1757,In_494);
and U2549 (N_2549,In_1513,In_1012);
or U2550 (N_2550,In_1691,In_1460);
nor U2551 (N_2551,In_383,In_430);
or U2552 (N_2552,In_1514,In_1114);
or U2553 (N_2553,In_714,In_1386);
nand U2554 (N_2554,In_155,In_1742);
and U2555 (N_2555,In_78,In_1017);
nor U2556 (N_2556,In_1619,In_489);
xor U2557 (N_2557,In_804,In_791);
nor U2558 (N_2558,In_1075,In_410);
nor U2559 (N_2559,In_1165,In_1220);
nand U2560 (N_2560,In_333,In_268);
nand U2561 (N_2561,In_1689,In_73);
or U2562 (N_2562,In_1327,In_1654);
and U2563 (N_2563,In_674,In_1391);
and U2564 (N_2564,In_417,In_1143);
xnor U2565 (N_2565,In_1805,In_636);
xor U2566 (N_2566,In_816,In_849);
and U2567 (N_2567,In_796,In_405);
nand U2568 (N_2568,In_291,In_88);
xor U2569 (N_2569,In_899,In_1944);
nor U2570 (N_2570,In_1117,In_767);
nor U2571 (N_2571,In_113,In_196);
nand U2572 (N_2572,In_87,In_1640);
xor U2573 (N_2573,In_257,In_484);
xor U2574 (N_2574,In_1354,In_1347);
and U2575 (N_2575,In_319,In_351);
nor U2576 (N_2576,In_1392,In_1022);
nand U2577 (N_2577,In_1370,In_378);
nand U2578 (N_2578,In_1224,In_419);
and U2579 (N_2579,In_1808,In_1954);
or U2580 (N_2580,In_466,In_1301);
or U2581 (N_2581,In_1566,In_1813);
nor U2582 (N_2582,In_1937,In_1417);
and U2583 (N_2583,In_322,In_1705);
and U2584 (N_2584,In_827,In_312);
xnor U2585 (N_2585,In_949,In_1529);
and U2586 (N_2586,In_210,In_832);
xnor U2587 (N_2587,In_477,In_1554);
nand U2588 (N_2588,In_185,In_482);
and U2589 (N_2589,In_457,In_498);
and U2590 (N_2590,In_747,In_1201);
or U2591 (N_2591,In_314,In_787);
nor U2592 (N_2592,In_7,In_692);
xor U2593 (N_2593,In_1871,In_866);
and U2594 (N_2594,In_779,In_277);
nand U2595 (N_2595,In_1169,In_1671);
nand U2596 (N_2596,In_1881,In_524);
nand U2597 (N_2597,In_1048,In_1772);
or U2598 (N_2598,In_1128,In_593);
xnor U2599 (N_2599,In_1577,In_1934);
nor U2600 (N_2600,In_912,In_1942);
and U2601 (N_2601,In_1261,In_125);
xnor U2602 (N_2602,In_240,In_371);
nor U2603 (N_2603,In_336,In_1131);
or U2604 (N_2604,In_644,In_1194);
nor U2605 (N_2605,In_647,In_1340);
nand U2606 (N_2606,In_1425,In_348);
nor U2607 (N_2607,In_1566,In_246);
nand U2608 (N_2608,In_991,In_1895);
xnor U2609 (N_2609,In_1266,In_539);
nand U2610 (N_2610,In_336,In_1129);
or U2611 (N_2611,In_1760,In_265);
and U2612 (N_2612,In_621,In_1091);
nand U2613 (N_2613,In_11,In_406);
xor U2614 (N_2614,In_78,In_1864);
or U2615 (N_2615,In_1677,In_636);
nand U2616 (N_2616,In_30,In_346);
and U2617 (N_2617,In_1214,In_1085);
and U2618 (N_2618,In_1237,In_1183);
nand U2619 (N_2619,In_1992,In_1231);
or U2620 (N_2620,In_637,In_548);
or U2621 (N_2621,In_1819,In_4);
xnor U2622 (N_2622,In_1209,In_426);
and U2623 (N_2623,In_81,In_1426);
nand U2624 (N_2624,In_1921,In_1833);
xor U2625 (N_2625,In_1624,In_105);
nor U2626 (N_2626,In_1520,In_1557);
xor U2627 (N_2627,In_1889,In_899);
nand U2628 (N_2628,In_438,In_179);
xnor U2629 (N_2629,In_1307,In_1057);
nand U2630 (N_2630,In_1356,In_1485);
nand U2631 (N_2631,In_827,In_568);
nand U2632 (N_2632,In_587,In_1298);
nand U2633 (N_2633,In_571,In_875);
or U2634 (N_2634,In_774,In_259);
or U2635 (N_2635,In_739,In_1249);
nand U2636 (N_2636,In_1039,In_26);
xnor U2637 (N_2637,In_690,In_1454);
and U2638 (N_2638,In_1588,In_1964);
nand U2639 (N_2639,In_211,In_808);
nand U2640 (N_2640,In_1749,In_1402);
xor U2641 (N_2641,In_177,In_628);
or U2642 (N_2642,In_545,In_1812);
nor U2643 (N_2643,In_1806,In_737);
and U2644 (N_2644,In_1804,In_1037);
and U2645 (N_2645,In_1818,In_589);
and U2646 (N_2646,In_759,In_1962);
nor U2647 (N_2647,In_349,In_217);
xor U2648 (N_2648,In_1425,In_1662);
and U2649 (N_2649,In_807,In_993);
nand U2650 (N_2650,In_547,In_1676);
xor U2651 (N_2651,In_965,In_640);
nand U2652 (N_2652,In_42,In_176);
xor U2653 (N_2653,In_1651,In_1566);
or U2654 (N_2654,In_1326,In_80);
and U2655 (N_2655,In_1911,In_243);
and U2656 (N_2656,In_1113,In_62);
nor U2657 (N_2657,In_1310,In_1356);
nor U2658 (N_2658,In_1378,In_1308);
xor U2659 (N_2659,In_1856,In_344);
xnor U2660 (N_2660,In_415,In_1982);
nand U2661 (N_2661,In_1047,In_1605);
nand U2662 (N_2662,In_355,In_1717);
or U2663 (N_2663,In_1494,In_1808);
and U2664 (N_2664,In_1555,In_1840);
nor U2665 (N_2665,In_192,In_404);
nand U2666 (N_2666,In_153,In_1725);
and U2667 (N_2667,In_1041,In_422);
and U2668 (N_2668,In_1698,In_453);
xor U2669 (N_2669,In_775,In_1773);
and U2670 (N_2670,In_1442,In_1153);
nor U2671 (N_2671,In_258,In_1084);
xnor U2672 (N_2672,In_230,In_1528);
xnor U2673 (N_2673,In_768,In_1703);
nor U2674 (N_2674,In_75,In_1804);
or U2675 (N_2675,In_948,In_1198);
or U2676 (N_2676,In_1596,In_1674);
nand U2677 (N_2677,In_1710,In_869);
xor U2678 (N_2678,In_287,In_760);
and U2679 (N_2679,In_424,In_642);
nand U2680 (N_2680,In_1015,In_113);
or U2681 (N_2681,In_1746,In_1561);
and U2682 (N_2682,In_1817,In_15);
nand U2683 (N_2683,In_1103,In_1327);
and U2684 (N_2684,In_623,In_1729);
or U2685 (N_2685,In_1307,In_438);
nand U2686 (N_2686,In_968,In_1835);
xor U2687 (N_2687,In_383,In_550);
nand U2688 (N_2688,In_1194,In_1971);
nand U2689 (N_2689,In_549,In_154);
nor U2690 (N_2690,In_1104,In_1276);
nor U2691 (N_2691,In_544,In_751);
nand U2692 (N_2692,In_522,In_1919);
xnor U2693 (N_2693,In_1985,In_1909);
nand U2694 (N_2694,In_1010,In_1090);
nor U2695 (N_2695,In_731,In_740);
xor U2696 (N_2696,In_984,In_1368);
and U2697 (N_2697,In_137,In_1913);
and U2698 (N_2698,In_1570,In_1174);
xnor U2699 (N_2699,In_719,In_1019);
nand U2700 (N_2700,In_1581,In_1636);
or U2701 (N_2701,In_258,In_393);
nand U2702 (N_2702,In_892,In_306);
or U2703 (N_2703,In_1250,In_1760);
and U2704 (N_2704,In_671,In_262);
nor U2705 (N_2705,In_647,In_183);
xnor U2706 (N_2706,In_906,In_1596);
and U2707 (N_2707,In_1049,In_373);
and U2708 (N_2708,In_984,In_1767);
xnor U2709 (N_2709,In_996,In_1266);
nand U2710 (N_2710,In_1968,In_967);
nor U2711 (N_2711,In_984,In_65);
nand U2712 (N_2712,In_1366,In_637);
nand U2713 (N_2713,In_1289,In_466);
nor U2714 (N_2714,In_566,In_1421);
or U2715 (N_2715,In_650,In_815);
xnor U2716 (N_2716,In_254,In_1225);
nand U2717 (N_2717,In_1275,In_1825);
and U2718 (N_2718,In_284,In_948);
xor U2719 (N_2719,In_338,In_896);
and U2720 (N_2720,In_1104,In_1709);
xor U2721 (N_2721,In_527,In_1814);
or U2722 (N_2722,In_984,In_1693);
and U2723 (N_2723,In_1300,In_741);
xor U2724 (N_2724,In_1917,In_399);
nor U2725 (N_2725,In_1352,In_1489);
and U2726 (N_2726,In_1082,In_1149);
nand U2727 (N_2727,In_378,In_1702);
or U2728 (N_2728,In_155,In_105);
nand U2729 (N_2729,In_1750,In_1385);
xnor U2730 (N_2730,In_1103,In_69);
nand U2731 (N_2731,In_1755,In_920);
or U2732 (N_2732,In_160,In_904);
or U2733 (N_2733,In_119,In_1226);
xnor U2734 (N_2734,In_68,In_10);
nor U2735 (N_2735,In_347,In_1576);
and U2736 (N_2736,In_1562,In_1938);
nor U2737 (N_2737,In_1718,In_1955);
xor U2738 (N_2738,In_1751,In_742);
xnor U2739 (N_2739,In_20,In_1236);
xor U2740 (N_2740,In_208,In_943);
and U2741 (N_2741,In_770,In_22);
xnor U2742 (N_2742,In_710,In_1252);
nor U2743 (N_2743,In_1471,In_767);
or U2744 (N_2744,In_284,In_914);
and U2745 (N_2745,In_1966,In_179);
xor U2746 (N_2746,In_737,In_110);
or U2747 (N_2747,In_119,In_452);
xor U2748 (N_2748,In_276,In_1456);
nor U2749 (N_2749,In_158,In_1003);
and U2750 (N_2750,In_555,In_1240);
nor U2751 (N_2751,In_1655,In_1904);
and U2752 (N_2752,In_1583,In_247);
and U2753 (N_2753,In_249,In_1764);
nor U2754 (N_2754,In_1562,In_1224);
xnor U2755 (N_2755,In_209,In_1760);
and U2756 (N_2756,In_1323,In_530);
or U2757 (N_2757,In_753,In_1031);
xnor U2758 (N_2758,In_69,In_1384);
xnor U2759 (N_2759,In_439,In_820);
nand U2760 (N_2760,In_1932,In_928);
nor U2761 (N_2761,In_395,In_235);
nand U2762 (N_2762,In_588,In_1177);
or U2763 (N_2763,In_1384,In_1509);
nor U2764 (N_2764,In_1677,In_915);
nand U2765 (N_2765,In_293,In_3);
and U2766 (N_2766,In_1964,In_720);
xor U2767 (N_2767,In_742,In_874);
nand U2768 (N_2768,In_1221,In_1515);
nor U2769 (N_2769,In_1304,In_1803);
and U2770 (N_2770,In_938,In_1509);
or U2771 (N_2771,In_1619,In_1944);
and U2772 (N_2772,In_1802,In_462);
xnor U2773 (N_2773,In_1402,In_551);
or U2774 (N_2774,In_393,In_1338);
nand U2775 (N_2775,In_866,In_1398);
xor U2776 (N_2776,In_20,In_788);
nand U2777 (N_2777,In_1369,In_178);
xor U2778 (N_2778,In_1724,In_1559);
nand U2779 (N_2779,In_980,In_1609);
or U2780 (N_2780,In_1254,In_1839);
nand U2781 (N_2781,In_1295,In_1476);
xor U2782 (N_2782,In_1314,In_436);
xor U2783 (N_2783,In_532,In_1072);
nand U2784 (N_2784,In_305,In_268);
or U2785 (N_2785,In_1237,In_1484);
xor U2786 (N_2786,In_1351,In_651);
and U2787 (N_2787,In_1313,In_1728);
or U2788 (N_2788,In_1524,In_1767);
or U2789 (N_2789,In_1268,In_1444);
xor U2790 (N_2790,In_316,In_1479);
or U2791 (N_2791,In_1043,In_401);
and U2792 (N_2792,In_796,In_468);
nor U2793 (N_2793,In_1983,In_1297);
xnor U2794 (N_2794,In_1002,In_916);
xnor U2795 (N_2795,In_836,In_1084);
nor U2796 (N_2796,In_1814,In_349);
and U2797 (N_2797,In_197,In_938);
and U2798 (N_2798,In_374,In_1966);
nand U2799 (N_2799,In_90,In_826);
nand U2800 (N_2800,In_179,In_1165);
xnor U2801 (N_2801,In_627,In_1849);
xnor U2802 (N_2802,In_48,In_1434);
or U2803 (N_2803,In_435,In_1417);
xor U2804 (N_2804,In_1565,In_1390);
nor U2805 (N_2805,In_1122,In_728);
xor U2806 (N_2806,In_21,In_569);
nor U2807 (N_2807,In_1313,In_920);
and U2808 (N_2808,In_484,In_1813);
nand U2809 (N_2809,In_783,In_1136);
or U2810 (N_2810,In_1993,In_295);
or U2811 (N_2811,In_908,In_210);
xnor U2812 (N_2812,In_1216,In_578);
and U2813 (N_2813,In_976,In_1276);
xor U2814 (N_2814,In_1629,In_1791);
xnor U2815 (N_2815,In_1391,In_1088);
xor U2816 (N_2816,In_572,In_1959);
and U2817 (N_2817,In_1252,In_1113);
or U2818 (N_2818,In_1084,In_1872);
nor U2819 (N_2819,In_679,In_1190);
nand U2820 (N_2820,In_1414,In_1329);
nand U2821 (N_2821,In_607,In_146);
xor U2822 (N_2822,In_1763,In_900);
and U2823 (N_2823,In_1004,In_941);
nor U2824 (N_2824,In_1638,In_1381);
xor U2825 (N_2825,In_894,In_1383);
or U2826 (N_2826,In_1104,In_843);
and U2827 (N_2827,In_1920,In_1932);
nor U2828 (N_2828,In_802,In_1648);
nor U2829 (N_2829,In_321,In_989);
nand U2830 (N_2830,In_1679,In_463);
nand U2831 (N_2831,In_56,In_992);
and U2832 (N_2832,In_909,In_1745);
and U2833 (N_2833,In_1664,In_1022);
xnor U2834 (N_2834,In_1582,In_1064);
or U2835 (N_2835,In_1396,In_860);
nand U2836 (N_2836,In_1900,In_617);
nand U2837 (N_2837,In_1157,In_1894);
xnor U2838 (N_2838,In_1807,In_1724);
nand U2839 (N_2839,In_1215,In_688);
and U2840 (N_2840,In_815,In_1817);
xor U2841 (N_2841,In_1383,In_231);
xor U2842 (N_2842,In_1193,In_966);
or U2843 (N_2843,In_1432,In_470);
and U2844 (N_2844,In_1821,In_964);
nor U2845 (N_2845,In_496,In_1171);
xnor U2846 (N_2846,In_1429,In_1977);
xor U2847 (N_2847,In_828,In_84);
nor U2848 (N_2848,In_564,In_1223);
xnor U2849 (N_2849,In_42,In_549);
or U2850 (N_2850,In_1767,In_1589);
nor U2851 (N_2851,In_801,In_1462);
or U2852 (N_2852,In_136,In_1739);
nand U2853 (N_2853,In_1507,In_244);
nor U2854 (N_2854,In_1588,In_357);
xnor U2855 (N_2855,In_643,In_1393);
nand U2856 (N_2856,In_1660,In_558);
nand U2857 (N_2857,In_503,In_869);
nor U2858 (N_2858,In_1993,In_1698);
and U2859 (N_2859,In_1268,In_1971);
nor U2860 (N_2860,In_774,In_533);
or U2861 (N_2861,In_1835,In_1420);
nand U2862 (N_2862,In_1389,In_170);
nand U2863 (N_2863,In_320,In_308);
or U2864 (N_2864,In_911,In_513);
nor U2865 (N_2865,In_1045,In_1690);
nor U2866 (N_2866,In_1939,In_271);
nor U2867 (N_2867,In_1854,In_1631);
and U2868 (N_2868,In_1626,In_567);
nand U2869 (N_2869,In_1620,In_1995);
and U2870 (N_2870,In_1275,In_578);
nor U2871 (N_2871,In_1515,In_1727);
and U2872 (N_2872,In_1452,In_544);
nand U2873 (N_2873,In_692,In_1946);
or U2874 (N_2874,In_898,In_59);
nor U2875 (N_2875,In_1873,In_1064);
xnor U2876 (N_2876,In_125,In_1420);
or U2877 (N_2877,In_196,In_1555);
nor U2878 (N_2878,In_1239,In_785);
or U2879 (N_2879,In_1660,In_378);
or U2880 (N_2880,In_1884,In_1806);
or U2881 (N_2881,In_899,In_1916);
or U2882 (N_2882,In_620,In_1853);
and U2883 (N_2883,In_626,In_304);
or U2884 (N_2884,In_34,In_148);
or U2885 (N_2885,In_1733,In_361);
nor U2886 (N_2886,In_104,In_231);
and U2887 (N_2887,In_825,In_1813);
xor U2888 (N_2888,In_399,In_432);
xor U2889 (N_2889,In_1995,In_191);
nor U2890 (N_2890,In_558,In_1530);
xnor U2891 (N_2891,In_893,In_642);
xnor U2892 (N_2892,In_1223,In_527);
xor U2893 (N_2893,In_1712,In_1229);
or U2894 (N_2894,In_1237,In_1449);
nand U2895 (N_2895,In_72,In_80);
nor U2896 (N_2896,In_1474,In_1306);
nand U2897 (N_2897,In_1980,In_1872);
and U2898 (N_2898,In_1761,In_1534);
xor U2899 (N_2899,In_1320,In_1121);
nand U2900 (N_2900,In_382,In_492);
and U2901 (N_2901,In_742,In_1523);
and U2902 (N_2902,In_1579,In_691);
and U2903 (N_2903,In_988,In_155);
nand U2904 (N_2904,In_1619,In_1939);
nor U2905 (N_2905,In_1341,In_1461);
and U2906 (N_2906,In_1184,In_1712);
nor U2907 (N_2907,In_529,In_600);
or U2908 (N_2908,In_142,In_811);
or U2909 (N_2909,In_1360,In_862);
nand U2910 (N_2910,In_1931,In_1292);
xnor U2911 (N_2911,In_118,In_142);
or U2912 (N_2912,In_114,In_940);
nand U2913 (N_2913,In_661,In_12);
nor U2914 (N_2914,In_699,In_1821);
and U2915 (N_2915,In_422,In_1339);
nor U2916 (N_2916,In_1583,In_722);
and U2917 (N_2917,In_1107,In_778);
and U2918 (N_2918,In_1507,In_1828);
and U2919 (N_2919,In_644,In_1269);
or U2920 (N_2920,In_1837,In_1067);
nand U2921 (N_2921,In_1874,In_27);
nand U2922 (N_2922,In_86,In_1064);
nor U2923 (N_2923,In_1174,In_1423);
nand U2924 (N_2924,In_1031,In_423);
nor U2925 (N_2925,In_1409,In_1571);
or U2926 (N_2926,In_615,In_328);
or U2927 (N_2927,In_948,In_1539);
nor U2928 (N_2928,In_1365,In_1198);
and U2929 (N_2929,In_592,In_586);
nand U2930 (N_2930,In_773,In_1695);
nor U2931 (N_2931,In_909,In_1643);
nand U2932 (N_2932,In_122,In_447);
nand U2933 (N_2933,In_789,In_824);
xnor U2934 (N_2934,In_1020,In_132);
and U2935 (N_2935,In_1536,In_108);
and U2936 (N_2936,In_1426,In_1187);
xnor U2937 (N_2937,In_1244,In_1798);
nand U2938 (N_2938,In_993,In_1354);
nor U2939 (N_2939,In_1833,In_257);
nand U2940 (N_2940,In_698,In_1637);
xnor U2941 (N_2941,In_1130,In_174);
nor U2942 (N_2942,In_201,In_419);
and U2943 (N_2943,In_364,In_1927);
nand U2944 (N_2944,In_639,In_1526);
nor U2945 (N_2945,In_872,In_547);
nor U2946 (N_2946,In_98,In_242);
nand U2947 (N_2947,In_954,In_1563);
xnor U2948 (N_2948,In_1289,In_1653);
or U2949 (N_2949,In_308,In_811);
or U2950 (N_2950,In_927,In_966);
xnor U2951 (N_2951,In_1215,In_1378);
and U2952 (N_2952,In_400,In_698);
nor U2953 (N_2953,In_961,In_400);
and U2954 (N_2954,In_68,In_742);
and U2955 (N_2955,In_563,In_666);
nand U2956 (N_2956,In_9,In_591);
xnor U2957 (N_2957,In_1983,In_556);
or U2958 (N_2958,In_1172,In_1232);
nand U2959 (N_2959,In_60,In_373);
nand U2960 (N_2960,In_427,In_533);
nand U2961 (N_2961,In_155,In_836);
nand U2962 (N_2962,In_304,In_859);
or U2963 (N_2963,In_430,In_227);
or U2964 (N_2964,In_284,In_225);
xnor U2965 (N_2965,In_1916,In_1304);
xnor U2966 (N_2966,In_1438,In_425);
nand U2967 (N_2967,In_1049,In_1830);
and U2968 (N_2968,In_294,In_1666);
nor U2969 (N_2969,In_295,In_332);
and U2970 (N_2970,In_162,In_958);
xor U2971 (N_2971,In_1946,In_705);
xor U2972 (N_2972,In_971,In_1906);
or U2973 (N_2973,In_1631,In_553);
xor U2974 (N_2974,In_1743,In_1867);
nand U2975 (N_2975,In_1229,In_1577);
and U2976 (N_2976,In_1332,In_59);
nor U2977 (N_2977,In_1587,In_161);
nand U2978 (N_2978,In_221,In_1871);
nand U2979 (N_2979,In_970,In_1413);
nand U2980 (N_2980,In_986,In_968);
and U2981 (N_2981,In_1766,In_1200);
nand U2982 (N_2982,In_650,In_599);
or U2983 (N_2983,In_418,In_515);
or U2984 (N_2984,In_943,In_261);
nand U2985 (N_2985,In_1547,In_1938);
and U2986 (N_2986,In_1,In_689);
xor U2987 (N_2987,In_1848,In_1019);
and U2988 (N_2988,In_1487,In_443);
xnor U2989 (N_2989,In_1953,In_896);
xnor U2990 (N_2990,In_5,In_419);
nand U2991 (N_2991,In_1616,In_1402);
xor U2992 (N_2992,In_826,In_783);
nand U2993 (N_2993,In_1677,In_811);
or U2994 (N_2994,In_550,In_1527);
xnor U2995 (N_2995,In_1767,In_114);
and U2996 (N_2996,In_686,In_1144);
nand U2997 (N_2997,In_838,In_1638);
xnor U2998 (N_2998,In_1951,In_392);
xor U2999 (N_2999,In_87,In_1319);
or U3000 (N_3000,In_1553,In_633);
xnor U3001 (N_3001,In_1044,In_160);
xnor U3002 (N_3002,In_1936,In_188);
xnor U3003 (N_3003,In_315,In_1629);
or U3004 (N_3004,In_356,In_397);
nand U3005 (N_3005,In_1905,In_914);
xnor U3006 (N_3006,In_610,In_442);
or U3007 (N_3007,In_1313,In_154);
or U3008 (N_3008,In_1283,In_1166);
or U3009 (N_3009,In_1136,In_1108);
nand U3010 (N_3010,In_1310,In_279);
nor U3011 (N_3011,In_1308,In_543);
or U3012 (N_3012,In_355,In_220);
or U3013 (N_3013,In_701,In_1872);
or U3014 (N_3014,In_1978,In_1774);
nand U3015 (N_3015,In_1872,In_479);
nand U3016 (N_3016,In_131,In_1414);
or U3017 (N_3017,In_266,In_1605);
nor U3018 (N_3018,In_908,In_1945);
and U3019 (N_3019,In_1499,In_138);
or U3020 (N_3020,In_1785,In_1920);
or U3021 (N_3021,In_240,In_1492);
nor U3022 (N_3022,In_1739,In_420);
nand U3023 (N_3023,In_547,In_1594);
and U3024 (N_3024,In_877,In_1679);
nor U3025 (N_3025,In_976,In_406);
xnor U3026 (N_3026,In_548,In_314);
and U3027 (N_3027,In_875,In_47);
and U3028 (N_3028,In_736,In_1633);
or U3029 (N_3029,In_304,In_1936);
or U3030 (N_3030,In_1980,In_635);
or U3031 (N_3031,In_701,In_1158);
or U3032 (N_3032,In_302,In_1547);
nor U3033 (N_3033,In_1352,In_226);
nand U3034 (N_3034,In_517,In_1801);
nor U3035 (N_3035,In_1280,In_1539);
xnor U3036 (N_3036,In_1985,In_1139);
nand U3037 (N_3037,In_1896,In_333);
nand U3038 (N_3038,In_380,In_5);
and U3039 (N_3039,In_551,In_17);
and U3040 (N_3040,In_855,In_580);
or U3041 (N_3041,In_1526,In_1969);
and U3042 (N_3042,In_66,In_624);
xnor U3043 (N_3043,In_1299,In_222);
xor U3044 (N_3044,In_1512,In_120);
xnor U3045 (N_3045,In_1652,In_643);
nor U3046 (N_3046,In_30,In_1165);
and U3047 (N_3047,In_477,In_1531);
nand U3048 (N_3048,In_1245,In_1169);
or U3049 (N_3049,In_708,In_365);
xor U3050 (N_3050,In_1730,In_998);
nand U3051 (N_3051,In_1887,In_1958);
and U3052 (N_3052,In_113,In_535);
or U3053 (N_3053,In_942,In_1926);
xnor U3054 (N_3054,In_1815,In_461);
nor U3055 (N_3055,In_1971,In_1196);
and U3056 (N_3056,In_1931,In_1535);
nand U3057 (N_3057,In_251,In_596);
nor U3058 (N_3058,In_644,In_531);
xor U3059 (N_3059,In_819,In_1011);
and U3060 (N_3060,In_1325,In_680);
and U3061 (N_3061,In_1475,In_219);
and U3062 (N_3062,In_1807,In_1283);
nand U3063 (N_3063,In_1391,In_343);
xnor U3064 (N_3064,In_1439,In_9);
nand U3065 (N_3065,In_1123,In_837);
xnor U3066 (N_3066,In_128,In_1680);
or U3067 (N_3067,In_1896,In_1910);
nand U3068 (N_3068,In_1580,In_560);
and U3069 (N_3069,In_427,In_239);
nand U3070 (N_3070,In_1122,In_1029);
xnor U3071 (N_3071,In_1957,In_533);
nand U3072 (N_3072,In_1127,In_1392);
nor U3073 (N_3073,In_1425,In_1915);
or U3074 (N_3074,In_1348,In_835);
or U3075 (N_3075,In_30,In_242);
nor U3076 (N_3076,In_28,In_1456);
or U3077 (N_3077,In_277,In_494);
nor U3078 (N_3078,In_1527,In_1002);
and U3079 (N_3079,In_1469,In_1459);
or U3080 (N_3080,In_1157,In_831);
nor U3081 (N_3081,In_257,In_344);
nor U3082 (N_3082,In_1921,In_1390);
xnor U3083 (N_3083,In_1238,In_939);
nand U3084 (N_3084,In_1008,In_1783);
xor U3085 (N_3085,In_90,In_1361);
or U3086 (N_3086,In_451,In_172);
nand U3087 (N_3087,In_1952,In_549);
and U3088 (N_3088,In_1406,In_1544);
nor U3089 (N_3089,In_840,In_1558);
and U3090 (N_3090,In_111,In_445);
or U3091 (N_3091,In_231,In_418);
or U3092 (N_3092,In_1186,In_412);
and U3093 (N_3093,In_847,In_1039);
and U3094 (N_3094,In_1470,In_1362);
nor U3095 (N_3095,In_770,In_257);
and U3096 (N_3096,In_1075,In_1829);
or U3097 (N_3097,In_1174,In_671);
xnor U3098 (N_3098,In_1696,In_7);
and U3099 (N_3099,In_1435,In_279);
or U3100 (N_3100,In_327,In_1911);
nor U3101 (N_3101,In_326,In_1885);
nor U3102 (N_3102,In_951,In_657);
or U3103 (N_3103,In_251,In_337);
and U3104 (N_3104,In_1039,In_543);
xor U3105 (N_3105,In_363,In_951);
or U3106 (N_3106,In_1126,In_1372);
xor U3107 (N_3107,In_1455,In_1694);
xor U3108 (N_3108,In_1274,In_154);
nor U3109 (N_3109,In_526,In_505);
nand U3110 (N_3110,In_1629,In_218);
or U3111 (N_3111,In_110,In_265);
xor U3112 (N_3112,In_1045,In_322);
or U3113 (N_3113,In_1099,In_1355);
nand U3114 (N_3114,In_602,In_555);
and U3115 (N_3115,In_770,In_1467);
xor U3116 (N_3116,In_1706,In_1417);
xor U3117 (N_3117,In_482,In_1555);
nor U3118 (N_3118,In_1284,In_234);
nand U3119 (N_3119,In_1729,In_106);
nand U3120 (N_3120,In_506,In_120);
nor U3121 (N_3121,In_1114,In_720);
or U3122 (N_3122,In_755,In_1445);
nor U3123 (N_3123,In_1446,In_756);
nand U3124 (N_3124,In_1574,In_1316);
nand U3125 (N_3125,In_1196,In_1672);
xor U3126 (N_3126,In_296,In_815);
or U3127 (N_3127,In_480,In_395);
and U3128 (N_3128,In_49,In_1436);
or U3129 (N_3129,In_1943,In_1247);
nor U3130 (N_3130,In_271,In_1656);
or U3131 (N_3131,In_440,In_1088);
and U3132 (N_3132,In_1895,In_1648);
nor U3133 (N_3133,In_1692,In_1977);
nand U3134 (N_3134,In_125,In_1869);
nor U3135 (N_3135,In_831,In_365);
nand U3136 (N_3136,In_1020,In_428);
and U3137 (N_3137,In_1591,In_427);
nor U3138 (N_3138,In_339,In_1223);
or U3139 (N_3139,In_1157,In_447);
or U3140 (N_3140,In_245,In_1747);
and U3141 (N_3141,In_985,In_368);
xnor U3142 (N_3142,In_151,In_13);
nor U3143 (N_3143,In_1892,In_382);
or U3144 (N_3144,In_690,In_164);
and U3145 (N_3145,In_720,In_489);
and U3146 (N_3146,In_1530,In_1856);
or U3147 (N_3147,In_1138,In_905);
nand U3148 (N_3148,In_1072,In_1431);
nand U3149 (N_3149,In_1368,In_1556);
nor U3150 (N_3150,In_491,In_1448);
or U3151 (N_3151,In_329,In_1153);
or U3152 (N_3152,In_1313,In_1717);
and U3153 (N_3153,In_1072,In_545);
xnor U3154 (N_3154,In_1245,In_21);
nand U3155 (N_3155,In_28,In_604);
and U3156 (N_3156,In_518,In_1283);
or U3157 (N_3157,In_717,In_1993);
or U3158 (N_3158,In_1305,In_470);
and U3159 (N_3159,In_1528,In_662);
and U3160 (N_3160,In_1303,In_1473);
and U3161 (N_3161,In_242,In_1103);
and U3162 (N_3162,In_838,In_1969);
xor U3163 (N_3163,In_200,In_1908);
xnor U3164 (N_3164,In_523,In_601);
xor U3165 (N_3165,In_270,In_222);
and U3166 (N_3166,In_1821,In_110);
nand U3167 (N_3167,In_228,In_1172);
nor U3168 (N_3168,In_1574,In_583);
xnor U3169 (N_3169,In_1645,In_486);
nand U3170 (N_3170,In_545,In_663);
nand U3171 (N_3171,In_79,In_1905);
xor U3172 (N_3172,In_257,In_648);
nor U3173 (N_3173,In_192,In_1158);
xnor U3174 (N_3174,In_723,In_1154);
nand U3175 (N_3175,In_1005,In_1348);
nand U3176 (N_3176,In_1887,In_255);
or U3177 (N_3177,In_1322,In_1820);
or U3178 (N_3178,In_497,In_1687);
or U3179 (N_3179,In_1238,In_251);
or U3180 (N_3180,In_868,In_1575);
nand U3181 (N_3181,In_710,In_1947);
nand U3182 (N_3182,In_1989,In_1799);
or U3183 (N_3183,In_848,In_1202);
and U3184 (N_3184,In_1598,In_1491);
or U3185 (N_3185,In_253,In_1313);
or U3186 (N_3186,In_443,In_1219);
or U3187 (N_3187,In_616,In_946);
or U3188 (N_3188,In_824,In_610);
xor U3189 (N_3189,In_109,In_1115);
or U3190 (N_3190,In_1478,In_130);
nand U3191 (N_3191,In_1236,In_921);
or U3192 (N_3192,In_256,In_503);
xnor U3193 (N_3193,In_1986,In_615);
and U3194 (N_3194,In_1446,In_1607);
nor U3195 (N_3195,In_1097,In_1323);
nand U3196 (N_3196,In_1541,In_1528);
nor U3197 (N_3197,In_1329,In_858);
and U3198 (N_3198,In_1992,In_765);
nor U3199 (N_3199,In_1261,In_851);
nor U3200 (N_3200,In_1296,In_211);
and U3201 (N_3201,In_1796,In_1462);
xnor U3202 (N_3202,In_618,In_603);
nor U3203 (N_3203,In_1101,In_891);
and U3204 (N_3204,In_786,In_1773);
xor U3205 (N_3205,In_1621,In_1907);
nand U3206 (N_3206,In_982,In_1419);
nand U3207 (N_3207,In_761,In_1929);
and U3208 (N_3208,In_1611,In_55);
nor U3209 (N_3209,In_460,In_711);
xnor U3210 (N_3210,In_810,In_1993);
nand U3211 (N_3211,In_1669,In_1859);
and U3212 (N_3212,In_904,In_137);
nand U3213 (N_3213,In_95,In_367);
nor U3214 (N_3214,In_1036,In_107);
and U3215 (N_3215,In_1229,In_1912);
nor U3216 (N_3216,In_915,In_676);
xnor U3217 (N_3217,In_400,In_1384);
nor U3218 (N_3218,In_1119,In_745);
or U3219 (N_3219,In_617,In_84);
and U3220 (N_3220,In_30,In_1854);
or U3221 (N_3221,In_1720,In_98);
and U3222 (N_3222,In_156,In_446);
or U3223 (N_3223,In_1768,In_1810);
and U3224 (N_3224,In_1910,In_1126);
nor U3225 (N_3225,In_904,In_595);
and U3226 (N_3226,In_1214,In_1221);
and U3227 (N_3227,In_1292,In_1744);
and U3228 (N_3228,In_1359,In_1954);
nor U3229 (N_3229,In_1491,In_547);
or U3230 (N_3230,In_1287,In_303);
and U3231 (N_3231,In_526,In_6);
and U3232 (N_3232,In_707,In_1178);
xor U3233 (N_3233,In_313,In_10);
nand U3234 (N_3234,In_233,In_1227);
nand U3235 (N_3235,In_329,In_1551);
nand U3236 (N_3236,In_371,In_82);
nand U3237 (N_3237,In_159,In_95);
or U3238 (N_3238,In_1045,In_373);
or U3239 (N_3239,In_1091,In_959);
xnor U3240 (N_3240,In_1805,In_678);
nand U3241 (N_3241,In_1359,In_181);
xor U3242 (N_3242,In_898,In_726);
or U3243 (N_3243,In_288,In_1608);
xor U3244 (N_3244,In_1549,In_1300);
nand U3245 (N_3245,In_75,In_925);
and U3246 (N_3246,In_153,In_1244);
or U3247 (N_3247,In_1677,In_1656);
and U3248 (N_3248,In_1085,In_1712);
and U3249 (N_3249,In_1443,In_1233);
or U3250 (N_3250,In_711,In_1406);
and U3251 (N_3251,In_1267,In_117);
nor U3252 (N_3252,In_916,In_1690);
nor U3253 (N_3253,In_545,In_1481);
nand U3254 (N_3254,In_600,In_1859);
or U3255 (N_3255,In_1150,In_965);
nand U3256 (N_3256,In_849,In_544);
nor U3257 (N_3257,In_1572,In_1796);
nand U3258 (N_3258,In_1513,In_1382);
nor U3259 (N_3259,In_1715,In_1642);
and U3260 (N_3260,In_1299,In_381);
xor U3261 (N_3261,In_370,In_883);
and U3262 (N_3262,In_1687,In_1111);
and U3263 (N_3263,In_1242,In_1727);
or U3264 (N_3264,In_79,In_1053);
xor U3265 (N_3265,In_1113,In_1620);
nor U3266 (N_3266,In_877,In_841);
nor U3267 (N_3267,In_1377,In_980);
xor U3268 (N_3268,In_1647,In_1466);
xnor U3269 (N_3269,In_945,In_1540);
and U3270 (N_3270,In_484,In_1375);
xor U3271 (N_3271,In_90,In_1590);
or U3272 (N_3272,In_962,In_667);
and U3273 (N_3273,In_465,In_1202);
xnor U3274 (N_3274,In_1185,In_1751);
and U3275 (N_3275,In_76,In_1619);
nand U3276 (N_3276,In_1730,In_628);
or U3277 (N_3277,In_939,In_1647);
nand U3278 (N_3278,In_1457,In_146);
or U3279 (N_3279,In_21,In_1392);
nor U3280 (N_3280,In_1500,In_32);
xnor U3281 (N_3281,In_1859,In_1207);
xor U3282 (N_3282,In_489,In_227);
nor U3283 (N_3283,In_1735,In_1464);
nand U3284 (N_3284,In_1196,In_573);
xor U3285 (N_3285,In_98,In_1989);
xor U3286 (N_3286,In_1671,In_1780);
xnor U3287 (N_3287,In_1554,In_1577);
nor U3288 (N_3288,In_1570,In_674);
nor U3289 (N_3289,In_109,In_1914);
xnor U3290 (N_3290,In_1986,In_1185);
nor U3291 (N_3291,In_86,In_791);
or U3292 (N_3292,In_1947,In_13);
xnor U3293 (N_3293,In_737,In_1977);
xor U3294 (N_3294,In_1023,In_1044);
and U3295 (N_3295,In_1262,In_968);
and U3296 (N_3296,In_1502,In_1270);
and U3297 (N_3297,In_1131,In_1329);
and U3298 (N_3298,In_592,In_496);
nand U3299 (N_3299,In_807,In_1620);
xnor U3300 (N_3300,In_90,In_299);
nor U3301 (N_3301,In_375,In_1433);
and U3302 (N_3302,In_896,In_328);
xnor U3303 (N_3303,In_1423,In_289);
and U3304 (N_3304,In_1595,In_336);
and U3305 (N_3305,In_273,In_415);
or U3306 (N_3306,In_50,In_546);
nand U3307 (N_3307,In_1072,In_742);
xnor U3308 (N_3308,In_369,In_23);
nand U3309 (N_3309,In_113,In_1828);
or U3310 (N_3310,In_1249,In_549);
and U3311 (N_3311,In_1391,In_1591);
nand U3312 (N_3312,In_25,In_936);
nor U3313 (N_3313,In_1972,In_1470);
and U3314 (N_3314,In_236,In_1070);
nor U3315 (N_3315,In_1340,In_835);
and U3316 (N_3316,In_1546,In_156);
nor U3317 (N_3317,In_560,In_1727);
xor U3318 (N_3318,In_1625,In_1282);
nor U3319 (N_3319,In_1322,In_1018);
xor U3320 (N_3320,In_131,In_728);
xnor U3321 (N_3321,In_162,In_1038);
and U3322 (N_3322,In_1104,In_1970);
and U3323 (N_3323,In_447,In_10);
nand U3324 (N_3324,In_489,In_19);
nand U3325 (N_3325,In_1239,In_1773);
and U3326 (N_3326,In_103,In_46);
or U3327 (N_3327,In_1203,In_192);
and U3328 (N_3328,In_454,In_1121);
xnor U3329 (N_3329,In_1045,In_425);
nand U3330 (N_3330,In_782,In_339);
nor U3331 (N_3331,In_817,In_1193);
or U3332 (N_3332,In_1784,In_1021);
xnor U3333 (N_3333,In_801,In_886);
nand U3334 (N_3334,In_1830,In_1574);
nand U3335 (N_3335,In_1892,In_431);
xor U3336 (N_3336,In_1193,In_1121);
xnor U3337 (N_3337,In_49,In_179);
xor U3338 (N_3338,In_1797,In_632);
xor U3339 (N_3339,In_899,In_711);
and U3340 (N_3340,In_1736,In_802);
nor U3341 (N_3341,In_1460,In_1393);
nor U3342 (N_3342,In_733,In_28);
xor U3343 (N_3343,In_1908,In_578);
nor U3344 (N_3344,In_842,In_506);
and U3345 (N_3345,In_275,In_425);
nor U3346 (N_3346,In_1226,In_546);
nor U3347 (N_3347,In_132,In_1197);
nand U3348 (N_3348,In_1380,In_424);
nand U3349 (N_3349,In_1676,In_414);
or U3350 (N_3350,In_1086,In_1294);
or U3351 (N_3351,In_1019,In_740);
xnor U3352 (N_3352,In_678,In_1539);
or U3353 (N_3353,In_1017,In_1374);
xnor U3354 (N_3354,In_1939,In_1044);
and U3355 (N_3355,In_1883,In_803);
nand U3356 (N_3356,In_390,In_679);
or U3357 (N_3357,In_18,In_401);
or U3358 (N_3358,In_1676,In_635);
and U3359 (N_3359,In_755,In_1444);
and U3360 (N_3360,In_1127,In_1801);
nor U3361 (N_3361,In_1729,In_1249);
and U3362 (N_3362,In_1761,In_1263);
nand U3363 (N_3363,In_1039,In_1824);
nand U3364 (N_3364,In_596,In_132);
nand U3365 (N_3365,In_1247,In_907);
or U3366 (N_3366,In_1188,In_1898);
and U3367 (N_3367,In_1358,In_979);
and U3368 (N_3368,In_1104,In_64);
nor U3369 (N_3369,In_1782,In_60);
nor U3370 (N_3370,In_1113,In_1306);
nor U3371 (N_3371,In_256,In_1866);
and U3372 (N_3372,In_499,In_161);
and U3373 (N_3373,In_1205,In_1947);
and U3374 (N_3374,In_13,In_694);
xor U3375 (N_3375,In_555,In_1570);
and U3376 (N_3376,In_356,In_1351);
and U3377 (N_3377,In_682,In_1347);
and U3378 (N_3378,In_552,In_734);
nand U3379 (N_3379,In_435,In_335);
xnor U3380 (N_3380,In_1317,In_1577);
nand U3381 (N_3381,In_419,In_1207);
nand U3382 (N_3382,In_1478,In_643);
xor U3383 (N_3383,In_1178,In_1047);
or U3384 (N_3384,In_1574,In_1061);
nor U3385 (N_3385,In_1275,In_1482);
nand U3386 (N_3386,In_1432,In_449);
xnor U3387 (N_3387,In_521,In_363);
or U3388 (N_3388,In_1871,In_513);
or U3389 (N_3389,In_893,In_1530);
nor U3390 (N_3390,In_84,In_1113);
nor U3391 (N_3391,In_232,In_1489);
xor U3392 (N_3392,In_1968,In_234);
or U3393 (N_3393,In_792,In_1545);
xnor U3394 (N_3394,In_854,In_896);
nand U3395 (N_3395,In_1715,In_1822);
or U3396 (N_3396,In_1510,In_513);
nor U3397 (N_3397,In_529,In_1244);
xor U3398 (N_3398,In_1213,In_1451);
xnor U3399 (N_3399,In_119,In_600);
nor U3400 (N_3400,In_1661,In_2);
xnor U3401 (N_3401,In_1327,In_990);
nand U3402 (N_3402,In_1358,In_7);
or U3403 (N_3403,In_883,In_657);
and U3404 (N_3404,In_1216,In_1769);
nor U3405 (N_3405,In_1537,In_935);
and U3406 (N_3406,In_988,In_1383);
nand U3407 (N_3407,In_1432,In_952);
nand U3408 (N_3408,In_377,In_108);
nor U3409 (N_3409,In_545,In_1677);
xor U3410 (N_3410,In_1273,In_650);
nand U3411 (N_3411,In_328,In_1255);
or U3412 (N_3412,In_1251,In_1869);
nand U3413 (N_3413,In_1350,In_845);
nand U3414 (N_3414,In_552,In_1510);
xor U3415 (N_3415,In_1428,In_1948);
xnor U3416 (N_3416,In_1373,In_1530);
or U3417 (N_3417,In_1901,In_281);
and U3418 (N_3418,In_389,In_1681);
and U3419 (N_3419,In_1469,In_777);
xnor U3420 (N_3420,In_1893,In_1061);
nor U3421 (N_3421,In_1998,In_1490);
nand U3422 (N_3422,In_495,In_319);
and U3423 (N_3423,In_1613,In_1683);
nand U3424 (N_3424,In_1451,In_914);
xor U3425 (N_3425,In_532,In_1744);
nand U3426 (N_3426,In_497,In_1785);
and U3427 (N_3427,In_1120,In_603);
xnor U3428 (N_3428,In_1116,In_1008);
and U3429 (N_3429,In_1135,In_1110);
nor U3430 (N_3430,In_1051,In_1491);
xor U3431 (N_3431,In_1469,In_1753);
nand U3432 (N_3432,In_1819,In_1409);
nand U3433 (N_3433,In_1254,In_1199);
nand U3434 (N_3434,In_1894,In_1890);
nor U3435 (N_3435,In_1211,In_1564);
nor U3436 (N_3436,In_1037,In_672);
or U3437 (N_3437,In_63,In_376);
nand U3438 (N_3438,In_876,In_1880);
nand U3439 (N_3439,In_323,In_173);
or U3440 (N_3440,In_573,In_1014);
xnor U3441 (N_3441,In_662,In_563);
or U3442 (N_3442,In_720,In_829);
xor U3443 (N_3443,In_979,In_584);
xnor U3444 (N_3444,In_914,In_765);
and U3445 (N_3445,In_333,In_1600);
and U3446 (N_3446,In_774,In_911);
and U3447 (N_3447,In_1425,In_954);
or U3448 (N_3448,In_279,In_1312);
and U3449 (N_3449,In_1599,In_1453);
xnor U3450 (N_3450,In_198,In_1720);
and U3451 (N_3451,In_1255,In_849);
nor U3452 (N_3452,In_1819,In_435);
and U3453 (N_3453,In_1332,In_36);
and U3454 (N_3454,In_1892,In_1623);
xor U3455 (N_3455,In_900,In_1783);
nand U3456 (N_3456,In_712,In_340);
or U3457 (N_3457,In_1813,In_1606);
nand U3458 (N_3458,In_179,In_916);
or U3459 (N_3459,In_1701,In_1732);
nor U3460 (N_3460,In_1187,In_484);
xnor U3461 (N_3461,In_1217,In_190);
and U3462 (N_3462,In_6,In_1263);
xnor U3463 (N_3463,In_922,In_886);
nor U3464 (N_3464,In_1396,In_213);
and U3465 (N_3465,In_35,In_211);
nor U3466 (N_3466,In_1433,In_441);
or U3467 (N_3467,In_1705,In_1191);
and U3468 (N_3468,In_344,In_1026);
nor U3469 (N_3469,In_1520,In_93);
nand U3470 (N_3470,In_191,In_1956);
or U3471 (N_3471,In_1,In_1745);
nand U3472 (N_3472,In_1083,In_1351);
and U3473 (N_3473,In_326,In_1950);
or U3474 (N_3474,In_1364,In_836);
or U3475 (N_3475,In_668,In_666);
nor U3476 (N_3476,In_1339,In_43);
and U3477 (N_3477,In_613,In_362);
nand U3478 (N_3478,In_1178,In_1145);
and U3479 (N_3479,In_1945,In_388);
nor U3480 (N_3480,In_893,In_514);
and U3481 (N_3481,In_1420,In_1013);
and U3482 (N_3482,In_1520,In_493);
nor U3483 (N_3483,In_1184,In_259);
nor U3484 (N_3484,In_1013,In_1584);
and U3485 (N_3485,In_1250,In_992);
or U3486 (N_3486,In_375,In_651);
or U3487 (N_3487,In_1096,In_46);
or U3488 (N_3488,In_1896,In_373);
xnor U3489 (N_3489,In_1970,In_925);
and U3490 (N_3490,In_987,In_1893);
xor U3491 (N_3491,In_360,In_693);
nand U3492 (N_3492,In_562,In_1623);
xnor U3493 (N_3493,In_1536,In_384);
xnor U3494 (N_3494,In_1554,In_1591);
xor U3495 (N_3495,In_401,In_856);
or U3496 (N_3496,In_48,In_696);
nor U3497 (N_3497,In_1497,In_850);
or U3498 (N_3498,In_1025,In_1163);
and U3499 (N_3499,In_477,In_1080);
or U3500 (N_3500,In_989,In_572);
nor U3501 (N_3501,In_1710,In_1499);
xnor U3502 (N_3502,In_848,In_1562);
or U3503 (N_3503,In_1133,In_400);
xor U3504 (N_3504,In_994,In_1394);
nand U3505 (N_3505,In_1782,In_87);
nand U3506 (N_3506,In_1869,In_1790);
and U3507 (N_3507,In_233,In_1631);
xnor U3508 (N_3508,In_1313,In_1928);
or U3509 (N_3509,In_1257,In_917);
xnor U3510 (N_3510,In_1164,In_1048);
nor U3511 (N_3511,In_945,In_363);
or U3512 (N_3512,In_208,In_251);
nor U3513 (N_3513,In_1754,In_770);
nor U3514 (N_3514,In_279,In_379);
and U3515 (N_3515,In_316,In_1430);
xnor U3516 (N_3516,In_381,In_1047);
nor U3517 (N_3517,In_1838,In_1252);
nor U3518 (N_3518,In_1915,In_223);
and U3519 (N_3519,In_1130,In_968);
xor U3520 (N_3520,In_1581,In_1158);
or U3521 (N_3521,In_691,In_1750);
nand U3522 (N_3522,In_243,In_1212);
nor U3523 (N_3523,In_1303,In_39);
nand U3524 (N_3524,In_747,In_800);
or U3525 (N_3525,In_1722,In_518);
or U3526 (N_3526,In_1195,In_1000);
nand U3527 (N_3527,In_1229,In_114);
or U3528 (N_3528,In_1045,In_647);
or U3529 (N_3529,In_600,In_790);
xnor U3530 (N_3530,In_1547,In_1062);
nor U3531 (N_3531,In_1059,In_1717);
nand U3532 (N_3532,In_1596,In_943);
or U3533 (N_3533,In_244,In_47);
xor U3534 (N_3534,In_1631,In_743);
or U3535 (N_3535,In_610,In_99);
and U3536 (N_3536,In_500,In_8);
or U3537 (N_3537,In_1678,In_229);
nor U3538 (N_3538,In_1518,In_1615);
and U3539 (N_3539,In_512,In_551);
or U3540 (N_3540,In_375,In_1402);
xnor U3541 (N_3541,In_161,In_53);
nand U3542 (N_3542,In_827,In_781);
nor U3543 (N_3543,In_263,In_1585);
nand U3544 (N_3544,In_280,In_650);
or U3545 (N_3545,In_808,In_437);
or U3546 (N_3546,In_614,In_1771);
nand U3547 (N_3547,In_522,In_1419);
or U3548 (N_3548,In_767,In_856);
xor U3549 (N_3549,In_1206,In_256);
nor U3550 (N_3550,In_1763,In_618);
nor U3551 (N_3551,In_121,In_1610);
nand U3552 (N_3552,In_1326,In_591);
and U3553 (N_3553,In_1921,In_945);
or U3554 (N_3554,In_1381,In_706);
nor U3555 (N_3555,In_1200,In_60);
xor U3556 (N_3556,In_561,In_1388);
and U3557 (N_3557,In_1588,In_1759);
xnor U3558 (N_3558,In_36,In_1802);
nand U3559 (N_3559,In_204,In_380);
and U3560 (N_3560,In_1983,In_567);
and U3561 (N_3561,In_219,In_1365);
xor U3562 (N_3562,In_768,In_76);
or U3563 (N_3563,In_280,In_700);
nand U3564 (N_3564,In_429,In_831);
or U3565 (N_3565,In_1784,In_16);
xor U3566 (N_3566,In_334,In_1100);
xnor U3567 (N_3567,In_1464,In_1975);
nor U3568 (N_3568,In_676,In_1396);
or U3569 (N_3569,In_1490,In_1767);
xnor U3570 (N_3570,In_527,In_1032);
and U3571 (N_3571,In_263,In_1717);
and U3572 (N_3572,In_645,In_1998);
nor U3573 (N_3573,In_200,In_766);
nor U3574 (N_3574,In_629,In_175);
nor U3575 (N_3575,In_1314,In_407);
and U3576 (N_3576,In_1732,In_646);
nand U3577 (N_3577,In_387,In_955);
nor U3578 (N_3578,In_1007,In_374);
or U3579 (N_3579,In_147,In_1205);
xor U3580 (N_3580,In_220,In_1335);
nor U3581 (N_3581,In_206,In_766);
nand U3582 (N_3582,In_16,In_71);
nand U3583 (N_3583,In_448,In_1106);
and U3584 (N_3584,In_1320,In_59);
xor U3585 (N_3585,In_1715,In_506);
and U3586 (N_3586,In_1891,In_560);
or U3587 (N_3587,In_1874,In_1445);
xnor U3588 (N_3588,In_1144,In_1812);
and U3589 (N_3589,In_1301,In_1894);
nor U3590 (N_3590,In_1482,In_728);
nor U3591 (N_3591,In_133,In_642);
xnor U3592 (N_3592,In_759,In_469);
xnor U3593 (N_3593,In_572,In_701);
nand U3594 (N_3594,In_1358,In_1667);
nand U3595 (N_3595,In_52,In_121);
nand U3596 (N_3596,In_1194,In_1739);
nor U3597 (N_3597,In_861,In_892);
or U3598 (N_3598,In_1219,In_584);
xnor U3599 (N_3599,In_1561,In_819);
nand U3600 (N_3600,In_157,In_1086);
nor U3601 (N_3601,In_1793,In_1979);
nor U3602 (N_3602,In_586,In_1883);
xnor U3603 (N_3603,In_470,In_325);
or U3604 (N_3604,In_1171,In_1450);
and U3605 (N_3605,In_684,In_656);
and U3606 (N_3606,In_817,In_1674);
nand U3607 (N_3607,In_1689,In_284);
and U3608 (N_3608,In_71,In_519);
nor U3609 (N_3609,In_1025,In_1863);
nand U3610 (N_3610,In_1796,In_205);
nor U3611 (N_3611,In_1739,In_1700);
nor U3612 (N_3612,In_885,In_1481);
and U3613 (N_3613,In_334,In_1348);
nor U3614 (N_3614,In_1132,In_915);
nor U3615 (N_3615,In_325,In_1470);
xor U3616 (N_3616,In_1089,In_1753);
nor U3617 (N_3617,In_432,In_211);
nor U3618 (N_3618,In_62,In_1047);
xnor U3619 (N_3619,In_1232,In_1856);
and U3620 (N_3620,In_1562,In_465);
nand U3621 (N_3621,In_763,In_1007);
nor U3622 (N_3622,In_1711,In_1011);
or U3623 (N_3623,In_1931,In_1712);
and U3624 (N_3624,In_222,In_897);
xnor U3625 (N_3625,In_598,In_1204);
and U3626 (N_3626,In_1752,In_347);
nand U3627 (N_3627,In_492,In_770);
or U3628 (N_3628,In_1502,In_30);
nand U3629 (N_3629,In_1095,In_1119);
or U3630 (N_3630,In_919,In_1964);
nor U3631 (N_3631,In_409,In_912);
xnor U3632 (N_3632,In_353,In_523);
xor U3633 (N_3633,In_472,In_840);
xor U3634 (N_3634,In_1588,In_867);
nor U3635 (N_3635,In_1687,In_1161);
xor U3636 (N_3636,In_887,In_443);
nor U3637 (N_3637,In_482,In_1977);
and U3638 (N_3638,In_747,In_1937);
xor U3639 (N_3639,In_641,In_1990);
or U3640 (N_3640,In_961,In_1145);
nand U3641 (N_3641,In_1249,In_1131);
xnor U3642 (N_3642,In_696,In_1213);
nand U3643 (N_3643,In_1208,In_1375);
xor U3644 (N_3644,In_998,In_816);
nor U3645 (N_3645,In_12,In_273);
nand U3646 (N_3646,In_1941,In_1026);
and U3647 (N_3647,In_1824,In_339);
nor U3648 (N_3648,In_1815,In_1989);
or U3649 (N_3649,In_1041,In_1866);
xnor U3650 (N_3650,In_1572,In_503);
and U3651 (N_3651,In_845,In_1829);
nand U3652 (N_3652,In_1112,In_11);
and U3653 (N_3653,In_1326,In_482);
or U3654 (N_3654,In_430,In_510);
or U3655 (N_3655,In_651,In_1245);
nor U3656 (N_3656,In_1799,In_872);
nor U3657 (N_3657,In_778,In_1424);
and U3658 (N_3658,In_1429,In_1559);
and U3659 (N_3659,In_1517,In_1336);
or U3660 (N_3660,In_908,In_1874);
nor U3661 (N_3661,In_784,In_257);
and U3662 (N_3662,In_1827,In_1875);
nor U3663 (N_3663,In_367,In_917);
nand U3664 (N_3664,In_379,In_1103);
and U3665 (N_3665,In_1647,In_1433);
and U3666 (N_3666,In_1348,In_205);
or U3667 (N_3667,In_1579,In_1619);
nor U3668 (N_3668,In_873,In_584);
xor U3669 (N_3669,In_1314,In_1657);
nand U3670 (N_3670,In_965,In_1402);
or U3671 (N_3671,In_846,In_1692);
or U3672 (N_3672,In_1693,In_1432);
xor U3673 (N_3673,In_1626,In_1166);
and U3674 (N_3674,In_1195,In_274);
nor U3675 (N_3675,In_1028,In_1786);
nor U3676 (N_3676,In_687,In_85);
and U3677 (N_3677,In_20,In_444);
and U3678 (N_3678,In_181,In_628);
xor U3679 (N_3679,In_1322,In_1289);
xor U3680 (N_3680,In_1914,In_1371);
or U3681 (N_3681,In_845,In_1489);
and U3682 (N_3682,In_1441,In_916);
nand U3683 (N_3683,In_1642,In_1063);
nor U3684 (N_3684,In_1638,In_115);
and U3685 (N_3685,In_286,In_1100);
nand U3686 (N_3686,In_968,In_535);
xnor U3687 (N_3687,In_573,In_217);
xor U3688 (N_3688,In_1026,In_1935);
or U3689 (N_3689,In_896,In_3);
and U3690 (N_3690,In_1829,In_1423);
or U3691 (N_3691,In_1849,In_798);
xnor U3692 (N_3692,In_299,In_868);
or U3693 (N_3693,In_877,In_1758);
and U3694 (N_3694,In_1952,In_798);
nor U3695 (N_3695,In_598,In_1627);
xor U3696 (N_3696,In_444,In_1252);
xnor U3697 (N_3697,In_1897,In_1433);
or U3698 (N_3698,In_1594,In_664);
xor U3699 (N_3699,In_1480,In_211);
nor U3700 (N_3700,In_81,In_1572);
and U3701 (N_3701,In_1396,In_477);
and U3702 (N_3702,In_1452,In_1541);
and U3703 (N_3703,In_47,In_593);
nor U3704 (N_3704,In_1527,In_1643);
and U3705 (N_3705,In_498,In_1706);
or U3706 (N_3706,In_98,In_402);
and U3707 (N_3707,In_281,In_1463);
xor U3708 (N_3708,In_372,In_79);
or U3709 (N_3709,In_1052,In_1068);
nor U3710 (N_3710,In_1577,In_194);
nand U3711 (N_3711,In_230,In_704);
xor U3712 (N_3712,In_496,In_1867);
xor U3713 (N_3713,In_1070,In_965);
and U3714 (N_3714,In_813,In_390);
nand U3715 (N_3715,In_1196,In_1066);
nand U3716 (N_3716,In_356,In_905);
or U3717 (N_3717,In_639,In_539);
nor U3718 (N_3718,In_1992,In_263);
nor U3719 (N_3719,In_1226,In_277);
xor U3720 (N_3720,In_1876,In_530);
or U3721 (N_3721,In_439,In_1773);
nor U3722 (N_3722,In_919,In_1166);
and U3723 (N_3723,In_1065,In_836);
xnor U3724 (N_3724,In_1272,In_30);
and U3725 (N_3725,In_1974,In_1826);
or U3726 (N_3726,In_1340,In_1419);
nand U3727 (N_3727,In_1447,In_118);
or U3728 (N_3728,In_328,In_1497);
xnor U3729 (N_3729,In_496,In_887);
xnor U3730 (N_3730,In_1105,In_1511);
nor U3731 (N_3731,In_1380,In_607);
and U3732 (N_3732,In_19,In_1386);
nand U3733 (N_3733,In_1755,In_1670);
nor U3734 (N_3734,In_1606,In_1271);
nor U3735 (N_3735,In_587,In_1179);
and U3736 (N_3736,In_1585,In_1586);
and U3737 (N_3737,In_1616,In_703);
or U3738 (N_3738,In_1559,In_798);
nand U3739 (N_3739,In_983,In_296);
xor U3740 (N_3740,In_1950,In_1399);
or U3741 (N_3741,In_1122,In_203);
nand U3742 (N_3742,In_101,In_271);
nand U3743 (N_3743,In_403,In_663);
nor U3744 (N_3744,In_1091,In_1999);
nand U3745 (N_3745,In_486,In_82);
nand U3746 (N_3746,In_1684,In_343);
or U3747 (N_3747,In_610,In_1229);
and U3748 (N_3748,In_183,In_1741);
nor U3749 (N_3749,In_416,In_1724);
or U3750 (N_3750,In_454,In_1049);
nand U3751 (N_3751,In_1397,In_138);
nor U3752 (N_3752,In_1977,In_1400);
or U3753 (N_3753,In_1940,In_1484);
nand U3754 (N_3754,In_1408,In_1393);
and U3755 (N_3755,In_1281,In_91);
nand U3756 (N_3756,In_1229,In_18);
nand U3757 (N_3757,In_1233,In_78);
or U3758 (N_3758,In_420,In_10);
nor U3759 (N_3759,In_1620,In_1673);
nand U3760 (N_3760,In_1935,In_747);
or U3761 (N_3761,In_930,In_1778);
or U3762 (N_3762,In_882,In_1492);
nor U3763 (N_3763,In_1339,In_1144);
nand U3764 (N_3764,In_505,In_88);
and U3765 (N_3765,In_274,In_1363);
or U3766 (N_3766,In_1162,In_1242);
nand U3767 (N_3767,In_373,In_487);
and U3768 (N_3768,In_259,In_1653);
and U3769 (N_3769,In_316,In_1771);
xnor U3770 (N_3770,In_713,In_1080);
nor U3771 (N_3771,In_962,In_7);
nor U3772 (N_3772,In_186,In_121);
nor U3773 (N_3773,In_1716,In_1723);
xnor U3774 (N_3774,In_1066,In_1580);
nand U3775 (N_3775,In_1406,In_1367);
and U3776 (N_3776,In_152,In_768);
and U3777 (N_3777,In_1230,In_1077);
nand U3778 (N_3778,In_359,In_1882);
xor U3779 (N_3779,In_430,In_1045);
xnor U3780 (N_3780,In_1302,In_1170);
xor U3781 (N_3781,In_762,In_1858);
and U3782 (N_3782,In_1436,In_1006);
and U3783 (N_3783,In_1170,In_1033);
and U3784 (N_3784,In_76,In_997);
or U3785 (N_3785,In_537,In_1576);
xnor U3786 (N_3786,In_1445,In_715);
nor U3787 (N_3787,In_121,In_1884);
nor U3788 (N_3788,In_1390,In_1205);
and U3789 (N_3789,In_1199,In_938);
xnor U3790 (N_3790,In_194,In_914);
nand U3791 (N_3791,In_858,In_1685);
nor U3792 (N_3792,In_449,In_1214);
nor U3793 (N_3793,In_1826,In_1669);
and U3794 (N_3794,In_124,In_967);
nor U3795 (N_3795,In_115,In_1355);
nand U3796 (N_3796,In_62,In_124);
nor U3797 (N_3797,In_1439,In_1270);
or U3798 (N_3798,In_1841,In_1506);
and U3799 (N_3799,In_1114,In_75);
xor U3800 (N_3800,In_716,In_143);
or U3801 (N_3801,In_887,In_1510);
nor U3802 (N_3802,In_377,In_1940);
or U3803 (N_3803,In_1536,In_1473);
or U3804 (N_3804,In_1960,In_1797);
xor U3805 (N_3805,In_1527,In_1594);
nor U3806 (N_3806,In_1914,In_1168);
nand U3807 (N_3807,In_1578,In_1952);
xor U3808 (N_3808,In_1906,In_1241);
nor U3809 (N_3809,In_1946,In_1308);
nand U3810 (N_3810,In_1128,In_1604);
nor U3811 (N_3811,In_426,In_1539);
or U3812 (N_3812,In_415,In_1733);
nor U3813 (N_3813,In_902,In_1861);
xor U3814 (N_3814,In_1984,In_1298);
nand U3815 (N_3815,In_51,In_1941);
xnor U3816 (N_3816,In_645,In_1952);
or U3817 (N_3817,In_1615,In_1850);
nor U3818 (N_3818,In_631,In_1485);
and U3819 (N_3819,In_1536,In_1730);
and U3820 (N_3820,In_1980,In_1697);
and U3821 (N_3821,In_844,In_1800);
xor U3822 (N_3822,In_345,In_164);
nand U3823 (N_3823,In_1076,In_806);
xor U3824 (N_3824,In_895,In_983);
or U3825 (N_3825,In_1316,In_328);
and U3826 (N_3826,In_1251,In_36);
nor U3827 (N_3827,In_1229,In_1167);
xnor U3828 (N_3828,In_1071,In_1279);
and U3829 (N_3829,In_1351,In_1566);
nor U3830 (N_3830,In_82,In_934);
nor U3831 (N_3831,In_869,In_1411);
nor U3832 (N_3832,In_343,In_767);
and U3833 (N_3833,In_1262,In_226);
or U3834 (N_3834,In_982,In_819);
or U3835 (N_3835,In_356,In_1700);
and U3836 (N_3836,In_626,In_486);
or U3837 (N_3837,In_315,In_363);
and U3838 (N_3838,In_1729,In_1830);
and U3839 (N_3839,In_1478,In_728);
xnor U3840 (N_3840,In_1775,In_1963);
xnor U3841 (N_3841,In_546,In_51);
or U3842 (N_3842,In_1705,In_1984);
nand U3843 (N_3843,In_1485,In_1669);
nor U3844 (N_3844,In_686,In_1338);
nand U3845 (N_3845,In_1629,In_1160);
or U3846 (N_3846,In_1554,In_721);
or U3847 (N_3847,In_1572,In_1271);
and U3848 (N_3848,In_901,In_815);
and U3849 (N_3849,In_377,In_352);
or U3850 (N_3850,In_1865,In_875);
nand U3851 (N_3851,In_1648,In_223);
nor U3852 (N_3852,In_1547,In_1998);
xor U3853 (N_3853,In_1130,In_954);
nand U3854 (N_3854,In_1087,In_1936);
nor U3855 (N_3855,In_1830,In_1025);
and U3856 (N_3856,In_1354,In_1071);
nand U3857 (N_3857,In_223,In_1779);
or U3858 (N_3858,In_1397,In_1723);
and U3859 (N_3859,In_1108,In_1584);
and U3860 (N_3860,In_1183,In_533);
nand U3861 (N_3861,In_606,In_505);
nand U3862 (N_3862,In_194,In_827);
nor U3863 (N_3863,In_0,In_1409);
and U3864 (N_3864,In_1521,In_43);
xnor U3865 (N_3865,In_195,In_906);
nor U3866 (N_3866,In_1659,In_1319);
xor U3867 (N_3867,In_305,In_1446);
and U3868 (N_3868,In_882,In_172);
nor U3869 (N_3869,In_108,In_420);
and U3870 (N_3870,In_563,In_1577);
xor U3871 (N_3871,In_827,In_1313);
xor U3872 (N_3872,In_1901,In_612);
or U3873 (N_3873,In_1813,In_47);
xor U3874 (N_3874,In_1905,In_1456);
xnor U3875 (N_3875,In_194,In_1810);
nand U3876 (N_3876,In_822,In_1036);
and U3877 (N_3877,In_457,In_1589);
and U3878 (N_3878,In_1386,In_1413);
or U3879 (N_3879,In_263,In_881);
nor U3880 (N_3880,In_1556,In_370);
xor U3881 (N_3881,In_1541,In_387);
and U3882 (N_3882,In_1672,In_1811);
nand U3883 (N_3883,In_124,In_1712);
xnor U3884 (N_3884,In_1628,In_515);
or U3885 (N_3885,In_450,In_894);
nor U3886 (N_3886,In_551,In_1997);
and U3887 (N_3887,In_385,In_285);
nand U3888 (N_3888,In_650,In_410);
and U3889 (N_3889,In_1883,In_753);
nand U3890 (N_3890,In_1713,In_582);
or U3891 (N_3891,In_714,In_26);
or U3892 (N_3892,In_162,In_1177);
and U3893 (N_3893,In_1066,In_236);
nand U3894 (N_3894,In_616,In_595);
nor U3895 (N_3895,In_554,In_87);
nor U3896 (N_3896,In_467,In_1528);
and U3897 (N_3897,In_1799,In_1428);
nand U3898 (N_3898,In_779,In_733);
or U3899 (N_3899,In_608,In_1335);
or U3900 (N_3900,In_1469,In_1985);
or U3901 (N_3901,In_1696,In_480);
or U3902 (N_3902,In_1666,In_268);
nor U3903 (N_3903,In_1017,In_1676);
nand U3904 (N_3904,In_1118,In_259);
nor U3905 (N_3905,In_119,In_1851);
nor U3906 (N_3906,In_214,In_790);
xor U3907 (N_3907,In_71,In_1397);
nor U3908 (N_3908,In_1385,In_152);
and U3909 (N_3909,In_328,In_1242);
xor U3910 (N_3910,In_1980,In_726);
xnor U3911 (N_3911,In_831,In_1128);
nor U3912 (N_3912,In_1106,In_518);
nor U3913 (N_3913,In_833,In_297);
xor U3914 (N_3914,In_752,In_1940);
xnor U3915 (N_3915,In_1317,In_1160);
or U3916 (N_3916,In_599,In_1555);
nor U3917 (N_3917,In_500,In_1302);
and U3918 (N_3918,In_604,In_520);
or U3919 (N_3919,In_135,In_409);
or U3920 (N_3920,In_942,In_1741);
xor U3921 (N_3921,In_1339,In_1704);
nor U3922 (N_3922,In_1969,In_1900);
or U3923 (N_3923,In_1023,In_1341);
xor U3924 (N_3924,In_739,In_1551);
nor U3925 (N_3925,In_949,In_1624);
xor U3926 (N_3926,In_465,In_179);
and U3927 (N_3927,In_1879,In_1295);
and U3928 (N_3928,In_623,In_1176);
nor U3929 (N_3929,In_773,In_1586);
nor U3930 (N_3930,In_1460,In_998);
nand U3931 (N_3931,In_1826,In_1856);
or U3932 (N_3932,In_172,In_1323);
xnor U3933 (N_3933,In_1355,In_168);
nand U3934 (N_3934,In_666,In_557);
xor U3935 (N_3935,In_623,In_753);
nor U3936 (N_3936,In_839,In_1011);
or U3937 (N_3937,In_550,In_681);
and U3938 (N_3938,In_1681,In_1573);
or U3939 (N_3939,In_125,In_954);
xnor U3940 (N_3940,In_737,In_1986);
or U3941 (N_3941,In_653,In_109);
xnor U3942 (N_3942,In_1024,In_1217);
nand U3943 (N_3943,In_1141,In_1071);
or U3944 (N_3944,In_696,In_1089);
xnor U3945 (N_3945,In_1098,In_1417);
xnor U3946 (N_3946,In_1343,In_98);
xnor U3947 (N_3947,In_159,In_307);
nor U3948 (N_3948,In_1015,In_1525);
xnor U3949 (N_3949,In_748,In_1570);
nand U3950 (N_3950,In_5,In_1582);
nand U3951 (N_3951,In_1303,In_1657);
and U3952 (N_3952,In_1778,In_558);
nand U3953 (N_3953,In_116,In_517);
or U3954 (N_3954,In_1665,In_1211);
and U3955 (N_3955,In_468,In_799);
and U3956 (N_3956,In_151,In_1188);
nand U3957 (N_3957,In_1315,In_982);
xnor U3958 (N_3958,In_1586,In_414);
nor U3959 (N_3959,In_937,In_1141);
xnor U3960 (N_3960,In_1,In_1425);
and U3961 (N_3961,In_1601,In_1358);
and U3962 (N_3962,In_1078,In_22);
nand U3963 (N_3963,In_803,In_1861);
xor U3964 (N_3964,In_1926,In_611);
or U3965 (N_3965,In_1030,In_1966);
nor U3966 (N_3966,In_414,In_658);
xnor U3967 (N_3967,In_1838,In_68);
xnor U3968 (N_3968,In_571,In_1307);
xor U3969 (N_3969,In_1032,In_808);
or U3970 (N_3970,In_739,In_476);
nand U3971 (N_3971,In_458,In_587);
nor U3972 (N_3972,In_1485,In_1196);
nand U3973 (N_3973,In_476,In_442);
nor U3974 (N_3974,In_228,In_1216);
and U3975 (N_3975,In_432,In_283);
nand U3976 (N_3976,In_283,In_1413);
or U3977 (N_3977,In_812,In_1554);
or U3978 (N_3978,In_1340,In_1224);
nor U3979 (N_3979,In_1949,In_352);
and U3980 (N_3980,In_1212,In_1044);
or U3981 (N_3981,In_1740,In_1560);
or U3982 (N_3982,In_104,In_658);
and U3983 (N_3983,In_210,In_1878);
nand U3984 (N_3984,In_1574,In_446);
nand U3985 (N_3985,In_1119,In_1709);
and U3986 (N_3986,In_1271,In_920);
xor U3987 (N_3987,In_1203,In_390);
nor U3988 (N_3988,In_512,In_1795);
xnor U3989 (N_3989,In_951,In_1260);
and U3990 (N_3990,In_1888,In_1491);
xor U3991 (N_3991,In_924,In_1605);
xor U3992 (N_3992,In_843,In_785);
xnor U3993 (N_3993,In_1846,In_212);
nand U3994 (N_3994,In_1122,In_1612);
or U3995 (N_3995,In_1805,In_677);
or U3996 (N_3996,In_1051,In_1101);
or U3997 (N_3997,In_1267,In_1803);
nor U3998 (N_3998,In_433,In_1872);
xnor U3999 (N_3999,In_1133,In_824);
nor U4000 (N_4000,N_3211,N_2280);
nor U4001 (N_4001,N_446,N_560);
and U4002 (N_4002,N_2357,N_1004);
or U4003 (N_4003,N_2894,N_3959);
and U4004 (N_4004,N_108,N_2942);
nor U4005 (N_4005,N_2835,N_2542);
and U4006 (N_4006,N_2897,N_3765);
and U4007 (N_4007,N_334,N_1255);
xnor U4008 (N_4008,N_601,N_2938);
and U4009 (N_4009,N_736,N_1054);
nand U4010 (N_4010,N_1641,N_1207);
xor U4011 (N_4011,N_1121,N_7);
nor U4012 (N_4012,N_2564,N_3213);
or U4013 (N_4013,N_336,N_478);
or U4014 (N_4014,N_2778,N_713);
or U4015 (N_4015,N_3667,N_424);
and U4016 (N_4016,N_1140,N_2220);
nand U4017 (N_4017,N_1378,N_452);
xor U4018 (N_4018,N_3849,N_2341);
nor U4019 (N_4019,N_2112,N_2201);
xnor U4020 (N_4020,N_1721,N_699);
and U4021 (N_4021,N_3463,N_2336);
and U4022 (N_4022,N_3989,N_2170);
nand U4023 (N_4023,N_2563,N_2781);
or U4024 (N_4024,N_3508,N_2538);
xor U4025 (N_4025,N_89,N_1489);
or U4026 (N_4026,N_2761,N_3963);
xor U4027 (N_4027,N_222,N_647);
or U4028 (N_4028,N_884,N_3200);
or U4029 (N_4029,N_1772,N_3399);
or U4030 (N_4030,N_145,N_241);
nand U4031 (N_4031,N_3680,N_724);
nand U4032 (N_4032,N_3859,N_2192);
nor U4033 (N_4033,N_1666,N_2);
and U4034 (N_4034,N_2382,N_2992);
nor U4035 (N_4035,N_2074,N_980);
or U4036 (N_4036,N_114,N_3591);
xnor U4037 (N_4037,N_1750,N_1153);
nand U4038 (N_4038,N_2474,N_2747);
xnor U4039 (N_4039,N_1598,N_956);
nand U4040 (N_4040,N_1946,N_3801);
nand U4041 (N_4041,N_3144,N_1711);
nand U4042 (N_4042,N_3044,N_2130);
nor U4043 (N_4043,N_1829,N_1484);
and U4044 (N_4044,N_252,N_213);
nor U4045 (N_4045,N_210,N_3363);
nand U4046 (N_4046,N_474,N_2369);
and U4047 (N_4047,N_3128,N_3109);
nand U4048 (N_4048,N_144,N_1234);
nor U4049 (N_4049,N_3819,N_1014);
and U4050 (N_4050,N_9,N_3013);
nand U4051 (N_4051,N_3600,N_1548);
nor U4052 (N_4052,N_3390,N_1842);
nand U4053 (N_4053,N_3284,N_3827);
and U4054 (N_4054,N_2375,N_3853);
nand U4055 (N_4055,N_2818,N_2719);
nand U4056 (N_4056,N_1016,N_47);
xor U4057 (N_4057,N_1464,N_3154);
and U4058 (N_4058,N_3504,N_2353);
and U4059 (N_4059,N_2775,N_624);
and U4060 (N_4060,N_2198,N_3650);
nor U4061 (N_4061,N_1863,N_3442);
nor U4062 (N_4062,N_303,N_2915);
nand U4063 (N_4063,N_1594,N_3522);
xnor U4064 (N_4064,N_357,N_1293);
or U4065 (N_4065,N_653,N_2588);
xor U4066 (N_4066,N_1786,N_1188);
or U4067 (N_4067,N_3655,N_3852);
nor U4068 (N_4068,N_3358,N_3876);
nand U4069 (N_4069,N_2326,N_1410);
nand U4070 (N_4070,N_754,N_543);
xor U4071 (N_4071,N_1189,N_1538);
nand U4072 (N_4072,N_3751,N_1569);
and U4073 (N_4073,N_1661,N_3325);
nor U4074 (N_4074,N_3550,N_2987);
nand U4075 (N_4075,N_1232,N_1689);
nor U4076 (N_4076,N_3884,N_2432);
and U4077 (N_4077,N_2872,N_3315);
or U4078 (N_4078,N_94,N_605);
xnor U4079 (N_4079,N_1011,N_1333);
nor U4080 (N_4080,N_3152,N_1555);
xnor U4081 (N_4081,N_3964,N_1197);
xor U4082 (N_4082,N_1665,N_3527);
or U4083 (N_4083,N_1698,N_273);
xor U4084 (N_4084,N_3294,N_3930);
or U4085 (N_4085,N_1107,N_522);
xor U4086 (N_4086,N_3967,N_2306);
or U4087 (N_4087,N_2355,N_1892);
nor U4088 (N_4088,N_1185,N_136);
xor U4089 (N_4089,N_1894,N_3398);
nor U4090 (N_4090,N_383,N_3245);
or U4091 (N_4091,N_3028,N_1804);
nand U4092 (N_4092,N_1568,N_2820);
nor U4093 (N_4093,N_2845,N_3259);
or U4094 (N_4094,N_323,N_3803);
or U4095 (N_4095,N_3632,N_3987);
and U4096 (N_4096,N_235,N_564);
nor U4097 (N_4097,N_3868,N_2299);
nand U4098 (N_4098,N_3924,N_990);
nor U4099 (N_4099,N_1298,N_2011);
and U4100 (N_4100,N_1431,N_1162);
nand U4101 (N_4101,N_1953,N_2420);
or U4102 (N_4102,N_1134,N_166);
nand U4103 (N_4103,N_2052,N_416);
nor U4104 (N_4104,N_3715,N_1768);
xnor U4105 (N_4105,N_2611,N_291);
or U4106 (N_4106,N_185,N_74);
and U4107 (N_4107,N_1270,N_3675);
xor U4108 (N_4108,N_2337,N_3047);
and U4109 (N_4109,N_2683,N_3186);
nand U4110 (N_4110,N_2970,N_860);
nand U4111 (N_4111,N_3922,N_81);
and U4112 (N_4112,N_1480,N_682);
and U4113 (N_4113,N_1691,N_338);
nor U4114 (N_4114,N_2486,N_3039);
nor U4115 (N_4115,N_2605,N_3572);
nand U4116 (N_4116,N_1334,N_1022);
xnor U4117 (N_4117,N_684,N_1356);
nor U4118 (N_4118,N_2493,N_2504);
and U4119 (N_4119,N_435,N_2748);
and U4120 (N_4120,N_2237,N_757);
or U4121 (N_4121,N_2904,N_3826);
nand U4122 (N_4122,N_422,N_1180);
or U4123 (N_4123,N_2986,N_70);
nand U4124 (N_4124,N_1025,N_3000);
nor U4125 (N_4125,N_3763,N_3906);
nand U4126 (N_4126,N_1890,N_2236);
or U4127 (N_4127,N_1936,N_2997);
nor U4128 (N_4128,N_1605,N_2230);
nor U4129 (N_4129,N_1531,N_831);
xor U4130 (N_4130,N_1530,N_3307);
nor U4131 (N_4131,N_401,N_1070);
and U4132 (N_4132,N_15,N_1311);
or U4133 (N_4133,N_1702,N_2955);
nor U4134 (N_4134,N_1460,N_302);
and U4135 (N_4135,N_2534,N_168);
or U4136 (N_4136,N_308,N_680);
and U4137 (N_4137,N_3085,N_343);
xnor U4138 (N_4138,N_3339,N_355);
or U4139 (N_4139,N_2557,N_2479);
or U4140 (N_4140,N_2892,N_2217);
nand U4141 (N_4141,N_1051,N_3753);
nand U4142 (N_4142,N_2741,N_24);
xor U4143 (N_4143,N_3770,N_3175);
or U4144 (N_4144,N_3203,N_3230);
and U4145 (N_4145,N_3406,N_763);
nand U4146 (N_4146,N_3419,N_2679);
nand U4147 (N_4147,N_756,N_1175);
nor U4148 (N_4148,N_3961,N_413);
nor U4149 (N_4149,N_2340,N_2949);
nor U4150 (N_4150,N_312,N_2405);
xnor U4151 (N_4151,N_1331,N_2789);
nand U4152 (N_4152,N_2971,N_2703);
xor U4153 (N_4153,N_2343,N_820);
and U4154 (N_4154,N_130,N_1554);
nand U4155 (N_4155,N_1821,N_2270);
nand U4156 (N_4156,N_1874,N_2169);
xnor U4157 (N_4157,N_2219,N_361);
or U4158 (N_4158,N_2017,N_3179);
or U4159 (N_4159,N_1727,N_1828);
or U4160 (N_4160,N_2529,N_228);
and U4161 (N_4161,N_854,N_481);
nor U4162 (N_4162,N_2762,N_1098);
nand U4163 (N_4163,N_1681,N_1583);
and U4164 (N_4164,N_72,N_2351);
nor U4165 (N_4165,N_1044,N_2344);
xnor U4166 (N_4166,N_1811,N_2332);
nand U4167 (N_4167,N_3180,N_1292);
or U4168 (N_4168,N_193,N_1013);
xnor U4169 (N_4169,N_322,N_1744);
xor U4170 (N_4170,N_784,N_3953);
and U4171 (N_4171,N_3617,N_1000);
nor U4172 (N_4172,N_1680,N_2587);
and U4173 (N_4173,N_2796,N_176);
xnor U4174 (N_4174,N_3124,N_3172);
nor U4175 (N_4175,N_945,N_2056);
nand U4176 (N_4176,N_491,N_760);
and U4177 (N_4177,N_472,N_2963);
nor U4178 (N_4178,N_1478,N_3764);
or U4179 (N_4179,N_3701,N_2846);
xor U4180 (N_4180,N_2144,N_5);
xor U4181 (N_4181,N_959,N_575);
nand U4182 (N_4182,N_3791,N_692);
nand U4183 (N_4183,N_1083,N_1254);
and U4184 (N_4184,N_2480,N_3666);
xor U4185 (N_4185,N_1622,N_1342);
and U4186 (N_4186,N_3931,N_2311);
or U4187 (N_4187,N_525,N_3240);
xor U4188 (N_4188,N_2559,N_910);
xor U4189 (N_4189,N_45,N_3225);
xnor U4190 (N_4190,N_3118,N_1852);
or U4191 (N_4191,N_3137,N_588);
nand U4192 (N_4192,N_3147,N_2126);
or U4193 (N_4193,N_1565,N_694);
nor U4194 (N_4194,N_1494,N_3705);
nand U4195 (N_4195,N_1048,N_1704);
and U4196 (N_4196,N_3596,N_3978);
or U4197 (N_4197,N_2395,N_3078);
xor U4198 (N_4198,N_419,N_3760);
nor U4199 (N_4199,N_3627,N_128);
nand U4200 (N_4200,N_3212,N_2798);
nor U4201 (N_4201,N_3829,N_1323);
nand U4202 (N_4202,N_2766,N_1700);
or U4203 (N_4203,N_3773,N_983);
or U4204 (N_4204,N_1558,N_129);
or U4205 (N_4205,N_3094,N_3816);
xor U4206 (N_4206,N_3539,N_236);
nand U4207 (N_4207,N_3703,N_3483);
or U4208 (N_4208,N_2252,N_3145);
nor U4209 (N_4209,N_567,N_2404);
and U4210 (N_4210,N_1145,N_589);
and U4211 (N_4211,N_2934,N_2460);
nand U4212 (N_4212,N_3707,N_2153);
xnor U4213 (N_4213,N_2046,N_3033);
xnor U4214 (N_4214,N_3559,N_2014);
nand U4215 (N_4215,N_986,N_2804);
or U4216 (N_4216,N_0,N_1424);
nand U4217 (N_4217,N_3811,N_86);
or U4218 (N_4218,N_1643,N_229);
and U4219 (N_4219,N_1682,N_3642);
nand U4220 (N_4220,N_1910,N_2799);
nand U4221 (N_4221,N_3725,N_3441);
nand U4222 (N_4222,N_3063,N_3415);
nor U4223 (N_4223,N_1642,N_2523);
nand U4224 (N_4224,N_2364,N_2216);
or U4225 (N_4225,N_121,N_2385);
nand U4226 (N_4226,N_845,N_3052);
xnor U4227 (N_4227,N_3165,N_1732);
or U4228 (N_4228,N_2854,N_3332);
nor U4229 (N_4229,N_1593,N_1461);
nand U4230 (N_4230,N_3834,N_873);
xor U4231 (N_4231,N_220,N_1944);
and U4232 (N_4232,N_1741,N_2419);
nor U4233 (N_4233,N_561,N_2589);
nand U4234 (N_4234,N_142,N_3335);
nor U4235 (N_4235,N_3322,N_181);
nor U4236 (N_4236,N_991,N_2288);
nor U4237 (N_4237,N_348,N_3302);
or U4238 (N_4238,N_1778,N_2547);
and U4239 (N_4239,N_1199,N_3251);
xnor U4240 (N_4240,N_1045,N_2768);
nand U4241 (N_4241,N_789,N_2359);
xor U4242 (N_4242,N_300,N_1168);
or U4243 (N_4243,N_2549,N_3818);
nor U4244 (N_4244,N_1644,N_2586);
nand U4245 (N_4245,N_1658,N_107);
nor U4246 (N_4246,N_2612,N_88);
and U4247 (N_4247,N_3936,N_2078);
and U4248 (N_4248,N_2195,N_2833);
or U4249 (N_4249,N_979,N_507);
nand U4250 (N_4250,N_1784,N_2541);
or U4251 (N_4251,N_1261,N_501);
or U4252 (N_4252,N_3523,N_1522);
and U4253 (N_4253,N_556,N_857);
nor U4254 (N_4254,N_3841,N_2304);
nor U4255 (N_4255,N_2965,N_1190);
nand U4256 (N_4256,N_1501,N_2993);
nand U4257 (N_4257,N_1922,N_3606);
nor U4258 (N_4258,N_3969,N_2654);
nor U4259 (N_4259,N_686,N_3288);
or U4260 (N_4260,N_1363,N_365);
xnor U4261 (N_4261,N_3379,N_61);
nand U4262 (N_4262,N_921,N_3439);
nor U4263 (N_4263,N_1348,N_731);
nand U4264 (N_4264,N_1679,N_2321);
or U4265 (N_4265,N_1792,N_2770);
nor U4266 (N_4266,N_151,N_2712);
nor U4267 (N_4267,N_2513,N_3757);
xor U4268 (N_4268,N_3243,N_1955);
or U4269 (N_4269,N_1135,N_2146);
and U4270 (N_4270,N_3222,N_270);
or U4271 (N_4271,N_1634,N_1653);
or U4272 (N_4272,N_1219,N_2810);
xor U4273 (N_4273,N_2642,N_170);
and U4274 (N_4274,N_1495,N_1649);
and U4275 (N_4275,N_3337,N_2035);
nand U4276 (N_4276,N_2805,N_1237);
xnor U4277 (N_4277,N_3955,N_3970);
or U4278 (N_4278,N_342,N_3656);
nand U4279 (N_4279,N_1079,N_3236);
nand U4280 (N_4280,N_1867,N_485);
nor U4281 (N_4281,N_2206,N_3531);
xor U4282 (N_4282,N_1984,N_2138);
xnor U4283 (N_4283,N_3050,N_1122);
xnor U4284 (N_4284,N_2692,N_3761);
or U4285 (N_4285,N_3326,N_263);
xor U4286 (N_4286,N_651,N_3329);
nand U4287 (N_4287,N_812,N_172);
or U4288 (N_4288,N_3939,N_3274);
nand U4289 (N_4289,N_3500,N_689);
or U4290 (N_4290,N_2196,N_3613);
nand U4291 (N_4291,N_2456,N_3330);
nor U4292 (N_4292,N_412,N_3071);
xnor U4293 (N_4293,N_664,N_1950);
xor U4294 (N_4294,N_1,N_1748);
nor U4295 (N_4295,N_883,N_60);
and U4296 (N_4296,N_3234,N_548);
xor U4297 (N_4297,N_1785,N_1918);
xor U4298 (N_4298,N_3120,N_1798);
nand U4299 (N_4299,N_3092,N_1796);
and U4300 (N_4300,N_2950,N_2828);
nand U4301 (N_4301,N_2840,N_480);
nor U4302 (N_4302,N_862,N_3110);
xnor U4303 (N_4303,N_197,N_3359);
nor U4304 (N_4304,N_251,N_2527);
or U4305 (N_4305,N_1940,N_3723);
or U4306 (N_4306,N_917,N_584);
nand U4307 (N_4307,N_1332,N_2576);
nor U4308 (N_4308,N_3995,N_3507);
nor U4309 (N_4309,N_3250,N_1765);
and U4310 (N_4310,N_2127,N_3608);
or U4311 (N_4311,N_1813,N_3425);
or U4312 (N_4312,N_2649,N_1305);
or U4313 (N_4313,N_3823,N_3233);
nor U4314 (N_4314,N_1755,N_3204);
and U4315 (N_4315,N_2621,N_2769);
nor U4316 (N_4316,N_1932,N_3355);
or U4317 (N_4317,N_3004,N_1817);
nor U4318 (N_4318,N_2763,N_238);
and U4319 (N_4319,N_75,N_3825);
nand U4320 (N_4320,N_2851,N_1154);
and U4321 (N_4321,N_2041,N_2173);
xor U4322 (N_4322,N_2390,N_3848);
and U4323 (N_4323,N_816,N_2086);
xnor U4324 (N_4324,N_3903,N_1490);
nand U4325 (N_4325,N_498,N_863);
nand U4326 (N_4326,N_2842,N_3331);
nand U4327 (N_4327,N_3889,N_3417);
nor U4328 (N_4328,N_965,N_943);
xor U4329 (N_4329,N_3453,N_2760);
nor U4330 (N_4330,N_1967,N_2994);
or U4331 (N_4331,N_1182,N_3985);
nand U4332 (N_4332,N_2881,N_1703);
xor U4333 (N_4333,N_2543,N_1878);
xor U4334 (N_4334,N_3347,N_1046);
xnor U4335 (N_4335,N_2537,N_3717);
or U4336 (N_4336,N_2289,N_2686);
or U4337 (N_4337,N_55,N_1393);
nand U4338 (N_4338,N_1758,N_2806);
xnor U4339 (N_4339,N_3045,N_1414);
and U4340 (N_4340,N_3865,N_1186);
and U4341 (N_4341,N_811,N_1043);
or U4342 (N_4342,N_1272,N_3652);
nand U4343 (N_4343,N_1344,N_1299);
and U4344 (N_4344,N_1971,N_661);
nand U4345 (N_4345,N_2607,N_1990);
and U4346 (N_4346,N_1080,N_2440);
xor U4347 (N_4347,N_379,N_1730);
and U4348 (N_4348,N_1656,N_173);
nand U4349 (N_4349,N_2874,N_3438);
and U4350 (N_4350,N_3863,N_1652);
and U4351 (N_4351,N_3007,N_3982);
xor U4352 (N_4352,N_3609,N_1169);
and U4353 (N_4353,N_704,N_1435);
and U4354 (N_4354,N_3575,N_3779);
and U4355 (N_4355,N_2862,N_78);
or U4356 (N_4356,N_415,N_1108);
or U4357 (N_4357,N_3173,N_349);
or U4358 (N_4358,N_1419,N_1877);
and U4359 (N_4359,N_3377,N_2147);
nor U4360 (N_4360,N_1542,N_592);
or U4361 (N_4361,N_2933,N_879);
or U4362 (N_4362,N_11,N_182);
nor U4363 (N_4363,N_518,N_2204);
xor U4364 (N_4364,N_146,N_1347);
nand U4365 (N_4365,N_3545,N_881);
and U4366 (N_4366,N_1525,N_2633);
and U4367 (N_4367,N_3843,N_1243);
nand U4368 (N_4368,N_3934,N_3221);
nor U4369 (N_4369,N_2227,N_1602);
nand U4370 (N_4370,N_2579,N_3919);
or U4371 (N_4371,N_2070,N_397);
or U4372 (N_4372,N_2313,N_1017);
nor U4373 (N_4373,N_420,N_1557);
nand U4374 (N_4374,N_3464,N_3114);
and U4375 (N_4375,N_10,N_818);
nand U4376 (N_4376,N_3475,N_2729);
nand U4377 (N_4377,N_558,N_475);
and U4378 (N_4378,N_1306,N_1581);
nor U4379 (N_4379,N_2439,N_3206);
nand U4380 (N_4380,N_3407,N_2831);
xor U4381 (N_4381,N_1773,N_712);
or U4382 (N_4382,N_1826,N_2455);
nor U4383 (N_4383,N_64,N_3719);
and U4384 (N_4384,N_368,N_1437);
nor U4385 (N_4385,N_1767,N_1577);
nand U4386 (N_4386,N_2210,N_3943);
nand U4387 (N_4387,N_2320,N_775);
nor U4388 (N_4388,N_1159,N_505);
xnor U4389 (N_4389,N_1650,N_3538);
nor U4390 (N_4390,N_2106,N_1449);
or U4391 (N_4391,N_3948,N_1274);
nand U4392 (N_4392,N_2389,N_1975);
nor U4393 (N_4393,N_2837,N_2454);
and U4394 (N_4394,N_3011,N_635);
and U4395 (N_4395,N_3309,N_1897);
xnor U4396 (N_4396,N_2451,N_3074);
nor U4397 (N_4397,N_51,N_2121);
xnor U4398 (N_4398,N_866,N_2852);
xor U4399 (N_4399,N_287,N_1835);
nand U4400 (N_4400,N_3401,N_685);
xnor U4401 (N_4401,N_2575,N_1756);
and U4402 (N_4402,N_1279,N_2421);
nor U4403 (N_4403,N_2241,N_3477);
or U4404 (N_4404,N_1409,N_2802);
nor U4405 (N_4405,N_48,N_3933);
and U4406 (N_4406,N_1761,N_369);
or U4407 (N_4407,N_1510,N_950);
nand U4408 (N_4408,N_1033,N_288);
and U4409 (N_4409,N_1336,N_1294);
nand U4410 (N_4410,N_2816,N_2923);
or U4411 (N_4411,N_998,N_604);
xor U4412 (N_4412,N_255,N_3893);
or U4413 (N_4413,N_2296,N_285);
nor U4414 (N_4414,N_1933,N_2136);
xor U4415 (N_4415,N_3228,N_1223);
xnor U4416 (N_4416,N_3083,N_3542);
nor U4417 (N_4417,N_3885,N_2316);
nand U4418 (N_4418,N_1533,N_586);
and U4419 (N_4419,N_809,N_1503);
and U4420 (N_4420,N_2941,N_3972);
or U4421 (N_4421,N_741,N_3295);
nand U4422 (N_4422,N_3008,N_3557);
or U4423 (N_4423,N_3878,N_2600);
and U4424 (N_4424,N_538,N_1969);
xnor U4425 (N_4425,N_3741,N_3014);
xor U4426 (N_4426,N_2032,N_3456);
nor U4427 (N_4427,N_62,N_3744);
or U4428 (N_4428,N_2279,N_1754);
nor U4429 (N_4429,N_1717,N_1405);
nand U4430 (N_4430,N_386,N_3730);
xnor U4431 (N_4431,N_3198,N_2723);
or U4432 (N_4432,N_566,N_852);
xor U4433 (N_4433,N_3605,N_8);
nand U4434 (N_4434,N_3368,N_1167);
xnor U4435 (N_4435,N_3663,N_98);
or U4436 (N_4436,N_2853,N_849);
or U4437 (N_4437,N_1091,N_2444);
xor U4438 (N_4438,N_3672,N_3537);
nor U4439 (N_4439,N_244,N_795);
nor U4440 (N_4440,N_769,N_2877);
and U4441 (N_4441,N_1442,N_780);
nor U4442 (N_4442,N_594,N_2757);
and U4443 (N_4443,N_1069,N_2096);
nand U4444 (N_4444,N_2660,N_722);
nor U4445 (N_4445,N_3001,N_2870);
xor U4446 (N_4446,N_721,N_3587);
and U4447 (N_4447,N_3755,N_2259);
xnor U4448 (N_4448,N_3595,N_2208);
and U4449 (N_4449,N_3266,N_3641);
and U4450 (N_4450,N_2267,N_2399);
and U4451 (N_4451,N_880,N_305);
and U4452 (N_4452,N_3817,N_620);
xnor U4453 (N_4453,N_90,N_974);
and U4454 (N_4454,N_3926,N_2223);
xnor U4455 (N_4455,N_2036,N_1352);
nor U4456 (N_4456,N_1908,N_1888);
xor U4457 (N_4457,N_727,N_3720);
nand U4458 (N_4458,N_384,N_753);
and U4459 (N_4459,N_3053,N_3285);
nor U4460 (N_4460,N_3750,N_3308);
and U4461 (N_4461,N_1328,N_2717);
xnor U4462 (N_4462,N_3030,N_1029);
xnor U4463 (N_4463,N_3857,N_904);
and U4464 (N_4464,N_3581,N_1321);
and U4465 (N_4465,N_3892,N_276);
or U4466 (N_4466,N_887,N_3556);
nand U4467 (N_4467,N_248,N_2638);
and U4468 (N_4468,N_3051,N_1992);
or U4469 (N_4469,N_2087,N_2393);
xnor U4470 (N_4470,N_1142,N_2500);
xor U4471 (N_4471,N_1313,N_3902);
nand U4472 (N_4472,N_2580,N_2975);
nand U4473 (N_4473,N_2373,N_2988);
and U4474 (N_4474,N_1064,N_2491);
nor U4475 (N_4475,N_1834,N_3090);
nand U4476 (N_4476,N_553,N_876);
xor U4477 (N_4477,N_1110,N_471);
xor U4478 (N_4478,N_484,N_3772);
and U4479 (N_4479,N_1042,N_1290);
and U4480 (N_4480,N_382,N_2715);
xor U4481 (N_4481,N_3423,N_3699);
or U4482 (N_4482,N_1858,N_1256);
xnor U4483 (N_4483,N_2260,N_1372);
and U4484 (N_4484,N_1286,N_815);
and U4485 (N_4485,N_1275,N_3769);
nand U4486 (N_4486,N_2569,N_499);
and U4487 (N_4487,N_377,N_1468);
or U4488 (N_4488,N_3684,N_394);
nor U4489 (N_4489,N_3260,N_3224);
nand U4490 (N_4490,N_83,N_2821);
or U4491 (N_4491,N_2166,N_3735);
nor U4492 (N_4492,N_3054,N_1585);
and U4493 (N_4493,N_3589,N_1304);
and U4494 (N_4494,N_3513,N_299);
xnor U4495 (N_4495,N_1841,N_3698);
nor U4496 (N_4496,N_2139,N_773);
and U4497 (N_4497,N_3383,N_681);
xnor U4498 (N_4498,N_3466,N_374);
xnor U4499 (N_4499,N_1493,N_660);
nor U4500 (N_4500,N_1928,N_2039);
nor U4501 (N_4501,N_2639,N_896);
and U4502 (N_4502,N_2619,N_2020);
xnor U4503 (N_4503,N_918,N_2108);
or U4504 (N_4504,N_3951,N_196);
nand U4505 (N_4505,N_3796,N_527);
xor U4506 (N_4506,N_1116,N_1505);
or U4507 (N_4507,N_317,N_985);
and U4508 (N_4508,N_639,N_3277);
or U4509 (N_4509,N_3143,N_791);
nor U4510 (N_4510,N_892,N_2908);
or U4511 (N_4511,N_3864,N_3839);
xor U4512 (N_4512,N_1850,N_2990);
or U4513 (N_4513,N_977,N_1760);
or U4514 (N_4514,N_3558,N_1898);
nand U4515 (N_4515,N_3536,N_551);
or U4516 (N_4516,N_1916,N_2961);
nor U4517 (N_4517,N_3357,N_3116);
or U4518 (N_4518,N_1158,N_191);
or U4519 (N_4519,N_2982,N_2782);
nand U4520 (N_4520,N_473,N_913);
and U4521 (N_4521,N_3202,N_824);
nand U4522 (N_4522,N_134,N_362);
and U4523 (N_4523,N_3866,N_137);
xor U4524 (N_4524,N_497,N_2516);
nand U4525 (N_4525,N_466,N_3578);
nand U4526 (N_4526,N_1229,N_899);
and U4527 (N_4527,N_2857,N_1889);
or U4528 (N_4528,N_3812,N_218);
nand U4529 (N_4529,N_2501,N_2978);
and U4530 (N_4530,N_2707,N_1545);
xor U4531 (N_4531,N_3544,N_3299);
nor U4532 (N_4532,N_2095,N_3977);
nand U4533 (N_4533,N_1638,N_1580);
or U4534 (N_4534,N_3758,N_859);
nor U4535 (N_4535,N_2765,N_1179);
nor U4536 (N_4536,N_735,N_3635);
nand U4537 (N_4537,N_3232,N_1608);
or U4538 (N_4538,N_2256,N_672);
nand U4539 (N_4539,N_1195,N_894);
nor U4540 (N_4540,N_396,N_1187);
and U4541 (N_4541,N_110,N_2644);
xnor U4542 (N_4542,N_1673,N_971);
xnor U4543 (N_4543,N_3336,N_2384);
nor U4544 (N_4544,N_2066,N_872);
or U4545 (N_4545,N_2531,N_1240);
nor U4546 (N_4546,N_2412,N_1636);
and U4547 (N_4547,N_3434,N_3104);
nand U4548 (N_4548,N_2625,N_3321);
or U4549 (N_4549,N_2680,N_3408);
and U4550 (N_4550,N_2135,N_2744);
xnor U4551 (N_4551,N_3626,N_1790);
and U4552 (N_4552,N_3688,N_449);
nand U4553 (N_4553,N_1287,N_33);
xnor U4554 (N_4554,N_1144,N_3320);
and U4555 (N_4555,N_666,N_674);
or U4556 (N_4556,N_25,N_279);
xor U4557 (N_4557,N_996,N_3365);
or U4558 (N_4558,N_2695,N_2142);
or U4559 (N_4559,N_3798,N_3182);
or U4560 (N_4560,N_1604,N_552);
and U4561 (N_4561,N_3940,N_427);
nand U4562 (N_4562,N_1962,N_2871);
nand U4563 (N_4563,N_1937,N_2566);
and U4564 (N_4564,N_243,N_1895);
or U4565 (N_4565,N_935,N_141);
nor U4566 (N_4566,N_954,N_3362);
nor U4567 (N_4567,N_3677,N_1672);
nor U4568 (N_4568,N_715,N_76);
nor U4569 (N_4569,N_3615,N_3831);
nor U4570 (N_4570,N_1855,N_1387);
nor U4571 (N_4571,N_3492,N_2302);
nor U4572 (N_4572,N_2409,N_1699);
nand U4573 (N_4573,N_3341,N_2794);
nand U4574 (N_4574,N_1483,N_2034);
nor U4575 (N_4575,N_2297,N_2793);
nor U4576 (N_4576,N_295,N_347);
nand U4577 (N_4577,N_1573,N_1961);
xor U4578 (N_4578,N_829,N_823);
and U4579 (N_4579,N_2333,N_1289);
nand U4580 (N_4580,N_2774,N_257);
xor U4581 (N_4581,N_494,N_375);
and U4582 (N_4582,N_245,N_1407);
or U4583 (N_4583,N_2613,N_3702);
nand U4584 (N_4584,N_178,N_2562);
xor U4585 (N_4585,N_2930,N_3886);
and U4586 (N_4586,N_1740,N_315);
and U4587 (N_4587,N_131,N_544);
xnor U4588 (N_4588,N_1635,N_2125);
nand U4589 (N_4589,N_309,N_3057);
xor U4590 (N_4590,N_2699,N_745);
and U4591 (N_4591,N_1671,N_3710);
nor U4592 (N_4592,N_3690,N_642);
nor U4593 (N_4593,N_3334,N_3112);
or U4594 (N_4594,N_455,N_333);
xor U4595 (N_4595,N_3634,N_3099);
nand U4596 (N_4596,N_1734,N_2255);
or U4597 (N_4597,N_2688,N_381);
and U4598 (N_4598,N_1020,N_3631);
and U4599 (N_4599,N_646,N_1719);
nor U4600 (N_4600,N_1165,N_2398);
and U4601 (N_4601,N_26,N_3681);
and U4602 (N_4602,N_3749,N_3311);
or U4603 (N_4603,N_258,N_3440);
nand U4604 (N_4604,N_3411,N_2593);
and U4605 (N_4605,N_2366,N_3235);
nand U4606 (N_4606,N_1739,N_2262);
xor U4607 (N_4607,N_842,N_462);
and U4608 (N_4608,N_559,N_3806);
and U4609 (N_4609,N_2807,N_310);
nor U4610 (N_4610,N_3343,N_1049);
nand U4611 (N_4611,N_2461,N_2488);
xnor U4612 (N_4612,N_1751,N_1938);
and U4613 (N_4613,N_1300,N_1859);
nor U4614 (N_4614,N_2515,N_3181);
and U4615 (N_4615,N_2043,N_2670);
nor U4616 (N_4616,N_2261,N_3709);
nand U4617 (N_4617,N_2293,N_640);
xor U4618 (N_4618,N_3444,N_3602);
xor U4619 (N_4619,N_720,N_2740);
or U4620 (N_4620,N_1619,N_2225);
xnor U4621 (N_4621,N_1511,N_3645);
xnor U4622 (N_4622,N_3686,N_1563);
xor U4623 (N_4623,N_669,N_2464);
nor U4624 (N_4624,N_1030,N_2272);
and U4625 (N_4625,N_3861,N_3020);
and U4626 (N_4626,N_1477,N_3306);
xor U4627 (N_4627,N_1239,N_3049);
nor U4628 (N_4628,N_636,N_1278);
nand U4629 (N_4629,N_2627,N_516);
and U4630 (N_4630,N_2864,N_3976);
nand U4631 (N_4631,N_286,N_2315);
nand U4632 (N_4632,N_1528,N_3214);
and U4633 (N_4633,N_1308,N_1854);
and U4634 (N_4634,N_433,N_1358);
nand U4635 (N_4635,N_3882,N_2379);
or U4636 (N_4636,N_3340,N_430);
nor U4637 (N_4637,N_1729,N_1102);
nor U4638 (N_4638,N_283,N_2466);
xor U4639 (N_4639,N_3879,N_1519);
nand U4640 (N_4640,N_1060,N_1226);
nor U4641 (N_4641,N_2338,N_20);
nand U4642 (N_4642,N_378,N_1757);
and U4643 (N_4643,N_1078,N_2468);
or U4644 (N_4644,N_2725,N_1815);
or U4645 (N_4645,N_1630,N_1418);
or U4646 (N_4646,N_2901,N_1720);
xnor U4647 (N_4647,N_1966,N_2080);
or U4648 (N_4648,N_1143,N_3514);
xnor U4649 (N_4649,N_509,N_1623);
nor U4650 (N_4650,N_957,N_1544);
nor U4651 (N_4651,N_2212,N_2457);
or U4652 (N_4652,N_3108,N_1627);
nor U4653 (N_4653,N_1900,N_2673);
nor U4654 (N_4654,N_2956,N_3679);
nor U4655 (N_4655,N_1769,N_765);
and U4656 (N_4656,N_2328,N_3724);
nand U4657 (N_4657,N_1903,N_2484);
and U4658 (N_4658,N_705,N_1201);
xnor U4659 (N_4659,N_737,N_776);
xor U4660 (N_4660,N_3776,N_2953);
and U4661 (N_4661,N_743,N_2072);
nor U4662 (N_4662,N_1191,N_1891);
and U4663 (N_4663,N_2064,N_1479);
and U4664 (N_4664,N_1915,N_2371);
nor U4665 (N_4665,N_1603,N_1283);
and U4666 (N_4666,N_2129,N_434);
or U4667 (N_4667,N_3984,N_630);
and U4668 (N_4668,N_3089,N_2641);
or U4669 (N_4669,N_2202,N_1365);
nand U4670 (N_4670,N_832,N_2116);
nor U4671 (N_4671,N_1596,N_3262);
nor U4672 (N_4672,N_1725,N_2331);
or U4673 (N_4673,N_278,N_189);
nor U4674 (N_4674,N_80,N_572);
and U4675 (N_4675,N_2182,N_1379);
and U4676 (N_4676,N_3086,N_1005);
xor U4677 (N_4677,N_1846,N_817);
and U4678 (N_4678,N_524,N_461);
xor U4679 (N_4679,N_116,N_180);
xor U4680 (N_4680,N_3125,N_2690);
nand U4681 (N_4681,N_1866,N_2510);
nand U4682 (N_4682,N_513,N_3217);
nor U4683 (N_4683,N_3255,N_1118);
xor U4684 (N_4684,N_1396,N_928);
and U4685 (N_4685,N_3654,N_2657);
xor U4686 (N_4686,N_1359,N_1475);
xor U4687 (N_4687,N_2913,N_1032);
nand U4688 (N_4688,N_1339,N_2860);
xnor U4689 (N_4689,N_1822,N_1248);
xor U4690 (N_4690,N_1231,N_3897);
nor U4691 (N_4691,N_939,N_3196);
xnor U4692 (N_4692,N_2777,N_3807);
and U4693 (N_4693,N_1427,N_978);
nor U4694 (N_4694,N_618,N_2697);
and U4695 (N_4695,N_3371,N_1968);
xnor U4696 (N_4696,N_392,N_833);
xnor U4697 (N_4697,N_2356,N_964);
and U4698 (N_4698,N_2927,N_3657);
or U4699 (N_4699,N_1376,N_1171);
nor U4700 (N_4700,N_1668,N_2661);
and U4701 (N_4701,N_3511,N_2345);
and U4702 (N_4702,N_3059,N_2181);
or U4703 (N_4703,N_306,N_755);
nand U4704 (N_4704,N_1099,N_3160);
xnor U4705 (N_4705,N_3388,N_1085);
nand U4706 (N_4706,N_1073,N_786);
nand U4707 (N_4707,N_2312,N_3356);
and U4708 (N_4708,N_1625,N_337);
nor U4709 (N_4709,N_470,N_1667);
nand U4710 (N_4710,N_1873,N_1612);
and U4711 (N_4711,N_631,N_3510);
xor U4712 (N_4712,N_1576,N_2505);
nand U4713 (N_4713,N_539,N_2776);
nand U4714 (N_4714,N_1853,N_2065);
and U4715 (N_4715,N_2131,N_297);
nand U4716 (N_4716,N_3046,N_535);
nand U4717 (N_4717,N_1139,N_1527);
xnor U4718 (N_4718,N_49,N_2868);
nor U4719 (N_4719,N_3253,N_2947);
xnor U4720 (N_4720,N_733,N_42);
or U4721 (N_4721,N_580,N_2422);
xor U4722 (N_4722,N_1211,N_52);
nor U4723 (N_4723,N_3430,N_1467);
and U4724 (N_4724,N_3949,N_650);
nor U4725 (N_4725,N_2246,N_3278);
nor U4726 (N_4726,N_1914,N_2785);
and U4727 (N_4727,N_99,N_1571);
or U4728 (N_4728,N_619,N_2736);
or U4729 (N_4729,N_2544,N_1759);
or U4730 (N_4730,N_3276,N_1128);
nand U4731 (N_4731,N_1205,N_3590);
nand U4732 (N_4732,N_3756,N_3875);
nand U4733 (N_4733,N_2669,N_3413);
or U4734 (N_4734,N_2386,N_407);
nand U4735 (N_4735,N_3888,N_2684);
and U4736 (N_4736,N_1354,N_1081);
nand U4737 (N_4737,N_1065,N_1807);
nor U4738 (N_4738,N_2022,N_1250);
nor U4739 (N_4739,N_2800,N_3474);
nand U4740 (N_4740,N_1722,N_3468);
and U4741 (N_4741,N_2791,N_387);
nor U4742 (N_4742,N_596,N_989);
nor U4743 (N_4743,N_3461,N_1052);
and U4744 (N_4744,N_1103,N_1566);
nand U4745 (N_4745,N_3954,N_1696);
xnor U4746 (N_4746,N_3637,N_1038);
or U4747 (N_4747,N_2152,N_3830);
and U4748 (N_4748,N_2083,N_830);
nand U4749 (N_4749,N_3478,N_3505);
nor U4750 (N_4750,N_3872,N_2573);
and U4751 (N_4751,N_1002,N_3979);
and U4752 (N_4752,N_1330,N_1087);
xnor U4753 (N_4753,N_869,N_2071);
nor U4754 (N_4754,N_1006,N_571);
and U4755 (N_4755,N_3041,N_3432);
or U4756 (N_4756,N_2783,N_2958);
xnor U4757 (N_4757,N_2582,N_354);
or U4758 (N_4758,N_1979,N_418);
or U4759 (N_4759,N_3226,N_3966);
xor U4760 (N_4760,N_3457,N_2092);
and U4761 (N_4761,N_875,N_2423);
and U4762 (N_4762,N_2075,N_2882);
nor U4763 (N_4763,N_3219,N_1374);
xor U4764 (N_4764,N_2843,N_1586);
xor U4765 (N_4765,N_2632,N_2425);
nor U4766 (N_4766,N_2038,N_2959);
or U4767 (N_4767,N_2618,N_2674);
nor U4768 (N_4768,N_280,N_1805);
and U4769 (N_4769,N_1389,N_1465);
nor U4770 (N_4770,N_1057,N_2838);
nor U4771 (N_4771,N_69,N_1438);
nor U4772 (N_4772,N_1382,N_2028);
nand U4773 (N_4773,N_1455,N_2507);
or U4774 (N_4774,N_3991,N_2496);
nand U4775 (N_4775,N_2539,N_1797);
nand U4776 (N_4776,N_901,N_577);
nand U4777 (N_4777,N_2890,N_1001);
nand U4778 (N_4778,N_38,N_718);
or U4779 (N_4779,N_615,N_3658);
and U4780 (N_4780,N_3366,N_1600);
nand U4781 (N_4781,N_467,N_2055);
and U4782 (N_4782,N_3115,N_3800);
xor U4783 (N_4783,N_622,N_758);
nor U4784 (N_4784,N_2590,N_3946);
or U4785 (N_4785,N_500,N_1268);
xor U4786 (N_4786,N_532,N_274);
nor U4787 (N_4787,N_1843,N_3743);
nor U4788 (N_4788,N_3069,N_225);
or U4789 (N_4789,N_1324,N_2433);
and U4790 (N_4790,N_3771,N_3990);
and U4791 (N_4791,N_1881,N_219);
nor U4792 (N_4792,N_1249,N_700);
or U4793 (N_4793,N_447,N_105);
and U4794 (N_4794,N_2298,N_282);
nand U4795 (N_4795,N_1670,N_3428);
nand U4796 (N_4796,N_2209,N_2335);
nand U4797 (N_4797,N_1244,N_1839);
and U4798 (N_4798,N_3697,N_3734);
or U4799 (N_4799,N_246,N_3737);
or U4800 (N_4800,N_1314,N_2520);
or U4801 (N_4801,N_2640,N_3091);
and U4802 (N_4802,N_3248,N_895);
xor U4803 (N_4803,N_2251,N_2554);
xnor U4804 (N_4804,N_3789,N_3065);
xnor U4805 (N_4805,N_3034,N_621);
and U4806 (N_4806,N_1082,N_2991);
nand U4807 (N_4807,N_3713,N_2085);
xnor U4808 (N_4808,N_2560,N_2485);
or U4809 (N_4809,N_66,N_2921);
or U4810 (N_4810,N_2449,N_582);
xnor U4811 (N_4811,N_2599,N_844);
nand U4812 (N_4812,N_706,N_2348);
xor U4813 (N_4813,N_429,N_2400);
nand U4814 (N_4814,N_1728,N_2896);
nor U4815 (N_4815,N_2430,N_3135);
nand U4816 (N_4816,N_1849,N_1327);
nand U4817 (N_4817,N_1325,N_1174);
nand U4818 (N_4818,N_1693,N_3774);
xnor U4819 (N_4819,N_3727,N_1485);
nand U4820 (N_4820,N_3103,N_112);
nor U4821 (N_4821,N_2102,N_1093);
and U4822 (N_4822,N_2040,N_2185);
xnor U4823 (N_4823,N_2624,N_35);
and U4824 (N_4824,N_3553,N_3267);
nor U4825 (N_4825,N_3992,N_2026);
xnor U4826 (N_4826,N_3562,N_3820);
xnor U4827 (N_4827,N_2561,N_2893);
xor U4828 (N_4828,N_611,N_2626);
nor U4829 (N_4829,N_2437,N_3426);
and U4830 (N_4830,N_521,N_2149);
nand U4831 (N_4831,N_2007,N_1203);
nor U4832 (N_4832,N_1486,N_3176);
xor U4833 (N_4833,N_1809,N_3400);
xnor U4834 (N_4834,N_2773,N_3777);
xor U4835 (N_4835,N_63,N_772);
and U4836 (N_4836,N_2242,N_3925);
nor U4837 (N_4837,N_868,N_856);
nor U4838 (N_4838,N_3944,N_3752);
and U4839 (N_4839,N_2899,N_2218);
or U4840 (N_4840,N_1905,N_655);
xor U4841 (N_4841,N_1280,N_1055);
or U4842 (N_4842,N_2743,N_2165);
nand U4843 (N_4843,N_649,N_3726);
nand U4844 (N_4844,N_217,N_1795);
nor U4845 (N_4845,N_1735,N_2658);
xnor U4846 (N_4846,N_3762,N_614);
nand U4847 (N_4847,N_3858,N_2067);
xnor U4848 (N_4848,N_1133,N_3700);
or U4849 (N_4849,N_1942,N_1183);
and U4850 (N_4850,N_2737,N_3670);
xnor U4851 (N_4851,N_1257,N_2647);
nand U4852 (N_4852,N_2228,N_1218);
or U4853 (N_4853,N_460,N_3031);
and U4854 (N_4854,N_1422,N_1247);
nor U4855 (N_4855,N_2924,N_3564);
and U4856 (N_4856,N_3210,N_2895);
nor U4857 (N_4857,N_889,N_1351);
and U4858 (N_4858,N_716,N_1217);
or U4859 (N_4859,N_3644,N_269);
or U4860 (N_4860,N_2458,N_3997);
or U4861 (N_4861,N_3372,N_696);
nand U4862 (N_4862,N_1301,N_388);
nor U4863 (N_4863,N_3612,N_638);
nand U4864 (N_4864,N_2758,N_506);
nand U4865 (N_4865,N_2025,N_623);
nand U4866 (N_4866,N_2000,N_3620);
and U4867 (N_4867,N_3901,N_202);
or U4868 (N_4868,N_2431,N_1491);
nor U4869 (N_4869,N_1119,N_1448);
and U4870 (N_4870,N_2200,N_3927);
and U4871 (N_4871,N_3923,N_714);
xor U4872 (N_4872,N_2967,N_1733);
nor U4873 (N_4873,N_1857,N_955);
and U4874 (N_4874,N_456,N_2681);
nand U4875 (N_4875,N_4,N_1007);
and U4876 (N_4876,N_1322,N_1076);
and U4877 (N_4877,N_806,N_2716);
xor U4878 (N_4878,N_2134,N_3237);
xor U4879 (N_4879,N_3142,N_2888);
nand U4880 (N_4880,N_1616,N_2667);
and U4881 (N_4881,N_1660,N_2509);
or U4882 (N_4882,N_2114,N_1958);
xnor U4883 (N_4883,N_3484,N_1800);
nand U4884 (N_4884,N_209,N_3106);
nand U4885 (N_4885,N_3449,N_821);
xnor U4886 (N_4886,N_3676,N_2727);
xnor U4887 (N_4887,N_742,N_3941);
nand U4888 (N_4888,N_1160,N_3096);
xor U4889 (N_4889,N_1262,N_533);
nand U4890 (N_4890,N_1810,N_1084);
xnor U4891 (N_4891,N_1381,N_2902);
xnor U4892 (N_4892,N_97,N_1646);
nand U4893 (N_4893,N_1056,N_19);
xnor U4894 (N_4894,N_610,N_221);
nand U4895 (N_4895,N_2054,N_2494);
nand U4896 (N_4896,N_2350,N_1504);
nor U4897 (N_4897,N_3019,N_652);
nand U4898 (N_4898,N_2850,N_2263);
or U4899 (N_4899,N_3733,N_2678);
or U4900 (N_4900,N_2111,N_827);
nand U4901 (N_4901,N_3291,N_3171);
nand U4902 (N_4902,N_3393,N_3646);
or U4903 (N_4903,N_207,N_547);
and U4904 (N_4904,N_1312,N_583);
and U4905 (N_4905,N_841,N_810);
or U4906 (N_4906,N_2578,N_2051);
nand U4907 (N_4907,N_1192,N_934);
nand U4908 (N_4908,N_2521,N_3155);
nor U4909 (N_4909,N_1063,N_3445);
xor U4910 (N_4910,N_2911,N_1851);
and U4911 (N_4911,N_2570,N_341);
or U4912 (N_4912,N_3480,N_3223);
nor U4913 (N_4913,N_1923,N_1579);
nand U4914 (N_4914,N_1907,N_3828);
and U4915 (N_4915,N_603,N_898);
xor U4916 (N_4916,N_2008,N_3822);
nand U4917 (N_4917,N_3824,N_2339);
nor U4918 (N_4918,N_1109,N_242);
xnor U4919 (N_4919,N_2478,N_21);
xor U4920 (N_4920,N_3996,N_3668);
nand U4921 (N_4921,N_325,N_2565);
xnor U4922 (N_4922,N_3319,N_3367);
or U4923 (N_4923,N_117,N_1803);
xnor U4924 (N_4924,N_808,N_3395);
xnor U4925 (N_4925,N_641,N_468);
and U4926 (N_4926,N_942,N_254);
xor U4927 (N_4927,N_27,N_3711);
xnor U4928 (N_4928,N_3844,N_1631);
and U4929 (N_4929,N_3072,N_2568);
nor U4930 (N_4930,N_224,N_2668);
nor U4931 (N_4931,N_2191,N_2604);
or U4932 (N_4932,N_2286,N_878);
or U4933 (N_4933,N_28,N_1193);
and U4934 (N_4934,N_2919,N_329);
nand U4935 (N_4935,N_2996,N_3123);
and U4936 (N_4936,N_947,N_1620);
or U4937 (N_4937,N_3082,N_2377);
nand U4938 (N_4938,N_3799,N_253);
nor U4939 (N_4939,N_266,N_2759);
nor U4940 (N_4940,N_3271,N_301);
nor U4941 (N_4941,N_2946,N_3649);
or U4942 (N_4942,N_1977,N_463);
and U4943 (N_4943,N_1595,N_3722);
nand U4944 (N_4944,N_944,N_3766);
nand U4945 (N_4945,N_156,N_3716);
xor U4946 (N_4946,N_3290,N_1657);
or U4947 (N_4947,N_1621,N_3519);
xnor U4948 (N_4948,N_3080,N_999);
nor U4949 (N_4949,N_138,N_226);
xnor U4950 (N_4950,N_2750,N_503);
and U4951 (N_4951,N_2698,N_3095);
xor U4952 (N_4952,N_1536,N_1369);
or U4953 (N_4953,N_2522,N_2664);
and U4954 (N_4954,N_1860,N_858);
and U4955 (N_4955,N_608,N_662);
or U4956 (N_4956,N_3404,N_428);
xnor U4957 (N_4957,N_2027,N_3874);
nor U4958 (N_4958,N_211,N_3671);
nor U4959 (N_4959,N_3521,N_1601);
xnor U4960 (N_4960,N_1152,N_3382);
xor U4961 (N_4961,N_3840,N_3148);
or U4962 (N_4962,N_3767,N_2918);
or U4963 (N_4963,N_1161,N_814);
nand U4964 (N_4964,N_3584,N_3561);
nor U4965 (N_4965,N_2167,N_1021);
or U4966 (N_4966,N_3242,N_1690);
nor U4967 (N_4967,N_126,N_625);
xor U4968 (N_4968,N_3164,N_3619);
or U4969 (N_4969,N_2952,N_445);
xnor U4970 (N_4970,N_351,N_2939);
and U4971 (N_4971,N_3543,N_442);
and U4972 (N_4972,N_1509,N_1731);
or U4973 (N_4973,N_3349,N_783);
xor U4974 (N_4974,N_3119,N_1819);
or U4975 (N_4975,N_372,N_2155);
or U4976 (N_4976,N_1213,N_3651);
and U4977 (N_4977,N_2691,N_459);
nand U4978 (N_4978,N_327,N_1488);
and U4979 (N_4979,N_597,N_3479);
or U4980 (N_4980,N_2084,N_3185);
nand U4981 (N_4981,N_3410,N_703);
nor U4982 (N_4982,N_1981,N_123);
or U4983 (N_4983,N_3403,N_932);
xor U4984 (N_4984,N_3517,N_3249);
and U4985 (N_4985,N_1077,N_3353);
nor U4986 (N_4986,N_2349,N_907);
nor U4987 (N_4987,N_335,N_1281);
and U4988 (N_4988,N_2577,N_3577);
nand U4989 (N_4989,N_2512,N_3497);
xor U4990 (N_4990,N_628,N_431);
xnor U4991 (N_4991,N_95,N_2631);
nor U4992 (N_4992,N_2859,N_1806);
nand U4993 (N_4993,N_3189,N_2651);
and U4994 (N_4994,N_1791,N_265);
and U4995 (N_4995,N_2672,N_1567);
xnor U4996 (N_4996,N_1973,N_3079);
xnor U4997 (N_4997,N_3728,N_1499);
or U4998 (N_4998,N_3003,N_3597);
and U4999 (N_4999,N_267,N_2844);
nand U5000 (N_5000,N_2995,N_2158);
nand U5001 (N_5001,N_2105,N_1875);
nor U5002 (N_5002,N_3130,N_2767);
and U5003 (N_5003,N_2352,N_3856);
nor U5004 (N_5004,N_1793,N_3813);
or U5005 (N_5005,N_2239,N_2002);
or U5006 (N_5006,N_1258,N_1259);
nand U5007 (N_5007,N_132,N_1976);
nor U5008 (N_5008,N_602,N_1825);
xnor U5009 (N_5009,N_825,N_670);
xnor U5010 (N_5010,N_1738,N_2001);
nand U5011 (N_5011,N_296,N_464);
xnor U5012 (N_5012,N_3786,N_637);
xor U5013 (N_5013,N_1716,N_331);
xor U5014 (N_5014,N_2506,N_2275);
or U5015 (N_5015,N_1264,N_1515);
and U5016 (N_5016,N_3541,N_3489);
nand U5017 (N_5017,N_688,N_2689);
nand U5018 (N_5018,N_124,N_1692);
xor U5019 (N_5019,N_2305,N_320);
xnor U5020 (N_5020,N_2880,N_3048);
nand U5021 (N_5021,N_2656,N_2645);
nor U5022 (N_5022,N_1238,N_1610);
xor U5023 (N_5023,N_982,N_948);
and U5024 (N_5024,N_593,N_187);
and U5025 (N_5025,N_2362,N_3981);
xnor U5026 (N_5026,N_2811,N_3006);
xor U5027 (N_5027,N_3583,N_3552);
nor U5028 (N_5028,N_3422,N_2372);
or U5029 (N_5029,N_2492,N_3896);
nor U5030 (N_5030,N_2780,N_2948);
or U5031 (N_5031,N_2462,N_993);
and U5032 (N_5032,N_1882,N_1708);
or U5033 (N_5033,N_1034,N_1628);
xnor U5034 (N_5034,N_120,N_1814);
nand U5035 (N_5035,N_2394,N_3193);
nand U5036 (N_5036,N_3488,N_408);
xnor U5037 (N_5037,N_3199,N_3794);
xor U5038 (N_5038,N_2803,N_1307);
nor U5039 (N_5039,N_1316,N_2254);
nand U5040 (N_5040,N_1529,N_1582);
xor U5041 (N_5041,N_3254,N_3345);
nor U5042 (N_5042,N_208,N_2053);
and U5043 (N_5043,N_3904,N_3847);
xor U5044 (N_5044,N_1556,N_2665);
xnor U5045 (N_5045,N_3167,N_364);
or U5046 (N_5046,N_405,N_3348);
xnor U5047 (N_5047,N_3691,N_2876);
nor U5048 (N_5048,N_2594,N_3501);
and U5049 (N_5049,N_1019,N_710);
and U5050 (N_5050,N_920,N_3506);
nand U5051 (N_5051,N_1540,N_520);
nor U5052 (N_5052,N_1282,N_1774);
or U5053 (N_5053,N_2221,N_3810);
xnor U5054 (N_5054,N_1997,N_360);
and U5055 (N_5055,N_1637,N_1959);
nor U5056 (N_5056,N_2137,N_984);
xnor U5057 (N_5057,N_3659,N_3446);
xnor U5058 (N_5058,N_2756,N_665);
xnor U5059 (N_5059,N_1310,N_232);
and U5060 (N_5060,N_3660,N_2003);
nand U5061 (N_5061,N_3986,N_1742);
and U5062 (N_5062,N_3360,N_1112);
and U5063 (N_5063,N_683,N_2211);
or U5064 (N_5064,N_1827,N_1452);
and U5065 (N_5065,N_3775,N_2849);
and U5066 (N_5066,N_2391,N_2323);
xnor U5067 (N_5067,N_1198,N_67);
xor U5068 (N_5068,N_3533,N_3804);
xnor U5069 (N_5069,N_2472,N_1870);
nor U5070 (N_5070,N_3673,N_861);
and U5071 (N_5071,N_1999,N_2528);
xor U5072 (N_5072,N_3653,N_440);
or U5073 (N_5073,N_79,N_2397);
or U5074 (N_5074,N_1302,N_2989);
nand U5075 (N_5075,N_3361,N_1400);
and U5076 (N_5076,N_3012,N_1086);
nor U5077 (N_5077,N_2718,N_1705);
nor U5078 (N_5078,N_2490,N_2477);
and U5079 (N_5079,N_557,N_877);
or U5080 (N_5080,N_2954,N_1597);
and U5081 (N_5081,N_2281,N_3746);
and U5082 (N_5082,N_3159,N_1876);
or U5083 (N_5083,N_1252,N_3389);
nor U5084 (N_5084,N_2608,N_2787);
xor U5085 (N_5085,N_2188,N_3376);
nor U5086 (N_5086,N_2945,N_1170);
xnor U5087 (N_5087,N_590,N_864);
nor U5088 (N_5088,N_2596,N_1206);
xor U5089 (N_5089,N_568,N_3633);
nor U5090 (N_5090,N_2693,N_940);
nor U5091 (N_5091,N_53,N_3391);
nand U5092 (N_5092,N_3067,N_271);
nand U5093 (N_5093,N_1415,N_96);
nor U5094 (N_5094,N_3630,N_3745);
and U5095 (N_5095,N_2163,N_1474);
nor U5096 (N_5096,N_3569,N_3016);
and U5097 (N_5097,N_453,N_1131);
nor U5098 (N_5098,N_3292,N_531);
nand U5099 (N_5099,N_1987,N_2489);
and U5100 (N_5100,N_402,N_2855);
and U5101 (N_5101,N_3554,N_457);
nand U5102 (N_5102,N_912,N_3101);
or U5103 (N_5103,N_1454,N_585);
and U5104 (N_5104,N_1677,N_951);
or U5105 (N_5105,N_1818,N_3971);
nor U5106 (N_5106,N_2314,N_1047);
nand U5107 (N_5107,N_2745,N_981);
and U5108 (N_5108,N_1364,N_591);
nand U5109 (N_5109,N_2830,N_1678);
nor U5110 (N_5110,N_3988,N_1184);
and U5111 (N_5111,N_2175,N_3177);
nand U5112 (N_5112,N_770,N_3344);
nor U5113 (N_5113,N_2514,N_486);
nor U5114 (N_5114,N_3392,N_2342);
or U5115 (N_5115,N_1902,N_1945);
and U5116 (N_5116,N_2922,N_648);
or U5117 (N_5117,N_122,N_2932);
xor U5118 (N_5118,N_3373,N_2060);
nand U5119 (N_5119,N_545,N_2964);
nor U5120 (N_5120,N_2176,N_2591);
and U5121 (N_5121,N_2546,N_1373);
nor U5122 (N_5122,N_750,N_3593);
xnor U5123 (N_5123,N_2754,N_2016);
xor U5124 (N_5124,N_1663,N_3141);
and U5125 (N_5125,N_3598,N_587);
and U5126 (N_5126,N_2931,N_3161);
nand U5127 (N_5127,N_321,N_1847);
nand U5128 (N_5128,N_1970,N_1089);
nand U5129 (N_5129,N_3370,N_3778);
nor U5130 (N_5130,N_2592,N_1633);
xnor U5131 (N_5131,N_2519,N_828);
xnor U5132 (N_5132,N_1426,N_2826);
and U5133 (N_5133,N_3460,N_690);
nor U5134 (N_5134,N_3421,N_436);
nor U5135 (N_5135,N_393,N_1456);
xnor U5136 (N_5136,N_1377,N_37);
xor U5137 (N_5137,N_1018,N_3021);
nor U5138 (N_5138,N_3729,N_2172);
xnor U5139 (N_5139,N_962,N_2848);
nor U5140 (N_5140,N_3802,N_2401);
nand U5141 (N_5141,N_1632,N_616);
and U5142 (N_5142,N_2571,N_3209);
nand U5143 (N_5143,N_2585,N_3231);
xnor U5144 (N_5144,N_1925,N_1639);
and U5145 (N_5145,N_3907,N_1695);
or U5146 (N_5146,N_2659,N_992);
or U5147 (N_5147,N_1546,N_3815);
nand U5148 (N_5148,N_1951,N_1513);
nand U5149 (N_5149,N_158,N_1177);
and U5150 (N_5150,N_1655,N_1930);
nor U5151 (N_5151,N_914,N_785);
or U5152 (N_5152,N_1482,N_3227);
and U5153 (N_5153,N_908,N_2746);
xnor U5154 (N_5154,N_1041,N_32);
and U5155 (N_5155,N_1764,N_1096);
nor U5156 (N_5156,N_1517,N_3314);
nor U5157 (N_5157,N_152,N_3056);
or U5158 (N_5158,N_702,N_2283);
xnor U5159 (N_5159,N_1589,N_149);
nand U5160 (N_5160,N_3149,N_385);
xor U5161 (N_5161,N_3201,N_293);
nand U5162 (N_5162,N_109,N_1451);
xnor U5163 (N_5163,N_2834,N_3281);
and U5164 (N_5164,N_3499,N_147);
and U5165 (N_5165,N_1413,N_1366);
or U5166 (N_5166,N_1512,N_2726);
nor U5167 (N_5167,N_855,N_3689);
xor U5168 (N_5168,N_2470,N_2903);
xor U5169 (N_5169,N_1572,N_2033);
nand U5170 (N_5170,N_2909,N_1885);
or U5171 (N_5171,N_1408,N_3880);
xor U5172 (N_5172,N_1291,N_2183);
and U5173 (N_5173,N_3084,N_1127);
or U5174 (N_5174,N_3117,N_1235);
nor U5175 (N_5175,N_34,N_2307);
nand U5176 (N_5176,N_425,N_1939);
and U5177 (N_5177,N_3957,N_2643);
and U5178 (N_5178,N_3405,N_3687);
or U5179 (N_5179,N_3397,N_834);
and U5180 (N_5180,N_2696,N_3905);
and U5181 (N_5181,N_262,N_1496);
and U5182 (N_5182,N_314,N_3695);
nor U5183 (N_5183,N_2524,N_1886);
nor U5184 (N_5184,N_3947,N_1927);
and U5185 (N_5185,N_2636,N_426);
nand U5186 (N_5186,N_911,N_2622);
and U5187 (N_5187,N_2309,N_119);
and U5188 (N_5188,N_2189,N_1457);
nor U5189 (N_5189,N_3867,N_1221);
nor U5190 (N_5190,N_1481,N_1222);
or U5191 (N_5191,N_708,N_3105);
and U5192 (N_5192,N_2556,N_3937);
and U5193 (N_5193,N_3785,N_1384);
and U5194 (N_5194,N_1883,N_2721);
or U5195 (N_5195,N_3163,N_1934);
xnor U5196 (N_5196,N_973,N_3714);
nand U5197 (N_5197,N_1236,N_1320);
nor U5198 (N_5198,N_719,N_888);
and U5199 (N_5199,N_3929,N_18);
nand U5200 (N_5200,N_1155,N_1260);
nand U5201 (N_5201,N_496,N_3409);
nand U5202 (N_5202,N_3487,N_2847);
nor U5203 (N_5203,N_2548,N_1253);
or U5204 (N_5204,N_1872,N_216);
xor U5205 (N_5205,N_3917,N_2708);
and U5206 (N_5206,N_746,N_1574);
and U5207 (N_5207,N_697,N_201);
or U5208 (N_5208,N_1972,N_3662);
nand U5209 (N_5209,N_1978,N_2981);
nor U5210 (N_5210,N_125,N_1766);
and U5211 (N_5211,N_836,N_2441);
or U5212 (N_5212,N_2438,N_3238);
and U5213 (N_5213,N_3437,N_85);
xor U5214 (N_5214,N_1088,N_3482);
or U5215 (N_5215,N_801,N_2671);
or U5216 (N_5216,N_1402,N_923);
and U5217 (N_5217,N_1156,N_2232);
xor U5218 (N_5218,N_514,N_56);
and U5219 (N_5219,N_843,N_1862);
and U5220 (N_5220,N_663,N_3396);
nand U5221 (N_5221,N_77,N_1624);
nand U5222 (N_5222,N_1753,N_3256);
nor U5223 (N_5223,N_406,N_1059);
and U5224 (N_5224,N_3075,N_1508);
or U5225 (N_5225,N_1094,N_2481);
or U5226 (N_5226,N_732,N_946);
nor U5227 (N_5227,N_687,N_3736);
or U5228 (N_5228,N_2467,N_800);
or U5229 (N_5229,N_2865,N_2184);
nor U5230 (N_5230,N_1749,N_3814);
and U5231 (N_5231,N_3024,N_3009);
nor U5232 (N_5232,N_43,N_1770);
or U5233 (N_5233,N_2050,N_1113);
nor U5234 (N_5234,N_2503,N_2920);
nand U5235 (N_5235,N_1115,N_3062);
xnor U5236 (N_5236,N_2257,N_2081);
nor U5237 (N_5237,N_3833,N_3184);
xor U5238 (N_5238,N_487,N_1921);
and U5239 (N_5239,N_3563,N_748);
or U5240 (N_5240,N_3265,N_3418);
or U5241 (N_5241,N_768,N_2885);
xor U5242 (N_5242,N_2606,N_1948);
or U5243 (N_5243,N_2190,N_2966);
nand U5244 (N_5244,N_73,N_949);
nor U5245 (N_5245,N_1404,N_3244);
or U5246 (N_5246,N_3420,N_2452);
and U5247 (N_5247,N_1104,N_3891);
xor U5248 (N_5248,N_2630,N_1762);
and U5249 (N_5249,N_3624,N_3077);
nor U5250 (N_5250,N_1911,N_2677);
nand U5251 (N_5251,N_3993,N_3832);
nand U5252 (N_5252,N_1309,N_802);
and U5253 (N_5253,N_1227,N_233);
nand U5254 (N_5254,N_2925,N_528);
xnor U5255 (N_5255,N_2250,N_2813);
nor U5256 (N_5256,N_3495,N_1472);
and U5257 (N_5257,N_2417,N_2162);
xnor U5258 (N_5258,N_3692,N_1267);
xnor U5259 (N_5259,N_2179,N_2709);
and U5260 (N_5260,N_40,N_1899);
and U5261 (N_5261,N_926,N_902);
nand U5262 (N_5262,N_2730,N_1909);
and U5263 (N_5263,N_540,N_565);
xnor U5264 (N_5264,N_903,N_3146);
xor U5265 (N_5265,N_3098,N_3241);
nor U5266 (N_5266,N_2551,N_3043);
or U5267 (N_5267,N_2160,N_3070);
or U5268 (N_5268,N_2856,N_2907);
nand U5269 (N_5269,N_1157,N_2310);
and U5270 (N_5270,N_1954,N_2414);
nand U5271 (N_5271,N_2735,N_2301);
nor U5272 (N_5272,N_1050,N_1233);
nor U5273 (N_5273,N_163,N_2023);
xnor U5274 (N_5274,N_113,N_546);
and U5275 (N_5275,N_3502,N_643);
and U5276 (N_5276,N_3066,N_3871);
and U5277 (N_5277,N_290,N_68);
nand U5278 (N_5278,N_1411,N_2687);
nor U5279 (N_5279,N_3129,N_3354);
xnor U5280 (N_5280,N_1659,N_3565);
nand U5281 (N_5281,N_1450,N_2274);
and U5282 (N_5282,N_2471,N_479);
nand U5283 (N_5283,N_2124,N_2614);
xnor U5284 (N_5284,N_3738,N_203);
xnor U5285 (N_5285,N_2361,N_2532);
xor U5286 (N_5286,N_1982,N_3918);
or U5287 (N_5287,N_798,N_3509);
and U5288 (N_5288,N_3317,N_1200);
nand U5289 (N_5289,N_2365,N_2005);
nand U5290 (N_5290,N_2099,N_534);
nor U5291 (N_5291,N_373,N_1090);
nand U5292 (N_5292,N_111,N_3327);
nand U5293 (N_5293,N_417,N_17);
xor U5294 (N_5294,N_2533,N_2617);
nor U5295 (N_5295,N_91,N_515);
xor U5296 (N_5296,N_2536,N_1931);
and U5297 (N_5297,N_3534,N_2595);
and U5298 (N_5298,N_1130,N_2418);
nor U5299 (N_5299,N_3068,N_1775);
nand U5300 (N_5300,N_3851,N_3369);
nand U5301 (N_5301,N_3381,N_2724);
xnor U5302 (N_5302,N_3566,N_2123);
xor U5303 (N_5303,N_2867,N_469);
xor U5304 (N_5304,N_3273,N_1329);
xnor U5305 (N_5305,N_1836,N_3289);
xor U5306 (N_5306,N_657,N_3252);
or U5307 (N_5307,N_929,N_3576);
and U5308 (N_5308,N_1550,N_1823);
nand U5309 (N_5309,N_3998,N_2097);
nand U5310 (N_5310,N_3394,N_192);
nand U5311 (N_5311,N_31,N_29);
or U5312 (N_5312,N_2540,N_925);
nand U5313 (N_5313,N_3318,N_1539);
nand U5314 (N_5314,N_1072,N_2972);
nor U5315 (N_5315,N_759,N_788);
xor U5316 (N_5316,N_2215,N_1225);
nand U5317 (N_5317,N_933,N_1535);
nor U5318 (N_5318,N_2245,N_3790);
or U5319 (N_5319,N_1723,N_1613);
nand U5320 (N_5320,N_1523,N_3915);
nor U5321 (N_5321,N_893,N_1027);
or U5322 (N_5322,N_2168,N_2792);
nor U5323 (N_5323,N_2610,N_1487);
nand U5324 (N_5324,N_2143,N_3433);
or U5325 (N_5325,N_1008,N_155);
or U5326 (N_5326,N_2795,N_1780);
nor U5327 (N_5327,N_2291,N_1777);
and U5328 (N_5328,N_3450,N_677);
nand U5329 (N_5329,N_1458,N_2278);
and U5330 (N_5330,N_1040,N_2199);
or U5331 (N_5331,N_264,N_796);
xor U5332 (N_5332,N_2910,N_2998);
and U5333 (N_5333,N_3580,N_3153);
and U5334 (N_5334,N_1214,N_3782);
and U5335 (N_5335,N_3191,N_1296);
or U5336 (N_5336,N_3038,N_3846);
or U5337 (N_5337,N_2823,N_2156);
or U5338 (N_5338,N_2044,N_3042);
xnor U5339 (N_5339,N_3890,N_199);
and U5340 (N_5340,N_2104,N_3100);
nand U5341 (N_5341,N_1430,N_115);
xor U5342 (N_5342,N_3994,N_840);
and U5343 (N_5343,N_1592,N_2714);
or U5344 (N_5344,N_2161,N_779);
or U5345 (N_5345,N_2233,N_632);
xor U5346 (N_5346,N_2518,N_2047);
nand U5347 (N_5347,N_3133,N_3132);
nand U5348 (N_5348,N_2801,N_2609);
and U5349 (N_5349,N_82,N_2133);
nand U5350 (N_5350,N_2704,N_93);
nor U5351 (N_5351,N_3037,N_1420);
and U5352 (N_5352,N_3795,N_3385);
and U5353 (N_5353,N_2113,N_2363);
and U5354 (N_5354,N_1340,N_905);
or U5355 (N_5355,N_104,N_3494);
xor U5356 (N_5356,N_495,N_391);
xor U5357 (N_5357,N_3452,N_3447);
or U5358 (N_5358,N_3076,N_3282);
xor U5359 (N_5359,N_667,N_54);
and U5360 (N_5360,N_353,N_1111);
and U5361 (N_5361,N_3974,N_316);
nor U5362 (N_5362,N_3740,N_1912);
xor U5363 (N_5363,N_2329,N_3845);
and U5364 (N_5364,N_1036,N_541);
and U5365 (N_5365,N_3324,N_2187);
nor U5366 (N_5366,N_1887,N_1714);
xnor U5367 (N_5367,N_1417,N_1212);
or U5368 (N_5368,N_3887,N_2287);
nand U5369 (N_5369,N_2628,N_3780);
xnor U5370 (N_5370,N_2545,N_3351);
nand U5371 (N_5371,N_3784,N_1263);
nor U5372 (N_5372,N_6,N_330);
xor U5373 (N_5373,N_867,N_576);
xnor U5374 (N_5374,N_2197,N_1590);
nand U5375 (N_5375,N_1129,N_675);
nand U5376 (N_5376,N_204,N_319);
nor U5377 (N_5377,N_332,N_644);
or U5378 (N_5378,N_441,N_2367);
and U5379 (N_5379,N_2243,N_1615);
nand U5380 (N_5380,N_3296,N_846);
nand U5381 (N_5381,N_135,N_1687);
xnor U5382 (N_5382,N_1391,N_2013);
xor U5383 (N_5383,N_968,N_2141);
nor U5384 (N_5384,N_2207,N_2869);
or U5385 (N_5385,N_2076,N_2663);
nand U5386 (N_5386,N_970,N_3187);
nor U5387 (N_5387,N_2705,N_2581);
nor U5388 (N_5388,N_1469,N_3682);
or U5389 (N_5389,N_1584,N_3683);
nand U5390 (N_5390,N_313,N_1215);
nor U5391 (N_5391,N_2118,N_230);
nand U5392 (N_5392,N_2720,N_529);
or U5393 (N_5393,N_2706,N_2983);
or U5394 (N_5394,N_2682,N_530);
nor U5395 (N_5395,N_3342,N_1952);
and U5396 (N_5396,N_3102,N_1463);
nand U5397 (N_5397,N_1242,N_1848);
nand U5398 (N_5398,N_3378,N_3518);
and U5399 (N_5399,N_835,N_1209);
nor U5400 (N_5400,N_822,N_633);
xor U5401 (N_5401,N_2240,N_2006);
or U5402 (N_5402,N_3064,N_3081);
and U5403 (N_5403,N_1514,N_952);
and U5404 (N_5404,N_2247,N_2940);
or U5405 (N_5405,N_1297,N_1917);
nor U5406 (N_5406,N_2388,N_2453);
nor U5407 (N_5407,N_2171,N_3708);
nor U5408 (N_5408,N_437,N_2482);
nor U5409 (N_5409,N_1763,N_1965);
or U5410 (N_5410,N_3567,N_3496);
or U5411 (N_5411,N_1737,N_1394);
xnor U5412 (N_5412,N_693,N_2334);
or U5413 (N_5413,N_1647,N_2413);
nor U5414 (N_5414,N_2205,N_2282);
and U5415 (N_5415,N_423,N_318);
nand U5416 (N_5416,N_2062,N_2957);
nand U5417 (N_5417,N_723,N_2815);
and U5418 (N_5418,N_439,N_2077);
nor U5419 (N_5419,N_2213,N_2059);
nand U5420 (N_5420,N_3528,N_2552);
and U5421 (N_5421,N_3809,N_837);
nand U5422 (N_5422,N_1552,N_2229);
nand U5423 (N_5423,N_778,N_3026);
nor U5424 (N_5424,N_1176,N_2049);
xnor U5425 (N_5425,N_3025,N_3458);
and U5426 (N_5426,N_2186,N_2912);
nand U5427 (N_5427,N_2231,N_3938);
xnor U5428 (N_5428,N_2906,N_2068);
nor U5429 (N_5429,N_2886,N_3850);
nor U5430 (N_5430,N_645,N_2752);
or U5431 (N_5431,N_1447,N_2322);
nand U5432 (N_5432,N_2276,N_1626);
xor U5433 (N_5433,N_1745,N_3573);
xor U5434 (N_5434,N_1591,N_1303);
or U5435 (N_5435,N_1216,N_782);
or U5436 (N_5436,N_976,N_1926);
or U5437 (N_5437,N_3469,N_2999);
xor U5438 (N_5438,N_599,N_3350);
or U5439 (N_5439,N_1706,N_1993);
nand U5440 (N_5440,N_924,N_1832);
and U5441 (N_5441,N_839,N_2583);
nor U5442 (N_5442,N_1553,N_2722);
xnor U5443 (N_5443,N_14,N_975);
xnor U5444 (N_5444,N_3002,N_1985);
or U5445 (N_5445,N_1879,N_969);
and U5446 (N_5446,N_2738,N_194);
nand U5447 (N_5447,N_2648,N_1164);
and U5448 (N_5448,N_937,N_3570);
nand U5449 (N_5449,N_1674,N_87);
xor U5450 (N_5450,N_2021,N_240);
and U5451 (N_5451,N_41,N_1575);
and U5452 (N_5452,N_1868,N_1401);
or U5453 (N_5453,N_3122,N_3178);
and U5454 (N_5454,N_3301,N_92);
nand U5455 (N_5455,N_3912,N_695);
and U5456 (N_5456,N_3968,N_1549);
or U5457 (N_5457,N_3134,N_3073);
and U5458 (N_5458,N_2031,N_1607);
or U5459 (N_5459,N_1747,N_1390);
nor U5460 (N_5460,N_2808,N_3207);
or U5461 (N_5461,N_3664,N_1147);
nand U5462 (N_5462,N_2122,N_162);
and U5463 (N_5463,N_3126,N_3582);
or U5464 (N_5464,N_3448,N_752);
or U5465 (N_5465,N_363,N_510);
nor U5466 (N_5466,N_2822,N_707);
and U5467 (N_5467,N_2601,N_1924);
or U5468 (N_5468,N_139,N_2442);
or U5469 (N_5469,N_1988,N_2861);
xnor U5470 (N_5470,N_2809,N_1151);
xnor U5471 (N_5471,N_2406,N_2103);
nand U5472 (N_5472,N_2148,N_2024);
nand U5473 (N_5473,N_3860,N_3748);
nor U5474 (N_5474,N_549,N_1856);
nor U5475 (N_5475,N_1349,N_1399);
nor U5476 (N_5476,N_493,N_294);
and U5477 (N_5477,N_1570,N_102);
or U5478 (N_5478,N_2327,N_740);
and U5479 (N_5479,N_3286,N_729);
or U5480 (N_5480,N_2753,N_562);
nor U5481 (N_5481,N_3618,N_1023);
or U5482 (N_5482,N_512,N_2048);
and U5483 (N_5483,N_1436,N_1906);
nor U5484 (N_5484,N_523,N_2082);
nand U5485 (N_5485,N_2602,N_44);
nand U5486 (N_5486,N_3183,N_3540);
nand U5487 (N_5487,N_3712,N_1265);
or U5488 (N_5488,N_1317,N_1106);
or U5489 (N_5489,N_1269,N_1588);
nand U5490 (N_5490,N_1208,N_819);
xnor U5491 (N_5491,N_1919,N_359);
or U5492 (N_5492,N_1869,N_165);
nand U5493 (N_5493,N_1039,N_3607);
nor U5494 (N_5494,N_2728,N_1371);
and U5495 (N_5495,N_214,N_3877);
xnor U5496 (N_5496,N_504,N_885);
nor U5497 (N_5497,N_3316,N_1675);
and U5498 (N_5498,N_1416,N_356);
xor U5499 (N_5499,N_626,N_2936);
nand U5500 (N_5500,N_260,N_133);
xnor U5501 (N_5501,N_519,N_2525);
and U5502 (N_5502,N_3485,N_658);
nand U5503 (N_5503,N_1204,N_3216);
nand U5504 (N_5504,N_3205,N_3731);
nand U5505 (N_5505,N_3040,N_963);
or U5506 (N_5506,N_2407,N_2100);
nand U5507 (N_5507,N_766,N_2277);
xor U5508 (N_5508,N_1996,N_1865);
xnor U5509 (N_5509,N_3855,N_2347);
or U5510 (N_5510,N_1466,N_324);
or U5511 (N_5511,N_2434,N_2637);
nor U5512 (N_5512,N_870,N_2951);
and U5513 (N_5513,N_2396,N_3017);
nor U5514 (N_5514,N_398,N_853);
and U5515 (N_5515,N_3374,N_3220);
or U5516 (N_5516,N_358,N_2266);
xnor U5517 (N_5517,N_3470,N_794);
or U5518 (N_5518,N_1629,N_1991);
or U5519 (N_5519,N_164,N_2879);
xnor U5520 (N_5520,N_2177,N_3380);
xnor U5521 (N_5521,N_3097,N_311);
nor U5522 (N_5522,N_2402,N_2812);
xnor U5523 (N_5523,N_2497,N_3674);
nand U5524 (N_5524,N_2535,N_613);
nand U5525 (N_5525,N_350,N_1124);
or U5526 (N_5526,N_2424,N_1009);
nand U5527 (N_5527,N_1035,N_578);
or U5528 (N_5528,N_2979,N_1315);
nand U5529 (N_5529,N_2891,N_3169);
nand U5530 (N_5530,N_3685,N_3429);
or U5531 (N_5531,N_3835,N_2511);
xnor U5532 (N_5532,N_3018,N_389);
and U5533 (N_5533,N_3718,N_725);
nor U5534 (N_5534,N_2447,N_404);
and U5535 (N_5535,N_2214,N_1701);
xor U5536 (N_5536,N_3704,N_2427);
nand U5537 (N_5537,N_1820,N_3869);
nor U5538 (N_5538,N_691,N_2416);
or U5539 (N_5539,N_1617,N_1246);
xnor U5540 (N_5540,N_3643,N_2711);
nand U5541 (N_5541,N_1343,N_1345);
xnor U5542 (N_5542,N_3694,N_1194);
xnor U5543 (N_5543,N_304,N_1380);
or U5544 (N_5544,N_2502,N_2685);
and U5545 (N_5545,N_2324,N_502);
nor U5546 (N_5546,N_1425,N_3808);
and U5547 (N_5547,N_1136,N_3678);
or U5548 (N_5548,N_1651,N_2249);
and U5549 (N_5549,N_717,N_3140);
or U5550 (N_5550,N_3208,N_2448);
nand U5551 (N_5551,N_3229,N_3170);
xnor U5552 (N_5552,N_1071,N_2984);
nor U5553 (N_5553,N_1341,N_328);
and U5554 (N_5554,N_3131,N_206);
nand U5555 (N_5555,N_2829,N_574);
or U5556 (N_5556,N_1497,N_200);
or U5557 (N_5557,N_2836,N_771);
nand U5558 (N_5558,N_3465,N_3287);
nand U5559 (N_5559,N_1120,N_1986);
nand U5560 (N_5560,N_915,N_153);
nand U5561 (N_5561,N_2061,N_3387);
nand U5562 (N_5562,N_511,N_3920);
and U5563 (N_5563,N_1686,N_3162);
xnor U5564 (N_5564,N_1150,N_2110);
and U5565 (N_5565,N_2508,N_3973);
xor U5566 (N_5566,N_421,N_994);
and U5567 (N_5567,N_272,N_2284);
and U5568 (N_5568,N_1444,N_3168);
and U5569 (N_5569,N_2117,N_1392);
or U5570 (N_5570,N_1782,N_3898);
nor U5571 (N_5571,N_2018,N_2010);
nand U5572 (N_5572,N_2629,N_3754);
and U5573 (N_5573,N_1500,N_3412);
xnor U5574 (N_5574,N_679,N_3157);
xor U5575 (N_5575,N_537,N_2814);
nand U5576 (N_5576,N_2884,N_1471);
or U5577 (N_5577,N_850,N_3883);
or U5578 (N_5578,N_2832,N_606);
xnor U5579 (N_5579,N_774,N_3983);
and U5580 (N_5580,N_3156,N_1957);
nor U5581 (N_5581,N_2866,N_1587);
and U5582 (N_5582,N_3648,N_2710);
nor U5583 (N_5583,N_1003,N_150);
nand U5584 (N_5584,N_3894,N_1713);
xor U5585 (N_5585,N_2914,N_762);
and U5586 (N_5586,N_961,N_2652);
xor U5587 (N_5587,N_2620,N_2030);
and U5588 (N_5588,N_1319,N_1061);
and U5589 (N_5589,N_3551,N_2019);
and U5590 (N_5590,N_2635,N_3911);
nand U5591 (N_5591,N_790,N_1833);
nor U5592 (N_5592,N_1473,N_268);
nor U5593 (N_5593,N_3055,N_2290);
xor U5594 (N_5594,N_1126,N_2650);
nand U5595 (N_5595,N_292,N_1024);
nand U5596 (N_5596,N_3781,N_488);
nand U5597 (N_5597,N_3916,N_340);
or U5598 (N_5598,N_1710,N_1337);
nand U5599 (N_5599,N_1534,N_1149);
xor U5600 (N_5600,N_1335,N_2292);
nand U5601 (N_5601,N_3960,N_3257);
nand U5602 (N_5602,N_1688,N_2093);
nand U5603 (N_5603,N_865,N_3258);
xnor U5604 (N_5604,N_3300,N_1228);
and U5605 (N_5605,N_2203,N_65);
xor U5606 (N_5606,N_897,N_454);
nor U5607 (N_5607,N_101,N_1492);
nor U5608 (N_5608,N_1611,N_1446);
or U5609 (N_5609,N_23,N_3616);
xor U5610 (N_5610,N_1526,N_1271);
and U5611 (N_5611,N_458,N_3239);
nand U5612 (N_5612,N_3956,N_159);
xor U5613 (N_5613,N_3107,N_100);
and U5614 (N_5614,N_1947,N_1476);
xor U5615 (N_5615,N_3215,N_1395);
and U5616 (N_5616,N_2898,N_2465);
nor U5617 (N_5617,N_1974,N_451);
nor U5618 (N_5618,N_1360,N_2969);
nor U5619 (N_5619,N_1685,N_1357);
and U5620 (N_5620,N_2700,N_2004);
nand U5621 (N_5621,N_1397,N_3268);
xnor U5622 (N_5622,N_2091,N_3304);
nand U5623 (N_5623,N_2702,N_3529);
or U5624 (N_5624,N_289,N_747);
or U5625 (N_5625,N_3279,N_2222);
and U5626 (N_5626,N_1830,N_2653);
nand U5627 (N_5627,N_2567,N_183);
xnor U5628 (N_5628,N_2317,N_2917);
or U5629 (N_5629,N_1920,N_1015);
nand U5630 (N_5630,N_179,N_1776);
and U5631 (N_5631,N_2749,N_3027);
xor U5632 (N_5632,N_3625,N_46);
and U5633 (N_5633,N_3263,N_609);
nand U5634 (N_5634,N_261,N_3805);
nand U5635 (N_5635,N_3870,N_2330);
nor U5636 (N_5636,N_3476,N_890);
and U5637 (N_5637,N_2253,N_346);
xor U5638 (N_5638,N_2786,N_3788);
nand U5639 (N_5639,N_307,N_916);
and U5640 (N_5640,N_2325,N_673);
or U5641 (N_5641,N_2194,N_1779);
xnor U5642 (N_5642,N_1062,N_3747);
xor U5643 (N_5643,N_443,N_1871);
or U5644 (N_5644,N_1010,N_1101);
and U5645 (N_5645,N_1202,N_960);
or U5646 (N_5646,N_277,N_678);
nor U5647 (N_5647,N_2553,N_3873);
nor U5648 (N_5648,N_3384,N_2109);
xor U5649 (N_5649,N_612,N_1541);
or U5650 (N_5650,N_3721,N_483);
or U5651 (N_5651,N_1707,N_3935);
xor U5652 (N_5652,N_777,N_3264);
nor U5653 (N_5653,N_2374,N_813);
and U5654 (N_5654,N_249,N_2285);
nand U5655 (N_5655,N_3471,N_2858);
and U5656 (N_5656,N_3139,N_1559);
and U5657 (N_5657,N_3174,N_3427);
and U5658 (N_5658,N_1284,N_542);
and U5659 (N_5659,N_2713,N_3585);
or U5660 (N_5660,N_886,N_1606);
or U5661 (N_5661,N_1163,N_1502);
xnor U5662 (N_5662,N_2294,N_3467);
nand U5663 (N_5663,N_1949,N_2180);
and U5664 (N_5664,N_1114,N_1067);
nand U5665 (N_5665,N_3190,N_1053);
nand U5666 (N_5666,N_2584,N_352);
and U5667 (N_5667,N_3601,N_2817);
xnor U5668 (N_5668,N_792,N_1273);
and U5669 (N_5669,N_1787,N_3375);
nor U5670 (N_5670,N_995,N_1736);
xor U5671 (N_5671,N_3136,N_3269);
xnor U5672 (N_5672,N_215,N_174);
xnor U5673 (N_5673,N_2495,N_414);
nor U5674 (N_5674,N_1532,N_1845);
or U5675 (N_5675,N_1838,N_1385);
nor U5676 (N_5676,N_1058,N_2354);
nor U5677 (N_5677,N_1983,N_882);
xor U5678 (N_5678,N_2473,N_930);
nor U5679 (N_5679,N_298,N_2446);
xnor U5680 (N_5680,N_2381,N_2463);
xnor U5681 (N_5681,N_1288,N_2751);
or U5682 (N_5682,N_3739,N_2887);
nor U5683 (N_5683,N_848,N_2603);
or U5684 (N_5684,N_3029,N_3333);
and U5685 (N_5685,N_2498,N_2878);
nor U5686 (N_5686,N_941,N_1440);
nand U5687 (N_5687,N_1609,N_16);
xor U5688 (N_5688,N_2732,N_936);
xor U5689 (N_5689,N_3023,N_3498);
nand U5690 (N_5690,N_3197,N_1423);
and U5691 (N_5691,N_938,N_555);
and U5692 (N_5692,N_1075,N_3462);
and U5693 (N_5693,N_140,N_1277);
and U5694 (N_5694,N_1506,N_3821);
nand U5695 (N_5695,N_2742,N_1123);
or U5696 (N_5696,N_2572,N_1694);
nor U5697 (N_5697,N_3574,N_2090);
and U5698 (N_5698,N_3490,N_2935);
nand U5699 (N_5699,N_1802,N_3303);
or U5700 (N_5700,N_184,N_2268);
or U5701 (N_5701,N_2403,N_1220);
and U5702 (N_5702,N_482,N_3035);
nand U5703 (N_5703,N_2788,N_1137);
and U5704 (N_5704,N_3913,N_1138);
nor U5705 (N_5705,N_3928,N_2779);
and U5706 (N_5706,N_1421,N_1543);
xnor U5707 (N_5707,N_2755,N_3414);
xnor U5708 (N_5708,N_3560,N_1346);
xor U5709 (N_5709,N_1844,N_826);
or U5710 (N_5710,N_1801,N_2841);
xnor U5711 (N_5711,N_3958,N_698);
nor U5712 (N_5712,N_2926,N_3061);
nor U5713 (N_5713,N_1386,N_797);
nand U5714 (N_5714,N_390,N_3431);
nand U5715 (N_5715,N_2174,N_1196);
and U5716 (N_5716,N_237,N_3732);
or U5717 (N_5717,N_1824,N_2733);
nor U5718 (N_5718,N_1406,N_3088);
and U5719 (N_5719,N_3473,N_931);
nand U5720 (N_5720,N_1224,N_659);
nand U5721 (N_5721,N_2731,N_3111);
nor U5722 (N_5722,N_734,N_411);
xor U5723 (N_5723,N_326,N_1724);
and U5724 (N_5724,N_987,N_84);
or U5725 (N_5725,N_205,N_570);
and U5726 (N_5726,N_3459,N_3900);
and U5727 (N_5727,N_2045,N_2968);
nand U5728 (N_5728,N_71,N_3032);
and U5729 (N_5729,N_1640,N_2244);
or U5730 (N_5730,N_550,N_1893);
nor U5731 (N_5731,N_1995,N_492);
xor U5732 (N_5732,N_367,N_972);
and U5733 (N_5733,N_3515,N_3472);
or U5734 (N_5734,N_376,N_2089);
nand U5735 (N_5735,N_3150,N_3549);
or U5736 (N_5736,N_1148,N_2555);
xor U5737 (N_5737,N_1428,N_1453);
nand U5738 (N_5738,N_2825,N_148);
and U5739 (N_5739,N_2392,N_275);
nor U5740 (N_5740,N_2308,N_1012);
and U5741 (N_5741,N_579,N_3127);
or U5742 (N_5742,N_2985,N_3548);
xnor U5743 (N_5743,N_2042,N_2598);
and U5744 (N_5744,N_1771,N_1783);
nand U5745 (N_5745,N_749,N_1361);
xor U5746 (N_5746,N_927,N_554);
nand U5747 (N_5747,N_3520,N_3622);
nand U5748 (N_5748,N_3313,N_3512);
and U5749 (N_5749,N_1516,N_2616);
nand U5750 (N_5750,N_3454,N_3058);
and U5751 (N_5751,N_1618,N_3797);
nand U5752 (N_5752,N_3338,N_3305);
xnor U5753 (N_5753,N_2655,N_3525);
nor U5754 (N_5754,N_2069,N_1441);
or U5755 (N_5755,N_1781,N_2094);
nor U5756 (N_5756,N_50,N_1788);
xor U5757 (N_5757,N_3838,N_1355);
nand U5758 (N_5758,N_1388,N_1068);
nand U5759 (N_5759,N_476,N_3665);
nor U5760 (N_5760,N_1956,N_3087);
xnor U5761 (N_5761,N_2426,N_2428);
nor U5762 (N_5762,N_2764,N_3486);
nor U5763 (N_5763,N_2883,N_2151);
nor U5764 (N_5764,N_3571,N_2387);
and U5765 (N_5765,N_526,N_2976);
and U5766 (N_5766,N_2662,N_1028);
xnor U5767 (N_5767,N_1896,N_3113);
and U5768 (N_5768,N_1507,N_1980);
or U5769 (N_5769,N_2269,N_3980);
nor U5770 (N_5770,N_2889,N_1172);
xor U5771 (N_5771,N_2944,N_2487);
or U5772 (N_5772,N_1285,N_169);
or U5773 (N_5773,N_1837,N_3640);
or U5774 (N_5774,N_2079,N_3283);
and U5775 (N_5775,N_1318,N_2318);
and U5776 (N_5776,N_2943,N_2526);
nor U5777 (N_5777,N_59,N_143);
nor U5778 (N_5778,N_767,N_1551);
xnor U5779 (N_5779,N_345,N_1368);
nand U5780 (N_5780,N_891,N_793);
and U5781 (N_5781,N_1789,N_3166);
nand U5782 (N_5782,N_2265,N_157);
xnor U5783 (N_5783,N_380,N_3546);
nand U5784 (N_5784,N_2226,N_803);
and U5785 (N_5785,N_3312,N_3530);
xnor U5786 (N_5786,N_2378,N_3364);
nor U5787 (N_5787,N_3293,N_1100);
or U5788 (N_5788,N_3455,N_654);
xor U5789 (N_5789,N_701,N_2646);
nor U5790 (N_5790,N_2098,N_2558);
and U5791 (N_5791,N_371,N_1537);
nand U5792 (N_5792,N_1799,N_1276);
xor U5793 (N_5793,N_2128,N_2157);
nand U5794 (N_5794,N_477,N_1398);
nor U5795 (N_5795,N_3588,N_988);
or U5796 (N_5796,N_1412,N_3610);
and U5797 (N_5797,N_2346,N_728);
and U5798 (N_5798,N_3628,N_738);
and U5799 (N_5799,N_2499,N_1808);
or U5800 (N_5800,N_1031,N_1353);
nor U5801 (N_5801,N_804,N_3792);
xnor U5802 (N_5802,N_399,N_2380);
and U5803 (N_5803,N_805,N_3416);
or U5804 (N_5804,N_3742,N_2303);
or U5805 (N_5805,N_871,N_1861);
nand U5806 (N_5806,N_600,N_2694);
or U5807 (N_5807,N_2819,N_1709);
and U5808 (N_5808,N_3942,N_1432);
and U5809 (N_5809,N_1676,N_2873);
and U5810 (N_5810,N_2771,N_3547);
xor U5811 (N_5811,N_634,N_2408);
nor U5812 (N_5812,N_2154,N_177);
nand U5813 (N_5813,N_2459,N_160);
and U5814 (N_5814,N_3298,N_3015);
nor U5815 (N_5815,N_3696,N_2119);
xnor U5816 (N_5816,N_1326,N_3424);
or U5817 (N_5817,N_3908,N_3592);
nand U5818 (N_5818,N_410,N_3451);
nor U5819 (N_5819,N_1614,N_2734);
and U5820 (N_5820,N_751,N_1654);
xnor U5821 (N_5821,N_227,N_3793);
or U5822 (N_5822,N_247,N_2383);
nor U5823 (N_5823,N_607,N_1715);
nand U5824 (N_5824,N_573,N_1941);
xor U5825 (N_5825,N_395,N_1683);
and U5826 (N_5826,N_250,N_671);
nor U5827 (N_5827,N_3759,N_2450);
and U5828 (N_5828,N_2875,N_490);
xnor U5829 (N_5829,N_256,N_1433);
nor U5830 (N_5830,N_13,N_195);
nand U5831 (N_5831,N_2436,N_3950);
nand U5832 (N_5832,N_171,N_1743);
nand U5833 (N_5833,N_3346,N_2012);
nand U5834 (N_5834,N_2145,N_2234);
or U5835 (N_5835,N_1884,N_1564);
nor U5836 (N_5836,N_1712,N_2905);
xnor U5837 (N_5837,N_3524,N_103);
nor U5838 (N_5838,N_1037,N_2193);
xor U5839 (N_5839,N_1173,N_1403);
or U5840 (N_5840,N_2415,N_1230);
xnor U5841 (N_5841,N_3036,N_629);
or U5842 (N_5842,N_1901,N_2300);
and U5843 (N_5843,N_900,N_127);
nor U5844 (N_5844,N_1518,N_3647);
or U5845 (N_5845,N_1963,N_444);
nor U5846 (N_5846,N_1092,N_2271);
or U5847 (N_5847,N_3436,N_2597);
nand U5848 (N_5848,N_3910,N_508);
nand U5849 (N_5849,N_1913,N_2517);
or U5850 (N_5850,N_807,N_1439);
or U5851 (N_5851,N_57,N_1026);
or U5852 (N_5852,N_3604,N_1669);
nand U5853 (N_5853,N_3060,N_1125);
nor U5854 (N_5854,N_3270,N_3328);
nand U5855 (N_5855,N_3310,N_3895);
or U5856 (N_5856,N_175,N_922);
nor U5857 (N_5857,N_1697,N_3914);
or U5858 (N_5858,N_239,N_595);
nand U5859 (N_5859,N_517,N_2676);
nor U5860 (N_5860,N_489,N_1662);
and U5861 (N_5861,N_3555,N_3);
nand U5862 (N_5862,N_2824,N_3526);
nor U5863 (N_5863,N_2370,N_2973);
and U5864 (N_5864,N_2159,N_1880);
or U5865 (N_5865,N_668,N_2088);
xnor U5866 (N_5866,N_1141,N_2974);
nand U5867 (N_5867,N_1964,N_1117);
xor U5868 (N_5868,N_3862,N_1470);
or U5869 (N_5869,N_1664,N_1726);
and U5870 (N_5870,N_764,N_1816);
or U5871 (N_5871,N_2107,N_2435);
nor U5872 (N_5872,N_2980,N_58);
and U5873 (N_5873,N_339,N_154);
or U5874 (N_5874,N_2178,N_3706);
or U5875 (N_5875,N_3952,N_2443);
nand U5876 (N_5876,N_2063,N_1684);
xnor U5877 (N_5877,N_1245,N_2483);
xnor U5878 (N_5878,N_761,N_2273);
xnor U5879 (N_5879,N_709,N_2360);
and U5880 (N_5880,N_3623,N_1434);
and U5881 (N_5881,N_2666,N_3352);
nor U5882 (N_5882,N_1498,N_2358);
or U5883 (N_5883,N_2476,N_536);
xnor U5884 (N_5884,N_919,N_400);
xor U5885 (N_5885,N_1241,N_366);
xor U5886 (N_5886,N_1904,N_617);
and U5887 (N_5887,N_1645,N_3638);
xor U5888 (N_5888,N_3611,N_39);
nand U5889 (N_5889,N_3599,N_3768);
and U5890 (N_5890,N_3158,N_3194);
xor U5891 (N_5891,N_2469,N_1362);
or U5892 (N_5892,N_3280,N_1998);
or U5893 (N_5893,N_966,N_1166);
nor U5894 (N_5894,N_2634,N_2140);
nor U5895 (N_5895,N_958,N_2248);
or U5896 (N_5896,N_906,N_190);
and U5897 (N_5897,N_1295,N_198);
and U5898 (N_5898,N_167,N_438);
or U5899 (N_5899,N_3218,N_3836);
xnor U5900 (N_5900,N_1375,N_234);
nor U5901 (N_5901,N_1831,N_2797);
nor U5902 (N_5902,N_188,N_231);
nand U5903 (N_5903,N_2238,N_3195);
xor U5904 (N_5904,N_2916,N_3639);
or U5905 (N_5905,N_730,N_1547);
xnor U5906 (N_5906,N_1521,N_3323);
xor U5907 (N_5907,N_3503,N_3661);
xnor U5908 (N_5908,N_2368,N_1181);
or U5909 (N_5909,N_1718,N_711);
and U5910 (N_5910,N_2772,N_2863);
xnor U5911 (N_5911,N_3261,N_3975);
nor U5912 (N_5912,N_281,N_3491);
xor U5913 (N_5913,N_1794,N_3138);
xor U5914 (N_5914,N_997,N_3247);
nor U5915 (N_5915,N_781,N_2962);
and U5916 (N_5916,N_847,N_1146);
xor U5917 (N_5917,N_344,N_2827);
nor U5918 (N_5918,N_118,N_3022);
nor U5919 (N_5919,N_2623,N_1599);
or U5920 (N_5920,N_851,N_2410);
or U5921 (N_5921,N_2101,N_2150);
xor U5922 (N_5922,N_2058,N_2115);
xnor U5923 (N_5923,N_2120,N_1459);
nor U5924 (N_5924,N_3603,N_3854);
or U5925 (N_5925,N_432,N_3532);
nand U5926 (N_5926,N_3693,N_1210);
or U5927 (N_5927,N_3443,N_3579);
nor U5928 (N_5928,N_2929,N_2960);
nor U5929 (N_5929,N_3899,N_3386);
or U5930 (N_5930,N_1097,N_2411);
or U5931 (N_5931,N_3402,N_627);
or U5932 (N_5932,N_1648,N_2445);
and U5933 (N_5933,N_1074,N_284);
nor U5934 (N_5934,N_3669,N_3535);
and U5935 (N_5935,N_1943,N_1445);
xor U5936 (N_5936,N_30,N_3783);
nand U5937 (N_5937,N_1429,N_1960);
nand U5938 (N_5938,N_3275,N_3093);
and U5939 (N_5939,N_2900,N_3921);
xor U5940 (N_5940,N_3192,N_106);
and U5941 (N_5941,N_3909,N_448);
xor U5942 (N_5942,N_3999,N_3962);
xor U5943 (N_5943,N_838,N_3837);
nand U5944 (N_5944,N_2029,N_450);
and U5945 (N_5945,N_953,N_3629);
or U5946 (N_5946,N_409,N_3188);
nor U5947 (N_5947,N_2224,N_1560);
or U5948 (N_5948,N_3516,N_370);
xor U5949 (N_5949,N_403,N_563);
or U5950 (N_5950,N_3121,N_2530);
and U5951 (N_5951,N_3945,N_1840);
xnor U5952 (N_5952,N_676,N_3586);
nor U5953 (N_5953,N_1524,N_1105);
and U5954 (N_5954,N_2429,N_1812);
nand U5955 (N_5955,N_1066,N_3435);
and U5956 (N_5956,N_2057,N_2295);
nor U5957 (N_5957,N_2701,N_2739);
nand U5958 (N_5958,N_3881,N_1520);
nand U5959 (N_5959,N_1251,N_2235);
or U5960 (N_5960,N_1989,N_3151);
and U5961 (N_5961,N_3568,N_1562);
xor U5962 (N_5962,N_3297,N_465);
nor U5963 (N_5963,N_1864,N_3493);
nand U5964 (N_5964,N_2009,N_3932);
nand U5965 (N_5965,N_874,N_744);
xor U5966 (N_5966,N_2073,N_726);
and U5967 (N_5967,N_1578,N_1350);
nor U5968 (N_5968,N_212,N_3621);
and U5969 (N_5969,N_3842,N_223);
nor U5970 (N_5970,N_2839,N_2615);
nand U5971 (N_5971,N_739,N_598);
or U5972 (N_5972,N_3246,N_581);
nor U5973 (N_5973,N_186,N_1383);
or U5974 (N_5974,N_569,N_1178);
or U5975 (N_5975,N_2790,N_3272);
or U5976 (N_5976,N_909,N_1443);
nand U5977 (N_5977,N_3010,N_2164);
and U5978 (N_5978,N_2037,N_1095);
and U5979 (N_5979,N_2928,N_2264);
xnor U5980 (N_5980,N_22,N_1561);
xnor U5981 (N_5981,N_1370,N_3787);
xnor U5982 (N_5982,N_12,N_259);
nor U5983 (N_5983,N_161,N_2574);
xor U5984 (N_5984,N_3636,N_2784);
nor U5985 (N_5985,N_3005,N_2132);
nor U5986 (N_5986,N_787,N_1929);
and U5987 (N_5987,N_2319,N_799);
xnor U5988 (N_5988,N_1367,N_2550);
and U5989 (N_5989,N_1994,N_1132);
xor U5990 (N_5990,N_2258,N_1752);
nand U5991 (N_5991,N_1935,N_1746);
nand U5992 (N_5992,N_3614,N_967);
or U5993 (N_5993,N_2977,N_3594);
or U5994 (N_5994,N_1338,N_1462);
or U5995 (N_5995,N_1266,N_656);
nor U5996 (N_5996,N_3481,N_2937);
or U5997 (N_5997,N_3965,N_2376);
nor U5998 (N_5998,N_2675,N_2475);
nor U5999 (N_5999,N_2015,N_36);
nand U6000 (N_6000,N_2005,N_579);
nand U6001 (N_6001,N_3746,N_2013);
or U6002 (N_6002,N_1933,N_1015);
xor U6003 (N_6003,N_3437,N_273);
nor U6004 (N_6004,N_1290,N_847);
or U6005 (N_6005,N_1044,N_1258);
and U6006 (N_6006,N_2623,N_2964);
or U6007 (N_6007,N_1347,N_3832);
nand U6008 (N_6008,N_2618,N_2567);
nand U6009 (N_6009,N_280,N_2152);
and U6010 (N_6010,N_102,N_2835);
xnor U6011 (N_6011,N_632,N_884);
and U6012 (N_6012,N_756,N_3435);
and U6013 (N_6013,N_1689,N_2969);
and U6014 (N_6014,N_1957,N_2240);
nor U6015 (N_6015,N_1574,N_1030);
nor U6016 (N_6016,N_1981,N_2695);
or U6017 (N_6017,N_1507,N_1247);
xnor U6018 (N_6018,N_1708,N_718);
or U6019 (N_6019,N_1382,N_114);
and U6020 (N_6020,N_2736,N_2415);
and U6021 (N_6021,N_3360,N_923);
nand U6022 (N_6022,N_2175,N_1711);
nor U6023 (N_6023,N_644,N_2451);
or U6024 (N_6024,N_2155,N_1739);
nor U6025 (N_6025,N_3362,N_322);
xnor U6026 (N_6026,N_2629,N_2354);
nor U6027 (N_6027,N_2978,N_3475);
or U6028 (N_6028,N_2473,N_2340);
xnor U6029 (N_6029,N_3915,N_1378);
nor U6030 (N_6030,N_2130,N_2283);
nor U6031 (N_6031,N_2545,N_2343);
and U6032 (N_6032,N_499,N_970);
xnor U6033 (N_6033,N_3266,N_2153);
xnor U6034 (N_6034,N_3699,N_618);
xor U6035 (N_6035,N_1753,N_2772);
nand U6036 (N_6036,N_2652,N_1936);
xnor U6037 (N_6037,N_3213,N_214);
nor U6038 (N_6038,N_507,N_1133);
and U6039 (N_6039,N_2052,N_304);
nand U6040 (N_6040,N_998,N_348);
and U6041 (N_6041,N_1823,N_668);
nand U6042 (N_6042,N_2497,N_802);
or U6043 (N_6043,N_563,N_2371);
nor U6044 (N_6044,N_3263,N_372);
xor U6045 (N_6045,N_3524,N_3509);
xor U6046 (N_6046,N_2482,N_702);
nor U6047 (N_6047,N_1,N_1230);
nor U6048 (N_6048,N_2637,N_3877);
or U6049 (N_6049,N_1543,N_1471);
xor U6050 (N_6050,N_2821,N_558);
nand U6051 (N_6051,N_2357,N_1200);
nor U6052 (N_6052,N_2411,N_2488);
nor U6053 (N_6053,N_507,N_1325);
nor U6054 (N_6054,N_2799,N_3938);
xor U6055 (N_6055,N_3576,N_2200);
nor U6056 (N_6056,N_2198,N_3285);
or U6057 (N_6057,N_2372,N_2149);
and U6058 (N_6058,N_3010,N_1313);
xor U6059 (N_6059,N_392,N_3750);
or U6060 (N_6060,N_1263,N_3702);
xor U6061 (N_6061,N_618,N_3410);
or U6062 (N_6062,N_1336,N_3412);
nor U6063 (N_6063,N_1041,N_40);
nor U6064 (N_6064,N_3377,N_2624);
xor U6065 (N_6065,N_3162,N_1805);
and U6066 (N_6066,N_3161,N_212);
xnor U6067 (N_6067,N_1401,N_2340);
xor U6068 (N_6068,N_2735,N_3766);
or U6069 (N_6069,N_1224,N_2931);
or U6070 (N_6070,N_3699,N_948);
nor U6071 (N_6071,N_901,N_2613);
nor U6072 (N_6072,N_3639,N_2367);
xnor U6073 (N_6073,N_2940,N_1965);
and U6074 (N_6074,N_864,N_410);
and U6075 (N_6075,N_3678,N_333);
nor U6076 (N_6076,N_259,N_1935);
or U6077 (N_6077,N_1318,N_3044);
nand U6078 (N_6078,N_2978,N_2484);
or U6079 (N_6079,N_514,N_1176);
or U6080 (N_6080,N_2940,N_392);
or U6081 (N_6081,N_2622,N_2642);
and U6082 (N_6082,N_1930,N_524);
or U6083 (N_6083,N_3779,N_1262);
and U6084 (N_6084,N_936,N_574);
or U6085 (N_6085,N_1506,N_210);
or U6086 (N_6086,N_2866,N_1296);
nand U6087 (N_6087,N_599,N_1414);
nor U6088 (N_6088,N_1971,N_1426);
nor U6089 (N_6089,N_2566,N_3108);
xor U6090 (N_6090,N_3564,N_2968);
nand U6091 (N_6091,N_209,N_2219);
and U6092 (N_6092,N_241,N_1612);
or U6093 (N_6093,N_2497,N_3441);
nand U6094 (N_6094,N_146,N_3251);
and U6095 (N_6095,N_224,N_2377);
or U6096 (N_6096,N_2491,N_2157);
nand U6097 (N_6097,N_674,N_929);
xnor U6098 (N_6098,N_1322,N_3411);
xnor U6099 (N_6099,N_1611,N_1496);
nand U6100 (N_6100,N_1232,N_1538);
nand U6101 (N_6101,N_1657,N_3860);
and U6102 (N_6102,N_2754,N_1707);
and U6103 (N_6103,N_3100,N_1714);
or U6104 (N_6104,N_3156,N_1605);
or U6105 (N_6105,N_3390,N_1435);
nand U6106 (N_6106,N_923,N_794);
and U6107 (N_6107,N_1613,N_718);
xnor U6108 (N_6108,N_1866,N_719);
nor U6109 (N_6109,N_1252,N_2909);
nor U6110 (N_6110,N_2342,N_3956);
nand U6111 (N_6111,N_2953,N_3138);
nand U6112 (N_6112,N_2248,N_2668);
nor U6113 (N_6113,N_2949,N_543);
or U6114 (N_6114,N_2752,N_2825);
and U6115 (N_6115,N_2405,N_2818);
and U6116 (N_6116,N_2056,N_991);
nor U6117 (N_6117,N_288,N_1795);
or U6118 (N_6118,N_1664,N_972);
nor U6119 (N_6119,N_272,N_2347);
nand U6120 (N_6120,N_2423,N_451);
xor U6121 (N_6121,N_616,N_2292);
xor U6122 (N_6122,N_3073,N_2496);
and U6123 (N_6123,N_437,N_1753);
nor U6124 (N_6124,N_3355,N_2547);
or U6125 (N_6125,N_1948,N_558);
xor U6126 (N_6126,N_609,N_2358);
xor U6127 (N_6127,N_894,N_795);
and U6128 (N_6128,N_2586,N_2824);
nor U6129 (N_6129,N_2765,N_912);
xnor U6130 (N_6130,N_1585,N_3689);
or U6131 (N_6131,N_1827,N_1860);
nand U6132 (N_6132,N_340,N_650);
or U6133 (N_6133,N_1761,N_2860);
xnor U6134 (N_6134,N_3116,N_237);
nor U6135 (N_6135,N_279,N_186);
and U6136 (N_6136,N_402,N_3483);
or U6137 (N_6137,N_2463,N_89);
nor U6138 (N_6138,N_913,N_1004);
nor U6139 (N_6139,N_2806,N_32);
or U6140 (N_6140,N_2652,N_739);
xnor U6141 (N_6141,N_1080,N_587);
or U6142 (N_6142,N_3941,N_2087);
xor U6143 (N_6143,N_2189,N_2245);
xnor U6144 (N_6144,N_562,N_24);
and U6145 (N_6145,N_1630,N_1793);
nand U6146 (N_6146,N_3801,N_2584);
or U6147 (N_6147,N_1554,N_975);
nand U6148 (N_6148,N_1694,N_2550);
nor U6149 (N_6149,N_478,N_2034);
and U6150 (N_6150,N_3243,N_2778);
and U6151 (N_6151,N_2216,N_539);
and U6152 (N_6152,N_3192,N_11);
and U6153 (N_6153,N_2686,N_2596);
xnor U6154 (N_6154,N_2745,N_2033);
nor U6155 (N_6155,N_2004,N_553);
xnor U6156 (N_6156,N_3425,N_884);
and U6157 (N_6157,N_2669,N_715);
and U6158 (N_6158,N_869,N_736);
and U6159 (N_6159,N_249,N_515);
xnor U6160 (N_6160,N_3398,N_750);
nor U6161 (N_6161,N_3904,N_1401);
xnor U6162 (N_6162,N_1811,N_1318);
nand U6163 (N_6163,N_2945,N_2539);
and U6164 (N_6164,N_1748,N_3025);
xor U6165 (N_6165,N_968,N_434);
nand U6166 (N_6166,N_1008,N_1028);
xor U6167 (N_6167,N_1575,N_3637);
or U6168 (N_6168,N_3720,N_3590);
xnor U6169 (N_6169,N_713,N_697);
and U6170 (N_6170,N_1815,N_2251);
nor U6171 (N_6171,N_3386,N_561);
and U6172 (N_6172,N_1111,N_3303);
nand U6173 (N_6173,N_2917,N_3740);
nand U6174 (N_6174,N_1921,N_3509);
xor U6175 (N_6175,N_904,N_2986);
xor U6176 (N_6176,N_2391,N_2753);
and U6177 (N_6177,N_1282,N_3103);
xnor U6178 (N_6178,N_1288,N_3812);
or U6179 (N_6179,N_771,N_432);
nand U6180 (N_6180,N_2849,N_3345);
xor U6181 (N_6181,N_2552,N_1951);
and U6182 (N_6182,N_3185,N_3539);
and U6183 (N_6183,N_3983,N_2407);
and U6184 (N_6184,N_3042,N_1080);
nand U6185 (N_6185,N_550,N_512);
xnor U6186 (N_6186,N_3886,N_3052);
and U6187 (N_6187,N_465,N_828);
nor U6188 (N_6188,N_448,N_3338);
and U6189 (N_6189,N_3934,N_1434);
xnor U6190 (N_6190,N_3424,N_3278);
nand U6191 (N_6191,N_1838,N_3639);
nand U6192 (N_6192,N_138,N_3977);
xor U6193 (N_6193,N_6,N_1426);
nor U6194 (N_6194,N_1995,N_1243);
and U6195 (N_6195,N_3026,N_1702);
nor U6196 (N_6196,N_1089,N_454);
or U6197 (N_6197,N_1341,N_1904);
and U6198 (N_6198,N_902,N_612);
and U6199 (N_6199,N_1639,N_1413);
nor U6200 (N_6200,N_2505,N_3309);
nand U6201 (N_6201,N_2732,N_616);
and U6202 (N_6202,N_1550,N_2121);
or U6203 (N_6203,N_3473,N_59);
nand U6204 (N_6204,N_3247,N_2796);
nor U6205 (N_6205,N_1474,N_1389);
or U6206 (N_6206,N_700,N_2032);
or U6207 (N_6207,N_2736,N_3822);
and U6208 (N_6208,N_1272,N_2858);
nor U6209 (N_6209,N_1874,N_2836);
nor U6210 (N_6210,N_2071,N_979);
and U6211 (N_6211,N_1147,N_2393);
and U6212 (N_6212,N_3276,N_2674);
xnor U6213 (N_6213,N_3579,N_2908);
xnor U6214 (N_6214,N_239,N_2397);
xnor U6215 (N_6215,N_2974,N_1683);
xor U6216 (N_6216,N_3806,N_2154);
and U6217 (N_6217,N_2644,N_1675);
and U6218 (N_6218,N_3651,N_2549);
and U6219 (N_6219,N_3057,N_425);
nor U6220 (N_6220,N_29,N_3713);
and U6221 (N_6221,N_1981,N_2693);
nand U6222 (N_6222,N_466,N_3316);
xnor U6223 (N_6223,N_2032,N_556);
xnor U6224 (N_6224,N_1176,N_1669);
nor U6225 (N_6225,N_1800,N_2078);
and U6226 (N_6226,N_2424,N_1944);
and U6227 (N_6227,N_979,N_1449);
or U6228 (N_6228,N_3906,N_31);
and U6229 (N_6229,N_2140,N_1127);
nor U6230 (N_6230,N_3561,N_1494);
xor U6231 (N_6231,N_1523,N_675);
nor U6232 (N_6232,N_3875,N_484);
xor U6233 (N_6233,N_2501,N_2755);
nand U6234 (N_6234,N_3845,N_3533);
nand U6235 (N_6235,N_3213,N_2941);
or U6236 (N_6236,N_3082,N_274);
nand U6237 (N_6237,N_1868,N_48);
xor U6238 (N_6238,N_3418,N_1886);
nor U6239 (N_6239,N_3794,N_1116);
or U6240 (N_6240,N_1960,N_1089);
or U6241 (N_6241,N_1007,N_3614);
nand U6242 (N_6242,N_870,N_290);
xnor U6243 (N_6243,N_3616,N_721);
xnor U6244 (N_6244,N_133,N_2513);
or U6245 (N_6245,N_3134,N_1766);
nor U6246 (N_6246,N_19,N_3572);
and U6247 (N_6247,N_1796,N_2786);
nand U6248 (N_6248,N_842,N_1210);
nor U6249 (N_6249,N_2468,N_2902);
or U6250 (N_6250,N_3709,N_2772);
and U6251 (N_6251,N_3312,N_749);
xor U6252 (N_6252,N_2248,N_956);
and U6253 (N_6253,N_1524,N_157);
nand U6254 (N_6254,N_1049,N_2659);
and U6255 (N_6255,N_2217,N_3120);
and U6256 (N_6256,N_1248,N_547);
or U6257 (N_6257,N_109,N_2700);
xor U6258 (N_6258,N_1020,N_3272);
and U6259 (N_6259,N_3304,N_453);
xnor U6260 (N_6260,N_3389,N_155);
or U6261 (N_6261,N_3865,N_893);
or U6262 (N_6262,N_510,N_386);
nand U6263 (N_6263,N_2422,N_2665);
nor U6264 (N_6264,N_2089,N_596);
and U6265 (N_6265,N_3782,N_3989);
nor U6266 (N_6266,N_2079,N_3758);
or U6267 (N_6267,N_347,N_1079);
xnor U6268 (N_6268,N_2097,N_2045);
or U6269 (N_6269,N_50,N_521);
nor U6270 (N_6270,N_2176,N_1535);
nand U6271 (N_6271,N_773,N_1052);
nand U6272 (N_6272,N_3966,N_3111);
and U6273 (N_6273,N_1343,N_1674);
nand U6274 (N_6274,N_1710,N_917);
and U6275 (N_6275,N_1165,N_3043);
nand U6276 (N_6276,N_1705,N_119);
and U6277 (N_6277,N_3844,N_2257);
and U6278 (N_6278,N_83,N_2436);
xnor U6279 (N_6279,N_872,N_1463);
and U6280 (N_6280,N_3498,N_2095);
or U6281 (N_6281,N_3796,N_2660);
or U6282 (N_6282,N_21,N_1124);
xnor U6283 (N_6283,N_3129,N_2157);
and U6284 (N_6284,N_2554,N_1285);
or U6285 (N_6285,N_3943,N_1754);
and U6286 (N_6286,N_2316,N_1628);
nor U6287 (N_6287,N_3405,N_3467);
xor U6288 (N_6288,N_1931,N_2832);
nor U6289 (N_6289,N_3806,N_3015);
and U6290 (N_6290,N_3086,N_2090);
and U6291 (N_6291,N_1752,N_2755);
and U6292 (N_6292,N_1998,N_1896);
xnor U6293 (N_6293,N_2838,N_249);
nor U6294 (N_6294,N_2851,N_282);
and U6295 (N_6295,N_344,N_2301);
xor U6296 (N_6296,N_1498,N_2634);
xnor U6297 (N_6297,N_499,N_410);
or U6298 (N_6298,N_541,N_2687);
nor U6299 (N_6299,N_584,N_2098);
nor U6300 (N_6300,N_2406,N_3405);
nand U6301 (N_6301,N_585,N_1859);
and U6302 (N_6302,N_3606,N_2939);
and U6303 (N_6303,N_1434,N_2100);
nor U6304 (N_6304,N_1054,N_568);
or U6305 (N_6305,N_1773,N_3911);
nor U6306 (N_6306,N_723,N_1390);
or U6307 (N_6307,N_294,N_1436);
or U6308 (N_6308,N_778,N_3590);
nor U6309 (N_6309,N_2417,N_2107);
or U6310 (N_6310,N_2380,N_1835);
nor U6311 (N_6311,N_3082,N_3293);
nor U6312 (N_6312,N_894,N_2439);
or U6313 (N_6313,N_779,N_909);
and U6314 (N_6314,N_3469,N_943);
and U6315 (N_6315,N_3843,N_1089);
nand U6316 (N_6316,N_2965,N_3665);
xor U6317 (N_6317,N_93,N_2748);
nand U6318 (N_6318,N_1572,N_2841);
xor U6319 (N_6319,N_1873,N_2976);
nor U6320 (N_6320,N_567,N_1039);
xnor U6321 (N_6321,N_246,N_1163);
and U6322 (N_6322,N_737,N_3279);
or U6323 (N_6323,N_298,N_2566);
nand U6324 (N_6324,N_368,N_3380);
or U6325 (N_6325,N_3479,N_2310);
or U6326 (N_6326,N_611,N_3747);
or U6327 (N_6327,N_1069,N_3522);
nand U6328 (N_6328,N_2311,N_2720);
or U6329 (N_6329,N_1681,N_1264);
or U6330 (N_6330,N_2213,N_3126);
nand U6331 (N_6331,N_2438,N_1908);
nand U6332 (N_6332,N_3977,N_47);
and U6333 (N_6333,N_1691,N_3419);
xor U6334 (N_6334,N_1220,N_2385);
or U6335 (N_6335,N_2583,N_2679);
nor U6336 (N_6336,N_2352,N_3122);
nand U6337 (N_6337,N_107,N_520);
xnor U6338 (N_6338,N_521,N_1974);
xor U6339 (N_6339,N_1777,N_3857);
and U6340 (N_6340,N_1477,N_3433);
and U6341 (N_6341,N_985,N_1968);
nand U6342 (N_6342,N_827,N_485);
nand U6343 (N_6343,N_1,N_2869);
or U6344 (N_6344,N_2206,N_3758);
xnor U6345 (N_6345,N_2741,N_3940);
and U6346 (N_6346,N_2010,N_586);
xor U6347 (N_6347,N_1305,N_2612);
xnor U6348 (N_6348,N_3527,N_1776);
nand U6349 (N_6349,N_1702,N_1060);
nand U6350 (N_6350,N_1301,N_3496);
nor U6351 (N_6351,N_1333,N_197);
xnor U6352 (N_6352,N_2357,N_1560);
nor U6353 (N_6353,N_1904,N_2838);
and U6354 (N_6354,N_3060,N_2585);
and U6355 (N_6355,N_387,N_2486);
xnor U6356 (N_6356,N_3061,N_2730);
nand U6357 (N_6357,N_1976,N_703);
nor U6358 (N_6358,N_1151,N_4);
xor U6359 (N_6359,N_2041,N_3161);
nor U6360 (N_6360,N_1622,N_2768);
xor U6361 (N_6361,N_2295,N_1922);
nor U6362 (N_6362,N_2482,N_1987);
xor U6363 (N_6363,N_2655,N_1133);
xor U6364 (N_6364,N_253,N_3959);
nand U6365 (N_6365,N_2913,N_1281);
xnor U6366 (N_6366,N_3771,N_3091);
or U6367 (N_6367,N_369,N_738);
nand U6368 (N_6368,N_3799,N_868);
nand U6369 (N_6369,N_2064,N_1600);
nand U6370 (N_6370,N_3507,N_3084);
nand U6371 (N_6371,N_1434,N_545);
xor U6372 (N_6372,N_2919,N_234);
or U6373 (N_6373,N_2036,N_3248);
or U6374 (N_6374,N_1395,N_38);
nor U6375 (N_6375,N_3985,N_1489);
nand U6376 (N_6376,N_2257,N_1264);
nand U6377 (N_6377,N_2512,N_872);
nor U6378 (N_6378,N_1319,N_1482);
and U6379 (N_6379,N_2850,N_3438);
xor U6380 (N_6380,N_637,N_81);
nor U6381 (N_6381,N_661,N_2540);
and U6382 (N_6382,N_2036,N_1344);
and U6383 (N_6383,N_3725,N_3693);
xor U6384 (N_6384,N_2263,N_2977);
or U6385 (N_6385,N_3256,N_1544);
and U6386 (N_6386,N_3804,N_1783);
nor U6387 (N_6387,N_1740,N_3917);
nand U6388 (N_6388,N_1804,N_1527);
nand U6389 (N_6389,N_2404,N_960);
or U6390 (N_6390,N_697,N_3909);
and U6391 (N_6391,N_2445,N_312);
xnor U6392 (N_6392,N_3731,N_213);
xnor U6393 (N_6393,N_698,N_187);
nand U6394 (N_6394,N_985,N_354);
and U6395 (N_6395,N_1144,N_1289);
nand U6396 (N_6396,N_3140,N_1400);
nor U6397 (N_6397,N_2237,N_1850);
xor U6398 (N_6398,N_797,N_21);
nor U6399 (N_6399,N_1997,N_1746);
xor U6400 (N_6400,N_2892,N_3756);
and U6401 (N_6401,N_1927,N_3160);
or U6402 (N_6402,N_1067,N_355);
and U6403 (N_6403,N_160,N_932);
nand U6404 (N_6404,N_3632,N_3215);
nand U6405 (N_6405,N_1377,N_2949);
or U6406 (N_6406,N_2294,N_3898);
nor U6407 (N_6407,N_801,N_2087);
or U6408 (N_6408,N_3199,N_3331);
nand U6409 (N_6409,N_1194,N_759);
nor U6410 (N_6410,N_3166,N_1980);
xnor U6411 (N_6411,N_2761,N_2472);
nor U6412 (N_6412,N_2012,N_112);
and U6413 (N_6413,N_2720,N_853);
xor U6414 (N_6414,N_2961,N_2674);
and U6415 (N_6415,N_472,N_2698);
xor U6416 (N_6416,N_734,N_3165);
nor U6417 (N_6417,N_3333,N_3035);
xnor U6418 (N_6418,N_3245,N_2588);
or U6419 (N_6419,N_721,N_1410);
nand U6420 (N_6420,N_2726,N_951);
or U6421 (N_6421,N_818,N_3692);
xnor U6422 (N_6422,N_3036,N_3697);
xnor U6423 (N_6423,N_317,N_1105);
and U6424 (N_6424,N_3320,N_1971);
or U6425 (N_6425,N_1486,N_2971);
and U6426 (N_6426,N_3412,N_1757);
nand U6427 (N_6427,N_3849,N_774);
nor U6428 (N_6428,N_2633,N_419);
and U6429 (N_6429,N_2928,N_2126);
nor U6430 (N_6430,N_1167,N_1873);
xnor U6431 (N_6431,N_2315,N_1832);
xor U6432 (N_6432,N_2666,N_1829);
or U6433 (N_6433,N_719,N_3324);
or U6434 (N_6434,N_2640,N_143);
or U6435 (N_6435,N_1366,N_3431);
xnor U6436 (N_6436,N_1131,N_1942);
and U6437 (N_6437,N_2050,N_2221);
nor U6438 (N_6438,N_2210,N_2863);
and U6439 (N_6439,N_2672,N_3257);
and U6440 (N_6440,N_3309,N_3441);
nand U6441 (N_6441,N_3245,N_3050);
nor U6442 (N_6442,N_41,N_3536);
or U6443 (N_6443,N_313,N_3825);
or U6444 (N_6444,N_359,N_1415);
nand U6445 (N_6445,N_3066,N_1004);
nor U6446 (N_6446,N_745,N_2563);
or U6447 (N_6447,N_2732,N_3878);
nor U6448 (N_6448,N_1660,N_2348);
or U6449 (N_6449,N_675,N_2772);
and U6450 (N_6450,N_1742,N_2287);
or U6451 (N_6451,N_1532,N_678);
nand U6452 (N_6452,N_100,N_3982);
nor U6453 (N_6453,N_1021,N_3103);
nor U6454 (N_6454,N_1048,N_3161);
xnor U6455 (N_6455,N_556,N_1139);
nor U6456 (N_6456,N_145,N_2289);
and U6457 (N_6457,N_2727,N_548);
or U6458 (N_6458,N_2535,N_3837);
xor U6459 (N_6459,N_1691,N_2509);
xnor U6460 (N_6460,N_2945,N_2198);
and U6461 (N_6461,N_1345,N_671);
nor U6462 (N_6462,N_3197,N_3675);
or U6463 (N_6463,N_3297,N_2404);
nand U6464 (N_6464,N_3423,N_2497);
xor U6465 (N_6465,N_782,N_737);
or U6466 (N_6466,N_3339,N_1300);
or U6467 (N_6467,N_2102,N_1549);
xnor U6468 (N_6468,N_185,N_2578);
nand U6469 (N_6469,N_2386,N_2334);
or U6470 (N_6470,N_3616,N_3477);
and U6471 (N_6471,N_3016,N_3261);
or U6472 (N_6472,N_1668,N_271);
xnor U6473 (N_6473,N_3302,N_1115);
or U6474 (N_6474,N_3985,N_2196);
nor U6475 (N_6475,N_1407,N_1020);
nand U6476 (N_6476,N_456,N_102);
nor U6477 (N_6477,N_319,N_141);
nor U6478 (N_6478,N_1697,N_1645);
or U6479 (N_6479,N_1052,N_1860);
nand U6480 (N_6480,N_1323,N_1591);
xor U6481 (N_6481,N_715,N_3803);
and U6482 (N_6482,N_1071,N_1447);
nand U6483 (N_6483,N_3016,N_2327);
and U6484 (N_6484,N_1475,N_2942);
and U6485 (N_6485,N_1622,N_821);
or U6486 (N_6486,N_1725,N_3090);
nand U6487 (N_6487,N_472,N_1987);
nor U6488 (N_6488,N_923,N_189);
nand U6489 (N_6489,N_764,N_79);
nor U6490 (N_6490,N_2342,N_3287);
xor U6491 (N_6491,N_3856,N_2392);
and U6492 (N_6492,N_368,N_678);
nor U6493 (N_6493,N_1422,N_992);
or U6494 (N_6494,N_1182,N_1251);
and U6495 (N_6495,N_2647,N_5);
nor U6496 (N_6496,N_1946,N_568);
xor U6497 (N_6497,N_2077,N_2433);
nor U6498 (N_6498,N_2073,N_1080);
and U6499 (N_6499,N_626,N_1634);
xor U6500 (N_6500,N_3962,N_617);
and U6501 (N_6501,N_1994,N_1109);
or U6502 (N_6502,N_3609,N_3360);
nand U6503 (N_6503,N_3319,N_634);
xor U6504 (N_6504,N_3450,N_225);
and U6505 (N_6505,N_2204,N_2217);
nand U6506 (N_6506,N_2739,N_3686);
xor U6507 (N_6507,N_162,N_1781);
or U6508 (N_6508,N_1653,N_452);
nor U6509 (N_6509,N_806,N_2556);
xor U6510 (N_6510,N_544,N_2822);
and U6511 (N_6511,N_402,N_488);
and U6512 (N_6512,N_493,N_2356);
nand U6513 (N_6513,N_601,N_1759);
and U6514 (N_6514,N_3133,N_3029);
or U6515 (N_6515,N_2477,N_2492);
and U6516 (N_6516,N_3299,N_2788);
nor U6517 (N_6517,N_2762,N_2);
nand U6518 (N_6518,N_2799,N_2805);
nor U6519 (N_6519,N_3084,N_3987);
nor U6520 (N_6520,N_1542,N_821);
or U6521 (N_6521,N_785,N_3058);
or U6522 (N_6522,N_3849,N_3860);
nand U6523 (N_6523,N_763,N_1410);
or U6524 (N_6524,N_2956,N_777);
nand U6525 (N_6525,N_3937,N_464);
or U6526 (N_6526,N_980,N_399);
nand U6527 (N_6527,N_2341,N_3791);
nand U6528 (N_6528,N_3639,N_2291);
nand U6529 (N_6529,N_3720,N_844);
and U6530 (N_6530,N_3555,N_3627);
xor U6531 (N_6531,N_1417,N_1421);
and U6532 (N_6532,N_1409,N_1276);
xnor U6533 (N_6533,N_1559,N_1754);
or U6534 (N_6534,N_3819,N_2220);
nand U6535 (N_6535,N_1286,N_2867);
nand U6536 (N_6536,N_2822,N_1071);
nor U6537 (N_6537,N_713,N_3904);
xnor U6538 (N_6538,N_2249,N_88);
nor U6539 (N_6539,N_494,N_991);
nand U6540 (N_6540,N_2200,N_76);
and U6541 (N_6541,N_2513,N_1546);
or U6542 (N_6542,N_1537,N_1059);
nand U6543 (N_6543,N_2148,N_896);
nor U6544 (N_6544,N_2831,N_3002);
xnor U6545 (N_6545,N_1053,N_342);
xor U6546 (N_6546,N_390,N_410);
and U6547 (N_6547,N_968,N_2565);
nand U6548 (N_6548,N_3718,N_3441);
or U6549 (N_6549,N_671,N_1941);
xnor U6550 (N_6550,N_3648,N_2779);
or U6551 (N_6551,N_1610,N_1776);
and U6552 (N_6552,N_2281,N_3758);
nand U6553 (N_6553,N_2802,N_3603);
and U6554 (N_6554,N_719,N_1798);
xnor U6555 (N_6555,N_1565,N_176);
nand U6556 (N_6556,N_686,N_2885);
and U6557 (N_6557,N_1086,N_3656);
nor U6558 (N_6558,N_3772,N_2040);
nor U6559 (N_6559,N_1784,N_618);
nand U6560 (N_6560,N_131,N_776);
nand U6561 (N_6561,N_1769,N_683);
or U6562 (N_6562,N_2702,N_1647);
nand U6563 (N_6563,N_1390,N_385);
and U6564 (N_6564,N_1418,N_3998);
nand U6565 (N_6565,N_226,N_3483);
nand U6566 (N_6566,N_2217,N_2751);
nand U6567 (N_6567,N_1157,N_2881);
nor U6568 (N_6568,N_901,N_1645);
nand U6569 (N_6569,N_3436,N_249);
xor U6570 (N_6570,N_3489,N_2445);
nor U6571 (N_6571,N_1885,N_516);
nand U6572 (N_6572,N_1451,N_1394);
nand U6573 (N_6573,N_3982,N_1016);
xnor U6574 (N_6574,N_326,N_3951);
nor U6575 (N_6575,N_106,N_2742);
and U6576 (N_6576,N_3248,N_1634);
xor U6577 (N_6577,N_3405,N_3714);
and U6578 (N_6578,N_95,N_2937);
and U6579 (N_6579,N_1669,N_2919);
nor U6580 (N_6580,N_1831,N_1635);
and U6581 (N_6581,N_1523,N_747);
nand U6582 (N_6582,N_1835,N_3152);
nor U6583 (N_6583,N_3730,N_3519);
xnor U6584 (N_6584,N_1029,N_3906);
or U6585 (N_6585,N_2373,N_1766);
and U6586 (N_6586,N_1675,N_3854);
and U6587 (N_6587,N_2378,N_1088);
and U6588 (N_6588,N_2909,N_2635);
xor U6589 (N_6589,N_3658,N_3168);
nor U6590 (N_6590,N_3258,N_2962);
and U6591 (N_6591,N_2111,N_2558);
or U6592 (N_6592,N_108,N_1685);
and U6593 (N_6593,N_474,N_2493);
xor U6594 (N_6594,N_583,N_2274);
xor U6595 (N_6595,N_2115,N_2446);
nand U6596 (N_6596,N_1666,N_2199);
nor U6597 (N_6597,N_1714,N_3075);
nor U6598 (N_6598,N_1699,N_2136);
or U6599 (N_6599,N_2139,N_1651);
nor U6600 (N_6600,N_188,N_3265);
xor U6601 (N_6601,N_196,N_976);
xnor U6602 (N_6602,N_3206,N_1769);
nand U6603 (N_6603,N_602,N_1530);
and U6604 (N_6604,N_95,N_479);
nor U6605 (N_6605,N_177,N_3512);
or U6606 (N_6606,N_2172,N_1748);
nand U6607 (N_6607,N_3347,N_3506);
or U6608 (N_6608,N_2628,N_3410);
nor U6609 (N_6609,N_77,N_2057);
or U6610 (N_6610,N_1102,N_1049);
or U6611 (N_6611,N_959,N_2734);
or U6612 (N_6612,N_2002,N_2021);
xor U6613 (N_6613,N_3021,N_3947);
or U6614 (N_6614,N_1796,N_1059);
and U6615 (N_6615,N_2680,N_739);
nor U6616 (N_6616,N_2162,N_667);
nor U6617 (N_6617,N_2379,N_2351);
xnor U6618 (N_6618,N_1907,N_3541);
or U6619 (N_6619,N_2048,N_827);
and U6620 (N_6620,N_909,N_1856);
xnor U6621 (N_6621,N_1944,N_2036);
nand U6622 (N_6622,N_1021,N_3829);
nand U6623 (N_6623,N_296,N_3617);
nand U6624 (N_6624,N_312,N_1724);
nor U6625 (N_6625,N_1340,N_1539);
and U6626 (N_6626,N_428,N_1154);
xnor U6627 (N_6627,N_3135,N_3370);
nand U6628 (N_6628,N_264,N_632);
nor U6629 (N_6629,N_45,N_2943);
nor U6630 (N_6630,N_3306,N_141);
xnor U6631 (N_6631,N_156,N_3667);
or U6632 (N_6632,N_2434,N_2852);
xnor U6633 (N_6633,N_2229,N_341);
nor U6634 (N_6634,N_3151,N_803);
nand U6635 (N_6635,N_2769,N_2749);
xor U6636 (N_6636,N_3997,N_660);
xor U6637 (N_6637,N_1136,N_1339);
and U6638 (N_6638,N_3449,N_3472);
nand U6639 (N_6639,N_589,N_1988);
or U6640 (N_6640,N_2956,N_39);
xnor U6641 (N_6641,N_3710,N_3936);
nand U6642 (N_6642,N_10,N_113);
and U6643 (N_6643,N_731,N_2828);
nor U6644 (N_6644,N_3343,N_3349);
and U6645 (N_6645,N_3777,N_2724);
and U6646 (N_6646,N_3653,N_1808);
or U6647 (N_6647,N_627,N_3600);
xnor U6648 (N_6648,N_2593,N_201);
nand U6649 (N_6649,N_3991,N_2513);
nand U6650 (N_6650,N_79,N_478);
nor U6651 (N_6651,N_2817,N_2088);
or U6652 (N_6652,N_1352,N_3190);
nor U6653 (N_6653,N_1654,N_1081);
and U6654 (N_6654,N_3654,N_2910);
or U6655 (N_6655,N_966,N_3338);
nand U6656 (N_6656,N_807,N_1597);
or U6657 (N_6657,N_846,N_1631);
or U6658 (N_6658,N_1904,N_611);
xor U6659 (N_6659,N_2201,N_2817);
xnor U6660 (N_6660,N_2263,N_3954);
and U6661 (N_6661,N_3928,N_2827);
or U6662 (N_6662,N_3843,N_6);
nor U6663 (N_6663,N_2678,N_2880);
or U6664 (N_6664,N_1384,N_735);
xor U6665 (N_6665,N_3636,N_204);
or U6666 (N_6666,N_2576,N_1845);
and U6667 (N_6667,N_3317,N_3561);
nor U6668 (N_6668,N_2163,N_2865);
and U6669 (N_6669,N_769,N_1206);
xnor U6670 (N_6670,N_410,N_1417);
nand U6671 (N_6671,N_533,N_3890);
or U6672 (N_6672,N_648,N_2951);
xor U6673 (N_6673,N_1963,N_1223);
and U6674 (N_6674,N_1794,N_3566);
nor U6675 (N_6675,N_2271,N_1140);
nand U6676 (N_6676,N_3959,N_2246);
and U6677 (N_6677,N_2879,N_2307);
or U6678 (N_6678,N_2934,N_643);
nor U6679 (N_6679,N_812,N_1865);
nand U6680 (N_6680,N_3237,N_478);
nor U6681 (N_6681,N_3869,N_1493);
nand U6682 (N_6682,N_1269,N_3857);
and U6683 (N_6683,N_3120,N_1292);
nor U6684 (N_6684,N_2897,N_2129);
and U6685 (N_6685,N_158,N_3786);
nor U6686 (N_6686,N_1250,N_184);
nor U6687 (N_6687,N_24,N_1438);
nor U6688 (N_6688,N_548,N_1907);
or U6689 (N_6689,N_1232,N_306);
nand U6690 (N_6690,N_2093,N_1353);
xnor U6691 (N_6691,N_2601,N_677);
nor U6692 (N_6692,N_1829,N_1957);
nor U6693 (N_6693,N_71,N_2839);
xnor U6694 (N_6694,N_2275,N_3033);
xor U6695 (N_6695,N_3338,N_2203);
xor U6696 (N_6696,N_820,N_2119);
xnor U6697 (N_6697,N_1648,N_3034);
xor U6698 (N_6698,N_1540,N_1114);
xor U6699 (N_6699,N_206,N_1912);
xnor U6700 (N_6700,N_882,N_3353);
or U6701 (N_6701,N_1577,N_770);
and U6702 (N_6702,N_380,N_3471);
nor U6703 (N_6703,N_2909,N_1799);
xor U6704 (N_6704,N_2324,N_1620);
xnor U6705 (N_6705,N_3635,N_2246);
nand U6706 (N_6706,N_179,N_316);
nand U6707 (N_6707,N_1068,N_224);
nand U6708 (N_6708,N_360,N_3420);
nor U6709 (N_6709,N_1127,N_706);
or U6710 (N_6710,N_505,N_101);
or U6711 (N_6711,N_1021,N_3725);
nor U6712 (N_6712,N_2078,N_1461);
nand U6713 (N_6713,N_3541,N_2319);
xnor U6714 (N_6714,N_2891,N_1948);
nor U6715 (N_6715,N_434,N_2233);
nor U6716 (N_6716,N_1239,N_609);
nor U6717 (N_6717,N_749,N_3127);
or U6718 (N_6718,N_1725,N_2263);
nand U6719 (N_6719,N_249,N_1242);
and U6720 (N_6720,N_2147,N_558);
xnor U6721 (N_6721,N_3857,N_2330);
nand U6722 (N_6722,N_508,N_685);
and U6723 (N_6723,N_3210,N_1634);
or U6724 (N_6724,N_149,N_2103);
xnor U6725 (N_6725,N_346,N_282);
and U6726 (N_6726,N_2283,N_2614);
nand U6727 (N_6727,N_2482,N_2243);
and U6728 (N_6728,N_1101,N_327);
and U6729 (N_6729,N_1905,N_3096);
nor U6730 (N_6730,N_2475,N_1909);
nor U6731 (N_6731,N_2475,N_409);
and U6732 (N_6732,N_740,N_2233);
and U6733 (N_6733,N_3566,N_1898);
and U6734 (N_6734,N_3151,N_3006);
xor U6735 (N_6735,N_3602,N_3523);
and U6736 (N_6736,N_623,N_282);
xnor U6737 (N_6737,N_2151,N_270);
nand U6738 (N_6738,N_3004,N_3810);
or U6739 (N_6739,N_3652,N_3130);
nand U6740 (N_6740,N_2886,N_2310);
xnor U6741 (N_6741,N_3357,N_390);
nor U6742 (N_6742,N_3025,N_3881);
nor U6743 (N_6743,N_2574,N_1668);
nor U6744 (N_6744,N_689,N_1464);
nor U6745 (N_6745,N_1112,N_2403);
and U6746 (N_6746,N_3906,N_3295);
or U6747 (N_6747,N_933,N_1877);
nand U6748 (N_6748,N_1675,N_3018);
nor U6749 (N_6749,N_3177,N_2444);
xnor U6750 (N_6750,N_2779,N_878);
nand U6751 (N_6751,N_1114,N_3396);
xor U6752 (N_6752,N_2056,N_1622);
and U6753 (N_6753,N_1826,N_1921);
and U6754 (N_6754,N_1475,N_3233);
or U6755 (N_6755,N_822,N_2388);
nand U6756 (N_6756,N_499,N_3199);
nor U6757 (N_6757,N_2590,N_2954);
or U6758 (N_6758,N_2121,N_1532);
or U6759 (N_6759,N_2809,N_3405);
xor U6760 (N_6760,N_1918,N_3166);
nor U6761 (N_6761,N_1592,N_1720);
nor U6762 (N_6762,N_3875,N_3888);
nand U6763 (N_6763,N_3907,N_3298);
and U6764 (N_6764,N_1433,N_1198);
xnor U6765 (N_6765,N_167,N_697);
or U6766 (N_6766,N_291,N_700);
nand U6767 (N_6767,N_3839,N_1009);
or U6768 (N_6768,N_1337,N_2087);
xnor U6769 (N_6769,N_1996,N_269);
nor U6770 (N_6770,N_1523,N_3694);
xor U6771 (N_6771,N_3109,N_2262);
nor U6772 (N_6772,N_2736,N_36);
and U6773 (N_6773,N_1299,N_2074);
xor U6774 (N_6774,N_1484,N_1044);
and U6775 (N_6775,N_2650,N_1669);
xnor U6776 (N_6776,N_1786,N_2000);
nand U6777 (N_6777,N_2929,N_3862);
or U6778 (N_6778,N_3403,N_1437);
and U6779 (N_6779,N_133,N_1459);
nand U6780 (N_6780,N_2922,N_1155);
or U6781 (N_6781,N_1755,N_3122);
nor U6782 (N_6782,N_975,N_3659);
and U6783 (N_6783,N_134,N_1486);
xor U6784 (N_6784,N_1316,N_1375);
nor U6785 (N_6785,N_1403,N_2548);
xnor U6786 (N_6786,N_2207,N_844);
or U6787 (N_6787,N_1535,N_3246);
xnor U6788 (N_6788,N_3787,N_232);
nand U6789 (N_6789,N_2869,N_1206);
nand U6790 (N_6790,N_3309,N_2120);
and U6791 (N_6791,N_347,N_3729);
and U6792 (N_6792,N_1177,N_2389);
or U6793 (N_6793,N_197,N_3041);
xor U6794 (N_6794,N_1456,N_348);
nand U6795 (N_6795,N_1814,N_2816);
nor U6796 (N_6796,N_3237,N_2803);
or U6797 (N_6797,N_3653,N_991);
nand U6798 (N_6798,N_1839,N_2366);
or U6799 (N_6799,N_927,N_2438);
nand U6800 (N_6800,N_3687,N_1110);
nand U6801 (N_6801,N_3218,N_612);
nor U6802 (N_6802,N_891,N_427);
and U6803 (N_6803,N_2738,N_2957);
xnor U6804 (N_6804,N_571,N_652);
and U6805 (N_6805,N_829,N_1124);
nor U6806 (N_6806,N_432,N_2830);
xnor U6807 (N_6807,N_2294,N_3403);
or U6808 (N_6808,N_1036,N_3534);
or U6809 (N_6809,N_3238,N_3802);
nor U6810 (N_6810,N_882,N_379);
and U6811 (N_6811,N_150,N_993);
or U6812 (N_6812,N_264,N_1977);
and U6813 (N_6813,N_1396,N_3602);
nor U6814 (N_6814,N_661,N_3644);
nand U6815 (N_6815,N_2603,N_1423);
or U6816 (N_6816,N_3766,N_132);
xnor U6817 (N_6817,N_2314,N_2794);
and U6818 (N_6818,N_1875,N_1991);
nand U6819 (N_6819,N_2634,N_2589);
xor U6820 (N_6820,N_3441,N_197);
nand U6821 (N_6821,N_1311,N_1702);
or U6822 (N_6822,N_2082,N_253);
and U6823 (N_6823,N_869,N_2270);
and U6824 (N_6824,N_1152,N_3950);
nor U6825 (N_6825,N_237,N_2604);
nor U6826 (N_6826,N_2596,N_2481);
nand U6827 (N_6827,N_2011,N_2769);
or U6828 (N_6828,N_1773,N_1584);
or U6829 (N_6829,N_300,N_3454);
nor U6830 (N_6830,N_2540,N_3349);
or U6831 (N_6831,N_1714,N_3277);
or U6832 (N_6832,N_2718,N_1898);
and U6833 (N_6833,N_3013,N_6);
nor U6834 (N_6834,N_1491,N_645);
nor U6835 (N_6835,N_524,N_2313);
xnor U6836 (N_6836,N_1862,N_2594);
nor U6837 (N_6837,N_2939,N_3674);
nor U6838 (N_6838,N_2485,N_2440);
or U6839 (N_6839,N_2989,N_520);
and U6840 (N_6840,N_661,N_3442);
and U6841 (N_6841,N_2564,N_3007);
nand U6842 (N_6842,N_464,N_3311);
nor U6843 (N_6843,N_756,N_3032);
or U6844 (N_6844,N_3020,N_1735);
xnor U6845 (N_6845,N_1124,N_2277);
and U6846 (N_6846,N_782,N_179);
nand U6847 (N_6847,N_2183,N_1615);
nor U6848 (N_6848,N_3317,N_819);
nor U6849 (N_6849,N_445,N_1489);
and U6850 (N_6850,N_1347,N_510);
nor U6851 (N_6851,N_2941,N_1710);
nand U6852 (N_6852,N_3331,N_1909);
nor U6853 (N_6853,N_1758,N_2413);
nand U6854 (N_6854,N_1785,N_3478);
nand U6855 (N_6855,N_626,N_240);
nand U6856 (N_6856,N_1425,N_1272);
nor U6857 (N_6857,N_561,N_3394);
nor U6858 (N_6858,N_3152,N_3572);
xnor U6859 (N_6859,N_3389,N_2908);
nor U6860 (N_6860,N_1486,N_2231);
nor U6861 (N_6861,N_3557,N_2055);
or U6862 (N_6862,N_1893,N_2906);
or U6863 (N_6863,N_1017,N_1738);
xor U6864 (N_6864,N_746,N_2332);
nor U6865 (N_6865,N_1510,N_1630);
nand U6866 (N_6866,N_950,N_3900);
xor U6867 (N_6867,N_686,N_1587);
nor U6868 (N_6868,N_307,N_1993);
and U6869 (N_6869,N_2664,N_1953);
and U6870 (N_6870,N_1757,N_3625);
nor U6871 (N_6871,N_1022,N_1283);
and U6872 (N_6872,N_493,N_240);
nand U6873 (N_6873,N_2353,N_1020);
nand U6874 (N_6874,N_358,N_1466);
nor U6875 (N_6875,N_65,N_1193);
and U6876 (N_6876,N_3850,N_98);
nor U6877 (N_6877,N_2556,N_3535);
xnor U6878 (N_6878,N_1153,N_355);
nor U6879 (N_6879,N_461,N_1329);
xnor U6880 (N_6880,N_3073,N_2825);
and U6881 (N_6881,N_2677,N_2120);
or U6882 (N_6882,N_2765,N_1301);
xnor U6883 (N_6883,N_1267,N_2656);
xnor U6884 (N_6884,N_837,N_3908);
or U6885 (N_6885,N_572,N_2645);
nand U6886 (N_6886,N_3397,N_1832);
nand U6887 (N_6887,N_2923,N_2124);
nand U6888 (N_6888,N_3103,N_664);
and U6889 (N_6889,N_2484,N_3043);
nand U6890 (N_6890,N_350,N_385);
nor U6891 (N_6891,N_280,N_3549);
or U6892 (N_6892,N_1910,N_3033);
nor U6893 (N_6893,N_716,N_1027);
xnor U6894 (N_6894,N_1101,N_815);
and U6895 (N_6895,N_3949,N_13);
or U6896 (N_6896,N_2711,N_2101);
nand U6897 (N_6897,N_1095,N_1527);
or U6898 (N_6898,N_2051,N_1399);
nand U6899 (N_6899,N_3267,N_2291);
nand U6900 (N_6900,N_1166,N_1049);
nor U6901 (N_6901,N_3060,N_3900);
or U6902 (N_6902,N_1796,N_2867);
xnor U6903 (N_6903,N_1957,N_3669);
xor U6904 (N_6904,N_2324,N_2801);
xnor U6905 (N_6905,N_3465,N_2501);
nand U6906 (N_6906,N_3997,N_759);
or U6907 (N_6907,N_3020,N_3614);
nor U6908 (N_6908,N_2060,N_3303);
or U6909 (N_6909,N_2619,N_287);
xnor U6910 (N_6910,N_1320,N_1607);
nor U6911 (N_6911,N_1195,N_2926);
and U6912 (N_6912,N_2774,N_2336);
xnor U6913 (N_6913,N_807,N_3680);
nand U6914 (N_6914,N_1434,N_3735);
or U6915 (N_6915,N_2646,N_3307);
nor U6916 (N_6916,N_3800,N_897);
xor U6917 (N_6917,N_1826,N_3296);
xor U6918 (N_6918,N_2276,N_3813);
or U6919 (N_6919,N_1653,N_390);
xor U6920 (N_6920,N_1917,N_3662);
and U6921 (N_6921,N_964,N_38);
xor U6922 (N_6922,N_900,N_60);
nand U6923 (N_6923,N_1734,N_2250);
nor U6924 (N_6924,N_2395,N_665);
nand U6925 (N_6925,N_1361,N_3542);
xor U6926 (N_6926,N_2788,N_1492);
nor U6927 (N_6927,N_2992,N_254);
and U6928 (N_6928,N_479,N_584);
and U6929 (N_6929,N_1158,N_2118);
nor U6930 (N_6930,N_204,N_3959);
or U6931 (N_6931,N_523,N_371);
nor U6932 (N_6932,N_3778,N_243);
or U6933 (N_6933,N_3821,N_31);
and U6934 (N_6934,N_3714,N_2805);
or U6935 (N_6935,N_3242,N_384);
nor U6936 (N_6936,N_1067,N_2460);
or U6937 (N_6937,N_3023,N_874);
or U6938 (N_6938,N_1330,N_3032);
and U6939 (N_6939,N_3537,N_3193);
xnor U6940 (N_6940,N_1900,N_3705);
and U6941 (N_6941,N_1032,N_573);
nand U6942 (N_6942,N_2138,N_3935);
xnor U6943 (N_6943,N_1473,N_732);
xnor U6944 (N_6944,N_2528,N_92);
nor U6945 (N_6945,N_3590,N_3712);
and U6946 (N_6946,N_3282,N_3355);
or U6947 (N_6947,N_2660,N_1339);
nor U6948 (N_6948,N_992,N_2198);
nor U6949 (N_6949,N_3770,N_1953);
nor U6950 (N_6950,N_3197,N_3127);
and U6951 (N_6951,N_101,N_2790);
and U6952 (N_6952,N_3937,N_1855);
xnor U6953 (N_6953,N_3804,N_2864);
nand U6954 (N_6954,N_1505,N_1876);
or U6955 (N_6955,N_3656,N_3665);
or U6956 (N_6956,N_2121,N_3292);
and U6957 (N_6957,N_2712,N_2224);
and U6958 (N_6958,N_146,N_3900);
xor U6959 (N_6959,N_2077,N_912);
or U6960 (N_6960,N_1797,N_1511);
or U6961 (N_6961,N_3346,N_3404);
nand U6962 (N_6962,N_1788,N_2744);
and U6963 (N_6963,N_2462,N_3501);
nand U6964 (N_6964,N_2817,N_187);
and U6965 (N_6965,N_1369,N_3011);
nand U6966 (N_6966,N_2897,N_349);
nand U6967 (N_6967,N_337,N_757);
nand U6968 (N_6968,N_1433,N_1209);
or U6969 (N_6969,N_2396,N_3242);
or U6970 (N_6970,N_3207,N_1486);
nand U6971 (N_6971,N_719,N_2839);
nand U6972 (N_6972,N_3030,N_2347);
xor U6973 (N_6973,N_3361,N_1287);
and U6974 (N_6974,N_727,N_3654);
nor U6975 (N_6975,N_2920,N_2018);
xnor U6976 (N_6976,N_2485,N_2861);
xor U6977 (N_6977,N_3399,N_1344);
or U6978 (N_6978,N_868,N_632);
or U6979 (N_6979,N_1956,N_2226);
xnor U6980 (N_6980,N_891,N_3581);
nand U6981 (N_6981,N_1241,N_333);
nor U6982 (N_6982,N_35,N_3490);
xor U6983 (N_6983,N_2913,N_1892);
xnor U6984 (N_6984,N_3332,N_2325);
or U6985 (N_6985,N_2004,N_1807);
and U6986 (N_6986,N_3427,N_2217);
nor U6987 (N_6987,N_2795,N_2356);
and U6988 (N_6988,N_3730,N_2800);
nand U6989 (N_6989,N_1259,N_494);
xor U6990 (N_6990,N_224,N_287);
or U6991 (N_6991,N_3292,N_1838);
or U6992 (N_6992,N_173,N_3991);
and U6993 (N_6993,N_1943,N_463);
nor U6994 (N_6994,N_2157,N_1529);
xor U6995 (N_6995,N_1944,N_3462);
nand U6996 (N_6996,N_2434,N_3167);
nand U6997 (N_6997,N_3834,N_3430);
nor U6998 (N_6998,N_3986,N_3218);
or U6999 (N_6999,N_2879,N_2556);
and U7000 (N_7000,N_3729,N_1533);
nand U7001 (N_7001,N_2492,N_972);
or U7002 (N_7002,N_366,N_2444);
nand U7003 (N_7003,N_1591,N_1117);
nand U7004 (N_7004,N_3022,N_3704);
nand U7005 (N_7005,N_2019,N_244);
or U7006 (N_7006,N_2793,N_358);
xor U7007 (N_7007,N_3104,N_1240);
or U7008 (N_7008,N_226,N_1723);
and U7009 (N_7009,N_1738,N_3706);
xnor U7010 (N_7010,N_999,N_2144);
xnor U7011 (N_7011,N_1952,N_2139);
or U7012 (N_7012,N_1142,N_2468);
nor U7013 (N_7013,N_3070,N_2117);
nor U7014 (N_7014,N_731,N_2621);
or U7015 (N_7015,N_2827,N_2008);
or U7016 (N_7016,N_2947,N_3243);
or U7017 (N_7017,N_2915,N_2440);
nand U7018 (N_7018,N_2717,N_1556);
nand U7019 (N_7019,N_1471,N_2947);
or U7020 (N_7020,N_3513,N_3946);
and U7021 (N_7021,N_384,N_1831);
nand U7022 (N_7022,N_3217,N_3223);
nor U7023 (N_7023,N_3406,N_3146);
nand U7024 (N_7024,N_1671,N_3958);
and U7025 (N_7025,N_3885,N_1942);
nor U7026 (N_7026,N_2870,N_1573);
xnor U7027 (N_7027,N_3361,N_1654);
nor U7028 (N_7028,N_2445,N_3844);
or U7029 (N_7029,N_2581,N_1883);
nor U7030 (N_7030,N_346,N_2984);
and U7031 (N_7031,N_1980,N_96);
nand U7032 (N_7032,N_693,N_1430);
and U7033 (N_7033,N_3070,N_1965);
nand U7034 (N_7034,N_1899,N_293);
and U7035 (N_7035,N_3926,N_1470);
xor U7036 (N_7036,N_1523,N_3354);
nor U7037 (N_7037,N_1024,N_3161);
nand U7038 (N_7038,N_901,N_1073);
or U7039 (N_7039,N_1468,N_2619);
nand U7040 (N_7040,N_2297,N_921);
and U7041 (N_7041,N_3069,N_3151);
or U7042 (N_7042,N_2331,N_3739);
or U7043 (N_7043,N_1282,N_1281);
xnor U7044 (N_7044,N_105,N_2162);
nor U7045 (N_7045,N_3837,N_626);
nand U7046 (N_7046,N_983,N_2150);
xor U7047 (N_7047,N_2305,N_3087);
xor U7048 (N_7048,N_1151,N_209);
nor U7049 (N_7049,N_1822,N_3722);
and U7050 (N_7050,N_1196,N_319);
nor U7051 (N_7051,N_2222,N_2658);
xnor U7052 (N_7052,N_3705,N_2617);
nor U7053 (N_7053,N_1943,N_674);
nand U7054 (N_7054,N_92,N_3941);
and U7055 (N_7055,N_2148,N_408);
and U7056 (N_7056,N_3982,N_3852);
or U7057 (N_7057,N_3590,N_924);
or U7058 (N_7058,N_3450,N_1001);
nor U7059 (N_7059,N_3550,N_2426);
and U7060 (N_7060,N_1569,N_3162);
and U7061 (N_7061,N_1738,N_458);
nand U7062 (N_7062,N_1534,N_1564);
nor U7063 (N_7063,N_2737,N_883);
and U7064 (N_7064,N_3152,N_3191);
nand U7065 (N_7065,N_1444,N_163);
nand U7066 (N_7066,N_219,N_2904);
nor U7067 (N_7067,N_3220,N_3810);
nor U7068 (N_7068,N_1118,N_2116);
and U7069 (N_7069,N_1774,N_2626);
or U7070 (N_7070,N_1477,N_1152);
xnor U7071 (N_7071,N_2784,N_3902);
xor U7072 (N_7072,N_1535,N_3371);
nor U7073 (N_7073,N_549,N_3707);
nand U7074 (N_7074,N_1919,N_2891);
nor U7075 (N_7075,N_2309,N_3800);
nand U7076 (N_7076,N_483,N_3285);
and U7077 (N_7077,N_3466,N_3418);
xnor U7078 (N_7078,N_3101,N_3142);
xor U7079 (N_7079,N_3436,N_2977);
or U7080 (N_7080,N_3668,N_3503);
nor U7081 (N_7081,N_2970,N_2107);
nor U7082 (N_7082,N_3795,N_2685);
nor U7083 (N_7083,N_3394,N_1948);
nand U7084 (N_7084,N_1957,N_2244);
nand U7085 (N_7085,N_3781,N_1141);
xnor U7086 (N_7086,N_3716,N_3053);
nor U7087 (N_7087,N_501,N_244);
xnor U7088 (N_7088,N_2658,N_1328);
xor U7089 (N_7089,N_3764,N_884);
nor U7090 (N_7090,N_1756,N_803);
nor U7091 (N_7091,N_3673,N_2096);
or U7092 (N_7092,N_3966,N_3665);
xnor U7093 (N_7093,N_3855,N_938);
nand U7094 (N_7094,N_88,N_729);
nor U7095 (N_7095,N_3768,N_718);
and U7096 (N_7096,N_2803,N_3928);
and U7097 (N_7097,N_3569,N_214);
nand U7098 (N_7098,N_1259,N_2061);
nand U7099 (N_7099,N_3154,N_2560);
nand U7100 (N_7100,N_2964,N_2279);
nor U7101 (N_7101,N_2556,N_3497);
nor U7102 (N_7102,N_2538,N_2236);
nor U7103 (N_7103,N_2966,N_2849);
or U7104 (N_7104,N_1923,N_1594);
and U7105 (N_7105,N_254,N_3672);
xnor U7106 (N_7106,N_3458,N_958);
or U7107 (N_7107,N_169,N_1119);
xor U7108 (N_7108,N_2867,N_3041);
xor U7109 (N_7109,N_1821,N_1315);
and U7110 (N_7110,N_228,N_424);
or U7111 (N_7111,N_2306,N_735);
xnor U7112 (N_7112,N_1346,N_403);
xnor U7113 (N_7113,N_2485,N_1145);
xnor U7114 (N_7114,N_3491,N_3641);
and U7115 (N_7115,N_981,N_3238);
nor U7116 (N_7116,N_2509,N_104);
nand U7117 (N_7117,N_3468,N_3084);
nor U7118 (N_7118,N_3026,N_199);
and U7119 (N_7119,N_3608,N_2989);
or U7120 (N_7120,N_3071,N_2621);
and U7121 (N_7121,N_2704,N_517);
nor U7122 (N_7122,N_3483,N_2290);
and U7123 (N_7123,N_209,N_3371);
nor U7124 (N_7124,N_3688,N_1770);
or U7125 (N_7125,N_2968,N_343);
nor U7126 (N_7126,N_631,N_82);
xnor U7127 (N_7127,N_1734,N_2592);
or U7128 (N_7128,N_822,N_3825);
xor U7129 (N_7129,N_2694,N_1092);
and U7130 (N_7130,N_1745,N_384);
nor U7131 (N_7131,N_447,N_3692);
xor U7132 (N_7132,N_595,N_3237);
or U7133 (N_7133,N_947,N_1140);
or U7134 (N_7134,N_1401,N_353);
and U7135 (N_7135,N_1480,N_769);
or U7136 (N_7136,N_1784,N_560);
or U7137 (N_7137,N_903,N_3318);
or U7138 (N_7138,N_2163,N_846);
or U7139 (N_7139,N_2030,N_2241);
and U7140 (N_7140,N_2284,N_2192);
and U7141 (N_7141,N_890,N_1971);
nand U7142 (N_7142,N_3024,N_1884);
nor U7143 (N_7143,N_1734,N_999);
xnor U7144 (N_7144,N_2959,N_2207);
and U7145 (N_7145,N_2755,N_3205);
nand U7146 (N_7146,N_1289,N_490);
nor U7147 (N_7147,N_2389,N_1464);
nor U7148 (N_7148,N_618,N_1831);
or U7149 (N_7149,N_1654,N_1425);
nor U7150 (N_7150,N_2787,N_80);
nor U7151 (N_7151,N_1759,N_522);
and U7152 (N_7152,N_2715,N_2950);
or U7153 (N_7153,N_1245,N_1405);
nor U7154 (N_7154,N_3450,N_2774);
nor U7155 (N_7155,N_2052,N_3990);
nor U7156 (N_7156,N_2018,N_3730);
nor U7157 (N_7157,N_1962,N_3813);
nor U7158 (N_7158,N_561,N_2963);
nand U7159 (N_7159,N_1806,N_96);
nor U7160 (N_7160,N_515,N_2422);
xor U7161 (N_7161,N_1482,N_566);
xnor U7162 (N_7162,N_3880,N_3721);
nor U7163 (N_7163,N_3480,N_2865);
xor U7164 (N_7164,N_1724,N_3336);
or U7165 (N_7165,N_479,N_700);
nand U7166 (N_7166,N_1045,N_705);
nor U7167 (N_7167,N_980,N_2745);
and U7168 (N_7168,N_22,N_823);
and U7169 (N_7169,N_3341,N_3132);
and U7170 (N_7170,N_269,N_211);
nor U7171 (N_7171,N_1897,N_1609);
nor U7172 (N_7172,N_44,N_3095);
and U7173 (N_7173,N_1146,N_3784);
xor U7174 (N_7174,N_2729,N_1127);
nand U7175 (N_7175,N_568,N_2500);
nor U7176 (N_7176,N_1209,N_1250);
nor U7177 (N_7177,N_923,N_3709);
nor U7178 (N_7178,N_929,N_2065);
nor U7179 (N_7179,N_21,N_1437);
nand U7180 (N_7180,N_3781,N_917);
and U7181 (N_7181,N_1204,N_2011);
and U7182 (N_7182,N_1907,N_2564);
or U7183 (N_7183,N_824,N_2456);
or U7184 (N_7184,N_2411,N_2652);
xnor U7185 (N_7185,N_2293,N_3765);
or U7186 (N_7186,N_1108,N_1008);
nor U7187 (N_7187,N_3298,N_3071);
or U7188 (N_7188,N_2751,N_2104);
nand U7189 (N_7189,N_1523,N_2666);
nor U7190 (N_7190,N_1243,N_3415);
xnor U7191 (N_7191,N_2585,N_1221);
and U7192 (N_7192,N_1944,N_3744);
or U7193 (N_7193,N_3605,N_2771);
and U7194 (N_7194,N_1455,N_1563);
or U7195 (N_7195,N_3837,N_837);
nor U7196 (N_7196,N_223,N_1126);
nor U7197 (N_7197,N_3744,N_2707);
nand U7198 (N_7198,N_702,N_477);
nor U7199 (N_7199,N_3887,N_1837);
nor U7200 (N_7200,N_1439,N_883);
and U7201 (N_7201,N_793,N_1408);
nor U7202 (N_7202,N_1088,N_3991);
nor U7203 (N_7203,N_3405,N_977);
nor U7204 (N_7204,N_803,N_2959);
nand U7205 (N_7205,N_3532,N_1987);
nand U7206 (N_7206,N_1885,N_753);
or U7207 (N_7207,N_2663,N_3234);
nand U7208 (N_7208,N_3225,N_2637);
xor U7209 (N_7209,N_3775,N_1921);
nand U7210 (N_7210,N_3403,N_1676);
xnor U7211 (N_7211,N_1840,N_559);
nor U7212 (N_7212,N_1173,N_835);
xor U7213 (N_7213,N_3343,N_2511);
xnor U7214 (N_7214,N_1750,N_3516);
nand U7215 (N_7215,N_1275,N_574);
and U7216 (N_7216,N_2444,N_535);
nand U7217 (N_7217,N_1371,N_3711);
xor U7218 (N_7218,N_3585,N_1017);
nor U7219 (N_7219,N_106,N_2210);
nand U7220 (N_7220,N_1889,N_3323);
and U7221 (N_7221,N_842,N_1169);
nand U7222 (N_7222,N_3773,N_3441);
nand U7223 (N_7223,N_1733,N_3099);
nand U7224 (N_7224,N_3970,N_1789);
xnor U7225 (N_7225,N_1916,N_2646);
xor U7226 (N_7226,N_2448,N_1800);
or U7227 (N_7227,N_3518,N_450);
nand U7228 (N_7228,N_2960,N_2607);
and U7229 (N_7229,N_1868,N_2583);
and U7230 (N_7230,N_3278,N_2998);
nor U7231 (N_7231,N_2553,N_1799);
and U7232 (N_7232,N_3754,N_1241);
or U7233 (N_7233,N_3708,N_2578);
xnor U7234 (N_7234,N_2950,N_2972);
nand U7235 (N_7235,N_436,N_1005);
or U7236 (N_7236,N_3948,N_252);
and U7237 (N_7237,N_3089,N_3805);
nor U7238 (N_7238,N_78,N_459);
nor U7239 (N_7239,N_2730,N_1031);
nor U7240 (N_7240,N_689,N_240);
nand U7241 (N_7241,N_3177,N_1483);
nor U7242 (N_7242,N_1039,N_3154);
xor U7243 (N_7243,N_1245,N_20);
and U7244 (N_7244,N_1083,N_2730);
or U7245 (N_7245,N_3156,N_824);
and U7246 (N_7246,N_3508,N_2818);
and U7247 (N_7247,N_3819,N_3112);
nand U7248 (N_7248,N_3434,N_874);
nor U7249 (N_7249,N_2252,N_2385);
nand U7250 (N_7250,N_404,N_813);
or U7251 (N_7251,N_1125,N_569);
nand U7252 (N_7252,N_2347,N_3368);
nand U7253 (N_7253,N_3976,N_240);
xnor U7254 (N_7254,N_1657,N_2803);
and U7255 (N_7255,N_2064,N_807);
and U7256 (N_7256,N_3528,N_903);
xor U7257 (N_7257,N_3901,N_3709);
nand U7258 (N_7258,N_653,N_551);
and U7259 (N_7259,N_872,N_3577);
xnor U7260 (N_7260,N_725,N_648);
nor U7261 (N_7261,N_3285,N_3841);
nor U7262 (N_7262,N_1341,N_2281);
nor U7263 (N_7263,N_3579,N_1584);
or U7264 (N_7264,N_3880,N_1035);
or U7265 (N_7265,N_1181,N_921);
or U7266 (N_7266,N_3942,N_959);
and U7267 (N_7267,N_3014,N_2740);
nand U7268 (N_7268,N_93,N_2534);
nand U7269 (N_7269,N_971,N_794);
xnor U7270 (N_7270,N_3586,N_3270);
and U7271 (N_7271,N_742,N_1308);
or U7272 (N_7272,N_3610,N_3775);
nand U7273 (N_7273,N_221,N_984);
or U7274 (N_7274,N_1488,N_2839);
nand U7275 (N_7275,N_918,N_2864);
nor U7276 (N_7276,N_3619,N_36);
xor U7277 (N_7277,N_2412,N_3835);
nand U7278 (N_7278,N_109,N_765);
nor U7279 (N_7279,N_3649,N_2638);
xor U7280 (N_7280,N_2011,N_2152);
nand U7281 (N_7281,N_1752,N_3097);
xor U7282 (N_7282,N_2302,N_3894);
nand U7283 (N_7283,N_630,N_3848);
and U7284 (N_7284,N_2662,N_981);
nand U7285 (N_7285,N_3066,N_997);
and U7286 (N_7286,N_1721,N_891);
nand U7287 (N_7287,N_1614,N_2527);
and U7288 (N_7288,N_2241,N_2506);
and U7289 (N_7289,N_927,N_1713);
xor U7290 (N_7290,N_891,N_1005);
and U7291 (N_7291,N_3093,N_2248);
or U7292 (N_7292,N_2441,N_3455);
and U7293 (N_7293,N_3658,N_3608);
and U7294 (N_7294,N_2006,N_1364);
or U7295 (N_7295,N_3126,N_3976);
and U7296 (N_7296,N_2296,N_2272);
and U7297 (N_7297,N_1924,N_1601);
nand U7298 (N_7298,N_1351,N_3968);
or U7299 (N_7299,N_3181,N_1286);
nor U7300 (N_7300,N_2294,N_2104);
xor U7301 (N_7301,N_1186,N_1616);
nor U7302 (N_7302,N_558,N_1773);
nor U7303 (N_7303,N_489,N_677);
nor U7304 (N_7304,N_1927,N_225);
and U7305 (N_7305,N_3728,N_2626);
nor U7306 (N_7306,N_981,N_3869);
nand U7307 (N_7307,N_654,N_58);
xnor U7308 (N_7308,N_2205,N_1231);
xor U7309 (N_7309,N_639,N_124);
or U7310 (N_7310,N_3663,N_3376);
nand U7311 (N_7311,N_2479,N_875);
xnor U7312 (N_7312,N_3604,N_2237);
nand U7313 (N_7313,N_1373,N_1055);
nand U7314 (N_7314,N_1794,N_2052);
nor U7315 (N_7315,N_2223,N_2919);
nand U7316 (N_7316,N_1151,N_3635);
or U7317 (N_7317,N_3368,N_3321);
and U7318 (N_7318,N_3339,N_2659);
xnor U7319 (N_7319,N_1279,N_387);
nand U7320 (N_7320,N_2642,N_788);
nor U7321 (N_7321,N_3495,N_3042);
and U7322 (N_7322,N_1627,N_2353);
nor U7323 (N_7323,N_1318,N_892);
xnor U7324 (N_7324,N_994,N_1562);
xor U7325 (N_7325,N_3766,N_1155);
nand U7326 (N_7326,N_2732,N_2132);
nor U7327 (N_7327,N_889,N_3697);
and U7328 (N_7328,N_2015,N_3659);
xor U7329 (N_7329,N_1554,N_3139);
nor U7330 (N_7330,N_486,N_2878);
and U7331 (N_7331,N_1980,N_1562);
nand U7332 (N_7332,N_2595,N_3764);
nand U7333 (N_7333,N_238,N_2749);
nor U7334 (N_7334,N_2579,N_407);
xnor U7335 (N_7335,N_1527,N_1606);
nand U7336 (N_7336,N_260,N_1650);
and U7337 (N_7337,N_532,N_1830);
and U7338 (N_7338,N_849,N_770);
nand U7339 (N_7339,N_3538,N_960);
nand U7340 (N_7340,N_3120,N_3646);
xor U7341 (N_7341,N_2703,N_1625);
nand U7342 (N_7342,N_938,N_2702);
or U7343 (N_7343,N_2959,N_3480);
nor U7344 (N_7344,N_2722,N_1281);
or U7345 (N_7345,N_1753,N_862);
nand U7346 (N_7346,N_1198,N_2529);
xor U7347 (N_7347,N_3373,N_2869);
or U7348 (N_7348,N_1498,N_921);
and U7349 (N_7349,N_3973,N_3939);
xor U7350 (N_7350,N_2425,N_3654);
or U7351 (N_7351,N_2730,N_491);
and U7352 (N_7352,N_2454,N_688);
or U7353 (N_7353,N_248,N_3996);
xor U7354 (N_7354,N_3525,N_1225);
nand U7355 (N_7355,N_911,N_972);
xnor U7356 (N_7356,N_2745,N_1300);
nor U7357 (N_7357,N_292,N_896);
or U7358 (N_7358,N_1352,N_3444);
xnor U7359 (N_7359,N_2834,N_438);
and U7360 (N_7360,N_370,N_2613);
xnor U7361 (N_7361,N_3351,N_280);
nand U7362 (N_7362,N_2914,N_78);
or U7363 (N_7363,N_1355,N_613);
and U7364 (N_7364,N_2808,N_3948);
nor U7365 (N_7365,N_1590,N_3482);
or U7366 (N_7366,N_1737,N_2341);
or U7367 (N_7367,N_1770,N_1118);
xor U7368 (N_7368,N_73,N_522);
xnor U7369 (N_7369,N_1054,N_1682);
nand U7370 (N_7370,N_686,N_1159);
nor U7371 (N_7371,N_64,N_935);
and U7372 (N_7372,N_1473,N_3240);
nor U7373 (N_7373,N_3927,N_359);
nand U7374 (N_7374,N_19,N_2852);
nand U7375 (N_7375,N_1452,N_2625);
xor U7376 (N_7376,N_82,N_1860);
and U7377 (N_7377,N_2037,N_3037);
nand U7378 (N_7378,N_286,N_1595);
xnor U7379 (N_7379,N_2759,N_2203);
nand U7380 (N_7380,N_3174,N_1919);
nor U7381 (N_7381,N_564,N_3627);
nand U7382 (N_7382,N_2934,N_99);
nand U7383 (N_7383,N_3651,N_1335);
nand U7384 (N_7384,N_3155,N_1843);
xnor U7385 (N_7385,N_3076,N_527);
nand U7386 (N_7386,N_3856,N_2385);
xnor U7387 (N_7387,N_508,N_2729);
nor U7388 (N_7388,N_1670,N_2305);
and U7389 (N_7389,N_901,N_1801);
xnor U7390 (N_7390,N_294,N_2810);
and U7391 (N_7391,N_2613,N_318);
or U7392 (N_7392,N_2846,N_2336);
nand U7393 (N_7393,N_1053,N_3405);
nor U7394 (N_7394,N_908,N_3789);
xnor U7395 (N_7395,N_854,N_1073);
xnor U7396 (N_7396,N_1393,N_3924);
xnor U7397 (N_7397,N_280,N_950);
and U7398 (N_7398,N_1947,N_3645);
and U7399 (N_7399,N_1702,N_3121);
nand U7400 (N_7400,N_3413,N_1303);
nand U7401 (N_7401,N_3821,N_3473);
nor U7402 (N_7402,N_1718,N_2581);
and U7403 (N_7403,N_2739,N_2878);
or U7404 (N_7404,N_692,N_3105);
nand U7405 (N_7405,N_2647,N_3120);
xor U7406 (N_7406,N_2502,N_2752);
nor U7407 (N_7407,N_3968,N_3681);
nand U7408 (N_7408,N_682,N_2308);
xnor U7409 (N_7409,N_793,N_835);
xor U7410 (N_7410,N_1819,N_3763);
and U7411 (N_7411,N_588,N_3508);
nand U7412 (N_7412,N_2254,N_2916);
and U7413 (N_7413,N_3854,N_2732);
and U7414 (N_7414,N_1978,N_100);
nor U7415 (N_7415,N_3359,N_497);
nor U7416 (N_7416,N_3083,N_2280);
or U7417 (N_7417,N_660,N_3160);
nand U7418 (N_7418,N_3389,N_3844);
nand U7419 (N_7419,N_1856,N_125);
nor U7420 (N_7420,N_220,N_3494);
nand U7421 (N_7421,N_558,N_3391);
nand U7422 (N_7422,N_2250,N_1496);
or U7423 (N_7423,N_2072,N_1667);
and U7424 (N_7424,N_1739,N_293);
nand U7425 (N_7425,N_104,N_2062);
nand U7426 (N_7426,N_1781,N_3783);
nor U7427 (N_7427,N_2603,N_543);
nand U7428 (N_7428,N_3292,N_426);
nand U7429 (N_7429,N_816,N_1833);
nor U7430 (N_7430,N_12,N_3906);
and U7431 (N_7431,N_999,N_93);
nor U7432 (N_7432,N_3652,N_1585);
nand U7433 (N_7433,N_1311,N_3810);
and U7434 (N_7434,N_3253,N_2984);
xor U7435 (N_7435,N_2021,N_1407);
nand U7436 (N_7436,N_3284,N_1627);
xor U7437 (N_7437,N_1316,N_1516);
or U7438 (N_7438,N_731,N_521);
nor U7439 (N_7439,N_3796,N_2021);
xnor U7440 (N_7440,N_286,N_4);
or U7441 (N_7441,N_2154,N_2548);
or U7442 (N_7442,N_3497,N_3827);
or U7443 (N_7443,N_306,N_1215);
nor U7444 (N_7444,N_3671,N_2120);
and U7445 (N_7445,N_2259,N_688);
xnor U7446 (N_7446,N_635,N_319);
nand U7447 (N_7447,N_1345,N_3685);
and U7448 (N_7448,N_375,N_48);
nand U7449 (N_7449,N_53,N_1037);
nor U7450 (N_7450,N_298,N_1728);
xor U7451 (N_7451,N_3590,N_2976);
xor U7452 (N_7452,N_2273,N_2525);
nand U7453 (N_7453,N_1077,N_2785);
nand U7454 (N_7454,N_2151,N_3182);
and U7455 (N_7455,N_67,N_1691);
xnor U7456 (N_7456,N_3544,N_1701);
nor U7457 (N_7457,N_1091,N_3414);
and U7458 (N_7458,N_987,N_2932);
nor U7459 (N_7459,N_2394,N_1097);
and U7460 (N_7460,N_1126,N_2170);
nor U7461 (N_7461,N_3818,N_330);
nor U7462 (N_7462,N_343,N_2141);
nand U7463 (N_7463,N_1025,N_3326);
nor U7464 (N_7464,N_3473,N_1187);
or U7465 (N_7465,N_480,N_3433);
nor U7466 (N_7466,N_1228,N_1162);
xnor U7467 (N_7467,N_633,N_2409);
nor U7468 (N_7468,N_1342,N_1005);
and U7469 (N_7469,N_3703,N_3989);
nor U7470 (N_7470,N_3915,N_2382);
or U7471 (N_7471,N_2313,N_2817);
nor U7472 (N_7472,N_3460,N_2332);
nor U7473 (N_7473,N_1164,N_1764);
or U7474 (N_7474,N_611,N_213);
nor U7475 (N_7475,N_3126,N_785);
or U7476 (N_7476,N_2803,N_144);
nor U7477 (N_7477,N_1378,N_3906);
and U7478 (N_7478,N_1959,N_2175);
nor U7479 (N_7479,N_1120,N_1690);
nand U7480 (N_7480,N_2376,N_3103);
nor U7481 (N_7481,N_3894,N_2143);
nand U7482 (N_7482,N_3860,N_956);
nor U7483 (N_7483,N_3299,N_2758);
xor U7484 (N_7484,N_1818,N_2705);
or U7485 (N_7485,N_2886,N_935);
nand U7486 (N_7486,N_733,N_3867);
nand U7487 (N_7487,N_894,N_164);
xor U7488 (N_7488,N_431,N_1050);
xnor U7489 (N_7489,N_3942,N_2581);
or U7490 (N_7490,N_3054,N_2295);
or U7491 (N_7491,N_630,N_1378);
nand U7492 (N_7492,N_2128,N_2341);
nand U7493 (N_7493,N_1938,N_2029);
nand U7494 (N_7494,N_3850,N_1352);
nor U7495 (N_7495,N_2811,N_1522);
nor U7496 (N_7496,N_3418,N_1834);
nor U7497 (N_7497,N_1462,N_3638);
nand U7498 (N_7498,N_1795,N_3920);
or U7499 (N_7499,N_1337,N_3266);
xnor U7500 (N_7500,N_2615,N_2010);
and U7501 (N_7501,N_3563,N_733);
or U7502 (N_7502,N_1024,N_2300);
xnor U7503 (N_7503,N_2622,N_3630);
nor U7504 (N_7504,N_508,N_717);
and U7505 (N_7505,N_549,N_3146);
xor U7506 (N_7506,N_446,N_1272);
nor U7507 (N_7507,N_3662,N_940);
nor U7508 (N_7508,N_1729,N_674);
xnor U7509 (N_7509,N_755,N_2835);
nor U7510 (N_7510,N_654,N_959);
nor U7511 (N_7511,N_338,N_2290);
nand U7512 (N_7512,N_2870,N_3794);
or U7513 (N_7513,N_2931,N_2826);
and U7514 (N_7514,N_203,N_2466);
xor U7515 (N_7515,N_2208,N_1680);
xor U7516 (N_7516,N_1456,N_1573);
or U7517 (N_7517,N_3967,N_542);
and U7518 (N_7518,N_3575,N_2276);
nor U7519 (N_7519,N_3514,N_533);
nor U7520 (N_7520,N_3118,N_1447);
or U7521 (N_7521,N_888,N_528);
or U7522 (N_7522,N_960,N_563);
nand U7523 (N_7523,N_2367,N_3989);
nor U7524 (N_7524,N_2018,N_3752);
nor U7525 (N_7525,N_1253,N_1760);
and U7526 (N_7526,N_2403,N_2508);
nand U7527 (N_7527,N_2668,N_2854);
xor U7528 (N_7528,N_1874,N_3250);
nand U7529 (N_7529,N_2366,N_1925);
nor U7530 (N_7530,N_2355,N_1265);
or U7531 (N_7531,N_962,N_72);
xor U7532 (N_7532,N_3708,N_1463);
nand U7533 (N_7533,N_666,N_3544);
or U7534 (N_7534,N_1044,N_3557);
or U7535 (N_7535,N_778,N_199);
and U7536 (N_7536,N_822,N_790);
xnor U7537 (N_7537,N_2418,N_2675);
nor U7538 (N_7538,N_2918,N_106);
xnor U7539 (N_7539,N_3165,N_2456);
xnor U7540 (N_7540,N_2630,N_3176);
nand U7541 (N_7541,N_3999,N_3548);
nor U7542 (N_7542,N_2569,N_3230);
and U7543 (N_7543,N_3493,N_637);
and U7544 (N_7544,N_1282,N_3034);
and U7545 (N_7545,N_3236,N_3880);
xor U7546 (N_7546,N_1456,N_3816);
or U7547 (N_7547,N_1729,N_2358);
or U7548 (N_7548,N_1371,N_1874);
nand U7549 (N_7549,N_1610,N_1235);
and U7550 (N_7550,N_3666,N_3715);
nor U7551 (N_7551,N_2828,N_914);
or U7552 (N_7552,N_1733,N_2068);
or U7553 (N_7553,N_3831,N_3385);
nor U7554 (N_7554,N_1977,N_3692);
nand U7555 (N_7555,N_2183,N_376);
xor U7556 (N_7556,N_1241,N_1831);
or U7557 (N_7557,N_3335,N_319);
nand U7558 (N_7558,N_3537,N_2832);
nand U7559 (N_7559,N_1916,N_2790);
xor U7560 (N_7560,N_2632,N_2451);
xor U7561 (N_7561,N_2030,N_1176);
or U7562 (N_7562,N_1940,N_3768);
or U7563 (N_7563,N_1996,N_2247);
nor U7564 (N_7564,N_2781,N_33);
nor U7565 (N_7565,N_863,N_1232);
xor U7566 (N_7566,N_1824,N_2945);
xor U7567 (N_7567,N_1823,N_3666);
xor U7568 (N_7568,N_1071,N_3120);
xnor U7569 (N_7569,N_1908,N_3565);
and U7570 (N_7570,N_944,N_2109);
and U7571 (N_7571,N_1787,N_459);
xor U7572 (N_7572,N_347,N_802);
nand U7573 (N_7573,N_1545,N_2153);
xnor U7574 (N_7574,N_886,N_2953);
or U7575 (N_7575,N_209,N_2844);
or U7576 (N_7576,N_1636,N_2128);
or U7577 (N_7577,N_109,N_3934);
and U7578 (N_7578,N_2525,N_911);
xor U7579 (N_7579,N_3550,N_2411);
nand U7580 (N_7580,N_3535,N_523);
xnor U7581 (N_7581,N_352,N_97);
and U7582 (N_7582,N_851,N_1330);
nor U7583 (N_7583,N_2710,N_3199);
or U7584 (N_7584,N_385,N_1447);
nand U7585 (N_7585,N_1608,N_2938);
nor U7586 (N_7586,N_1794,N_2799);
nand U7587 (N_7587,N_1474,N_1504);
nand U7588 (N_7588,N_1028,N_3964);
and U7589 (N_7589,N_505,N_3012);
and U7590 (N_7590,N_3717,N_3923);
xnor U7591 (N_7591,N_2113,N_3946);
and U7592 (N_7592,N_2472,N_1797);
nor U7593 (N_7593,N_94,N_2844);
xnor U7594 (N_7594,N_610,N_2890);
and U7595 (N_7595,N_1830,N_1158);
and U7596 (N_7596,N_1452,N_113);
or U7597 (N_7597,N_2847,N_1726);
and U7598 (N_7598,N_3741,N_3450);
or U7599 (N_7599,N_1828,N_3022);
xor U7600 (N_7600,N_2237,N_1588);
and U7601 (N_7601,N_3297,N_3123);
and U7602 (N_7602,N_199,N_388);
nand U7603 (N_7603,N_2290,N_3108);
nand U7604 (N_7604,N_2739,N_1869);
nand U7605 (N_7605,N_476,N_2714);
or U7606 (N_7606,N_213,N_2271);
xor U7607 (N_7607,N_3515,N_2810);
nand U7608 (N_7608,N_2758,N_484);
or U7609 (N_7609,N_3235,N_1264);
and U7610 (N_7610,N_3064,N_2525);
or U7611 (N_7611,N_3217,N_3725);
and U7612 (N_7612,N_2835,N_992);
nor U7613 (N_7613,N_1185,N_595);
nand U7614 (N_7614,N_542,N_3696);
nand U7615 (N_7615,N_2981,N_3708);
xnor U7616 (N_7616,N_3846,N_3832);
nand U7617 (N_7617,N_2888,N_2498);
nand U7618 (N_7618,N_3233,N_1150);
and U7619 (N_7619,N_1527,N_3483);
nand U7620 (N_7620,N_2585,N_3619);
nand U7621 (N_7621,N_657,N_1553);
and U7622 (N_7622,N_1674,N_755);
or U7623 (N_7623,N_1684,N_3484);
and U7624 (N_7624,N_2631,N_803);
or U7625 (N_7625,N_7,N_1722);
nor U7626 (N_7626,N_3034,N_1119);
xnor U7627 (N_7627,N_585,N_3273);
nand U7628 (N_7628,N_1910,N_3702);
nor U7629 (N_7629,N_3767,N_2623);
nand U7630 (N_7630,N_1509,N_3281);
or U7631 (N_7631,N_3496,N_3002);
and U7632 (N_7632,N_303,N_914);
and U7633 (N_7633,N_2262,N_504);
and U7634 (N_7634,N_205,N_3720);
xnor U7635 (N_7635,N_151,N_1950);
nor U7636 (N_7636,N_1743,N_268);
xor U7637 (N_7637,N_2509,N_3144);
or U7638 (N_7638,N_2254,N_2891);
or U7639 (N_7639,N_572,N_1312);
or U7640 (N_7640,N_433,N_1018);
or U7641 (N_7641,N_1847,N_3740);
and U7642 (N_7642,N_1888,N_3700);
nand U7643 (N_7643,N_828,N_3845);
or U7644 (N_7644,N_3090,N_1767);
xnor U7645 (N_7645,N_518,N_744);
xnor U7646 (N_7646,N_3020,N_303);
or U7647 (N_7647,N_2192,N_3685);
nor U7648 (N_7648,N_3089,N_1280);
and U7649 (N_7649,N_3889,N_3306);
and U7650 (N_7650,N_1789,N_3028);
or U7651 (N_7651,N_242,N_670);
nand U7652 (N_7652,N_1817,N_642);
and U7653 (N_7653,N_2550,N_1449);
or U7654 (N_7654,N_3692,N_1805);
nor U7655 (N_7655,N_2061,N_617);
nor U7656 (N_7656,N_1662,N_2790);
or U7657 (N_7657,N_3780,N_1243);
and U7658 (N_7658,N_2283,N_3617);
or U7659 (N_7659,N_1398,N_334);
xnor U7660 (N_7660,N_3251,N_2022);
and U7661 (N_7661,N_2030,N_413);
nor U7662 (N_7662,N_367,N_1875);
nand U7663 (N_7663,N_1620,N_2618);
and U7664 (N_7664,N_1254,N_1637);
or U7665 (N_7665,N_3103,N_1736);
nor U7666 (N_7666,N_2652,N_1661);
nor U7667 (N_7667,N_2977,N_536);
nor U7668 (N_7668,N_1297,N_978);
and U7669 (N_7669,N_3573,N_1934);
or U7670 (N_7670,N_2186,N_97);
nand U7671 (N_7671,N_3,N_789);
nand U7672 (N_7672,N_1477,N_1347);
nor U7673 (N_7673,N_3428,N_267);
and U7674 (N_7674,N_800,N_1811);
nand U7675 (N_7675,N_1880,N_2094);
xnor U7676 (N_7676,N_839,N_831);
nor U7677 (N_7677,N_1264,N_664);
and U7678 (N_7678,N_1064,N_2698);
and U7679 (N_7679,N_264,N_2195);
nor U7680 (N_7680,N_3225,N_3638);
nor U7681 (N_7681,N_90,N_3052);
nor U7682 (N_7682,N_1769,N_1367);
nand U7683 (N_7683,N_2862,N_1226);
or U7684 (N_7684,N_2910,N_3751);
xnor U7685 (N_7685,N_1217,N_1868);
and U7686 (N_7686,N_1482,N_2247);
or U7687 (N_7687,N_3857,N_3381);
and U7688 (N_7688,N_3115,N_1492);
and U7689 (N_7689,N_3022,N_2334);
nand U7690 (N_7690,N_3666,N_873);
and U7691 (N_7691,N_3253,N_1983);
or U7692 (N_7692,N_219,N_1090);
or U7693 (N_7693,N_1931,N_2981);
xor U7694 (N_7694,N_514,N_229);
xnor U7695 (N_7695,N_2566,N_498);
or U7696 (N_7696,N_17,N_114);
and U7697 (N_7697,N_722,N_1502);
or U7698 (N_7698,N_2299,N_2176);
nor U7699 (N_7699,N_1469,N_330);
and U7700 (N_7700,N_811,N_1004);
and U7701 (N_7701,N_1868,N_854);
xor U7702 (N_7702,N_1112,N_1175);
nand U7703 (N_7703,N_1033,N_1427);
nor U7704 (N_7704,N_3983,N_974);
xnor U7705 (N_7705,N_251,N_3043);
or U7706 (N_7706,N_3573,N_2225);
nand U7707 (N_7707,N_1523,N_3743);
or U7708 (N_7708,N_3002,N_3985);
or U7709 (N_7709,N_1230,N_3312);
xor U7710 (N_7710,N_2157,N_1132);
nor U7711 (N_7711,N_2190,N_3696);
and U7712 (N_7712,N_3576,N_2482);
nor U7713 (N_7713,N_1784,N_2522);
xor U7714 (N_7714,N_2052,N_1813);
and U7715 (N_7715,N_1191,N_3084);
nand U7716 (N_7716,N_3409,N_1090);
and U7717 (N_7717,N_2798,N_1686);
or U7718 (N_7718,N_20,N_3035);
and U7719 (N_7719,N_1227,N_3978);
or U7720 (N_7720,N_1600,N_3193);
or U7721 (N_7721,N_1613,N_3800);
or U7722 (N_7722,N_3580,N_1242);
or U7723 (N_7723,N_1176,N_2473);
nor U7724 (N_7724,N_851,N_791);
xor U7725 (N_7725,N_722,N_1102);
or U7726 (N_7726,N_1978,N_1614);
nand U7727 (N_7727,N_1940,N_172);
xor U7728 (N_7728,N_402,N_1958);
nand U7729 (N_7729,N_2877,N_1572);
xnor U7730 (N_7730,N_270,N_3565);
or U7731 (N_7731,N_194,N_3355);
xnor U7732 (N_7732,N_2668,N_2524);
nor U7733 (N_7733,N_3231,N_69);
or U7734 (N_7734,N_3268,N_3531);
and U7735 (N_7735,N_2299,N_2774);
nor U7736 (N_7736,N_1655,N_2667);
xnor U7737 (N_7737,N_430,N_871);
and U7738 (N_7738,N_3818,N_2099);
nor U7739 (N_7739,N_1735,N_2258);
xnor U7740 (N_7740,N_1777,N_646);
and U7741 (N_7741,N_772,N_832);
nor U7742 (N_7742,N_2987,N_967);
nand U7743 (N_7743,N_1841,N_918);
or U7744 (N_7744,N_3104,N_2426);
xnor U7745 (N_7745,N_1085,N_3429);
xnor U7746 (N_7746,N_3317,N_3280);
nand U7747 (N_7747,N_311,N_1011);
and U7748 (N_7748,N_1122,N_473);
nand U7749 (N_7749,N_1373,N_217);
and U7750 (N_7750,N_2639,N_2756);
or U7751 (N_7751,N_216,N_3518);
xnor U7752 (N_7752,N_3159,N_1601);
nand U7753 (N_7753,N_2736,N_3439);
nand U7754 (N_7754,N_943,N_1456);
nor U7755 (N_7755,N_2279,N_2385);
nand U7756 (N_7756,N_3807,N_511);
xnor U7757 (N_7757,N_1362,N_1652);
xnor U7758 (N_7758,N_1747,N_110);
nand U7759 (N_7759,N_3769,N_2720);
xor U7760 (N_7760,N_2003,N_927);
nand U7761 (N_7761,N_3538,N_3806);
xor U7762 (N_7762,N_2190,N_1901);
or U7763 (N_7763,N_2154,N_246);
or U7764 (N_7764,N_142,N_3699);
nand U7765 (N_7765,N_1677,N_2143);
and U7766 (N_7766,N_3420,N_3823);
nand U7767 (N_7767,N_3319,N_2687);
or U7768 (N_7768,N_3070,N_1904);
nand U7769 (N_7769,N_1821,N_847);
and U7770 (N_7770,N_1273,N_1907);
and U7771 (N_7771,N_3458,N_2125);
nor U7772 (N_7772,N_2268,N_3879);
or U7773 (N_7773,N_84,N_767);
and U7774 (N_7774,N_2106,N_657);
or U7775 (N_7775,N_3158,N_1752);
or U7776 (N_7776,N_1543,N_3924);
nor U7777 (N_7777,N_511,N_3914);
or U7778 (N_7778,N_3601,N_2352);
xor U7779 (N_7779,N_3543,N_3303);
xnor U7780 (N_7780,N_3810,N_488);
nor U7781 (N_7781,N_581,N_2280);
xor U7782 (N_7782,N_3472,N_1426);
nand U7783 (N_7783,N_1879,N_1555);
and U7784 (N_7784,N_2207,N_3690);
nor U7785 (N_7785,N_787,N_1234);
and U7786 (N_7786,N_1816,N_1352);
nor U7787 (N_7787,N_115,N_651);
xnor U7788 (N_7788,N_645,N_398);
nor U7789 (N_7789,N_1066,N_2776);
or U7790 (N_7790,N_2313,N_3257);
and U7791 (N_7791,N_881,N_1676);
nand U7792 (N_7792,N_297,N_1545);
and U7793 (N_7793,N_1026,N_343);
or U7794 (N_7794,N_1730,N_2686);
nor U7795 (N_7795,N_734,N_3229);
xnor U7796 (N_7796,N_411,N_1151);
xor U7797 (N_7797,N_2196,N_3025);
nor U7798 (N_7798,N_1570,N_1952);
nand U7799 (N_7799,N_2752,N_320);
xnor U7800 (N_7800,N_620,N_2917);
xnor U7801 (N_7801,N_1200,N_1234);
nor U7802 (N_7802,N_1164,N_1913);
or U7803 (N_7803,N_1571,N_760);
nor U7804 (N_7804,N_2789,N_2493);
nor U7805 (N_7805,N_464,N_1852);
nand U7806 (N_7806,N_38,N_1300);
and U7807 (N_7807,N_2771,N_2436);
xor U7808 (N_7808,N_3135,N_3456);
nand U7809 (N_7809,N_2649,N_3392);
nor U7810 (N_7810,N_841,N_3606);
xnor U7811 (N_7811,N_1829,N_431);
xor U7812 (N_7812,N_1478,N_3561);
xnor U7813 (N_7813,N_2430,N_3082);
or U7814 (N_7814,N_2017,N_1538);
or U7815 (N_7815,N_3838,N_2816);
nand U7816 (N_7816,N_2523,N_2743);
and U7817 (N_7817,N_116,N_2354);
nand U7818 (N_7818,N_3574,N_2098);
and U7819 (N_7819,N_1103,N_3266);
or U7820 (N_7820,N_1087,N_2823);
xnor U7821 (N_7821,N_3873,N_3942);
and U7822 (N_7822,N_2809,N_3526);
nor U7823 (N_7823,N_2643,N_3989);
nand U7824 (N_7824,N_2216,N_3036);
nor U7825 (N_7825,N_1849,N_3550);
nor U7826 (N_7826,N_1312,N_194);
or U7827 (N_7827,N_1678,N_2124);
nand U7828 (N_7828,N_3221,N_1710);
nor U7829 (N_7829,N_2008,N_1008);
nand U7830 (N_7830,N_2799,N_2844);
nor U7831 (N_7831,N_3131,N_565);
and U7832 (N_7832,N_2746,N_1067);
nor U7833 (N_7833,N_3508,N_2879);
nand U7834 (N_7834,N_3156,N_1858);
or U7835 (N_7835,N_1219,N_1311);
or U7836 (N_7836,N_3398,N_3161);
nor U7837 (N_7837,N_337,N_1917);
nand U7838 (N_7838,N_2749,N_3763);
xor U7839 (N_7839,N_2809,N_2544);
xor U7840 (N_7840,N_1180,N_3465);
or U7841 (N_7841,N_2649,N_2771);
nand U7842 (N_7842,N_2362,N_264);
and U7843 (N_7843,N_1806,N_843);
or U7844 (N_7844,N_3588,N_3628);
nor U7845 (N_7845,N_1898,N_3429);
and U7846 (N_7846,N_2726,N_1041);
nor U7847 (N_7847,N_3334,N_938);
nand U7848 (N_7848,N_2353,N_865);
nor U7849 (N_7849,N_1638,N_717);
nor U7850 (N_7850,N_3140,N_3725);
and U7851 (N_7851,N_1235,N_3933);
nor U7852 (N_7852,N_2750,N_3468);
or U7853 (N_7853,N_1017,N_2872);
nor U7854 (N_7854,N_1250,N_766);
nand U7855 (N_7855,N_1289,N_3245);
nand U7856 (N_7856,N_3565,N_2145);
or U7857 (N_7857,N_361,N_3166);
nand U7858 (N_7858,N_2491,N_2616);
nor U7859 (N_7859,N_2897,N_3348);
and U7860 (N_7860,N_2760,N_1955);
and U7861 (N_7861,N_3679,N_1452);
and U7862 (N_7862,N_1414,N_228);
nor U7863 (N_7863,N_1706,N_414);
nor U7864 (N_7864,N_1363,N_133);
nand U7865 (N_7865,N_1989,N_2294);
nand U7866 (N_7866,N_2527,N_3751);
nand U7867 (N_7867,N_1981,N_166);
or U7868 (N_7868,N_638,N_3616);
xor U7869 (N_7869,N_787,N_144);
nor U7870 (N_7870,N_1106,N_1208);
and U7871 (N_7871,N_1898,N_1796);
and U7872 (N_7872,N_701,N_3419);
nand U7873 (N_7873,N_2226,N_3352);
and U7874 (N_7874,N_2379,N_2953);
nand U7875 (N_7875,N_3954,N_2617);
xnor U7876 (N_7876,N_516,N_201);
xor U7877 (N_7877,N_1468,N_3091);
nand U7878 (N_7878,N_443,N_2791);
nor U7879 (N_7879,N_3082,N_1025);
and U7880 (N_7880,N_2029,N_1801);
and U7881 (N_7881,N_110,N_1169);
xor U7882 (N_7882,N_3387,N_2701);
xnor U7883 (N_7883,N_1568,N_124);
xor U7884 (N_7884,N_1734,N_725);
and U7885 (N_7885,N_2749,N_2006);
nor U7886 (N_7886,N_50,N_1086);
or U7887 (N_7887,N_2175,N_3056);
nand U7888 (N_7888,N_846,N_2460);
xnor U7889 (N_7889,N_570,N_738);
xor U7890 (N_7890,N_3148,N_2424);
xnor U7891 (N_7891,N_2139,N_2482);
nor U7892 (N_7892,N_2430,N_3120);
nand U7893 (N_7893,N_1987,N_2533);
xor U7894 (N_7894,N_1361,N_1863);
and U7895 (N_7895,N_1727,N_339);
xnor U7896 (N_7896,N_3749,N_1166);
nand U7897 (N_7897,N_62,N_2746);
or U7898 (N_7898,N_16,N_1610);
and U7899 (N_7899,N_3867,N_1672);
and U7900 (N_7900,N_1616,N_336);
nand U7901 (N_7901,N_3655,N_2332);
nand U7902 (N_7902,N_1732,N_605);
or U7903 (N_7903,N_285,N_2808);
nor U7904 (N_7904,N_2266,N_816);
or U7905 (N_7905,N_990,N_2233);
and U7906 (N_7906,N_2204,N_718);
nor U7907 (N_7907,N_1330,N_736);
xnor U7908 (N_7908,N_3691,N_874);
nor U7909 (N_7909,N_2432,N_2606);
nor U7910 (N_7910,N_2812,N_3151);
or U7911 (N_7911,N_3250,N_696);
xor U7912 (N_7912,N_67,N_3467);
or U7913 (N_7913,N_1531,N_1721);
nand U7914 (N_7914,N_3428,N_551);
nor U7915 (N_7915,N_2102,N_623);
and U7916 (N_7916,N_1502,N_2039);
nand U7917 (N_7917,N_426,N_3372);
xnor U7918 (N_7918,N_2787,N_409);
nand U7919 (N_7919,N_727,N_51);
xor U7920 (N_7920,N_346,N_3885);
nor U7921 (N_7921,N_1139,N_3237);
or U7922 (N_7922,N_1901,N_2876);
or U7923 (N_7923,N_3611,N_1252);
nand U7924 (N_7924,N_3369,N_3462);
or U7925 (N_7925,N_841,N_364);
nand U7926 (N_7926,N_3839,N_241);
nand U7927 (N_7927,N_3869,N_3097);
and U7928 (N_7928,N_3561,N_2618);
nand U7929 (N_7929,N_1174,N_2440);
or U7930 (N_7930,N_3717,N_2093);
nor U7931 (N_7931,N_66,N_3426);
or U7932 (N_7932,N_3981,N_590);
xnor U7933 (N_7933,N_45,N_2136);
nor U7934 (N_7934,N_1138,N_3351);
and U7935 (N_7935,N_2156,N_3426);
xnor U7936 (N_7936,N_1669,N_283);
or U7937 (N_7937,N_2105,N_3834);
nand U7938 (N_7938,N_741,N_1880);
nor U7939 (N_7939,N_2185,N_2815);
xnor U7940 (N_7940,N_1049,N_1525);
or U7941 (N_7941,N_2213,N_773);
nor U7942 (N_7942,N_1569,N_946);
nand U7943 (N_7943,N_3044,N_92);
xor U7944 (N_7944,N_1467,N_3797);
nor U7945 (N_7945,N_3670,N_271);
or U7946 (N_7946,N_2367,N_605);
nor U7947 (N_7947,N_3602,N_1580);
nor U7948 (N_7948,N_2471,N_3410);
nor U7949 (N_7949,N_3536,N_263);
and U7950 (N_7950,N_2636,N_3350);
nand U7951 (N_7951,N_3594,N_1933);
nand U7952 (N_7952,N_2791,N_1284);
nor U7953 (N_7953,N_1393,N_329);
nor U7954 (N_7954,N_153,N_2040);
or U7955 (N_7955,N_3280,N_720);
nand U7956 (N_7956,N_1085,N_2184);
and U7957 (N_7957,N_2855,N_3876);
nand U7958 (N_7958,N_2417,N_2873);
and U7959 (N_7959,N_263,N_2281);
nor U7960 (N_7960,N_256,N_459);
nor U7961 (N_7961,N_601,N_1347);
xor U7962 (N_7962,N_496,N_2902);
and U7963 (N_7963,N_3585,N_998);
nor U7964 (N_7964,N_1495,N_685);
nor U7965 (N_7965,N_132,N_284);
xnor U7966 (N_7966,N_1009,N_1359);
xnor U7967 (N_7967,N_1739,N_3104);
nor U7968 (N_7968,N_2349,N_2159);
xor U7969 (N_7969,N_264,N_1346);
xor U7970 (N_7970,N_3163,N_1628);
xor U7971 (N_7971,N_3637,N_432);
nand U7972 (N_7972,N_1582,N_2162);
xor U7973 (N_7973,N_1492,N_3009);
nand U7974 (N_7974,N_1525,N_2884);
and U7975 (N_7975,N_2308,N_1338);
and U7976 (N_7976,N_1320,N_54);
xor U7977 (N_7977,N_3210,N_3134);
and U7978 (N_7978,N_3113,N_2015);
and U7979 (N_7979,N_2553,N_2384);
and U7980 (N_7980,N_645,N_740);
nand U7981 (N_7981,N_2750,N_316);
nand U7982 (N_7982,N_3020,N_3787);
and U7983 (N_7983,N_1245,N_382);
xnor U7984 (N_7984,N_2131,N_287);
nor U7985 (N_7985,N_1337,N_1464);
nand U7986 (N_7986,N_3684,N_276);
or U7987 (N_7987,N_1216,N_583);
xor U7988 (N_7988,N_1611,N_1478);
and U7989 (N_7989,N_3521,N_334);
nand U7990 (N_7990,N_3517,N_504);
nor U7991 (N_7991,N_1746,N_2923);
xnor U7992 (N_7992,N_2333,N_1230);
nor U7993 (N_7993,N_3482,N_39);
xor U7994 (N_7994,N_2063,N_1865);
or U7995 (N_7995,N_1935,N_2386);
and U7996 (N_7996,N_3678,N_738);
xor U7997 (N_7997,N_1207,N_59);
xnor U7998 (N_7998,N_731,N_2551);
or U7999 (N_7999,N_1784,N_1326);
nor U8000 (N_8000,N_4962,N_4050);
xnor U8001 (N_8001,N_5154,N_5746);
nand U8002 (N_8002,N_4145,N_4289);
nand U8003 (N_8003,N_6839,N_6979);
and U8004 (N_8004,N_6812,N_4335);
nor U8005 (N_8005,N_7287,N_7441);
nor U8006 (N_8006,N_7588,N_6648);
nand U8007 (N_8007,N_7820,N_6793);
or U8008 (N_8008,N_7270,N_4445);
nand U8009 (N_8009,N_6003,N_4800);
nand U8010 (N_8010,N_6036,N_6700);
nor U8011 (N_8011,N_4498,N_4879);
or U8012 (N_8012,N_4294,N_6930);
xor U8013 (N_8013,N_4201,N_5434);
nor U8014 (N_8014,N_5617,N_4029);
or U8015 (N_8015,N_4493,N_6267);
xor U8016 (N_8016,N_6370,N_6223);
nand U8017 (N_8017,N_7426,N_6496);
xnor U8018 (N_8018,N_6637,N_5881);
and U8019 (N_8019,N_5357,N_6257);
xnor U8020 (N_8020,N_4228,N_6950);
xor U8021 (N_8021,N_5808,N_7973);
nor U8022 (N_8022,N_4684,N_5900);
and U8023 (N_8023,N_5728,N_4739);
nor U8024 (N_8024,N_6269,N_7126);
nand U8025 (N_8025,N_6270,N_5195);
xnor U8026 (N_8026,N_5918,N_5114);
nor U8027 (N_8027,N_6408,N_7558);
xnor U8028 (N_8028,N_4302,N_6818);
xor U8029 (N_8029,N_6701,N_7541);
nand U8030 (N_8030,N_7004,N_6449);
xnor U8031 (N_8031,N_4326,N_4956);
or U8032 (N_8032,N_7615,N_4621);
and U8033 (N_8033,N_6880,N_4542);
or U8034 (N_8034,N_6507,N_5879);
nor U8035 (N_8035,N_6155,N_6992);
xnor U8036 (N_8036,N_4417,N_6946);
and U8037 (N_8037,N_7302,N_4339);
and U8038 (N_8038,N_7942,N_7041);
or U8039 (N_8039,N_7540,N_4790);
and U8040 (N_8040,N_6090,N_6233);
xnor U8041 (N_8041,N_5903,N_4546);
or U8042 (N_8042,N_6712,N_7634);
or U8043 (N_8043,N_7711,N_7339);
xor U8044 (N_8044,N_7662,N_4617);
and U8045 (N_8045,N_4644,N_4926);
nand U8046 (N_8046,N_5796,N_5749);
or U8047 (N_8047,N_5963,N_5669);
xnor U8048 (N_8048,N_5361,N_5852);
or U8049 (N_8049,N_5200,N_5572);
or U8050 (N_8050,N_7611,N_5291);
or U8051 (N_8051,N_7969,N_5094);
nor U8052 (N_8052,N_4931,N_5787);
and U8053 (N_8053,N_7629,N_4081);
xor U8054 (N_8054,N_7485,N_5237);
nand U8055 (N_8055,N_7188,N_7111);
and U8056 (N_8056,N_4647,N_4924);
and U8057 (N_8057,N_6931,N_7781);
nand U8058 (N_8058,N_7534,N_6580);
and U8059 (N_8059,N_6834,N_5546);
xor U8060 (N_8060,N_7354,N_7581);
nand U8061 (N_8061,N_6253,N_7345);
nor U8062 (N_8062,N_5709,N_4844);
and U8063 (N_8063,N_7084,N_6088);
or U8064 (N_8064,N_7018,N_5487);
xor U8065 (N_8065,N_4950,N_5172);
xor U8066 (N_8066,N_4311,N_6190);
and U8067 (N_8067,N_4325,N_4393);
xor U8068 (N_8068,N_5255,N_7067);
nor U8069 (N_8069,N_7187,N_5671);
nand U8070 (N_8070,N_4783,N_5547);
and U8071 (N_8071,N_7587,N_7161);
nand U8072 (N_8072,N_7065,N_7199);
and U8073 (N_8073,N_5998,N_4487);
xnor U8074 (N_8074,N_4401,N_5066);
or U8075 (N_8075,N_4168,N_7395);
or U8076 (N_8076,N_4723,N_7136);
or U8077 (N_8077,N_5090,N_4855);
xnor U8078 (N_8078,N_5424,N_7455);
nor U8079 (N_8079,N_7192,N_6897);
nand U8080 (N_8080,N_4492,N_5327);
or U8081 (N_8081,N_4020,N_4589);
nand U8082 (N_8082,N_4305,N_7543);
nand U8083 (N_8083,N_4390,N_5651);
xor U8084 (N_8084,N_5920,N_4922);
and U8085 (N_8085,N_6396,N_6431);
and U8086 (N_8086,N_4270,N_5486);
or U8087 (N_8087,N_6693,N_6969);
and U8088 (N_8088,N_4259,N_4491);
or U8089 (N_8089,N_4109,N_7022);
and U8090 (N_8090,N_5839,N_6334);
nand U8091 (N_8091,N_4164,N_4613);
nand U8092 (N_8092,N_7821,N_6160);
and U8093 (N_8093,N_5049,N_6591);
and U8094 (N_8094,N_4345,N_6705);
nand U8095 (N_8095,N_7656,N_6288);
and U8096 (N_8096,N_6464,N_6632);
nand U8097 (N_8097,N_4406,N_6216);
nand U8098 (N_8098,N_5444,N_5987);
or U8099 (N_8099,N_5199,N_4687);
nand U8100 (N_8100,N_7382,N_7379);
xnor U8101 (N_8101,N_4628,N_4843);
xor U8102 (N_8102,N_4659,N_5176);
nand U8103 (N_8103,N_5054,N_4072);
nor U8104 (N_8104,N_7025,N_7113);
nor U8105 (N_8105,N_7058,N_4720);
or U8106 (N_8106,N_5641,N_4984);
nand U8107 (N_8107,N_4980,N_4362);
nand U8108 (N_8108,N_7974,N_7515);
xnor U8109 (N_8109,N_7612,N_4527);
xnor U8110 (N_8110,N_7862,N_5134);
nor U8111 (N_8111,N_4928,N_7882);
nor U8112 (N_8112,N_4781,N_7191);
xnor U8113 (N_8113,N_4229,N_5609);
or U8114 (N_8114,N_7059,N_6696);
and U8115 (N_8115,N_5028,N_5699);
and U8116 (N_8116,N_7181,N_7823);
nor U8117 (N_8117,N_6644,N_6602);
and U8118 (N_8118,N_6013,N_5904);
nand U8119 (N_8119,N_7357,N_6366);
and U8120 (N_8120,N_6792,N_5296);
or U8121 (N_8121,N_6400,N_6323);
nor U8122 (N_8122,N_4566,N_6862);
and U8123 (N_8123,N_5785,N_4529);
xor U8124 (N_8124,N_7367,N_4773);
xnor U8125 (N_8125,N_6666,N_7854);
and U8126 (N_8126,N_6775,N_6219);
and U8127 (N_8127,N_7529,N_7036);
nand U8128 (N_8128,N_4933,N_4836);
or U8129 (N_8129,N_6441,N_4338);
xor U8130 (N_8130,N_6035,N_7519);
nand U8131 (N_8131,N_6709,N_7933);
xor U8132 (N_8132,N_5734,N_4422);
nor U8133 (N_8133,N_7403,N_7457);
nor U8134 (N_8134,N_6577,N_6776);
nand U8135 (N_8135,N_6654,N_4707);
xnor U8136 (N_8136,N_4948,N_7490);
and U8137 (N_8137,N_6029,N_5123);
nor U8138 (N_8138,N_6587,N_4601);
or U8139 (N_8139,N_4175,N_4102);
xnor U8140 (N_8140,N_6405,N_4795);
xnor U8141 (N_8141,N_5425,N_4640);
and U8142 (N_8142,N_6402,N_5443);
xnor U8143 (N_8143,N_6807,N_5849);
and U8144 (N_8144,N_7647,N_6867);
and U8145 (N_8145,N_6061,N_7369);
xnor U8146 (N_8146,N_4196,N_6312);
nand U8147 (N_8147,N_5618,N_7848);
nor U8148 (N_8148,N_5056,N_4643);
nand U8149 (N_8149,N_4301,N_6111);
nand U8150 (N_8150,N_6806,N_6749);
nor U8151 (N_8151,N_6528,N_5589);
xor U8152 (N_8152,N_5704,N_7996);
and U8153 (N_8153,N_6306,N_5191);
and U8154 (N_8154,N_4955,N_5845);
or U8155 (N_8155,N_6418,N_4633);
nand U8156 (N_8156,N_7262,N_4389);
or U8157 (N_8157,N_4346,N_7238);
xnor U8158 (N_8158,N_4280,N_4112);
xor U8159 (N_8159,N_7796,N_7806);
nor U8160 (N_8160,N_7771,N_7591);
xor U8161 (N_8161,N_6538,N_5445);
nor U8162 (N_8162,N_5750,N_5403);
or U8163 (N_8163,N_6081,N_5768);
nand U8164 (N_8164,N_6935,N_7704);
nor U8165 (N_8165,N_4988,N_7673);
and U8166 (N_8166,N_4363,N_4384);
nand U8167 (N_8167,N_4600,N_6857);
nor U8168 (N_8168,N_7177,N_4411);
nor U8169 (N_8169,N_5912,N_7316);
nor U8170 (N_8170,N_4025,N_5454);
nor U8171 (N_8171,N_7589,N_6801);
xor U8172 (N_8172,N_5418,N_4322);
nand U8173 (N_8173,N_6653,N_6256);
and U8174 (N_8174,N_6611,N_5645);
xor U8175 (N_8175,N_4920,N_4897);
and U8176 (N_8176,N_7003,N_4155);
nor U8177 (N_8177,N_5874,N_6546);
or U8178 (N_8178,N_7994,N_6064);
xor U8179 (N_8179,N_6033,N_7331);
or U8180 (N_8180,N_5924,N_6665);
or U8181 (N_8181,N_7907,N_7722);
and U8182 (N_8182,N_7350,N_7202);
or U8183 (N_8183,N_7987,N_7211);
xor U8184 (N_8184,N_7028,N_6584);
nand U8185 (N_8185,N_5107,N_4638);
nand U8186 (N_8186,N_7697,N_4908);
and U8187 (N_8187,N_4121,N_6631);
or U8188 (N_8188,N_6572,N_4130);
nand U8189 (N_8189,N_5745,N_6137);
nor U8190 (N_8190,N_5364,N_5220);
nor U8191 (N_8191,N_4887,N_5722);
or U8192 (N_8192,N_4975,N_7105);
nand U8193 (N_8193,N_4446,N_7842);
nand U8194 (N_8194,N_7135,N_7073);
nor U8195 (N_8195,N_4544,N_4923);
nand U8196 (N_8196,N_6852,N_5214);
nor U8197 (N_8197,N_7416,N_6926);
nand U8198 (N_8198,N_6905,N_6170);
and U8199 (N_8199,N_6565,N_4991);
nand U8200 (N_8200,N_7653,N_5062);
or U8201 (N_8201,N_7183,N_4021);
and U8202 (N_8202,N_7583,N_4063);
or U8203 (N_8203,N_4724,N_4483);
nor U8204 (N_8204,N_5398,N_6173);
xnor U8205 (N_8205,N_6854,N_5106);
nand U8206 (N_8206,N_4059,N_6413);
xnor U8207 (N_8207,N_5401,N_4892);
and U8208 (N_8208,N_4431,N_5690);
or U8209 (N_8209,N_6467,N_6645);
and U8210 (N_8210,N_4796,N_4833);
or U8211 (N_8211,N_5600,N_5544);
nor U8212 (N_8212,N_5450,N_7929);
and U8213 (N_8213,N_4710,N_5126);
nor U8214 (N_8214,N_6704,N_4022);
nand U8215 (N_8215,N_5503,N_4375);
nor U8216 (N_8216,N_7840,N_4986);
and U8217 (N_8217,N_7010,N_4750);
nor U8218 (N_8218,N_6130,N_7738);
nand U8219 (N_8219,N_7305,N_5073);
xor U8220 (N_8220,N_4144,N_5095);
or U8221 (N_8221,N_5708,N_5657);
or U8222 (N_8222,N_7048,N_6622);
nand U8223 (N_8223,N_5339,N_4917);
nor U8224 (N_8224,N_5777,N_4952);
nor U8225 (N_8225,N_4578,N_7503);
nand U8226 (N_8226,N_7780,N_7535);
nand U8227 (N_8227,N_4142,N_6833);
and U8228 (N_8228,N_6985,N_5701);
and U8229 (N_8229,N_6322,N_7635);
nand U8230 (N_8230,N_4910,N_7982);
nor U8231 (N_8231,N_6077,N_5356);
nand U8232 (N_8232,N_7865,N_7215);
nand U8233 (N_8233,N_5775,N_7916);
xnor U8234 (N_8234,N_7463,N_4263);
or U8235 (N_8235,N_4191,N_4009);
or U8236 (N_8236,N_4309,N_7364);
and U8237 (N_8237,N_5165,N_7739);
or U8238 (N_8238,N_6049,N_4891);
nor U8239 (N_8239,N_4475,N_7857);
xnor U8240 (N_8240,N_4011,N_6607);
nor U8241 (N_8241,N_5001,N_6915);
or U8242 (N_8242,N_6641,N_6615);
nor U8243 (N_8243,N_5579,N_6026);
xor U8244 (N_8244,N_7246,N_4616);
xor U8245 (N_8245,N_6119,N_4571);
xor U8246 (N_8246,N_5504,N_6768);
and U8247 (N_8247,N_4014,N_4451);
and U8248 (N_8248,N_5637,N_5584);
xnor U8249 (N_8249,N_6180,N_6357);
nor U8250 (N_8250,N_6660,N_4173);
xor U8251 (N_8251,N_6001,N_4805);
nand U8252 (N_8252,N_4568,N_7616);
xnor U8253 (N_8253,N_5737,N_6011);
and U8254 (N_8254,N_5212,N_7110);
and U8255 (N_8255,N_7908,N_7822);
and U8256 (N_8256,N_5921,N_7828);
nand U8257 (N_8257,N_4005,N_4013);
nand U8258 (N_8258,N_7712,N_5917);
nor U8259 (N_8259,N_7934,N_7404);
nand U8260 (N_8260,N_5674,N_4661);
and U8261 (N_8261,N_7198,N_6224);
nand U8262 (N_8262,N_6475,N_4224);
and U8263 (N_8263,N_7706,N_4114);
xor U8264 (N_8264,N_7243,N_7687);
xor U8265 (N_8265,N_7143,N_6238);
or U8266 (N_8266,N_4627,N_5529);
xnor U8267 (N_8267,N_6059,N_6633);
and U8268 (N_8268,N_7768,N_6674);
nor U8269 (N_8269,N_6347,N_4106);
or U8270 (N_8270,N_7193,N_7983);
or U8271 (N_8271,N_6045,N_7329);
nor U8272 (N_8272,N_6629,N_7154);
nor U8273 (N_8273,N_4500,N_7894);
xnor U8274 (N_8274,N_5875,N_5192);
nand U8275 (N_8275,N_6780,N_5520);
xnor U8276 (N_8276,N_5160,N_6490);
xor U8277 (N_8277,N_6291,N_7317);
or U8278 (N_8278,N_7391,N_5112);
nand U8279 (N_8279,N_7650,N_4650);
or U8280 (N_8280,N_6582,N_5412);
nor U8281 (N_8281,N_5556,N_6018);
or U8282 (N_8282,N_6516,N_6827);
xor U8283 (N_8283,N_5307,N_7850);
and U8284 (N_8284,N_5536,N_5452);
nand U8285 (N_8285,N_6535,N_7201);
and U8286 (N_8286,N_4605,N_6682);
nor U8287 (N_8287,N_4579,N_7225);
nand U8288 (N_8288,N_4337,N_5366);
nand U8289 (N_8289,N_6429,N_4245);
nor U8290 (N_8290,N_5116,N_4727);
nor U8291 (N_8291,N_4695,N_6175);
xnor U8292 (N_8292,N_6530,N_4176);
nor U8293 (N_8293,N_5866,N_6848);
or U8294 (N_8294,N_5990,N_5740);
or U8295 (N_8295,N_6786,N_6095);
or U8296 (N_8296,N_4026,N_6140);
nor U8297 (N_8297,N_7748,N_6922);
nand U8298 (N_8298,N_7985,N_5449);
and U8299 (N_8299,N_5014,N_6363);
nand U8300 (N_8300,N_4458,N_4745);
nand U8301 (N_8301,N_4299,N_5896);
nor U8302 (N_8302,N_6715,N_7568);
or U8303 (N_8303,N_4671,N_7346);
and U8304 (N_8304,N_4747,N_6755);
or U8305 (N_8305,N_6748,N_5610);
or U8306 (N_8306,N_7251,N_4157);
and U8307 (N_8307,N_6203,N_4698);
nand U8308 (N_8308,N_6714,N_5314);
nand U8309 (N_8309,N_6122,N_5431);
nand U8310 (N_8310,N_7565,N_7280);
nand U8311 (N_8311,N_6390,N_6681);
and U8312 (N_8312,N_7469,N_5906);
and U8313 (N_8313,N_6252,N_7260);
nor U8314 (N_8314,N_7909,N_4027);
or U8315 (N_8315,N_5125,N_4992);
nor U8316 (N_8316,N_7125,N_6575);
or U8317 (N_8317,N_5260,N_6943);
nand U8318 (N_8318,N_5332,N_5862);
or U8319 (N_8319,N_5269,N_7434);
nor U8320 (N_8320,N_5002,N_6157);
or U8321 (N_8321,N_6196,N_6784);
xor U8322 (N_8322,N_6285,N_5502);
nand U8323 (N_8323,N_6016,N_4754);
xor U8324 (N_8324,N_4126,N_5784);
and U8325 (N_8325,N_6638,N_4878);
nand U8326 (N_8326,N_6427,N_6966);
and U8327 (N_8327,N_7265,N_7120);
nand U8328 (N_8328,N_6903,N_5238);
xnor U8329 (N_8329,N_6826,N_5612);
or U8330 (N_8330,N_7789,N_5773);
nor U8331 (N_8331,N_4782,N_6782);
nor U8332 (N_8332,N_6249,N_5940);
and U8333 (N_8333,N_7217,N_4612);
or U8334 (N_8334,N_4039,N_4881);
nor U8335 (N_8335,N_7524,N_5267);
nor U8336 (N_8336,N_5029,N_5938);
and U8337 (N_8337,N_4610,N_7066);
nand U8338 (N_8338,N_5231,N_4430);
nor U8339 (N_8339,N_4798,N_5872);
nor U8340 (N_8340,N_7186,N_7679);
and U8341 (N_8341,N_6191,N_5826);
nor U8342 (N_8342,N_4420,N_6022);
xnor U8343 (N_8343,N_6286,N_5086);
and U8344 (N_8344,N_6015,N_6142);
nor U8345 (N_8345,N_7286,N_6916);
nor U8346 (N_8346,N_7702,N_4258);
nand U8347 (N_8347,N_6614,N_6840);
or U8348 (N_8348,N_7684,N_7536);
and U8349 (N_8349,N_6103,N_4381);
or U8350 (N_8350,N_5204,N_4847);
or U8351 (N_8351,N_7365,N_5654);
nand U8352 (N_8352,N_6900,N_5156);
xnor U8353 (N_8353,N_7306,N_7918);
nand U8354 (N_8354,N_6127,N_5076);
and U8355 (N_8355,N_4110,N_7952);
xnor U8356 (N_8356,N_7049,N_7880);
or U8357 (N_8357,N_4001,N_6139);
or U8358 (N_8358,N_6940,N_4653);
or U8359 (N_8359,N_6978,N_4062);
or U8360 (N_8360,N_7756,N_4036);
and U8361 (N_8361,N_7671,N_7374);
nor U8362 (N_8362,N_4221,N_5170);
and U8363 (N_8363,N_6236,N_4906);
xor U8364 (N_8364,N_5718,N_5816);
xor U8365 (N_8365,N_5281,N_7509);
nor U8366 (N_8366,N_5039,N_5621);
xnor U8367 (N_8367,N_5194,N_5102);
and U8368 (N_8368,N_6330,N_6934);
nor U8369 (N_8369,N_6673,N_5495);
nor U8370 (N_8370,N_7319,N_5128);
nor U8371 (N_8371,N_7026,N_4737);
nor U8372 (N_8372,N_4332,N_7531);
or U8373 (N_8373,N_4995,N_7229);
xnor U8374 (N_8374,N_5496,N_5869);
xnor U8375 (N_8375,N_7851,N_4635);
and U8376 (N_8376,N_7641,N_5697);
nand U8377 (N_8377,N_4961,N_7632);
xor U8378 (N_8378,N_6412,N_5349);
nand U8379 (N_8379,N_6723,N_7131);
and U8380 (N_8380,N_5000,N_4954);
nand U8381 (N_8381,N_4075,N_5455);
nand U8382 (N_8382,N_6961,N_7601);
nor U8383 (N_8383,N_7745,N_6525);
xor U8384 (N_8384,N_5736,N_5760);
nor U8385 (N_8385,N_5227,N_7868);
nor U8386 (N_8386,N_5757,N_5447);
xnor U8387 (N_8387,N_7134,N_6708);
nor U8388 (N_8388,N_7945,N_4748);
nand U8389 (N_8389,N_6845,N_4731);
xnor U8390 (N_8390,N_7995,N_6711);
nor U8391 (N_8391,N_5018,N_4324);
or U8392 (N_8392,N_6918,N_7686);
or U8393 (N_8393,N_7377,N_5535);
nand U8394 (N_8394,N_5135,N_6986);
nand U8395 (N_8395,N_5138,N_4706);
nor U8396 (N_8396,N_7567,N_5139);
or U8397 (N_8397,N_4143,N_6382);
or U8398 (N_8398,N_4348,N_4996);
and U8399 (N_8399,N_4333,N_5350);
xnor U8400 (N_8400,N_6433,N_7257);
nand U8401 (N_8401,N_4207,N_4403);
nor U8402 (N_8402,N_4031,N_5553);
and U8403 (N_8403,N_6866,N_7948);
and U8404 (N_8404,N_7902,N_5995);
xnor U8405 (N_8405,N_6817,N_6042);
or U8406 (N_8406,N_5967,N_4018);
and U8407 (N_8407,N_7166,N_6624);
nor U8408 (N_8408,N_5949,N_5567);
or U8409 (N_8409,N_5333,N_5942);
xor U8410 (N_8410,N_6020,N_6320);
and U8411 (N_8411,N_4738,N_5221);
nor U8412 (N_8412,N_7905,N_7578);
xnor U8413 (N_8413,N_6529,N_6948);
nand U8414 (N_8414,N_5252,N_6885);
xor U8415 (N_8415,N_7083,N_4077);
nand U8416 (N_8416,N_5010,N_7207);
and U8417 (N_8417,N_5646,N_7849);
nand U8418 (N_8418,N_6729,N_5604);
xor U8419 (N_8419,N_7413,N_7569);
or U8420 (N_8420,N_6855,N_7414);
nor U8421 (N_8421,N_7023,N_5347);
or U8422 (N_8422,N_7576,N_5328);
or U8423 (N_8423,N_7362,N_6576);
or U8424 (N_8424,N_4392,N_7843);
nor U8425 (N_8425,N_5402,N_5955);
nand U8426 (N_8426,N_6994,N_7799);
nor U8427 (N_8427,N_6295,N_7677);
nor U8428 (N_8428,N_5429,N_5515);
and U8429 (N_8429,N_4515,N_5488);
nand U8430 (N_8430,N_7294,N_6126);
nor U8431 (N_8431,N_6171,N_5545);
and U8432 (N_8432,N_4456,N_7838);
nor U8433 (N_8433,N_6469,N_7087);
xor U8434 (N_8434,N_6851,N_7011);
nand U8435 (N_8435,N_6461,N_6025);
nor U8436 (N_8436,N_7920,N_6343);
and U8437 (N_8437,N_6774,N_6192);
or U8438 (N_8438,N_5457,N_7459);
xnor U8439 (N_8439,N_4312,N_6933);
nand U8440 (N_8440,N_5490,N_6415);
and U8441 (N_8441,N_6054,N_4669);
nor U8442 (N_8442,N_6129,N_6822);
nor U8443 (N_8443,N_5422,N_7385);
nand U8444 (N_8444,N_6805,N_4539);
and U8445 (N_8445,N_5470,N_7770);
nand U8446 (N_8446,N_7932,N_6892);
xnor U8447 (N_8447,N_6006,N_6371);
nand U8448 (N_8448,N_6232,N_5365);
nor U8449 (N_8449,N_5019,N_6761);
and U8450 (N_8450,N_5691,N_4107);
nor U8451 (N_8451,N_5415,N_4885);
nand U8452 (N_8452,N_6965,N_5038);
or U8453 (N_8453,N_7206,N_7016);
nor U8454 (N_8454,N_6437,N_7728);
xnor U8455 (N_8455,N_5428,N_7168);
nand U8456 (N_8456,N_7866,N_5289);
and U8457 (N_8457,N_7222,N_5819);
or U8458 (N_8458,N_7388,N_4524);
nand U8459 (N_8459,N_7348,N_5119);
nor U8460 (N_8460,N_5363,N_4496);
and U8461 (N_8461,N_4436,N_4386);
nand U8462 (N_8462,N_5044,N_4414);
and U8463 (N_8463,N_6778,N_6471);
and U8464 (N_8464,N_6031,N_4983);
and U8465 (N_8465,N_5310,N_5295);
and U8466 (N_8466,N_6562,N_4876);
xnor U8467 (N_8467,N_6802,N_7658);
or U8468 (N_8468,N_6713,N_6387);
or U8469 (N_8469,N_4052,N_6581);
nor U8470 (N_8470,N_5414,N_4098);
xnor U8471 (N_8471,N_4793,N_4208);
and U8472 (N_8472,N_7245,N_5925);
and U8473 (N_8473,N_5177,N_4407);
nor U8474 (N_8474,N_4851,N_7130);
nor U8475 (N_8475,N_7645,N_7574);
xnor U8476 (N_8476,N_7250,N_4134);
xor U8477 (N_8477,N_5877,N_4394);
or U8478 (N_8478,N_5141,N_6456);
xor U8479 (N_8479,N_4410,N_7274);
and U8480 (N_8480,N_7147,N_4169);
nor U8481 (N_8481,N_5005,N_7846);
and U8482 (N_8482,N_6647,N_7887);
nor U8483 (N_8483,N_7743,N_6113);
or U8484 (N_8484,N_5275,N_5206);
nor U8485 (N_8485,N_7924,N_4148);
or U8486 (N_8486,N_5313,N_5132);
nand U8487 (N_8487,N_6166,N_6968);
nor U8488 (N_8488,N_6895,N_5224);
nand U8489 (N_8489,N_5725,N_6958);
and U8490 (N_8490,N_6255,N_5466);
and U8491 (N_8491,N_6702,N_7400);
xnor U8492 (N_8492,N_6554,N_7812);
or U8493 (N_8493,N_6215,N_5929);
or U8494 (N_8494,N_7035,N_5277);
nor U8495 (N_8495,N_5246,N_7228);
nand U8496 (N_8496,N_5263,N_7742);
xnor U8497 (N_8497,N_7078,N_7736);
nor U8498 (N_8498,N_7440,N_4167);
or U8499 (N_8499,N_7213,N_4771);
and U8500 (N_8500,N_5097,N_5059);
or U8501 (N_8501,N_4463,N_7514);
nor U8502 (N_8502,N_4321,N_7696);
or U8503 (N_8503,N_4718,N_4835);
nand U8504 (N_8504,N_5249,N_7203);
nor U8505 (N_8505,N_7387,N_5175);
nand U8506 (N_8506,N_5109,N_6838);
and U8507 (N_8507,N_5435,N_5025);
or U8508 (N_8508,N_6762,N_7546);
or U8509 (N_8509,N_4067,N_4815);
nand U8510 (N_8510,N_4286,N_6517);
or U8511 (N_8511,N_7839,N_6416);
and U8512 (N_8512,N_5331,N_5926);
and U8513 (N_8513,N_7096,N_5984);
or U8514 (N_8514,N_5404,N_6181);
and U8515 (N_8515,N_5345,N_7127);
nand U8516 (N_8516,N_6519,N_7182);
nand U8517 (N_8517,N_5055,N_7454);
nor U8518 (N_8518,N_7644,N_4146);
nand U8519 (N_8519,N_5635,N_6634);
or U8520 (N_8520,N_5492,N_7427);
or U8521 (N_8521,N_6272,N_4040);
or U8522 (N_8522,N_5812,N_6410);
xor U8523 (N_8523,N_6842,N_4901);
or U8524 (N_8524,N_4351,N_4846);
xnor U8525 (N_8525,N_7330,N_5625);
and U8526 (N_8526,N_6495,N_5779);
or U8527 (N_8527,N_4136,N_7944);
and U8528 (N_8528,N_5322,N_5712);
nor U8529 (N_8529,N_7984,N_7584);
nand U8530 (N_8530,N_7235,N_6853);
and U8531 (N_8531,N_6053,N_5223);
or U8532 (N_8532,N_6763,N_6603);
or U8533 (N_8533,N_5299,N_4559);
and U8534 (N_8534,N_4104,N_4383);
nand U8535 (N_8535,N_5799,N_7885);
nor U8536 (N_8536,N_7779,N_4076);
and U8537 (N_8537,N_4866,N_6726);
nand U8538 (N_8538,N_5348,N_5975);
nor U8539 (N_8539,N_5440,N_6104);
nand U8540 (N_8540,N_5052,N_6071);
and U8541 (N_8541,N_6571,N_4794);
nand U8542 (N_8542,N_6789,N_4606);
xnor U8543 (N_8543,N_7077,N_4287);
nor U8544 (N_8544,N_7140,N_5163);
and U8545 (N_8545,N_5655,N_5105);
xnor U8546 (N_8546,N_4034,N_4903);
xor U8547 (N_8547,N_4281,N_7815);
nor U8548 (N_8548,N_5048,N_4696);
nand U8549 (N_8549,N_5675,N_7361);
nand U8550 (N_8550,N_4665,N_5292);
or U8551 (N_8551,N_6212,N_6860);
and U8552 (N_8552,N_6823,N_4517);
nor U8553 (N_8553,N_7776,N_6980);
or U8554 (N_8554,N_5541,N_4651);
and U8555 (N_8555,N_4115,N_4083);
nand U8556 (N_8556,N_4839,N_7499);
xor U8557 (N_8557,N_5776,N_4911);
nand U8558 (N_8558,N_6294,N_6664);
nor U8559 (N_8559,N_7408,N_7070);
or U8560 (N_8560,N_7542,N_4257);
xnor U8561 (N_8561,N_4829,N_6947);
nor U8562 (N_8562,N_7977,N_7383);
nor U8563 (N_8563,N_6428,N_5886);
nor U8564 (N_8564,N_6010,N_7640);
nand U8565 (N_8565,N_6896,N_7972);
and U8566 (N_8566,N_7335,N_5744);
nand U8567 (N_8567,N_4197,N_5828);
nand U8568 (N_8568,N_7695,N_6351);
nor U8569 (N_8569,N_7000,N_6375);
xnor U8570 (N_8570,N_6555,N_7626);
and U8571 (N_8571,N_7804,N_5525);
or U8572 (N_8572,N_5187,N_4268);
and U8573 (N_8573,N_5136,N_7705);
xnor U8574 (N_8574,N_5432,N_4183);
xor U8575 (N_8575,N_4220,N_5070);
nor U8576 (N_8576,N_7941,N_4251);
and U8577 (N_8577,N_6785,N_5247);
nor U8578 (N_8578,N_5489,N_6639);
or U8579 (N_8579,N_6096,N_7392);
xor U8580 (N_8580,N_7772,N_6656);
nor U8581 (N_8581,N_5876,N_4654);
nand U8582 (N_8582,N_4320,N_7356);
xor U8583 (N_8583,N_6767,N_5285);
xor U8584 (N_8584,N_7513,N_5371);
nor U8585 (N_8585,N_5323,N_7919);
nand U8586 (N_8586,N_6891,N_6542);
and U8587 (N_8587,N_7877,N_6108);
nand U8588 (N_8588,N_5325,N_5847);
nor U8589 (N_8589,N_6338,N_7156);
or U8590 (N_8590,N_5950,N_5518);
nor U8591 (N_8591,N_6116,N_7721);
and U8592 (N_8592,N_7167,N_5894);
nand U8593 (N_8593,N_4117,N_7352);
and U8594 (N_8594,N_5210,N_4740);
or U8595 (N_8595,N_7795,N_7744);
and U8596 (N_8596,N_7107,N_4060);
or U8597 (N_8597,N_5608,N_7394);
or U8598 (N_8598,N_4441,N_5959);
nand U8599 (N_8599,N_4946,N_6888);
nand U8600 (N_8600,N_5882,N_5117);
or U8601 (N_8601,N_6829,N_6076);
or U8602 (N_8602,N_7299,N_6987);
nand U8603 (N_8603,N_6446,N_6339);
nor U8604 (N_8604,N_5794,N_4365);
xor U8605 (N_8605,N_5756,N_6289);
xor U8606 (N_8606,N_6589,N_4959);
xnor U8607 (N_8607,N_6277,N_6172);
and U8608 (N_8608,N_4214,N_4803);
or U8609 (N_8609,N_5509,N_5597);
nand U8610 (N_8610,N_5481,N_5763);
or U8611 (N_8611,N_5902,N_5146);
nor U8612 (N_8612,N_5408,N_4217);
nor U8613 (N_8613,N_4283,N_4927);
xnor U8614 (N_8614,N_4085,N_6613);
nand U8615 (N_8615,N_4770,N_4797);
nand U8616 (N_8616,N_6697,N_4577);
nand U8617 (N_8617,N_6744,N_6569);
xnor U8618 (N_8618,N_6678,N_6964);
or U8619 (N_8619,N_7458,N_6319);
or U8620 (N_8620,N_6152,N_6041);
nand U8621 (N_8621,N_7153,N_4824);
nand U8622 (N_8622,N_5382,N_4567);
nor U8623 (N_8623,N_4079,N_5911);
nor U8624 (N_8624,N_6963,N_7518);
nand U8625 (N_8625,N_5113,N_7639);
xnor U8626 (N_8626,N_6133,N_5484);
xnor U8627 (N_8627,N_7442,N_5517);
xor U8628 (N_8628,N_4973,N_7376);
or U8629 (N_8629,N_7980,N_7472);
nand U8630 (N_8630,N_6929,N_7654);
nor U8631 (N_8631,N_7579,N_5992);
or U8632 (N_8632,N_5863,N_7236);
nor U8633 (N_8633,N_6942,N_6163);
and U8634 (N_8634,N_7683,N_5976);
nand U8635 (N_8635,N_5219,N_5483);
or U8636 (N_8636,N_7963,N_6376);
nand U8637 (N_8637,N_5372,N_7617);
nor U8638 (N_8638,N_5870,N_6178);
nand U8639 (N_8639,N_6560,N_6019);
and U8640 (N_8640,N_7212,N_4055);
or U8641 (N_8641,N_6953,N_6734);
or U8642 (N_8642,N_6597,N_5803);
xor U8643 (N_8643,N_6193,N_5164);
or U8644 (N_8644,N_7308,N_5985);
nand U8645 (N_8645,N_6717,N_5672);
nor U8646 (N_8646,N_7314,N_4867);
nand U8647 (N_8647,N_4611,N_7415);
nor U8648 (N_8648,N_5815,N_7888);
or U8649 (N_8649,N_5036,N_7560);
and U8650 (N_8650,N_5652,N_4632);
and U8651 (N_8651,N_4921,N_4254);
xor U8652 (N_8652,N_7253,N_7052);
and U8653 (N_8653,N_6904,N_5417);
nand U8654 (N_8654,N_7807,N_7947);
xnor U8655 (N_8655,N_7190,N_7278);
nor U8656 (N_8656,N_5268,N_6406);
and U8657 (N_8657,N_6278,N_7668);
nand U8658 (N_8658,N_7753,N_6688);
nand U8659 (N_8659,N_6598,N_5179);
nand U8660 (N_8660,N_5391,N_4038);
and U8661 (N_8661,N_7132,N_5539);
and U8662 (N_8662,N_6799,N_4494);
nand U8663 (N_8663,N_4570,N_5387);
nor U8664 (N_8664,N_4425,N_4473);
and U8665 (N_8665,N_7449,N_7360);
nand U8666 (N_8666,N_4331,N_6009);
nand U8667 (N_8667,N_4787,N_6242);
or U8668 (N_8668,N_6932,N_7486);
nor U8669 (N_8669,N_5264,N_7912);
and U8670 (N_8670,N_4080,N_7242);
nand U8671 (N_8671,N_5868,N_6752);
and U8672 (N_8672,N_4049,N_4360);
or U8673 (N_8673,N_5931,N_5851);
nor U8674 (N_8674,N_7600,N_4202);
and U8675 (N_8675,N_7091,N_7298);
nand U8676 (N_8676,N_4206,N_6194);
xnor U8677 (N_8677,N_7498,N_5013);
nand U8678 (N_8678,N_4652,N_4862);
xor U8679 (N_8679,N_4532,N_7923);
nand U8680 (N_8680,N_7883,N_6549);
nor U8681 (N_8681,N_7571,N_4285);
nor U8682 (N_8682,N_5898,N_6566);
nand U8683 (N_8683,N_5592,N_7968);
nand U8684 (N_8684,N_5396,N_6765);
xor U8685 (N_8685,N_4474,N_4615);
xor U8686 (N_8686,N_6329,N_7700);
nor U8687 (N_8687,N_7593,N_4497);
xor U8688 (N_8688,N_4823,N_4634);
or U8689 (N_8689,N_5511,N_5168);
and U8690 (N_8690,N_4247,N_6498);
nor U8691 (N_8691,N_5695,N_6691);
xnor U8692 (N_8692,N_7210,N_7962);
nand U8693 (N_8693,N_4447,N_4998);
or U8694 (N_8694,N_4472,N_7055);
xor U8695 (N_8695,N_5892,N_7715);
and U8696 (N_8696,N_4935,N_5475);
nor U8697 (N_8697,N_7200,N_5578);
and U8698 (N_8698,N_6526,N_4664);
nand U8699 (N_8699,N_4689,N_5311);
nand U8700 (N_8700,N_4541,N_6386);
nor U8701 (N_8701,N_7802,N_6694);
nand U8702 (N_8702,N_4602,N_4678);
or U8703 (N_8703,N_6315,N_6975);
nor U8704 (N_8704,N_7466,N_6491);
nor U8705 (N_8705,N_4806,N_5344);
nand U8706 (N_8706,N_5276,N_6539);
xor U8707 (N_8707,N_7320,N_4941);
nand U8708 (N_8708,N_7101,N_4113);
or U8709 (N_8709,N_6476,N_7368);
nor U8710 (N_8710,N_7218,N_7526);
nor U8711 (N_8711,N_4658,N_5827);
nand U8712 (N_8712,N_7620,N_7676);
nand U8713 (N_8713,N_7324,N_7740);
nor U8714 (N_8714,N_4093,N_5622);
nand U8715 (N_8715,N_6220,N_6439);
nor U8716 (N_8716,N_4788,N_4188);
xnor U8717 (N_8717,N_5061,N_7648);
xor U8718 (N_8718,N_7691,N_7643);
nor U8719 (N_8719,N_6949,N_4010);
xnor U8720 (N_8720,N_5421,N_6630);
or U8721 (N_8721,N_4404,N_5469);
and U8722 (N_8722,N_4387,N_7792);
and U8723 (N_8723,N_6524,N_6070);
nor U8724 (N_8724,N_4869,N_7836);
xnor U8725 (N_8725,N_7505,N_5390);
nor U8726 (N_8726,N_6132,N_6457);
and U8727 (N_8727,N_6385,N_7405);
xor U8728 (N_8728,N_6512,N_5051);
xor U8729 (N_8729,N_4704,N_5732);
and U8730 (N_8730,N_4275,N_6797);
and U8731 (N_8731,N_7480,N_7195);
nor U8732 (N_8732,N_4976,N_6676);
xnor U8733 (N_8733,N_4677,N_5969);
and U8734 (N_8734,N_5947,N_4019);
nor U8735 (N_8735,N_5272,N_4174);
or U8736 (N_8736,N_6850,N_5648);
and U8737 (N_8737,N_4682,N_5037);
and U8738 (N_8738,N_7230,N_6460);
nand U8739 (N_8739,N_7876,N_4930);
or U8740 (N_8740,N_6199,N_4812);
nor U8741 (N_8741,N_4032,N_6738);
nand U8742 (N_8742,N_7765,N_7266);
or U8743 (N_8743,N_7790,N_7321);
nor U8744 (N_8744,N_6595,N_6865);
nor U8745 (N_8745,N_6902,N_4453);
nor U8746 (N_8746,N_5788,N_5989);
xnor U8747 (N_8747,N_5273,N_4203);
and U8748 (N_8748,N_4637,N_7272);
nor U8749 (N_8749,N_6621,N_4507);
xor U8750 (N_8750,N_6235,N_4967);
nand U8751 (N_8751,N_4697,N_5715);
nor U8752 (N_8752,N_4128,N_7599);
nor U8753 (N_8753,N_5270,N_4900);
or U8754 (N_8754,N_7826,N_7863);
and U8755 (N_8755,N_6534,N_4303);
and U8756 (N_8756,N_7598,N_6800);
and U8757 (N_8757,N_7527,N_6048);
nor U8758 (N_8758,N_6228,N_5817);
xnor U8759 (N_8759,N_5607,N_4535);
nand U8760 (N_8760,N_6796,N_5914);
or U8761 (N_8761,N_7910,N_4118);
or U8762 (N_8762,N_7412,N_5823);
or U8763 (N_8763,N_4525,N_6091);
nand U8764 (N_8764,N_7495,N_6411);
or U8765 (N_8765,N_6254,N_7152);
or U8766 (N_8766,N_4334,N_6409);
nand U8767 (N_8767,N_6532,N_7090);
or U8768 (N_8768,N_6506,N_6079);
nand U8769 (N_8769,N_4636,N_6268);
nor U8770 (N_8770,N_5359,N_7886);
xnor U8771 (N_8771,N_5710,N_4170);
nor U8772 (N_8772,N_7614,N_6585);
nor U8773 (N_8773,N_4477,N_7553);
xnor U8774 (N_8774,N_7359,N_7162);
xnor U8775 (N_8775,N_7327,N_5772);
nand U8776 (N_8776,N_6145,N_5441);
nor U8777 (N_8777,N_7473,N_6422);
or U8778 (N_8778,N_4550,N_7050);
nor U8779 (N_8779,N_4396,N_6149);
or U8780 (N_8780,N_4909,N_4646);
nor U8781 (N_8781,N_4502,N_7680);
nand U8782 (N_8782,N_6989,N_7197);
xnor U8783 (N_8783,N_4971,N_6814);
and U8784 (N_8784,N_4158,N_5278);
nor U8785 (N_8785,N_6318,N_4421);
nor U8786 (N_8786,N_4536,N_7284);
and U8787 (N_8787,N_7766,N_5563);
and U8788 (N_8788,N_4951,N_6783);
and U8789 (N_8789,N_4631,N_4757);
nor U8790 (N_8790,N_4035,N_5754);
xnor U8791 (N_8791,N_5171,N_5793);
or U8792 (N_8792,N_6677,N_6039);
nand U8793 (N_8793,N_5373,N_4124);
and U8794 (N_8794,N_6651,N_6276);
nand U8795 (N_8795,N_7597,N_7891);
nand U8796 (N_8796,N_5243,N_4053);
nand U8797 (N_8797,N_4629,N_7148);
xor U8798 (N_8798,N_7295,N_5538);
nor U8799 (N_8799,N_5145,N_5384);
or U8800 (N_8800,N_7303,N_6044);
nor U8801 (N_8801,N_4882,N_7718);
xor U8802 (N_8802,N_4162,N_7609);
and U8803 (N_8803,N_5185,N_5936);
xnor U8804 (N_8804,N_4218,N_5298);
nand U8805 (N_8805,N_5889,N_5067);
nor U8806 (N_8806,N_7724,N_4947);
nand U8807 (N_8807,N_6692,N_4728);
and U8808 (N_8808,N_6809,N_5742);
or U8809 (N_8809,N_6583,N_7661);
nor U8810 (N_8810,N_4756,N_5588);
and U8811 (N_8811,N_6533,N_6007);
nand U8812 (N_8812,N_5201,N_6485);
and U8813 (N_8813,N_6162,N_4070);
and U8814 (N_8814,N_4681,N_7027);
nor U8815 (N_8815,N_7479,N_7904);
and U8816 (N_8816,N_6159,N_4057);
and U8817 (N_8817,N_5807,N_7755);
and U8818 (N_8818,N_7268,N_7304);
and U8819 (N_8819,N_5155,N_4185);
xnor U8820 (N_8820,N_4683,N_7834);
and U8821 (N_8821,N_6047,N_7709);
and U8822 (N_8822,N_5748,N_4732);
or U8823 (N_8823,N_6135,N_4814);
and U8824 (N_8824,N_4105,N_6040);
and U8825 (N_8825,N_5964,N_5979);
xor U8826 (N_8826,N_5820,N_6293);
nand U8827 (N_8827,N_6890,N_5406);
xor U8828 (N_8828,N_5362,N_6690);
nand U8829 (N_8829,N_4703,N_5551);
nor U8830 (N_8830,N_5790,N_5626);
or U8831 (N_8831,N_6474,N_6970);
or U8832 (N_8832,N_5684,N_4744);
xor U8833 (N_8833,N_6308,N_7701);
nand U8834 (N_8834,N_6609,N_5381);
nor U8835 (N_8835,N_7138,N_5887);
nor U8836 (N_8836,N_6017,N_4213);
and U8837 (N_8837,N_5091,N_6395);
and U8838 (N_8838,N_7595,N_5587);
or U8839 (N_8839,N_7476,N_4046);
nor U8840 (N_8840,N_4041,N_5593);
and U8841 (N_8841,N_5636,N_6144);
nor U8842 (N_8842,N_4645,N_6545);
nor U8843 (N_8843,N_5679,N_6661);
or U8844 (N_8844,N_6497,N_6623);
or U8845 (N_8845,N_6552,N_6182);
xor U8846 (N_8846,N_5355,N_7911);
or U8847 (N_8847,N_4811,N_4767);
nand U8848 (N_8848,N_5526,N_7056);
xor U8849 (N_8849,N_5008,N_5880);
and U8850 (N_8850,N_7398,N_6923);
and U8851 (N_8851,N_5640,N_6202);
xor U8852 (N_8852,N_7053,N_6509);
or U8853 (N_8853,N_4368,N_7922);
or U8854 (N_8854,N_7547,N_6341);
nor U8855 (N_8855,N_4769,N_7118);
nand U8856 (N_8856,N_6307,N_4216);
nand U8857 (N_8857,N_7906,N_6425);
and U8858 (N_8858,N_4101,N_4266);
xor U8859 (N_8859,N_6195,N_6881);
or U8860 (N_8860,N_4760,N_6058);
nand U8861 (N_8861,N_7114,N_7500);
xnor U8862 (N_8862,N_4813,N_6924);
nand U8863 (N_8863,N_4593,N_5015);
xnor U8864 (N_8864,N_4435,N_5993);
nand U8865 (N_8865,N_4449,N_4003);
and U8866 (N_8866,N_6240,N_6815);
nor U8867 (N_8867,N_7630,N_7573);
or U8868 (N_8868,N_4061,N_4553);
nor U8869 (N_8869,N_5997,N_6056);
and U8870 (N_8870,N_4448,N_7689);
xor U8871 (N_8871,N_4915,N_7223);
nor U8872 (N_8872,N_7899,N_4310);
or U8873 (N_8873,N_5326,N_7562);
nor U8874 (N_8874,N_4426,N_7275);
xor U8875 (N_8875,N_6668,N_5034);
nand U8876 (N_8876,N_4886,N_7725);
and U8877 (N_8877,N_7508,N_7310);
xor U8878 (N_8878,N_6372,N_5996);
nand U8879 (N_8879,N_7045,N_7402);
nor U8880 (N_8880,N_7334,N_5743);
and U8881 (N_8881,N_5405,N_5181);
nor U8882 (N_8882,N_7037,N_4232);
nand U8883 (N_8883,N_7502,N_6472);
or U8884 (N_8884,N_4511,N_7642);
and U8885 (N_8885,N_6899,N_4587);
nor U8886 (N_8886,N_7497,N_7520);
and U8887 (N_8887,N_7219,N_6292);
xor U8888 (N_8888,N_4304,N_4716);
xor U8889 (N_8889,N_5129,N_5262);
nor U8890 (N_8890,N_4555,N_7988);
xnor U8891 (N_8891,N_6508,N_7410);
xor U8892 (N_8892,N_7549,N_5603);
or U8893 (N_8893,N_7106,N_5841);
xnor U8894 (N_8894,N_7019,N_7528);
nor U8895 (N_8895,N_5184,N_7861);
nand U8896 (N_8896,N_4152,N_7489);
nand U8897 (N_8897,N_7544,N_4166);
xor U8898 (N_8898,N_4506,N_4327);
or U8899 (N_8899,N_6578,N_4741);
or U8900 (N_8900,N_4236,N_7898);
and U8901 (N_8901,N_4753,N_6808);
and U8902 (N_8902,N_5075,N_5683);
nor U8903 (N_8903,N_6771,N_6099);
xor U8904 (N_8904,N_5735,N_5189);
xnor U8905 (N_8905,N_4630,N_4253);
or U8906 (N_8906,N_7008,N_7602);
xor U8907 (N_8907,N_5897,N_4488);
or U8908 (N_8908,N_6301,N_5068);
or U8909 (N_8909,N_7669,N_7184);
and U8910 (N_8910,N_5664,N_4852);
nor U8911 (N_8911,N_7884,N_4150);
nor U8912 (N_8912,N_4242,N_4358);
and U8913 (N_8913,N_4402,N_7063);
and U8914 (N_8914,N_7824,N_5512);
and U8915 (N_8915,N_7116,N_6698);
nand U8916 (N_8916,N_7936,N_7554);
nor U8917 (N_8917,N_4925,N_4932);
and U8918 (N_8918,N_6393,N_4736);
or U8919 (N_8919,N_7961,N_5031);
and U8920 (N_8920,N_7428,N_6165);
nor U8921 (N_8921,N_4234,N_5676);
nand U8922 (N_8922,N_7729,N_5498);
nor U8923 (N_8923,N_7102,N_7068);
or U8924 (N_8924,N_6628,N_7971);
nor U8925 (N_8925,N_7355,N_4291);
and U8926 (N_8926,N_4149,N_5197);
nor U8927 (N_8927,N_5680,N_7717);
or U8928 (N_8928,N_7749,N_7845);
and U8929 (N_8929,N_7089,N_7890);
nor U8930 (N_8930,N_7057,N_7456);
or U8931 (N_8931,N_5423,N_4347);
nand U8932 (N_8932,N_7064,N_4341);
nor U8933 (N_8933,N_4693,N_7782);
and U8934 (N_8934,N_6417,N_6197);
nand U8935 (N_8935,N_4692,N_6421);
nand U8936 (N_8936,N_7949,N_6080);
nand U8937 (N_8937,N_5813,N_4974);
and U8938 (N_8938,N_5133,N_4023);
and U8939 (N_8939,N_5127,N_7692);
or U8940 (N_8940,N_5527,N_7778);
xnor U8941 (N_8941,N_7791,N_4821);
nor U8942 (N_8942,N_5283,N_6444);
and U8943 (N_8943,N_4252,N_6513);
nand U8944 (N_8944,N_5271,N_5753);
or U8945 (N_8945,N_5161,N_4936);
or U8946 (N_8946,N_4153,N_6618);
nand U8947 (N_8947,N_7216,N_7425);
nor U8948 (N_8948,N_6680,N_5236);
nor U8949 (N_8949,N_7585,N_5822);
nor U8950 (N_8950,N_7046,N_4415);
or U8951 (N_8951,N_5098,N_6573);
nand U8952 (N_8952,N_4765,N_5662);
xor U8953 (N_8953,N_6686,N_4830);
xor U8954 (N_8954,N_4452,N_5933);
and U8955 (N_8955,N_7551,N_5688);
nand U8956 (N_8956,N_5353,N_5392);
and U8957 (N_8957,N_5078,N_5686);
xnor U8958 (N_8958,N_6913,N_5150);
or U8959 (N_8959,N_5956,N_5304);
nor U8960 (N_8960,N_5478,N_6154);
nor U8961 (N_8961,N_5568,N_4017);
nand U8962 (N_8962,N_4370,N_4997);
nand U8963 (N_8963,N_4953,N_5514);
nand U8964 (N_8964,N_6164,N_5810);
or U8965 (N_8965,N_4212,N_5650);
or U8966 (N_8966,N_4573,N_7446);
xnor U8967 (N_8967,N_5282,N_4256);
and U8968 (N_8968,N_6290,N_4752);
nand U8969 (N_8969,N_4429,N_4685);
nor U8970 (N_8970,N_4316,N_5560);
nand U8971 (N_8971,N_4822,N_4859);
xnor U8972 (N_8972,N_4766,N_5004);
nor U8973 (N_8973,N_5040,N_6161);
nand U8974 (N_8974,N_5665,N_7108);
xnor U8975 (N_8975,N_4874,N_4082);
or U8976 (N_8976,N_7232,N_5064);
and U8977 (N_8977,N_5602,N_5374);
nand U8978 (N_8978,N_6073,N_7351);
nand U8979 (N_8979,N_6296,N_6988);
xnor U8980 (N_8980,N_6084,N_6087);
nand U8981 (N_8981,N_6420,N_7155);
nand U8982 (N_8982,N_7313,N_5716);
nor U8983 (N_8983,N_6443,N_4356);
nand U8984 (N_8984,N_5436,N_5557);
nor U8985 (N_8985,N_4700,N_4825);
xnor U8986 (N_8986,N_6075,N_7393);
and U8987 (N_8987,N_4340,N_5542);
or U8988 (N_8988,N_6520,N_7775);
nor U8989 (N_8989,N_7659,N_6739);
nor U8990 (N_8990,N_4364,N_6745);
nor U8991 (N_8991,N_4521,N_5456);
nand U8992 (N_8992,N_5948,N_6662);
or U8993 (N_8993,N_7703,N_4721);
nand U8994 (N_8994,N_7805,N_6184);
or U8995 (N_8995,N_4308,N_6453);
and U8996 (N_8996,N_5446,N_5835);
nor U8997 (N_8997,N_6174,N_4295);
nand U8998 (N_8998,N_4015,N_5856);
nor U8999 (N_8999,N_5217,N_5581);
nand U9000 (N_9000,N_5324,N_4854);
xnor U9001 (N_9001,N_7993,N_6596);
nor U9002 (N_9002,N_4288,N_7990);
xnor U9003 (N_9003,N_6365,N_4726);
nor U9004 (N_9004,N_5682,N_5497);
or U9005 (N_9005,N_5463,N_5783);
nor U9006 (N_9006,N_7103,N_4139);
nor U9007 (N_9007,N_6863,N_4008);
xnor U9008 (N_9008,N_4171,N_4178);
xnor U9009 (N_9009,N_6251,N_6424);
and U9010 (N_9010,N_4966,N_5152);
xor U9011 (N_9011,N_6321,N_4226);
xnor U9012 (N_9012,N_4875,N_6859);
and U9013 (N_9013,N_4397,N_4184);
nor U9014 (N_9014,N_6672,N_7340);
and U9015 (N_9015,N_4194,N_6990);
nor U9016 (N_9016,N_5528,N_7550);
nor U9017 (N_9017,N_7798,N_5047);
and U9018 (N_9018,N_4328,N_5319);
xnor U9019 (N_9019,N_6504,N_5534);
nor U9020 (N_9020,N_7094,N_6586);
xnor U9021 (N_9021,N_5727,N_6311);
nor U9022 (N_9022,N_6706,N_6757);
xnor U9023 (N_9023,N_4584,N_7737);
xor U9024 (N_9024,N_6089,N_6394);
nand U9025 (N_9025,N_6898,N_5213);
or U9026 (N_9026,N_7389,N_4772);
and U9027 (N_9027,N_4504,N_5703);
xor U9028 (N_9028,N_4755,N_6284);
xor U9029 (N_9029,N_5821,N_7013);
nand U9030 (N_9030,N_7145,N_7233);
nand U9031 (N_9031,N_5169,N_7690);
nor U9032 (N_9032,N_4780,N_6310);
nor U9033 (N_9033,N_4427,N_5287);
or U9034 (N_9034,N_5375,N_5792);
nand U9035 (N_9035,N_5506,N_4454);
or U9036 (N_9036,N_7109,N_5395);
or U9037 (N_9037,N_7517,N_7381);
xor U9038 (N_9038,N_5121,N_5303);
or U9039 (N_9039,N_6663,N_5016);
xnor U9040 (N_9040,N_4133,N_5376);
and U9041 (N_9041,N_4701,N_5286);
or U9042 (N_9042,N_5594,N_4580);
and U9043 (N_9043,N_6540,N_4729);
nor U9044 (N_9044,N_4768,N_6564);
nor U9045 (N_9045,N_5569,N_4481);
xnor U9046 (N_9046,N_5765,N_5801);
nor U9047 (N_9047,N_4172,N_4330);
nor U9048 (N_9048,N_6134,N_4423);
xnor U9049 (N_9049,N_4762,N_7735);
nor U9050 (N_9050,N_5798,N_6325);
nor U9051 (N_9051,N_4799,N_6101);
and U9052 (N_9052,N_5026,N_7610);
and U9053 (N_9053,N_4265,N_7814);
xor U9054 (N_9054,N_7411,N_7819);
or U9055 (N_9055,N_7014,N_6014);
nor U9056 (N_9056,N_7179,N_4306);
xnor U9057 (N_9057,N_5759,N_4200);
or U9058 (N_9058,N_7146,N_7522);
xnor U9059 (N_9059,N_7175,N_4357);
and U9060 (N_9060,N_5312,N_4465);
and U9061 (N_9061,N_5907,N_5340);
or U9062 (N_9062,N_7224,N_7196);
nand U9063 (N_9063,N_5901,N_6710);
or U9064 (N_9064,N_7436,N_4033);
nand U9065 (N_9065,N_6333,N_6742);
nor U9066 (N_9066,N_5524,N_4861);
or U9067 (N_9067,N_7478,N_6102);
nor U9068 (N_9068,N_4138,N_7239);
nand U9069 (N_9069,N_4845,N_5717);
or U9070 (N_9070,N_5101,N_4276);
and U9071 (N_9071,N_4442,N_7129);
or U9072 (N_9072,N_4211,N_6448);
or U9073 (N_9073,N_4235,N_5256);
nand U9074 (N_9074,N_6669,N_4439);
or U9075 (N_9075,N_7227,N_6886);
nand U9076 (N_9076,N_4670,N_7682);
xnor U9077 (N_9077,N_6414,N_7422);
xor U9078 (N_9078,N_4722,N_4399);
and U9079 (N_9079,N_6462,N_5860);
xor U9080 (N_9080,N_6234,N_7510);
xor U9081 (N_9081,N_5797,N_5230);
nor U9082 (N_9082,N_5668,N_5582);
or U9083 (N_9083,N_4789,N_6340);
or U9084 (N_9084,N_4490,N_4648);
or U9085 (N_9085,N_7259,N_6689);
nor U9086 (N_9086,N_6358,N_5590);
or U9087 (N_9087,N_5057,N_6401);
xor U9088 (N_9088,N_4620,N_4462);
nand U9089 (N_9089,N_6065,N_7556);
xor U9090 (N_9090,N_4871,N_4889);
xor U9091 (N_9091,N_7007,N_6477);
and U9092 (N_9092,N_5824,N_5895);
nand U9093 (N_9093,N_4091,N_6751);
xor U9094 (N_9094,N_7951,N_4161);
nand U9095 (N_9095,N_6737,N_6936);
xor U9096 (N_9096,N_5234,N_6486);
or U9097 (N_9097,N_4899,N_4819);
nand U9098 (N_9098,N_5074,N_5968);
nor U9099 (N_9099,N_6684,N_4120);
nor U9100 (N_9100,N_5099,N_5843);
nor U9101 (N_9101,N_4561,N_5458);
xor U9102 (N_9102,N_4791,N_7185);
nand U9103 (N_9103,N_5696,N_5186);
and U9104 (N_9104,N_4271,N_7879);
nor U9105 (N_9105,N_6835,N_5030);
xnor U9106 (N_9106,N_5724,N_7176);
or U9107 (N_9107,N_7950,N_4108);
and U9108 (N_9108,N_5088,N_7521);
nand U9109 (N_9109,N_4734,N_4940);
nor U9110 (N_9110,N_4478,N_5367);
xnor U9111 (N_9111,N_7992,N_6502);
or U9112 (N_9112,N_5595,N_7960);
nand U9113 (N_9113,N_7869,N_7205);
xnor U9114 (N_9114,N_5060,N_6368);
and U9115 (N_9115,N_4043,N_6169);
or U9116 (N_9116,N_6125,N_6260);
and U9117 (N_9117,N_4860,N_7165);
nor U9118 (N_9118,N_7638,N_7750);
or U9119 (N_9119,N_5248,N_4470);
xnor U9120 (N_9120,N_6820,N_4890);
nand U9121 (N_9121,N_4443,N_4141);
or U9122 (N_9122,N_4604,N_4893);
or U9123 (N_9123,N_4904,N_4460);
nor U9124 (N_9124,N_4914,N_7927);
or U9125 (N_9125,N_4526,N_6998);
or U9126 (N_9126,N_4711,N_7935);
nand U9127 (N_9127,N_6057,N_7144);
or U9128 (N_9128,N_4160,N_7226);
nand U9129 (N_9129,N_7817,N_5738);
or U9130 (N_9130,N_6758,N_7900);
nor U9131 (N_9131,N_7076,N_4520);
or U9132 (N_9132,N_5624,N_4204);
nor U9133 (N_9133,N_4219,N_6407);
and U9134 (N_9134,N_5216,N_7966);
and U9135 (N_9135,N_7619,N_5462);
nor U9136 (N_9136,N_6488,N_4499);
nor U9137 (N_9137,N_7783,N_4329);
and U9138 (N_9138,N_5570,N_6733);
and U9139 (N_9139,N_6974,N_5468);
and U9140 (N_9140,N_7649,N_7160);
nand U9141 (N_9141,N_7561,N_4434);
nand U9142 (N_9142,N_4323,N_5846);
and U9143 (N_9143,N_6907,N_6741);
or U9144 (N_9144,N_6052,N_4514);
nand U9145 (N_9145,N_7998,N_7342);
nand U9146 (N_9146,N_7100,N_6092);
and U9147 (N_9147,N_4624,N_7082);
and U9148 (N_9148,N_7061,N_6505);
nor U9149 (N_9149,N_6068,N_5142);
and U9150 (N_9150,N_7435,N_4895);
xnor U9151 (N_9151,N_7637,N_7123);
xor U9152 (N_9152,N_7627,N_7437);
xor U9153 (N_9153,N_6109,N_5566);
nand U9154 (N_9154,N_4868,N_6553);
xor U9155 (N_9155,N_6643,N_4090);
nor U9156 (N_9156,N_7938,N_4225);
nand U9157 (N_9157,N_4709,N_7811);
and U9158 (N_9158,N_4412,N_5315);
and U9159 (N_9159,N_6350,N_7261);
xor U9160 (N_9160,N_4802,N_5505);
nor U9161 (N_9161,N_4129,N_4778);
nor U9162 (N_9162,N_4804,N_4512);
nor U9163 (N_9163,N_7423,N_5079);
and U9164 (N_9164,N_5442,N_5491);
nand U9165 (N_9165,N_6227,N_7491);
and U9166 (N_9166,N_7621,N_7788);
or U9167 (N_9167,N_4549,N_7871);
and U9168 (N_9168,N_6309,N_5941);
and U9169 (N_9169,N_4293,N_6773);
xor U9170 (N_9170,N_6695,N_4047);
nand U9171 (N_9171,N_5666,N_4137);
or U9172 (N_9172,N_5253,N_7511);
or U9173 (N_9173,N_7318,N_7439);
xnor U9174 (N_9174,N_6012,N_4590);
and U9175 (N_9175,N_7847,N_7248);
xnor U9176 (N_9176,N_7752,N_4215);
xor U9177 (N_9177,N_7774,N_5555);
or U9178 (N_9178,N_4816,N_4459);
and U9179 (N_9179,N_6069,N_6201);
xnor U9180 (N_9180,N_5755,N_6743);
nand U9181 (N_9181,N_5644,N_4820);
or U9182 (N_9182,N_4051,N_5218);
and U9183 (N_9183,N_5531,N_4457);
nor U9184 (N_9184,N_4094,N_6759);
nor U9185 (N_9185,N_5198,N_6995);
or U9186 (N_9186,N_4818,N_6521);
or U9187 (N_9187,N_5786,N_4210);
or U9188 (N_9188,N_7917,N_5685);
xor U9189 (N_9189,N_4641,N_6352);
and U9190 (N_9190,N_5188,N_5011);
or U9191 (N_9191,N_6262,N_7586);
nand U9192 (N_9192,N_6685,N_6649);
nand U9193 (N_9193,N_6503,N_6136);
or U9194 (N_9194,N_5166,N_7837);
and U9195 (N_9195,N_4842,N_5180);
or U9196 (N_9196,N_5279,N_4471);
xnor U9197 (N_9197,N_4199,N_4246);
and U9198 (N_9198,N_6362,N_6732);
nand U9199 (N_9199,N_6870,N_7970);
xor U9200 (N_9200,N_6066,N_5053);
nand U9201 (N_9201,N_6388,N_4548);
or U9202 (N_9202,N_4657,N_5632);
nor U9203 (N_9203,N_5731,N_7386);
nand U9204 (N_9204,N_4686,N_4545);
and U9205 (N_9205,N_6983,N_4938);
xor U9206 (N_9206,N_7832,N_4668);
nand U9207 (N_9207,N_5733,N_5678);
nor U9208 (N_9208,N_5811,N_6579);
nor U9209 (N_9209,N_6266,N_6046);
nand U9210 (N_9210,N_6211,N_4065);
nor U9211 (N_9211,N_6082,N_4888);
and U9212 (N_9212,N_5806,N_4250);
xor U9213 (N_9213,N_4004,N_7492);
nor U9214 (N_9214,N_5354,N_7501);
xnor U9215 (N_9215,N_5305,N_4759);
and U9216 (N_9216,N_6213,N_6118);
nand U9217 (N_9217,N_4100,N_6151);
and U9218 (N_9218,N_6206,N_4503);
or U9219 (N_9219,N_4779,N_6959);
nor U9220 (N_9220,N_4187,N_4742);
xor U9221 (N_9221,N_4378,N_7461);
nand U9222 (N_9222,N_5388,N_4523);
xor U9223 (N_9223,N_6844,N_5453);
xnor U9224 (N_9224,N_6050,N_6264);
nor U9225 (N_9225,N_6332,N_4674);
xor U9226 (N_9226,N_6008,N_4977);
or U9227 (N_9227,N_5081,N_7301);
nand U9228 (N_9228,N_4349,N_6828);
and U9229 (N_9229,N_5471,N_5523);
xor U9230 (N_9230,N_4455,N_4277);
nor U9231 (N_9231,N_7981,N_5103);
nand U9232 (N_9232,N_6954,N_4314);
nor U9233 (N_9233,N_5747,N_7484);
nand U9234 (N_9234,N_6731,N_4273);
xor U9235 (N_9235,N_4942,N_6177);
or U9236 (N_9236,N_5427,N_6484);
nor U9237 (N_9237,N_4227,N_6183);
nand U9238 (N_9238,N_5448,N_5337);
and U9239 (N_9239,N_5071,N_7164);
nor U9240 (N_9240,N_5689,N_6207);
nor U9241 (N_9241,N_7956,N_5032);
nand U9242 (N_9242,N_5196,N_4763);
and U9243 (N_9243,N_5855,N_7288);
or U9244 (N_9244,N_7159,N_5494);
nand U9245 (N_9245,N_5601,N_4391);
xor U9246 (N_9246,N_7892,N_6383);
nor U9247 (N_9247,N_6635,N_6556);
nand U9248 (N_9248,N_5369,N_5317);
nor U9249 (N_9249,N_6543,N_5084);
nand U9250 (N_9250,N_5611,N_7079);
nand U9251 (N_9251,N_6636,N_4840);
or U9252 (N_9252,N_7133,N_4853);
xor U9253 (N_9253,N_5140,N_7688);
nand U9254 (N_9254,N_6982,N_4585);
nor U9255 (N_9255,N_5854,N_4588);
and U9256 (N_9256,N_4848,N_4419);
xor U9257 (N_9257,N_4828,N_7353);
xnor U9258 (N_9258,N_5700,N_7667);
xor U9259 (N_9259,N_5082,N_5631);
nor U9260 (N_9260,N_5338,N_5576);
nor U9261 (N_9261,N_6074,N_6658);
xor U9262 (N_9262,N_6282,N_5899);
and U9263 (N_9263,N_7204,N_6523);
xor U9264 (N_9264,N_6841,N_5620);
or U9265 (N_9265,N_4905,N_5420);
and U9266 (N_9266,N_5974,N_4963);
nand U9267 (N_9267,N_7719,N_5884);
nor U9268 (N_9268,N_5825,N_5153);
nand U9269 (N_9269,N_4509,N_7366);
nand U9270 (N_9270,N_4717,N_6728);
xnor U9271 (N_9271,N_4599,N_6657);
nor U9272 (N_9272,N_5087,N_6106);
nor U9273 (N_9273,N_6374,N_7557);
and U9274 (N_9274,N_5151,N_5393);
xor U9275 (N_9275,N_4894,N_4597);
or U9276 (N_9276,N_5459,N_4480);
and U9277 (N_9277,N_7606,N_5226);
nor U9278 (N_9278,N_4361,N_5522);
and U9279 (N_9279,N_5980,N_6440);
xnor U9280 (N_9280,N_7946,N_6098);
xnor U9281 (N_9281,N_6716,N_7281);
nor U9282 (N_9282,N_7372,N_4468);
xor U9283 (N_9283,N_4382,N_5687);
nand U9284 (N_9284,N_6237,N_6028);
and U9285 (N_9285,N_6847,N_7853);
and U9286 (N_9286,N_4140,N_5780);
nand U9287 (N_9287,N_7137,N_4958);
nand U9288 (N_9288,N_6230,N_6250);
nand U9289 (N_9289,N_6606,N_4068);
or U9290 (N_9290,N_7290,N_7841);
and U9291 (N_9291,N_7062,N_5829);
nand U9292 (N_9292,N_5190,N_7800);
nor U9293 (N_9293,N_6720,N_7475);
or U9294 (N_9294,N_6086,N_5966);
nand U9295 (N_9295,N_5482,N_7699);
nor U9296 (N_9296,N_7040,N_4495);
or U9297 (N_9297,N_5297,N_4131);
xnor U9298 (N_9298,N_6707,N_7420);
and U9299 (N_9299,N_6359,N_7856);
xor U9300 (N_9300,N_4785,N_4450);
or U9301 (N_9301,N_4135,N_5222);
nor U9302 (N_9302,N_6760,N_6198);
or U9303 (N_9303,N_7655,N_4379);
xnor U9304 (N_9304,N_6683,N_6150);
nor U9305 (N_9305,N_5961,N_6984);
nand U9306 (N_9306,N_6921,N_6670);
and U9307 (N_9307,N_4989,N_6280);
nor U9308 (N_9308,N_7594,N_5571);
nand U9309 (N_9309,N_7424,N_7315);
nor U9310 (N_9310,N_5118,N_4826);
nand U9311 (N_9311,N_4307,N_6399);
and U9312 (N_9312,N_7283,N_6055);
and U9313 (N_9313,N_6777,N_5501);
nor U9314 (N_9314,N_5663,N_7663);
or U9315 (N_9315,N_6034,N_7833);
xnor U9316 (N_9316,N_4489,N_4979);
nor U9317 (N_9317,N_5508,N_7282);
nor U9318 (N_9318,N_5352,N_4284);
and U9319 (N_9319,N_6541,N_7397);
xnor U9320 (N_9320,N_7786,N_5368);
nand U9321 (N_9321,N_5193,N_4792);
and U9322 (N_9322,N_7431,N_7889);
xor U9323 (N_9323,N_6241,N_7957);
or U9324 (N_9324,N_6967,N_4827);
nand U9325 (N_9325,N_5335,N_6302);
and U9326 (N_9326,N_4865,N_7470);
or U9327 (N_9327,N_6981,N_5386);
nand U9328 (N_9328,N_5865,N_7371);
nand U9329 (N_9329,N_7343,N_5629);
xnor U9330 (N_9330,N_6550,N_5702);
or U9331 (N_9331,N_5944,N_5519);
or U9332 (N_9332,N_7564,N_7810);
and U9333 (N_9333,N_7015,N_4388);
and U9334 (N_9334,N_7605,N_7092);
and U9335 (N_9335,N_4563,N_5122);
nand U9336 (N_9336,N_5537,N_4088);
or U9337 (N_9337,N_5461,N_5965);
xnor U9338 (N_9338,N_4939,N_6893);
xor U9339 (N_9339,N_4999,N_5507);
nor U9340 (N_9340,N_5859,N_4159);
or U9341 (N_9341,N_6167,N_6501);
nand U9342 (N_9342,N_7928,N_6819);
nor U9343 (N_9343,N_7444,N_7042);
xor U9344 (N_9344,N_5713,N_6204);
nor U9345 (N_9345,N_4964,N_6617);
nand U9346 (N_9346,N_5334,N_7603);
and U9347 (N_9347,N_5042,N_7012);
nor U9348 (N_9348,N_6141,N_4775);
and U9349 (N_9349,N_7864,N_6032);
nand U9350 (N_9350,N_4119,N_6831);
and U9351 (N_9351,N_7380,N_4776);
xnor U9352 (N_9352,N_5642,N_6559);
nand U9353 (N_9353,N_7483,N_6083);
or U9354 (N_9354,N_6100,N_5550);
or U9355 (N_9355,N_6021,N_5864);
nor U9356 (N_9356,N_5946,N_4012);
nand U9357 (N_9357,N_4864,N_4675);
xnor U9358 (N_9358,N_6466,N_4918);
nand U9359 (N_9359,N_5410,N_7453);
or U9360 (N_9360,N_5250,N_6722);
or U9361 (N_9361,N_5430,N_5596);
or U9362 (N_9362,N_6356,N_6646);
or U9363 (N_9363,N_6642,N_6794);
or U9364 (N_9364,N_7830,N_4817);
and U9365 (N_9365,N_7681,N_4609);
and U9366 (N_9366,N_4902,N_7504);
nor U9367 (N_9367,N_6023,N_5477);
xor U9368 (N_9368,N_5789,N_5035);
and U9369 (N_9369,N_7915,N_5861);
nand U9370 (N_9370,N_6114,N_6218);
nand U9371 (N_9371,N_7421,N_4154);
xor U9372 (N_9372,N_5043,N_6781);
nor U9373 (N_9373,N_7657,N_4125);
nor U9374 (N_9374,N_5982,N_5767);
nand U9375 (N_9375,N_5972,N_7818);
nand U9376 (N_9376,N_4238,N_4528);
nor U9377 (N_9377,N_6002,N_4344);
nor U9378 (N_9378,N_4534,N_4395);
xor U9379 (N_9379,N_4192,N_6482);
or U9380 (N_9380,N_5530,N_5730);
xnor U9381 (N_9381,N_5782,N_4672);
xnor U9382 (N_9382,N_5714,N_6327);
nor U9383 (N_9383,N_5719,N_4467);
nand U9384 (N_9384,N_4870,N_5548);
or U9385 (N_9385,N_6349,N_4177);
nand U9386 (N_9386,N_5416,N_4949);
or U9387 (N_9387,N_7978,N_4156);
nand U9388 (N_9388,N_6887,N_5473);
or U9389 (N_9389,N_6483,N_4181);
xnor U9390 (N_9390,N_7030,N_6430);
nor U9391 (N_9391,N_5358,N_5962);
nand U9392 (N_9392,N_6105,N_4513);
or U9393 (N_9393,N_4735,N_7099);
nand U9394 (N_9394,N_4663,N_7825);
nor U9395 (N_9395,N_5063,N_4376);
nor U9396 (N_9396,N_4074,N_4619);
xor U9397 (N_9397,N_4557,N_4058);
nand U9398 (N_9398,N_7875,N_4558);
nand U9399 (N_9399,N_4369,N_7872);
or U9400 (N_9400,N_4595,N_5379);
nor U9401 (N_9401,N_5540,N_5293);
and U9402 (N_9402,N_6200,N_5294);
nor U9403 (N_9403,N_7271,N_5007);
or U9404 (N_9404,N_6051,N_6769);
xor U9405 (N_9405,N_6531,N_5451);
and U9406 (N_9406,N_7297,N_7881);
xor U9407 (N_9407,N_7081,N_4260);
nand U9408 (N_9408,N_6355,N_7903);
nand U9409 (N_9409,N_6830,N_6874);
nand U9410 (N_9410,N_4071,N_4244);
and U9411 (N_9411,N_5183,N_6703);
nor U9412 (N_9412,N_7685,N_6450);
and U9413 (N_9413,N_7707,N_6451);
nand U9414 (N_9414,N_4856,N_7095);
xor U9415 (N_9415,N_4279,N_7097);
nand U9416 (N_9416,N_7341,N_7432);
and U9417 (N_9417,N_5516,N_4656);
xnor U9418 (N_9418,N_5202,N_6906);
nor U9419 (N_9419,N_4708,N_7665);
nand U9420 (N_9420,N_6659,N_4064);
and U9421 (N_9421,N_7997,N_6188);
and U9422 (N_9422,N_5659,N_6156);
or U9423 (N_9423,N_5476,N_5720);
or U9424 (N_9424,N_7577,N_4030);
or U9425 (N_9425,N_6493,N_5574);
or U9426 (N_9426,N_6209,N_6747);
or U9427 (N_9427,N_7481,N_7279);
xor U9428 (N_9428,N_5083,N_6843);
xor U9429 (N_9429,N_6753,N_5809);
nor U9430 (N_9430,N_7512,N_6447);
nor U9431 (N_9431,N_6616,N_4510);
or U9432 (N_9432,N_5580,N_7914);
and U9433 (N_9433,N_5235,N_6821);
or U9434 (N_9434,N_5288,N_5108);
or U9435 (N_9435,N_6335,N_6938);
nor U9436 (N_9436,N_7572,N_5958);
nand U9437 (N_9437,N_5627,N_6248);
or U9438 (N_9438,N_4603,N_5905);
xnor U9439 (N_9439,N_7021,N_7622);
nand U9440 (N_9440,N_4919,N_6861);
or U9441 (N_9441,N_6085,N_6920);
and U9442 (N_9442,N_4981,N_4066);
xor U9443 (N_9443,N_6481,N_4714);
and U9444 (N_9444,N_5957,N_4466);
or U9445 (N_9445,N_5922,N_6458);
or U9446 (N_9446,N_7732,N_5999);
or U9447 (N_9447,N_7172,N_5041);
nand U9448 (N_9448,N_5284,N_5769);
nor U9449 (N_9449,N_4608,N_4832);
and U9450 (N_9450,N_6210,N_6470);
nand U9451 (N_9451,N_7005,N_5935);
nor U9452 (N_9452,N_6117,N_6246);
nand U9453 (N_9453,N_7979,N_5837);
nand U9454 (N_9454,N_7338,N_5024);
nor U9455 (N_9455,N_6265,N_4596);
xor U9456 (N_9456,N_5085,N_6093);
or U9457 (N_9457,N_6380,N_5158);
nand U9458 (N_9458,N_6779,N_7953);
xor U9459 (N_9459,N_4044,N_6605);
or U9460 (N_9460,N_4476,N_5050);
nor U9461 (N_9461,N_4373,N_6945);
xnor U9462 (N_9462,N_4884,N_6787);
or U9463 (N_9463,N_5766,N_7523);
or U9464 (N_9464,N_5493,N_4440);
nand U9465 (N_9465,N_5888,N_5460);
nand U9466 (N_9466,N_4965,N_7396);
xnor U9467 (N_9467,N_4002,N_4313);
xor U9468 (N_9468,N_6879,N_6912);
and U9469 (N_9469,N_5833,N_5438);
or U9470 (N_9470,N_5009,N_6480);
or U9471 (N_9471,N_6331,N_7149);
nor U9472 (N_9472,N_6699,N_6419);
and U9473 (N_9473,N_7592,N_4315);
nor U9474 (N_9474,N_7006,N_7462);
xor U9475 (N_9475,N_6072,N_6561);
nor U9476 (N_9476,N_5439,N_6919);
nand U9477 (N_9477,N_7375,N_4807);
nor U9478 (N_9478,N_7764,N_5225);
and U9479 (N_9479,N_6455,N_4437);
nor U9480 (N_9480,N_5619,N_4103);
nand U9481 (N_9481,N_6991,N_7031);
xor U9482 (N_9482,N_4428,N_5850);
or U9483 (N_9483,N_5308,N_5873);
nand U9484 (N_9484,N_5583,N_7009);
or U9485 (N_9485,N_6138,N_4508);
or U9486 (N_9486,N_4622,N_5309);
or U9487 (N_9487,N_7773,N_7169);
or U9488 (N_9488,N_4625,N_5147);
nand U9489 (N_9489,N_7954,N_6810);
or U9490 (N_9490,N_6875,N_6570);
and U9491 (N_9491,N_5834,N_4655);
xnor U9492 (N_9492,N_5378,N_5614);
nor U9493 (N_9493,N_5215,N_4898);
nand U9494 (N_9494,N_5257,N_4180);
xnor U9495 (N_9495,N_6097,N_4551);
and U9496 (N_9496,N_4751,N_7150);
and U9497 (N_9497,N_6962,N_7582);
nand U9498 (N_9498,N_4317,N_6590);
or U9499 (N_9499,N_6037,N_5020);
xnor U9500 (N_9500,N_6354,N_4809);
and U9501 (N_9501,N_4056,N_6515);
nor U9502 (N_9502,N_5913,N_7370);
nand U9503 (N_9503,N_4758,N_4582);
xnor U9504 (N_9504,N_7575,N_4552);
or U9505 (N_9505,N_6824,N_7258);
nand U9506 (N_9506,N_6846,N_4850);
xnor U9507 (N_9507,N_5945,N_6544);
and U9508 (N_9508,N_5647,N_7157);
and U9509 (N_9509,N_7477,N_5065);
nand U9510 (N_9510,N_5173,N_7443);
or U9511 (N_9511,N_5692,N_4554);
nand U9512 (N_9512,N_7525,N_6381);
xor U9513 (N_9513,N_6229,N_6273);
and U9514 (N_9514,N_6000,N_4978);
and U9515 (N_9515,N_4649,N_7747);
or U9516 (N_9516,N_4416,N_6604);
nor U9517 (N_9517,N_4233,N_5883);
nand U9518 (N_9518,N_4614,N_4944);
nor U9519 (N_9519,N_6217,N_7029);
nand U9520 (N_9520,N_6187,N_6788);
or U9521 (N_9521,N_6956,N_6258);
nor U9522 (N_9522,N_7844,N_5543);
and U9523 (N_9523,N_4300,N_6955);
and U9524 (N_9524,N_5613,N_7255);
nand U9525 (N_9525,N_4538,N_5266);
and U9526 (N_9526,N_5360,N_4623);
xor U9527 (N_9527,N_5241,N_7803);
xnor U9528 (N_9528,N_7855,N_4591);
or U9529 (N_9529,N_5802,N_5245);
nand U9530 (N_9530,N_4424,N_6377);
xnor U9531 (N_9531,N_4516,N_5842);
xnor U9532 (N_9532,N_4298,N_6871);
xnor U9533 (N_9533,N_7921,N_6231);
nand U9534 (N_9534,N_5814,N_5137);
nor U9535 (N_9535,N_6972,N_4858);
xnor U9536 (N_9536,N_4087,N_5464);
nand U9537 (N_9537,N_7112,N_4222);
nor U9538 (N_9538,N_5124,N_7002);
xnor U9539 (N_9539,N_6463,N_5909);
nand U9540 (N_9540,N_6608,N_5575);
and U9541 (N_9541,N_5885,N_7384);
nand U9542 (N_9542,N_6868,N_5385);
xnor U9543 (N_9543,N_4575,N_6917);
xor U9544 (N_9544,N_6627,N_4095);
and U9545 (N_9545,N_7580,N_6123);
xor U9546 (N_9546,N_7552,N_7194);
or U9547 (N_9547,N_4282,N_4838);
or U9548 (N_9548,N_4123,N_4372);
nand U9549 (N_9549,N_5658,N_7539);
xor U9550 (N_9550,N_7333,N_6908);
nand U9551 (N_9551,N_6361,N_6107);
nor U9552 (N_9552,N_6510,N_7328);
or U9553 (N_9553,N_7874,N_7895);
or U9554 (N_9554,N_7730,N_7760);
nor U9555 (N_9555,N_7860,N_7069);
xor U9556 (N_9556,N_6960,N_7189);
nand U9557 (N_9557,N_7300,N_5981);
nor U9558 (N_9558,N_7231,N_4985);
xnor U9559 (N_9559,N_5994,N_4241);
nand U9560 (N_9560,N_4239,N_6927);
nor U9561 (N_9561,N_4849,N_5089);
nor U9562 (N_9562,N_4486,N_6300);
nor U9563 (N_9563,N_4127,N_5960);
or U9564 (N_9564,N_4943,N_6514);
and U9565 (N_9565,N_4209,N_5499);
or U9566 (N_9566,N_7901,N_4262);
or U9567 (N_9567,N_6977,N_7633);
xor U9568 (N_9568,N_4877,N_6214);
nand U9569 (N_9569,N_6813,N_6952);
or U9570 (N_9570,N_6996,N_4367);
nand U9571 (N_9571,N_7785,N_7269);
xor U9572 (N_9572,N_7273,N_6271);
and U9573 (N_9573,N_4352,N_7893);
nand U9574 (N_9574,N_7835,N_4240);
and U9575 (N_9575,N_6281,N_4409);
or U9576 (N_9576,N_5673,N_4078);
xnor U9577 (N_9577,N_6479,N_7852);
or U9578 (N_9578,N_6601,N_7034);
xnor U9579 (N_9579,N_6367,N_4248);
xor U9580 (N_9580,N_6245,N_6303);
and U9581 (N_9581,N_4000,N_4198);
nor U9582 (N_9582,N_5419,N_5159);
nor U9583 (N_9583,N_5033,N_4097);
and U9584 (N_9584,N_6957,N_6884);
nor U9585 (N_9585,N_6432,N_4990);
nor U9586 (N_9586,N_6146,N_5670);
or U9587 (N_9587,N_6971,N_4377);
nor U9588 (N_9588,N_5409,N_6205);
nor U9589 (N_9589,N_5342,N_6094);
nand U9590 (N_9590,N_6718,N_5805);
or U9591 (N_9591,N_7624,N_4024);
or U9592 (N_9592,N_4564,N_7664);
and U9593 (N_9593,N_5149,N_4581);
and U9594 (N_9594,N_4485,N_6625);
and U9595 (N_9595,N_7931,N_6494);
or U9596 (N_9596,N_7151,N_7158);
or U9597 (N_9597,N_7797,N_5397);
nand U9598 (N_9598,N_5919,N_7989);
and U9599 (N_9599,N_4116,N_7494);
and U9600 (N_9600,N_6650,N_7267);
nand U9601 (N_9601,N_7590,N_6226);
or U9602 (N_9602,N_7758,N_5336);
nand U9603 (N_9603,N_4243,N_4537);
xor U9604 (N_9604,N_7430,N_7244);
or U9605 (N_9605,N_5970,N_5205);
nand U9606 (N_9606,N_6944,N_4355);
and U9607 (N_9607,N_5480,N_6110);
nor U9608 (N_9608,N_4712,N_6222);
and U9609 (N_9609,N_5585,N_4366);
xnor U9610 (N_9610,N_6687,N_4743);
nand U9611 (N_9611,N_4970,N_7651);
or U9612 (N_9612,N_4522,N_5157);
nor U9613 (N_9613,N_6465,N_4810);
nand U9614 (N_9614,N_7264,N_5012);
or U9615 (N_9615,N_4896,N_7292);
nor U9616 (N_9616,N_4761,N_5857);
xor U9617 (N_9617,N_4042,N_5254);
nand U9618 (N_9618,N_5077,N_7024);
and U9619 (N_9619,N_6914,N_7043);
nand U9620 (N_9620,N_7964,N_4342);
or U9621 (N_9621,N_4719,N_7221);
and U9622 (N_9622,N_4841,N_5586);
nand U9623 (N_9623,N_6030,N_6435);
nor U9624 (N_9624,N_4987,N_7751);
nand U9625 (N_9625,N_7256,N_6725);
or U9626 (N_9626,N_7409,N_5795);
nand U9627 (N_9627,N_6121,N_7608);
nor U9628 (N_9628,N_5558,N_7625);
or U9629 (N_9629,N_4501,N_4715);
or U9630 (N_9630,N_5472,N_7618);
nor U9631 (N_9631,N_7975,N_5208);
nand U9632 (N_9632,N_5770,N_7496);
xnor U9633 (N_9633,N_4479,N_7965);
xor U9634 (N_9634,N_6522,N_7460);
xor U9635 (N_9635,N_5027,N_6811);
nand U9636 (N_9636,N_6724,N_5711);
nand U9637 (N_9637,N_7344,N_5301);
xor U9638 (N_9638,N_7967,N_5174);
nor U9639 (N_9639,N_4660,N_6883);
nand U9640 (N_9640,N_4667,N_7337);
nand U9641 (N_9641,N_6024,N_7263);
and U9642 (N_9642,N_7119,N_7088);
nand U9643 (N_9643,N_7285,N_7171);
and U9644 (N_9644,N_7646,N_7636);
or U9645 (N_9645,N_4945,N_7017);
nor U9646 (N_9646,N_4913,N_7674);
xnor U9647 (N_9647,N_7548,N_5228);
xnor U9648 (N_9648,N_4957,N_5694);
nand U9649 (N_9649,N_7358,N_7487);
and U9650 (N_9650,N_4464,N_5800);
or U9651 (N_9651,N_6837,N_7468);
and U9652 (N_9652,N_6297,N_7808);
or U9653 (N_9653,N_4530,N_4264);
nand U9654 (N_9654,N_5513,N_4694);
xnor U9655 (N_9655,N_6423,N_7939);
or U9656 (N_9656,N_6721,N_6951);
nor U9657 (N_9657,N_5058,N_4576);
nand U9658 (N_9658,N_4863,N_6304);
or U9659 (N_9659,N_6973,N_7793);
nand U9660 (N_9660,N_6557,N_5729);
nor U9661 (N_9661,N_6937,N_6445);
and U9662 (N_9662,N_4968,N_5656);
and U9663 (N_9663,N_4249,N_4592);
and U9664 (N_9664,N_7976,N_7829);
or U9665 (N_9665,N_5244,N_4084);
and U9666 (N_9666,N_6671,N_6115);
nand U9667 (N_9667,N_6869,N_4916);
or U9668 (N_9668,N_4255,N_4680);
or U9669 (N_9669,N_5758,N_5380);
nand U9670 (N_9670,N_7429,N_6326);
nor U9671 (N_9671,N_6313,N_6518);
xnor U9672 (N_9672,N_7532,N_5639);
and U9673 (N_9673,N_7121,N_6112);
nor U9674 (N_9674,N_4099,N_6305);
and U9675 (N_9675,N_5093,N_6143);
or U9676 (N_9676,N_6459,N_6027);
and U9677 (N_9677,N_4359,N_7401);
or U9678 (N_9678,N_7115,N_7293);
xnor U9679 (N_9679,N_7085,N_5554);
xnor U9680 (N_9680,N_6876,N_7178);
nor U9681 (N_9681,N_4274,N_7128);
or U9682 (N_9682,N_6397,N_7714);
nor U9683 (N_9683,N_6626,N_6619);
nand U9684 (N_9684,N_7390,N_7727);
and U9685 (N_9685,N_7325,N_7438);
or U9686 (N_9686,N_5774,N_5831);
xor U9687 (N_9687,N_6259,N_4073);
nand U9688 (N_9688,N_6436,N_6993);
and U9689 (N_9689,N_6337,N_6389);
and U9690 (N_9690,N_7122,N_5661);
or U9691 (N_9691,N_6317,N_7827);
xnor U9692 (N_9692,N_5329,N_5561);
xnor U9693 (N_9693,N_6189,N_4092);
xnor U9694 (N_9694,N_5437,N_6816);
xor U9695 (N_9695,N_4433,N_4929);
and U9696 (N_9696,N_5565,N_5239);
or U9697 (N_9697,N_4784,N_6836);
nand U9698 (N_9698,N_6736,N_6858);
xnor U9699 (N_9699,N_7060,N_4290);
nand U9700 (N_9700,N_4777,N_5021);
and U9701 (N_9701,N_6567,N_7926);
or U9702 (N_9702,N_4774,N_6594);
nor U9703 (N_9703,N_7180,N_5778);
and U9704 (N_9704,N_4469,N_7958);
nand U9705 (N_9705,N_6364,N_5616);
xnor U9706 (N_9706,N_7723,N_4122);
and U9707 (N_9707,N_7047,N_6941);
nor U9708 (N_9708,N_6620,N_7418);
or U9709 (N_9709,N_6746,N_7623);
xor U9710 (N_9710,N_7001,N_6849);
xor U9711 (N_9711,N_5698,N_7080);
nor U9712 (N_9712,N_6798,N_6473);
xor U9713 (N_9713,N_6261,N_4662);
or U9714 (N_9714,N_6148,N_5069);
and U9715 (N_9715,N_6314,N_5300);
or U9716 (N_9716,N_4831,N_6378);
or U9717 (N_9717,N_7214,N_7311);
and U9718 (N_9718,N_7086,N_6928);
nand U9719 (N_9719,N_6391,N_6346);
nor U9720 (N_9720,N_6610,N_5844);
nand U9721 (N_9721,N_4353,N_6274);
nor U9722 (N_9722,N_4398,N_6750);
and U9723 (N_9723,N_7363,N_5932);
or U9724 (N_9724,N_4190,N_5092);
nand U9725 (N_9725,N_6360,N_4531);
nand U9726 (N_9726,N_7784,N_5080);
and U9727 (N_9727,N_6221,N_5045);
and U9728 (N_9728,N_5951,N_4230);
nor U9729 (N_9729,N_7943,N_4937);
and U9730 (N_9730,N_5407,N_6754);
nand U9731 (N_9731,N_5930,N_6791);
or U9732 (N_9732,N_5893,N_4543);
xor U9733 (N_9733,N_4380,N_5377);
or U9734 (N_9734,N_6124,N_5115);
or U9735 (N_9735,N_7675,N_7754);
or U9736 (N_9736,N_7559,N_5521);
nand U9737 (N_9737,N_5500,N_7249);
nand U9738 (N_9738,N_5804,N_7859);
xnor U9739 (N_9739,N_5306,N_7693);
nor U9740 (N_9740,N_6452,N_6384);
xnor U9741 (N_9741,N_4147,N_4934);
or U9742 (N_9742,N_4069,N_5346);
xnor U9743 (N_9743,N_4179,N_6078);
xor U9744 (N_9744,N_6005,N_7093);
or U9745 (N_9745,N_7757,N_6336);
nor U9746 (N_9746,N_6599,N_5971);
nor U9747 (N_9747,N_5341,N_7347);
nor U9748 (N_9748,N_4565,N_7769);
nand U9749 (N_9749,N_4642,N_7897);
and U9750 (N_9750,N_7670,N_6403);
nor U9751 (N_9751,N_6547,N_5182);
or U9752 (N_9752,N_6299,N_4907);
and U9753 (N_9753,N_6527,N_4730);
and U9754 (N_9754,N_5923,N_4560);
nand U9755 (N_9755,N_5764,N_7220);
nand U9756 (N_9756,N_4336,N_7252);
and U9757 (N_9757,N_6179,N_6120);
and U9758 (N_9758,N_6243,N_4400);
nor U9759 (N_9759,N_7925,N_7124);
nand U9760 (N_9760,N_5003,N_7098);
xnor U9761 (N_9761,N_5046,N_5681);
and U9762 (N_9762,N_6832,N_7516);
xnor U9763 (N_9763,N_6153,N_5667);
xnor U9764 (N_9764,N_7809,N_5939);
or U9765 (N_9765,N_7467,N_5131);
or U9766 (N_9766,N_5104,N_7051);
or U9767 (N_9767,N_7896,N_5927);
and U9768 (N_9768,N_6489,N_6730);
nor U9769 (N_9769,N_6287,N_5148);
nor U9770 (N_9770,N_4569,N_6454);
nand U9771 (N_9771,N_6158,N_4418);
or U9772 (N_9772,N_7322,N_7474);
xnor U9773 (N_9773,N_7170,N_4163);
nand U9774 (N_9774,N_4872,N_7054);
nand U9775 (N_9775,N_5203,N_4343);
xnor U9776 (N_9776,N_6225,N_5330);
nor U9777 (N_9777,N_7465,N_5916);
nand U9778 (N_9778,N_6600,N_7858);
and U9779 (N_9779,N_7698,N_6558);
or U9780 (N_9780,N_4691,N_7450);
and U9781 (N_9781,N_7209,N_5351);
or U9782 (N_9782,N_7761,N_7373);
nand U9783 (N_9783,N_7530,N_7417);
and U9784 (N_9784,N_7247,N_6756);
xor U9785 (N_9785,N_4319,N_5890);
nand U9786 (N_9786,N_7937,N_5474);
or U9787 (N_9787,N_5605,N_5643);
nand U9788 (N_9788,N_4037,N_5943);
nand U9789 (N_9789,N_4562,N_6764);
or U9790 (N_9790,N_6766,N_5623);
xor U9791 (N_9791,N_6279,N_4045);
xnor U9792 (N_9792,N_7312,N_4292);
or U9793 (N_9793,N_7867,N_5853);
and U9794 (N_9794,N_5143,N_6536);
and U9795 (N_9795,N_6803,N_4272);
xnor U9796 (N_9796,N_7074,N_6328);
and U9797 (N_9797,N_4583,N_4834);
and U9798 (N_9798,N_4048,N_7139);
nor U9799 (N_9799,N_7596,N_7660);
nand U9800 (N_9800,N_6679,N_5564);
nor U9801 (N_9801,N_6062,N_7406);
xor U9802 (N_9802,N_4676,N_4408);
or U9803 (N_9803,N_5261,N_5634);
xor U9804 (N_9804,N_4607,N_4132);
nor U9805 (N_9805,N_4054,N_4261);
or U9806 (N_9806,N_6612,N_4518);
nand U9807 (N_9807,N_7746,N_7075);
nand U9808 (N_9808,N_7794,N_5791);
nor U9809 (N_9809,N_7831,N_6640);
xnor U9810 (N_9810,N_5752,N_7631);
nor U9811 (N_9811,N_4883,N_7141);
or U9812 (N_9812,N_5726,N_5830);
xor U9813 (N_9813,N_5399,N_6442);
nor U9814 (N_9814,N_5858,N_5751);
nor U9815 (N_9815,N_7763,N_5394);
and U9816 (N_9816,N_5211,N_6038);
xor U9817 (N_9817,N_5908,N_7033);
xnor U9818 (N_9818,N_5771,N_4688);
and U9819 (N_9819,N_5144,N_4540);
xor U9820 (N_9820,N_5598,N_5891);
nand U9821 (N_9821,N_6353,N_7787);
and U9822 (N_9822,N_6548,N_5370);
xnor U9823 (N_9823,N_6298,N_7613);
or U9824 (N_9824,N_5832,N_7991);
or U9825 (N_9825,N_5162,N_5400);
nor U9826 (N_9826,N_7986,N_7296);
and U9827 (N_9827,N_7652,N_7451);
nor U9828 (N_9828,N_6537,N_6478);
and U9829 (N_9829,N_6185,N_7163);
nor U9830 (N_9830,N_4994,N_4679);
or U9831 (N_9831,N_7734,N_7307);
nor U9832 (N_9832,N_7072,N_4533);
nor U9833 (N_9833,N_6147,N_4702);
xnor U9834 (N_9834,N_7326,N_4556);
xnor U9835 (N_9835,N_7955,N_6373);
xor U9836 (N_9836,N_7254,N_5707);
and U9837 (N_9837,N_6511,N_5302);
nand U9838 (N_9838,N_5577,N_5660);
nor U9839 (N_9839,N_5653,N_5562);
nand U9840 (N_9840,N_5533,N_5274);
nor U9841 (N_9841,N_6999,N_7452);
nand U9842 (N_9842,N_5096,N_7349);
or U9843 (N_9843,N_5413,N_4598);
xnor U9844 (N_9844,N_7570,N_7628);
or U9845 (N_9845,N_4371,N_7801);
xnor U9846 (N_9846,N_4237,N_4808);
nand U9847 (N_9847,N_7323,N_5721);
and U9848 (N_9848,N_4705,N_4725);
nor U9849 (N_9849,N_7237,N_6551);
or U9850 (N_9850,N_5836,N_7545);
nor U9851 (N_9851,N_6247,N_5762);
nand U9852 (N_9852,N_5953,N_5426);
xnor U9853 (N_9853,N_7930,N_4519);
or U9854 (N_9854,N_4982,N_5838);
and U9855 (N_9855,N_6588,N_5207);
and U9856 (N_9856,N_5910,N_6772);
and U9857 (N_9857,N_7234,N_5100);
nor U9858 (N_9858,N_7488,N_7708);
and U9859 (N_9859,N_6316,N_5265);
or U9860 (N_9860,N_4786,N_6176);
xor U9861 (N_9861,N_4960,N_4007);
nor U9862 (N_9862,N_5259,N_4482);
nand U9863 (N_9863,N_6369,N_6877);
xnor U9864 (N_9864,N_7020,N_5485);
xor U9865 (N_9865,N_6804,N_4028);
xnor U9866 (N_9866,N_4297,N_5615);
nand U9867 (N_9867,N_6392,N_4223);
nor U9868 (N_9868,N_7399,N_4873);
and U9869 (N_9869,N_6244,N_5705);
xnor U9870 (N_9870,N_4572,N_6889);
and U9871 (N_9871,N_7759,N_7940);
and U9872 (N_9872,N_6128,N_6168);
or U9873 (N_9873,N_7336,N_4269);
or U9874 (N_9874,N_5022,N_4618);
xnor U9875 (N_9875,N_4267,N_6675);
or U9876 (N_9876,N_4837,N_5167);
nand U9877 (N_9877,N_6324,N_6910);
or U9878 (N_9878,N_4189,N_5977);
or U9879 (N_9879,N_4413,N_7726);
nor U9880 (N_9880,N_5120,N_4857);
xor U9881 (N_9881,N_7767,N_7038);
nor U9882 (N_9882,N_7142,N_6882);
nor U9883 (N_9883,N_6655,N_7506);
nand U9884 (N_9884,N_6345,N_7694);
and U9885 (N_9885,N_4505,N_7332);
or U9886 (N_9886,N_7733,N_5178);
nand U9887 (N_9887,N_5258,N_5290);
nor U9888 (N_9888,N_4186,N_6344);
or U9889 (N_9889,N_4182,N_7482);
or U9890 (N_9890,N_4438,N_6770);
or U9891 (N_9891,N_5130,N_4690);
nor U9892 (N_9892,N_5573,N_7741);
and U9893 (N_9893,N_4096,N_7104);
or U9894 (N_9894,N_4484,N_6727);
xnor U9895 (N_9895,N_7378,N_6735);
xor U9896 (N_9896,N_5549,N_6499);
or U9897 (N_9897,N_5017,N_5630);
nor U9898 (N_9898,N_5934,N_5633);
nand U9899 (N_9899,N_5383,N_4713);
xnor U9900 (N_9900,N_5467,N_5006);
or U9901 (N_9901,N_5591,N_5638);
xnor U9902 (N_9902,N_7241,N_5878);
or U9903 (N_9903,N_7407,N_5552);
and U9904 (N_9904,N_4086,N_7716);
or U9905 (N_9905,N_7720,N_6825);
and U9906 (N_9906,N_4444,N_5510);
xnor U9907 (N_9907,N_6568,N_7713);
nor U9908 (N_9908,N_6593,N_6894);
and U9909 (N_9909,N_6740,N_5318);
and U9910 (N_9910,N_4574,N_6404);
xnor U9911 (N_9911,N_7731,N_4385);
nor U9912 (N_9912,N_4764,N_4354);
nor U9913 (N_9913,N_4350,N_4151);
nand U9914 (N_9914,N_7289,N_5023);
and U9915 (N_9915,N_7309,N_7277);
nor U9916 (N_9916,N_5321,N_7208);
nor U9917 (N_9917,N_7999,N_5251);
or U9918 (N_9918,N_6790,N_6976);
and U9919 (N_9919,N_6873,N_7873);
xnor U9920 (N_9920,N_4746,N_5233);
xor U9921 (N_9921,N_4006,N_5739);
xnor U9922 (N_9922,N_7710,N_6487);
nand U9923 (N_9923,N_4673,N_7173);
nand U9924 (N_9924,N_5973,N_4278);
nand U9925 (N_9925,N_4016,N_6856);
and U9926 (N_9926,N_4193,N_5928);
or U9927 (N_9927,N_4912,N_6208);
or U9928 (N_9928,N_7445,N_6795);
and U9929 (N_9929,N_5465,N_7666);
xnor U9930 (N_9930,N_6434,N_5954);
nand U9931 (N_9931,N_6925,N_4586);
xnor U9932 (N_9932,N_4461,N_6997);
or U9933 (N_9933,N_5316,N_6574);
nor U9934 (N_9934,N_5628,N_6719);
or U9935 (N_9935,N_6667,N_7604);
or U9936 (N_9936,N_5242,N_7555);
nor U9937 (N_9937,N_5559,N_5693);
nand U9938 (N_9938,N_6468,N_6500);
and U9939 (N_9939,N_6067,N_5741);
xnor U9940 (N_9940,N_6348,N_4639);
nor U9941 (N_9941,N_7913,N_5677);
and U9942 (N_9942,N_7447,N_6939);
nand U9943 (N_9943,N_7816,N_6872);
and U9944 (N_9944,N_7044,N_5072);
nand U9945 (N_9945,N_6438,N_4165);
and U9946 (N_9946,N_5240,N_4195);
or U9947 (N_9947,N_5411,N_6426);
nand U9948 (N_9948,N_4969,N_6275);
and U9949 (N_9949,N_7507,N_7039);
or U9950 (N_9950,N_7678,N_6901);
and U9951 (N_9951,N_6878,N_5867);
or U9952 (N_9952,N_6563,N_6379);
or U9953 (N_9953,N_4547,N_5781);
and U9954 (N_9954,N_6283,N_4432);
xor U9955 (N_9955,N_7607,N_7419);
xnor U9956 (N_9956,N_6652,N_5761);
and U9957 (N_9957,N_5988,N_5532);
nor U9958 (N_9958,N_5818,N_5986);
or U9959 (N_9959,N_5937,N_4296);
xor U9960 (N_9960,N_5343,N_7538);
xnor U9961 (N_9961,N_7471,N_7813);
and U9962 (N_9962,N_4594,N_5111);
or U9963 (N_9963,N_4089,N_7672);
or U9964 (N_9964,N_5229,N_4231);
or U9965 (N_9965,N_6909,N_5389);
nor U9966 (N_9966,N_6004,N_4318);
or U9967 (N_9967,N_7533,N_5209);
or U9968 (N_9968,N_4666,N_5649);
or U9969 (N_9969,N_6398,N_6342);
xnor U9970 (N_9970,N_5232,N_7566);
and U9971 (N_9971,N_6592,N_4626);
or U9972 (N_9972,N_6131,N_7448);
xor U9973 (N_9973,N_4972,N_6864);
and U9974 (N_9974,N_7959,N_7291);
nor U9975 (N_9975,N_5723,N_6063);
and U9976 (N_9976,N_6060,N_5599);
or U9977 (N_9977,N_5848,N_7878);
xor U9978 (N_9978,N_6492,N_4374);
or U9979 (N_9979,N_4111,N_7174);
nand U9980 (N_9980,N_7032,N_5280);
or U9981 (N_9981,N_5991,N_7117);
nor U9982 (N_9982,N_5110,N_5840);
nand U9983 (N_9983,N_5606,N_4801);
xnor U9984 (N_9984,N_7433,N_7537);
nor U9985 (N_9985,N_7762,N_5871);
xor U9986 (N_9986,N_5952,N_7071);
nor U9987 (N_9987,N_6263,N_4405);
and U9988 (N_9988,N_4880,N_7563);
and U9989 (N_9989,N_5433,N_7240);
and U9990 (N_9990,N_7493,N_7777);
or U9991 (N_9991,N_6239,N_7870);
nor U9992 (N_9992,N_4993,N_5983);
or U9993 (N_9993,N_6186,N_5978);
and U9994 (N_9994,N_7276,N_5915);
nor U9995 (N_9995,N_5706,N_4749);
or U9996 (N_9996,N_4733,N_5320);
nand U9997 (N_9997,N_6911,N_4699);
nand U9998 (N_9998,N_6043,N_5479);
nor U9999 (N_9999,N_7464,N_4205);
nand U10000 (N_10000,N_5486,N_6646);
nand U10001 (N_10001,N_6987,N_4335);
or U10002 (N_10002,N_7332,N_7934);
nor U10003 (N_10003,N_7428,N_7037);
or U10004 (N_10004,N_7961,N_5807);
nor U10005 (N_10005,N_5037,N_7307);
and U10006 (N_10006,N_6130,N_5188);
xor U10007 (N_10007,N_4447,N_7551);
nand U10008 (N_10008,N_6035,N_6699);
nand U10009 (N_10009,N_4470,N_5641);
nor U10010 (N_10010,N_5593,N_5942);
xor U10011 (N_10011,N_7288,N_6346);
and U10012 (N_10012,N_5451,N_6900);
xor U10013 (N_10013,N_7352,N_5568);
or U10014 (N_10014,N_5013,N_5639);
xnor U10015 (N_10015,N_4709,N_4105);
xor U10016 (N_10016,N_7510,N_7404);
nand U10017 (N_10017,N_5475,N_7895);
xor U10018 (N_10018,N_5875,N_5619);
nand U10019 (N_10019,N_4805,N_6042);
nand U10020 (N_10020,N_4034,N_5929);
or U10021 (N_10021,N_4009,N_6079);
and U10022 (N_10022,N_5756,N_4355);
xnor U10023 (N_10023,N_6446,N_7768);
and U10024 (N_10024,N_6785,N_5315);
or U10025 (N_10025,N_4616,N_4120);
nor U10026 (N_10026,N_4314,N_7345);
xor U10027 (N_10027,N_6581,N_6691);
and U10028 (N_10028,N_6700,N_7272);
xnor U10029 (N_10029,N_6554,N_4006);
and U10030 (N_10030,N_4967,N_7630);
and U10031 (N_10031,N_4246,N_4429);
nor U10032 (N_10032,N_5201,N_4025);
xnor U10033 (N_10033,N_7876,N_5867);
or U10034 (N_10034,N_5371,N_4854);
nand U10035 (N_10035,N_7347,N_4134);
or U10036 (N_10036,N_7978,N_6837);
nand U10037 (N_10037,N_7315,N_5471);
and U10038 (N_10038,N_5736,N_5710);
or U10039 (N_10039,N_5256,N_4905);
nand U10040 (N_10040,N_5942,N_5805);
and U10041 (N_10041,N_4491,N_5717);
nor U10042 (N_10042,N_5835,N_5432);
xnor U10043 (N_10043,N_4416,N_6415);
nor U10044 (N_10044,N_7634,N_5095);
nand U10045 (N_10045,N_5541,N_4697);
and U10046 (N_10046,N_6370,N_4411);
or U10047 (N_10047,N_7124,N_4740);
xor U10048 (N_10048,N_6504,N_5023);
xor U10049 (N_10049,N_5430,N_4944);
or U10050 (N_10050,N_7220,N_5038);
or U10051 (N_10051,N_5802,N_4957);
nand U10052 (N_10052,N_7946,N_7396);
nand U10053 (N_10053,N_6054,N_7382);
nor U10054 (N_10054,N_5801,N_5475);
nor U10055 (N_10055,N_6517,N_6220);
or U10056 (N_10056,N_4883,N_4648);
nand U10057 (N_10057,N_6662,N_4484);
and U10058 (N_10058,N_7302,N_4091);
nand U10059 (N_10059,N_4142,N_4092);
nand U10060 (N_10060,N_6414,N_5047);
and U10061 (N_10061,N_4318,N_6825);
or U10062 (N_10062,N_5009,N_6808);
or U10063 (N_10063,N_7711,N_4868);
xor U10064 (N_10064,N_4467,N_7065);
and U10065 (N_10065,N_4922,N_5779);
or U10066 (N_10066,N_4782,N_4164);
nand U10067 (N_10067,N_4745,N_7262);
xnor U10068 (N_10068,N_6141,N_7247);
nand U10069 (N_10069,N_5045,N_5318);
or U10070 (N_10070,N_4124,N_5111);
or U10071 (N_10071,N_7141,N_5550);
and U10072 (N_10072,N_5443,N_5892);
nor U10073 (N_10073,N_5487,N_6108);
nand U10074 (N_10074,N_7439,N_7444);
xnor U10075 (N_10075,N_7488,N_7258);
or U10076 (N_10076,N_6678,N_5547);
xnor U10077 (N_10077,N_7971,N_6710);
and U10078 (N_10078,N_7837,N_7116);
nand U10079 (N_10079,N_7093,N_5609);
or U10080 (N_10080,N_7735,N_5273);
nand U10081 (N_10081,N_6294,N_4620);
or U10082 (N_10082,N_6210,N_7917);
xor U10083 (N_10083,N_5316,N_7924);
nand U10084 (N_10084,N_4084,N_7449);
xnor U10085 (N_10085,N_6906,N_7304);
or U10086 (N_10086,N_4748,N_7950);
xor U10087 (N_10087,N_6252,N_4526);
and U10088 (N_10088,N_7934,N_7732);
nand U10089 (N_10089,N_7638,N_7682);
nand U10090 (N_10090,N_4267,N_6041);
or U10091 (N_10091,N_4609,N_6983);
nand U10092 (N_10092,N_4445,N_6346);
or U10093 (N_10093,N_4952,N_5843);
nor U10094 (N_10094,N_4816,N_6701);
nor U10095 (N_10095,N_7048,N_7181);
and U10096 (N_10096,N_7452,N_4522);
and U10097 (N_10097,N_5781,N_6959);
nor U10098 (N_10098,N_5840,N_5561);
and U10099 (N_10099,N_6045,N_7959);
nand U10100 (N_10100,N_5605,N_6226);
and U10101 (N_10101,N_6106,N_5086);
or U10102 (N_10102,N_4702,N_6780);
nand U10103 (N_10103,N_7702,N_4749);
nor U10104 (N_10104,N_4762,N_6792);
or U10105 (N_10105,N_6396,N_6314);
nand U10106 (N_10106,N_6737,N_7833);
xor U10107 (N_10107,N_5053,N_7651);
xnor U10108 (N_10108,N_5984,N_5392);
and U10109 (N_10109,N_7353,N_6304);
xnor U10110 (N_10110,N_4964,N_4298);
and U10111 (N_10111,N_6801,N_7107);
nor U10112 (N_10112,N_7757,N_5540);
and U10113 (N_10113,N_6292,N_7713);
and U10114 (N_10114,N_6385,N_5925);
xor U10115 (N_10115,N_6276,N_5973);
nand U10116 (N_10116,N_7138,N_6022);
xnor U10117 (N_10117,N_6750,N_4120);
xnor U10118 (N_10118,N_6127,N_6049);
xnor U10119 (N_10119,N_7658,N_7212);
and U10120 (N_10120,N_4066,N_6108);
nor U10121 (N_10121,N_4104,N_5663);
nor U10122 (N_10122,N_4345,N_7771);
and U10123 (N_10123,N_6095,N_4967);
nand U10124 (N_10124,N_4024,N_6478);
and U10125 (N_10125,N_5147,N_7207);
nand U10126 (N_10126,N_7664,N_6934);
nor U10127 (N_10127,N_7723,N_5875);
nor U10128 (N_10128,N_5500,N_6295);
or U10129 (N_10129,N_6469,N_6997);
and U10130 (N_10130,N_5907,N_6459);
nor U10131 (N_10131,N_5628,N_4688);
xor U10132 (N_10132,N_7312,N_4920);
nand U10133 (N_10133,N_6585,N_5406);
and U10134 (N_10134,N_5399,N_7630);
or U10135 (N_10135,N_4613,N_7811);
or U10136 (N_10136,N_6426,N_5110);
xnor U10137 (N_10137,N_4023,N_5344);
and U10138 (N_10138,N_4373,N_5999);
xnor U10139 (N_10139,N_7364,N_6010);
xnor U10140 (N_10140,N_6313,N_6682);
nor U10141 (N_10141,N_6510,N_5798);
and U10142 (N_10142,N_5854,N_6348);
xnor U10143 (N_10143,N_4421,N_4340);
xnor U10144 (N_10144,N_4391,N_5826);
xnor U10145 (N_10145,N_5282,N_4597);
nand U10146 (N_10146,N_7635,N_4798);
xnor U10147 (N_10147,N_4459,N_4371);
xnor U10148 (N_10148,N_7244,N_5104);
or U10149 (N_10149,N_4565,N_7779);
nor U10150 (N_10150,N_4926,N_7368);
and U10151 (N_10151,N_7937,N_5195);
or U10152 (N_10152,N_4728,N_6487);
nor U10153 (N_10153,N_4057,N_5702);
xnor U10154 (N_10154,N_6647,N_7994);
or U10155 (N_10155,N_5108,N_5456);
nor U10156 (N_10156,N_5077,N_4725);
nand U10157 (N_10157,N_5890,N_6861);
nand U10158 (N_10158,N_6312,N_4530);
and U10159 (N_10159,N_5135,N_7111);
nor U10160 (N_10160,N_7533,N_4434);
or U10161 (N_10161,N_4824,N_7699);
xor U10162 (N_10162,N_7776,N_5178);
and U10163 (N_10163,N_5665,N_4305);
or U10164 (N_10164,N_6665,N_4247);
nor U10165 (N_10165,N_5243,N_7043);
nor U10166 (N_10166,N_7908,N_4650);
or U10167 (N_10167,N_7676,N_6018);
nand U10168 (N_10168,N_7254,N_7533);
nand U10169 (N_10169,N_4352,N_5557);
nor U10170 (N_10170,N_6562,N_7889);
nor U10171 (N_10171,N_6892,N_5665);
or U10172 (N_10172,N_4427,N_4588);
nand U10173 (N_10173,N_7763,N_4805);
or U10174 (N_10174,N_5809,N_6354);
xnor U10175 (N_10175,N_6618,N_4505);
nor U10176 (N_10176,N_6978,N_5827);
nand U10177 (N_10177,N_5071,N_7911);
and U10178 (N_10178,N_5046,N_5168);
xnor U10179 (N_10179,N_4157,N_6754);
or U10180 (N_10180,N_5238,N_7284);
nor U10181 (N_10181,N_4821,N_5042);
nor U10182 (N_10182,N_6943,N_5257);
and U10183 (N_10183,N_5649,N_7635);
xnor U10184 (N_10184,N_5935,N_7166);
nand U10185 (N_10185,N_5739,N_4032);
nand U10186 (N_10186,N_6582,N_6437);
or U10187 (N_10187,N_6791,N_4721);
or U10188 (N_10188,N_5818,N_7730);
nand U10189 (N_10189,N_6806,N_4923);
nor U10190 (N_10190,N_6048,N_5729);
xor U10191 (N_10191,N_5604,N_4088);
and U10192 (N_10192,N_7534,N_5979);
nand U10193 (N_10193,N_7311,N_6934);
and U10194 (N_10194,N_7231,N_7941);
nand U10195 (N_10195,N_7945,N_7469);
nand U10196 (N_10196,N_6024,N_6115);
xor U10197 (N_10197,N_4241,N_5906);
nand U10198 (N_10198,N_5236,N_7375);
xor U10199 (N_10199,N_4338,N_4579);
or U10200 (N_10200,N_4253,N_4596);
or U10201 (N_10201,N_4045,N_6708);
xnor U10202 (N_10202,N_4418,N_6093);
and U10203 (N_10203,N_7901,N_5748);
nand U10204 (N_10204,N_4529,N_4500);
and U10205 (N_10205,N_4286,N_4246);
or U10206 (N_10206,N_7328,N_7806);
nor U10207 (N_10207,N_7426,N_4159);
xor U10208 (N_10208,N_6244,N_5935);
nand U10209 (N_10209,N_4971,N_5495);
nor U10210 (N_10210,N_4569,N_6004);
nand U10211 (N_10211,N_5594,N_6491);
and U10212 (N_10212,N_7967,N_6969);
and U10213 (N_10213,N_6056,N_6338);
or U10214 (N_10214,N_5007,N_5486);
nand U10215 (N_10215,N_7205,N_6183);
or U10216 (N_10216,N_4681,N_5003);
nor U10217 (N_10217,N_4719,N_6189);
or U10218 (N_10218,N_4222,N_4008);
and U10219 (N_10219,N_5204,N_5987);
nor U10220 (N_10220,N_7311,N_4202);
nand U10221 (N_10221,N_7903,N_7691);
nor U10222 (N_10222,N_7494,N_4224);
or U10223 (N_10223,N_7072,N_6527);
nor U10224 (N_10224,N_6470,N_4874);
or U10225 (N_10225,N_5531,N_5542);
nor U10226 (N_10226,N_6921,N_6963);
or U10227 (N_10227,N_4584,N_7580);
nand U10228 (N_10228,N_5612,N_5720);
nand U10229 (N_10229,N_6751,N_7708);
xnor U10230 (N_10230,N_7437,N_7327);
nand U10231 (N_10231,N_6602,N_7879);
and U10232 (N_10232,N_4057,N_7439);
and U10233 (N_10233,N_7072,N_5691);
nor U10234 (N_10234,N_5701,N_4556);
and U10235 (N_10235,N_5974,N_5830);
xnor U10236 (N_10236,N_7963,N_5258);
or U10237 (N_10237,N_6046,N_4162);
or U10238 (N_10238,N_7411,N_5450);
and U10239 (N_10239,N_5112,N_6206);
nand U10240 (N_10240,N_4083,N_5772);
nor U10241 (N_10241,N_7298,N_7134);
or U10242 (N_10242,N_5853,N_4980);
or U10243 (N_10243,N_4892,N_4764);
or U10244 (N_10244,N_4304,N_4393);
nand U10245 (N_10245,N_5625,N_4498);
or U10246 (N_10246,N_6835,N_6160);
or U10247 (N_10247,N_6521,N_5107);
and U10248 (N_10248,N_7243,N_4101);
and U10249 (N_10249,N_5178,N_4963);
and U10250 (N_10250,N_5687,N_4474);
and U10251 (N_10251,N_4057,N_7162);
nand U10252 (N_10252,N_4482,N_6522);
nand U10253 (N_10253,N_5393,N_6254);
nor U10254 (N_10254,N_6726,N_6512);
and U10255 (N_10255,N_5997,N_5759);
or U10256 (N_10256,N_5508,N_5425);
xor U10257 (N_10257,N_5889,N_4341);
or U10258 (N_10258,N_5453,N_5866);
nor U10259 (N_10259,N_4787,N_4590);
nor U10260 (N_10260,N_4750,N_6413);
nand U10261 (N_10261,N_7752,N_6821);
nor U10262 (N_10262,N_5440,N_4532);
xor U10263 (N_10263,N_4658,N_4441);
nand U10264 (N_10264,N_5021,N_4104);
and U10265 (N_10265,N_7555,N_4867);
nand U10266 (N_10266,N_5794,N_5421);
or U10267 (N_10267,N_6871,N_4709);
nor U10268 (N_10268,N_4957,N_7276);
or U10269 (N_10269,N_4022,N_6001);
and U10270 (N_10270,N_5535,N_5918);
nor U10271 (N_10271,N_6458,N_7782);
nand U10272 (N_10272,N_4142,N_7241);
and U10273 (N_10273,N_4464,N_6992);
xor U10274 (N_10274,N_4233,N_4730);
or U10275 (N_10275,N_5216,N_5407);
or U10276 (N_10276,N_7532,N_4446);
xnor U10277 (N_10277,N_7899,N_4374);
and U10278 (N_10278,N_6451,N_6728);
nor U10279 (N_10279,N_5060,N_7465);
nor U10280 (N_10280,N_7700,N_6957);
and U10281 (N_10281,N_6665,N_6087);
nor U10282 (N_10282,N_6557,N_4146);
and U10283 (N_10283,N_4782,N_6545);
nor U10284 (N_10284,N_5454,N_5273);
nand U10285 (N_10285,N_4180,N_6930);
nand U10286 (N_10286,N_6146,N_5146);
or U10287 (N_10287,N_7980,N_6085);
xor U10288 (N_10288,N_4997,N_4731);
nor U10289 (N_10289,N_4795,N_5148);
nor U10290 (N_10290,N_6409,N_5718);
nand U10291 (N_10291,N_6555,N_7609);
and U10292 (N_10292,N_5043,N_4110);
nor U10293 (N_10293,N_5748,N_6096);
nand U10294 (N_10294,N_7061,N_4968);
or U10295 (N_10295,N_6827,N_6578);
and U10296 (N_10296,N_6568,N_7126);
xnor U10297 (N_10297,N_6925,N_7181);
or U10298 (N_10298,N_5266,N_4549);
and U10299 (N_10299,N_6796,N_5835);
or U10300 (N_10300,N_6151,N_7568);
xnor U10301 (N_10301,N_5865,N_4370);
nor U10302 (N_10302,N_4933,N_5373);
and U10303 (N_10303,N_7116,N_6983);
nand U10304 (N_10304,N_5765,N_6322);
nor U10305 (N_10305,N_5418,N_5813);
and U10306 (N_10306,N_6638,N_6296);
nand U10307 (N_10307,N_4631,N_7284);
xor U10308 (N_10308,N_4661,N_5424);
nand U10309 (N_10309,N_4872,N_4976);
nand U10310 (N_10310,N_4470,N_4059);
xnor U10311 (N_10311,N_4425,N_5720);
nor U10312 (N_10312,N_7418,N_7277);
and U10313 (N_10313,N_6337,N_5149);
xor U10314 (N_10314,N_7607,N_6460);
or U10315 (N_10315,N_6953,N_4417);
nor U10316 (N_10316,N_5740,N_5632);
xnor U10317 (N_10317,N_4580,N_4623);
and U10318 (N_10318,N_5885,N_6026);
xnor U10319 (N_10319,N_7543,N_4291);
nor U10320 (N_10320,N_7632,N_6621);
nand U10321 (N_10321,N_4149,N_6073);
xnor U10322 (N_10322,N_5841,N_4323);
and U10323 (N_10323,N_4616,N_5826);
and U10324 (N_10324,N_6637,N_5610);
xnor U10325 (N_10325,N_7062,N_6859);
xnor U10326 (N_10326,N_4647,N_5426);
nor U10327 (N_10327,N_5343,N_5404);
xnor U10328 (N_10328,N_7850,N_5554);
nor U10329 (N_10329,N_7257,N_7915);
and U10330 (N_10330,N_7380,N_7786);
nand U10331 (N_10331,N_4232,N_6254);
nand U10332 (N_10332,N_6132,N_5234);
and U10333 (N_10333,N_5578,N_5594);
and U10334 (N_10334,N_6029,N_5472);
and U10335 (N_10335,N_6769,N_5575);
or U10336 (N_10336,N_6314,N_6531);
nand U10337 (N_10337,N_4188,N_6829);
xnor U10338 (N_10338,N_6227,N_6264);
xnor U10339 (N_10339,N_4159,N_5406);
and U10340 (N_10340,N_4983,N_7764);
or U10341 (N_10341,N_4996,N_7364);
nor U10342 (N_10342,N_5425,N_4084);
xnor U10343 (N_10343,N_7149,N_5231);
and U10344 (N_10344,N_5599,N_4426);
or U10345 (N_10345,N_7339,N_4156);
and U10346 (N_10346,N_6728,N_7441);
and U10347 (N_10347,N_6555,N_6592);
xnor U10348 (N_10348,N_4741,N_4765);
nand U10349 (N_10349,N_5432,N_4545);
or U10350 (N_10350,N_5205,N_7858);
xnor U10351 (N_10351,N_5146,N_7532);
nor U10352 (N_10352,N_6624,N_4173);
and U10353 (N_10353,N_6506,N_6416);
and U10354 (N_10354,N_7278,N_5169);
nor U10355 (N_10355,N_5006,N_7482);
nor U10356 (N_10356,N_7626,N_5345);
and U10357 (N_10357,N_5543,N_6266);
nand U10358 (N_10358,N_5518,N_7550);
or U10359 (N_10359,N_5184,N_7455);
or U10360 (N_10360,N_7360,N_4531);
nand U10361 (N_10361,N_5946,N_6939);
nand U10362 (N_10362,N_4119,N_5504);
or U10363 (N_10363,N_7193,N_4203);
or U10364 (N_10364,N_7120,N_4310);
nor U10365 (N_10365,N_7530,N_5999);
nand U10366 (N_10366,N_6984,N_7016);
or U10367 (N_10367,N_7813,N_6061);
nand U10368 (N_10368,N_5239,N_7364);
and U10369 (N_10369,N_7710,N_4935);
xnor U10370 (N_10370,N_4218,N_5901);
nand U10371 (N_10371,N_6924,N_7087);
xnor U10372 (N_10372,N_6142,N_4364);
nand U10373 (N_10373,N_5694,N_5514);
nand U10374 (N_10374,N_6528,N_6167);
nand U10375 (N_10375,N_7232,N_5866);
nand U10376 (N_10376,N_6382,N_7730);
xnor U10377 (N_10377,N_4954,N_7256);
and U10378 (N_10378,N_4115,N_5356);
nor U10379 (N_10379,N_7104,N_4515);
or U10380 (N_10380,N_4297,N_7782);
or U10381 (N_10381,N_6957,N_5932);
xor U10382 (N_10382,N_7364,N_5335);
xor U10383 (N_10383,N_7787,N_5809);
nand U10384 (N_10384,N_5572,N_7797);
nor U10385 (N_10385,N_5905,N_7328);
and U10386 (N_10386,N_7402,N_4320);
nor U10387 (N_10387,N_6907,N_7654);
xor U10388 (N_10388,N_6774,N_5603);
or U10389 (N_10389,N_6449,N_4290);
xor U10390 (N_10390,N_5251,N_7633);
xnor U10391 (N_10391,N_5211,N_4853);
and U10392 (N_10392,N_5691,N_5913);
nand U10393 (N_10393,N_7201,N_6959);
nor U10394 (N_10394,N_5041,N_7887);
nand U10395 (N_10395,N_6963,N_4401);
xnor U10396 (N_10396,N_4194,N_4017);
nand U10397 (N_10397,N_4061,N_6338);
nor U10398 (N_10398,N_5468,N_6605);
and U10399 (N_10399,N_6679,N_4740);
or U10400 (N_10400,N_6342,N_6338);
and U10401 (N_10401,N_5976,N_7469);
nand U10402 (N_10402,N_5911,N_6197);
or U10403 (N_10403,N_7510,N_5612);
nor U10404 (N_10404,N_6215,N_5020);
nand U10405 (N_10405,N_5520,N_7835);
or U10406 (N_10406,N_6361,N_5892);
and U10407 (N_10407,N_4461,N_7317);
nand U10408 (N_10408,N_6750,N_5749);
and U10409 (N_10409,N_6418,N_6853);
nor U10410 (N_10410,N_4997,N_7823);
and U10411 (N_10411,N_4583,N_4679);
or U10412 (N_10412,N_7669,N_7491);
nor U10413 (N_10413,N_4659,N_4685);
or U10414 (N_10414,N_5810,N_6062);
nor U10415 (N_10415,N_4458,N_6057);
nor U10416 (N_10416,N_6433,N_7656);
nor U10417 (N_10417,N_5984,N_5326);
nand U10418 (N_10418,N_4901,N_7844);
and U10419 (N_10419,N_7117,N_5875);
or U10420 (N_10420,N_7664,N_4492);
nor U10421 (N_10421,N_5739,N_6341);
or U10422 (N_10422,N_7609,N_4582);
xor U10423 (N_10423,N_4572,N_4807);
xor U10424 (N_10424,N_4512,N_6902);
or U10425 (N_10425,N_7883,N_7707);
and U10426 (N_10426,N_4161,N_4480);
xor U10427 (N_10427,N_4297,N_7928);
nor U10428 (N_10428,N_4524,N_4871);
or U10429 (N_10429,N_7492,N_7053);
nand U10430 (N_10430,N_4010,N_5258);
nand U10431 (N_10431,N_7980,N_7006);
xnor U10432 (N_10432,N_4887,N_6226);
or U10433 (N_10433,N_4560,N_5981);
or U10434 (N_10434,N_6505,N_4016);
and U10435 (N_10435,N_5652,N_5961);
nor U10436 (N_10436,N_7695,N_4149);
nand U10437 (N_10437,N_4040,N_7825);
nand U10438 (N_10438,N_7733,N_5230);
and U10439 (N_10439,N_7901,N_6595);
or U10440 (N_10440,N_4603,N_7377);
xnor U10441 (N_10441,N_4127,N_4190);
xnor U10442 (N_10442,N_4680,N_5696);
and U10443 (N_10443,N_7854,N_4271);
or U10444 (N_10444,N_7383,N_4302);
and U10445 (N_10445,N_7637,N_6540);
or U10446 (N_10446,N_5394,N_5035);
xor U10447 (N_10447,N_7571,N_5347);
xor U10448 (N_10448,N_5460,N_5547);
or U10449 (N_10449,N_7223,N_4818);
or U10450 (N_10450,N_4895,N_6036);
or U10451 (N_10451,N_6212,N_6207);
nand U10452 (N_10452,N_6659,N_7019);
nand U10453 (N_10453,N_4351,N_4390);
nand U10454 (N_10454,N_7925,N_5428);
xor U10455 (N_10455,N_4584,N_5024);
xnor U10456 (N_10456,N_5868,N_6874);
or U10457 (N_10457,N_7753,N_5930);
nor U10458 (N_10458,N_4599,N_7232);
nor U10459 (N_10459,N_6469,N_6652);
or U10460 (N_10460,N_4153,N_4718);
or U10461 (N_10461,N_7165,N_7751);
or U10462 (N_10462,N_4716,N_7564);
or U10463 (N_10463,N_7626,N_7589);
and U10464 (N_10464,N_5469,N_7125);
nor U10465 (N_10465,N_4407,N_5444);
or U10466 (N_10466,N_4210,N_4816);
nor U10467 (N_10467,N_7202,N_7886);
and U10468 (N_10468,N_4831,N_4259);
and U10469 (N_10469,N_7474,N_4736);
nand U10470 (N_10470,N_5366,N_4230);
or U10471 (N_10471,N_5104,N_6712);
xor U10472 (N_10472,N_7242,N_7687);
nand U10473 (N_10473,N_6467,N_5408);
or U10474 (N_10474,N_6057,N_6920);
nand U10475 (N_10475,N_7242,N_4576);
nand U10476 (N_10476,N_7115,N_4322);
and U10477 (N_10477,N_7938,N_4063);
or U10478 (N_10478,N_4501,N_5703);
nand U10479 (N_10479,N_6928,N_6694);
or U10480 (N_10480,N_6418,N_7846);
xnor U10481 (N_10481,N_6813,N_5631);
nor U10482 (N_10482,N_4021,N_4299);
and U10483 (N_10483,N_6883,N_4310);
and U10484 (N_10484,N_4585,N_4258);
or U10485 (N_10485,N_5092,N_6649);
or U10486 (N_10486,N_5906,N_6198);
and U10487 (N_10487,N_7450,N_4927);
xor U10488 (N_10488,N_4792,N_6133);
xnor U10489 (N_10489,N_6021,N_4298);
or U10490 (N_10490,N_4266,N_6685);
nand U10491 (N_10491,N_7069,N_6768);
xor U10492 (N_10492,N_4405,N_6314);
nor U10493 (N_10493,N_6931,N_6401);
and U10494 (N_10494,N_4304,N_4649);
and U10495 (N_10495,N_4707,N_7646);
or U10496 (N_10496,N_6191,N_4481);
nand U10497 (N_10497,N_5582,N_5830);
and U10498 (N_10498,N_5414,N_6544);
nand U10499 (N_10499,N_5887,N_7953);
xnor U10500 (N_10500,N_5822,N_6934);
nand U10501 (N_10501,N_4719,N_4152);
and U10502 (N_10502,N_6318,N_6636);
nor U10503 (N_10503,N_7541,N_7015);
and U10504 (N_10504,N_4456,N_5610);
xor U10505 (N_10505,N_4524,N_4938);
nand U10506 (N_10506,N_5766,N_7335);
xnor U10507 (N_10507,N_5138,N_5344);
or U10508 (N_10508,N_4284,N_4540);
and U10509 (N_10509,N_6124,N_4594);
and U10510 (N_10510,N_7908,N_5676);
nor U10511 (N_10511,N_6666,N_5602);
nor U10512 (N_10512,N_5997,N_6543);
nand U10513 (N_10513,N_7974,N_6077);
nand U10514 (N_10514,N_4116,N_6291);
nand U10515 (N_10515,N_5173,N_7562);
or U10516 (N_10516,N_6484,N_6212);
nor U10517 (N_10517,N_7197,N_6658);
xor U10518 (N_10518,N_6990,N_7420);
and U10519 (N_10519,N_6641,N_4775);
nand U10520 (N_10520,N_4033,N_6608);
or U10521 (N_10521,N_5091,N_7440);
xor U10522 (N_10522,N_4198,N_4182);
nor U10523 (N_10523,N_6030,N_4129);
nand U10524 (N_10524,N_4259,N_5334);
nor U10525 (N_10525,N_6227,N_5826);
nand U10526 (N_10526,N_6460,N_5946);
xor U10527 (N_10527,N_6746,N_6271);
and U10528 (N_10528,N_4162,N_7824);
xnor U10529 (N_10529,N_5843,N_5328);
and U10530 (N_10530,N_4569,N_7087);
xor U10531 (N_10531,N_7262,N_6661);
nand U10532 (N_10532,N_7647,N_4181);
xor U10533 (N_10533,N_4847,N_5474);
nor U10534 (N_10534,N_5968,N_6384);
or U10535 (N_10535,N_6968,N_4102);
or U10536 (N_10536,N_6116,N_7490);
xor U10537 (N_10537,N_5184,N_7863);
and U10538 (N_10538,N_7256,N_4795);
or U10539 (N_10539,N_7545,N_4938);
or U10540 (N_10540,N_7660,N_4754);
and U10541 (N_10541,N_7641,N_6855);
or U10542 (N_10542,N_6532,N_4480);
or U10543 (N_10543,N_5810,N_5287);
and U10544 (N_10544,N_6899,N_4868);
or U10545 (N_10545,N_5343,N_4407);
and U10546 (N_10546,N_5379,N_7632);
nand U10547 (N_10547,N_4586,N_7202);
or U10548 (N_10548,N_4639,N_4552);
and U10549 (N_10549,N_5688,N_7365);
and U10550 (N_10550,N_5411,N_4610);
and U10551 (N_10551,N_4603,N_6167);
or U10552 (N_10552,N_7803,N_4777);
and U10553 (N_10553,N_7105,N_4496);
nand U10554 (N_10554,N_4134,N_7466);
nand U10555 (N_10555,N_7766,N_6345);
nor U10556 (N_10556,N_7090,N_7867);
xnor U10557 (N_10557,N_5103,N_6449);
and U10558 (N_10558,N_7514,N_4527);
and U10559 (N_10559,N_7104,N_5910);
and U10560 (N_10560,N_4008,N_7268);
nor U10561 (N_10561,N_7541,N_4755);
nor U10562 (N_10562,N_6752,N_7779);
nand U10563 (N_10563,N_4905,N_5605);
xnor U10564 (N_10564,N_4818,N_6675);
nand U10565 (N_10565,N_5146,N_6197);
and U10566 (N_10566,N_4427,N_5582);
nor U10567 (N_10567,N_5936,N_7330);
nand U10568 (N_10568,N_6316,N_7243);
nor U10569 (N_10569,N_6092,N_7129);
xor U10570 (N_10570,N_6484,N_6972);
nand U10571 (N_10571,N_6391,N_5741);
nand U10572 (N_10572,N_6664,N_7907);
or U10573 (N_10573,N_4285,N_7618);
or U10574 (N_10574,N_6518,N_7662);
and U10575 (N_10575,N_5033,N_4174);
or U10576 (N_10576,N_5605,N_4108);
and U10577 (N_10577,N_6818,N_5894);
nand U10578 (N_10578,N_4081,N_7366);
nand U10579 (N_10579,N_4618,N_6036);
nor U10580 (N_10580,N_4649,N_6193);
nor U10581 (N_10581,N_6723,N_5803);
nand U10582 (N_10582,N_5418,N_6897);
and U10583 (N_10583,N_4347,N_6455);
xor U10584 (N_10584,N_4180,N_5449);
or U10585 (N_10585,N_7131,N_5372);
xnor U10586 (N_10586,N_5654,N_5379);
nor U10587 (N_10587,N_4268,N_5832);
or U10588 (N_10588,N_4515,N_4297);
and U10589 (N_10589,N_4691,N_4630);
nor U10590 (N_10590,N_7928,N_4245);
or U10591 (N_10591,N_7258,N_4948);
and U10592 (N_10592,N_7192,N_4999);
and U10593 (N_10593,N_4848,N_4499);
or U10594 (N_10594,N_4599,N_5117);
nor U10595 (N_10595,N_7337,N_4517);
nand U10596 (N_10596,N_6601,N_7335);
xor U10597 (N_10597,N_7068,N_6914);
and U10598 (N_10598,N_7165,N_7338);
xor U10599 (N_10599,N_7676,N_7817);
xnor U10600 (N_10600,N_7448,N_7184);
nand U10601 (N_10601,N_6755,N_6668);
or U10602 (N_10602,N_6145,N_5970);
nor U10603 (N_10603,N_6111,N_5775);
nor U10604 (N_10604,N_6935,N_5740);
xnor U10605 (N_10605,N_7937,N_5512);
and U10606 (N_10606,N_7650,N_4112);
nand U10607 (N_10607,N_7613,N_7260);
and U10608 (N_10608,N_5147,N_4285);
or U10609 (N_10609,N_4698,N_6048);
nand U10610 (N_10610,N_4336,N_7670);
or U10611 (N_10611,N_4927,N_5848);
xnor U10612 (N_10612,N_7987,N_5902);
nor U10613 (N_10613,N_5185,N_5788);
xnor U10614 (N_10614,N_5657,N_6574);
and U10615 (N_10615,N_7234,N_4386);
xnor U10616 (N_10616,N_4161,N_4846);
and U10617 (N_10617,N_4212,N_6357);
nor U10618 (N_10618,N_5778,N_7975);
and U10619 (N_10619,N_5291,N_7248);
nor U10620 (N_10620,N_7743,N_5998);
and U10621 (N_10621,N_6782,N_6067);
and U10622 (N_10622,N_5668,N_5065);
and U10623 (N_10623,N_6657,N_7785);
or U10624 (N_10624,N_6385,N_4855);
nor U10625 (N_10625,N_7568,N_4442);
and U10626 (N_10626,N_4732,N_7281);
or U10627 (N_10627,N_6311,N_6119);
and U10628 (N_10628,N_7001,N_4894);
and U10629 (N_10629,N_6290,N_6642);
or U10630 (N_10630,N_4834,N_7023);
xor U10631 (N_10631,N_5849,N_4420);
xor U10632 (N_10632,N_4820,N_4169);
nor U10633 (N_10633,N_4886,N_7021);
nor U10634 (N_10634,N_6271,N_5078);
xnor U10635 (N_10635,N_4361,N_5019);
xnor U10636 (N_10636,N_4162,N_7601);
xnor U10637 (N_10637,N_4179,N_4201);
xnor U10638 (N_10638,N_7433,N_7802);
xor U10639 (N_10639,N_5537,N_4877);
and U10640 (N_10640,N_5759,N_5870);
and U10641 (N_10641,N_7346,N_4428);
nor U10642 (N_10642,N_4106,N_7637);
nand U10643 (N_10643,N_7983,N_7708);
or U10644 (N_10644,N_4255,N_6624);
and U10645 (N_10645,N_4760,N_7402);
xnor U10646 (N_10646,N_6704,N_5532);
xor U10647 (N_10647,N_7871,N_5371);
or U10648 (N_10648,N_6200,N_6878);
and U10649 (N_10649,N_4828,N_7172);
xor U10650 (N_10650,N_6074,N_7872);
and U10651 (N_10651,N_4374,N_7321);
xnor U10652 (N_10652,N_4379,N_4138);
xor U10653 (N_10653,N_4688,N_5186);
or U10654 (N_10654,N_7234,N_7121);
and U10655 (N_10655,N_7931,N_6448);
xor U10656 (N_10656,N_5690,N_5600);
xor U10657 (N_10657,N_5139,N_6509);
nand U10658 (N_10658,N_7216,N_4382);
nand U10659 (N_10659,N_6889,N_5826);
nand U10660 (N_10660,N_6355,N_6487);
xnor U10661 (N_10661,N_6405,N_7140);
xnor U10662 (N_10662,N_7117,N_5603);
nor U10663 (N_10663,N_7762,N_6255);
nand U10664 (N_10664,N_5908,N_7104);
xor U10665 (N_10665,N_5560,N_7183);
nand U10666 (N_10666,N_4289,N_5008);
xnor U10667 (N_10667,N_4734,N_7153);
and U10668 (N_10668,N_4661,N_5060);
xor U10669 (N_10669,N_6540,N_5556);
nand U10670 (N_10670,N_7552,N_6173);
nand U10671 (N_10671,N_7637,N_4846);
nor U10672 (N_10672,N_7186,N_7202);
or U10673 (N_10673,N_4180,N_6912);
nor U10674 (N_10674,N_7935,N_6128);
xor U10675 (N_10675,N_4141,N_7533);
xor U10676 (N_10676,N_5837,N_5607);
xnor U10677 (N_10677,N_4242,N_5521);
nand U10678 (N_10678,N_5112,N_7237);
nor U10679 (N_10679,N_7928,N_4572);
and U10680 (N_10680,N_6254,N_4450);
nor U10681 (N_10681,N_6315,N_7554);
or U10682 (N_10682,N_7262,N_6071);
nor U10683 (N_10683,N_4207,N_6744);
nor U10684 (N_10684,N_5785,N_5948);
nor U10685 (N_10685,N_5571,N_7115);
xor U10686 (N_10686,N_6673,N_4434);
or U10687 (N_10687,N_6488,N_5376);
or U10688 (N_10688,N_7233,N_4096);
nand U10689 (N_10689,N_4762,N_7196);
nand U10690 (N_10690,N_7536,N_5100);
nor U10691 (N_10691,N_4368,N_5158);
and U10692 (N_10692,N_4074,N_6945);
and U10693 (N_10693,N_5671,N_4298);
and U10694 (N_10694,N_5474,N_5836);
and U10695 (N_10695,N_6841,N_6312);
xnor U10696 (N_10696,N_4791,N_7549);
and U10697 (N_10697,N_5699,N_4860);
or U10698 (N_10698,N_7755,N_5248);
or U10699 (N_10699,N_4632,N_7543);
xor U10700 (N_10700,N_6633,N_4517);
or U10701 (N_10701,N_5972,N_7886);
or U10702 (N_10702,N_6605,N_7055);
nor U10703 (N_10703,N_5194,N_7095);
and U10704 (N_10704,N_7491,N_7903);
xor U10705 (N_10705,N_7475,N_5607);
or U10706 (N_10706,N_6017,N_7923);
or U10707 (N_10707,N_6752,N_6545);
and U10708 (N_10708,N_4756,N_6057);
nor U10709 (N_10709,N_4168,N_6051);
nor U10710 (N_10710,N_7196,N_7851);
and U10711 (N_10711,N_4883,N_5149);
or U10712 (N_10712,N_5849,N_5852);
and U10713 (N_10713,N_5392,N_6725);
and U10714 (N_10714,N_5248,N_7929);
and U10715 (N_10715,N_4702,N_5214);
xnor U10716 (N_10716,N_4202,N_4364);
or U10717 (N_10717,N_6780,N_5893);
nand U10718 (N_10718,N_5431,N_4620);
and U10719 (N_10719,N_4726,N_7723);
or U10720 (N_10720,N_6297,N_6946);
or U10721 (N_10721,N_4136,N_6083);
or U10722 (N_10722,N_6099,N_4332);
nor U10723 (N_10723,N_4991,N_6969);
or U10724 (N_10724,N_6379,N_7791);
and U10725 (N_10725,N_6876,N_4315);
and U10726 (N_10726,N_6632,N_5087);
nand U10727 (N_10727,N_7530,N_7458);
xor U10728 (N_10728,N_6024,N_4373);
nand U10729 (N_10729,N_6589,N_6234);
xnor U10730 (N_10730,N_4662,N_5231);
nor U10731 (N_10731,N_4688,N_5380);
or U10732 (N_10732,N_7860,N_4183);
nor U10733 (N_10733,N_4040,N_7105);
xnor U10734 (N_10734,N_5966,N_7254);
nand U10735 (N_10735,N_6929,N_4066);
nand U10736 (N_10736,N_5822,N_6034);
nor U10737 (N_10737,N_4435,N_5182);
nor U10738 (N_10738,N_6755,N_7773);
and U10739 (N_10739,N_4130,N_6966);
or U10740 (N_10740,N_4468,N_5379);
or U10741 (N_10741,N_6059,N_6116);
nor U10742 (N_10742,N_5823,N_6062);
nand U10743 (N_10743,N_7710,N_6930);
and U10744 (N_10744,N_6004,N_7795);
or U10745 (N_10745,N_5725,N_6954);
or U10746 (N_10746,N_6229,N_5363);
or U10747 (N_10747,N_7050,N_7087);
nor U10748 (N_10748,N_7878,N_6739);
or U10749 (N_10749,N_7119,N_5574);
nand U10750 (N_10750,N_5709,N_7751);
xor U10751 (N_10751,N_5335,N_5918);
nand U10752 (N_10752,N_4180,N_6654);
or U10753 (N_10753,N_4532,N_5097);
and U10754 (N_10754,N_6060,N_4614);
and U10755 (N_10755,N_7073,N_5717);
nand U10756 (N_10756,N_4360,N_6717);
and U10757 (N_10757,N_7860,N_5731);
nand U10758 (N_10758,N_6135,N_6775);
or U10759 (N_10759,N_5081,N_4122);
xor U10760 (N_10760,N_7504,N_6107);
nand U10761 (N_10761,N_5928,N_5308);
and U10762 (N_10762,N_5328,N_6034);
nand U10763 (N_10763,N_7089,N_6167);
or U10764 (N_10764,N_6533,N_4205);
and U10765 (N_10765,N_5198,N_4747);
nand U10766 (N_10766,N_5340,N_7905);
nand U10767 (N_10767,N_6517,N_4155);
nor U10768 (N_10768,N_4693,N_7336);
nand U10769 (N_10769,N_7597,N_6625);
nand U10770 (N_10770,N_5957,N_5105);
nor U10771 (N_10771,N_7001,N_6967);
and U10772 (N_10772,N_7522,N_7932);
nor U10773 (N_10773,N_4884,N_6902);
nand U10774 (N_10774,N_4953,N_5346);
xnor U10775 (N_10775,N_6787,N_6958);
nand U10776 (N_10776,N_5991,N_4495);
nor U10777 (N_10777,N_4333,N_5448);
xor U10778 (N_10778,N_5824,N_6123);
nor U10779 (N_10779,N_6912,N_4269);
nand U10780 (N_10780,N_6499,N_6338);
nand U10781 (N_10781,N_5268,N_6531);
or U10782 (N_10782,N_5708,N_6146);
xnor U10783 (N_10783,N_7667,N_5316);
or U10784 (N_10784,N_7026,N_5792);
xor U10785 (N_10785,N_7160,N_5205);
and U10786 (N_10786,N_7094,N_6376);
nor U10787 (N_10787,N_4578,N_5152);
xnor U10788 (N_10788,N_5249,N_6514);
or U10789 (N_10789,N_4059,N_5331);
xnor U10790 (N_10790,N_7662,N_6320);
nand U10791 (N_10791,N_5615,N_6838);
or U10792 (N_10792,N_4202,N_4013);
or U10793 (N_10793,N_4532,N_5319);
xnor U10794 (N_10794,N_7844,N_4427);
and U10795 (N_10795,N_5634,N_6900);
nor U10796 (N_10796,N_4418,N_5453);
or U10797 (N_10797,N_6258,N_4108);
and U10798 (N_10798,N_7822,N_5513);
nand U10799 (N_10799,N_7490,N_4399);
xor U10800 (N_10800,N_4041,N_6154);
nor U10801 (N_10801,N_5571,N_6258);
and U10802 (N_10802,N_5622,N_7973);
xor U10803 (N_10803,N_7184,N_5690);
nand U10804 (N_10804,N_7365,N_6867);
or U10805 (N_10805,N_7180,N_5163);
nor U10806 (N_10806,N_4737,N_7825);
nand U10807 (N_10807,N_4302,N_5119);
or U10808 (N_10808,N_6525,N_4704);
nor U10809 (N_10809,N_4147,N_5749);
xor U10810 (N_10810,N_4746,N_5364);
or U10811 (N_10811,N_5803,N_4556);
or U10812 (N_10812,N_7146,N_4103);
nor U10813 (N_10813,N_4157,N_5528);
nor U10814 (N_10814,N_7959,N_5074);
and U10815 (N_10815,N_6835,N_6336);
xnor U10816 (N_10816,N_5735,N_5442);
nand U10817 (N_10817,N_5190,N_6177);
and U10818 (N_10818,N_7342,N_5488);
nor U10819 (N_10819,N_5347,N_5282);
and U10820 (N_10820,N_6808,N_6988);
and U10821 (N_10821,N_7668,N_7851);
nand U10822 (N_10822,N_4595,N_5828);
or U10823 (N_10823,N_4401,N_7856);
xnor U10824 (N_10824,N_6266,N_4453);
nand U10825 (N_10825,N_4573,N_7442);
xnor U10826 (N_10826,N_6382,N_5080);
xnor U10827 (N_10827,N_5963,N_6410);
or U10828 (N_10828,N_7929,N_5723);
or U10829 (N_10829,N_4804,N_6398);
or U10830 (N_10830,N_6726,N_5706);
nand U10831 (N_10831,N_6146,N_7677);
nor U10832 (N_10832,N_7457,N_6637);
nor U10833 (N_10833,N_7713,N_6508);
and U10834 (N_10834,N_6758,N_7104);
nor U10835 (N_10835,N_6849,N_5154);
and U10836 (N_10836,N_5195,N_4493);
nor U10837 (N_10837,N_5442,N_7777);
or U10838 (N_10838,N_4114,N_6942);
and U10839 (N_10839,N_6598,N_4215);
and U10840 (N_10840,N_6453,N_4689);
nor U10841 (N_10841,N_6382,N_7404);
xor U10842 (N_10842,N_6801,N_7572);
nor U10843 (N_10843,N_7204,N_7399);
nand U10844 (N_10844,N_5464,N_5670);
nor U10845 (N_10845,N_4126,N_7949);
and U10846 (N_10846,N_4979,N_5576);
xor U10847 (N_10847,N_5443,N_5161);
or U10848 (N_10848,N_4820,N_6024);
nor U10849 (N_10849,N_4335,N_5303);
or U10850 (N_10850,N_7134,N_7386);
nor U10851 (N_10851,N_7516,N_4111);
xor U10852 (N_10852,N_7577,N_7321);
or U10853 (N_10853,N_5465,N_7089);
and U10854 (N_10854,N_4343,N_7391);
nor U10855 (N_10855,N_5835,N_4698);
or U10856 (N_10856,N_5507,N_4188);
nand U10857 (N_10857,N_7566,N_7764);
xor U10858 (N_10858,N_5837,N_4102);
nor U10859 (N_10859,N_5740,N_5335);
nand U10860 (N_10860,N_4587,N_4371);
xor U10861 (N_10861,N_4010,N_7566);
or U10862 (N_10862,N_7054,N_7145);
nand U10863 (N_10863,N_4880,N_4432);
xor U10864 (N_10864,N_5464,N_4170);
or U10865 (N_10865,N_6881,N_4629);
and U10866 (N_10866,N_4159,N_5210);
or U10867 (N_10867,N_4850,N_4043);
xor U10868 (N_10868,N_7202,N_5378);
nand U10869 (N_10869,N_6563,N_4654);
nor U10870 (N_10870,N_5621,N_4922);
and U10871 (N_10871,N_6332,N_5184);
nand U10872 (N_10872,N_7880,N_7405);
xor U10873 (N_10873,N_5331,N_4084);
or U10874 (N_10874,N_4323,N_4359);
nand U10875 (N_10875,N_7840,N_4174);
xor U10876 (N_10876,N_7181,N_4273);
and U10877 (N_10877,N_4245,N_6261);
or U10878 (N_10878,N_5371,N_7473);
nand U10879 (N_10879,N_7700,N_4666);
nand U10880 (N_10880,N_7264,N_5758);
nand U10881 (N_10881,N_7437,N_7396);
and U10882 (N_10882,N_6471,N_5450);
nand U10883 (N_10883,N_4632,N_5214);
or U10884 (N_10884,N_5222,N_5770);
and U10885 (N_10885,N_4841,N_6688);
or U10886 (N_10886,N_5419,N_6941);
xnor U10887 (N_10887,N_4836,N_6860);
nand U10888 (N_10888,N_6582,N_7495);
nand U10889 (N_10889,N_5568,N_4207);
xor U10890 (N_10890,N_6204,N_5752);
nand U10891 (N_10891,N_7685,N_4894);
and U10892 (N_10892,N_7078,N_4570);
nor U10893 (N_10893,N_6444,N_6206);
nor U10894 (N_10894,N_6958,N_5584);
and U10895 (N_10895,N_7326,N_7468);
xnor U10896 (N_10896,N_7215,N_4425);
xor U10897 (N_10897,N_5139,N_7357);
nand U10898 (N_10898,N_7898,N_6230);
or U10899 (N_10899,N_6638,N_6683);
or U10900 (N_10900,N_6090,N_4591);
and U10901 (N_10901,N_5206,N_5835);
nor U10902 (N_10902,N_7993,N_5429);
xor U10903 (N_10903,N_7272,N_4648);
or U10904 (N_10904,N_6093,N_7445);
nor U10905 (N_10905,N_4766,N_7147);
nor U10906 (N_10906,N_7066,N_5487);
or U10907 (N_10907,N_7245,N_7540);
xor U10908 (N_10908,N_7281,N_7945);
xor U10909 (N_10909,N_5564,N_5424);
nor U10910 (N_10910,N_6025,N_6530);
nor U10911 (N_10911,N_5226,N_7372);
and U10912 (N_10912,N_5825,N_7146);
and U10913 (N_10913,N_5937,N_7561);
nand U10914 (N_10914,N_5825,N_7179);
nand U10915 (N_10915,N_7391,N_6425);
xnor U10916 (N_10916,N_6664,N_6813);
xnor U10917 (N_10917,N_7682,N_4502);
or U10918 (N_10918,N_6987,N_4781);
and U10919 (N_10919,N_5687,N_5355);
nor U10920 (N_10920,N_5457,N_4096);
xnor U10921 (N_10921,N_4533,N_6596);
xor U10922 (N_10922,N_4355,N_7104);
or U10923 (N_10923,N_5451,N_4743);
xnor U10924 (N_10924,N_5075,N_7999);
nor U10925 (N_10925,N_5674,N_5973);
nor U10926 (N_10926,N_5511,N_4277);
xor U10927 (N_10927,N_7452,N_6431);
xnor U10928 (N_10928,N_7712,N_5329);
xor U10929 (N_10929,N_4422,N_5779);
or U10930 (N_10930,N_5494,N_4426);
and U10931 (N_10931,N_7518,N_4052);
nor U10932 (N_10932,N_6107,N_6934);
nor U10933 (N_10933,N_4751,N_7386);
nand U10934 (N_10934,N_7836,N_5443);
or U10935 (N_10935,N_4730,N_7530);
nand U10936 (N_10936,N_6911,N_4626);
nand U10937 (N_10937,N_7188,N_5660);
xnor U10938 (N_10938,N_6709,N_6649);
and U10939 (N_10939,N_6675,N_7086);
or U10940 (N_10940,N_7416,N_6096);
or U10941 (N_10941,N_6144,N_6895);
or U10942 (N_10942,N_6950,N_7905);
xor U10943 (N_10943,N_6812,N_6493);
or U10944 (N_10944,N_5816,N_4975);
nand U10945 (N_10945,N_4222,N_4998);
xor U10946 (N_10946,N_7471,N_6791);
and U10947 (N_10947,N_6151,N_4202);
nand U10948 (N_10948,N_5249,N_4138);
or U10949 (N_10949,N_5467,N_7265);
nor U10950 (N_10950,N_6525,N_7127);
and U10951 (N_10951,N_4648,N_7980);
and U10952 (N_10952,N_7893,N_4377);
nor U10953 (N_10953,N_4986,N_4114);
and U10954 (N_10954,N_5255,N_6447);
nand U10955 (N_10955,N_4605,N_7690);
nor U10956 (N_10956,N_4603,N_7980);
nand U10957 (N_10957,N_4968,N_7422);
nor U10958 (N_10958,N_7939,N_7643);
and U10959 (N_10959,N_7486,N_7941);
nor U10960 (N_10960,N_6090,N_6707);
xor U10961 (N_10961,N_6539,N_7119);
and U10962 (N_10962,N_5435,N_6695);
or U10963 (N_10963,N_5342,N_7200);
xnor U10964 (N_10964,N_6277,N_4498);
xor U10965 (N_10965,N_6084,N_7872);
xor U10966 (N_10966,N_4709,N_5549);
nor U10967 (N_10967,N_7262,N_5637);
and U10968 (N_10968,N_5698,N_4586);
nand U10969 (N_10969,N_5534,N_4293);
and U10970 (N_10970,N_7945,N_6216);
nor U10971 (N_10971,N_7868,N_6893);
nor U10972 (N_10972,N_6751,N_6280);
nor U10973 (N_10973,N_5938,N_4811);
xor U10974 (N_10974,N_6900,N_6981);
xnor U10975 (N_10975,N_4351,N_4175);
xnor U10976 (N_10976,N_5845,N_5258);
nor U10977 (N_10977,N_7009,N_5478);
xnor U10978 (N_10978,N_4833,N_5653);
nand U10979 (N_10979,N_6375,N_4233);
and U10980 (N_10980,N_5041,N_4371);
xnor U10981 (N_10981,N_5093,N_6940);
nand U10982 (N_10982,N_7251,N_4539);
nor U10983 (N_10983,N_4282,N_4619);
nor U10984 (N_10984,N_7811,N_6146);
and U10985 (N_10985,N_5311,N_6492);
or U10986 (N_10986,N_5008,N_4258);
xnor U10987 (N_10987,N_7787,N_7853);
and U10988 (N_10988,N_7115,N_6921);
nor U10989 (N_10989,N_4169,N_6842);
nor U10990 (N_10990,N_7973,N_5157);
and U10991 (N_10991,N_7652,N_4892);
and U10992 (N_10992,N_4240,N_7315);
xnor U10993 (N_10993,N_6054,N_5239);
nor U10994 (N_10994,N_6495,N_5034);
xnor U10995 (N_10995,N_5362,N_4218);
nor U10996 (N_10996,N_7250,N_6135);
or U10997 (N_10997,N_6741,N_7187);
nor U10998 (N_10998,N_5495,N_7801);
xnor U10999 (N_10999,N_7016,N_6805);
xnor U11000 (N_11000,N_4363,N_7927);
nand U11001 (N_11001,N_7045,N_7744);
nand U11002 (N_11002,N_6061,N_5895);
or U11003 (N_11003,N_6957,N_4097);
nand U11004 (N_11004,N_7140,N_6220);
and U11005 (N_11005,N_5581,N_6527);
or U11006 (N_11006,N_5848,N_5306);
and U11007 (N_11007,N_6917,N_6722);
and U11008 (N_11008,N_6467,N_6308);
and U11009 (N_11009,N_5246,N_4474);
nand U11010 (N_11010,N_4309,N_5825);
and U11011 (N_11011,N_7135,N_6716);
xor U11012 (N_11012,N_6413,N_7442);
or U11013 (N_11013,N_7420,N_6579);
nor U11014 (N_11014,N_7976,N_7671);
and U11015 (N_11015,N_7503,N_6689);
nand U11016 (N_11016,N_4731,N_5272);
and U11017 (N_11017,N_6917,N_4634);
nand U11018 (N_11018,N_5119,N_5407);
nand U11019 (N_11019,N_7804,N_6788);
and U11020 (N_11020,N_6817,N_4463);
and U11021 (N_11021,N_7061,N_7047);
or U11022 (N_11022,N_7677,N_7882);
and U11023 (N_11023,N_6439,N_4045);
and U11024 (N_11024,N_4127,N_6933);
nand U11025 (N_11025,N_5279,N_6998);
nand U11026 (N_11026,N_4219,N_4772);
and U11027 (N_11027,N_5179,N_6872);
nor U11028 (N_11028,N_6143,N_4330);
and U11029 (N_11029,N_6534,N_5647);
and U11030 (N_11030,N_4368,N_4423);
or U11031 (N_11031,N_6866,N_7460);
or U11032 (N_11032,N_7013,N_4657);
nor U11033 (N_11033,N_6014,N_5183);
nand U11034 (N_11034,N_6014,N_7829);
and U11035 (N_11035,N_7377,N_7455);
xnor U11036 (N_11036,N_6988,N_6401);
nor U11037 (N_11037,N_5917,N_4922);
xnor U11038 (N_11038,N_7690,N_4473);
xor U11039 (N_11039,N_6685,N_4638);
nor U11040 (N_11040,N_4691,N_4679);
xor U11041 (N_11041,N_4165,N_7601);
nor U11042 (N_11042,N_6983,N_4721);
or U11043 (N_11043,N_7997,N_4611);
and U11044 (N_11044,N_5550,N_6692);
or U11045 (N_11045,N_6690,N_5322);
xnor U11046 (N_11046,N_6205,N_4787);
nor U11047 (N_11047,N_5355,N_5784);
xor U11048 (N_11048,N_4500,N_4221);
and U11049 (N_11049,N_4536,N_5539);
nand U11050 (N_11050,N_6233,N_5181);
and U11051 (N_11051,N_6943,N_6013);
nor U11052 (N_11052,N_5355,N_6793);
xor U11053 (N_11053,N_7634,N_7118);
nand U11054 (N_11054,N_5156,N_6054);
nor U11055 (N_11055,N_6494,N_4376);
or U11056 (N_11056,N_7106,N_5706);
and U11057 (N_11057,N_7631,N_4216);
nand U11058 (N_11058,N_7752,N_7193);
nor U11059 (N_11059,N_7701,N_6775);
or U11060 (N_11060,N_7865,N_7889);
and U11061 (N_11061,N_6763,N_7461);
nor U11062 (N_11062,N_7210,N_5669);
and U11063 (N_11063,N_7691,N_6446);
nand U11064 (N_11064,N_5309,N_6413);
nand U11065 (N_11065,N_6623,N_6279);
and U11066 (N_11066,N_6769,N_6847);
nand U11067 (N_11067,N_5372,N_7641);
nor U11068 (N_11068,N_4098,N_6069);
nand U11069 (N_11069,N_5219,N_5006);
nor U11070 (N_11070,N_4437,N_5247);
xor U11071 (N_11071,N_6992,N_4428);
nand U11072 (N_11072,N_6532,N_4150);
xnor U11073 (N_11073,N_6168,N_7969);
or U11074 (N_11074,N_7701,N_4012);
nor U11075 (N_11075,N_7278,N_7960);
and U11076 (N_11076,N_6143,N_6645);
xor U11077 (N_11077,N_6767,N_6303);
nand U11078 (N_11078,N_5096,N_6979);
nand U11079 (N_11079,N_7379,N_6975);
xor U11080 (N_11080,N_6214,N_4144);
nand U11081 (N_11081,N_7329,N_4276);
or U11082 (N_11082,N_4540,N_4650);
and U11083 (N_11083,N_4165,N_6327);
xnor U11084 (N_11084,N_5746,N_6847);
nor U11085 (N_11085,N_4674,N_7396);
or U11086 (N_11086,N_6508,N_6605);
xnor U11087 (N_11087,N_5357,N_6403);
nand U11088 (N_11088,N_6097,N_5634);
nand U11089 (N_11089,N_6486,N_7885);
or U11090 (N_11090,N_6156,N_7924);
nor U11091 (N_11091,N_4195,N_4778);
nor U11092 (N_11092,N_5475,N_7209);
xor U11093 (N_11093,N_6729,N_4447);
nor U11094 (N_11094,N_4611,N_4431);
or U11095 (N_11095,N_6947,N_7959);
or U11096 (N_11096,N_7048,N_6774);
xor U11097 (N_11097,N_7067,N_7494);
nand U11098 (N_11098,N_7495,N_6439);
xor U11099 (N_11099,N_5707,N_5878);
or U11100 (N_11100,N_6061,N_6228);
nand U11101 (N_11101,N_5383,N_5378);
or U11102 (N_11102,N_6638,N_5845);
xor U11103 (N_11103,N_7854,N_5744);
nor U11104 (N_11104,N_4106,N_6537);
and U11105 (N_11105,N_4072,N_7398);
nor U11106 (N_11106,N_7927,N_6963);
nor U11107 (N_11107,N_7902,N_4267);
nand U11108 (N_11108,N_6278,N_4267);
or U11109 (N_11109,N_7169,N_4406);
nand U11110 (N_11110,N_4867,N_7399);
nand U11111 (N_11111,N_6618,N_4551);
and U11112 (N_11112,N_7697,N_7823);
or U11113 (N_11113,N_7506,N_7502);
or U11114 (N_11114,N_5123,N_7183);
xor U11115 (N_11115,N_7995,N_5401);
or U11116 (N_11116,N_6198,N_6127);
or U11117 (N_11117,N_4930,N_5555);
nand U11118 (N_11118,N_5333,N_4964);
nor U11119 (N_11119,N_7824,N_6161);
nor U11120 (N_11120,N_6739,N_5499);
and U11121 (N_11121,N_7783,N_4564);
nor U11122 (N_11122,N_4219,N_6849);
xor U11123 (N_11123,N_7044,N_5369);
and U11124 (N_11124,N_4062,N_5937);
xor U11125 (N_11125,N_4809,N_6792);
or U11126 (N_11126,N_4672,N_6855);
xnor U11127 (N_11127,N_4154,N_5028);
nor U11128 (N_11128,N_7780,N_6290);
nor U11129 (N_11129,N_5076,N_6940);
nor U11130 (N_11130,N_6556,N_6275);
and U11131 (N_11131,N_5018,N_7716);
xor U11132 (N_11132,N_4740,N_6576);
nor U11133 (N_11133,N_5052,N_7489);
nor U11134 (N_11134,N_7204,N_7866);
and U11135 (N_11135,N_5838,N_6163);
or U11136 (N_11136,N_5036,N_7438);
nand U11137 (N_11137,N_6151,N_6731);
xnor U11138 (N_11138,N_7700,N_6568);
xnor U11139 (N_11139,N_7168,N_4628);
and U11140 (N_11140,N_4276,N_7387);
nor U11141 (N_11141,N_7389,N_4366);
nand U11142 (N_11142,N_4310,N_6251);
or U11143 (N_11143,N_5405,N_4505);
xor U11144 (N_11144,N_7781,N_5377);
xnor U11145 (N_11145,N_4061,N_6749);
or U11146 (N_11146,N_4281,N_5270);
or U11147 (N_11147,N_4311,N_4730);
nand U11148 (N_11148,N_6109,N_5813);
or U11149 (N_11149,N_7511,N_6781);
or U11150 (N_11150,N_7873,N_6693);
and U11151 (N_11151,N_4165,N_5039);
nand U11152 (N_11152,N_4766,N_7452);
and U11153 (N_11153,N_4602,N_7928);
nor U11154 (N_11154,N_7593,N_6897);
or U11155 (N_11155,N_6540,N_6280);
nand U11156 (N_11156,N_5227,N_7213);
xnor U11157 (N_11157,N_5323,N_5050);
nand U11158 (N_11158,N_6743,N_4429);
nand U11159 (N_11159,N_6255,N_7490);
and U11160 (N_11160,N_6051,N_5574);
nor U11161 (N_11161,N_5650,N_7398);
and U11162 (N_11162,N_7380,N_5516);
or U11163 (N_11163,N_5456,N_5289);
or U11164 (N_11164,N_4385,N_7214);
xnor U11165 (N_11165,N_5953,N_4134);
nor U11166 (N_11166,N_6295,N_6707);
and U11167 (N_11167,N_7532,N_5256);
and U11168 (N_11168,N_6019,N_7494);
or U11169 (N_11169,N_5283,N_4094);
nand U11170 (N_11170,N_4630,N_4535);
or U11171 (N_11171,N_6458,N_7987);
nand U11172 (N_11172,N_7421,N_6660);
or U11173 (N_11173,N_4289,N_6750);
and U11174 (N_11174,N_6204,N_4619);
and U11175 (N_11175,N_7278,N_6592);
and U11176 (N_11176,N_5286,N_7323);
xnor U11177 (N_11177,N_4669,N_6553);
xnor U11178 (N_11178,N_4104,N_4691);
or U11179 (N_11179,N_5399,N_4913);
nand U11180 (N_11180,N_7810,N_6371);
or U11181 (N_11181,N_5363,N_7379);
nand U11182 (N_11182,N_6124,N_5573);
xnor U11183 (N_11183,N_4499,N_6651);
xnor U11184 (N_11184,N_5398,N_7781);
and U11185 (N_11185,N_5862,N_6819);
xor U11186 (N_11186,N_5666,N_5806);
nor U11187 (N_11187,N_7515,N_6337);
nand U11188 (N_11188,N_6239,N_5898);
and U11189 (N_11189,N_6082,N_4420);
xnor U11190 (N_11190,N_7899,N_5716);
or U11191 (N_11191,N_4723,N_4032);
xor U11192 (N_11192,N_7492,N_5776);
or U11193 (N_11193,N_4487,N_6132);
or U11194 (N_11194,N_4398,N_5903);
xnor U11195 (N_11195,N_7406,N_6929);
nand U11196 (N_11196,N_5287,N_6335);
xnor U11197 (N_11197,N_4134,N_7815);
xnor U11198 (N_11198,N_7784,N_5093);
and U11199 (N_11199,N_4304,N_4010);
nor U11200 (N_11200,N_4708,N_7656);
nor U11201 (N_11201,N_6458,N_4747);
nor U11202 (N_11202,N_6815,N_6148);
and U11203 (N_11203,N_7175,N_4740);
nor U11204 (N_11204,N_6456,N_6266);
xor U11205 (N_11205,N_4319,N_6435);
and U11206 (N_11206,N_6749,N_4190);
nor U11207 (N_11207,N_7301,N_7750);
and U11208 (N_11208,N_6015,N_7648);
and U11209 (N_11209,N_7694,N_5822);
nor U11210 (N_11210,N_6832,N_5624);
or U11211 (N_11211,N_5821,N_5802);
nor U11212 (N_11212,N_6773,N_4823);
or U11213 (N_11213,N_4318,N_4292);
nand U11214 (N_11214,N_5763,N_6465);
and U11215 (N_11215,N_5085,N_7726);
or U11216 (N_11216,N_6624,N_4512);
xor U11217 (N_11217,N_5616,N_7372);
nor U11218 (N_11218,N_7575,N_4175);
xor U11219 (N_11219,N_7252,N_4571);
xor U11220 (N_11220,N_4053,N_6235);
nor U11221 (N_11221,N_6565,N_5980);
and U11222 (N_11222,N_7310,N_4228);
or U11223 (N_11223,N_5036,N_7833);
or U11224 (N_11224,N_4987,N_7923);
nor U11225 (N_11225,N_7046,N_5367);
or U11226 (N_11226,N_5616,N_4815);
nor U11227 (N_11227,N_7574,N_4232);
and U11228 (N_11228,N_7483,N_6483);
nor U11229 (N_11229,N_5533,N_5375);
or U11230 (N_11230,N_6241,N_7229);
nand U11231 (N_11231,N_4046,N_4981);
nor U11232 (N_11232,N_4263,N_4288);
nor U11233 (N_11233,N_6308,N_5869);
and U11234 (N_11234,N_6161,N_4882);
or U11235 (N_11235,N_7492,N_7770);
or U11236 (N_11236,N_6900,N_5462);
or U11237 (N_11237,N_5996,N_4748);
nor U11238 (N_11238,N_4723,N_4035);
xor U11239 (N_11239,N_6643,N_4551);
nand U11240 (N_11240,N_6104,N_4659);
nor U11241 (N_11241,N_7051,N_5481);
xor U11242 (N_11242,N_7152,N_4950);
and U11243 (N_11243,N_6823,N_4278);
and U11244 (N_11244,N_7707,N_4127);
or U11245 (N_11245,N_4514,N_5340);
xnor U11246 (N_11246,N_6262,N_5520);
nor U11247 (N_11247,N_5743,N_5875);
nand U11248 (N_11248,N_7240,N_6008);
nor U11249 (N_11249,N_6379,N_7211);
nor U11250 (N_11250,N_5190,N_7787);
nand U11251 (N_11251,N_7082,N_4790);
xor U11252 (N_11252,N_7885,N_5613);
and U11253 (N_11253,N_6123,N_4981);
xnor U11254 (N_11254,N_7003,N_6250);
xnor U11255 (N_11255,N_7556,N_4202);
nor U11256 (N_11256,N_6886,N_5954);
or U11257 (N_11257,N_6985,N_5875);
and U11258 (N_11258,N_7111,N_4508);
xor U11259 (N_11259,N_7782,N_4109);
or U11260 (N_11260,N_4611,N_5690);
nor U11261 (N_11261,N_4251,N_7124);
or U11262 (N_11262,N_6326,N_7006);
xnor U11263 (N_11263,N_4392,N_6275);
xnor U11264 (N_11264,N_6779,N_5044);
nor U11265 (N_11265,N_6374,N_6810);
nand U11266 (N_11266,N_6177,N_6790);
xnor U11267 (N_11267,N_5693,N_5726);
nand U11268 (N_11268,N_7515,N_7239);
nand U11269 (N_11269,N_6723,N_7172);
xor U11270 (N_11270,N_7158,N_5399);
xnor U11271 (N_11271,N_6655,N_4334);
and U11272 (N_11272,N_7689,N_5485);
nand U11273 (N_11273,N_6678,N_4501);
and U11274 (N_11274,N_6761,N_7767);
nand U11275 (N_11275,N_4561,N_4141);
nand U11276 (N_11276,N_5174,N_5429);
nor U11277 (N_11277,N_5025,N_6548);
or U11278 (N_11278,N_6554,N_4744);
xor U11279 (N_11279,N_7057,N_6220);
or U11280 (N_11280,N_7000,N_6183);
xor U11281 (N_11281,N_5331,N_4533);
xnor U11282 (N_11282,N_7103,N_4134);
nor U11283 (N_11283,N_4533,N_4073);
nand U11284 (N_11284,N_7119,N_4581);
or U11285 (N_11285,N_6247,N_4754);
nor U11286 (N_11286,N_7330,N_5624);
nor U11287 (N_11287,N_4822,N_5688);
nor U11288 (N_11288,N_4523,N_6271);
nor U11289 (N_11289,N_5148,N_6353);
or U11290 (N_11290,N_7066,N_6788);
xor U11291 (N_11291,N_7696,N_5293);
xor U11292 (N_11292,N_5816,N_7537);
nand U11293 (N_11293,N_6875,N_7762);
and U11294 (N_11294,N_6491,N_5175);
and U11295 (N_11295,N_7292,N_5630);
nand U11296 (N_11296,N_6351,N_5148);
nand U11297 (N_11297,N_6903,N_7982);
nor U11298 (N_11298,N_7533,N_5377);
and U11299 (N_11299,N_7727,N_6019);
or U11300 (N_11300,N_6572,N_7339);
nor U11301 (N_11301,N_7180,N_6796);
xor U11302 (N_11302,N_4234,N_4257);
xor U11303 (N_11303,N_6204,N_6856);
and U11304 (N_11304,N_7254,N_6568);
nor U11305 (N_11305,N_5143,N_5702);
xor U11306 (N_11306,N_5480,N_4676);
nand U11307 (N_11307,N_7192,N_7195);
nand U11308 (N_11308,N_4109,N_4574);
xnor U11309 (N_11309,N_4272,N_5346);
nand U11310 (N_11310,N_4210,N_7233);
or U11311 (N_11311,N_6119,N_6884);
and U11312 (N_11312,N_6153,N_4021);
or U11313 (N_11313,N_5984,N_5114);
nand U11314 (N_11314,N_4153,N_6992);
nand U11315 (N_11315,N_7186,N_7484);
nor U11316 (N_11316,N_5946,N_6961);
or U11317 (N_11317,N_6615,N_4730);
and U11318 (N_11318,N_7997,N_6915);
nand U11319 (N_11319,N_4783,N_6888);
nor U11320 (N_11320,N_7492,N_7890);
or U11321 (N_11321,N_7190,N_4286);
xor U11322 (N_11322,N_5213,N_6566);
nand U11323 (N_11323,N_7839,N_7221);
xor U11324 (N_11324,N_5786,N_5348);
nand U11325 (N_11325,N_6861,N_6926);
xnor U11326 (N_11326,N_5939,N_5793);
xnor U11327 (N_11327,N_5820,N_5409);
nand U11328 (N_11328,N_4625,N_7855);
nand U11329 (N_11329,N_6657,N_6813);
or U11330 (N_11330,N_4112,N_5135);
and U11331 (N_11331,N_7340,N_7480);
and U11332 (N_11332,N_7303,N_5213);
nand U11333 (N_11333,N_4717,N_5772);
nor U11334 (N_11334,N_5736,N_4088);
and U11335 (N_11335,N_6815,N_6180);
or U11336 (N_11336,N_4879,N_5533);
xor U11337 (N_11337,N_7177,N_5407);
or U11338 (N_11338,N_5328,N_6430);
or U11339 (N_11339,N_4313,N_5627);
xnor U11340 (N_11340,N_6474,N_4650);
nand U11341 (N_11341,N_7396,N_7246);
or U11342 (N_11342,N_5827,N_4347);
xor U11343 (N_11343,N_6086,N_6602);
nor U11344 (N_11344,N_6270,N_5467);
xnor U11345 (N_11345,N_5557,N_7143);
and U11346 (N_11346,N_5550,N_7129);
and U11347 (N_11347,N_6184,N_4545);
and U11348 (N_11348,N_5308,N_7264);
nor U11349 (N_11349,N_4523,N_5490);
xor U11350 (N_11350,N_6029,N_5893);
and U11351 (N_11351,N_7802,N_4517);
nor U11352 (N_11352,N_4977,N_7770);
or U11353 (N_11353,N_7905,N_5544);
xor U11354 (N_11354,N_7341,N_5628);
and U11355 (N_11355,N_6220,N_4553);
nand U11356 (N_11356,N_7590,N_6052);
nor U11357 (N_11357,N_4181,N_7426);
nand U11358 (N_11358,N_5721,N_4625);
or U11359 (N_11359,N_7298,N_7334);
nor U11360 (N_11360,N_4057,N_5850);
and U11361 (N_11361,N_7197,N_6169);
and U11362 (N_11362,N_6590,N_6079);
or U11363 (N_11363,N_4245,N_6148);
xnor U11364 (N_11364,N_5131,N_7370);
and U11365 (N_11365,N_5199,N_5101);
nand U11366 (N_11366,N_7258,N_4173);
and U11367 (N_11367,N_4998,N_5813);
or U11368 (N_11368,N_6722,N_7538);
or U11369 (N_11369,N_7584,N_7831);
or U11370 (N_11370,N_7910,N_4610);
nor U11371 (N_11371,N_7126,N_6522);
or U11372 (N_11372,N_6997,N_4427);
nor U11373 (N_11373,N_4907,N_5120);
or U11374 (N_11374,N_5422,N_5839);
or U11375 (N_11375,N_5664,N_7529);
and U11376 (N_11376,N_5460,N_5025);
and U11377 (N_11377,N_6706,N_4774);
or U11378 (N_11378,N_4212,N_7108);
xnor U11379 (N_11379,N_5565,N_5840);
or U11380 (N_11380,N_4738,N_5085);
nand U11381 (N_11381,N_7659,N_7921);
xor U11382 (N_11382,N_5865,N_7284);
nor U11383 (N_11383,N_4902,N_5887);
and U11384 (N_11384,N_4675,N_4238);
and U11385 (N_11385,N_4584,N_4010);
xnor U11386 (N_11386,N_7821,N_4286);
nand U11387 (N_11387,N_6058,N_6374);
nand U11388 (N_11388,N_7376,N_7229);
and U11389 (N_11389,N_5528,N_7213);
nand U11390 (N_11390,N_7843,N_4268);
or U11391 (N_11391,N_4955,N_5017);
nand U11392 (N_11392,N_7833,N_6819);
nor U11393 (N_11393,N_5260,N_4834);
or U11394 (N_11394,N_6058,N_6371);
nor U11395 (N_11395,N_4412,N_6594);
or U11396 (N_11396,N_6156,N_4056);
or U11397 (N_11397,N_6387,N_5138);
or U11398 (N_11398,N_7579,N_4054);
and U11399 (N_11399,N_7831,N_4450);
and U11400 (N_11400,N_4267,N_6465);
and U11401 (N_11401,N_6324,N_7102);
nor U11402 (N_11402,N_6854,N_4692);
nor U11403 (N_11403,N_6055,N_6162);
or U11404 (N_11404,N_7032,N_6535);
xor U11405 (N_11405,N_4700,N_7090);
xnor U11406 (N_11406,N_6368,N_4725);
xnor U11407 (N_11407,N_5583,N_7114);
and U11408 (N_11408,N_7578,N_6040);
and U11409 (N_11409,N_6572,N_6771);
nor U11410 (N_11410,N_4276,N_5037);
nor U11411 (N_11411,N_7336,N_4241);
or U11412 (N_11412,N_4559,N_6279);
or U11413 (N_11413,N_7013,N_4721);
nor U11414 (N_11414,N_5778,N_6444);
xor U11415 (N_11415,N_7871,N_6285);
nor U11416 (N_11416,N_7471,N_4394);
and U11417 (N_11417,N_4130,N_6725);
nor U11418 (N_11418,N_5783,N_7410);
and U11419 (N_11419,N_5242,N_6274);
and U11420 (N_11420,N_6149,N_7183);
nand U11421 (N_11421,N_5650,N_6861);
xnor U11422 (N_11422,N_6038,N_4195);
xor U11423 (N_11423,N_7996,N_7874);
xor U11424 (N_11424,N_4013,N_6576);
nor U11425 (N_11425,N_6142,N_7334);
xor U11426 (N_11426,N_5269,N_4010);
xnor U11427 (N_11427,N_6312,N_5867);
or U11428 (N_11428,N_6521,N_4894);
nor U11429 (N_11429,N_7540,N_6109);
nand U11430 (N_11430,N_5726,N_7046);
and U11431 (N_11431,N_6156,N_5186);
nor U11432 (N_11432,N_6372,N_7850);
or U11433 (N_11433,N_7822,N_5704);
nor U11434 (N_11434,N_4378,N_5027);
xor U11435 (N_11435,N_5150,N_6576);
nand U11436 (N_11436,N_7073,N_6332);
or U11437 (N_11437,N_5527,N_4916);
nor U11438 (N_11438,N_5823,N_6645);
or U11439 (N_11439,N_6210,N_7295);
or U11440 (N_11440,N_4106,N_4614);
nor U11441 (N_11441,N_5413,N_7331);
nand U11442 (N_11442,N_4322,N_5496);
nand U11443 (N_11443,N_4950,N_5927);
or U11444 (N_11444,N_5834,N_6712);
or U11445 (N_11445,N_5176,N_4690);
nand U11446 (N_11446,N_5986,N_4627);
or U11447 (N_11447,N_4903,N_6368);
nor U11448 (N_11448,N_5316,N_5304);
nand U11449 (N_11449,N_4892,N_6665);
xnor U11450 (N_11450,N_7233,N_7828);
nor U11451 (N_11451,N_5759,N_4125);
and U11452 (N_11452,N_4957,N_4400);
xor U11453 (N_11453,N_5070,N_4529);
and U11454 (N_11454,N_5342,N_6138);
or U11455 (N_11455,N_4121,N_5232);
xnor U11456 (N_11456,N_4321,N_5636);
and U11457 (N_11457,N_7049,N_6416);
nand U11458 (N_11458,N_6494,N_4147);
nand U11459 (N_11459,N_7773,N_4620);
nor U11460 (N_11460,N_6490,N_5775);
xnor U11461 (N_11461,N_5857,N_7030);
nand U11462 (N_11462,N_5216,N_6988);
xnor U11463 (N_11463,N_7863,N_4892);
xor U11464 (N_11464,N_7986,N_7992);
nand U11465 (N_11465,N_6836,N_4219);
nand U11466 (N_11466,N_7430,N_7407);
or U11467 (N_11467,N_7242,N_4194);
or U11468 (N_11468,N_6989,N_6524);
and U11469 (N_11469,N_5088,N_6078);
and U11470 (N_11470,N_4031,N_7961);
nand U11471 (N_11471,N_5863,N_5626);
nand U11472 (N_11472,N_7790,N_6129);
nor U11473 (N_11473,N_6136,N_6604);
and U11474 (N_11474,N_7777,N_5259);
nor U11475 (N_11475,N_7466,N_4819);
nand U11476 (N_11476,N_4778,N_5733);
nand U11477 (N_11477,N_7331,N_6696);
or U11478 (N_11478,N_7477,N_7955);
and U11479 (N_11479,N_7172,N_7236);
nand U11480 (N_11480,N_6531,N_4076);
and U11481 (N_11481,N_5457,N_5051);
and U11482 (N_11482,N_4175,N_7987);
xnor U11483 (N_11483,N_7247,N_7896);
and U11484 (N_11484,N_4559,N_7909);
xnor U11485 (N_11485,N_5527,N_6364);
nor U11486 (N_11486,N_4628,N_6456);
xor U11487 (N_11487,N_6951,N_6335);
nor U11488 (N_11488,N_6892,N_4405);
and U11489 (N_11489,N_7595,N_5497);
or U11490 (N_11490,N_7317,N_4540);
xor U11491 (N_11491,N_5318,N_7247);
and U11492 (N_11492,N_5646,N_7227);
xor U11493 (N_11493,N_4614,N_4366);
nor U11494 (N_11494,N_6937,N_5525);
or U11495 (N_11495,N_7678,N_5157);
nand U11496 (N_11496,N_5321,N_7393);
and U11497 (N_11497,N_7911,N_7061);
nor U11498 (N_11498,N_7298,N_7297);
or U11499 (N_11499,N_6780,N_5513);
xnor U11500 (N_11500,N_7300,N_4501);
or U11501 (N_11501,N_6805,N_5577);
nor U11502 (N_11502,N_6651,N_6106);
nand U11503 (N_11503,N_4672,N_5703);
nor U11504 (N_11504,N_5343,N_7129);
and U11505 (N_11505,N_4907,N_7331);
and U11506 (N_11506,N_4183,N_4969);
xnor U11507 (N_11507,N_4121,N_7361);
xnor U11508 (N_11508,N_5065,N_7233);
xor U11509 (N_11509,N_6502,N_6081);
nor U11510 (N_11510,N_5103,N_7857);
and U11511 (N_11511,N_7027,N_4340);
xor U11512 (N_11512,N_6951,N_4536);
and U11513 (N_11513,N_7458,N_5644);
xor U11514 (N_11514,N_5794,N_4043);
nor U11515 (N_11515,N_5076,N_7054);
and U11516 (N_11516,N_6168,N_6069);
or U11517 (N_11517,N_6030,N_6021);
and U11518 (N_11518,N_4933,N_4204);
or U11519 (N_11519,N_5377,N_5287);
xor U11520 (N_11520,N_6064,N_7305);
nand U11521 (N_11521,N_7567,N_7622);
xnor U11522 (N_11522,N_7029,N_7807);
xor U11523 (N_11523,N_6354,N_4267);
nor U11524 (N_11524,N_6833,N_6064);
and U11525 (N_11525,N_6171,N_7350);
and U11526 (N_11526,N_7959,N_5361);
nand U11527 (N_11527,N_5595,N_7095);
and U11528 (N_11528,N_4616,N_4290);
or U11529 (N_11529,N_5371,N_4088);
nor U11530 (N_11530,N_4580,N_6929);
nor U11531 (N_11531,N_5849,N_4562);
nand U11532 (N_11532,N_6834,N_5921);
or U11533 (N_11533,N_4865,N_7483);
nor U11534 (N_11534,N_6948,N_6317);
nor U11535 (N_11535,N_6071,N_5422);
or U11536 (N_11536,N_7347,N_7271);
xor U11537 (N_11537,N_7384,N_7100);
or U11538 (N_11538,N_4380,N_6167);
and U11539 (N_11539,N_6905,N_6436);
and U11540 (N_11540,N_5791,N_4959);
and U11541 (N_11541,N_4864,N_6936);
xor U11542 (N_11542,N_5815,N_7963);
xnor U11543 (N_11543,N_5095,N_4936);
nand U11544 (N_11544,N_4318,N_4446);
xor U11545 (N_11545,N_7265,N_5062);
xnor U11546 (N_11546,N_5560,N_4885);
and U11547 (N_11547,N_7580,N_6720);
nand U11548 (N_11548,N_6625,N_6683);
xor U11549 (N_11549,N_6505,N_4309);
xor U11550 (N_11550,N_4695,N_5791);
nor U11551 (N_11551,N_6741,N_4877);
and U11552 (N_11552,N_5053,N_5454);
xor U11553 (N_11553,N_5626,N_6534);
xor U11554 (N_11554,N_7584,N_7941);
and U11555 (N_11555,N_5133,N_7173);
or U11556 (N_11556,N_5957,N_7582);
nand U11557 (N_11557,N_7153,N_4442);
nor U11558 (N_11558,N_6248,N_6815);
and U11559 (N_11559,N_5682,N_5227);
xnor U11560 (N_11560,N_6388,N_5869);
and U11561 (N_11561,N_6327,N_6445);
xor U11562 (N_11562,N_6896,N_4640);
nand U11563 (N_11563,N_7301,N_5131);
or U11564 (N_11564,N_7312,N_4298);
or U11565 (N_11565,N_5663,N_4011);
nor U11566 (N_11566,N_4010,N_6682);
and U11567 (N_11567,N_6113,N_6355);
nor U11568 (N_11568,N_6143,N_4163);
nand U11569 (N_11569,N_7645,N_4540);
and U11570 (N_11570,N_7765,N_7157);
xor U11571 (N_11571,N_6959,N_4442);
nor U11572 (N_11572,N_4892,N_5667);
and U11573 (N_11573,N_5888,N_4504);
xnor U11574 (N_11574,N_7015,N_4080);
and U11575 (N_11575,N_7462,N_7558);
nor U11576 (N_11576,N_6959,N_6311);
or U11577 (N_11577,N_5750,N_6997);
xor U11578 (N_11578,N_5871,N_4874);
xnor U11579 (N_11579,N_5727,N_5029);
xnor U11580 (N_11580,N_4903,N_5867);
nand U11581 (N_11581,N_7577,N_4796);
and U11582 (N_11582,N_6542,N_6684);
or U11583 (N_11583,N_5369,N_7261);
or U11584 (N_11584,N_7418,N_7859);
xnor U11585 (N_11585,N_6675,N_5857);
nand U11586 (N_11586,N_4947,N_7107);
and U11587 (N_11587,N_6962,N_7849);
or U11588 (N_11588,N_5513,N_5334);
nand U11589 (N_11589,N_7523,N_7143);
and U11590 (N_11590,N_4439,N_4969);
and U11591 (N_11591,N_4550,N_5518);
or U11592 (N_11592,N_6067,N_7585);
nand U11593 (N_11593,N_4566,N_5681);
or U11594 (N_11594,N_7489,N_4219);
nor U11595 (N_11595,N_5999,N_4386);
or U11596 (N_11596,N_4881,N_6641);
nor U11597 (N_11597,N_6017,N_4836);
nor U11598 (N_11598,N_6125,N_4303);
nor U11599 (N_11599,N_6608,N_6538);
or U11600 (N_11600,N_4317,N_5536);
and U11601 (N_11601,N_4761,N_5432);
or U11602 (N_11602,N_7137,N_7427);
or U11603 (N_11603,N_6615,N_5771);
and U11604 (N_11604,N_5222,N_7108);
xnor U11605 (N_11605,N_5057,N_5136);
nand U11606 (N_11606,N_5209,N_4383);
or U11607 (N_11607,N_6628,N_5938);
and U11608 (N_11608,N_5698,N_4241);
nand U11609 (N_11609,N_4645,N_4970);
and U11610 (N_11610,N_5552,N_7754);
and U11611 (N_11611,N_5286,N_4354);
and U11612 (N_11612,N_4594,N_6798);
nand U11613 (N_11613,N_5273,N_7985);
nor U11614 (N_11614,N_4886,N_5632);
and U11615 (N_11615,N_6489,N_7568);
and U11616 (N_11616,N_6867,N_6023);
and U11617 (N_11617,N_5983,N_7652);
nor U11618 (N_11618,N_7419,N_4718);
nand U11619 (N_11619,N_4670,N_7205);
or U11620 (N_11620,N_5055,N_6413);
nand U11621 (N_11621,N_7299,N_5100);
xnor U11622 (N_11622,N_4086,N_4413);
and U11623 (N_11623,N_4064,N_7185);
or U11624 (N_11624,N_5498,N_6506);
xor U11625 (N_11625,N_4562,N_6780);
or U11626 (N_11626,N_4412,N_4632);
nor U11627 (N_11627,N_5698,N_6762);
xor U11628 (N_11628,N_5405,N_6701);
nor U11629 (N_11629,N_7568,N_5553);
and U11630 (N_11630,N_7737,N_6663);
or U11631 (N_11631,N_6497,N_4755);
nor U11632 (N_11632,N_6189,N_7715);
xnor U11633 (N_11633,N_5762,N_4167);
or U11634 (N_11634,N_4949,N_5632);
and U11635 (N_11635,N_7660,N_4614);
or U11636 (N_11636,N_4048,N_5604);
nand U11637 (N_11637,N_4523,N_6566);
or U11638 (N_11638,N_6615,N_7106);
and U11639 (N_11639,N_4826,N_6038);
and U11640 (N_11640,N_6066,N_7860);
xnor U11641 (N_11641,N_4630,N_4171);
nor U11642 (N_11642,N_4566,N_5867);
nand U11643 (N_11643,N_6891,N_6419);
nand U11644 (N_11644,N_4008,N_6466);
xnor U11645 (N_11645,N_4216,N_7522);
and U11646 (N_11646,N_5677,N_6316);
or U11647 (N_11647,N_6176,N_5051);
nor U11648 (N_11648,N_4505,N_6678);
nor U11649 (N_11649,N_4302,N_7546);
nand U11650 (N_11650,N_5447,N_6308);
xor U11651 (N_11651,N_4866,N_6470);
or U11652 (N_11652,N_6099,N_4861);
xor U11653 (N_11653,N_7912,N_5152);
and U11654 (N_11654,N_7990,N_5348);
nor U11655 (N_11655,N_4815,N_5915);
nand U11656 (N_11656,N_7341,N_5572);
xor U11657 (N_11657,N_4986,N_6135);
or U11658 (N_11658,N_5406,N_5665);
and U11659 (N_11659,N_6853,N_7306);
nand U11660 (N_11660,N_4937,N_6386);
nand U11661 (N_11661,N_6885,N_5127);
or U11662 (N_11662,N_4599,N_6367);
nand U11663 (N_11663,N_7875,N_4938);
xor U11664 (N_11664,N_5805,N_6477);
nand U11665 (N_11665,N_4227,N_4965);
and U11666 (N_11666,N_5707,N_5525);
or U11667 (N_11667,N_7919,N_7945);
or U11668 (N_11668,N_7358,N_4733);
and U11669 (N_11669,N_6910,N_4902);
and U11670 (N_11670,N_6664,N_6849);
nor U11671 (N_11671,N_6485,N_6525);
nand U11672 (N_11672,N_7127,N_6337);
xor U11673 (N_11673,N_5331,N_6640);
nor U11674 (N_11674,N_6683,N_6137);
or U11675 (N_11675,N_7223,N_6848);
nor U11676 (N_11676,N_5716,N_4003);
nor U11677 (N_11677,N_5155,N_4482);
and U11678 (N_11678,N_5260,N_5077);
and U11679 (N_11679,N_7818,N_5625);
and U11680 (N_11680,N_5029,N_6253);
or U11681 (N_11681,N_6504,N_5903);
or U11682 (N_11682,N_6690,N_7606);
xor U11683 (N_11683,N_5576,N_7874);
nor U11684 (N_11684,N_7696,N_6520);
or U11685 (N_11685,N_5556,N_5445);
nand U11686 (N_11686,N_7640,N_6454);
xnor U11687 (N_11687,N_6056,N_6738);
nand U11688 (N_11688,N_7341,N_5972);
xnor U11689 (N_11689,N_7437,N_4809);
and U11690 (N_11690,N_4260,N_7829);
and U11691 (N_11691,N_6403,N_4323);
and U11692 (N_11692,N_7261,N_7126);
xnor U11693 (N_11693,N_7300,N_5442);
nand U11694 (N_11694,N_4795,N_4483);
and U11695 (N_11695,N_7236,N_4231);
xor U11696 (N_11696,N_5829,N_6717);
or U11697 (N_11697,N_4776,N_5320);
nor U11698 (N_11698,N_5285,N_6858);
and U11699 (N_11699,N_5088,N_4350);
or U11700 (N_11700,N_5645,N_7051);
xnor U11701 (N_11701,N_4478,N_6993);
or U11702 (N_11702,N_7938,N_5386);
nand U11703 (N_11703,N_4717,N_4884);
xor U11704 (N_11704,N_5824,N_5374);
xnor U11705 (N_11705,N_5436,N_6065);
xnor U11706 (N_11706,N_6359,N_5082);
or U11707 (N_11707,N_5616,N_6274);
or U11708 (N_11708,N_7632,N_4663);
or U11709 (N_11709,N_5247,N_7909);
nand U11710 (N_11710,N_4382,N_5862);
nand U11711 (N_11711,N_4123,N_7288);
nor U11712 (N_11712,N_6788,N_7951);
and U11713 (N_11713,N_5827,N_4333);
nor U11714 (N_11714,N_4415,N_5294);
nand U11715 (N_11715,N_7582,N_6234);
nor U11716 (N_11716,N_6004,N_6377);
xnor U11717 (N_11717,N_4956,N_7836);
and U11718 (N_11718,N_7074,N_5903);
xnor U11719 (N_11719,N_7526,N_6277);
nand U11720 (N_11720,N_4346,N_5650);
xnor U11721 (N_11721,N_4280,N_7715);
nand U11722 (N_11722,N_5620,N_6004);
nand U11723 (N_11723,N_5899,N_6141);
nor U11724 (N_11724,N_4845,N_7845);
nand U11725 (N_11725,N_7625,N_5392);
and U11726 (N_11726,N_6546,N_6561);
and U11727 (N_11727,N_4717,N_5374);
xnor U11728 (N_11728,N_6283,N_4208);
xor U11729 (N_11729,N_6164,N_4467);
nor U11730 (N_11730,N_6561,N_4254);
nand U11731 (N_11731,N_5018,N_4308);
nand U11732 (N_11732,N_6739,N_7227);
xnor U11733 (N_11733,N_6897,N_4822);
nor U11734 (N_11734,N_6541,N_4555);
and U11735 (N_11735,N_5993,N_5442);
and U11736 (N_11736,N_4881,N_5314);
nand U11737 (N_11737,N_4837,N_4788);
or U11738 (N_11738,N_4951,N_5742);
xor U11739 (N_11739,N_6551,N_4960);
and U11740 (N_11740,N_5396,N_5714);
xnor U11741 (N_11741,N_5068,N_5979);
nand U11742 (N_11742,N_6370,N_5239);
xor U11743 (N_11743,N_4834,N_6968);
nand U11744 (N_11744,N_7266,N_6761);
or U11745 (N_11745,N_5446,N_5644);
and U11746 (N_11746,N_7983,N_7764);
or U11747 (N_11747,N_4166,N_4767);
or U11748 (N_11748,N_5243,N_4936);
or U11749 (N_11749,N_4056,N_5285);
xnor U11750 (N_11750,N_7498,N_4391);
xnor U11751 (N_11751,N_4747,N_4572);
and U11752 (N_11752,N_5297,N_6638);
nand U11753 (N_11753,N_7199,N_6167);
nand U11754 (N_11754,N_5674,N_6178);
nand U11755 (N_11755,N_5896,N_7522);
xor U11756 (N_11756,N_4370,N_7407);
nand U11757 (N_11757,N_7949,N_6625);
and U11758 (N_11758,N_5111,N_7587);
nand U11759 (N_11759,N_7055,N_7995);
xor U11760 (N_11760,N_4318,N_7551);
or U11761 (N_11761,N_7179,N_7480);
xor U11762 (N_11762,N_5611,N_4698);
and U11763 (N_11763,N_6472,N_4397);
nand U11764 (N_11764,N_4937,N_5626);
and U11765 (N_11765,N_6199,N_5042);
or U11766 (N_11766,N_4115,N_7404);
xnor U11767 (N_11767,N_4347,N_5753);
nand U11768 (N_11768,N_5884,N_4058);
or U11769 (N_11769,N_6399,N_4394);
nand U11770 (N_11770,N_5017,N_5586);
or U11771 (N_11771,N_4651,N_5224);
xnor U11772 (N_11772,N_4591,N_7792);
nor U11773 (N_11773,N_4800,N_7606);
nand U11774 (N_11774,N_6639,N_5088);
nor U11775 (N_11775,N_4997,N_4984);
and U11776 (N_11776,N_4648,N_5491);
and U11777 (N_11777,N_6612,N_4158);
nand U11778 (N_11778,N_5436,N_6766);
xnor U11779 (N_11779,N_4174,N_5862);
nor U11780 (N_11780,N_4874,N_5917);
and U11781 (N_11781,N_6473,N_7360);
and U11782 (N_11782,N_6518,N_7723);
or U11783 (N_11783,N_7639,N_4021);
nor U11784 (N_11784,N_5132,N_5601);
or U11785 (N_11785,N_5867,N_4803);
nor U11786 (N_11786,N_6462,N_6194);
or U11787 (N_11787,N_5921,N_7195);
nor U11788 (N_11788,N_7569,N_6812);
nor U11789 (N_11789,N_4117,N_4876);
xor U11790 (N_11790,N_4162,N_6502);
nand U11791 (N_11791,N_7746,N_6026);
nand U11792 (N_11792,N_5333,N_5339);
xnor U11793 (N_11793,N_7642,N_6078);
nand U11794 (N_11794,N_6391,N_7543);
xor U11795 (N_11795,N_4763,N_4827);
nor U11796 (N_11796,N_5646,N_5456);
nand U11797 (N_11797,N_4316,N_4667);
nand U11798 (N_11798,N_4614,N_6077);
nor U11799 (N_11799,N_4560,N_7838);
nor U11800 (N_11800,N_7062,N_6162);
nor U11801 (N_11801,N_5813,N_7344);
nand U11802 (N_11802,N_7587,N_7325);
and U11803 (N_11803,N_7947,N_7172);
nor U11804 (N_11804,N_4883,N_7691);
or U11805 (N_11805,N_6346,N_4661);
xor U11806 (N_11806,N_6656,N_5226);
and U11807 (N_11807,N_7171,N_4179);
nor U11808 (N_11808,N_6823,N_6057);
nor U11809 (N_11809,N_5523,N_5810);
nand U11810 (N_11810,N_7124,N_5891);
and U11811 (N_11811,N_6282,N_6164);
xnor U11812 (N_11812,N_6436,N_4298);
nor U11813 (N_11813,N_7004,N_4988);
nor U11814 (N_11814,N_5174,N_6178);
nor U11815 (N_11815,N_6872,N_6102);
nor U11816 (N_11816,N_4685,N_6184);
and U11817 (N_11817,N_4568,N_5203);
and U11818 (N_11818,N_6112,N_4335);
nand U11819 (N_11819,N_5915,N_4995);
nand U11820 (N_11820,N_4206,N_7925);
or U11821 (N_11821,N_7176,N_5590);
or U11822 (N_11822,N_7115,N_5451);
nand U11823 (N_11823,N_7275,N_4487);
or U11824 (N_11824,N_7289,N_5293);
nor U11825 (N_11825,N_4914,N_5152);
nor U11826 (N_11826,N_4081,N_7934);
nand U11827 (N_11827,N_7107,N_6518);
nand U11828 (N_11828,N_6774,N_5992);
xnor U11829 (N_11829,N_7967,N_4769);
and U11830 (N_11830,N_5950,N_6301);
nand U11831 (N_11831,N_5636,N_7219);
nor U11832 (N_11832,N_4642,N_5290);
xnor U11833 (N_11833,N_7689,N_5345);
or U11834 (N_11834,N_4539,N_7153);
nand U11835 (N_11835,N_4771,N_6752);
and U11836 (N_11836,N_5339,N_7648);
nor U11837 (N_11837,N_7343,N_6499);
nand U11838 (N_11838,N_4546,N_7429);
nand U11839 (N_11839,N_7108,N_7718);
nand U11840 (N_11840,N_6265,N_6365);
nor U11841 (N_11841,N_7850,N_6403);
nor U11842 (N_11842,N_4304,N_7944);
nor U11843 (N_11843,N_5719,N_5186);
or U11844 (N_11844,N_4367,N_6472);
xor U11845 (N_11845,N_6826,N_4473);
nor U11846 (N_11846,N_6805,N_7919);
or U11847 (N_11847,N_7383,N_7080);
xnor U11848 (N_11848,N_7865,N_7067);
and U11849 (N_11849,N_4525,N_6134);
nand U11850 (N_11850,N_6407,N_7877);
nand U11851 (N_11851,N_7504,N_7087);
and U11852 (N_11852,N_6899,N_4661);
xor U11853 (N_11853,N_7532,N_7714);
and U11854 (N_11854,N_6349,N_6959);
or U11855 (N_11855,N_7508,N_6165);
xor U11856 (N_11856,N_5104,N_5764);
and U11857 (N_11857,N_5714,N_7818);
and U11858 (N_11858,N_6134,N_7712);
nor U11859 (N_11859,N_5300,N_7454);
and U11860 (N_11860,N_7429,N_6553);
or U11861 (N_11861,N_7416,N_6463);
nand U11862 (N_11862,N_5847,N_5480);
nor U11863 (N_11863,N_5657,N_4170);
and U11864 (N_11864,N_4850,N_5182);
nand U11865 (N_11865,N_5867,N_7022);
or U11866 (N_11866,N_4371,N_5619);
nand U11867 (N_11867,N_5954,N_4473);
nand U11868 (N_11868,N_6601,N_7916);
nor U11869 (N_11869,N_7348,N_4295);
nand U11870 (N_11870,N_4887,N_5782);
nand U11871 (N_11871,N_4295,N_4496);
xnor U11872 (N_11872,N_7017,N_4116);
nand U11873 (N_11873,N_4398,N_6218);
xor U11874 (N_11874,N_7866,N_7043);
and U11875 (N_11875,N_6241,N_4608);
nor U11876 (N_11876,N_7316,N_6876);
nor U11877 (N_11877,N_7395,N_5938);
nand U11878 (N_11878,N_7595,N_4149);
or U11879 (N_11879,N_4267,N_4977);
nor U11880 (N_11880,N_4430,N_4268);
nand U11881 (N_11881,N_4888,N_5699);
nor U11882 (N_11882,N_4358,N_4908);
nand U11883 (N_11883,N_5754,N_4680);
xor U11884 (N_11884,N_4625,N_5377);
nor U11885 (N_11885,N_7616,N_6445);
xor U11886 (N_11886,N_4828,N_4217);
nor U11887 (N_11887,N_5665,N_4031);
nand U11888 (N_11888,N_6159,N_6465);
xnor U11889 (N_11889,N_4829,N_7634);
nor U11890 (N_11890,N_4183,N_7696);
or U11891 (N_11891,N_6962,N_5588);
or U11892 (N_11892,N_6515,N_7407);
nand U11893 (N_11893,N_6994,N_7395);
and U11894 (N_11894,N_6744,N_5063);
xnor U11895 (N_11895,N_6526,N_4271);
or U11896 (N_11896,N_4757,N_7820);
xnor U11897 (N_11897,N_5239,N_7788);
nor U11898 (N_11898,N_5625,N_7716);
xor U11899 (N_11899,N_5723,N_4508);
or U11900 (N_11900,N_4193,N_5055);
xor U11901 (N_11901,N_5574,N_7618);
nand U11902 (N_11902,N_7262,N_6547);
nor U11903 (N_11903,N_5524,N_6613);
nand U11904 (N_11904,N_4321,N_6992);
nand U11905 (N_11905,N_4487,N_4892);
nor U11906 (N_11906,N_6887,N_5643);
nor U11907 (N_11907,N_5778,N_7021);
and U11908 (N_11908,N_7477,N_6536);
xnor U11909 (N_11909,N_5904,N_4317);
xor U11910 (N_11910,N_4643,N_7685);
and U11911 (N_11911,N_4145,N_6562);
and U11912 (N_11912,N_6444,N_7378);
and U11913 (N_11913,N_7761,N_7444);
or U11914 (N_11914,N_6171,N_5643);
and U11915 (N_11915,N_5067,N_5170);
nand U11916 (N_11916,N_5071,N_5181);
or U11917 (N_11917,N_5740,N_7958);
xnor U11918 (N_11918,N_7067,N_5727);
nand U11919 (N_11919,N_4053,N_7009);
nor U11920 (N_11920,N_4622,N_5441);
xnor U11921 (N_11921,N_7192,N_6953);
and U11922 (N_11922,N_4732,N_7918);
and U11923 (N_11923,N_6277,N_7888);
or U11924 (N_11924,N_4869,N_6437);
nor U11925 (N_11925,N_6675,N_6732);
nand U11926 (N_11926,N_7882,N_6500);
or U11927 (N_11927,N_4315,N_5289);
and U11928 (N_11928,N_5920,N_7637);
nand U11929 (N_11929,N_4941,N_7056);
nand U11930 (N_11930,N_7531,N_5791);
xnor U11931 (N_11931,N_6150,N_5921);
and U11932 (N_11932,N_4690,N_7933);
nor U11933 (N_11933,N_4781,N_4820);
and U11934 (N_11934,N_5458,N_7701);
nand U11935 (N_11935,N_5342,N_7902);
or U11936 (N_11936,N_7937,N_6045);
and U11937 (N_11937,N_5274,N_7532);
nor U11938 (N_11938,N_7544,N_5452);
and U11939 (N_11939,N_4259,N_6933);
and U11940 (N_11940,N_4459,N_5561);
or U11941 (N_11941,N_4315,N_5366);
nor U11942 (N_11942,N_5836,N_7251);
or U11943 (N_11943,N_6759,N_4125);
and U11944 (N_11944,N_4841,N_5104);
and U11945 (N_11945,N_7465,N_5641);
and U11946 (N_11946,N_5373,N_5743);
or U11947 (N_11947,N_4773,N_6251);
and U11948 (N_11948,N_5265,N_6901);
xor U11949 (N_11949,N_6244,N_7580);
nor U11950 (N_11950,N_7059,N_5467);
nor U11951 (N_11951,N_5406,N_6736);
nand U11952 (N_11952,N_6015,N_7592);
and U11953 (N_11953,N_6745,N_6706);
or U11954 (N_11954,N_7895,N_6825);
xnor U11955 (N_11955,N_5863,N_7606);
or U11956 (N_11956,N_4346,N_4711);
nor U11957 (N_11957,N_6606,N_7549);
xnor U11958 (N_11958,N_7110,N_5499);
or U11959 (N_11959,N_5547,N_5595);
nand U11960 (N_11960,N_4979,N_4804);
and U11961 (N_11961,N_4752,N_5083);
and U11962 (N_11962,N_6377,N_4018);
or U11963 (N_11963,N_5947,N_5871);
xor U11964 (N_11964,N_6564,N_5286);
xor U11965 (N_11965,N_6959,N_7915);
nor U11966 (N_11966,N_4127,N_7530);
xor U11967 (N_11967,N_4660,N_7021);
or U11968 (N_11968,N_4873,N_4104);
xor U11969 (N_11969,N_6603,N_4406);
nor U11970 (N_11970,N_5876,N_6571);
xor U11971 (N_11971,N_7129,N_6715);
and U11972 (N_11972,N_6962,N_4567);
nand U11973 (N_11973,N_4233,N_5903);
nor U11974 (N_11974,N_6917,N_4869);
nor U11975 (N_11975,N_6375,N_5408);
and U11976 (N_11976,N_5727,N_4788);
and U11977 (N_11977,N_5300,N_7977);
and U11978 (N_11978,N_6592,N_7878);
nor U11979 (N_11979,N_5872,N_7199);
and U11980 (N_11980,N_7335,N_5697);
and U11981 (N_11981,N_6599,N_4882);
or U11982 (N_11982,N_4892,N_6379);
or U11983 (N_11983,N_6285,N_4514);
nand U11984 (N_11984,N_4619,N_5431);
nor U11985 (N_11985,N_6782,N_5342);
xnor U11986 (N_11986,N_7197,N_7460);
nor U11987 (N_11987,N_6598,N_6225);
nor U11988 (N_11988,N_6427,N_5441);
xor U11989 (N_11989,N_7641,N_4138);
and U11990 (N_11990,N_5355,N_6538);
nor U11991 (N_11991,N_5658,N_4266);
or U11992 (N_11992,N_7616,N_5320);
or U11993 (N_11993,N_7513,N_5938);
nand U11994 (N_11994,N_5229,N_6245);
nor U11995 (N_11995,N_6805,N_6549);
or U11996 (N_11996,N_6711,N_7886);
or U11997 (N_11997,N_5430,N_5973);
or U11998 (N_11998,N_6350,N_4131);
nand U11999 (N_11999,N_6524,N_7799);
xnor U12000 (N_12000,N_9210,N_11879);
or U12001 (N_12001,N_8752,N_9810);
xor U12002 (N_12002,N_10858,N_11644);
nand U12003 (N_12003,N_9305,N_11771);
xor U12004 (N_12004,N_8213,N_10189);
nand U12005 (N_12005,N_8854,N_10853);
or U12006 (N_12006,N_10210,N_8682);
or U12007 (N_12007,N_9191,N_9819);
nor U12008 (N_12008,N_9877,N_10876);
or U12009 (N_12009,N_10218,N_9226);
or U12010 (N_12010,N_11254,N_9738);
or U12011 (N_12011,N_9044,N_9826);
and U12012 (N_12012,N_9295,N_9190);
and U12013 (N_12013,N_11448,N_9055);
nand U12014 (N_12014,N_8039,N_8830);
xor U12015 (N_12015,N_9591,N_8360);
or U12016 (N_12016,N_8327,N_9304);
and U12017 (N_12017,N_11616,N_10840);
xor U12018 (N_12018,N_11760,N_9776);
nand U12019 (N_12019,N_10751,N_10983);
and U12020 (N_12020,N_10686,N_9629);
xnor U12021 (N_12021,N_9575,N_11449);
nor U12022 (N_12022,N_9496,N_10208);
and U12023 (N_12023,N_8340,N_9025);
and U12024 (N_12024,N_11047,N_10545);
and U12025 (N_12025,N_9759,N_8399);
nor U12026 (N_12026,N_11208,N_10167);
and U12027 (N_12027,N_8933,N_9834);
xor U12028 (N_12028,N_8126,N_8827);
xnor U12029 (N_12029,N_9925,N_9288);
nand U12030 (N_12030,N_11442,N_10359);
xnor U12031 (N_12031,N_8432,N_9658);
xnor U12032 (N_12032,N_10364,N_9660);
and U12033 (N_12033,N_9988,N_10395);
nand U12034 (N_12034,N_11728,N_11375);
nor U12035 (N_12035,N_9214,N_10910);
xnor U12036 (N_12036,N_10258,N_10644);
nor U12037 (N_12037,N_11466,N_9487);
nand U12038 (N_12038,N_8942,N_11832);
xnor U12039 (N_12039,N_11193,N_11532);
xor U12040 (N_12040,N_8685,N_10382);
and U12041 (N_12041,N_11994,N_11107);
nor U12042 (N_12042,N_9987,N_10112);
xor U12043 (N_12043,N_10308,N_9897);
or U12044 (N_12044,N_8008,N_8531);
nand U12045 (N_12045,N_11389,N_10367);
and U12046 (N_12046,N_8655,N_9884);
and U12047 (N_12047,N_10078,N_8634);
nand U12048 (N_12048,N_11020,N_10832);
nor U12049 (N_12049,N_9491,N_10997);
nor U12050 (N_12050,N_10544,N_10996);
nor U12051 (N_12051,N_11735,N_10214);
nand U12052 (N_12052,N_8737,N_8012);
xnor U12053 (N_12053,N_8461,N_9871);
and U12054 (N_12054,N_11804,N_11428);
xor U12055 (N_12055,N_8811,N_8603);
nand U12056 (N_12056,N_9346,N_8601);
nand U12057 (N_12057,N_9708,N_10192);
or U12058 (N_12058,N_9493,N_10804);
xnor U12059 (N_12059,N_8688,N_11534);
nand U12060 (N_12060,N_11516,N_8349);
nor U12061 (N_12061,N_10135,N_8224);
nor U12062 (N_12062,N_11163,N_11624);
nand U12063 (N_12063,N_8810,N_8179);
nand U12064 (N_12064,N_11109,N_10877);
xor U12065 (N_12065,N_10689,N_10289);
or U12066 (N_12066,N_10375,N_10119);
xor U12067 (N_12067,N_11517,N_11803);
nand U12068 (N_12068,N_11656,N_8951);
or U12069 (N_12069,N_11553,N_8333);
nor U12070 (N_12070,N_8540,N_11768);
and U12071 (N_12071,N_8211,N_8476);
nor U12072 (N_12072,N_8772,N_10620);
nor U12073 (N_12073,N_11403,N_10727);
or U12074 (N_12074,N_8185,N_11593);
or U12075 (N_12075,N_8734,N_9456);
or U12076 (N_12076,N_8940,N_8521);
xnor U12077 (N_12077,N_11826,N_10144);
nor U12078 (N_12078,N_10764,N_8938);
nor U12079 (N_12079,N_10777,N_8516);
nor U12080 (N_12080,N_10496,N_8896);
xnor U12081 (N_12081,N_8394,N_10940);
or U12082 (N_12082,N_10589,N_8163);
nor U12083 (N_12083,N_9771,N_9885);
or U12084 (N_12084,N_9447,N_11342);
nand U12085 (N_12085,N_8803,N_8853);
nand U12086 (N_12086,N_10455,N_10046);
xor U12087 (N_12087,N_8209,N_8716);
nand U12088 (N_12088,N_8985,N_10713);
nand U12089 (N_12089,N_10965,N_8554);
xor U12090 (N_12090,N_8496,N_11506);
nand U12091 (N_12091,N_11155,N_11789);
nand U12092 (N_12092,N_8148,N_11078);
nor U12093 (N_12093,N_11296,N_11714);
or U12094 (N_12094,N_8373,N_9898);
nand U12095 (N_12095,N_11695,N_10153);
or U12096 (N_12096,N_10197,N_8868);
xnor U12097 (N_12097,N_11142,N_10328);
xnor U12098 (N_12098,N_9281,N_10216);
or U12099 (N_12099,N_11810,N_11878);
nand U12100 (N_12100,N_10401,N_8460);
xor U12101 (N_12101,N_9704,N_8676);
and U12102 (N_12102,N_9382,N_9809);
or U12103 (N_12103,N_11373,N_10571);
and U12104 (N_12104,N_9169,N_11190);
and U12105 (N_12105,N_11625,N_9015);
and U12106 (N_12106,N_10019,N_11858);
and U12107 (N_12107,N_8296,N_9774);
xor U12108 (N_12108,N_10986,N_8489);
nand U12109 (N_12109,N_9541,N_11010);
xnor U12110 (N_12110,N_10896,N_9912);
or U12111 (N_12111,N_8992,N_8654);
and U12112 (N_12112,N_9034,N_11178);
nand U12113 (N_12113,N_11212,N_9260);
xor U12114 (N_12114,N_10150,N_9934);
or U12115 (N_12115,N_8721,N_10419);
nor U12116 (N_12116,N_10411,N_11834);
or U12117 (N_12117,N_8825,N_9802);
xor U12118 (N_12118,N_8692,N_11259);
nand U12119 (N_12119,N_11673,N_11014);
and U12120 (N_12120,N_10169,N_10176);
nor U12121 (N_12121,N_11898,N_11774);
xor U12122 (N_12122,N_8826,N_11947);
and U12123 (N_12123,N_9749,N_11817);
nor U12124 (N_12124,N_9383,N_10662);
and U12125 (N_12125,N_8695,N_11585);
and U12126 (N_12126,N_9948,N_10259);
or U12127 (N_12127,N_11577,N_10861);
nand U12128 (N_12128,N_10528,N_11042);
nor U12129 (N_12129,N_11022,N_9828);
nand U12130 (N_12130,N_11393,N_9961);
nor U12131 (N_12131,N_9065,N_8573);
nor U12132 (N_12132,N_11647,N_10323);
or U12133 (N_12133,N_8819,N_11380);
nand U12134 (N_12134,N_9110,N_11230);
nor U12135 (N_12135,N_10392,N_11753);
or U12136 (N_12136,N_11521,N_8212);
nor U12137 (N_12137,N_9521,N_10527);
xnor U12138 (N_12138,N_10475,N_11678);
or U12139 (N_12139,N_8608,N_11362);
xor U12140 (N_12140,N_11173,N_10386);
or U12141 (N_12141,N_11750,N_10533);
nor U12142 (N_12142,N_10261,N_10546);
xor U12143 (N_12143,N_10989,N_9113);
or U12144 (N_12144,N_10498,N_8999);
xnor U12145 (N_12145,N_11037,N_10802);
xor U12146 (N_12146,N_10909,N_9402);
xnor U12147 (N_12147,N_9659,N_11475);
nand U12148 (N_12148,N_11043,N_11946);
nor U12149 (N_12149,N_8059,N_8511);
and U12150 (N_12150,N_10449,N_10124);
and U12151 (N_12151,N_11836,N_9098);
or U12152 (N_12152,N_11901,N_11361);
nand U12153 (N_12153,N_8917,N_9911);
xor U12154 (N_12154,N_11665,N_8108);
nor U12155 (N_12155,N_9276,N_8323);
or U12156 (N_12156,N_11662,N_8606);
xor U12157 (N_12157,N_9822,N_11162);
nand U12158 (N_12158,N_10347,N_10785);
xnor U12159 (N_12159,N_11443,N_9378);
or U12160 (N_12160,N_10915,N_11036);
nor U12161 (N_12161,N_11423,N_11351);
nand U12162 (N_12162,N_9931,N_8863);
nor U12163 (N_12163,N_8056,N_10302);
and U12164 (N_12164,N_8989,N_11346);
xor U12165 (N_12165,N_10211,N_9386);
nor U12166 (N_12166,N_9202,N_11217);
nand U12167 (N_12167,N_9365,N_10201);
xnor U12168 (N_12168,N_11387,N_11120);
xor U12169 (N_12169,N_9435,N_8892);
nand U12170 (N_12170,N_8096,N_9976);
or U12171 (N_12171,N_11811,N_8230);
or U12172 (N_12172,N_11830,N_8534);
nor U12173 (N_12173,N_9620,N_11893);
nand U12174 (N_12174,N_11089,N_11374);
xnor U12175 (N_12175,N_8062,N_10241);
nand U12176 (N_12176,N_11298,N_10806);
or U12177 (N_12177,N_9886,N_10735);
and U12178 (N_12178,N_8034,N_8283);
and U12179 (N_12179,N_8684,N_10405);
or U12180 (N_12180,N_8481,N_10518);
nand U12181 (N_12181,N_10280,N_9020);
and U12182 (N_12182,N_10768,N_9263);
nor U12183 (N_12183,N_10358,N_11177);
and U12184 (N_12184,N_11667,N_9547);
nor U12185 (N_12185,N_8229,N_8488);
xor U12186 (N_12186,N_10257,N_10038);
and U12187 (N_12187,N_8404,N_8510);
xnor U12188 (N_12188,N_10672,N_9322);
nor U12189 (N_12189,N_9280,N_10604);
xnor U12190 (N_12190,N_8932,N_10174);
xor U12191 (N_12191,N_11936,N_8262);
nand U12192 (N_12192,N_10142,N_11966);
and U12193 (N_12193,N_10331,N_8670);
xor U12194 (N_12194,N_8272,N_10959);
and U12195 (N_12195,N_8709,N_9565);
xnor U12196 (N_12196,N_11454,N_11397);
or U12197 (N_12197,N_11845,N_10229);
nand U12198 (N_12198,N_11228,N_8016);
xnor U12199 (N_12199,N_9852,N_8468);
nand U12200 (N_12200,N_11145,N_9520);
nor U12201 (N_12201,N_9782,N_10605);
nand U12202 (N_12202,N_10015,N_10775);
nand U12203 (N_12203,N_11911,N_9067);
or U12204 (N_12204,N_9985,N_11694);
and U12205 (N_12205,N_11088,N_8547);
and U12206 (N_12206,N_11158,N_10456);
and U12207 (N_12207,N_8828,N_9615);
xor U12208 (N_12208,N_9082,N_10140);
or U12209 (N_12209,N_8395,N_9395);
nand U12210 (N_12210,N_11824,N_8382);
xor U12211 (N_12211,N_8028,N_8623);
nor U12212 (N_12212,N_8733,N_11045);
or U12213 (N_12213,N_10512,N_10776);
nand U12214 (N_12214,N_8894,N_9361);
nand U12215 (N_12215,N_9740,N_9939);
nand U12216 (N_12216,N_8440,N_10937);
xor U12217 (N_12217,N_8485,N_10948);
xor U12218 (N_12218,N_11666,N_8385);
xnor U12219 (N_12219,N_10998,N_8639);
nand U12220 (N_12220,N_10137,N_8638);
nor U12221 (N_12221,N_8741,N_8015);
or U12222 (N_12222,N_8788,N_9194);
and U12223 (N_12223,N_10579,N_8832);
nor U12224 (N_12224,N_10324,N_8313);
nand U12225 (N_12225,N_8881,N_8591);
or U12226 (N_12226,N_8282,N_10575);
or U12227 (N_12227,N_11295,N_9879);
and U12228 (N_12228,N_9420,N_9794);
nand U12229 (N_12229,N_11419,N_8033);
or U12230 (N_12230,N_9061,N_10227);
nand U12231 (N_12231,N_9176,N_10326);
or U12232 (N_12232,N_10924,N_10655);
and U12233 (N_12233,N_11823,N_8689);
nor U12234 (N_12234,N_8957,N_11251);
and U12235 (N_12235,N_11060,N_10875);
nand U12236 (N_12236,N_10685,N_8928);
or U12237 (N_12237,N_8668,N_10251);
nand U12238 (N_12238,N_10509,N_8533);
nor U12239 (N_12239,N_10448,N_11490);
or U12240 (N_12240,N_11535,N_10946);
and U12241 (N_12241,N_10616,N_10103);
nor U12242 (N_12242,N_11725,N_11329);
or U12243 (N_12243,N_9648,N_11359);
xor U12244 (N_12244,N_10559,N_8646);
nand U12245 (N_12245,N_8783,N_8414);
xnor U12246 (N_12246,N_11659,N_11336);
or U12247 (N_12247,N_9423,N_9422);
nand U12248 (N_12248,N_8030,N_8377);
xor U12249 (N_12249,N_8982,N_11224);
nand U12250 (N_12250,N_9144,N_9803);
nor U12251 (N_12251,N_9882,N_11438);
xnor U12252 (N_12252,N_8746,N_11341);
nand U12253 (N_12253,N_9369,N_8838);
xnor U12254 (N_12254,N_8066,N_9303);
nor U12255 (N_12255,N_10893,N_10346);
or U12256 (N_12256,N_8870,N_9631);
xor U12257 (N_12257,N_8268,N_9392);
or U12258 (N_12258,N_10995,N_11791);
nor U12259 (N_12259,N_9237,N_11460);
or U12260 (N_12260,N_9855,N_10511);
xor U12261 (N_12261,N_8437,N_11903);
nand U12262 (N_12262,N_10584,N_8374);
nor U12263 (N_12263,N_9559,N_9696);
nand U12264 (N_12264,N_11222,N_10851);
nand U12265 (N_12265,N_10220,N_9998);
nor U12266 (N_12266,N_8107,N_10154);
or U12267 (N_12267,N_10428,N_11703);
xor U12268 (N_12268,N_10637,N_11692);
xnor U12269 (N_12269,N_10580,N_9503);
nand U12270 (N_12270,N_8072,N_8890);
or U12271 (N_12271,N_11793,N_9319);
nand U12272 (N_12272,N_8605,N_9117);
xor U12273 (N_12273,N_10706,N_9846);
or U12274 (N_12274,N_9690,N_11052);
and U12275 (N_12275,N_8088,N_8009);
or U12276 (N_12276,N_8543,N_10157);
nand U12277 (N_12277,N_10325,N_10415);
xnor U12278 (N_12278,N_9108,N_8402);
nor U12279 (N_12279,N_8233,N_11900);
xor U12280 (N_12280,N_8356,N_8666);
nor U12281 (N_12281,N_10636,N_8998);
or U12282 (N_12282,N_8273,N_10809);
xnor U12283 (N_12283,N_8883,N_9761);
or U12284 (N_12284,N_8473,N_9120);
or U12285 (N_12285,N_8410,N_10994);
nand U12286 (N_12286,N_10118,N_8791);
nor U12287 (N_12287,N_8934,N_10178);
nor U12288 (N_12288,N_9730,N_10281);
xnor U12289 (N_12289,N_11256,N_8344);
xor U12290 (N_12290,N_8099,N_10502);
or U12291 (N_12291,N_8845,N_10856);
xor U12292 (N_12292,N_10705,N_11323);
nor U12293 (N_12293,N_10837,N_9011);
xnor U12294 (N_12294,N_10035,N_11431);
xnor U12295 (N_12295,N_10606,N_8627);
xor U12296 (N_12296,N_10357,N_10477);
nand U12297 (N_12297,N_10868,N_11710);
and U12298 (N_12298,N_9125,N_8659);
or U12299 (N_12299,N_9849,N_10133);
xnor U12300 (N_12300,N_11634,N_9012);
nor U12301 (N_12301,N_10671,N_10440);
or U12302 (N_12302,N_11343,N_10481);
nand U12303 (N_12303,N_10447,N_11300);
or U12304 (N_12304,N_10129,N_10017);
or U12305 (N_12305,N_9760,N_10731);
xnor U12306 (N_12306,N_11123,N_9607);
or U12307 (N_12307,N_9285,N_9102);
nor U12308 (N_12308,N_10060,N_8095);
nand U12309 (N_12309,N_10245,N_11927);
nor U12310 (N_12310,N_11138,N_8071);
nor U12311 (N_12311,N_10435,N_9236);
and U12312 (N_12312,N_8271,N_9376);
and U12313 (N_12313,N_10399,N_11648);
xnor U12314 (N_12314,N_8937,N_10563);
nor U12315 (N_12315,N_8119,N_9189);
nand U12316 (N_12316,N_10212,N_11497);
nor U12317 (N_12317,N_10618,N_11627);
and U12318 (N_12318,N_11481,N_9890);
and U12319 (N_12319,N_11675,N_8831);
or U12320 (N_12320,N_8795,N_8816);
and U12321 (N_12321,N_8002,N_8541);
xnor U12322 (N_12322,N_10075,N_8875);
and U12323 (N_12323,N_9235,N_9996);
or U12324 (N_12324,N_10188,N_8156);
xnor U12325 (N_12325,N_10491,N_10539);
nand U12326 (N_12326,N_10792,N_8352);
xor U12327 (N_12327,N_10478,N_8723);
or U12328 (N_12328,N_11701,N_8031);
and U12329 (N_12329,N_8117,N_9397);
xnor U12330 (N_12330,N_11087,N_11776);
xnor U12331 (N_12331,N_11463,N_10221);
or U12332 (N_12332,N_10404,N_9045);
xor U12333 (N_12333,N_10132,N_8140);
and U12334 (N_12334,N_9465,N_9657);
and U12335 (N_12335,N_11595,N_8434);
and U12336 (N_12336,N_9875,N_10818);
and U12337 (N_12337,N_9406,N_11621);
xor U12338 (N_12338,N_10143,N_8864);
or U12339 (N_12339,N_11293,N_8103);
nand U12340 (N_12340,N_10950,N_9843);
nand U12341 (N_12341,N_11513,N_10973);
and U12342 (N_12342,N_11842,N_11320);
xor U12343 (N_12343,N_8758,N_9311);
nor U12344 (N_12344,N_11603,N_11289);
or U12345 (N_12345,N_10101,N_11896);
nand U12346 (N_12346,N_9043,N_9229);
xnor U12347 (N_12347,N_9059,N_10508);
nor U12348 (N_12348,N_8181,N_9078);
nor U12349 (N_12349,N_11887,N_9312);
or U12350 (N_12350,N_10391,N_9531);
xnor U12351 (N_12351,N_8426,N_8368);
or U12352 (N_12352,N_8898,N_9825);
nor U12353 (N_12353,N_10005,N_11097);
xor U12354 (N_12354,N_10473,N_9715);
or U12355 (N_12355,N_11924,N_9164);
and U12356 (N_12356,N_8529,N_10844);
nor U12357 (N_12357,N_11294,N_8930);
nand U12358 (N_12358,N_11417,N_9789);
and U12359 (N_12359,N_9293,N_10433);
nor U12360 (N_12360,N_10901,N_9743);
or U12361 (N_12361,N_9056,N_8701);
nor U12362 (N_12362,N_11129,N_9146);
nand U12363 (N_12363,N_8401,N_10138);
xor U12364 (N_12364,N_11827,N_8202);
or U12365 (N_12365,N_11040,N_9734);
or U12366 (N_12366,N_9244,N_8435);
xor U12367 (N_12367,N_8077,N_10656);
xor U12368 (N_12368,N_8051,N_11649);
nor U12369 (N_12369,N_11007,N_8680);
nor U12370 (N_12370,N_8157,N_10013);
xnor U12371 (N_12371,N_8580,N_8790);
nand U12372 (N_12372,N_10369,N_8593);
or U12373 (N_12373,N_10532,N_9112);
and U12374 (N_12374,N_8495,N_10457);
nor U12375 (N_12375,N_10388,N_9905);
nor U12376 (N_12376,N_10266,N_8466);
or U12377 (N_12377,N_10665,N_11070);
or U12378 (N_12378,N_11274,N_10865);
and U12379 (N_12379,N_11591,N_11169);
nor U12380 (N_12380,N_11601,N_11670);
nand U12381 (N_12381,N_10761,N_9997);
xnor U12382 (N_12382,N_8455,N_8923);
and U12383 (N_12383,N_10315,N_11385);
xor U12384 (N_12384,N_11058,N_9798);
nor U12385 (N_12385,N_11050,N_10554);
nand U12386 (N_12386,N_9611,N_8147);
and U12387 (N_12387,N_10343,N_10814);
nand U12388 (N_12388,N_9929,N_10413);
nor U12389 (N_12389,N_11574,N_8208);
xor U12390 (N_12390,N_11583,N_10274);
nor U12391 (N_12391,N_8472,N_8199);
nand U12392 (N_12392,N_10161,N_10849);
and U12393 (N_12393,N_8740,N_11566);
or U12394 (N_12394,N_11757,N_10933);
xor U12395 (N_12395,N_10892,N_8755);
and U12396 (N_12396,N_10106,N_10085);
xnor U12397 (N_12397,N_8082,N_10847);
xnor U12398 (N_12398,N_8537,N_11871);
nor U12399 (N_12399,N_8149,N_11849);
xnor U12400 (N_12400,N_9616,N_11524);
and U12401 (N_12401,N_11889,N_8170);
and U12402 (N_12402,N_8508,N_8607);
or U12403 (N_12403,N_9141,N_9324);
nand U12404 (N_12404,N_8326,N_9536);
nand U12405 (N_12405,N_10757,N_8754);
and U12406 (N_12406,N_10065,N_10898);
nor U12407 (N_12407,N_9859,N_9507);
or U12408 (N_12408,N_11734,N_11555);
nor U12409 (N_12409,N_11415,N_10904);
nor U12410 (N_12410,N_9662,N_8579);
xnor U12411 (N_12411,N_10592,N_9564);
nand U12412 (N_12412,N_8876,N_11370);
or U12413 (N_12413,N_11962,N_8338);
nand U12414 (N_12414,N_11983,N_11143);
or U12415 (N_12415,N_9153,N_8941);
nand U12416 (N_12416,N_9954,N_11510);
or U12417 (N_12417,N_8256,N_11242);
or U12418 (N_12418,N_8443,N_10052);
nor U12419 (N_12419,N_10094,N_9571);
or U12420 (N_12420,N_8642,N_10993);
and U12421 (N_12421,N_9649,N_9463);
nand U12422 (N_12422,N_11004,N_8144);
nand U12423 (N_12423,N_8064,N_11557);
xor U12424 (N_12424,N_11921,N_11780);
and U12425 (N_12425,N_8503,N_10363);
and U12426 (N_12426,N_9003,N_9778);
and U12427 (N_12427,N_11018,N_8973);
xor U12428 (N_12428,N_11762,N_9687);
xor U12429 (N_12429,N_10230,N_9980);
or U12430 (N_12430,N_8652,N_11210);
and U12431 (N_12431,N_9838,N_11737);
nor U12432 (N_12432,N_10287,N_11700);
nand U12433 (N_12433,N_9323,N_9372);
or U12434 (N_12434,N_11693,N_10410);
nand U12435 (N_12435,N_9396,N_11681);
nor U12436 (N_12436,N_11498,N_10416);
nand U12437 (N_12437,N_9470,N_11874);
nand U12438 (N_12438,N_11005,N_10614);
or U12439 (N_12439,N_9551,N_8306);
xor U12440 (N_12440,N_8409,N_9727);
and U12441 (N_12441,N_9167,N_11032);
nor U12442 (N_12442,N_10531,N_10234);
nand U12443 (N_12443,N_10774,N_10882);
or U12444 (N_12444,N_11794,N_11372);
and U12445 (N_12445,N_9437,N_10928);
or U12446 (N_12446,N_9509,N_9197);
or U12447 (N_12447,N_11597,N_8169);
xnor U12448 (N_12448,N_10400,N_8128);
or U12449 (N_12449,N_8196,N_8806);
or U12450 (N_12450,N_9910,N_8724);
and U12451 (N_12451,N_11392,N_9593);
nor U12452 (N_12452,N_10918,N_9861);
and U12453 (N_12453,N_9000,N_8303);
nor U12454 (N_12454,N_8697,N_11157);
and U12455 (N_12455,N_10203,N_11997);
or U12456 (N_12456,N_11612,N_8058);
xnor U12457 (N_12457,N_9384,N_9561);
xor U12458 (N_12458,N_9400,N_8546);
or U12459 (N_12459,N_11316,N_8965);
nand U12460 (N_12460,N_10513,N_8478);
xnor U12461 (N_12461,N_11282,N_10902);
or U12462 (N_12462,N_9816,N_9313);
or U12463 (N_12463,N_11944,N_11699);
or U12464 (N_12464,N_9143,N_10408);
or U12465 (N_12465,N_9477,N_11055);
xnor U12466 (N_12466,N_10762,N_8092);
and U12467 (N_12467,N_10223,N_8247);
or U12468 (N_12468,N_8674,N_11929);
xor U12469 (N_12469,N_11069,N_9255);
and U12470 (N_12470,N_10352,N_9206);
or U12471 (N_12471,N_8921,N_10228);
or U12472 (N_12472,N_11306,N_9450);
and U12473 (N_12473,N_9156,N_9518);
nor U12474 (N_12474,N_9728,N_10504);
and U12475 (N_12475,N_11550,N_10903);
xnor U12476 (N_12476,N_9274,N_10155);
nor U12477 (N_12477,N_8728,N_8195);
nand U12478 (N_12478,N_9804,N_9736);
nor U12479 (N_12479,N_9339,N_9950);
and U12480 (N_12480,N_11713,N_8017);
nor U12481 (N_12481,N_8782,N_10767);
nor U12482 (N_12482,N_10383,N_9414);
nand U12483 (N_12483,N_11729,N_8744);
or U12484 (N_12484,N_8269,N_9357);
nor U12485 (N_12485,N_9941,N_10022);
or U12486 (N_12486,N_10424,N_9718);
or U12487 (N_12487,N_8158,N_11100);
and U12488 (N_12488,N_11767,N_9844);
nand U12489 (N_12489,N_11486,N_8635);
xor U12490 (N_12490,N_9667,N_8004);
or U12491 (N_12491,N_11895,N_11334);
and U12492 (N_12492,N_10332,N_11548);
nor U12493 (N_12493,N_10914,N_9284);
and U12494 (N_12494,N_10716,N_9368);
nand U12495 (N_12495,N_10414,N_8559);
nor U12496 (N_12496,N_8348,N_8742);
xor U12497 (N_12497,N_10704,N_10517);
and U12498 (N_12498,N_9483,N_11908);
xor U12499 (N_12499,N_11639,N_9514);
nor U12500 (N_12500,N_11515,N_8812);
and U12501 (N_12501,N_10734,N_10417);
and U12502 (N_12502,N_11395,N_11839);
or U12503 (N_12503,N_9026,N_8221);
or U12504 (N_12504,N_11679,N_9184);
nor U12505 (N_12505,N_8052,N_9083);
nor U12506 (N_12506,N_9779,N_8526);
or U12507 (N_12507,N_8244,N_8364);
nor U12508 (N_12508,N_10687,N_9702);
and U12509 (N_12509,N_9375,N_10187);
nand U12510 (N_12510,N_9138,N_10763);
or U12511 (N_12511,N_9103,N_11002);
nor U12512 (N_12512,N_9023,N_11992);
and U12513 (N_12513,N_10680,N_9426);
nand U12514 (N_12514,N_11056,N_10967);
xor U12515 (N_12515,N_9101,N_10285);
xor U12516 (N_12516,N_11743,N_8166);
nand U12517 (N_12517,N_9587,N_8966);
nor U12518 (N_12518,N_10674,N_8249);
xnor U12519 (N_12519,N_11608,N_9027);
or U12520 (N_12520,N_9090,N_10270);
nand U12521 (N_12521,N_11331,N_9380);
nor U12522 (N_12522,N_9927,N_10884);
nor U12523 (N_12523,N_9717,N_8922);
xnor U12524 (N_12524,N_11880,N_8430);
nand U12525 (N_12525,N_10173,N_11473);
xnor U12526 (N_12526,N_8357,N_9216);
xnor U12527 (N_12527,N_8512,N_8636);
nand U12528 (N_12528,N_11628,N_10871);
xnor U12529 (N_12529,N_8569,N_8703);
xor U12530 (N_12530,N_9532,N_9863);
nand U12531 (N_12531,N_11411,N_11867);
or U12532 (N_12532,N_9873,N_11434);
nor U12533 (N_12533,N_8873,N_8778);
xnor U12534 (N_12534,N_10862,N_8188);
nor U12535 (N_12535,N_9172,N_10535);
or U12536 (N_12536,N_8969,N_11781);
nand U12537 (N_12537,N_11607,N_11066);
nor U12538 (N_12538,N_8719,N_9349);
xor U12539 (N_12539,N_9606,N_9490);
xor U12540 (N_12540,N_8036,N_11352);
xor U12541 (N_12541,N_11716,N_10529);
xor U12542 (N_12542,N_10048,N_11046);
or U12543 (N_12543,N_8613,N_9192);
or U12544 (N_12544,N_11668,N_9902);
xor U12545 (N_12545,N_8000,N_9497);
nor U12546 (N_12546,N_8785,N_8959);
or U12547 (N_12547,N_10193,N_9343);
xor U12548 (N_12548,N_10235,N_11023);
nand U12549 (N_12549,N_9452,N_11868);
xnor U12550 (N_12550,N_10123,N_11501);
nor U12551 (N_12551,N_9458,N_10649);
or U12552 (N_12552,N_9706,N_10596);
nor U12553 (N_12553,N_10020,N_10926);
nor U12554 (N_12554,N_9637,N_10336);
xor U12555 (N_12555,N_8189,N_9517);
xnor U12556 (N_12556,N_10126,N_10314);
nor U12557 (N_12557,N_10209,N_11815);
and U12558 (N_12558,N_8997,N_8846);
xnor U12559 (N_12559,N_10275,N_11977);
nand U12560 (N_12560,N_8690,N_11030);
or U12561 (N_12561,N_8415,N_10585);
or U12562 (N_12562,N_8532,N_10372);
nand U12563 (N_12563,N_9524,N_9107);
nand U12564 (N_12564,N_11925,N_10450);
and U12565 (N_12565,N_9198,N_8771);
xor U12566 (N_12566,N_11586,N_9122);
nor U12567 (N_12567,N_10368,N_9168);
and U12568 (N_12568,N_8903,N_11326);
xor U12569 (N_12569,N_11741,N_10784);
xnor U12570 (N_12570,N_8774,N_8312);
and U12571 (N_12571,N_8182,N_11697);
nand U12572 (N_12572,N_9182,N_10453);
xor U12573 (N_12573,N_8228,N_10682);
xnor U12574 (N_12574,N_10353,N_9633);
and U12575 (N_12575,N_11174,N_11077);
xnor U12576 (N_12576,N_11090,N_8612);
xnor U12577 (N_12577,N_8954,N_11064);
nor U12578 (N_12578,N_11820,N_9824);
or U12579 (N_12579,N_9327,N_9781);
nand U12580 (N_12580,N_11226,N_8145);
or U12581 (N_12581,N_9675,N_8237);
or U12582 (N_12582,N_9664,N_9552);
xor U12583 (N_12583,N_10756,N_8935);
xnor U12584 (N_12584,N_8594,N_11049);
or U12585 (N_12585,N_8242,N_8704);
nand U12586 (N_12586,N_10170,N_11221);
xnor U12587 (N_12587,N_10711,N_10854);
and U12588 (N_12588,N_11796,N_10597);
and U12589 (N_12589,N_11850,N_8367);
and U12590 (N_12590,N_9010,N_8904);
or U12591 (N_12591,N_11688,N_9294);
nand U12592 (N_12592,N_11132,N_9353);
xor U12593 (N_12593,N_9992,N_9165);
and U12594 (N_12594,N_10224,N_8055);
nor U12595 (N_12595,N_10377,N_11297);
nor U12596 (N_12596,N_9290,N_10841);
and U12597 (N_12597,N_8867,N_10788);
xor U12598 (N_12598,N_10202,N_9309);
nand U12599 (N_12599,N_10200,N_11008);
and U12600 (N_12600,N_9482,N_8037);
nand U12601 (N_12601,N_8729,N_8378);
nand U12602 (N_12602,N_8585,N_11538);
nand U12603 (N_12603,N_11773,N_11290);
nor U12604 (N_12604,N_9434,N_10217);
and U12605 (N_12605,N_9752,N_8888);
xor U12606 (N_12606,N_11537,N_9693);
or U12607 (N_12607,N_8528,N_10607);
nor U12608 (N_12608,N_11930,N_11539);
or U12609 (N_12609,N_9094,N_11565);
nor U12610 (N_12610,N_11386,N_10881);
and U12611 (N_12611,N_8193,N_8371);
nor U12612 (N_12612,N_11399,N_9087);
nor U12613 (N_12613,N_11764,N_8425);
or U12614 (N_12614,N_11215,N_9903);
nand U12615 (N_12615,N_11890,N_8599);
and U12616 (N_12616,N_8236,N_9364);
nand U12617 (N_12617,N_11035,N_9746);
and U12618 (N_12618,N_8265,N_10938);
and U12619 (N_12619,N_8029,N_9457);
nand U12620 (N_12620,N_10487,N_10811);
and U12621 (N_12621,N_10072,N_10268);
nand U12622 (N_12622,N_9054,N_10679);
and U12623 (N_12623,N_10873,N_8445);
nand U12624 (N_12624,N_11048,N_10667);
or U12625 (N_12625,N_8611,N_9800);
or U12626 (N_12626,N_10828,N_10582);
xnor U12627 (N_12627,N_9334,N_11919);
or U12628 (N_12628,N_8264,N_11814);
and U12629 (N_12629,N_9241,N_9287);
nand U12630 (N_12630,N_11184,N_9105);
nand U12631 (N_12631,N_10093,N_10099);
and U12632 (N_12632,N_11663,N_9820);
and U12633 (N_12633,N_9937,N_8960);
nor U12634 (N_12634,N_10233,N_11592);
nor U12635 (N_12635,N_8660,N_10501);
xnor U12636 (N_12636,N_11785,N_10026);
nor U12637 (N_12637,N_9530,N_9865);
xor U12638 (N_12638,N_8644,N_10934);
nor U12639 (N_12639,N_8981,N_9239);
nand U12640 (N_12640,N_11134,N_10798);
nand U12641 (N_12641,N_11928,N_10522);
and U12642 (N_12642,N_8961,N_11115);
nor U12643 (N_12643,N_10720,N_10322);
or U12644 (N_12644,N_10069,N_11749);
nor U12645 (N_12645,N_9317,N_9537);
xnor U12646 (N_12646,N_9013,N_8254);
and U12647 (N_12647,N_10839,N_10262);
nor U12648 (N_12648,N_11472,N_9455);
and U12649 (N_12649,N_9767,N_8280);
xnor U12650 (N_12650,N_10817,N_10891);
xor U12651 (N_12651,N_10199,N_10747);
or U12652 (N_12652,N_8952,N_8289);
nand U12653 (N_12653,N_10848,N_8469);
nor U12654 (N_12654,N_8070,N_11324);
nand U12655 (N_12655,N_10855,N_10742);
or U12656 (N_12656,N_8160,N_8524);
nand U12657 (N_12657,N_11398,N_9131);
or U12658 (N_12658,N_11740,N_11453);
and U12659 (N_12659,N_9259,N_9526);
or U12660 (N_12660,N_8350,N_10082);
or U12661 (N_12661,N_8041,N_11179);
nor U12662 (N_12662,N_10736,N_10499);
xor U12663 (N_12663,N_9926,N_8962);
or U12664 (N_12664,N_8735,N_10722);
and U12665 (N_12665,N_8550,N_8046);
nand U12666 (N_12666,N_10394,N_11972);
and U12667 (N_12667,N_11238,N_11281);
or U12668 (N_12668,N_8102,N_8797);
xnor U12669 (N_12669,N_11732,N_9399);
or U12670 (N_12670,N_10952,N_11831);
and U12671 (N_12671,N_10087,N_9563);
nor U12672 (N_12672,N_10317,N_11436);
nand U12673 (N_12673,N_10247,N_11027);
xnor U12674 (N_12674,N_10050,N_11261);
or U12675 (N_12675,N_11365,N_11562);
nand U12676 (N_12676,N_9175,N_9268);
nor U12677 (N_12677,N_10808,N_9757);
or U12678 (N_12678,N_11413,N_11367);
or U12679 (N_12679,N_9033,N_9655);
or U12680 (N_12680,N_11382,N_11926);
nand U12681 (N_12681,N_11637,N_9200);
and U12682 (N_12682,N_10962,N_11988);
nand U12683 (N_12683,N_11958,N_10617);
xor U12684 (N_12684,N_8451,N_9246);
or U12685 (N_12685,N_11358,N_8515);
xnor U12686 (N_12686,N_11655,N_11795);
nor U12687 (N_12687,N_10141,N_9965);
or U12688 (N_12688,N_8325,N_11484);
nand U12689 (N_12689,N_9449,N_8944);
and U12690 (N_12690,N_9747,N_11797);
nor U12691 (N_12691,N_9516,N_11390);
and U12692 (N_12692,N_10696,N_8625);
nand U12693 (N_12693,N_10943,N_10030);
and U12694 (N_12694,N_8743,N_8309);
nor U12695 (N_12695,N_9831,N_10821);
nor U12696 (N_12696,N_11219,N_9697);
xnor U12697 (N_12697,N_11275,N_8539);
or U12698 (N_12698,N_9240,N_11396);
nor U12699 (N_12699,N_8164,N_9974);
and U12700 (N_12700,N_10009,N_11602);
and U12701 (N_12701,N_9163,N_9772);
or U12702 (N_12702,N_10345,N_11747);
nor U12703 (N_12703,N_10292,N_10953);
xnor U12704 (N_12704,N_10439,N_8859);
nor U12705 (N_12705,N_8712,N_11126);
nor U12706 (N_12706,N_10843,N_11204);
and U12707 (N_12707,N_11068,N_9109);
or U12708 (N_12708,N_9036,N_10536);
nor U12709 (N_12709,N_8420,N_8779);
nor U12710 (N_12710,N_11235,N_9351);
nand U12711 (N_12711,N_11402,N_11477);
nand U12712 (N_12712,N_8809,N_9123);
nor U12713 (N_12713,N_11579,N_8760);
nand U12714 (N_12714,N_10772,N_11711);
nor U12715 (N_12715,N_8328,N_8491);
and U12716 (N_12716,N_9654,N_9971);
and U12717 (N_12717,N_11945,N_11188);
nor U12718 (N_12718,N_10787,N_11404);
xnor U12719 (N_12719,N_11432,N_10701);
or U12720 (N_12720,N_11474,N_8548);
nor U12721 (N_12721,N_9186,N_10669);
or U12722 (N_12722,N_11322,N_9581);
nor U12723 (N_12723,N_8699,N_9515);
or U12724 (N_12724,N_9813,N_11303);
or U12725 (N_12725,N_8347,N_11523);
nor U12726 (N_12726,N_8899,N_11410);
xor U12727 (N_12727,N_10360,N_11086);
xnor U12728 (N_12728,N_11491,N_8243);
nor U12729 (N_12729,N_8207,N_9196);
nand U12730 (N_12730,N_9075,N_10590);
nand U12731 (N_12731,N_10668,N_8807);
nor U12732 (N_12732,N_11345,N_10958);
nand U12733 (N_12733,N_11709,N_11001);
and U12734 (N_12734,N_9628,N_10115);
xor U12735 (N_12735,N_11576,N_9972);
or U12736 (N_12736,N_10653,N_9510);
or U12737 (N_12737,N_11556,N_8315);
nand U12738 (N_12738,N_9858,N_9986);
or U12739 (N_12739,N_11606,N_10746);
and U12740 (N_12740,N_8136,N_11025);
and U12741 (N_12741,N_10423,N_9599);
xor U12742 (N_12742,N_9793,N_9982);
nand U12743 (N_12743,N_10307,N_9264);
xnor U12744 (N_12744,N_11652,N_8141);
nand U12745 (N_12745,N_8101,N_11313);
nand U12746 (N_12746,N_8987,N_11257);
or U12747 (N_12747,N_10699,N_10670);
or U12748 (N_12748,N_10341,N_9207);
or U12749 (N_12749,N_11960,N_11920);
or U12750 (N_12750,N_11130,N_10745);
and U12751 (N_12751,N_8633,N_11340);
and U12752 (N_12752,N_8829,N_9049);
nor U12753 (N_12753,N_11578,N_11287);
nor U12754 (N_12754,N_8974,N_9983);
nand U12755 (N_12755,N_10459,N_11429);
or U12756 (N_12756,N_9215,N_11822);
xnor U12757 (N_12757,N_9362,N_10016);
or U12758 (N_12758,N_9250,N_9930);
nor U12759 (N_12759,N_11967,N_10623);
nand U12760 (N_12760,N_9851,N_10460);
or U12761 (N_12761,N_10625,N_10588);
xor U12762 (N_12762,N_8596,N_11554);
xor U12763 (N_12763,N_8505,N_8200);
and U12764 (N_12764,N_8977,N_9069);
nor U12765 (N_12765,N_8452,N_11509);
or U12766 (N_12766,N_9097,N_8400);
or U12767 (N_12767,N_8023,N_9428);
nor U12768 (N_12768,N_10520,N_11514);
and U12769 (N_12769,N_10730,N_9193);
or U12770 (N_12770,N_11819,N_10182);
or U12771 (N_12771,N_11394,N_11376);
and U12772 (N_12772,N_10578,N_11407);
xor U12773 (N_12773,N_8925,N_9204);
nor U12774 (N_12774,N_8106,N_9433);
nand U12775 (N_12775,N_9314,N_8765);
nor U12776 (N_12776,N_11651,N_10162);
xor U12777 (N_12777,N_9005,N_8302);
or U12778 (N_12778,N_10602,N_9119);
nand U12779 (N_12779,N_11746,N_9609);
and U12780 (N_12780,N_9817,N_11338);
nand U12781 (N_12781,N_10156,N_9957);
nand U12782 (N_12782,N_10702,N_8336);
nor U12783 (N_12783,N_11425,N_9840);
and U12784 (N_12784,N_10466,N_8412);
and U12785 (N_12785,N_8084,N_8218);
and U12786 (N_12786,N_11201,N_8858);
or U12787 (N_12787,N_9254,N_8386);
nor U12788 (N_12788,N_9258,N_11563);
nand U12789 (N_12789,N_9523,N_8860);
nand U12790 (N_12790,N_8615,N_11074);
or U12791 (N_12791,N_11205,N_9896);
xnor U12792 (N_12792,N_10880,N_10384);
nand U12793 (N_12793,N_8010,N_11883);
nand U12794 (N_12794,N_10963,N_8180);
or U12795 (N_12795,N_10054,N_8570);
nand U12796 (N_12796,N_11039,N_8295);
nand U12797 (N_12797,N_9769,N_11119);
xor U12798 (N_12798,N_11339,N_8150);
nand U12799 (N_12799,N_8759,N_11485);
xor U12800 (N_12800,N_9681,N_10758);
nand U12801 (N_12801,N_10271,N_10885);
or U12802 (N_12802,N_8542,N_11745);
and U12803 (N_12803,N_8026,N_8219);
nor U12804 (N_12804,N_10385,N_8844);
xor U12805 (N_12805,N_10820,N_8234);
xnor U12806 (N_12806,N_8284,N_9945);
xor U12807 (N_12807,N_10801,N_10601);
xnor U12808 (N_12808,N_11469,N_8135);
nand U12809 (N_12809,N_11191,N_11742);
nand U12810 (N_12810,N_10374,N_9643);
xnor U12811 (N_12811,N_10083,N_8700);
and U12812 (N_12812,N_8614,N_10626);
nand U12813 (N_12813,N_11718,N_8129);
or U12814 (N_12814,N_9642,N_8518);
or U12815 (N_12815,N_9297,N_11891);
xor U12816 (N_12816,N_10429,N_11733);
or U12817 (N_12817,N_9498,N_9676);
and U12818 (N_12818,N_8556,N_8259);
xor U12819 (N_12819,N_10766,N_9578);
nor U12820 (N_12820,N_11937,N_10389);
and U12821 (N_12821,N_11263,N_11938);
and U12822 (N_12822,N_9238,N_11164);
nand U12823 (N_12823,N_11167,N_11271);
or U12824 (N_12824,N_11551,N_11696);
and U12825 (N_12825,N_10743,N_9074);
and U12826 (N_12826,N_9062,N_9333);
nand U12827 (N_12827,N_8916,N_8458);
xor U12828 (N_12828,N_11103,N_10273);
nor U12829 (N_12829,N_10894,N_11851);
nand U12830 (N_12830,N_10737,N_11715);
xor U12831 (N_12831,N_10479,N_9505);
and U12832 (N_12832,N_9568,N_10014);
or U12833 (N_12833,N_11104,N_9944);
nor U12834 (N_12834,N_10248,N_9095);
and U12835 (N_12835,N_10011,N_8848);
xnor U12836 (N_12836,N_10232,N_11197);
xor U12837 (N_12837,N_8079,N_8630);
or U12838 (N_12838,N_10754,N_8808);
nand U12839 (N_12839,N_8427,N_10648);
xnor U12840 (N_12840,N_9442,N_9485);
or U12841 (N_12841,N_9823,N_9550);
or U12842 (N_12842,N_10293,N_10296);
nand U12843 (N_12843,N_10889,N_11912);
xnor U12844 (N_12844,N_9481,N_11755);
xor U12845 (N_12845,N_10778,N_8467);
and U12846 (N_12846,N_11307,N_8619);
nor U12847 (N_12847,N_9719,N_10198);
or U12848 (N_12848,N_8939,N_9161);
or U12849 (N_12849,N_11529,N_8525);
xnor U12850 (N_12850,N_9572,N_11975);
and U12851 (N_12851,N_11098,N_10008);
xor U12852 (N_12852,N_8065,N_11526);
nand U12853 (N_12853,N_11384,N_11759);
xor U12854 (N_12854,N_10309,N_9751);
or U12855 (N_12855,N_10272,N_9811);
xnor U12856 (N_12856,N_8227,N_9421);
nand U12857 (N_12857,N_9177,N_8183);
or U12858 (N_12858,N_11280,N_8851);
and U12859 (N_12859,N_9703,N_10313);
and U12860 (N_12860,N_11512,N_10562);
or U12861 (N_12861,N_8279,N_10944);
xor U12862 (N_12862,N_9038,N_8986);
nor U12863 (N_12863,N_10600,N_8931);
and U12864 (N_12864,N_10988,N_10652);
or U12865 (N_12865,N_10104,N_8459);
and U12866 (N_12866,N_10432,N_11721);
or U12867 (N_12867,N_9230,N_10780);
nor U12868 (N_12868,N_8494,N_10181);
or U12869 (N_12869,N_8824,N_10834);
nor U12870 (N_12870,N_10927,N_9600);
xor U12871 (N_12871,N_8389,N_10269);
or U12872 (N_12872,N_11333,N_10066);
nand U12873 (N_12873,N_9958,N_9569);
xor U12874 (N_12874,N_8475,N_11249);
nand U12875 (N_12875,N_11799,N_9019);
nand U12876 (N_12876,N_9350,N_11113);
nand U12877 (N_12877,N_9410,N_8318);
and U12878 (N_12878,N_11674,N_10045);
or U12879 (N_12879,N_11181,N_11769);
and U12880 (N_12880,N_8291,N_9116);
and U12881 (N_12881,N_9488,N_11752);
nand U12882 (N_12882,N_11082,N_9443);
and U12883 (N_12883,N_10397,N_10098);
nor U12884 (N_12884,N_9801,N_10646);
xor U12885 (N_12885,N_11128,N_9721);
and U12886 (N_12886,N_8311,N_11932);
nand U12887 (N_12887,N_8813,N_8621);
nor U12888 (N_12888,N_8563,N_10062);
xor U12889 (N_12889,N_8286,N_8125);
and U12890 (N_12890,N_10654,N_9909);
nor U12891 (N_12891,N_11645,N_11033);
nor U12892 (N_12892,N_10781,N_8672);
nand U12893 (N_12893,N_9806,N_8216);
and U12894 (N_12894,N_8918,N_11465);
xor U12895 (N_12895,N_8121,N_10080);
and U12896 (N_12896,N_10446,N_8578);
and U12897 (N_12897,N_10642,N_10282);
nand U12898 (N_12898,N_11479,N_8397);
or U12899 (N_12899,N_11168,N_8936);
xnor U12900 (N_12900,N_11011,N_9256);
nor U12901 (N_12901,N_8781,N_8855);
nor U12902 (N_12902,N_10548,N_9933);
nand U12903 (N_12903,N_9522,N_9092);
nor U12904 (N_12904,N_8372,N_11790);
or U12905 (N_12905,N_11232,N_8222);
nor U12906 (N_12906,N_11941,N_8748);
nand U12907 (N_12907,N_10759,N_11570);
xnor U12908 (N_12908,N_9278,N_10311);
nand U12909 (N_12909,N_11470,N_11543);
and U12910 (N_12910,N_8739,N_10515);
or U12911 (N_12911,N_9848,N_9533);
or U12912 (N_12912,N_9080,N_9699);
nor U12913 (N_12913,N_11658,N_10470);
and U12914 (N_12914,N_10819,N_8011);
xor U12915 (N_12915,N_8281,N_11493);
nor U12916 (N_12916,N_11435,N_9756);
or U12917 (N_12917,N_11876,N_11582);
nand U12918 (N_12918,N_10025,N_10673);
nor U12919 (N_12919,N_11439,N_8346);
nor U12920 (N_12920,N_9385,N_11327);
nor U12921 (N_12921,N_11065,N_11573);
nand U12922 (N_12922,N_11642,N_9975);
xor U12923 (N_12923,N_9341,N_11260);
and U12924 (N_12924,N_11558,N_11272);
nor U12925 (N_12925,N_9389,N_11459);
nand U12926 (N_12926,N_11239,N_11951);
xnor U12927 (N_12927,N_8993,N_9242);
nor U12928 (N_12928,N_11467,N_11258);
xnor U12929 (N_12929,N_9940,N_9951);
xnor U12930 (N_12930,N_11489,N_10318);
or U12931 (N_12931,N_10076,N_10621);
nor U12932 (N_12932,N_8945,N_8566);
or U12933 (N_12933,N_11897,N_10688);
or U12934 (N_12934,N_9022,N_9814);
nor U12935 (N_12935,N_8363,N_11229);
nand U12936 (N_12936,N_11984,N_11317);
and U12937 (N_12937,N_9932,N_8984);
or U12938 (N_12938,N_10010,N_11482);
nor U12939 (N_12939,N_9325,N_9529);
or U12940 (N_12940,N_9199,N_11114);
or U12941 (N_12941,N_10980,N_10036);
nand U12942 (N_12942,N_11569,N_11231);
or U12943 (N_12943,N_9770,N_11125);
or U12944 (N_12944,N_9306,N_11855);
nand U12945 (N_12945,N_10255,N_11541);
nor U12946 (N_12946,N_9712,N_11643);
nor U12947 (N_12947,N_8307,N_10609);
nand U12948 (N_12948,N_8086,N_8449);
xor U12949 (N_12949,N_8317,N_8882);
and U12950 (N_12950,N_9352,N_10857);
nor U12951 (N_12951,N_11038,N_10864);
nor U12952 (N_12952,N_11784,N_9233);
or U12953 (N_12953,N_10184,N_10692);
and U12954 (N_12954,N_10560,N_9081);
nor U12955 (N_12955,N_8761,N_11349);
nand U12956 (N_12956,N_9977,N_11147);
xor U12957 (N_12957,N_10583,N_8698);
nor U12958 (N_12958,N_8080,N_9283);
nor U12959 (N_12959,N_10895,N_10047);
and U12960 (N_12960,N_11650,N_10120);
xor U12961 (N_12961,N_9627,N_11246);
nand U12962 (N_12962,N_10859,N_11522);
or U12963 (N_12963,N_8667,N_8131);
or U12964 (N_12964,N_10207,N_10631);
and U12965 (N_12965,N_10134,N_10298);
or U12966 (N_12966,N_10921,N_8177);
xnor U12967 (N_12967,N_11854,N_11422);
and U12968 (N_12968,N_8507,N_9289);
and U12969 (N_12969,N_10561,N_10330);
nand U12970 (N_12970,N_11487,N_10081);
nor U12971 (N_12971,N_8725,N_8720);
xnor U12972 (N_12972,N_10252,N_8408);
nor U12973 (N_12973,N_8834,N_8305);
nand U12974 (N_12974,N_8866,N_10148);
xnor U12975 (N_12975,N_8134,N_9713);
xnor U12976 (N_12976,N_8581,N_9666);
xor U12977 (N_12977,N_9780,N_11671);
xnor U12978 (N_12978,N_8886,N_10725);
and U12979 (N_12979,N_9008,N_11705);
xor U12980 (N_12980,N_8250,N_8087);
xor U12981 (N_12981,N_8293,N_9994);
nand U12982 (N_12982,N_8996,N_11350);
and U12983 (N_12983,N_11253,N_10406);
and U12984 (N_12984,N_9596,N_9900);
and U12985 (N_12985,N_11633,N_8175);
nand U12986 (N_12986,N_9614,N_8560);
and U12987 (N_12987,N_10327,N_9411);
nand U12988 (N_12988,N_11379,N_9468);
nor U12989 (N_12989,N_9671,N_10480);
nor U12990 (N_12990,N_9624,N_11829);
or U12991 (N_12991,N_11717,N_8335);
nand U12992 (N_12992,N_8345,N_8517);
nor U12993 (N_12993,N_11220,N_9640);
nand U12994 (N_12994,N_10244,N_10319);
nand U12995 (N_12995,N_11953,N_9137);
or U12996 (N_12996,N_10102,N_10955);
or U12997 (N_12997,N_9454,N_10657);
and U12998 (N_12998,N_10683,N_8314);
nor U12999 (N_12999,N_10393,N_9479);
or U13000 (N_13000,N_8276,N_11159);
nor U13001 (N_13001,N_10116,N_11108);
or U13002 (N_13002,N_9335,N_11445);
or U13003 (N_13003,N_9279,N_8802);
xor U13004 (N_13004,N_8887,N_10907);
xnor U13005 (N_13005,N_10018,N_9050);
nor U13006 (N_13006,N_9680,N_11305);
xor U13007 (N_13007,N_10294,N_10634);
and U13008 (N_13008,N_9394,N_9739);
and U13009 (N_13009,N_8976,N_11206);
nor U13010 (N_13010,N_8805,N_10976);
nor U13011 (N_13011,N_10681,N_9726);
nor U13012 (N_13012,N_11319,N_9245);
and U13013 (N_13013,N_11180,N_8776);
xnor U13014 (N_13014,N_11600,N_8626);
or U13015 (N_13015,N_10825,N_10733);
and U13016 (N_13016,N_8091,N_8203);
nand U13017 (N_13017,N_8407,N_8255);
xnor U13018 (N_13018,N_8251,N_8901);
xor U13019 (N_13019,N_9585,N_10939);
nand U13020 (N_13020,N_9445,N_8649);
nor U13021 (N_13021,N_11614,N_8490);
and U13022 (N_13022,N_10236,N_10813);
xnor U13023 (N_13023,N_8837,N_10845);
nor U13024 (N_13024,N_10402,N_9286);
nor U13025 (N_13025,N_9525,N_11031);
nand U13026 (N_13026,N_10949,N_8320);
nand U13027 (N_13027,N_9300,N_8598);
xnor U13028 (N_13028,N_8561,N_10651);
nand U13029 (N_13029,N_11006,N_10610);
nor U13030 (N_13030,N_9104,N_8905);
and U13031 (N_13031,N_9500,N_9051);
or U13032 (N_13032,N_11135,N_9248);
nand U13033 (N_13033,N_8021,N_11835);
and U13034 (N_13034,N_9673,N_11809);
xor U13035 (N_13035,N_10916,N_11026);
nand U13036 (N_13036,N_10493,N_8705);
or U13037 (N_13037,N_9622,N_10053);
or U13038 (N_13038,N_10537,N_8133);
nor U13039 (N_13039,N_9251,N_9296);
nand U13040 (N_13040,N_11596,N_10231);
nor U13041 (N_13041,N_11886,N_11933);
nor U13042 (N_13042,N_11866,N_10344);
or U13043 (N_13043,N_10122,N_10534);
and U13044 (N_13044,N_11092,N_9914);
or U13045 (N_13045,N_8201,N_8429);
or U13046 (N_13046,N_9880,N_11660);
and U13047 (N_13047,N_8075,N_10105);
and U13048 (N_13048,N_11682,N_9603);
xor U13049 (N_13049,N_11724,N_9506);
nor U13050 (N_13050,N_11369,N_10516);
xnor U13051 (N_13051,N_10945,N_9473);
nand U13052 (N_13052,N_9595,N_8339);
or U13053 (N_13053,N_10721,N_10822);
or U13054 (N_13054,N_10557,N_10301);
and U13055 (N_13055,N_10693,N_10846);
xor U13056 (N_13056,N_9874,N_9876);
nand U13057 (N_13057,N_11687,N_9864);
xor U13058 (N_13058,N_8730,N_9812);
nand U13059 (N_13059,N_10691,N_11315);
xnor U13060 (N_13060,N_11444,N_8536);
and U13061 (N_13061,N_9942,N_10748);
nand U13062 (N_13062,N_11216,N_11186);
nor U13063 (N_13063,N_11841,N_9832);
and U13064 (N_13064,N_11171,N_9185);
xnor U13065 (N_13065,N_9636,N_8127);
nor U13066 (N_13066,N_9878,N_10381);
xnor U13067 (N_13067,N_10444,N_11588);
xor U13068 (N_13068,N_8260,N_8877);
or U13069 (N_13069,N_9218,N_9583);
xnor U13070 (N_13070,N_10242,N_8050);
nand U13071 (N_13071,N_8602,N_9174);
and U13072 (N_13072,N_10186,N_8814);
or U13073 (N_13073,N_11187,N_11476);
nor U13074 (N_13074,N_9678,N_9430);
or U13075 (N_13075,N_11575,N_9461);
or U13076 (N_13076,N_8912,N_10086);
and U13077 (N_13077,N_8111,N_10678);
xnor U13078 (N_13078,N_11615,N_11133);
nand U13079 (N_13079,N_11223,N_11378);
or U13080 (N_13080,N_11892,N_9298);
and U13081 (N_13081,N_8297,N_9438);
nor U13082 (N_13082,N_9698,N_10732);
nor U13083 (N_13083,N_10966,N_8889);
or U13084 (N_13084,N_11085,N_9070);
nor U13085 (N_13085,N_11777,N_11726);
nand U13086 (N_13086,N_8775,N_8786);
or U13087 (N_13087,N_10521,N_8990);
or U13088 (N_13088,N_9792,N_8076);
xor U13089 (N_13089,N_8801,N_9594);
nor U13090 (N_13090,N_11154,N_11355);
nor U13091 (N_13091,N_9785,N_11599);
or U13092 (N_13092,N_11838,N_11291);
xnor U13093 (N_13093,N_11739,N_11203);
nor U13094 (N_13094,N_8789,N_9358);
xnor U13095 (N_13095,N_9574,N_11141);
and U13096 (N_13096,N_8662,N_11447);
nor U13097 (N_13097,N_8217,N_9128);
or U13098 (N_13098,N_10125,N_9035);
and U13099 (N_13099,N_10740,N_11813);
or U13100 (N_13100,N_8343,N_11520);
xnor U13101 (N_13101,N_11408,N_9630);
nor U13102 (N_13102,N_8545,N_9431);
nand U13103 (N_13103,N_11198,N_10288);
nor U13104 (N_13104,N_8391,N_10666);
nor U13105 (N_13105,N_8081,N_11034);
nor U13106 (N_13106,N_9077,N_9271);
or U13107 (N_13107,N_8909,N_8304);
nor U13108 (N_13108,N_9744,N_11051);
or U13109 (N_13109,N_11840,N_11457);
nand U13110 (N_13110,N_11196,N_10321);
or U13111 (N_13111,N_11455,N_9441);
nor U13112 (N_13112,N_11800,N_8610);
nand U13113 (N_13113,N_10593,N_9057);
and U13114 (N_13114,N_10664,N_10291);
xor U13115 (N_13115,N_10887,N_10490);
nand U13116 (N_13116,N_8862,N_9588);
and U13117 (N_13117,N_11416,N_10260);
and U13118 (N_13118,N_11234,N_9617);
nor U13119 (N_13119,N_11657,N_8007);
xnor U13120 (N_13120,N_11243,N_11860);
nor U13121 (N_13121,N_11959,N_8358);
xor U13122 (N_13122,N_10744,N_8043);
nor U13123 (N_13123,N_8753,N_10403);
nand U13124 (N_13124,N_8691,N_9887);
or U13125 (N_13125,N_8727,N_8661);
nand U13126 (N_13126,N_8717,N_9920);
xnor U13127 (N_13127,N_9894,N_11961);
nor U13128 (N_13128,N_10629,N_9374);
and U13129 (N_13129,N_9835,N_9732);
nor U13130 (N_13130,N_11730,N_9195);
and U13131 (N_13131,N_10628,N_8995);
or U13132 (N_13132,N_8514,N_11763);
nor U13133 (N_13133,N_11561,N_11712);
or U13134 (N_13134,N_8571,N_8155);
nor U13135 (N_13135,N_9208,N_10179);
and U13136 (N_13136,N_10984,N_11872);
nor U13137 (N_13137,N_10147,N_8198);
and U13138 (N_13138,N_10300,N_8151);
nand U13139 (N_13139,N_11916,N_10071);
xnor U13140 (N_13140,N_9535,N_11110);
nand U13141 (N_13141,N_8768,N_8375);
or U13142 (N_13142,N_10823,N_11792);
and U13143 (N_13143,N_10239,N_9818);
or U13144 (N_13144,N_11949,N_8538);
nand U13145 (N_13145,N_9650,N_10724);
nand U13146 (N_13146,N_8821,N_10969);
nand U13147 (N_13147,N_11604,N_9962);
or U13148 (N_13148,N_8097,N_10426);
or U13149 (N_13149,N_11250,N_10278);
xor U13150 (N_13150,N_9612,N_9149);
nand U13151 (N_13151,N_11433,N_10860);
xnor U13152 (N_13152,N_8575,N_11636);
and U13153 (N_13153,N_10340,N_11015);
and U13154 (N_13154,N_9841,N_11029);
xnor U13155 (N_13155,N_9459,N_10947);
xnor U13156 (N_13156,N_11175,N_11344);
and U13157 (N_13157,N_8631,N_9646);
or U13158 (N_13158,N_10599,N_9212);
or U13159 (N_13159,N_11189,N_8384);
xnor U13160 (N_13160,N_11426,N_8694);
nand U13161 (N_13161,N_8277,N_8506);
nor U13162 (N_13162,N_10974,N_9883);
or U13163 (N_13163,N_10569,N_8069);
xor U13164 (N_13164,N_9231,N_9597);
and U13165 (N_13165,N_9342,N_8910);
or U13166 (N_13166,N_9916,N_8003);
xnor U13167 (N_13167,N_9635,N_8643);
xor U13168 (N_13168,N_8632,N_10306);
xor U13169 (N_13169,N_9765,N_9504);
or U13170 (N_13170,N_11172,N_8618);
and U13171 (N_13171,N_10553,N_8462);
xnor U13172 (N_13172,N_11775,N_9417);
and U13173 (N_13173,N_11995,N_8552);
and U13174 (N_13174,N_11989,N_9528);
or U13175 (N_13175,N_11149,N_11686);
and U13176 (N_13176,N_8756,N_8906);
and U13177 (N_13177,N_11400,N_8387);
nand U13178 (N_13178,N_8920,N_10485);
and U13179 (N_13179,N_10929,N_11985);
xnor U13180 (N_13180,N_11041,N_10770);
nor U13181 (N_13181,N_11495,N_11942);
nand U13182 (N_13182,N_11751,N_9347);
or U13183 (N_13183,N_9639,N_11504);
or U13184 (N_13184,N_11571,N_11499);
nor U13185 (N_13185,N_9978,N_10526);
or U13186 (N_13186,N_10936,N_11072);
or U13187 (N_13187,N_8191,N_11406);
nand U13188 (N_13188,N_8850,N_8687);
xor U13189 (N_13189,N_9173,N_8968);
xnor U13190 (N_13190,N_10356,N_11214);
nand U13191 (N_13191,N_8161,N_9096);
or U13192 (N_13192,N_10613,N_8331);
xor U13193 (N_13193,N_11852,N_8943);
and U13194 (N_13194,N_10961,N_10900);
or U13195 (N_13195,N_10422,N_11099);
nand U13196 (N_13196,N_10542,N_8955);
xnor U13197 (N_13197,N_11948,N_10451);
nor U13198 (N_13198,N_8116,N_9205);
nand U13199 (N_13199,N_10488,N_11503);
nand U13200 (N_13200,N_9694,N_8365);
nor U13201 (N_13201,N_10335,N_11904);
nor U13202 (N_13202,N_9527,N_11405);
nand U13203 (N_13203,N_11062,N_11964);
nor U13204 (N_13204,N_9682,N_10530);
and U13205 (N_13205,N_10695,N_11299);
nor U13206 (N_13206,N_9145,N_9130);
xnor U13207 (N_13207,N_8398,N_8732);
or U13208 (N_13208,N_11268,N_11106);
xnor U13209 (N_13209,N_9566,N_9534);
nand U13210 (N_13210,N_10205,N_9791);
or U13211 (N_13211,N_10591,N_8849);
and U13212 (N_13212,N_10149,N_9653);
or U13213 (N_13213,N_9539,N_9724);
xnor U13214 (N_13214,N_8590,N_9356);
nor U13215 (N_13215,N_11304,N_9956);
and U13216 (N_13216,N_11166,N_11683);
and U13217 (N_13217,N_11862,N_9419);
nand U13218 (N_13218,N_10568,N_11605);
nor U13219 (N_13219,N_8215,N_8822);
xor U13220 (N_13220,N_11691,N_10194);
or U13221 (N_13221,N_10127,N_10070);
and U13222 (N_13222,N_11437,N_9674);
nand U13223 (N_13223,N_9072,N_10339);
xor U13224 (N_13224,N_10932,N_8971);
xnor U13225 (N_13225,N_11309,N_10136);
nor U13226 (N_13226,N_10040,N_9222);
nand U13227 (N_13227,N_11248,N_11638);
or U13228 (N_13228,N_9567,N_9990);
and U13229 (N_13229,N_11931,N_9330);
and U13230 (N_13230,N_11312,N_9651);
nor U13231 (N_13231,N_9467,N_11265);
or U13232 (N_13232,N_8584,N_8044);
nand U13233 (N_13233,N_10111,N_8780);
xnor U13234 (N_13234,N_10985,N_10107);
nand U13235 (N_13235,N_8310,N_11227);
nand U13236 (N_13236,N_8978,N_10044);
nor U13237 (N_13237,N_11821,N_11905);
xnor U13238 (N_13238,N_8479,N_10710);
nor U13239 (N_13239,N_8261,N_9707);
xnor U13240 (N_13240,N_11073,N_8063);
xnor U13241 (N_13241,N_9100,N_11121);
or U13242 (N_13242,N_9969,N_11744);
and U13243 (N_13243,N_8991,N_8564);
nor U13244 (N_13244,N_8622,N_11247);
nor U13245 (N_13245,N_10055,N_8187);
nand U13246 (N_13246,N_11084,N_10800);
or U13247 (N_13247,N_10964,N_10551);
xnor U13248 (N_13248,N_8750,N_8418);
nand U13249 (N_13249,N_11286,N_11200);
xor U13250 (N_13250,N_10635,N_11360);
nand U13251 (N_13251,N_8167,N_8763);
nand U13252 (N_13252,N_9388,N_9888);
and U13253 (N_13253,N_9344,N_11952);
nand U13254 (N_13254,N_9085,N_10500);
nand U13255 (N_13255,N_11288,N_9460);
and U13256 (N_13256,N_10723,N_11818);
xnor U13257 (N_13257,N_10510,N_10002);
or U13258 (N_13258,N_8804,N_9573);
or U13259 (N_13259,N_10152,N_8073);
or U13260 (N_13260,N_10337,N_10092);
nor U13261 (N_13261,N_10708,N_9321);
xnor U13262 (N_13262,N_9115,N_9140);
xnor U13263 (N_13263,N_9355,N_11677);
nand U13264 (N_13264,N_9007,N_9764);
or U13265 (N_13265,N_11292,N_8231);
xnor U13266 (N_13266,N_10970,N_8558);
or U13267 (N_13267,N_9862,N_8843);
nor U13268 (N_13268,N_10057,N_9418);
nand U13269 (N_13269,N_10525,N_10799);
xor U13270 (N_13270,N_11383,N_10838);
xnor U13271 (N_13271,N_10304,N_10549);
or U13272 (N_13272,N_9709,N_8645);
nor U13273 (N_13273,N_8210,N_11618);
or U13274 (N_13274,N_11464,N_11505);
nor U13275 (N_13275,N_10206,N_10935);
or U13276 (N_13276,N_11518,N_8522);
nand U13277 (N_13277,N_10779,N_10034);
xnor U13278 (N_13278,N_10835,N_10803);
xnor U13279 (N_13279,N_9827,N_10586);
and U13280 (N_13280,N_11758,N_11552);
nor U13281 (N_13281,N_8060,N_11182);
and U13282 (N_13282,N_10249,N_8767);
xnor U13283 (N_13283,N_8544,N_8722);
nor U13284 (N_13284,N_9589,N_10420);
or U13285 (N_13285,N_10445,N_9710);
nand U13286 (N_13286,N_10067,N_10254);
and U13287 (N_13287,N_8355,N_9243);
nand U13288 (N_13288,N_11328,N_8366);
nor U13289 (N_13289,N_10246,N_10264);
and U13290 (N_13290,N_8871,N_11846);
or U13291 (N_13291,N_9340,N_9893);
xor U13292 (N_13292,N_11956,N_8232);
nand U13293 (N_13293,N_10021,N_9720);
xnor U13294 (N_13294,N_10765,N_8501);
or U13295 (N_13295,N_10442,N_8671);
nor U13296 (N_13296,N_11782,N_10833);
and U13297 (N_13297,N_11348,N_9512);
xor U13298 (N_13298,N_8045,N_11302);
and U13299 (N_13299,N_9166,N_11124);
nor U13300 (N_13300,N_9924,N_8530);
nor U13301 (N_13301,N_8061,N_10815);
nor U13302 (N_13302,N_11864,N_10827);
nand U13303 (N_13303,N_8500,N_10333);
nand U13304 (N_13304,N_9560,N_10443);
nor U13305 (N_13305,N_11009,N_10942);
or U13306 (N_13306,N_8926,N_10486);
or U13307 (N_13307,N_11356,N_11519);
nor U13308 (N_13308,N_9601,N_9282);
nand U13309 (N_13309,N_10427,N_11183);
and U13310 (N_13310,N_10919,N_9857);
nor U13311 (N_13311,N_8956,N_10760);
xor U13312 (N_13312,N_9187,N_9393);
and U13313 (N_13313,N_10981,N_10004);
nor U13314 (N_13314,N_10773,N_10168);
or U13315 (N_13315,N_8301,N_9018);
nor U13316 (N_13316,N_11451,N_9830);
nor U13317 (N_13317,N_10279,N_9786);
nand U13318 (N_13318,N_8246,N_8153);
and U13319 (N_13319,N_8681,N_9332);
nor U13320 (N_13320,N_8523,N_8112);
nand U13321 (N_13321,N_8245,N_11533);
and U13322 (N_13322,N_11641,N_9379);
or U13323 (N_13323,N_10139,N_8983);
nand U13324 (N_13324,N_9292,N_8379);
and U13325 (N_13325,N_9139,N_8392);
and U13326 (N_13326,N_11568,N_10703);
xnor U13327 (N_13327,N_9928,N_8184);
xor U13328 (N_13328,N_8049,N_11754);
xor U13329 (N_13329,N_9247,N_10842);
nand U13330 (N_13330,N_9562,N_11704);
or U13331 (N_13331,N_10041,N_9923);
or U13332 (N_13332,N_8679,N_10503);
or U13333 (N_13333,N_10729,N_10712);
nor U13334 (N_13334,N_9318,N_8419);
and U13335 (N_13335,N_11902,N_9755);
and U13336 (N_13336,N_8390,N_10495);
xnor U13337 (N_13337,N_11083,N_11194);
nand U13338 (N_13338,N_11494,N_8025);
xnor U13339 (N_13339,N_8686,N_9359);
and U13340 (N_13340,N_10366,N_9448);
and U13341 (N_13341,N_10029,N_9179);
or U13342 (N_13342,N_8880,N_11863);
xor U13343 (N_13343,N_8911,N_10755);
nor U13344 (N_13344,N_11368,N_9002);
xor U13345 (N_13345,N_8799,N_9444);
and U13346 (N_13346,N_11478,N_9171);
xnor U13347 (N_13347,N_10650,N_9091);
and U13348 (N_13348,N_10088,N_10555);
nand U13349 (N_13349,N_11267,N_10472);
xor U13350 (N_13350,N_8024,N_8438);
or U13351 (N_13351,N_8946,N_9656);
xor U13352 (N_13352,N_8252,N_10012);
xor U13353 (N_13353,N_11914,N_10172);
xor U13354 (N_13354,N_10750,N_10305);
nand U13355 (N_13355,N_8527,N_9188);
nor U13356 (N_13356,N_8900,N_10978);
and U13357 (N_13357,N_10407,N_9227);
or U13358 (N_13358,N_11770,N_9048);
nor U13359 (N_13359,N_8994,N_9683);
nor U13360 (N_13360,N_10816,N_9360);
nor U13361 (N_13361,N_9063,N_9089);
nand U13362 (N_13362,N_9232,N_9068);
or U13363 (N_13363,N_9501,N_10064);
or U13364 (N_13364,N_11527,N_10899);
nor U13365 (N_13365,N_11024,N_11779);
or U13366 (N_13366,N_9989,N_10371);
and U13367 (N_13367,N_10566,N_11723);
nand U13368 (N_13368,N_9492,N_11325);
and U13369 (N_13369,N_10836,N_10574);
nand U13370 (N_13370,N_9964,N_9669);
nand U13371 (N_13371,N_8132,N_10023);
nor U13372 (N_13372,N_9598,N_11012);
nor U13373 (N_13373,N_9542,N_8949);
or U13374 (N_13374,N_11802,N_11689);
or U13375 (N_13375,N_9913,N_8369);
xor U13376 (N_13376,N_11594,N_10878);
xnor U13377 (N_13377,N_8205,N_8032);
nor U13378 (N_13378,N_9677,N_9403);
nand U13379 (N_13379,N_8787,N_11237);
nand U13380 (N_13380,N_11847,N_8769);
or U13381 (N_13381,N_10000,N_11971);
xnor U13382 (N_13382,N_11646,N_10024);
xnor U13383 (N_13383,N_8815,N_9291);
xor U13384 (N_13384,N_9966,N_10425);
and U13385 (N_13385,N_10329,N_9582);
and U13386 (N_13386,N_10237,N_10850);
nand U13387 (N_13387,N_9158,N_8396);
nor U13388 (N_13388,N_10524,N_9797);
nand U13389 (N_13389,N_8620,N_8257);
and U13390 (N_13390,N_11922,N_10003);
and U13391 (N_13391,N_11017,N_9796);
nor U13392 (N_13392,N_8499,N_8321);
nor U13393 (N_13393,N_11581,N_10378);
nor U13394 (N_13394,N_11805,N_8138);
and U13395 (N_13395,N_11075,N_9466);
and U13396 (N_13396,N_9150,N_10793);
nand U13397 (N_13397,N_11207,N_9970);
and U13398 (N_13398,N_9647,N_9272);
nor U13399 (N_13399,N_11278,N_10968);
nor U13400 (N_13400,N_9265,N_9748);
nor U13401 (N_13401,N_11441,N_9042);
nor U13402 (N_13402,N_8354,N_10108);
and U13403 (N_13403,N_9266,N_8519);
and U13404 (N_13404,N_9895,N_9645);
nand U13405 (N_13405,N_11653,N_11560);
xnor U13406 (N_13406,N_9127,N_8047);
nor U13407 (N_13407,N_9952,N_11894);
nand U13408 (N_13408,N_11308,N_11131);
and U13409 (N_13409,N_9147,N_11877);
or U13410 (N_13410,N_9413,N_9060);
nand U13411 (N_13411,N_10913,N_8562);
and U13412 (N_13412,N_8520,N_9904);
xnor U13413 (N_13413,N_9866,N_8869);
and U13414 (N_13414,N_9133,N_11003);
nand U13415 (N_13415,N_8278,N_10185);
and U13416 (N_13416,N_9787,N_9947);
nand U13417 (N_13417,N_11963,N_8884);
and U13418 (N_13418,N_10243,N_11127);
xor U13419 (N_13419,N_8793,N_11071);
nor U13420 (N_13420,N_11825,N_10497);
nor U13421 (N_13421,N_10869,N_8204);
xor U13422 (N_13422,N_8714,N_10519);
xnor U13423 (N_13423,N_10715,N_10031);
and U13424 (N_13424,N_8504,N_8270);
nor U13425 (N_13425,N_8576,N_8702);
nand U13426 (N_13426,N_11899,N_11843);
xor U13427 (N_13427,N_9553,N_10922);
and U13428 (N_13428,N_8083,N_11160);
xnor U13429 (N_13429,N_11917,N_9679);
and U13430 (N_13430,N_9478,N_9114);
or U13431 (N_13431,N_9540,N_9464);
or U13432 (N_13432,N_10752,N_11430);
nand U13433 (N_13433,N_10196,N_11456);
nor U13434 (N_13434,N_10316,N_10073);
or U13435 (N_13435,N_9731,N_9486);
nand U13436 (N_13436,N_11337,N_9348);
nand U13437 (N_13437,N_8557,N_10941);
nor U13438 (N_13438,N_11080,N_9316);
and U13439 (N_13439,N_11170,N_8574);
xor U13440 (N_13440,N_8535,N_10810);
nor U13441 (N_13441,N_11424,N_9519);
xnor U13442 (N_13442,N_9733,N_11979);
or U13443 (N_13443,N_10564,N_10166);
xnor U13444 (N_13444,N_8241,N_11059);
xor U13445 (N_13445,N_10059,N_9695);
nor U13446 (N_13446,N_8388,N_11152);
and U13447 (N_13447,N_8948,N_8334);
or U13448 (N_13448,N_9213,N_10982);
nor U13449 (N_13449,N_9009,N_11680);
and U13450 (N_13450,N_9310,N_10430);
xor U13451 (N_13451,N_9833,N_8747);
xnor U13452 (N_13452,N_8857,N_8298);
nand U13453 (N_13453,N_10222,N_8852);
or U13454 (N_13454,N_11418,N_8847);
nand U13455 (N_13455,N_9084,N_8154);
nand U13456 (N_13456,N_10611,N_8104);
or U13457 (N_13457,N_9762,N_8411);
xnor U13458 (N_13458,N_10660,N_11094);
nand U13459 (N_13459,N_9839,N_10709);
or U13460 (N_13460,N_8833,N_10476);
or U13461 (N_13461,N_11353,N_10888);
or U13462 (N_13462,N_9915,N_8239);
nand U13463 (N_13463,N_9472,N_10863);
xnor U13464 (N_13464,N_9354,N_11452);
and U13465 (N_13465,N_11105,N_8146);
or U13466 (N_13466,N_10295,N_10039);
xor U13467 (N_13467,N_8020,N_9148);
nor U13468 (N_13468,N_10615,N_9716);
xor U13469 (N_13469,N_9579,N_11906);
nand U13470 (N_13470,N_9407,N_11471);
nor U13471 (N_13471,N_9688,N_10576);
nand U13472 (N_13472,N_9004,N_10350);
xor U13473 (N_13473,N_10897,N_8176);
nand U13474 (N_13474,N_9111,N_10690);
or U13475 (N_13475,N_11061,N_8332);
or U13476 (N_13476,N_9224,N_11270);
and U13477 (N_13477,N_11986,N_8592);
xor U13478 (N_13478,N_9668,N_10977);
or U13479 (N_13479,N_8446,N_8914);
and U13480 (N_13480,N_11028,N_8664);
xnor U13481 (N_13481,N_10362,N_8553);
nand U13482 (N_13482,N_11965,N_8403);
or U13483 (N_13483,N_8192,N_9338);
or U13484 (N_13484,N_9270,N_8484);
and U13485 (N_13485,N_11722,N_8105);
xnor U13486 (N_13486,N_9079,N_10786);
and U13487 (N_13487,N_11016,N_11969);
xnor U13488 (N_13488,N_10263,N_10719);
nand U13489 (N_13489,N_10431,N_9017);
and U13490 (N_13490,N_9474,N_9126);
xor U13491 (N_13491,N_8647,N_11153);
nor U13492 (N_13492,N_11885,N_8492);
and U13493 (N_13493,N_8089,N_8329);
xnor U13494 (N_13494,N_10441,N_9946);
and U13495 (N_13495,N_8006,N_10714);
xnor U13496 (N_13496,N_9592,N_11427);
nand U13497 (N_13497,N_10351,N_10630);
or U13498 (N_13498,N_11870,N_8673);
or U13499 (N_13499,N_10908,N_10297);
or U13500 (N_13500,N_11702,N_9577);
and U13501 (N_13501,N_9155,N_10547);
or U13502 (N_13502,N_8463,N_11093);
nand U13503 (N_13503,N_10130,N_8300);
and U13504 (N_13504,N_9160,N_10867);
or U13505 (N_13505,N_8588,N_8416);
and U13506 (N_13506,N_10095,N_9366);
and U13507 (N_13507,N_10151,N_9415);
and U13508 (N_13508,N_8683,N_8120);
or U13509 (N_13509,N_8258,N_11719);
nor U13510 (N_13510,N_8376,N_10718);
xor U13511 (N_13511,N_9993,N_9494);
and U13512 (N_13512,N_9557,N_11672);
or U13513 (N_13513,N_8757,N_10240);
nand U13514 (N_13514,N_9499,N_8710);
and U13515 (N_13515,N_9405,N_11598);
and U13516 (N_13516,N_9028,N_11934);
xnor U13517 (N_13517,N_8798,N_11778);
or U13518 (N_13518,N_10398,N_10068);
or U13519 (N_13519,N_8950,N_9963);
xnor U13520 (N_13520,N_10474,N_10177);
xnor U13521 (N_13521,N_11139,N_9955);
nand U13522 (N_13522,N_9302,N_9641);
or U13523 (N_13523,N_9032,N_10992);
xnor U13524 (N_13524,N_8927,N_11857);
nor U13525 (N_13525,N_8924,N_8483);
xor U13526 (N_13526,N_9129,N_11255);
xor U13527 (N_13527,N_11736,N_10567);
or U13528 (N_13528,N_10215,N_8465);
nor U13529 (N_13529,N_10923,N_11923);
or U13530 (N_13530,N_9700,N_11572);
nand U13531 (N_13531,N_8749,N_10146);
or U13532 (N_13532,N_10795,N_8197);
xnor U13533 (N_13533,N_9037,N_10096);
nor U13534 (N_13534,N_9041,N_9784);
and U13535 (N_13535,N_8708,N_9722);
and U13536 (N_13536,N_11262,N_8958);
nor U13537 (N_13537,N_8353,N_8565);
nand U13538 (N_13538,N_8122,N_10697);
xnor U13539 (N_13539,N_10387,N_8152);
nor U13540 (N_13540,N_10905,N_9984);
or U13541 (N_13541,N_8263,N_8651);
or U13542 (N_13542,N_9881,N_10638);
or U13543 (N_13543,N_8442,N_11266);
xor U13544 (N_13544,N_9867,N_9326);
nand U13545 (N_13545,N_11252,N_10489);
nor U13546 (N_13546,N_11021,N_9892);
xor U13547 (N_13547,N_8370,N_10627);
nand U13548 (N_13548,N_9093,N_11067);
and U13549 (N_13549,N_10355,N_9723);
nand U13550 (N_13550,N_11765,N_8696);
nand U13551 (N_13551,N_8970,N_9401);
xor U13552 (N_13552,N_11982,N_11664);
xnor U13553 (N_13553,N_11209,N_8194);
nand U13554 (N_13554,N_9917,N_9269);
nor U13555 (N_13555,N_8975,N_10183);
nand U13556 (N_13556,N_8405,N_10412);
nand U13557 (N_13557,N_11019,N_8919);
xnor U13558 (N_13558,N_11720,N_9872);
nor U13559 (N_13559,N_9973,N_11136);
xnor U13560 (N_13560,N_10492,N_8628);
xnor U13561 (N_13561,N_11939,N_9086);
nor U13562 (N_13562,N_11388,N_8330);
nand U13563 (N_13563,N_8572,N_9576);
and U13564 (N_13564,N_10091,N_11812);
nand U13565 (N_13565,N_11144,N_8493);
xor U13566 (N_13566,N_10109,N_11391);
xor U13567 (N_13567,N_9446,N_8137);
and U13568 (N_13568,N_10250,N_10700);
xnor U13569 (N_13569,N_11996,N_11053);
and U13570 (N_13570,N_8142,N_11137);
xor U13571 (N_13571,N_8393,N_9918);
nand U13572 (N_13572,N_8115,N_8823);
xnor U13573 (N_13573,N_8718,N_8287);
nor U13574 (N_13574,N_9829,N_9040);
and U13575 (N_13575,N_8777,N_9850);
and U13576 (N_13576,N_8454,N_10379);
or U13577 (N_13577,N_9014,N_10484);
nand U13578 (N_13578,N_10027,N_8040);
or U13579 (N_13579,N_8842,N_9412);
nand U13580 (N_13580,N_11335,N_11623);
and U13581 (N_13581,N_10694,N_8042);
and U13582 (N_13582,N_11567,N_10783);
xor U13583 (N_13583,N_8929,N_9546);
and U13584 (N_13584,N_11146,N_10051);
nor U13585 (N_13585,N_11156,N_10061);
and U13586 (N_13586,N_11150,N_11844);
and U13587 (N_13587,N_11192,N_8299);
and U13588 (N_13588,N_10791,N_9331);
nand U13589 (N_13589,N_10951,N_8322);
xnor U13590 (N_13590,N_9142,N_9209);
nor U13591 (N_13591,N_8953,N_8487);
or U13592 (N_13592,N_10276,N_8839);
nor U13593 (N_13593,N_8168,N_10789);
nor U13594 (N_13594,N_9729,N_9652);
and U13595 (N_13595,N_9432,N_9249);
nor U13596 (N_13596,N_11613,N_9047);
xnor U13597 (N_13597,N_11332,N_11853);
nor U13598 (N_13598,N_11377,N_10469);
or U13599 (N_13599,N_8657,N_9538);
or U13600 (N_13600,N_10145,N_11492);
and U13601 (N_13601,N_8477,N_10972);
nand U13602 (N_13602,N_8113,N_10538);
and U13603 (N_13603,N_8433,N_9686);
xnor U13604 (N_13604,N_11409,N_9705);
or U13605 (N_13605,N_10805,N_9178);
nand U13606 (N_13606,N_10160,N_10771);
nor U13607 (N_13607,N_11101,N_8979);
or U13608 (N_13608,N_9076,N_11511);
nand U13609 (N_13609,N_10312,N_11544);
xnor U13610 (N_13610,N_9001,N_8577);
nand U13611 (N_13611,N_10506,N_9935);
nor U13612 (N_13612,N_8159,N_9590);
nor U13613 (N_13613,N_8707,N_11140);
xor U13614 (N_13614,N_8587,N_10219);
and U13615 (N_13615,N_9995,N_11788);
or U13616 (N_13616,N_9632,N_9949);
and U13617 (N_13617,N_9618,N_10195);
nor U13618 (N_13618,N_10110,N_11756);
nor U13619 (N_13619,N_9408,N_9570);
nand U13620 (N_13620,N_9429,N_9742);
nand U13621 (N_13621,N_9106,N_10277);
nor U13622 (N_13622,N_10290,N_10505);
nor U13623 (N_13623,N_8162,N_11727);
and U13624 (N_13624,N_9252,N_11381);
or U13625 (N_13625,N_10089,N_8893);
and U13626 (N_13626,N_9328,N_11364);
and U13627 (N_13627,N_10619,N_8656);
or U13628 (N_13628,N_10556,N_9745);
nand U13629 (N_13629,N_10612,N_11806);
and U13630 (N_13630,N_10467,N_8629);
or U13631 (N_13631,N_11277,N_11013);
nor U13632 (N_13632,N_10954,N_11264);
or U13633 (N_13633,N_8422,N_11508);
xnor U13634 (N_13634,N_11063,N_9427);
and U13635 (N_13635,N_8861,N_11640);
nor U13636 (N_13636,N_9480,N_10594);
nand U13637 (N_13637,N_10677,N_8223);
nand U13638 (N_13638,N_9701,N_10074);
or U13639 (N_13639,N_9157,N_9136);
nor U13640 (N_13640,N_11500,N_11279);
xnor U13641 (N_13641,N_11111,N_9159);
nor U13642 (N_13642,N_8341,N_9953);
xor U13643 (N_13643,N_9670,N_11461);
nand U13644 (N_13644,N_8226,N_9511);
nor U13645 (N_13645,N_11978,N_11981);
nor U13646 (N_13646,N_10826,N_9320);
nand U13647 (N_13647,N_11999,N_10283);
and U13648 (N_13648,N_11631,N_11480);
nor U13649 (N_13649,N_8190,N_8711);
nor U13650 (N_13650,N_10676,N_10338);
or U13651 (N_13651,N_8171,N_11241);
nand U13652 (N_13652,N_10684,N_10879);
or U13653 (N_13653,N_10552,N_9183);
nor U13654 (N_13654,N_9763,N_11507);
and U13655 (N_13655,N_8100,N_9836);
xor U13656 (N_13656,N_11213,N_10349);
and U13657 (N_13657,N_9363,N_9558);
xor U13658 (N_13658,N_10421,N_11909);
or U13659 (N_13659,N_8762,N_11276);
nand U13660 (N_13660,N_10056,N_9217);
nand U13661 (N_13661,N_9162,N_8800);
or U13662 (N_13662,N_9046,N_10049);
and U13663 (N_13663,N_11285,N_11609);
or U13664 (N_13664,N_8292,N_10647);
nand U13665 (N_13665,N_8342,N_8486);
and U13666 (N_13666,N_9853,N_8054);
and U13667 (N_13667,N_8078,N_9424);
nor U13668 (N_13668,N_8648,N_10462);
and U13669 (N_13669,N_10640,N_10925);
and U13670 (N_13670,N_8650,N_10409);
xnor U13671 (N_13671,N_10830,N_11301);
nor U13672 (N_13672,N_9031,N_8450);
and U13673 (N_13673,N_8098,N_11240);
nand U13674 (N_13674,N_8509,N_8018);
and U13675 (N_13675,N_9223,N_8013);
or U13676 (N_13676,N_11635,N_8448);
nand U13677 (N_13677,N_9262,N_8751);
nand U13678 (N_13678,N_9030,N_9261);
nor U13679 (N_13679,N_8665,N_8640);
nor U13680 (N_13680,N_10253,N_9211);
xnor U13681 (N_13681,N_11684,N_9555);
or U13682 (N_13682,N_10348,N_11731);
or U13683 (N_13683,N_10171,N_10999);
or U13684 (N_13684,N_11496,N_10541);
and U13685 (N_13685,N_9024,N_11095);
nand U13686 (N_13686,N_8513,N_10717);
nor U13687 (N_13687,N_9623,N_10570);
nor U13688 (N_13688,N_9919,N_8165);
nor U13689 (N_13689,N_10659,N_11202);
nor U13690 (N_13690,N_10299,N_10286);
nand U13691 (N_13691,N_11910,N_9908);
or U13692 (N_13692,N_10507,N_10225);
xor U13693 (N_13693,N_9016,N_8874);
xor U13694 (N_13694,N_10001,N_9967);
and U13695 (N_13695,N_9943,N_11218);
nand U13696 (N_13696,N_8879,N_11873);
or U13697 (N_13697,N_10373,N_11420);
nor U13698 (N_13698,N_9228,N_10883);
xnor U13699 (N_13699,N_11707,N_11865);
nand U13700 (N_13700,N_11076,N_9854);
nor U13701 (N_13701,N_8856,N_11244);
xor U13702 (N_13702,N_8967,N_8005);
nand U13703 (N_13703,N_9921,N_9315);
nand U13704 (N_13704,N_9692,N_8818);
xnor U13705 (N_13705,N_11118,N_10639);
xor U13706 (N_13706,N_9619,N_9425);
and U13707 (N_13707,N_11525,N_8715);
nor U13708 (N_13708,N_9870,N_11881);
and U13709 (N_13709,N_8266,N_8294);
or U13710 (N_13710,N_11968,N_8597);
and U13711 (N_13711,N_10204,N_10645);
and U13712 (N_13712,N_11273,N_11787);
xnor U13713 (N_13713,N_9118,N_9257);
nand U13714 (N_13714,N_8693,N_10100);
or U13715 (N_13715,N_11913,N_11318);
xor U13716 (N_13716,N_9544,N_10163);
and U13717 (N_13717,N_9899,N_9610);
nor U13718 (N_13718,N_11446,N_9901);
nor U13719 (N_13719,N_8820,N_8796);
xor U13720 (N_13720,N_8555,N_8359);
xnor U13721 (N_13721,N_8022,N_9462);
nor U13722 (N_13722,N_10726,N_8130);
and U13723 (N_13723,N_8027,N_9891);
or U13724 (N_13724,N_8380,N_9856);
xnor U13725 (N_13725,N_11531,N_8048);
and U13726 (N_13726,N_10006,N_10468);
xor U13727 (N_13727,N_8604,N_9626);
xor U13728 (N_13728,N_9842,N_8637);
or U13729 (N_13729,N_9968,N_8038);
and U13730 (N_13730,N_9805,N_8770);
nand U13731 (N_13731,N_8947,N_8275);
nand U13732 (N_13732,N_10987,N_10158);
nand U13733 (N_13733,N_10084,N_11542);
nor U13734 (N_13734,N_11993,N_8964);
and U13735 (N_13735,N_8431,N_9053);
nand U13736 (N_13736,N_8908,N_9453);
or U13737 (N_13737,N_9170,N_10797);
xnor U13738 (N_13738,N_9815,N_8624);
and U13739 (N_13739,N_11589,N_9621);
nand U13740 (N_13740,N_9066,N_8424);
xor U13741 (N_13741,N_8235,N_9134);
or U13742 (N_13742,N_9754,N_9807);
and U13743 (N_13743,N_10267,N_9625);
nand U13744 (N_13744,N_8817,N_11176);
nand U13745 (N_13745,N_9845,N_9684);
xor U13746 (N_13746,N_11000,N_8053);
xnor U13747 (N_13747,N_10956,N_8068);
xnor U13748 (N_13748,N_10796,N_9387);
or U13749 (N_13749,N_11869,N_8362);
and U13750 (N_13750,N_11748,N_8019);
and U13751 (N_13751,N_9750,N_8474);
or U13752 (N_13752,N_8214,N_11546);
nor U13753 (N_13753,N_10159,N_11970);
xnor U13754 (N_13754,N_9795,N_11611);
or U13755 (N_13755,N_9991,N_9981);
nor U13756 (N_13756,N_8658,N_10090);
or U13757 (N_13757,N_10376,N_9377);
xnor U13758 (N_13758,N_9220,N_11859);
nand U13759 (N_13759,N_9476,N_10543);
nor U13760 (N_13760,N_8290,N_9152);
nor U13761 (N_13761,N_8316,N_8206);
nand U13762 (N_13762,N_9513,N_8457);
nand U13763 (N_13763,N_11738,N_10738);
or U13764 (N_13764,N_8220,N_8436);
and U13765 (N_13765,N_10434,N_10790);
nand U13766 (N_13766,N_9275,N_9860);
or U13767 (N_13767,N_11661,N_10361);
or U13768 (N_13768,N_8678,N_8726);
nand U13769 (N_13769,N_8663,N_11540);
and U13770 (N_13770,N_8288,N_8551);
nor U13771 (N_13771,N_10824,N_8351);
nor U13772 (N_13772,N_9181,N_11632);
or U13773 (N_13773,N_11622,N_8988);
xnor U13774 (N_13774,N_10960,N_11211);
or U13775 (N_13775,N_10641,N_8143);
nand U13776 (N_13776,N_9753,N_11440);
and U13777 (N_13777,N_8907,N_10370);
and U13778 (N_13778,N_10365,N_11102);
and U13779 (N_13779,N_10931,N_9021);
and U13780 (N_13780,N_9436,N_10749);
nand U13781 (N_13781,N_10396,N_8178);
nor U13782 (N_13782,N_9391,N_11549);
or U13783 (N_13783,N_11950,N_9922);
nand U13784 (N_13784,N_8963,N_11987);
nor U13785 (N_13785,N_9906,N_10482);
or U13786 (N_13786,N_8653,N_8439);
and U13787 (N_13787,N_10175,N_10971);
nor U13788 (N_13788,N_9644,N_10256);
or U13789 (N_13789,N_11283,N_8470);
and U13790 (N_13790,N_8319,N_8586);
nor U13791 (N_13791,N_11081,N_8174);
xnor U13792 (N_13792,N_11079,N_11955);
or U13793 (N_13793,N_9451,N_8784);
xnor U13794 (N_13794,N_10180,N_8836);
nand U13795 (N_13795,N_11245,N_8736);
or U13796 (N_13796,N_8428,N_9554);
nand U13797 (N_13797,N_11096,N_10632);
nor U13798 (N_13798,N_10284,N_11772);
and U13799 (N_13799,N_11676,N_11882);
nor U13800 (N_13800,N_10438,N_10957);
nor U13801 (N_13801,N_11547,N_10191);
xor U13802 (N_13802,N_9638,N_9821);
nand U13803 (N_13803,N_9661,N_10911);
nor U13804 (N_13804,N_9273,N_9556);
xnor U13805 (N_13805,N_10042,N_9367);
and U13806 (N_13806,N_8123,N_8308);
nand U13807 (N_13807,N_11943,N_9234);
nand U13808 (N_13808,N_8706,N_8980);
or U13809 (N_13809,N_10707,N_10303);
nor U13810 (N_13810,N_11907,N_10975);
nand U13811 (N_13811,N_9088,N_9799);
nand U13812 (N_13812,N_11314,N_8456);
nand U13813 (N_13813,N_8897,N_10624);
nand U13814 (N_13814,N_10573,N_8447);
and U13815 (N_13815,N_11371,N_10930);
and U13816 (N_13816,N_11330,N_9907);
nand U13817 (N_13817,N_10661,N_11195);
xnor U13818 (N_13818,N_9071,N_10991);
or U13819 (N_13819,N_8090,N_10458);
or U13820 (N_13820,N_9735,N_10565);
or U13821 (N_13821,N_8677,N_10190);
and U13822 (N_13822,N_8057,N_8383);
and U13823 (N_13823,N_8267,N_11054);
nor U13824 (N_13824,N_11584,N_10079);
or U13825 (N_13825,N_8766,N_10310);
nor U13826 (N_13826,N_8567,N_9711);
nand U13827 (N_13827,N_11148,N_10874);
and U13828 (N_13828,N_10165,N_9495);
nand U13829 (N_13829,N_11590,N_11462);
nand U13830 (N_13830,N_11357,N_8085);
and U13831 (N_13831,N_8094,N_8139);
nor U13832 (N_13832,N_10917,N_9741);
nor U13833 (N_13833,N_11620,N_9277);
nand U13834 (N_13834,N_11915,N_11976);
or U13835 (N_13835,N_10581,N_10550);
nand U13836 (N_13836,N_9201,N_9889);
nor U13837 (N_13837,N_9337,N_10643);
xor U13838 (N_13838,N_8240,N_11848);
or U13839 (N_13839,N_9225,N_9808);
nand U13840 (N_13840,N_9398,N_10741);
nor U13841 (N_13841,N_11310,N_11888);
nor U13842 (N_13842,N_11117,N_10979);
or U13843 (N_13843,N_9777,N_9151);
xnor U13844 (N_13844,N_10812,N_11833);
xnor U13845 (N_13845,N_8738,N_9584);
xnor U13846 (N_13846,N_9768,N_8878);
xnor U13847 (N_13847,N_11580,N_11940);
xnor U13848 (N_13848,N_11998,N_9508);
nand U13849 (N_13849,N_9605,N_9219);
nor U13850 (N_13850,N_10043,N_10320);
nand U13851 (N_13851,N_11483,N_10698);
nor U13852 (N_13852,N_8186,N_11884);
xor U13853 (N_13853,N_10117,N_9979);
and U13854 (N_13854,N_9548,N_10463);
or U13855 (N_13855,N_10121,N_11321);
xor U13856 (N_13856,N_10587,N_8773);
xor U13857 (N_13857,N_10058,N_11610);
nand U13858 (N_13858,N_10063,N_10494);
and U13859 (N_13859,N_8413,N_10226);
nor U13860 (N_13860,N_9121,N_10033);
and U13861 (N_13861,N_10436,N_9689);
and U13862 (N_13862,N_9775,N_9602);
nor U13863 (N_13863,N_10465,N_11690);
and U13864 (N_13864,N_9685,N_10572);
nand U13865 (N_13865,N_9307,N_10028);
nand U13866 (N_13866,N_11151,N_10113);
nor U13867 (N_13867,N_8745,N_9837);
or U13868 (N_13868,N_10890,N_9064);
or U13869 (N_13869,N_10461,N_9154);
nor U13870 (N_13870,N_8444,N_11708);
nor U13871 (N_13871,N_9006,N_10437);
nand U13872 (N_13872,N_9132,N_9725);
xnor U13873 (N_13873,N_10354,N_8381);
xor U13874 (N_13874,N_10342,N_11468);
nor U13875 (N_13875,N_8253,N_11488);
xor U13876 (N_13876,N_11980,N_11057);
nand U13877 (N_13877,N_9336,N_9936);
nor U13878 (N_13878,N_8915,N_9329);
nor U13879 (N_13879,N_11233,N_9124);
or U13880 (N_13880,N_9029,N_9371);
nand U13881 (N_13881,N_11619,N_9960);
nor U13882 (N_13882,N_8118,N_8617);
xnor U13883 (N_13883,N_9475,N_10990);
nand U13884 (N_13884,N_8337,N_10558);
nand U13885 (N_13885,N_8114,N_8891);
xor U13886 (N_13886,N_11856,N_8225);
xor U13887 (N_13887,N_9663,N_8417);
nor U13888 (N_13888,N_11161,N_11654);
nor U13889 (N_13889,N_11816,N_9381);
nor U13890 (N_13890,N_8502,N_11536);
or U13891 (N_13891,N_9502,N_9999);
and U13892 (N_13892,N_8109,N_10675);
and U13893 (N_13893,N_8841,N_9580);
nand U13894 (N_13894,N_11091,N_11783);
and U13895 (N_13895,N_10514,N_9604);
nor U13896 (N_13896,N_9586,N_9058);
and U13897 (N_13897,N_8582,N_8669);
nor U13898 (N_13898,N_11808,N_11801);
or U13899 (N_13899,N_8595,N_10540);
nor U13900 (N_13900,N_10097,N_11284);
and U13901 (N_13901,N_10886,N_11786);
nand U13902 (N_13902,N_10739,N_8453);
or U13903 (N_13903,N_10128,N_8441);
nor U13904 (N_13904,N_9938,N_10452);
or U13905 (N_13905,N_10769,N_8172);
nand U13906 (N_13906,N_8406,N_9489);
and U13907 (N_13907,N_11918,N_9484);
xor U13908 (N_13908,N_11458,N_8972);
nor U13909 (N_13909,N_8583,N_10032);
and U13910 (N_13910,N_8471,N_8497);
xnor U13911 (N_13911,N_11412,N_11991);
or U13912 (N_13912,N_8285,N_9608);
nand U13913 (N_13913,N_11798,N_11875);
and U13914 (N_13914,N_8616,N_11973);
or U13915 (N_13915,N_10753,N_11685);
xnor U13916 (N_13916,N_8074,N_10807);
nand U13917 (N_13917,N_10872,N_8764);
nand U13918 (N_13918,N_9847,N_11185);
and U13919 (N_13919,N_11450,N_11530);
xnor U13920 (N_13920,N_11617,N_11122);
xnor U13921 (N_13921,N_8589,N_8248);
and U13922 (N_13922,N_9672,N_9543);
or U13923 (N_13923,N_8498,N_9788);
nor U13924 (N_13924,N_10603,N_8324);
nand U13925 (N_13925,N_9634,N_9299);
nor U13926 (N_13926,N_9665,N_8423);
or U13927 (N_13927,N_11116,N_8093);
nand U13928 (N_13928,N_11401,N_9253);
xor U13929 (N_13929,N_8840,N_10131);
nand U13930 (N_13930,N_10622,N_8480);
or U13931 (N_13931,N_11629,N_9691);
and U13932 (N_13932,N_8885,N_10831);
nand U13933 (N_13933,N_10633,N_10523);
xor U13934 (N_13934,N_9868,N_8794);
xor U13935 (N_13935,N_9783,N_9052);
xnor U13936 (N_13936,N_11837,N_11044);
xnor U13937 (N_13937,N_8173,N_9390);
nand U13938 (N_13938,N_10728,N_10870);
nor U13939 (N_13939,N_10912,N_9471);
xor U13940 (N_13940,N_11354,N_8421);
and U13941 (N_13941,N_10663,N_9404);
xor U13942 (N_13942,N_10852,N_11626);
nor U13943 (N_13943,N_9073,N_11974);
nand U13944 (N_13944,N_10265,N_10577);
nand U13945 (N_13945,N_8902,N_11828);
or U13946 (N_13946,N_8641,N_10595);
nor U13947 (N_13947,N_11502,N_11587);
or U13948 (N_13948,N_11311,N_8872);
nand U13949 (N_13949,N_9869,N_10213);
or U13950 (N_13950,N_9345,N_9180);
nor U13951 (N_13951,N_8238,N_8110);
or U13952 (N_13952,N_10114,N_10380);
nor U13953 (N_13953,N_9373,N_9370);
nor U13954 (N_13954,N_11861,N_9416);
nand U13955 (N_13955,N_10454,N_8549);
and U13956 (N_13956,N_11414,N_8865);
or U13957 (N_13957,N_11669,N_8361);
and U13958 (N_13958,N_11957,N_9613);
or U13959 (N_13959,N_9959,N_11564);
nand U13960 (N_13960,N_10077,N_9766);
xor U13961 (N_13961,N_10794,N_11199);
and U13962 (N_13962,N_9440,N_11528);
nand U13963 (N_13963,N_11954,N_10334);
and U13964 (N_13964,N_10598,N_9439);
nand U13965 (N_13965,N_10418,N_10238);
xor U13966 (N_13966,N_9790,N_9714);
xnor U13967 (N_13967,N_9267,N_9549);
and U13968 (N_13968,N_8035,N_9221);
xor U13969 (N_13969,N_10829,N_9301);
or U13970 (N_13970,N_11366,N_11990);
and U13971 (N_13971,N_8792,N_9758);
and U13972 (N_13972,N_11165,N_9099);
and U13973 (N_13973,N_8482,N_10866);
xor U13974 (N_13974,N_10164,N_8274);
nor U13975 (N_13975,N_8124,N_11706);
xnor U13976 (N_13976,N_10464,N_11559);
xnor U13977 (N_13977,N_11112,N_11236);
nor U13978 (N_13978,N_10608,N_8895);
nor U13979 (N_13979,N_10920,N_9773);
nor U13980 (N_13980,N_10658,N_10007);
or U13981 (N_13981,N_9203,N_8675);
and U13982 (N_13982,N_8014,N_11761);
and U13983 (N_13983,N_11766,N_10390);
xnor U13984 (N_13984,N_8713,N_9039);
nor U13985 (N_13985,N_11807,N_8568);
or U13986 (N_13986,N_11698,N_11421);
nor U13987 (N_13987,N_10471,N_11630);
xor U13988 (N_13988,N_8913,N_9737);
or U13989 (N_13989,N_9409,N_9545);
nor U13990 (N_13990,N_10037,N_8835);
xor U13991 (N_13991,N_11225,N_10483);
nand U13992 (N_13992,N_11363,N_9135);
xor U13993 (N_13993,N_10782,N_9469);
or U13994 (N_13994,N_8609,N_11347);
xor U13995 (N_13995,N_11269,N_8731);
xor U13996 (N_13996,N_8464,N_11935);
nand U13997 (N_13997,N_11545,N_8600);
nor U13998 (N_13998,N_10906,N_9308);
nand U13999 (N_13999,N_8001,N_8067);
and U14000 (N_14000,N_11778,N_11202);
nor U14001 (N_14001,N_10197,N_11394);
nand U14002 (N_14002,N_8963,N_10143);
and U14003 (N_14003,N_10592,N_8378);
xnor U14004 (N_14004,N_8185,N_9670);
nand U14005 (N_14005,N_10200,N_9188);
and U14006 (N_14006,N_11460,N_9095);
nand U14007 (N_14007,N_11127,N_10900);
xnor U14008 (N_14008,N_11449,N_8312);
and U14009 (N_14009,N_8236,N_10858);
or U14010 (N_14010,N_11465,N_8170);
and U14011 (N_14011,N_11750,N_8168);
and U14012 (N_14012,N_9736,N_8530);
nand U14013 (N_14013,N_11079,N_11961);
or U14014 (N_14014,N_11293,N_10635);
nor U14015 (N_14015,N_11996,N_8118);
xnor U14016 (N_14016,N_8084,N_8346);
nor U14017 (N_14017,N_9081,N_8198);
nand U14018 (N_14018,N_9837,N_10594);
or U14019 (N_14019,N_8098,N_11388);
or U14020 (N_14020,N_11357,N_9956);
or U14021 (N_14021,N_11659,N_11462);
xor U14022 (N_14022,N_10309,N_9074);
or U14023 (N_14023,N_9620,N_8406);
and U14024 (N_14024,N_8580,N_8770);
and U14025 (N_14025,N_9472,N_11229);
xnor U14026 (N_14026,N_11102,N_10008);
nor U14027 (N_14027,N_9679,N_9115);
xor U14028 (N_14028,N_9711,N_11836);
xor U14029 (N_14029,N_11780,N_9181);
or U14030 (N_14030,N_10647,N_9660);
and U14031 (N_14031,N_8339,N_11874);
xor U14032 (N_14032,N_11969,N_8161);
nor U14033 (N_14033,N_10230,N_8825);
and U14034 (N_14034,N_8081,N_11096);
xor U14035 (N_14035,N_11881,N_11724);
or U14036 (N_14036,N_9517,N_9627);
and U14037 (N_14037,N_11715,N_9823);
and U14038 (N_14038,N_9999,N_9410);
or U14039 (N_14039,N_10465,N_9518);
and U14040 (N_14040,N_11381,N_11943);
nand U14041 (N_14041,N_8936,N_11780);
nand U14042 (N_14042,N_9074,N_10205);
and U14043 (N_14043,N_10901,N_11924);
xnor U14044 (N_14044,N_11819,N_10771);
nor U14045 (N_14045,N_11185,N_10304);
nor U14046 (N_14046,N_10114,N_8495);
or U14047 (N_14047,N_9452,N_8942);
and U14048 (N_14048,N_10347,N_8004);
nor U14049 (N_14049,N_11776,N_8211);
and U14050 (N_14050,N_9623,N_9880);
xor U14051 (N_14051,N_9641,N_9217);
nand U14052 (N_14052,N_9086,N_8224);
xnor U14053 (N_14053,N_10191,N_11176);
xor U14054 (N_14054,N_8620,N_10769);
nor U14055 (N_14055,N_11948,N_11899);
xor U14056 (N_14056,N_10609,N_11031);
nor U14057 (N_14057,N_11836,N_9872);
and U14058 (N_14058,N_11412,N_8326);
nand U14059 (N_14059,N_10064,N_9710);
and U14060 (N_14060,N_10202,N_8647);
or U14061 (N_14061,N_9260,N_8612);
xor U14062 (N_14062,N_9490,N_8234);
xnor U14063 (N_14063,N_10745,N_10285);
nand U14064 (N_14064,N_10861,N_9559);
nand U14065 (N_14065,N_8775,N_9523);
nand U14066 (N_14066,N_11012,N_11246);
or U14067 (N_14067,N_8373,N_10795);
or U14068 (N_14068,N_9879,N_9911);
xnor U14069 (N_14069,N_11426,N_11938);
nor U14070 (N_14070,N_9297,N_10308);
xor U14071 (N_14071,N_9027,N_9130);
or U14072 (N_14072,N_8579,N_10168);
nor U14073 (N_14073,N_10519,N_11459);
or U14074 (N_14074,N_10993,N_9151);
nand U14075 (N_14075,N_8022,N_8471);
or U14076 (N_14076,N_9347,N_11284);
xor U14077 (N_14077,N_9792,N_8662);
nand U14078 (N_14078,N_10446,N_11686);
and U14079 (N_14079,N_8479,N_9369);
xor U14080 (N_14080,N_10393,N_8843);
nor U14081 (N_14081,N_9710,N_8307);
xnor U14082 (N_14082,N_10149,N_11635);
and U14083 (N_14083,N_9248,N_8630);
nand U14084 (N_14084,N_8907,N_9693);
or U14085 (N_14085,N_9361,N_8060);
nand U14086 (N_14086,N_11512,N_8396);
and U14087 (N_14087,N_8303,N_10832);
xnor U14088 (N_14088,N_8770,N_10827);
and U14089 (N_14089,N_9010,N_9888);
nand U14090 (N_14090,N_9795,N_11285);
nor U14091 (N_14091,N_8137,N_9174);
and U14092 (N_14092,N_10097,N_8288);
nor U14093 (N_14093,N_8202,N_8615);
xor U14094 (N_14094,N_11904,N_8224);
xor U14095 (N_14095,N_10093,N_11055);
nor U14096 (N_14096,N_9405,N_11144);
nand U14097 (N_14097,N_11700,N_11177);
and U14098 (N_14098,N_9693,N_9488);
nor U14099 (N_14099,N_10694,N_10825);
nor U14100 (N_14100,N_9355,N_9906);
xnor U14101 (N_14101,N_9997,N_9438);
and U14102 (N_14102,N_11725,N_10655);
xor U14103 (N_14103,N_8985,N_10102);
nor U14104 (N_14104,N_9957,N_9403);
nand U14105 (N_14105,N_10464,N_9637);
nor U14106 (N_14106,N_9296,N_10793);
xnor U14107 (N_14107,N_9520,N_10233);
xnor U14108 (N_14108,N_9267,N_8364);
nor U14109 (N_14109,N_11371,N_11872);
xnor U14110 (N_14110,N_11568,N_8711);
nand U14111 (N_14111,N_9290,N_8112);
and U14112 (N_14112,N_8452,N_11081);
and U14113 (N_14113,N_9048,N_11289);
and U14114 (N_14114,N_9255,N_11877);
nor U14115 (N_14115,N_8257,N_10073);
xnor U14116 (N_14116,N_10179,N_8448);
nor U14117 (N_14117,N_8360,N_8840);
or U14118 (N_14118,N_9824,N_9880);
and U14119 (N_14119,N_9311,N_8593);
nand U14120 (N_14120,N_11675,N_10694);
and U14121 (N_14121,N_8247,N_11045);
or U14122 (N_14122,N_8557,N_11718);
xor U14123 (N_14123,N_11854,N_9231);
nand U14124 (N_14124,N_11872,N_10298);
nand U14125 (N_14125,N_9983,N_9635);
nand U14126 (N_14126,N_8307,N_9263);
nor U14127 (N_14127,N_11239,N_8243);
nand U14128 (N_14128,N_8499,N_11200);
nand U14129 (N_14129,N_10958,N_9639);
and U14130 (N_14130,N_8107,N_9566);
nor U14131 (N_14131,N_8441,N_10208);
or U14132 (N_14132,N_11630,N_9737);
nor U14133 (N_14133,N_9809,N_8523);
nor U14134 (N_14134,N_8764,N_8171);
and U14135 (N_14135,N_9335,N_11896);
nor U14136 (N_14136,N_8113,N_10168);
nand U14137 (N_14137,N_10393,N_11607);
xor U14138 (N_14138,N_8069,N_9372);
nand U14139 (N_14139,N_8755,N_8771);
or U14140 (N_14140,N_10088,N_8505);
xnor U14141 (N_14141,N_11293,N_11321);
and U14142 (N_14142,N_9250,N_10528);
nand U14143 (N_14143,N_11257,N_8893);
xnor U14144 (N_14144,N_8531,N_8680);
xor U14145 (N_14145,N_8959,N_9053);
nor U14146 (N_14146,N_11443,N_8393);
nor U14147 (N_14147,N_10449,N_9495);
xnor U14148 (N_14148,N_10287,N_10632);
nor U14149 (N_14149,N_9566,N_8169);
and U14150 (N_14150,N_10964,N_10364);
and U14151 (N_14151,N_10251,N_9403);
xnor U14152 (N_14152,N_11606,N_9386);
and U14153 (N_14153,N_8384,N_11911);
nand U14154 (N_14154,N_8352,N_10252);
or U14155 (N_14155,N_9819,N_10516);
or U14156 (N_14156,N_11494,N_11632);
xnor U14157 (N_14157,N_9815,N_9183);
nor U14158 (N_14158,N_10330,N_11331);
nand U14159 (N_14159,N_8536,N_8800);
nand U14160 (N_14160,N_11313,N_10391);
nor U14161 (N_14161,N_9383,N_9922);
nand U14162 (N_14162,N_8062,N_11320);
nor U14163 (N_14163,N_10381,N_11665);
nand U14164 (N_14164,N_10213,N_8085);
nor U14165 (N_14165,N_9636,N_11073);
or U14166 (N_14166,N_10952,N_10604);
nor U14167 (N_14167,N_10373,N_10290);
or U14168 (N_14168,N_8385,N_8621);
xnor U14169 (N_14169,N_11572,N_10025);
xor U14170 (N_14170,N_11569,N_11373);
nand U14171 (N_14171,N_11187,N_8631);
and U14172 (N_14172,N_10182,N_10157);
and U14173 (N_14173,N_10494,N_8035);
xor U14174 (N_14174,N_8793,N_10584);
and U14175 (N_14175,N_8846,N_8671);
nand U14176 (N_14176,N_11526,N_8262);
nor U14177 (N_14177,N_11377,N_9646);
xnor U14178 (N_14178,N_9007,N_11905);
or U14179 (N_14179,N_10849,N_11158);
and U14180 (N_14180,N_9456,N_8276);
nand U14181 (N_14181,N_9678,N_9714);
nand U14182 (N_14182,N_10312,N_8950);
or U14183 (N_14183,N_10565,N_9157);
and U14184 (N_14184,N_11058,N_8892);
xnor U14185 (N_14185,N_9988,N_8585);
nor U14186 (N_14186,N_9617,N_10542);
nand U14187 (N_14187,N_8762,N_11336);
nor U14188 (N_14188,N_11137,N_11799);
and U14189 (N_14189,N_11444,N_11310);
or U14190 (N_14190,N_11954,N_8525);
or U14191 (N_14191,N_11440,N_9424);
xnor U14192 (N_14192,N_11152,N_10303);
xnor U14193 (N_14193,N_10813,N_11647);
nor U14194 (N_14194,N_9518,N_9177);
and U14195 (N_14195,N_10799,N_8545);
nor U14196 (N_14196,N_9234,N_9946);
or U14197 (N_14197,N_10309,N_8482);
nor U14198 (N_14198,N_8829,N_8203);
nand U14199 (N_14199,N_10545,N_9875);
xnor U14200 (N_14200,N_11816,N_11402);
nand U14201 (N_14201,N_9036,N_10603);
or U14202 (N_14202,N_8445,N_10900);
nand U14203 (N_14203,N_9809,N_8687);
nor U14204 (N_14204,N_10997,N_8833);
nand U14205 (N_14205,N_10730,N_9983);
nor U14206 (N_14206,N_10674,N_8146);
nor U14207 (N_14207,N_10032,N_10800);
and U14208 (N_14208,N_11219,N_10668);
nor U14209 (N_14209,N_8233,N_9785);
nor U14210 (N_14210,N_11266,N_9985);
nand U14211 (N_14211,N_11946,N_11087);
nor U14212 (N_14212,N_8003,N_9271);
nor U14213 (N_14213,N_8249,N_9944);
nand U14214 (N_14214,N_10194,N_9727);
nand U14215 (N_14215,N_8116,N_11720);
nand U14216 (N_14216,N_8462,N_8041);
and U14217 (N_14217,N_9884,N_10445);
nor U14218 (N_14218,N_11204,N_8982);
nor U14219 (N_14219,N_11624,N_8386);
nor U14220 (N_14220,N_10230,N_10853);
or U14221 (N_14221,N_9654,N_11957);
xor U14222 (N_14222,N_8251,N_8009);
nor U14223 (N_14223,N_10204,N_11822);
and U14224 (N_14224,N_9674,N_10331);
or U14225 (N_14225,N_8875,N_10150);
and U14226 (N_14226,N_11261,N_8653);
nand U14227 (N_14227,N_11448,N_10961);
xnor U14228 (N_14228,N_8220,N_11406);
and U14229 (N_14229,N_10051,N_8458);
and U14230 (N_14230,N_10381,N_9804);
xnor U14231 (N_14231,N_8313,N_9907);
and U14232 (N_14232,N_9777,N_10322);
nor U14233 (N_14233,N_10936,N_10026);
nor U14234 (N_14234,N_11686,N_9647);
and U14235 (N_14235,N_8677,N_10644);
and U14236 (N_14236,N_8038,N_9386);
or U14237 (N_14237,N_10940,N_9547);
or U14238 (N_14238,N_8160,N_8395);
nand U14239 (N_14239,N_9463,N_11879);
xor U14240 (N_14240,N_10312,N_9664);
xnor U14241 (N_14241,N_8901,N_11310);
nand U14242 (N_14242,N_9404,N_10129);
or U14243 (N_14243,N_10289,N_10345);
nor U14244 (N_14244,N_11684,N_10457);
nor U14245 (N_14245,N_11387,N_11692);
xor U14246 (N_14246,N_9654,N_9492);
nor U14247 (N_14247,N_9865,N_10517);
nand U14248 (N_14248,N_9489,N_11231);
nor U14249 (N_14249,N_10147,N_9118);
nor U14250 (N_14250,N_10616,N_8786);
nand U14251 (N_14251,N_9111,N_8803);
xor U14252 (N_14252,N_10228,N_8792);
xor U14253 (N_14253,N_8087,N_8412);
xor U14254 (N_14254,N_11368,N_9119);
nand U14255 (N_14255,N_8988,N_9380);
or U14256 (N_14256,N_8776,N_11335);
or U14257 (N_14257,N_8342,N_8598);
xnor U14258 (N_14258,N_8674,N_9017);
and U14259 (N_14259,N_9606,N_9564);
and U14260 (N_14260,N_8179,N_10656);
nand U14261 (N_14261,N_9725,N_11828);
xor U14262 (N_14262,N_11857,N_9441);
xnor U14263 (N_14263,N_9560,N_11656);
xnor U14264 (N_14264,N_11717,N_8233);
xor U14265 (N_14265,N_11846,N_11623);
and U14266 (N_14266,N_9277,N_11925);
xnor U14267 (N_14267,N_8655,N_10730);
nand U14268 (N_14268,N_9967,N_9046);
or U14269 (N_14269,N_10484,N_9293);
and U14270 (N_14270,N_10041,N_9864);
nand U14271 (N_14271,N_8948,N_9379);
nand U14272 (N_14272,N_8923,N_10939);
nand U14273 (N_14273,N_10209,N_11239);
nor U14274 (N_14274,N_11159,N_10184);
and U14275 (N_14275,N_10104,N_9237);
and U14276 (N_14276,N_11713,N_8645);
xor U14277 (N_14277,N_9097,N_10991);
or U14278 (N_14278,N_11786,N_10433);
and U14279 (N_14279,N_10696,N_11249);
nor U14280 (N_14280,N_8160,N_8418);
xor U14281 (N_14281,N_9702,N_10167);
and U14282 (N_14282,N_9829,N_8173);
xnor U14283 (N_14283,N_9054,N_9082);
and U14284 (N_14284,N_9680,N_11785);
and U14285 (N_14285,N_8990,N_9343);
xnor U14286 (N_14286,N_8732,N_10218);
or U14287 (N_14287,N_11835,N_9162);
xnor U14288 (N_14288,N_8419,N_8796);
nor U14289 (N_14289,N_8781,N_8483);
and U14290 (N_14290,N_9497,N_10005);
xnor U14291 (N_14291,N_9957,N_9874);
or U14292 (N_14292,N_8995,N_10130);
xnor U14293 (N_14293,N_11945,N_11476);
nor U14294 (N_14294,N_9853,N_11117);
or U14295 (N_14295,N_11276,N_11390);
or U14296 (N_14296,N_10436,N_11119);
nor U14297 (N_14297,N_10320,N_11595);
or U14298 (N_14298,N_9947,N_9864);
or U14299 (N_14299,N_11178,N_11007);
nand U14300 (N_14300,N_10284,N_8375);
nand U14301 (N_14301,N_10598,N_9387);
xnor U14302 (N_14302,N_10123,N_8731);
nor U14303 (N_14303,N_11232,N_10453);
nand U14304 (N_14304,N_11820,N_10697);
nand U14305 (N_14305,N_9250,N_8705);
nor U14306 (N_14306,N_8999,N_9431);
nand U14307 (N_14307,N_11934,N_10732);
nand U14308 (N_14308,N_10732,N_8581);
or U14309 (N_14309,N_9222,N_11680);
nand U14310 (N_14310,N_9373,N_9884);
xor U14311 (N_14311,N_9468,N_8882);
and U14312 (N_14312,N_10719,N_11016);
or U14313 (N_14313,N_9643,N_10034);
xor U14314 (N_14314,N_8976,N_10335);
xnor U14315 (N_14315,N_10772,N_8968);
nand U14316 (N_14316,N_11606,N_8293);
or U14317 (N_14317,N_10908,N_8096);
nand U14318 (N_14318,N_11044,N_9043);
nor U14319 (N_14319,N_11730,N_9957);
and U14320 (N_14320,N_11047,N_11135);
xnor U14321 (N_14321,N_9382,N_10647);
nor U14322 (N_14322,N_11697,N_10200);
xnor U14323 (N_14323,N_9198,N_11715);
or U14324 (N_14324,N_11243,N_11400);
nor U14325 (N_14325,N_9252,N_10237);
or U14326 (N_14326,N_11011,N_9394);
xnor U14327 (N_14327,N_8903,N_9814);
and U14328 (N_14328,N_9697,N_11996);
or U14329 (N_14329,N_11206,N_10433);
xor U14330 (N_14330,N_9606,N_10622);
or U14331 (N_14331,N_10619,N_9549);
nand U14332 (N_14332,N_8569,N_11661);
nor U14333 (N_14333,N_8617,N_10618);
or U14334 (N_14334,N_10494,N_9934);
or U14335 (N_14335,N_11442,N_8882);
xnor U14336 (N_14336,N_10489,N_9324);
and U14337 (N_14337,N_11750,N_8314);
xor U14338 (N_14338,N_8509,N_11152);
xnor U14339 (N_14339,N_10374,N_10378);
or U14340 (N_14340,N_9341,N_10788);
nand U14341 (N_14341,N_11103,N_11723);
nand U14342 (N_14342,N_11055,N_11048);
nand U14343 (N_14343,N_9583,N_8446);
and U14344 (N_14344,N_8969,N_9909);
and U14345 (N_14345,N_11635,N_8051);
nand U14346 (N_14346,N_11063,N_8515);
nand U14347 (N_14347,N_10075,N_11276);
or U14348 (N_14348,N_10409,N_10189);
nand U14349 (N_14349,N_10145,N_10361);
nor U14350 (N_14350,N_9760,N_9683);
and U14351 (N_14351,N_8360,N_9685);
or U14352 (N_14352,N_10696,N_9913);
and U14353 (N_14353,N_9113,N_9603);
xor U14354 (N_14354,N_10170,N_9506);
and U14355 (N_14355,N_8897,N_8016);
nor U14356 (N_14356,N_10773,N_8862);
and U14357 (N_14357,N_10646,N_8183);
or U14358 (N_14358,N_9571,N_10234);
nand U14359 (N_14359,N_10600,N_10760);
xnor U14360 (N_14360,N_9323,N_8148);
or U14361 (N_14361,N_11404,N_8753);
nand U14362 (N_14362,N_10242,N_9503);
or U14363 (N_14363,N_8814,N_11817);
xor U14364 (N_14364,N_8857,N_10322);
nand U14365 (N_14365,N_10262,N_10413);
nand U14366 (N_14366,N_9153,N_11669);
or U14367 (N_14367,N_10960,N_10741);
xor U14368 (N_14368,N_9119,N_10793);
nor U14369 (N_14369,N_8526,N_10956);
xnor U14370 (N_14370,N_8902,N_9630);
nor U14371 (N_14371,N_9850,N_8447);
nor U14372 (N_14372,N_9397,N_9015);
xor U14373 (N_14373,N_10096,N_8632);
and U14374 (N_14374,N_10374,N_10308);
nor U14375 (N_14375,N_10484,N_10898);
nor U14376 (N_14376,N_8343,N_9480);
and U14377 (N_14377,N_11896,N_8883);
nor U14378 (N_14378,N_11603,N_11865);
and U14379 (N_14379,N_9036,N_11920);
xnor U14380 (N_14380,N_10758,N_8158);
and U14381 (N_14381,N_9739,N_11970);
nand U14382 (N_14382,N_11061,N_8002);
and U14383 (N_14383,N_11617,N_9973);
and U14384 (N_14384,N_9977,N_9998);
and U14385 (N_14385,N_11613,N_11441);
xor U14386 (N_14386,N_10169,N_9259);
xnor U14387 (N_14387,N_9743,N_10279);
or U14388 (N_14388,N_9553,N_10811);
xnor U14389 (N_14389,N_9331,N_10292);
nand U14390 (N_14390,N_10715,N_8347);
xnor U14391 (N_14391,N_11809,N_10738);
and U14392 (N_14392,N_11085,N_9576);
xor U14393 (N_14393,N_11043,N_9556);
nor U14394 (N_14394,N_10671,N_9270);
xor U14395 (N_14395,N_8759,N_9966);
xnor U14396 (N_14396,N_9654,N_10930);
and U14397 (N_14397,N_8037,N_8036);
and U14398 (N_14398,N_9514,N_9681);
and U14399 (N_14399,N_9829,N_8888);
and U14400 (N_14400,N_9215,N_8124);
nand U14401 (N_14401,N_9568,N_8684);
nand U14402 (N_14402,N_8686,N_9035);
nand U14403 (N_14403,N_9602,N_10779);
and U14404 (N_14404,N_8655,N_11872);
nor U14405 (N_14405,N_10891,N_9314);
or U14406 (N_14406,N_10436,N_8027);
nor U14407 (N_14407,N_8052,N_9942);
or U14408 (N_14408,N_8184,N_11466);
nor U14409 (N_14409,N_11172,N_8075);
nand U14410 (N_14410,N_9494,N_10377);
or U14411 (N_14411,N_11045,N_8691);
nor U14412 (N_14412,N_11171,N_9528);
or U14413 (N_14413,N_10331,N_8570);
xor U14414 (N_14414,N_11215,N_11355);
or U14415 (N_14415,N_11264,N_8680);
or U14416 (N_14416,N_8142,N_10220);
and U14417 (N_14417,N_11047,N_9796);
or U14418 (N_14418,N_11182,N_9457);
and U14419 (N_14419,N_8713,N_8371);
nor U14420 (N_14420,N_8817,N_9589);
nand U14421 (N_14421,N_10883,N_10517);
or U14422 (N_14422,N_11033,N_9071);
nand U14423 (N_14423,N_8685,N_9648);
and U14424 (N_14424,N_9582,N_11883);
or U14425 (N_14425,N_9834,N_9608);
or U14426 (N_14426,N_9269,N_9876);
and U14427 (N_14427,N_10604,N_11907);
or U14428 (N_14428,N_8457,N_10846);
and U14429 (N_14429,N_11880,N_11637);
nand U14430 (N_14430,N_11877,N_10365);
xnor U14431 (N_14431,N_11729,N_11239);
or U14432 (N_14432,N_10318,N_9515);
xor U14433 (N_14433,N_11064,N_8323);
nand U14434 (N_14434,N_11937,N_8484);
xor U14435 (N_14435,N_8883,N_8216);
or U14436 (N_14436,N_11880,N_8965);
and U14437 (N_14437,N_10425,N_9947);
and U14438 (N_14438,N_8157,N_10004);
or U14439 (N_14439,N_8616,N_11190);
or U14440 (N_14440,N_8971,N_10054);
nor U14441 (N_14441,N_8703,N_10251);
or U14442 (N_14442,N_11552,N_8725);
nand U14443 (N_14443,N_11887,N_11659);
xor U14444 (N_14444,N_10646,N_11557);
and U14445 (N_14445,N_8776,N_10866);
nor U14446 (N_14446,N_11139,N_10697);
xor U14447 (N_14447,N_11712,N_10149);
nand U14448 (N_14448,N_10419,N_11662);
nor U14449 (N_14449,N_8926,N_8142);
nor U14450 (N_14450,N_8471,N_11217);
nor U14451 (N_14451,N_8661,N_10080);
xnor U14452 (N_14452,N_9870,N_11299);
and U14453 (N_14453,N_10970,N_11140);
and U14454 (N_14454,N_8352,N_8416);
nor U14455 (N_14455,N_9801,N_11924);
nor U14456 (N_14456,N_10333,N_11131);
nor U14457 (N_14457,N_9320,N_10583);
and U14458 (N_14458,N_11103,N_10633);
nor U14459 (N_14459,N_8529,N_8427);
xor U14460 (N_14460,N_10147,N_8212);
or U14461 (N_14461,N_11324,N_11696);
xnor U14462 (N_14462,N_11587,N_8660);
xor U14463 (N_14463,N_9060,N_11575);
nand U14464 (N_14464,N_9970,N_10951);
nor U14465 (N_14465,N_11061,N_10406);
or U14466 (N_14466,N_10218,N_11642);
and U14467 (N_14467,N_11482,N_10353);
nand U14468 (N_14468,N_9854,N_11443);
or U14469 (N_14469,N_11425,N_10452);
xor U14470 (N_14470,N_8249,N_11377);
nand U14471 (N_14471,N_10827,N_8920);
xor U14472 (N_14472,N_8192,N_11182);
xor U14473 (N_14473,N_8412,N_11463);
xnor U14474 (N_14474,N_9533,N_10244);
and U14475 (N_14475,N_9319,N_11875);
and U14476 (N_14476,N_9263,N_10743);
xor U14477 (N_14477,N_11061,N_8557);
and U14478 (N_14478,N_11659,N_8911);
nor U14479 (N_14479,N_8651,N_11179);
and U14480 (N_14480,N_11551,N_10870);
xor U14481 (N_14481,N_8807,N_11364);
xnor U14482 (N_14482,N_11462,N_8048);
or U14483 (N_14483,N_10662,N_9327);
nor U14484 (N_14484,N_10856,N_9463);
and U14485 (N_14485,N_11272,N_9109);
xor U14486 (N_14486,N_11570,N_9430);
xor U14487 (N_14487,N_9864,N_10578);
and U14488 (N_14488,N_9551,N_8098);
nand U14489 (N_14489,N_9496,N_9234);
nor U14490 (N_14490,N_11514,N_9176);
xnor U14491 (N_14491,N_9530,N_8340);
and U14492 (N_14492,N_8869,N_9580);
and U14493 (N_14493,N_8044,N_10602);
nand U14494 (N_14494,N_10119,N_8355);
or U14495 (N_14495,N_8145,N_8625);
and U14496 (N_14496,N_10383,N_8798);
xnor U14497 (N_14497,N_11803,N_10128);
and U14498 (N_14498,N_10224,N_10140);
nand U14499 (N_14499,N_10557,N_8818);
nand U14500 (N_14500,N_10004,N_10937);
and U14501 (N_14501,N_11665,N_11350);
xnor U14502 (N_14502,N_11162,N_10742);
and U14503 (N_14503,N_10124,N_8328);
nor U14504 (N_14504,N_10123,N_11746);
nor U14505 (N_14505,N_10137,N_8428);
nand U14506 (N_14506,N_8001,N_9718);
xnor U14507 (N_14507,N_10123,N_11111);
nor U14508 (N_14508,N_9695,N_8774);
nand U14509 (N_14509,N_8854,N_11628);
nor U14510 (N_14510,N_11116,N_11490);
and U14511 (N_14511,N_10932,N_9157);
or U14512 (N_14512,N_9298,N_9735);
nor U14513 (N_14513,N_10532,N_11696);
nand U14514 (N_14514,N_9983,N_11375);
nand U14515 (N_14515,N_10984,N_9210);
or U14516 (N_14516,N_11242,N_11528);
nand U14517 (N_14517,N_10426,N_8609);
xor U14518 (N_14518,N_8841,N_8719);
xnor U14519 (N_14519,N_9754,N_8326);
xnor U14520 (N_14520,N_8183,N_8475);
and U14521 (N_14521,N_9596,N_9390);
nor U14522 (N_14522,N_8327,N_10997);
xnor U14523 (N_14523,N_9164,N_10443);
nor U14524 (N_14524,N_10805,N_8359);
nor U14525 (N_14525,N_11363,N_8865);
or U14526 (N_14526,N_9090,N_9936);
nor U14527 (N_14527,N_11166,N_8016);
nor U14528 (N_14528,N_9764,N_11106);
nand U14529 (N_14529,N_11164,N_10874);
xnor U14530 (N_14530,N_9357,N_9238);
nor U14531 (N_14531,N_11052,N_9928);
or U14532 (N_14532,N_9762,N_8542);
and U14533 (N_14533,N_9842,N_8154);
or U14534 (N_14534,N_10124,N_9151);
xor U14535 (N_14535,N_11053,N_11272);
and U14536 (N_14536,N_9851,N_10028);
nor U14537 (N_14537,N_10983,N_9936);
and U14538 (N_14538,N_8760,N_10196);
nor U14539 (N_14539,N_11649,N_11492);
or U14540 (N_14540,N_10369,N_10792);
nor U14541 (N_14541,N_9281,N_9209);
nor U14542 (N_14542,N_11625,N_8465);
or U14543 (N_14543,N_10146,N_10107);
or U14544 (N_14544,N_9319,N_10402);
xnor U14545 (N_14545,N_11558,N_10243);
and U14546 (N_14546,N_10497,N_10793);
or U14547 (N_14547,N_8613,N_9687);
or U14548 (N_14548,N_8213,N_11462);
nand U14549 (N_14549,N_11538,N_10450);
xnor U14550 (N_14550,N_8198,N_10024);
and U14551 (N_14551,N_11366,N_10692);
nor U14552 (N_14552,N_9593,N_10745);
nand U14553 (N_14553,N_11981,N_9823);
nor U14554 (N_14554,N_8924,N_10503);
and U14555 (N_14555,N_8949,N_10139);
nor U14556 (N_14556,N_8830,N_8401);
nor U14557 (N_14557,N_9352,N_9645);
nor U14558 (N_14558,N_8075,N_8316);
xnor U14559 (N_14559,N_8867,N_11926);
or U14560 (N_14560,N_8258,N_11367);
nor U14561 (N_14561,N_10498,N_8141);
nand U14562 (N_14562,N_10433,N_10756);
and U14563 (N_14563,N_9361,N_9369);
or U14564 (N_14564,N_10100,N_9406);
nand U14565 (N_14565,N_11480,N_10631);
nand U14566 (N_14566,N_11614,N_11180);
and U14567 (N_14567,N_8141,N_8126);
and U14568 (N_14568,N_8194,N_11721);
nor U14569 (N_14569,N_10500,N_8326);
xnor U14570 (N_14570,N_10936,N_10138);
xnor U14571 (N_14571,N_10027,N_10258);
xor U14572 (N_14572,N_11545,N_8118);
xor U14573 (N_14573,N_8853,N_9742);
nor U14574 (N_14574,N_8541,N_8967);
xor U14575 (N_14575,N_11007,N_8150);
or U14576 (N_14576,N_11596,N_8266);
nand U14577 (N_14577,N_9179,N_8447);
nor U14578 (N_14578,N_10781,N_11988);
or U14579 (N_14579,N_10496,N_9005);
nor U14580 (N_14580,N_11864,N_10680);
xor U14581 (N_14581,N_10833,N_8736);
nor U14582 (N_14582,N_10718,N_11411);
and U14583 (N_14583,N_10287,N_11426);
nor U14584 (N_14584,N_10921,N_9113);
xnor U14585 (N_14585,N_10662,N_11903);
nand U14586 (N_14586,N_9475,N_10862);
nor U14587 (N_14587,N_11114,N_11833);
nand U14588 (N_14588,N_9935,N_10234);
nor U14589 (N_14589,N_8363,N_11640);
nor U14590 (N_14590,N_10497,N_11733);
nand U14591 (N_14591,N_10610,N_11124);
and U14592 (N_14592,N_8231,N_8003);
and U14593 (N_14593,N_11520,N_10053);
xnor U14594 (N_14594,N_11748,N_11901);
xnor U14595 (N_14595,N_8581,N_9426);
or U14596 (N_14596,N_9670,N_8295);
or U14597 (N_14597,N_9253,N_8906);
nand U14598 (N_14598,N_8706,N_11478);
and U14599 (N_14599,N_10281,N_9095);
and U14600 (N_14600,N_10145,N_9126);
nand U14601 (N_14601,N_10868,N_10531);
and U14602 (N_14602,N_9281,N_8254);
nor U14603 (N_14603,N_10405,N_11182);
and U14604 (N_14604,N_8477,N_10306);
xor U14605 (N_14605,N_10402,N_8725);
and U14606 (N_14606,N_8653,N_9314);
xnor U14607 (N_14607,N_9921,N_8415);
and U14608 (N_14608,N_8890,N_11676);
nor U14609 (N_14609,N_9022,N_9410);
and U14610 (N_14610,N_11763,N_10456);
nor U14611 (N_14611,N_10107,N_9552);
or U14612 (N_14612,N_9488,N_10187);
or U14613 (N_14613,N_11035,N_11259);
and U14614 (N_14614,N_10288,N_8809);
nand U14615 (N_14615,N_8842,N_10202);
nand U14616 (N_14616,N_11262,N_8540);
nor U14617 (N_14617,N_11240,N_10652);
or U14618 (N_14618,N_9919,N_11579);
and U14619 (N_14619,N_11742,N_8084);
or U14620 (N_14620,N_10177,N_9075);
nor U14621 (N_14621,N_8267,N_10796);
or U14622 (N_14622,N_10058,N_10919);
xnor U14623 (N_14623,N_8782,N_9109);
or U14624 (N_14624,N_11751,N_9984);
nand U14625 (N_14625,N_9589,N_8356);
and U14626 (N_14626,N_9537,N_9094);
or U14627 (N_14627,N_8256,N_11275);
nand U14628 (N_14628,N_10670,N_8488);
nor U14629 (N_14629,N_11417,N_8910);
xnor U14630 (N_14630,N_11632,N_11353);
and U14631 (N_14631,N_8269,N_10290);
nor U14632 (N_14632,N_10681,N_11806);
nand U14633 (N_14633,N_10836,N_9794);
and U14634 (N_14634,N_9459,N_8866);
nand U14635 (N_14635,N_10967,N_10457);
and U14636 (N_14636,N_11094,N_11622);
nand U14637 (N_14637,N_10153,N_8149);
or U14638 (N_14638,N_10521,N_11712);
nand U14639 (N_14639,N_8998,N_8367);
or U14640 (N_14640,N_9137,N_10073);
xor U14641 (N_14641,N_10485,N_10956);
or U14642 (N_14642,N_9164,N_8222);
and U14643 (N_14643,N_10729,N_9475);
and U14644 (N_14644,N_9900,N_10559);
nand U14645 (N_14645,N_9974,N_9636);
and U14646 (N_14646,N_10260,N_8448);
nor U14647 (N_14647,N_9617,N_10335);
nand U14648 (N_14648,N_9637,N_9063);
nand U14649 (N_14649,N_8144,N_11655);
nor U14650 (N_14650,N_11544,N_9097);
nand U14651 (N_14651,N_11600,N_11117);
or U14652 (N_14652,N_9668,N_10178);
nand U14653 (N_14653,N_11543,N_10804);
or U14654 (N_14654,N_9081,N_8959);
nor U14655 (N_14655,N_8877,N_10933);
or U14656 (N_14656,N_11049,N_10494);
xnor U14657 (N_14657,N_8179,N_8049);
nor U14658 (N_14658,N_8042,N_10070);
nor U14659 (N_14659,N_10409,N_8503);
nand U14660 (N_14660,N_8925,N_11198);
or U14661 (N_14661,N_11250,N_9137);
xnor U14662 (N_14662,N_9668,N_9329);
and U14663 (N_14663,N_11182,N_11606);
nand U14664 (N_14664,N_10597,N_8164);
nand U14665 (N_14665,N_10111,N_10991);
nor U14666 (N_14666,N_10089,N_8267);
or U14667 (N_14667,N_8153,N_8411);
and U14668 (N_14668,N_9886,N_8041);
nor U14669 (N_14669,N_8331,N_11806);
xor U14670 (N_14670,N_9386,N_11750);
nand U14671 (N_14671,N_9134,N_9540);
xnor U14672 (N_14672,N_10051,N_9442);
xor U14673 (N_14673,N_10261,N_11675);
nand U14674 (N_14674,N_9292,N_10084);
nor U14675 (N_14675,N_11316,N_8538);
xor U14676 (N_14676,N_11481,N_9889);
or U14677 (N_14677,N_8173,N_9437);
nand U14678 (N_14678,N_11048,N_11231);
nand U14679 (N_14679,N_8956,N_10969);
xnor U14680 (N_14680,N_10049,N_10968);
and U14681 (N_14681,N_11724,N_10186);
xor U14682 (N_14682,N_8760,N_9048);
and U14683 (N_14683,N_9130,N_9937);
or U14684 (N_14684,N_9554,N_9821);
and U14685 (N_14685,N_9550,N_10411);
xor U14686 (N_14686,N_8337,N_8973);
xnor U14687 (N_14687,N_9931,N_10735);
or U14688 (N_14688,N_10879,N_9524);
or U14689 (N_14689,N_9881,N_8866);
nor U14690 (N_14690,N_10398,N_10683);
xnor U14691 (N_14691,N_9955,N_8936);
or U14692 (N_14692,N_9242,N_8514);
or U14693 (N_14693,N_11931,N_9763);
and U14694 (N_14694,N_8402,N_9382);
nor U14695 (N_14695,N_8256,N_11180);
nand U14696 (N_14696,N_9733,N_9147);
and U14697 (N_14697,N_9461,N_10657);
and U14698 (N_14698,N_11548,N_8509);
xor U14699 (N_14699,N_11045,N_11922);
nand U14700 (N_14700,N_9845,N_8120);
and U14701 (N_14701,N_10699,N_9856);
and U14702 (N_14702,N_8340,N_10194);
xor U14703 (N_14703,N_9201,N_9807);
and U14704 (N_14704,N_9344,N_10981);
nor U14705 (N_14705,N_8222,N_11821);
xnor U14706 (N_14706,N_10770,N_10908);
xnor U14707 (N_14707,N_11674,N_9514);
xor U14708 (N_14708,N_8506,N_9509);
nor U14709 (N_14709,N_8367,N_10594);
or U14710 (N_14710,N_10742,N_11446);
or U14711 (N_14711,N_11310,N_11173);
and U14712 (N_14712,N_9956,N_8949);
and U14713 (N_14713,N_10471,N_10937);
nor U14714 (N_14714,N_10185,N_11965);
nand U14715 (N_14715,N_11327,N_8034);
nor U14716 (N_14716,N_8449,N_11924);
or U14717 (N_14717,N_11792,N_11485);
nor U14718 (N_14718,N_11369,N_10902);
or U14719 (N_14719,N_10384,N_11041);
xnor U14720 (N_14720,N_11260,N_11008);
xnor U14721 (N_14721,N_8561,N_9551);
or U14722 (N_14722,N_9629,N_8500);
or U14723 (N_14723,N_9676,N_9202);
xor U14724 (N_14724,N_9062,N_10221);
xor U14725 (N_14725,N_8614,N_10410);
nand U14726 (N_14726,N_10283,N_9541);
or U14727 (N_14727,N_9197,N_9589);
and U14728 (N_14728,N_10198,N_8003);
xnor U14729 (N_14729,N_10954,N_10246);
nor U14730 (N_14730,N_11066,N_9539);
xor U14731 (N_14731,N_8578,N_9229);
xnor U14732 (N_14732,N_11313,N_9130);
xor U14733 (N_14733,N_10993,N_11613);
or U14734 (N_14734,N_9797,N_9851);
nor U14735 (N_14735,N_10830,N_11585);
nor U14736 (N_14736,N_10509,N_8328);
and U14737 (N_14737,N_10965,N_10658);
and U14738 (N_14738,N_9859,N_9093);
and U14739 (N_14739,N_11227,N_9824);
nand U14740 (N_14740,N_10843,N_9039);
and U14741 (N_14741,N_10241,N_9344);
nor U14742 (N_14742,N_9211,N_11319);
nor U14743 (N_14743,N_9492,N_9247);
or U14744 (N_14744,N_10618,N_9483);
xnor U14745 (N_14745,N_10847,N_8790);
xor U14746 (N_14746,N_8762,N_8410);
nor U14747 (N_14747,N_11988,N_10793);
or U14748 (N_14748,N_9060,N_11155);
nand U14749 (N_14749,N_8523,N_9502);
nor U14750 (N_14750,N_9119,N_9756);
xnor U14751 (N_14751,N_10038,N_8654);
xor U14752 (N_14752,N_11015,N_10840);
nand U14753 (N_14753,N_10789,N_10529);
nand U14754 (N_14754,N_8350,N_9483);
xor U14755 (N_14755,N_9325,N_11728);
and U14756 (N_14756,N_9799,N_9633);
nand U14757 (N_14757,N_8992,N_10161);
or U14758 (N_14758,N_11534,N_9062);
xor U14759 (N_14759,N_9277,N_11332);
xnor U14760 (N_14760,N_9569,N_8579);
nor U14761 (N_14761,N_9420,N_8190);
nand U14762 (N_14762,N_9582,N_9297);
xnor U14763 (N_14763,N_11546,N_8662);
or U14764 (N_14764,N_11108,N_11360);
or U14765 (N_14765,N_8706,N_8825);
nor U14766 (N_14766,N_9394,N_9736);
or U14767 (N_14767,N_9189,N_9213);
and U14768 (N_14768,N_10315,N_8542);
nor U14769 (N_14769,N_10583,N_8661);
and U14770 (N_14770,N_11743,N_10022);
nand U14771 (N_14771,N_10597,N_9808);
nand U14772 (N_14772,N_8330,N_9347);
and U14773 (N_14773,N_8003,N_9874);
xor U14774 (N_14774,N_9938,N_8057);
xnor U14775 (N_14775,N_10609,N_11208);
nor U14776 (N_14776,N_11432,N_8898);
xor U14777 (N_14777,N_8498,N_9964);
nor U14778 (N_14778,N_11688,N_11644);
nor U14779 (N_14779,N_8106,N_9123);
and U14780 (N_14780,N_8405,N_9246);
nand U14781 (N_14781,N_10014,N_10689);
nor U14782 (N_14782,N_11695,N_9361);
or U14783 (N_14783,N_9907,N_10890);
nand U14784 (N_14784,N_10565,N_9266);
or U14785 (N_14785,N_10986,N_9416);
or U14786 (N_14786,N_8506,N_8732);
xor U14787 (N_14787,N_8587,N_9118);
nand U14788 (N_14788,N_9800,N_8150);
nand U14789 (N_14789,N_9938,N_9275);
and U14790 (N_14790,N_11423,N_8296);
nand U14791 (N_14791,N_8802,N_8789);
and U14792 (N_14792,N_10692,N_11477);
nor U14793 (N_14793,N_8001,N_9373);
nor U14794 (N_14794,N_10328,N_10502);
and U14795 (N_14795,N_9830,N_10068);
and U14796 (N_14796,N_9058,N_9768);
nand U14797 (N_14797,N_10795,N_11106);
nand U14798 (N_14798,N_8480,N_8923);
nand U14799 (N_14799,N_8007,N_8369);
nand U14800 (N_14800,N_10817,N_10512);
nand U14801 (N_14801,N_11899,N_9655);
xor U14802 (N_14802,N_8025,N_11893);
nor U14803 (N_14803,N_11625,N_8207);
xor U14804 (N_14804,N_9817,N_8978);
or U14805 (N_14805,N_11033,N_11806);
xor U14806 (N_14806,N_8596,N_9871);
and U14807 (N_14807,N_10890,N_8994);
and U14808 (N_14808,N_11753,N_11908);
or U14809 (N_14809,N_9017,N_11357);
or U14810 (N_14810,N_9292,N_8369);
nor U14811 (N_14811,N_9698,N_11231);
and U14812 (N_14812,N_9431,N_9821);
nor U14813 (N_14813,N_9818,N_8545);
or U14814 (N_14814,N_8762,N_8315);
nor U14815 (N_14815,N_8811,N_10353);
nor U14816 (N_14816,N_8064,N_8737);
nor U14817 (N_14817,N_9121,N_9802);
or U14818 (N_14818,N_9723,N_10208);
or U14819 (N_14819,N_10129,N_11098);
xor U14820 (N_14820,N_10665,N_11712);
nand U14821 (N_14821,N_8559,N_10751);
or U14822 (N_14822,N_10816,N_8574);
and U14823 (N_14823,N_8886,N_11108);
or U14824 (N_14824,N_11705,N_11413);
nor U14825 (N_14825,N_11833,N_11932);
or U14826 (N_14826,N_11941,N_8957);
xnor U14827 (N_14827,N_11540,N_8964);
and U14828 (N_14828,N_9417,N_10354);
nand U14829 (N_14829,N_11130,N_10056);
nor U14830 (N_14830,N_11177,N_11995);
and U14831 (N_14831,N_10369,N_10022);
or U14832 (N_14832,N_10979,N_11315);
nor U14833 (N_14833,N_10611,N_10357);
xor U14834 (N_14834,N_10288,N_9449);
nor U14835 (N_14835,N_10989,N_8528);
and U14836 (N_14836,N_11871,N_8344);
xnor U14837 (N_14837,N_8324,N_9297);
nand U14838 (N_14838,N_11832,N_11905);
or U14839 (N_14839,N_9303,N_9912);
and U14840 (N_14840,N_8192,N_11507);
nand U14841 (N_14841,N_9024,N_11982);
nand U14842 (N_14842,N_8298,N_11884);
nand U14843 (N_14843,N_8085,N_11737);
nand U14844 (N_14844,N_10510,N_11484);
and U14845 (N_14845,N_10544,N_11723);
or U14846 (N_14846,N_11468,N_9264);
and U14847 (N_14847,N_8068,N_10051);
nor U14848 (N_14848,N_9051,N_9982);
nor U14849 (N_14849,N_8813,N_10607);
xor U14850 (N_14850,N_11541,N_9980);
nand U14851 (N_14851,N_10116,N_10480);
xor U14852 (N_14852,N_11497,N_11148);
nor U14853 (N_14853,N_9202,N_8229);
nor U14854 (N_14854,N_8724,N_10167);
or U14855 (N_14855,N_9313,N_9203);
nand U14856 (N_14856,N_11732,N_8950);
or U14857 (N_14857,N_10769,N_11433);
and U14858 (N_14858,N_10936,N_10604);
or U14859 (N_14859,N_9970,N_9545);
xor U14860 (N_14860,N_9001,N_11380);
nand U14861 (N_14861,N_11919,N_9382);
and U14862 (N_14862,N_11316,N_8151);
nor U14863 (N_14863,N_9979,N_8155);
and U14864 (N_14864,N_9445,N_10410);
and U14865 (N_14865,N_11812,N_11846);
and U14866 (N_14866,N_9607,N_10225);
xor U14867 (N_14867,N_10168,N_11648);
nand U14868 (N_14868,N_9792,N_9292);
nor U14869 (N_14869,N_10176,N_10253);
xor U14870 (N_14870,N_10480,N_10785);
nand U14871 (N_14871,N_9658,N_11100);
xnor U14872 (N_14872,N_11975,N_10500);
and U14873 (N_14873,N_10752,N_11537);
nor U14874 (N_14874,N_11915,N_9998);
nand U14875 (N_14875,N_10381,N_9428);
nor U14876 (N_14876,N_9438,N_8836);
or U14877 (N_14877,N_10542,N_11408);
and U14878 (N_14878,N_9115,N_9795);
or U14879 (N_14879,N_10691,N_10436);
nand U14880 (N_14880,N_8098,N_10132);
xor U14881 (N_14881,N_11793,N_10153);
nor U14882 (N_14882,N_10977,N_10127);
or U14883 (N_14883,N_10923,N_11880);
nor U14884 (N_14884,N_8918,N_9738);
and U14885 (N_14885,N_8878,N_8439);
and U14886 (N_14886,N_8390,N_11650);
or U14887 (N_14887,N_9461,N_9039);
xnor U14888 (N_14888,N_11739,N_10120);
xor U14889 (N_14889,N_8801,N_8412);
and U14890 (N_14890,N_11413,N_8463);
and U14891 (N_14891,N_11813,N_10298);
and U14892 (N_14892,N_9574,N_11200);
or U14893 (N_14893,N_9402,N_9455);
and U14894 (N_14894,N_11106,N_10647);
nor U14895 (N_14895,N_9403,N_10197);
and U14896 (N_14896,N_11433,N_11030);
nor U14897 (N_14897,N_11119,N_9543);
nand U14898 (N_14898,N_8496,N_11729);
nand U14899 (N_14899,N_9135,N_11885);
nand U14900 (N_14900,N_9392,N_11724);
xor U14901 (N_14901,N_9541,N_9627);
nand U14902 (N_14902,N_10024,N_8510);
xor U14903 (N_14903,N_9275,N_8878);
or U14904 (N_14904,N_9663,N_8137);
xnor U14905 (N_14905,N_9334,N_9564);
nand U14906 (N_14906,N_10090,N_10551);
and U14907 (N_14907,N_8697,N_10216);
and U14908 (N_14908,N_9626,N_9400);
or U14909 (N_14909,N_9927,N_9926);
or U14910 (N_14910,N_8404,N_11325);
nor U14911 (N_14911,N_11075,N_9812);
or U14912 (N_14912,N_11641,N_8667);
xor U14913 (N_14913,N_10034,N_9957);
nor U14914 (N_14914,N_10782,N_11893);
xnor U14915 (N_14915,N_11655,N_10995);
nand U14916 (N_14916,N_10152,N_8511);
nor U14917 (N_14917,N_8266,N_8740);
nor U14918 (N_14918,N_11090,N_8707);
nand U14919 (N_14919,N_10604,N_10677);
nand U14920 (N_14920,N_8347,N_11218);
and U14921 (N_14921,N_10327,N_8080);
or U14922 (N_14922,N_9012,N_8641);
and U14923 (N_14923,N_9185,N_11526);
xnor U14924 (N_14924,N_8599,N_10054);
nor U14925 (N_14925,N_10413,N_9762);
nand U14926 (N_14926,N_8946,N_10425);
nor U14927 (N_14927,N_11226,N_10453);
nand U14928 (N_14928,N_8177,N_10804);
nand U14929 (N_14929,N_8090,N_11699);
or U14930 (N_14930,N_9371,N_11860);
or U14931 (N_14931,N_9071,N_11464);
and U14932 (N_14932,N_8504,N_8077);
or U14933 (N_14933,N_8585,N_11360);
or U14934 (N_14934,N_10089,N_9586);
nand U14935 (N_14935,N_11874,N_9970);
nor U14936 (N_14936,N_9988,N_8527);
or U14937 (N_14937,N_11806,N_11681);
nor U14938 (N_14938,N_11736,N_9166);
or U14939 (N_14939,N_10810,N_10125);
or U14940 (N_14940,N_10634,N_11784);
or U14941 (N_14941,N_8298,N_10544);
xor U14942 (N_14942,N_8251,N_8245);
xnor U14943 (N_14943,N_11661,N_11059);
or U14944 (N_14944,N_10095,N_10019);
and U14945 (N_14945,N_10199,N_11724);
or U14946 (N_14946,N_11533,N_8306);
xnor U14947 (N_14947,N_8428,N_11032);
and U14948 (N_14948,N_11971,N_8259);
and U14949 (N_14949,N_8310,N_8954);
nand U14950 (N_14950,N_8037,N_9063);
or U14951 (N_14951,N_11668,N_10053);
nor U14952 (N_14952,N_10789,N_9967);
nor U14953 (N_14953,N_10551,N_10361);
and U14954 (N_14954,N_10199,N_11424);
xor U14955 (N_14955,N_9198,N_9999);
or U14956 (N_14956,N_11815,N_8712);
nor U14957 (N_14957,N_9571,N_10544);
or U14958 (N_14958,N_10911,N_8072);
and U14959 (N_14959,N_9384,N_10520);
or U14960 (N_14960,N_9469,N_8724);
nand U14961 (N_14961,N_10140,N_10335);
or U14962 (N_14962,N_11457,N_10634);
nor U14963 (N_14963,N_10663,N_8782);
nand U14964 (N_14964,N_8702,N_10907);
nor U14965 (N_14965,N_10484,N_9710);
and U14966 (N_14966,N_8953,N_10189);
nor U14967 (N_14967,N_8676,N_11407);
and U14968 (N_14968,N_10663,N_10282);
xor U14969 (N_14969,N_9246,N_10823);
xnor U14970 (N_14970,N_8078,N_11358);
or U14971 (N_14971,N_8747,N_9354);
nand U14972 (N_14972,N_11403,N_9149);
or U14973 (N_14973,N_8956,N_8466);
nor U14974 (N_14974,N_9128,N_10354);
xor U14975 (N_14975,N_11036,N_9545);
nand U14976 (N_14976,N_11593,N_11274);
nand U14977 (N_14977,N_9356,N_9849);
nor U14978 (N_14978,N_11954,N_11842);
or U14979 (N_14979,N_10907,N_10458);
and U14980 (N_14980,N_9605,N_11303);
and U14981 (N_14981,N_11936,N_9652);
and U14982 (N_14982,N_8413,N_8894);
and U14983 (N_14983,N_8855,N_9056);
xnor U14984 (N_14984,N_11766,N_11784);
or U14985 (N_14985,N_10588,N_10874);
nand U14986 (N_14986,N_8324,N_10058);
nand U14987 (N_14987,N_9605,N_9814);
or U14988 (N_14988,N_11147,N_10213);
nand U14989 (N_14989,N_10560,N_8754);
nor U14990 (N_14990,N_11157,N_8256);
nor U14991 (N_14991,N_10033,N_9099);
and U14992 (N_14992,N_9393,N_11719);
nand U14993 (N_14993,N_8453,N_11398);
and U14994 (N_14994,N_9319,N_9133);
nand U14995 (N_14995,N_8631,N_10436);
nand U14996 (N_14996,N_8444,N_11860);
nand U14997 (N_14997,N_11042,N_9922);
xor U14998 (N_14998,N_10133,N_10662);
or U14999 (N_14999,N_9814,N_10533);
nand U15000 (N_15000,N_11815,N_8119);
and U15001 (N_15001,N_9618,N_9136);
xor U15002 (N_15002,N_10476,N_9461);
or U15003 (N_15003,N_8447,N_9933);
xnor U15004 (N_15004,N_10293,N_10582);
nor U15005 (N_15005,N_10413,N_10759);
and U15006 (N_15006,N_9472,N_9884);
nor U15007 (N_15007,N_8235,N_10514);
and U15008 (N_15008,N_9856,N_9328);
nand U15009 (N_15009,N_10224,N_9593);
and U15010 (N_15010,N_11694,N_8756);
xor U15011 (N_15011,N_9788,N_11897);
xnor U15012 (N_15012,N_11216,N_10916);
and U15013 (N_15013,N_8838,N_10050);
or U15014 (N_15014,N_8461,N_10273);
or U15015 (N_15015,N_10485,N_11957);
or U15016 (N_15016,N_10382,N_10208);
and U15017 (N_15017,N_10841,N_11669);
and U15018 (N_15018,N_9442,N_9759);
or U15019 (N_15019,N_10010,N_8352);
nand U15020 (N_15020,N_11481,N_11409);
or U15021 (N_15021,N_8890,N_11373);
nor U15022 (N_15022,N_9655,N_11329);
and U15023 (N_15023,N_9122,N_9609);
nor U15024 (N_15024,N_11638,N_9683);
nand U15025 (N_15025,N_9886,N_9235);
xor U15026 (N_15026,N_9129,N_10509);
or U15027 (N_15027,N_11571,N_9037);
and U15028 (N_15028,N_11929,N_10329);
or U15029 (N_15029,N_9293,N_10432);
and U15030 (N_15030,N_8323,N_10985);
nand U15031 (N_15031,N_11832,N_9728);
or U15032 (N_15032,N_10333,N_11954);
or U15033 (N_15033,N_10360,N_8757);
nand U15034 (N_15034,N_11761,N_8397);
nand U15035 (N_15035,N_9568,N_11567);
or U15036 (N_15036,N_11246,N_9773);
nor U15037 (N_15037,N_11054,N_11578);
and U15038 (N_15038,N_10457,N_8459);
or U15039 (N_15039,N_11194,N_9549);
nor U15040 (N_15040,N_10676,N_9879);
xnor U15041 (N_15041,N_10154,N_10006);
xor U15042 (N_15042,N_9473,N_11493);
xor U15043 (N_15043,N_8918,N_9458);
nor U15044 (N_15044,N_9403,N_9287);
xor U15045 (N_15045,N_11419,N_8617);
xnor U15046 (N_15046,N_8732,N_8885);
or U15047 (N_15047,N_10501,N_10567);
nor U15048 (N_15048,N_11157,N_11425);
nor U15049 (N_15049,N_9991,N_10126);
nor U15050 (N_15050,N_11043,N_11160);
nor U15051 (N_15051,N_10329,N_10909);
xor U15052 (N_15052,N_11428,N_10726);
or U15053 (N_15053,N_8571,N_8347);
and U15054 (N_15054,N_11658,N_8879);
xor U15055 (N_15055,N_11451,N_10698);
xor U15056 (N_15056,N_9995,N_11975);
nor U15057 (N_15057,N_8537,N_11966);
nand U15058 (N_15058,N_10817,N_10019);
nand U15059 (N_15059,N_11424,N_8948);
or U15060 (N_15060,N_8052,N_11454);
nand U15061 (N_15061,N_11423,N_8465);
xor U15062 (N_15062,N_9101,N_11107);
xnor U15063 (N_15063,N_11274,N_10502);
nand U15064 (N_15064,N_8146,N_11025);
xor U15065 (N_15065,N_11721,N_11161);
nor U15066 (N_15066,N_9221,N_8975);
or U15067 (N_15067,N_10026,N_11586);
or U15068 (N_15068,N_8450,N_10753);
or U15069 (N_15069,N_9797,N_9388);
and U15070 (N_15070,N_9043,N_10050);
nand U15071 (N_15071,N_8947,N_8892);
xnor U15072 (N_15072,N_10189,N_8495);
or U15073 (N_15073,N_10205,N_9984);
nor U15074 (N_15074,N_10312,N_9145);
or U15075 (N_15075,N_8035,N_9430);
nor U15076 (N_15076,N_8280,N_9684);
nand U15077 (N_15077,N_11322,N_8084);
xor U15078 (N_15078,N_9949,N_11703);
nand U15079 (N_15079,N_9826,N_8684);
or U15080 (N_15080,N_8080,N_11535);
nand U15081 (N_15081,N_9180,N_11646);
or U15082 (N_15082,N_9673,N_8834);
nand U15083 (N_15083,N_10104,N_11332);
or U15084 (N_15084,N_9553,N_8954);
or U15085 (N_15085,N_10823,N_11664);
xor U15086 (N_15086,N_9570,N_10372);
nor U15087 (N_15087,N_9082,N_10533);
or U15088 (N_15088,N_8848,N_9408);
and U15089 (N_15089,N_9812,N_11622);
nand U15090 (N_15090,N_11773,N_9044);
or U15091 (N_15091,N_10288,N_10908);
xor U15092 (N_15092,N_10596,N_8605);
nand U15093 (N_15093,N_8622,N_8919);
or U15094 (N_15094,N_8357,N_11666);
nand U15095 (N_15095,N_9452,N_11880);
or U15096 (N_15096,N_10374,N_9482);
or U15097 (N_15097,N_8414,N_8848);
or U15098 (N_15098,N_11743,N_8789);
or U15099 (N_15099,N_11983,N_9457);
nand U15100 (N_15100,N_9512,N_8361);
or U15101 (N_15101,N_11972,N_10111);
nor U15102 (N_15102,N_9981,N_9499);
nor U15103 (N_15103,N_10020,N_10035);
nand U15104 (N_15104,N_9846,N_11826);
and U15105 (N_15105,N_11014,N_8670);
nand U15106 (N_15106,N_9409,N_8855);
or U15107 (N_15107,N_9394,N_9052);
xnor U15108 (N_15108,N_11681,N_9731);
or U15109 (N_15109,N_11691,N_11706);
or U15110 (N_15110,N_9152,N_8918);
xor U15111 (N_15111,N_8583,N_8174);
nand U15112 (N_15112,N_11917,N_8205);
nand U15113 (N_15113,N_9160,N_11214);
nor U15114 (N_15114,N_8081,N_11470);
xor U15115 (N_15115,N_8092,N_8809);
xor U15116 (N_15116,N_9078,N_11952);
xnor U15117 (N_15117,N_11215,N_10184);
xnor U15118 (N_15118,N_10418,N_9861);
and U15119 (N_15119,N_9083,N_9605);
or U15120 (N_15120,N_11434,N_8542);
nand U15121 (N_15121,N_10675,N_11123);
nor U15122 (N_15122,N_9898,N_8331);
nor U15123 (N_15123,N_11908,N_9537);
or U15124 (N_15124,N_9303,N_8576);
and U15125 (N_15125,N_11420,N_8028);
nor U15126 (N_15126,N_11331,N_8152);
and U15127 (N_15127,N_10934,N_11176);
nand U15128 (N_15128,N_11786,N_9943);
nor U15129 (N_15129,N_11863,N_11263);
or U15130 (N_15130,N_9107,N_8027);
and U15131 (N_15131,N_10426,N_9392);
nor U15132 (N_15132,N_8061,N_9858);
xor U15133 (N_15133,N_10562,N_8123);
xnor U15134 (N_15134,N_8369,N_8560);
and U15135 (N_15135,N_10070,N_11053);
or U15136 (N_15136,N_11835,N_8472);
and U15137 (N_15137,N_8299,N_11590);
nand U15138 (N_15138,N_10664,N_10366);
xnor U15139 (N_15139,N_8335,N_8900);
nand U15140 (N_15140,N_11150,N_8359);
xnor U15141 (N_15141,N_8987,N_9428);
nand U15142 (N_15142,N_8295,N_9188);
or U15143 (N_15143,N_9427,N_10907);
and U15144 (N_15144,N_11307,N_11778);
nand U15145 (N_15145,N_9939,N_11868);
xor U15146 (N_15146,N_8258,N_11620);
xnor U15147 (N_15147,N_11573,N_8752);
nor U15148 (N_15148,N_9260,N_8329);
nor U15149 (N_15149,N_8505,N_8789);
or U15150 (N_15150,N_10578,N_10401);
and U15151 (N_15151,N_10552,N_8108);
and U15152 (N_15152,N_11807,N_10446);
nor U15153 (N_15153,N_10345,N_11968);
and U15154 (N_15154,N_8145,N_11686);
nand U15155 (N_15155,N_10528,N_9550);
xnor U15156 (N_15156,N_8921,N_9491);
xnor U15157 (N_15157,N_11490,N_8044);
or U15158 (N_15158,N_11867,N_11789);
and U15159 (N_15159,N_8609,N_9129);
nor U15160 (N_15160,N_10517,N_9190);
nand U15161 (N_15161,N_9682,N_9556);
or U15162 (N_15162,N_10608,N_11524);
nand U15163 (N_15163,N_10636,N_9763);
nor U15164 (N_15164,N_9432,N_11641);
nor U15165 (N_15165,N_9876,N_11865);
and U15166 (N_15166,N_10853,N_8389);
nor U15167 (N_15167,N_11723,N_10548);
xnor U15168 (N_15168,N_8738,N_8663);
and U15169 (N_15169,N_11768,N_10124);
or U15170 (N_15170,N_9762,N_11810);
and U15171 (N_15171,N_10678,N_8180);
and U15172 (N_15172,N_9880,N_11500);
xor U15173 (N_15173,N_8590,N_8057);
nor U15174 (N_15174,N_11758,N_11880);
or U15175 (N_15175,N_9607,N_10353);
xnor U15176 (N_15176,N_8111,N_11629);
nand U15177 (N_15177,N_10416,N_9387);
xor U15178 (N_15178,N_9363,N_11989);
or U15179 (N_15179,N_9330,N_10745);
nand U15180 (N_15180,N_10905,N_9125);
nor U15181 (N_15181,N_9791,N_9398);
or U15182 (N_15182,N_11037,N_10614);
and U15183 (N_15183,N_11530,N_10081);
xnor U15184 (N_15184,N_9529,N_9948);
nand U15185 (N_15185,N_8047,N_9473);
xnor U15186 (N_15186,N_9916,N_8904);
xor U15187 (N_15187,N_10595,N_10289);
and U15188 (N_15188,N_9094,N_8696);
nand U15189 (N_15189,N_9862,N_8855);
xor U15190 (N_15190,N_11299,N_9143);
nand U15191 (N_15191,N_10763,N_11272);
nor U15192 (N_15192,N_8451,N_11874);
xnor U15193 (N_15193,N_11618,N_8473);
and U15194 (N_15194,N_8271,N_10109);
or U15195 (N_15195,N_9932,N_9066);
xnor U15196 (N_15196,N_8371,N_11818);
or U15197 (N_15197,N_11511,N_10489);
nand U15198 (N_15198,N_11296,N_9814);
xnor U15199 (N_15199,N_11296,N_11246);
nand U15200 (N_15200,N_8268,N_10926);
and U15201 (N_15201,N_10134,N_8436);
nor U15202 (N_15202,N_9885,N_11915);
nand U15203 (N_15203,N_9228,N_10707);
xor U15204 (N_15204,N_9188,N_10969);
xor U15205 (N_15205,N_10068,N_10878);
nand U15206 (N_15206,N_9517,N_10015);
or U15207 (N_15207,N_8684,N_10744);
or U15208 (N_15208,N_11546,N_9987);
or U15209 (N_15209,N_9659,N_8879);
or U15210 (N_15210,N_10016,N_9936);
or U15211 (N_15211,N_8867,N_11082);
nor U15212 (N_15212,N_9836,N_9504);
xnor U15213 (N_15213,N_11070,N_11547);
and U15214 (N_15214,N_9755,N_9938);
nand U15215 (N_15215,N_9259,N_11788);
or U15216 (N_15216,N_8745,N_10152);
xnor U15217 (N_15217,N_9403,N_10315);
and U15218 (N_15218,N_8764,N_11336);
xnor U15219 (N_15219,N_10144,N_9115);
nor U15220 (N_15220,N_9853,N_10818);
or U15221 (N_15221,N_8545,N_10250);
nand U15222 (N_15222,N_9311,N_11915);
nand U15223 (N_15223,N_11555,N_8162);
xnor U15224 (N_15224,N_8243,N_10201);
and U15225 (N_15225,N_11302,N_9081);
and U15226 (N_15226,N_11590,N_8761);
nor U15227 (N_15227,N_9520,N_9957);
or U15228 (N_15228,N_10554,N_10277);
nand U15229 (N_15229,N_8623,N_11572);
nor U15230 (N_15230,N_11682,N_10123);
nor U15231 (N_15231,N_9584,N_8610);
nor U15232 (N_15232,N_10104,N_8763);
and U15233 (N_15233,N_9998,N_10468);
xor U15234 (N_15234,N_11729,N_11553);
nor U15235 (N_15235,N_10777,N_10097);
xnor U15236 (N_15236,N_11600,N_9671);
and U15237 (N_15237,N_9709,N_11282);
nand U15238 (N_15238,N_10361,N_8788);
or U15239 (N_15239,N_9256,N_8344);
and U15240 (N_15240,N_8919,N_11265);
nand U15241 (N_15241,N_9539,N_9272);
and U15242 (N_15242,N_9611,N_9655);
or U15243 (N_15243,N_9306,N_11323);
nor U15244 (N_15244,N_8494,N_11841);
and U15245 (N_15245,N_11288,N_9856);
nor U15246 (N_15246,N_9268,N_11059);
nand U15247 (N_15247,N_8274,N_8987);
nand U15248 (N_15248,N_8749,N_10999);
or U15249 (N_15249,N_11513,N_11917);
nand U15250 (N_15250,N_9219,N_10001);
nand U15251 (N_15251,N_11098,N_8862);
nor U15252 (N_15252,N_10741,N_8238);
nand U15253 (N_15253,N_8459,N_10823);
nand U15254 (N_15254,N_11633,N_9914);
and U15255 (N_15255,N_9189,N_9760);
xor U15256 (N_15256,N_11873,N_11153);
nor U15257 (N_15257,N_9021,N_10110);
nand U15258 (N_15258,N_11319,N_11019);
or U15259 (N_15259,N_8681,N_10600);
and U15260 (N_15260,N_8107,N_11898);
or U15261 (N_15261,N_11812,N_10055);
or U15262 (N_15262,N_9557,N_9421);
or U15263 (N_15263,N_9283,N_9718);
and U15264 (N_15264,N_10230,N_8102);
nand U15265 (N_15265,N_8706,N_8436);
nor U15266 (N_15266,N_11018,N_8587);
nor U15267 (N_15267,N_11719,N_8965);
nand U15268 (N_15268,N_10479,N_10074);
or U15269 (N_15269,N_8987,N_8476);
nor U15270 (N_15270,N_8440,N_9857);
and U15271 (N_15271,N_11317,N_11056);
nand U15272 (N_15272,N_10951,N_11173);
and U15273 (N_15273,N_9218,N_10674);
nor U15274 (N_15274,N_8321,N_10956);
and U15275 (N_15275,N_10812,N_10603);
and U15276 (N_15276,N_11047,N_10669);
nor U15277 (N_15277,N_10211,N_9107);
nand U15278 (N_15278,N_9319,N_9580);
nor U15279 (N_15279,N_11825,N_10645);
or U15280 (N_15280,N_10811,N_9494);
and U15281 (N_15281,N_10408,N_8031);
xnor U15282 (N_15282,N_8181,N_10209);
nor U15283 (N_15283,N_10572,N_11952);
xor U15284 (N_15284,N_9685,N_9032);
xnor U15285 (N_15285,N_11614,N_10454);
nand U15286 (N_15286,N_10145,N_10204);
nor U15287 (N_15287,N_10862,N_11001);
nand U15288 (N_15288,N_11757,N_8562);
xnor U15289 (N_15289,N_8174,N_11986);
nor U15290 (N_15290,N_11016,N_11844);
nor U15291 (N_15291,N_8499,N_11403);
nand U15292 (N_15292,N_8388,N_10746);
nor U15293 (N_15293,N_8331,N_10504);
or U15294 (N_15294,N_9717,N_11011);
nand U15295 (N_15295,N_9102,N_11505);
and U15296 (N_15296,N_8674,N_10305);
xnor U15297 (N_15297,N_11936,N_9126);
and U15298 (N_15298,N_9123,N_10221);
or U15299 (N_15299,N_11005,N_8696);
xor U15300 (N_15300,N_11288,N_9246);
nand U15301 (N_15301,N_8633,N_8564);
nor U15302 (N_15302,N_11375,N_10908);
nor U15303 (N_15303,N_11363,N_10373);
nor U15304 (N_15304,N_10961,N_10810);
and U15305 (N_15305,N_8268,N_8513);
nor U15306 (N_15306,N_8571,N_8512);
nor U15307 (N_15307,N_11676,N_10360);
nor U15308 (N_15308,N_8040,N_11008);
and U15309 (N_15309,N_10165,N_11616);
xor U15310 (N_15310,N_8981,N_8184);
or U15311 (N_15311,N_8703,N_8114);
and U15312 (N_15312,N_11988,N_8305);
nand U15313 (N_15313,N_8468,N_8679);
nand U15314 (N_15314,N_11399,N_10256);
nand U15315 (N_15315,N_9779,N_10630);
xor U15316 (N_15316,N_9833,N_10476);
or U15317 (N_15317,N_9388,N_8610);
xnor U15318 (N_15318,N_10799,N_9578);
and U15319 (N_15319,N_11180,N_10273);
xnor U15320 (N_15320,N_8158,N_8852);
xnor U15321 (N_15321,N_8196,N_11107);
xor U15322 (N_15322,N_10883,N_8855);
nand U15323 (N_15323,N_9921,N_8558);
xor U15324 (N_15324,N_9553,N_11748);
nand U15325 (N_15325,N_11039,N_8732);
nand U15326 (N_15326,N_11198,N_9578);
xor U15327 (N_15327,N_10719,N_10253);
and U15328 (N_15328,N_9979,N_9617);
nor U15329 (N_15329,N_8071,N_9651);
xnor U15330 (N_15330,N_10948,N_9668);
or U15331 (N_15331,N_8978,N_11333);
xor U15332 (N_15332,N_11025,N_11935);
nand U15333 (N_15333,N_10037,N_10493);
nand U15334 (N_15334,N_11756,N_10376);
xnor U15335 (N_15335,N_9356,N_11654);
or U15336 (N_15336,N_8235,N_9961);
nor U15337 (N_15337,N_9525,N_10399);
nor U15338 (N_15338,N_9222,N_8203);
nand U15339 (N_15339,N_9257,N_9099);
or U15340 (N_15340,N_10690,N_11652);
xor U15341 (N_15341,N_8061,N_9020);
nor U15342 (N_15342,N_10836,N_8395);
nor U15343 (N_15343,N_10181,N_9408);
nor U15344 (N_15344,N_10408,N_8139);
or U15345 (N_15345,N_11613,N_10117);
xnor U15346 (N_15346,N_8017,N_11212);
nand U15347 (N_15347,N_9891,N_10991);
xor U15348 (N_15348,N_8534,N_8177);
xor U15349 (N_15349,N_11611,N_10716);
and U15350 (N_15350,N_11266,N_11853);
nand U15351 (N_15351,N_8865,N_8029);
or U15352 (N_15352,N_10863,N_9117);
or U15353 (N_15353,N_10395,N_8984);
nor U15354 (N_15354,N_9292,N_10487);
and U15355 (N_15355,N_8362,N_10567);
nor U15356 (N_15356,N_8895,N_8197);
nor U15357 (N_15357,N_9836,N_11718);
xor U15358 (N_15358,N_11279,N_9043);
xnor U15359 (N_15359,N_9866,N_8447);
or U15360 (N_15360,N_9845,N_11555);
nand U15361 (N_15361,N_10701,N_10143);
nand U15362 (N_15362,N_9564,N_10584);
nand U15363 (N_15363,N_9007,N_8267);
xnor U15364 (N_15364,N_9785,N_11558);
and U15365 (N_15365,N_11063,N_9739);
xor U15366 (N_15366,N_11891,N_11522);
nand U15367 (N_15367,N_11793,N_8098);
or U15368 (N_15368,N_10714,N_10988);
nand U15369 (N_15369,N_10087,N_8089);
nand U15370 (N_15370,N_8954,N_9159);
nand U15371 (N_15371,N_10307,N_11483);
nor U15372 (N_15372,N_8062,N_10709);
nor U15373 (N_15373,N_9412,N_8190);
nor U15374 (N_15374,N_9599,N_10851);
nor U15375 (N_15375,N_9314,N_10649);
nor U15376 (N_15376,N_11179,N_11174);
and U15377 (N_15377,N_11793,N_10486);
xor U15378 (N_15378,N_10448,N_11138);
xor U15379 (N_15379,N_9320,N_10700);
nand U15380 (N_15380,N_9360,N_10541);
or U15381 (N_15381,N_9493,N_10761);
nand U15382 (N_15382,N_8887,N_9856);
or U15383 (N_15383,N_9269,N_11080);
nor U15384 (N_15384,N_9650,N_10510);
and U15385 (N_15385,N_8770,N_11112);
or U15386 (N_15386,N_11503,N_9004);
and U15387 (N_15387,N_11908,N_9616);
and U15388 (N_15388,N_8972,N_9562);
nand U15389 (N_15389,N_9557,N_8469);
or U15390 (N_15390,N_8796,N_11504);
nand U15391 (N_15391,N_11122,N_11624);
nor U15392 (N_15392,N_8554,N_11404);
xor U15393 (N_15393,N_9833,N_11910);
and U15394 (N_15394,N_11018,N_9316);
and U15395 (N_15395,N_9212,N_9236);
nand U15396 (N_15396,N_9048,N_9863);
xor U15397 (N_15397,N_11903,N_10774);
xor U15398 (N_15398,N_8303,N_10227);
nand U15399 (N_15399,N_9351,N_10953);
xor U15400 (N_15400,N_8051,N_10577);
nor U15401 (N_15401,N_11718,N_8735);
nor U15402 (N_15402,N_10942,N_11992);
xor U15403 (N_15403,N_10907,N_8074);
and U15404 (N_15404,N_8042,N_9501);
xor U15405 (N_15405,N_8049,N_10653);
xor U15406 (N_15406,N_9504,N_8978);
nor U15407 (N_15407,N_11707,N_10541);
xor U15408 (N_15408,N_10575,N_10059);
nand U15409 (N_15409,N_10252,N_10952);
and U15410 (N_15410,N_11832,N_11765);
nand U15411 (N_15411,N_11171,N_9146);
xnor U15412 (N_15412,N_9906,N_9297);
xor U15413 (N_15413,N_11611,N_8350);
xor U15414 (N_15414,N_9145,N_9511);
and U15415 (N_15415,N_9769,N_11896);
and U15416 (N_15416,N_8741,N_8970);
xor U15417 (N_15417,N_10030,N_11295);
and U15418 (N_15418,N_10172,N_11841);
nand U15419 (N_15419,N_9209,N_11102);
xnor U15420 (N_15420,N_10942,N_10586);
xnor U15421 (N_15421,N_8864,N_10676);
and U15422 (N_15422,N_9257,N_11693);
nand U15423 (N_15423,N_8453,N_10409);
nand U15424 (N_15424,N_8829,N_10587);
xor U15425 (N_15425,N_9582,N_8196);
xnor U15426 (N_15426,N_10669,N_10612);
xnor U15427 (N_15427,N_9762,N_10101);
and U15428 (N_15428,N_11756,N_8665);
and U15429 (N_15429,N_11558,N_11642);
nor U15430 (N_15430,N_10185,N_10413);
xor U15431 (N_15431,N_8547,N_9431);
or U15432 (N_15432,N_8852,N_10671);
nand U15433 (N_15433,N_8814,N_11690);
and U15434 (N_15434,N_10350,N_9564);
and U15435 (N_15435,N_10788,N_8692);
or U15436 (N_15436,N_11183,N_8520);
nor U15437 (N_15437,N_10229,N_8414);
and U15438 (N_15438,N_9406,N_10942);
xnor U15439 (N_15439,N_9390,N_9773);
nand U15440 (N_15440,N_10575,N_9417);
and U15441 (N_15441,N_10654,N_11615);
and U15442 (N_15442,N_10834,N_10893);
xor U15443 (N_15443,N_10735,N_8927);
nand U15444 (N_15444,N_8482,N_9587);
and U15445 (N_15445,N_8889,N_10336);
nor U15446 (N_15446,N_11112,N_10224);
and U15447 (N_15447,N_11505,N_10236);
and U15448 (N_15448,N_10239,N_9557);
xnor U15449 (N_15449,N_9072,N_11086);
and U15450 (N_15450,N_9087,N_9947);
and U15451 (N_15451,N_10162,N_10785);
xnor U15452 (N_15452,N_8379,N_9171);
nand U15453 (N_15453,N_11162,N_10141);
or U15454 (N_15454,N_10152,N_11598);
xor U15455 (N_15455,N_10326,N_9366);
nor U15456 (N_15456,N_11628,N_9305);
nand U15457 (N_15457,N_8619,N_10847);
nand U15458 (N_15458,N_10841,N_9265);
xor U15459 (N_15459,N_11075,N_8424);
and U15460 (N_15460,N_8423,N_9919);
and U15461 (N_15461,N_11606,N_10447);
xor U15462 (N_15462,N_8643,N_9536);
nor U15463 (N_15463,N_9365,N_8194);
nand U15464 (N_15464,N_11116,N_11678);
or U15465 (N_15465,N_11842,N_8659);
xor U15466 (N_15466,N_11885,N_11114);
nor U15467 (N_15467,N_9109,N_10021);
nand U15468 (N_15468,N_11777,N_8847);
and U15469 (N_15469,N_11922,N_8994);
nor U15470 (N_15470,N_10592,N_10613);
or U15471 (N_15471,N_10979,N_9918);
nand U15472 (N_15472,N_9172,N_11165);
nor U15473 (N_15473,N_9493,N_9859);
xnor U15474 (N_15474,N_9303,N_10599);
nor U15475 (N_15475,N_10880,N_9634);
nor U15476 (N_15476,N_9812,N_8722);
nand U15477 (N_15477,N_8889,N_8323);
xor U15478 (N_15478,N_10112,N_10824);
nand U15479 (N_15479,N_8102,N_11383);
nand U15480 (N_15480,N_11888,N_11056);
nand U15481 (N_15481,N_8962,N_11009);
nand U15482 (N_15482,N_8137,N_11126);
nor U15483 (N_15483,N_8789,N_11221);
and U15484 (N_15484,N_9974,N_9079);
nor U15485 (N_15485,N_9240,N_11165);
nor U15486 (N_15486,N_11196,N_9319);
nand U15487 (N_15487,N_9865,N_8120);
or U15488 (N_15488,N_9012,N_8382);
nor U15489 (N_15489,N_8980,N_9025);
nor U15490 (N_15490,N_10070,N_11681);
or U15491 (N_15491,N_10114,N_9760);
nand U15492 (N_15492,N_9596,N_9063);
xor U15493 (N_15493,N_10192,N_11619);
nor U15494 (N_15494,N_9587,N_8339);
and U15495 (N_15495,N_11229,N_9757);
and U15496 (N_15496,N_11049,N_9706);
or U15497 (N_15497,N_9892,N_8972);
or U15498 (N_15498,N_10896,N_11644);
or U15499 (N_15499,N_9765,N_11728);
xnor U15500 (N_15500,N_10603,N_11198);
nand U15501 (N_15501,N_10884,N_8519);
xnor U15502 (N_15502,N_10100,N_8640);
and U15503 (N_15503,N_11325,N_10816);
nor U15504 (N_15504,N_11984,N_9636);
and U15505 (N_15505,N_8637,N_8071);
nand U15506 (N_15506,N_9976,N_9458);
or U15507 (N_15507,N_8269,N_10842);
nor U15508 (N_15508,N_8132,N_10306);
xnor U15509 (N_15509,N_9221,N_10062);
nand U15510 (N_15510,N_9606,N_9056);
or U15511 (N_15511,N_8132,N_11297);
nand U15512 (N_15512,N_8720,N_8889);
nand U15513 (N_15513,N_9479,N_8129);
nand U15514 (N_15514,N_8682,N_9993);
nor U15515 (N_15515,N_8666,N_10375);
or U15516 (N_15516,N_11280,N_11203);
xnor U15517 (N_15517,N_8025,N_9004);
nor U15518 (N_15518,N_11796,N_11672);
nand U15519 (N_15519,N_11154,N_10773);
nor U15520 (N_15520,N_8026,N_11536);
nand U15521 (N_15521,N_11599,N_10101);
or U15522 (N_15522,N_11502,N_9954);
and U15523 (N_15523,N_9845,N_11891);
nand U15524 (N_15524,N_11201,N_9053);
nor U15525 (N_15525,N_8403,N_8310);
nand U15526 (N_15526,N_9347,N_11172);
xor U15527 (N_15527,N_11270,N_9272);
nor U15528 (N_15528,N_10032,N_10657);
or U15529 (N_15529,N_11394,N_9751);
xnor U15530 (N_15530,N_11862,N_9713);
xor U15531 (N_15531,N_10578,N_11741);
nand U15532 (N_15532,N_11279,N_8845);
xor U15533 (N_15533,N_11140,N_10531);
nand U15534 (N_15534,N_8268,N_10973);
or U15535 (N_15535,N_10536,N_8996);
or U15536 (N_15536,N_11525,N_10976);
nand U15537 (N_15537,N_8540,N_11515);
nand U15538 (N_15538,N_8785,N_11746);
or U15539 (N_15539,N_8605,N_11955);
nor U15540 (N_15540,N_9548,N_8556);
nor U15541 (N_15541,N_9768,N_8947);
xor U15542 (N_15542,N_9196,N_9572);
nand U15543 (N_15543,N_10665,N_11802);
and U15544 (N_15544,N_11416,N_10542);
nand U15545 (N_15545,N_9045,N_10908);
or U15546 (N_15546,N_9515,N_10691);
and U15547 (N_15547,N_10671,N_11905);
xnor U15548 (N_15548,N_10069,N_9043);
or U15549 (N_15549,N_10280,N_8415);
or U15550 (N_15550,N_9436,N_8826);
nor U15551 (N_15551,N_8090,N_10605);
xor U15552 (N_15552,N_8007,N_8344);
nand U15553 (N_15553,N_8933,N_11411);
xor U15554 (N_15554,N_9400,N_11237);
nor U15555 (N_15555,N_8949,N_10828);
nand U15556 (N_15556,N_11597,N_9704);
xor U15557 (N_15557,N_9327,N_9858);
or U15558 (N_15558,N_8203,N_10114);
or U15559 (N_15559,N_8851,N_10667);
nand U15560 (N_15560,N_10520,N_11632);
and U15561 (N_15561,N_10828,N_11113);
nand U15562 (N_15562,N_10038,N_11989);
or U15563 (N_15563,N_8842,N_11019);
and U15564 (N_15564,N_11773,N_11035);
xor U15565 (N_15565,N_9746,N_8839);
or U15566 (N_15566,N_11193,N_9990);
and U15567 (N_15567,N_11507,N_9834);
and U15568 (N_15568,N_10263,N_8167);
or U15569 (N_15569,N_10831,N_11724);
nand U15570 (N_15570,N_8757,N_8629);
nor U15571 (N_15571,N_11440,N_8464);
nand U15572 (N_15572,N_9940,N_11216);
and U15573 (N_15573,N_8146,N_11815);
xnor U15574 (N_15574,N_10165,N_11217);
and U15575 (N_15575,N_8649,N_8826);
or U15576 (N_15576,N_11326,N_10475);
xor U15577 (N_15577,N_9004,N_10671);
nor U15578 (N_15578,N_8094,N_8583);
xnor U15579 (N_15579,N_8561,N_9324);
and U15580 (N_15580,N_10233,N_10696);
nand U15581 (N_15581,N_10328,N_9029);
xor U15582 (N_15582,N_9710,N_9957);
nand U15583 (N_15583,N_9090,N_9657);
or U15584 (N_15584,N_11866,N_10136);
xnor U15585 (N_15585,N_9810,N_11911);
nand U15586 (N_15586,N_8215,N_9294);
nand U15587 (N_15587,N_10418,N_11865);
or U15588 (N_15588,N_8939,N_11215);
xor U15589 (N_15589,N_10892,N_11191);
nand U15590 (N_15590,N_11895,N_9868);
nand U15591 (N_15591,N_10070,N_9074);
xor U15592 (N_15592,N_8650,N_9273);
nor U15593 (N_15593,N_10253,N_11943);
and U15594 (N_15594,N_10705,N_9071);
nand U15595 (N_15595,N_10022,N_11398);
and U15596 (N_15596,N_8138,N_9401);
and U15597 (N_15597,N_11542,N_11912);
nor U15598 (N_15598,N_9800,N_11871);
and U15599 (N_15599,N_9657,N_10166);
xor U15600 (N_15600,N_10660,N_9624);
nand U15601 (N_15601,N_8103,N_10106);
or U15602 (N_15602,N_10346,N_8539);
nand U15603 (N_15603,N_11408,N_10165);
and U15604 (N_15604,N_10455,N_8637);
xor U15605 (N_15605,N_10757,N_8207);
nor U15606 (N_15606,N_9059,N_10710);
nor U15607 (N_15607,N_11652,N_10665);
nor U15608 (N_15608,N_8373,N_11646);
nor U15609 (N_15609,N_8975,N_10353);
xnor U15610 (N_15610,N_10263,N_8452);
nand U15611 (N_15611,N_11820,N_9683);
xnor U15612 (N_15612,N_9286,N_11654);
and U15613 (N_15613,N_8614,N_8048);
and U15614 (N_15614,N_10014,N_11047);
or U15615 (N_15615,N_10689,N_10154);
xnor U15616 (N_15616,N_8058,N_8154);
nand U15617 (N_15617,N_10722,N_9619);
xor U15618 (N_15618,N_9451,N_8797);
xnor U15619 (N_15619,N_9841,N_8754);
nor U15620 (N_15620,N_10925,N_11718);
and U15621 (N_15621,N_9164,N_9606);
xnor U15622 (N_15622,N_11726,N_8402);
or U15623 (N_15623,N_11293,N_8608);
nand U15624 (N_15624,N_10892,N_8148);
and U15625 (N_15625,N_11394,N_9755);
xnor U15626 (N_15626,N_8892,N_10450);
or U15627 (N_15627,N_8758,N_10620);
nand U15628 (N_15628,N_11354,N_11672);
and U15629 (N_15629,N_10747,N_9160);
nor U15630 (N_15630,N_10300,N_9328);
and U15631 (N_15631,N_9430,N_11648);
or U15632 (N_15632,N_8921,N_10993);
xnor U15633 (N_15633,N_9508,N_11345);
nand U15634 (N_15634,N_10474,N_9696);
or U15635 (N_15635,N_8176,N_10566);
xor U15636 (N_15636,N_8303,N_11709);
nor U15637 (N_15637,N_11820,N_10149);
nor U15638 (N_15638,N_11895,N_10664);
or U15639 (N_15639,N_11984,N_9720);
nor U15640 (N_15640,N_11035,N_8802);
or U15641 (N_15641,N_11009,N_10128);
or U15642 (N_15642,N_8602,N_11393);
or U15643 (N_15643,N_10863,N_9482);
nor U15644 (N_15644,N_9078,N_10161);
xnor U15645 (N_15645,N_8017,N_10872);
xor U15646 (N_15646,N_9854,N_8102);
nor U15647 (N_15647,N_9492,N_8874);
and U15648 (N_15648,N_8593,N_10871);
nor U15649 (N_15649,N_11059,N_8697);
or U15650 (N_15650,N_8661,N_10699);
or U15651 (N_15651,N_9180,N_11100);
nor U15652 (N_15652,N_10851,N_11175);
and U15653 (N_15653,N_11189,N_10938);
nand U15654 (N_15654,N_8386,N_8859);
nand U15655 (N_15655,N_11302,N_10128);
xnor U15656 (N_15656,N_11323,N_10414);
or U15657 (N_15657,N_9464,N_9879);
nand U15658 (N_15658,N_8102,N_11390);
or U15659 (N_15659,N_11759,N_10977);
xnor U15660 (N_15660,N_11110,N_10643);
and U15661 (N_15661,N_8342,N_11714);
and U15662 (N_15662,N_11441,N_10497);
or U15663 (N_15663,N_10403,N_8932);
or U15664 (N_15664,N_8995,N_8938);
or U15665 (N_15665,N_9029,N_11727);
xnor U15666 (N_15666,N_8383,N_11782);
and U15667 (N_15667,N_9951,N_11357);
and U15668 (N_15668,N_11521,N_10374);
and U15669 (N_15669,N_8883,N_8208);
and U15670 (N_15670,N_8712,N_11070);
nand U15671 (N_15671,N_10668,N_11285);
and U15672 (N_15672,N_11214,N_9151);
xnor U15673 (N_15673,N_9113,N_10499);
or U15674 (N_15674,N_9466,N_9053);
nor U15675 (N_15675,N_11231,N_8650);
xnor U15676 (N_15676,N_10685,N_9979);
nand U15677 (N_15677,N_10027,N_8170);
or U15678 (N_15678,N_10096,N_8031);
nor U15679 (N_15679,N_8082,N_9431);
xnor U15680 (N_15680,N_8679,N_9996);
and U15681 (N_15681,N_8224,N_8697);
xor U15682 (N_15682,N_11853,N_8552);
xor U15683 (N_15683,N_11273,N_8518);
nand U15684 (N_15684,N_10239,N_11932);
nand U15685 (N_15685,N_9048,N_8875);
and U15686 (N_15686,N_8146,N_8308);
nand U15687 (N_15687,N_11924,N_8982);
or U15688 (N_15688,N_10381,N_10652);
and U15689 (N_15689,N_11521,N_10556);
xor U15690 (N_15690,N_9889,N_11082);
and U15691 (N_15691,N_11739,N_9369);
nor U15692 (N_15692,N_10522,N_8306);
nand U15693 (N_15693,N_11276,N_8068);
nor U15694 (N_15694,N_10436,N_9520);
or U15695 (N_15695,N_10144,N_8141);
nand U15696 (N_15696,N_10047,N_8615);
nand U15697 (N_15697,N_10353,N_8761);
nand U15698 (N_15698,N_10037,N_8483);
and U15699 (N_15699,N_10189,N_9508);
nand U15700 (N_15700,N_10157,N_8688);
and U15701 (N_15701,N_8973,N_9990);
xnor U15702 (N_15702,N_8487,N_10458);
and U15703 (N_15703,N_11405,N_8029);
and U15704 (N_15704,N_11069,N_10063);
nor U15705 (N_15705,N_9622,N_10513);
nor U15706 (N_15706,N_11308,N_8792);
and U15707 (N_15707,N_9778,N_9816);
nor U15708 (N_15708,N_11232,N_9077);
or U15709 (N_15709,N_10771,N_8434);
and U15710 (N_15710,N_11750,N_8085);
nand U15711 (N_15711,N_11289,N_8525);
nor U15712 (N_15712,N_11703,N_11888);
nand U15713 (N_15713,N_8055,N_11190);
nor U15714 (N_15714,N_8895,N_8686);
nor U15715 (N_15715,N_8324,N_11460);
nor U15716 (N_15716,N_10911,N_8598);
and U15717 (N_15717,N_11771,N_9576);
xor U15718 (N_15718,N_11690,N_8343);
nand U15719 (N_15719,N_10773,N_9855);
xnor U15720 (N_15720,N_9177,N_8397);
xor U15721 (N_15721,N_9850,N_9179);
nor U15722 (N_15722,N_8643,N_8108);
nand U15723 (N_15723,N_8921,N_11271);
nand U15724 (N_15724,N_11397,N_10422);
nor U15725 (N_15725,N_8236,N_9843);
nor U15726 (N_15726,N_11751,N_11066);
and U15727 (N_15727,N_9419,N_9270);
nand U15728 (N_15728,N_9564,N_9664);
and U15729 (N_15729,N_11699,N_10690);
and U15730 (N_15730,N_11677,N_10415);
xor U15731 (N_15731,N_9085,N_11446);
xor U15732 (N_15732,N_9910,N_11079);
or U15733 (N_15733,N_9595,N_8698);
nor U15734 (N_15734,N_11321,N_8709);
or U15735 (N_15735,N_9906,N_11126);
or U15736 (N_15736,N_11230,N_8645);
or U15737 (N_15737,N_9731,N_10778);
nor U15738 (N_15738,N_11930,N_9645);
and U15739 (N_15739,N_11973,N_10039);
and U15740 (N_15740,N_10587,N_9987);
nor U15741 (N_15741,N_9894,N_9083);
xnor U15742 (N_15742,N_10571,N_11402);
or U15743 (N_15743,N_8498,N_9421);
and U15744 (N_15744,N_9051,N_9531);
nand U15745 (N_15745,N_8378,N_9218);
nor U15746 (N_15746,N_8217,N_8108);
nand U15747 (N_15747,N_9931,N_8982);
and U15748 (N_15748,N_8949,N_8557);
nand U15749 (N_15749,N_10470,N_11789);
or U15750 (N_15750,N_10115,N_10029);
xor U15751 (N_15751,N_8514,N_8037);
nor U15752 (N_15752,N_11621,N_11060);
nand U15753 (N_15753,N_10273,N_8443);
nand U15754 (N_15754,N_10752,N_8165);
and U15755 (N_15755,N_10494,N_10465);
xor U15756 (N_15756,N_9787,N_9121);
or U15757 (N_15757,N_11655,N_8184);
xnor U15758 (N_15758,N_9157,N_10573);
or U15759 (N_15759,N_11339,N_10277);
or U15760 (N_15760,N_9809,N_8067);
xor U15761 (N_15761,N_11699,N_9286);
and U15762 (N_15762,N_8306,N_10193);
nor U15763 (N_15763,N_10745,N_10501);
xor U15764 (N_15764,N_10410,N_11395);
nor U15765 (N_15765,N_11316,N_9084);
nor U15766 (N_15766,N_9330,N_8364);
xor U15767 (N_15767,N_9604,N_9900);
nand U15768 (N_15768,N_8231,N_9379);
nor U15769 (N_15769,N_8784,N_11976);
or U15770 (N_15770,N_8223,N_9346);
xnor U15771 (N_15771,N_11633,N_8939);
xnor U15772 (N_15772,N_11885,N_10073);
nand U15773 (N_15773,N_8427,N_9196);
xnor U15774 (N_15774,N_8218,N_8567);
nand U15775 (N_15775,N_10708,N_10714);
nor U15776 (N_15776,N_9282,N_11459);
xnor U15777 (N_15777,N_8884,N_9550);
nand U15778 (N_15778,N_10111,N_10284);
nand U15779 (N_15779,N_9928,N_9762);
nor U15780 (N_15780,N_11586,N_10574);
and U15781 (N_15781,N_11764,N_8449);
nor U15782 (N_15782,N_8123,N_11838);
nor U15783 (N_15783,N_8631,N_8865);
nand U15784 (N_15784,N_10295,N_9440);
xnor U15785 (N_15785,N_10183,N_11341);
nor U15786 (N_15786,N_8375,N_11383);
or U15787 (N_15787,N_9144,N_11918);
xor U15788 (N_15788,N_8996,N_9101);
and U15789 (N_15789,N_8704,N_8223);
xor U15790 (N_15790,N_8826,N_10015);
nor U15791 (N_15791,N_8594,N_9703);
and U15792 (N_15792,N_8460,N_11443);
or U15793 (N_15793,N_8326,N_9285);
nand U15794 (N_15794,N_9416,N_11177);
nand U15795 (N_15795,N_9964,N_8961);
nand U15796 (N_15796,N_11788,N_11074);
xnor U15797 (N_15797,N_9208,N_9191);
or U15798 (N_15798,N_11758,N_11012);
xor U15799 (N_15799,N_9485,N_10040);
xnor U15800 (N_15800,N_8792,N_10777);
nand U15801 (N_15801,N_9775,N_10990);
or U15802 (N_15802,N_9117,N_11323);
nand U15803 (N_15803,N_8541,N_10467);
and U15804 (N_15804,N_8109,N_8902);
xor U15805 (N_15805,N_8530,N_8110);
and U15806 (N_15806,N_9660,N_10128);
nand U15807 (N_15807,N_9117,N_11595);
or U15808 (N_15808,N_11150,N_8488);
nand U15809 (N_15809,N_10650,N_9048);
xnor U15810 (N_15810,N_9906,N_9432);
nor U15811 (N_15811,N_9635,N_11221);
xnor U15812 (N_15812,N_8496,N_8557);
or U15813 (N_15813,N_11605,N_11390);
nor U15814 (N_15814,N_8841,N_11357);
or U15815 (N_15815,N_8088,N_11918);
and U15816 (N_15816,N_10147,N_10735);
or U15817 (N_15817,N_9105,N_8645);
and U15818 (N_15818,N_11790,N_8933);
nand U15819 (N_15819,N_9537,N_10675);
and U15820 (N_15820,N_9868,N_9478);
xnor U15821 (N_15821,N_9517,N_11544);
and U15822 (N_15822,N_9881,N_11063);
and U15823 (N_15823,N_9966,N_8692);
nor U15824 (N_15824,N_8933,N_9397);
or U15825 (N_15825,N_9179,N_10788);
and U15826 (N_15826,N_9623,N_10240);
nor U15827 (N_15827,N_8098,N_9966);
nand U15828 (N_15828,N_10910,N_8967);
or U15829 (N_15829,N_9229,N_8563);
or U15830 (N_15830,N_11170,N_8676);
and U15831 (N_15831,N_8645,N_8037);
nor U15832 (N_15832,N_8494,N_8001);
or U15833 (N_15833,N_9632,N_10637);
or U15834 (N_15834,N_9531,N_11159);
xnor U15835 (N_15835,N_9946,N_9526);
xor U15836 (N_15836,N_11107,N_11888);
and U15837 (N_15837,N_11796,N_11987);
xnor U15838 (N_15838,N_8886,N_8906);
nor U15839 (N_15839,N_10031,N_11562);
xnor U15840 (N_15840,N_10491,N_11714);
xnor U15841 (N_15841,N_8988,N_11921);
nand U15842 (N_15842,N_10508,N_10742);
xor U15843 (N_15843,N_9102,N_9051);
nand U15844 (N_15844,N_10709,N_8626);
and U15845 (N_15845,N_9438,N_9215);
or U15846 (N_15846,N_11894,N_11098);
or U15847 (N_15847,N_8757,N_10458);
xnor U15848 (N_15848,N_11604,N_9466);
nand U15849 (N_15849,N_9593,N_8164);
nor U15850 (N_15850,N_9328,N_11412);
or U15851 (N_15851,N_11710,N_11764);
nor U15852 (N_15852,N_9178,N_10407);
nor U15853 (N_15853,N_11827,N_8736);
nor U15854 (N_15854,N_11477,N_8942);
nor U15855 (N_15855,N_10870,N_11406);
or U15856 (N_15856,N_11332,N_10835);
and U15857 (N_15857,N_11172,N_11896);
or U15858 (N_15858,N_10228,N_10264);
nand U15859 (N_15859,N_10633,N_11677);
nand U15860 (N_15860,N_11228,N_10336);
and U15861 (N_15861,N_11231,N_11219);
xnor U15862 (N_15862,N_10484,N_10997);
or U15863 (N_15863,N_10806,N_11553);
xnor U15864 (N_15864,N_10463,N_9277);
and U15865 (N_15865,N_9804,N_8912);
xor U15866 (N_15866,N_8243,N_11039);
xnor U15867 (N_15867,N_9727,N_10774);
and U15868 (N_15868,N_9286,N_9217);
nor U15869 (N_15869,N_9723,N_9785);
nor U15870 (N_15870,N_11435,N_10611);
nor U15871 (N_15871,N_11015,N_8436);
and U15872 (N_15872,N_8799,N_9014);
and U15873 (N_15873,N_9064,N_11982);
xnor U15874 (N_15874,N_10985,N_11791);
nor U15875 (N_15875,N_10416,N_11733);
and U15876 (N_15876,N_10499,N_10264);
and U15877 (N_15877,N_8348,N_11654);
xnor U15878 (N_15878,N_11071,N_10111);
xor U15879 (N_15879,N_8304,N_11041);
or U15880 (N_15880,N_10470,N_9564);
xnor U15881 (N_15881,N_10800,N_9772);
nor U15882 (N_15882,N_9113,N_8053);
and U15883 (N_15883,N_9911,N_11574);
or U15884 (N_15884,N_9954,N_10646);
nor U15885 (N_15885,N_10688,N_10250);
or U15886 (N_15886,N_11365,N_10577);
and U15887 (N_15887,N_10695,N_8844);
and U15888 (N_15888,N_8279,N_9722);
nor U15889 (N_15889,N_11575,N_8388);
nor U15890 (N_15890,N_10471,N_8357);
nor U15891 (N_15891,N_11727,N_11500);
or U15892 (N_15892,N_10966,N_8746);
or U15893 (N_15893,N_9138,N_11269);
xnor U15894 (N_15894,N_10392,N_11007);
nor U15895 (N_15895,N_8689,N_9402);
or U15896 (N_15896,N_9880,N_11008);
xor U15897 (N_15897,N_9635,N_8415);
nor U15898 (N_15898,N_10156,N_8566);
nand U15899 (N_15899,N_8961,N_11505);
nand U15900 (N_15900,N_8980,N_9277);
nor U15901 (N_15901,N_11709,N_9458);
nand U15902 (N_15902,N_9189,N_10353);
or U15903 (N_15903,N_8441,N_8292);
or U15904 (N_15904,N_11648,N_8482);
or U15905 (N_15905,N_8101,N_8639);
and U15906 (N_15906,N_8777,N_8721);
xnor U15907 (N_15907,N_9826,N_10530);
or U15908 (N_15908,N_9397,N_8878);
nor U15909 (N_15909,N_11299,N_9012);
nand U15910 (N_15910,N_9144,N_8792);
xnor U15911 (N_15911,N_8099,N_8182);
or U15912 (N_15912,N_11996,N_9833);
and U15913 (N_15913,N_8455,N_11511);
and U15914 (N_15914,N_10531,N_10237);
nand U15915 (N_15915,N_10625,N_8652);
nand U15916 (N_15916,N_10503,N_11692);
or U15917 (N_15917,N_10340,N_8593);
xor U15918 (N_15918,N_11163,N_11977);
or U15919 (N_15919,N_11666,N_10323);
and U15920 (N_15920,N_11674,N_11734);
nand U15921 (N_15921,N_10309,N_8378);
and U15922 (N_15922,N_8983,N_9436);
or U15923 (N_15923,N_8808,N_8714);
nor U15924 (N_15924,N_10068,N_8963);
and U15925 (N_15925,N_11155,N_8413);
and U15926 (N_15926,N_10645,N_10272);
nor U15927 (N_15927,N_11333,N_8331);
nand U15928 (N_15928,N_9272,N_9587);
nand U15929 (N_15929,N_10731,N_11422);
and U15930 (N_15930,N_10934,N_9216);
or U15931 (N_15931,N_9537,N_11267);
nand U15932 (N_15932,N_9149,N_10700);
or U15933 (N_15933,N_11244,N_9368);
xnor U15934 (N_15934,N_10663,N_11275);
nand U15935 (N_15935,N_11356,N_9472);
xnor U15936 (N_15936,N_8889,N_11182);
nand U15937 (N_15937,N_10500,N_10344);
or U15938 (N_15938,N_11560,N_8908);
nor U15939 (N_15939,N_9062,N_8901);
xor U15940 (N_15940,N_9697,N_10262);
nor U15941 (N_15941,N_10138,N_8202);
and U15942 (N_15942,N_11653,N_10216);
xor U15943 (N_15943,N_8270,N_8359);
or U15944 (N_15944,N_8822,N_11153);
and U15945 (N_15945,N_11322,N_11089);
nor U15946 (N_15946,N_11742,N_11516);
xor U15947 (N_15947,N_9815,N_8343);
or U15948 (N_15948,N_11216,N_8415);
and U15949 (N_15949,N_9656,N_10010);
xor U15950 (N_15950,N_11744,N_11241);
or U15951 (N_15951,N_9397,N_9560);
and U15952 (N_15952,N_9201,N_9023);
nor U15953 (N_15953,N_9096,N_9525);
xor U15954 (N_15954,N_9718,N_8685);
nand U15955 (N_15955,N_11541,N_10203);
nand U15956 (N_15956,N_8662,N_11844);
nand U15957 (N_15957,N_11673,N_11589);
or U15958 (N_15958,N_11657,N_8194);
or U15959 (N_15959,N_8864,N_8972);
and U15960 (N_15960,N_10171,N_11711);
and U15961 (N_15961,N_10910,N_9994);
xor U15962 (N_15962,N_10900,N_10387);
xor U15963 (N_15963,N_9310,N_10193);
xnor U15964 (N_15964,N_10327,N_11662);
xor U15965 (N_15965,N_10919,N_8692);
nor U15966 (N_15966,N_11062,N_11233);
nand U15967 (N_15967,N_11085,N_10480);
nor U15968 (N_15968,N_8140,N_11301);
xor U15969 (N_15969,N_11563,N_11727);
nor U15970 (N_15970,N_10461,N_11495);
or U15971 (N_15971,N_10960,N_11916);
and U15972 (N_15972,N_9408,N_10638);
or U15973 (N_15973,N_11677,N_10028);
xnor U15974 (N_15974,N_9896,N_10153);
or U15975 (N_15975,N_9465,N_10488);
xor U15976 (N_15976,N_11664,N_8647);
or U15977 (N_15977,N_8485,N_8869);
xnor U15978 (N_15978,N_11959,N_10614);
or U15979 (N_15979,N_11650,N_8720);
nor U15980 (N_15980,N_9796,N_8683);
nor U15981 (N_15981,N_9690,N_9141);
nand U15982 (N_15982,N_9899,N_9165);
nand U15983 (N_15983,N_8353,N_11149);
xor U15984 (N_15984,N_10342,N_10743);
nand U15985 (N_15985,N_10171,N_11025);
nor U15986 (N_15986,N_11932,N_9103);
or U15987 (N_15987,N_8116,N_10506);
nor U15988 (N_15988,N_11878,N_11929);
nor U15989 (N_15989,N_8666,N_11561);
nor U15990 (N_15990,N_11932,N_10867);
xnor U15991 (N_15991,N_9461,N_10391);
nor U15992 (N_15992,N_10315,N_9634);
xor U15993 (N_15993,N_11285,N_10129);
xor U15994 (N_15994,N_9781,N_8054);
xor U15995 (N_15995,N_9663,N_11901);
and U15996 (N_15996,N_11874,N_8151);
and U15997 (N_15997,N_11738,N_10806);
nor U15998 (N_15998,N_11024,N_8481);
nor U15999 (N_15999,N_10750,N_11811);
and U16000 (N_16000,N_12534,N_14961);
nand U16001 (N_16001,N_14028,N_12543);
and U16002 (N_16002,N_13930,N_14639);
nor U16003 (N_16003,N_15039,N_15404);
or U16004 (N_16004,N_13898,N_12131);
or U16005 (N_16005,N_13596,N_13748);
and U16006 (N_16006,N_13801,N_15619);
xor U16007 (N_16007,N_15721,N_15104);
and U16008 (N_16008,N_13462,N_13319);
nand U16009 (N_16009,N_14108,N_13450);
or U16010 (N_16010,N_13443,N_14192);
and U16011 (N_16011,N_15422,N_15548);
xnor U16012 (N_16012,N_14363,N_14796);
nor U16013 (N_16013,N_14749,N_13533);
and U16014 (N_16014,N_15597,N_12774);
or U16015 (N_16015,N_12233,N_12448);
or U16016 (N_16016,N_15003,N_12752);
nand U16017 (N_16017,N_12686,N_14465);
or U16018 (N_16018,N_15752,N_15972);
nand U16019 (N_16019,N_14853,N_12865);
nor U16020 (N_16020,N_12362,N_14246);
nand U16021 (N_16021,N_12620,N_15711);
nor U16022 (N_16022,N_12129,N_13142);
xor U16023 (N_16023,N_14279,N_15198);
nor U16024 (N_16024,N_12381,N_12922);
nand U16025 (N_16025,N_14384,N_15906);
and U16026 (N_16026,N_15055,N_15199);
or U16027 (N_16027,N_14197,N_13239);
nand U16028 (N_16028,N_15970,N_15608);
or U16029 (N_16029,N_15434,N_15320);
nand U16030 (N_16030,N_15505,N_14349);
nand U16031 (N_16031,N_15487,N_13904);
nand U16032 (N_16032,N_14615,N_14631);
xor U16033 (N_16033,N_15694,N_12301);
or U16034 (N_16034,N_13640,N_14797);
xnor U16035 (N_16035,N_14560,N_13112);
nand U16036 (N_16036,N_12683,N_13000);
and U16037 (N_16037,N_13136,N_12216);
or U16038 (N_16038,N_14259,N_13742);
xnor U16039 (N_16039,N_15601,N_15478);
and U16040 (N_16040,N_14202,N_13297);
or U16041 (N_16041,N_14308,N_15835);
xnor U16042 (N_16042,N_14479,N_12291);
xor U16043 (N_16043,N_14158,N_13526);
nor U16044 (N_16044,N_12294,N_12570);
or U16045 (N_16045,N_14078,N_15354);
xor U16046 (N_16046,N_14050,N_15468);
or U16047 (N_16047,N_15379,N_13939);
nand U16048 (N_16048,N_12529,N_13288);
and U16049 (N_16049,N_14643,N_12626);
or U16050 (N_16050,N_12147,N_12780);
nand U16051 (N_16051,N_15025,N_12115);
nand U16052 (N_16052,N_12361,N_12152);
nand U16053 (N_16053,N_14449,N_14871);
and U16054 (N_16054,N_13090,N_14657);
or U16055 (N_16055,N_12082,N_14293);
nor U16056 (N_16056,N_15890,N_14032);
and U16057 (N_16057,N_12897,N_15408);
nor U16058 (N_16058,N_14404,N_15451);
and U16059 (N_16059,N_14154,N_12642);
or U16060 (N_16060,N_12271,N_14885);
nor U16061 (N_16061,N_12662,N_13960);
nand U16062 (N_16062,N_12071,N_14589);
xor U16063 (N_16063,N_12490,N_13964);
or U16064 (N_16064,N_15265,N_12128);
and U16065 (N_16065,N_15357,N_15576);
xor U16066 (N_16066,N_12306,N_13353);
or U16067 (N_16067,N_12622,N_13461);
nor U16068 (N_16068,N_12015,N_14025);
xor U16069 (N_16069,N_15334,N_13582);
or U16070 (N_16070,N_13900,N_14237);
nor U16071 (N_16071,N_12067,N_13950);
or U16072 (N_16072,N_15131,N_15176);
nand U16073 (N_16073,N_12196,N_15174);
nor U16074 (N_16074,N_12026,N_12459);
nand U16075 (N_16075,N_14642,N_13943);
xor U16076 (N_16076,N_13238,N_14566);
or U16077 (N_16077,N_13361,N_12045);
or U16078 (N_16078,N_15564,N_15460);
xnor U16079 (N_16079,N_14710,N_13671);
nand U16080 (N_16080,N_12770,N_13209);
or U16081 (N_16081,N_14618,N_15258);
nor U16082 (N_16082,N_14133,N_13468);
or U16083 (N_16083,N_15062,N_15290);
nor U16084 (N_16084,N_14283,N_12278);
nand U16085 (N_16085,N_14802,N_15660);
xor U16086 (N_16086,N_12215,N_12458);
nand U16087 (N_16087,N_14581,N_15403);
nor U16088 (N_16088,N_15923,N_14641);
nand U16089 (N_16089,N_15851,N_15538);
nand U16090 (N_16090,N_13798,N_14408);
or U16091 (N_16091,N_14607,N_13338);
xor U16092 (N_16092,N_12682,N_13255);
nand U16093 (N_16093,N_13169,N_13089);
nand U16094 (N_16094,N_13663,N_13860);
nand U16095 (N_16095,N_14896,N_12438);
nor U16096 (N_16096,N_15206,N_15935);
xnor U16097 (N_16097,N_14570,N_14811);
nor U16098 (N_16098,N_12224,N_15859);
and U16099 (N_16099,N_14357,N_14594);
xnor U16100 (N_16100,N_13464,N_13638);
xnor U16101 (N_16101,N_13863,N_12899);
or U16102 (N_16102,N_12533,N_15742);
nand U16103 (N_16103,N_12731,N_14650);
nand U16104 (N_16104,N_13689,N_14172);
nand U16105 (N_16105,N_14105,N_14272);
nand U16106 (N_16106,N_15778,N_13008);
or U16107 (N_16107,N_15223,N_12892);
and U16108 (N_16108,N_13481,N_14022);
xor U16109 (N_16109,N_15894,N_12228);
nor U16110 (N_16110,N_15042,N_14191);
xnor U16111 (N_16111,N_14280,N_14561);
xor U16112 (N_16112,N_12947,N_12343);
or U16113 (N_16113,N_15579,N_15847);
nand U16114 (N_16114,N_13507,N_12332);
xor U16115 (N_16115,N_14556,N_12065);
xnor U16116 (N_16116,N_12681,N_12424);
nor U16117 (N_16117,N_12334,N_13466);
xor U16118 (N_16118,N_13884,N_15433);
and U16119 (N_16119,N_13315,N_13454);
nand U16120 (N_16120,N_15865,N_12603);
or U16121 (N_16121,N_13349,N_13124);
or U16122 (N_16122,N_12217,N_13746);
xnor U16123 (N_16123,N_12698,N_14416);
nand U16124 (N_16124,N_12646,N_15498);
or U16125 (N_16125,N_15339,N_15627);
xnor U16126 (N_16126,N_15572,N_15236);
nor U16127 (N_16127,N_15382,N_15109);
nor U16128 (N_16128,N_12392,N_13809);
and U16129 (N_16129,N_13324,N_12193);
xnor U16130 (N_16130,N_14458,N_15232);
nand U16131 (N_16131,N_14957,N_13376);
nand U16132 (N_16132,N_13852,N_13535);
and U16133 (N_16133,N_15748,N_12333);
nor U16134 (N_16134,N_14413,N_12613);
nand U16135 (N_16135,N_14296,N_15183);
and U16136 (N_16136,N_15336,N_13757);
or U16137 (N_16137,N_14292,N_13325);
or U16138 (N_16138,N_13848,N_14997);
nand U16139 (N_16139,N_13267,N_15080);
and U16140 (N_16140,N_14793,N_13761);
xnor U16141 (N_16141,N_14966,N_14276);
or U16142 (N_16142,N_14524,N_15910);
nor U16143 (N_16143,N_14894,N_12755);
xnor U16144 (N_16144,N_12804,N_12862);
xnor U16145 (N_16145,N_13573,N_12275);
and U16146 (N_16146,N_13151,N_14623);
nand U16147 (N_16147,N_15998,N_14247);
or U16148 (N_16148,N_14313,N_12208);
nor U16149 (N_16149,N_14654,N_12888);
xor U16150 (N_16150,N_13052,N_15364);
nand U16151 (N_16151,N_14668,N_15209);
or U16152 (N_16152,N_13992,N_13684);
nor U16153 (N_16153,N_13694,N_12001);
nand U16154 (N_16154,N_15973,N_15361);
nand U16155 (N_16155,N_12076,N_12408);
xnor U16156 (N_16156,N_15896,N_15803);
and U16157 (N_16157,N_15056,N_14096);
and U16158 (N_16158,N_13605,N_12000);
nor U16159 (N_16159,N_15776,N_13143);
or U16160 (N_16160,N_15327,N_12996);
or U16161 (N_16161,N_14095,N_15014);
nor U16162 (N_16162,N_13666,N_12195);
nand U16163 (N_16163,N_14728,N_14175);
or U16164 (N_16164,N_14598,N_13038);
nor U16165 (N_16165,N_12644,N_12696);
or U16166 (N_16166,N_13816,N_15292);
nand U16167 (N_16167,N_15749,N_13808);
and U16168 (N_16168,N_14018,N_14778);
xor U16169 (N_16169,N_15402,N_15848);
xnor U16170 (N_16170,N_14083,N_14489);
or U16171 (N_16171,N_12016,N_13201);
xor U16172 (N_16172,N_13682,N_12905);
and U16173 (N_16173,N_15204,N_12759);
xnor U16174 (N_16174,N_13956,N_13426);
and U16175 (N_16175,N_13429,N_12474);
nand U16176 (N_16176,N_15815,N_12492);
xor U16177 (N_16177,N_13773,N_14635);
and U16178 (N_16178,N_15775,N_13381);
or U16179 (N_16179,N_12461,N_15846);
nand U16180 (N_16180,N_12403,N_12024);
nand U16181 (N_16181,N_15344,N_14249);
nor U16182 (N_16182,N_14010,N_12087);
and U16183 (N_16183,N_14300,N_12563);
nand U16184 (N_16184,N_13911,N_13487);
and U16185 (N_16185,N_13036,N_15479);
nand U16186 (N_16186,N_14502,N_12327);
and U16187 (N_16187,N_13252,N_13827);
xor U16188 (N_16188,N_14141,N_15149);
nand U16189 (N_16189,N_12859,N_13147);
and U16190 (N_16190,N_14161,N_14490);
xor U16191 (N_16191,N_14117,N_14858);
xor U16192 (N_16192,N_12803,N_14400);
nor U16193 (N_16193,N_13336,N_12842);
and U16194 (N_16194,N_12638,N_14454);
nor U16195 (N_16195,N_13404,N_12337);
xor U16196 (N_16196,N_13849,N_13519);
or U16197 (N_16197,N_12480,N_13735);
nand U16198 (N_16198,N_15872,N_12191);
nor U16199 (N_16199,N_12818,N_14774);
nand U16200 (N_16200,N_15684,N_14721);
nor U16201 (N_16201,N_12039,N_13921);
xor U16202 (N_16202,N_13790,N_15172);
xnor U16203 (N_16203,N_14850,N_14186);
nor U16204 (N_16204,N_15822,N_15448);
nand U16205 (N_16205,N_12468,N_12744);
nand U16206 (N_16206,N_12860,N_14697);
nor U16207 (N_16207,N_13562,N_12732);
nand U16208 (N_16208,N_12733,N_12265);
or U16209 (N_16209,N_15366,N_13722);
nand U16210 (N_16210,N_12421,N_14281);
xor U16211 (N_16211,N_12767,N_14829);
xnor U16212 (N_16212,N_13411,N_13138);
or U16213 (N_16213,N_15850,N_12876);
nor U16214 (N_16214,N_15637,N_14052);
and U16215 (N_16215,N_14744,N_13345);
and U16216 (N_16216,N_14763,N_12930);
and U16217 (N_16217,N_15255,N_12336);
nor U16218 (N_16218,N_12573,N_15351);
nand U16219 (N_16219,N_14859,N_15567);
nor U16220 (N_16220,N_12054,N_13941);
xor U16221 (N_16221,N_14346,N_12541);
or U16222 (N_16222,N_13776,N_14143);
xor U16223 (N_16223,N_14015,N_14146);
nand U16224 (N_16224,N_14954,N_13784);
or U16225 (N_16225,N_12237,N_13980);
xnor U16226 (N_16226,N_15770,N_13926);
nor U16227 (N_16227,N_13734,N_13044);
xnor U16228 (N_16228,N_15575,N_14717);
xor U16229 (N_16229,N_12377,N_12126);
xnor U16230 (N_16230,N_12820,N_12238);
nor U16231 (N_16231,N_15342,N_14203);
and U16232 (N_16232,N_13854,N_13300);
nand U16233 (N_16233,N_15086,N_15257);
nor U16234 (N_16234,N_13009,N_14890);
nor U16235 (N_16235,N_12349,N_15490);
or U16236 (N_16236,N_13914,N_15671);
and U16237 (N_16237,N_12560,N_12510);
xnor U16238 (N_16238,N_12960,N_15173);
xnor U16239 (N_16239,N_15501,N_15921);
xnor U16240 (N_16240,N_13749,N_12070);
nor U16241 (N_16241,N_13826,N_15115);
and U16242 (N_16242,N_14358,N_15667);
and U16243 (N_16243,N_12198,N_12887);
xor U16244 (N_16244,N_12599,N_14538);
and U16245 (N_16245,N_13831,N_13316);
and U16246 (N_16246,N_13499,N_15124);
nor U16247 (N_16247,N_12398,N_15069);
nand U16248 (N_16248,N_15283,N_14628);
and U16249 (N_16249,N_13740,N_15496);
xor U16250 (N_16250,N_14945,N_12629);
or U16251 (N_16251,N_13385,N_12371);
xor U16252 (N_16252,N_13447,N_15182);
or U16253 (N_16253,N_14433,N_13357);
or U16254 (N_16254,N_13818,N_13341);
nand U16255 (N_16255,N_15560,N_14208);
nor U16256 (N_16256,N_15881,N_13227);
and U16257 (N_16257,N_13417,N_15277);
nand U16258 (N_16258,N_13212,N_15866);
nand U16259 (N_16259,N_15833,N_14658);
xor U16260 (N_16260,N_13160,N_12589);
nand U16261 (N_16261,N_14244,N_13543);
nand U16262 (N_16262,N_15338,N_14646);
or U16263 (N_16263,N_12906,N_12898);
or U16264 (N_16264,N_15603,N_12261);
nand U16265 (N_16265,N_12307,N_14719);
nor U16266 (N_16266,N_13929,N_13503);
and U16267 (N_16267,N_13245,N_15882);
nand U16268 (N_16268,N_12410,N_14196);
nand U16269 (N_16269,N_13966,N_14911);
and U16270 (N_16270,N_15934,N_15303);
and U16271 (N_16271,N_13177,N_12754);
nor U16272 (N_16272,N_14810,N_12486);
xnor U16273 (N_16273,N_15860,N_13842);
xnor U16274 (N_16274,N_13728,N_12192);
or U16275 (N_16275,N_12360,N_12565);
nor U16276 (N_16276,N_14807,N_12795);
nand U16277 (N_16277,N_14394,N_13115);
nand U16278 (N_16278,N_15125,N_13862);
nor U16279 (N_16279,N_14974,N_13393);
xor U16280 (N_16280,N_13494,N_12548);
nand U16281 (N_16281,N_14227,N_14873);
nand U16282 (N_16282,N_12197,N_13584);
or U16283 (N_16283,N_12553,N_13775);
and U16284 (N_16284,N_13681,N_14068);
nand U16285 (N_16285,N_13579,N_12157);
or U16286 (N_16286,N_12978,N_14152);
and U16287 (N_16287,N_14434,N_15904);
xnor U16288 (N_16288,N_14330,N_14423);
nand U16289 (N_16289,N_12608,N_13667);
nor U16290 (N_16290,N_13785,N_13019);
xnor U16291 (N_16291,N_12673,N_14903);
nor U16292 (N_16292,N_14526,N_15485);
xor U16293 (N_16293,N_14824,N_12882);
nor U16294 (N_16294,N_14684,N_14150);
and U16295 (N_16295,N_14225,N_13386);
nor U16296 (N_16296,N_14705,N_15526);
nand U16297 (N_16297,N_13403,N_15240);
nand U16298 (N_16298,N_15816,N_13318);
xor U16299 (N_16299,N_15286,N_14073);
xor U16300 (N_16300,N_12231,N_12385);
nor U16301 (N_16301,N_12837,N_15628);
xnor U16302 (N_16302,N_15927,N_15502);
nor U16303 (N_16303,N_12075,N_13161);
and U16304 (N_16304,N_12436,N_15317);
or U16305 (N_16305,N_13745,N_14901);
nor U16306 (N_16306,N_15453,N_14459);
xor U16307 (N_16307,N_14417,N_13289);
or U16308 (N_16308,N_13232,N_15296);
nor U16309 (N_16309,N_12050,N_13083);
nor U16310 (N_16310,N_14981,N_12394);
or U16311 (N_16311,N_12810,N_12987);
or U16312 (N_16312,N_13768,N_12063);
and U16313 (N_16313,N_15461,N_14801);
or U16314 (N_16314,N_15251,N_12011);
or U16315 (N_16315,N_15962,N_12777);
nor U16316 (N_16316,N_15826,N_14552);
or U16317 (N_16317,N_13226,N_12132);
or U16318 (N_16318,N_14616,N_14179);
and U16319 (N_16319,N_13576,N_15365);
or U16320 (N_16320,N_15233,N_14884);
and U16321 (N_16321,N_12223,N_15585);
and U16322 (N_16322,N_15372,N_12220);
xor U16323 (N_16323,N_12494,N_12870);
nand U16324 (N_16324,N_13216,N_15150);
and U16325 (N_16325,N_15380,N_15511);
or U16326 (N_16326,N_12304,N_12847);
nand U16327 (N_16327,N_13034,N_15216);
nand U16328 (N_16328,N_13538,N_12679);
and U16329 (N_16329,N_15713,N_15612);
xor U16330 (N_16330,N_13732,N_15699);
or U16331 (N_16331,N_14764,N_13591);
nor U16332 (N_16332,N_12954,N_14307);
xor U16333 (N_16333,N_13037,N_12415);
nand U16334 (N_16334,N_14878,N_14070);
and U16335 (N_16335,N_12124,N_13597);
or U16336 (N_16336,N_12321,N_15337);
or U16337 (N_16337,N_13056,N_13537);
xnor U16338 (N_16338,N_15982,N_15712);
and U16339 (N_16339,N_12109,N_14597);
and U16340 (N_16340,N_14941,N_14483);
and U16341 (N_16341,N_15542,N_15989);
xnor U16342 (N_16342,N_12049,N_12708);
nand U16343 (N_16343,N_15340,N_15590);
or U16344 (N_16344,N_12684,N_13713);
xnor U16345 (N_16345,N_15444,N_13223);
nand U16346 (N_16346,N_14204,N_13332);
nor U16347 (N_16347,N_12479,N_13269);
or U16348 (N_16348,N_12339,N_14427);
nand U16349 (N_16349,N_12260,N_15659);
nand U16350 (N_16350,N_12040,N_15215);
nor U16351 (N_16351,N_12583,N_14026);
nand U16352 (N_16352,N_12704,N_13737);
xnor U16353 (N_16353,N_15429,N_14014);
nor U16354 (N_16354,N_12566,N_14780);
and U16355 (N_16355,N_12427,N_14462);
xnor U16356 (N_16356,N_15727,N_13182);
and U16357 (N_16357,N_15394,N_14439);
nand U16358 (N_16358,N_13259,N_12460);
nor U16359 (N_16359,N_14484,N_13355);
nor U16360 (N_16360,N_15274,N_12739);
or U16361 (N_16361,N_13982,N_13938);
nor U16362 (N_16362,N_14285,N_14933);
nor U16363 (N_16363,N_13840,N_15745);
nor U16364 (N_16364,N_15486,N_12580);
nor U16365 (N_16365,N_13159,N_13476);
xnor U16366 (N_16366,N_15166,N_13190);
nand U16367 (N_16367,N_12077,N_13889);
or U16368 (N_16368,N_13933,N_14021);
nor U16369 (N_16369,N_15836,N_14979);
nor U16370 (N_16370,N_12748,N_15008);
xnor U16371 (N_16371,N_15152,N_14841);
or U16372 (N_16372,N_15722,N_13726);
nor U16373 (N_16373,N_15643,N_12648);
nand U16374 (N_16374,N_14232,N_13120);
and U16375 (N_16375,N_13716,N_15581);
and U16376 (N_16376,N_13793,N_12868);
xnor U16377 (N_16377,N_12771,N_15877);
and U16378 (N_16378,N_14722,N_13770);
nor U16379 (N_16379,N_13780,N_14826);
nor U16380 (N_16380,N_15774,N_14482);
xor U16381 (N_16381,N_13354,N_14337);
nand U16382 (N_16382,N_13396,N_15864);
nand U16383 (N_16383,N_12358,N_14596);
nand U16384 (N_16384,N_14231,N_15958);
and U16385 (N_16385,N_13528,N_12655);
xnor U16386 (N_16386,N_13890,N_12359);
xnor U16387 (N_16387,N_15858,N_14235);
or U16388 (N_16388,N_13063,N_13719);
or U16389 (N_16389,N_12068,N_12105);
nand U16390 (N_16390,N_14266,N_15110);
and U16391 (N_16391,N_15550,N_13804);
or U16392 (N_16392,N_12502,N_14002);
and U16393 (N_16393,N_14752,N_12959);
or U16394 (N_16394,N_12137,N_13850);
nor U16395 (N_16395,N_14924,N_13474);
or U16396 (N_16396,N_12043,N_14061);
or U16397 (N_16397,N_13024,N_14737);
nor U16398 (N_16398,N_12276,N_14575);
nor U16399 (N_16399,N_15767,N_14239);
nor U16400 (N_16400,N_15800,N_12952);
and U16401 (N_16401,N_14532,N_13917);
nand U16402 (N_16402,N_12852,N_13328);
nor U16403 (N_16403,N_14121,N_15464);
xor U16404 (N_16404,N_12760,N_15799);
xnor U16405 (N_16405,N_14112,N_13137);
nor U16406 (N_16406,N_15097,N_13086);
and U16407 (N_16407,N_13696,N_14604);
or U16408 (N_16408,N_13028,N_14855);
nand U16409 (N_16409,N_14323,N_15992);
nand U16410 (N_16410,N_14881,N_15301);
nor U16411 (N_16411,N_15798,N_13683);
and U16412 (N_16412,N_13184,N_14891);
xnor U16413 (N_16413,N_12538,N_13942);
xnor U16414 (N_16414,N_14543,N_12440);
and U16415 (N_16415,N_14487,N_15527);
nor U16416 (N_16416,N_13265,N_13032);
xnor U16417 (N_16417,N_12179,N_15928);
nor U16418 (N_16418,N_15557,N_15462);
and U16419 (N_16419,N_13651,N_12728);
nand U16420 (N_16420,N_15672,N_14113);
nand U16421 (N_16421,N_13910,N_15687);
or U16422 (N_16422,N_14830,N_15533);
nor U16423 (N_16423,N_13119,N_13413);
xnor U16424 (N_16424,N_14390,N_12667);
or U16425 (N_16425,N_12849,N_14666);
nand U16426 (N_16426,N_15544,N_14064);
or U16427 (N_16427,N_15259,N_15222);
nor U16428 (N_16428,N_15054,N_15137);
xnor U16429 (N_16429,N_13428,N_14441);
nand U16430 (N_16430,N_14019,N_15611);
nor U16431 (N_16431,N_13859,N_13794);
nand U16432 (N_16432,N_14403,N_15041);
or U16433 (N_16433,N_12251,N_12807);
nor U16434 (N_16434,N_14261,N_15878);
nor U16435 (N_16435,N_13313,N_13158);
nor U16436 (N_16436,N_13278,N_14360);
or U16437 (N_16437,N_12155,N_13983);
nor U16438 (N_16438,N_13408,N_15680);
nor U16439 (N_16439,N_14522,N_14291);
or U16440 (N_16440,N_13058,N_13676);
or U16441 (N_16441,N_12725,N_15578);
or U16442 (N_16442,N_14382,N_15163);
and U16443 (N_16443,N_15640,N_13834);
nor U16444 (N_16444,N_15294,N_14724);
nand U16445 (N_16445,N_12211,N_12450);
and U16446 (N_16446,N_12712,N_15371);
and U16447 (N_16447,N_12832,N_14030);
or U16448 (N_16448,N_13645,N_13026);
nor U16449 (N_16449,N_12250,N_14212);
nor U16450 (N_16450,N_14410,N_15539);
and U16451 (N_16451,N_14055,N_14111);
nand U16452 (N_16452,N_14745,N_15105);
or U16453 (N_16453,N_14844,N_13122);
nand U16454 (N_16454,N_13327,N_12975);
nand U16455 (N_16455,N_13331,N_14516);
nor U16456 (N_16456,N_14518,N_13451);
or U16457 (N_16457,N_13935,N_13449);
nand U16458 (N_16458,N_13639,N_14688);
xnor U16459 (N_16459,N_14971,N_13883);
or U16460 (N_16460,N_12446,N_12625);
and U16461 (N_16461,N_13060,N_14601);
nand U16462 (N_16462,N_15683,N_12724);
or U16463 (N_16463,N_14707,N_15599);
or U16464 (N_16464,N_14284,N_13751);
xor U16465 (N_16465,N_12853,N_13249);
xnor U16466 (N_16466,N_12758,N_15756);
nor U16467 (N_16467,N_13303,N_13358);
or U16468 (N_16468,N_13629,N_15378);
and U16469 (N_16469,N_13673,N_15794);
or U16470 (N_16470,N_15029,N_15996);
and U16471 (N_16471,N_15295,N_15980);
nand U16472 (N_16472,N_14980,N_12503);
xnor U16473 (N_16473,N_15200,N_14007);
and U16474 (N_16474,N_12258,N_14286);
nand U16475 (N_16475,N_13471,N_15503);
and U16476 (N_16476,N_12595,N_14573);
nor U16477 (N_16477,N_13766,N_14372);
or U16478 (N_16478,N_14367,N_13373);
nand U16479 (N_16479,N_14910,N_13599);
or U16480 (N_16480,N_13087,N_13435);
or U16481 (N_16481,N_13192,N_13545);
and U16482 (N_16482,N_14751,N_12914);
nor U16483 (N_16483,N_15268,N_14593);
or U16484 (N_16484,N_14438,N_12692);
or U16485 (N_16485,N_14275,N_12805);
or U16486 (N_16486,N_14219,N_15717);
nand U16487 (N_16487,N_15734,N_15061);
and U16488 (N_16488,N_15447,N_15078);
nand U16489 (N_16489,N_12004,N_12230);
xor U16490 (N_16490,N_15117,N_13590);
and U16491 (N_16491,N_12312,N_14299);
nand U16492 (N_16492,N_15673,N_13071);
xor U16493 (N_16493,N_12229,N_13181);
nor U16494 (N_16494,N_12469,N_12800);
xor U16495 (N_16495,N_13166,N_12279);
and U16496 (N_16496,N_14466,N_15537);
xor U16497 (N_16497,N_15210,N_12598);
or U16498 (N_16498,N_12632,N_13479);
xor U16499 (N_16499,N_13200,N_15059);
xnor U16500 (N_16500,N_15281,N_12036);
xor U16501 (N_16501,N_15315,N_12735);
xor U16502 (N_16502,N_12609,N_15554);
or U16503 (N_16503,N_13536,N_13175);
nor U16504 (N_16504,N_14265,N_13779);
and U16505 (N_16505,N_13687,N_14294);
xnor U16506 (N_16506,N_15589,N_14877);
nand U16507 (N_16507,N_14887,N_13424);
and U16508 (N_16508,N_12815,N_13207);
and U16509 (N_16509,N_12059,N_13575);
or U16510 (N_16510,N_14016,N_14156);
and U16511 (N_16511,N_14600,N_12055);
nor U16512 (N_16512,N_15467,N_14968);
xnor U16513 (N_16513,N_15616,N_14270);
xor U16514 (N_16514,N_13438,N_13825);
nand U16515 (N_16515,N_13572,N_13755);
or U16516 (N_16516,N_14726,N_15474);
nand U16517 (N_16517,N_14488,N_15543);
or U16518 (N_16518,N_12341,N_15026);
or U16519 (N_16519,N_14925,N_12869);
and U16520 (N_16520,N_15761,N_12348);
xor U16521 (N_16521,N_15027,N_12579);
and U16522 (N_16522,N_14897,N_12156);
or U16523 (N_16523,N_15239,N_12710);
and U16524 (N_16524,N_14426,N_15108);
nor U16525 (N_16525,N_13241,N_15964);
and U16526 (N_16526,N_15497,N_13743);
nand U16527 (N_16527,N_14723,N_12628);
nor U16528 (N_16528,N_12647,N_12829);
and U16529 (N_16529,N_12738,N_14804);
nand U16530 (N_16530,N_15751,N_13510);
and U16531 (N_16531,N_15346,N_13727);
and U16532 (N_16532,N_14066,N_13231);
nand U16533 (N_16533,N_15688,N_14808);
xnor U16534 (N_16534,N_12021,N_14678);
nor U16535 (N_16535,N_14775,N_12025);
and U16536 (N_16536,N_15823,N_15050);
xor U16537 (N_16537,N_15991,N_14765);
nand U16538 (N_16538,N_14076,N_12791);
or U16539 (N_16539,N_12133,N_15993);
and U16540 (N_16540,N_15949,N_14645);
and U16541 (N_16541,N_13551,N_12093);
nor U16542 (N_16542,N_13668,N_14361);
and U16543 (N_16543,N_15450,N_15977);
or U16544 (N_16544,N_13940,N_12005);
xnor U16545 (N_16545,N_13778,N_15985);
nand U16546 (N_16546,N_15235,N_15261);
and U16547 (N_16547,N_13070,N_14332);
nor U16548 (N_16548,N_15179,N_15057);
nand U16549 (N_16549,N_12222,N_15884);
nand U16550 (N_16550,N_13901,N_15735);
or U16551 (N_16551,N_15142,N_15647);
and U16552 (N_16552,N_15999,N_12639);
and U16553 (N_16553,N_13379,N_14044);
nand U16554 (N_16554,N_12956,N_15249);
xnor U16555 (N_16555,N_13544,N_14770);
or U16556 (N_16556,N_15285,N_15813);
nor U16557 (N_16557,N_12325,N_15623);
and U16558 (N_16558,N_15409,N_13628);
or U16559 (N_16559,N_13453,N_13944);
xnor U16560 (N_16560,N_14861,N_12064);
nand U16561 (N_16561,N_15838,N_13348);
or U16562 (N_16562,N_13981,N_15482);
nand U16563 (N_16563,N_14936,N_14714);
xor U16564 (N_16564,N_15308,N_12799);
xor U16565 (N_16565,N_13364,N_14514);
nand U16566 (N_16566,N_12096,N_14036);
nor U16567 (N_16567,N_13796,N_14736);
or U16568 (N_16568,N_13362,N_12443);
and U16569 (N_16569,N_14712,N_13523);
and U16570 (N_16570,N_15755,N_12722);
nor U16571 (N_16571,N_12300,N_15390);
nor U16572 (N_16572,N_13875,N_12426);
nand U16573 (N_16573,N_15370,N_15602);
and U16574 (N_16574,N_14799,N_15411);
nor U16575 (N_16575,N_13876,N_15704);
or U16576 (N_16576,N_13763,N_12516);
and U16577 (N_16577,N_12509,N_14000);
or U16578 (N_16578,N_13627,N_12582);
xnor U16579 (N_16579,N_15957,N_14260);
and U16580 (N_16580,N_14398,N_14769);
or U16581 (N_16581,N_14165,N_14210);
or U16582 (N_16582,N_12500,N_13703);
nor U16583 (N_16583,N_12395,N_12287);
nor U16584 (N_16584,N_13626,N_14568);
xor U16585 (N_16585,N_13984,N_12383);
and U16586 (N_16586,N_14200,N_15121);
nand U16587 (N_16587,N_12255,N_13172);
nor U16588 (N_16588,N_15809,N_13493);
or U16589 (N_16589,N_12422,N_14610);
xnor U16590 (N_16590,N_15103,N_12788);
xor U16591 (N_16591,N_12969,N_15347);
nand U16592 (N_16592,N_15410,N_14004);
nor U16593 (N_16593,N_14402,N_14035);
and U16594 (N_16594,N_12861,N_14137);
or U16595 (N_16595,N_12232,N_15898);
xnor U16596 (N_16596,N_12988,N_12941);
or U16597 (N_16597,N_13144,N_12122);
nor U16598 (N_16598,N_15430,N_15046);
and U16599 (N_16599,N_12591,N_13592);
nor U16600 (N_16600,N_15588,N_13416);
xnor U16601 (N_16601,N_12154,N_12575);
xor U16602 (N_16602,N_14760,N_15060);
or U16603 (N_16603,N_15568,N_13853);
xnor U16604 (N_16604,N_14148,N_12564);
and U16605 (N_16605,N_13769,N_12148);
xor U16606 (N_16606,N_14930,N_14776);
nand U16607 (N_16607,N_13210,N_14655);
nor U16608 (N_16608,N_12835,N_15737);
nor U16609 (N_16609,N_12209,N_14768);
xor U16610 (N_16610,N_12848,N_12958);
or U16611 (N_16611,N_15875,N_12449);
xnor U16612 (N_16612,N_14084,N_15413);
xnor U16613 (N_16613,N_13887,N_14325);
nand U16614 (N_16614,N_12578,N_15570);
xnor U16615 (N_16615,N_13228,N_12615);
nor U16616 (N_16616,N_14695,N_12114);
or U16617 (N_16617,N_15574,N_13650);
or U16618 (N_16618,N_13296,N_15698);
xnor U16619 (N_16619,N_14343,N_13637);
and U16620 (N_16620,N_13155,N_13511);
nand U16621 (N_16621,N_12412,N_13174);
nand U16622 (N_16622,N_12239,N_15990);
xor U16623 (N_16623,N_15610,N_12904);
and U16624 (N_16624,N_12813,N_13618);
nor U16625 (N_16625,N_15534,N_13243);
and U16626 (N_16626,N_15473,N_12850);
xnor U16627 (N_16627,N_14889,N_12496);
nor U16628 (N_16628,N_14023,N_13797);
nand U16629 (N_16629,N_14772,N_13084);
or U16630 (N_16630,N_12296,N_13475);
or U16631 (N_16631,N_13061,N_14521);
nor U16632 (N_16632,N_15128,N_15652);
nand U16633 (N_16633,N_15065,N_15714);
or U16634 (N_16634,N_13855,N_15772);
nand U16635 (N_16635,N_12828,N_14194);
or U16636 (N_16636,N_15493,N_13412);
xnor U16637 (N_16637,N_12685,N_15076);
nand U16638 (N_16638,N_15983,N_14511);
xor U16639 (N_16639,N_13079,N_14233);
xor U16640 (N_16640,N_13350,N_13907);
xnor U16641 (N_16641,N_13015,N_14213);
nand U16642 (N_16642,N_12163,N_13167);
and U16643 (N_16643,N_14908,N_14672);
xor U16644 (N_16644,N_15155,N_15897);
nor U16645 (N_16645,N_14304,N_15677);
xor U16646 (N_16646,N_12263,N_13099);
and U16647 (N_16647,N_13047,N_13491);
or U16648 (N_16648,N_14428,N_12245);
nand U16649 (N_16649,N_15401,N_12473);
and U16650 (N_16650,N_12676,N_12113);
nand U16651 (N_16651,N_15837,N_12083);
or U16652 (N_16652,N_12159,N_15819);
nand U16653 (N_16653,N_12019,N_13811);
and U16654 (N_16654,N_14943,N_12962);
nand U16655 (N_16655,N_14253,N_13678);
xor U16656 (N_16656,N_15976,N_12046);
nor U16657 (N_16657,N_15252,N_14288);
or U16658 (N_16658,N_14366,N_13445);
nand U16659 (N_16659,N_13022,N_14094);
nand U16660 (N_16660,N_15242,N_12768);
xor U16661 (N_16661,N_13415,N_13053);
nor U16662 (N_16662,N_15626,N_13039);
and U16663 (N_16663,N_13490,N_15019);
xnor U16664 (N_16664,N_12928,N_14101);
nor U16665 (N_16665,N_12984,N_14734);
nor U16666 (N_16666,N_15270,N_15386);
xor U16667 (N_16667,N_15618,N_13286);
and U16668 (N_16668,N_12607,N_12621);
and U16669 (N_16669,N_15948,N_14781);
nand U16670 (N_16670,N_13540,N_13598);
and U16671 (N_16671,N_12207,N_14882);
nand U16672 (N_16672,N_12792,N_14762);
and U16673 (N_16673,N_14740,N_12072);
nor U16674 (N_16674,N_12544,N_12491);
and U16675 (N_16675,N_14129,N_12176);
or U16676 (N_16676,N_13430,N_14031);
nor U16677 (N_16677,N_13139,N_15495);
nand U16678 (N_16678,N_14883,N_15333);
and U16679 (N_16679,N_15869,N_15186);
and U16680 (N_16680,N_13867,N_15143);
nor U16681 (N_16681,N_14674,N_12401);
nor U16682 (N_16682,N_15801,N_14037);
or U16683 (N_16683,N_15786,N_14351);
nand U16684 (N_16684,N_15929,N_14756);
nand U16685 (N_16685,N_15556,N_14188);
nand U16686 (N_16686,N_15322,N_13515);
or U16687 (N_16687,N_15571,N_13273);
nand U16688 (N_16688,N_15318,N_15419);
nor U16689 (N_16689,N_14879,N_15420);
and U16690 (N_16690,N_15540,N_13632);
xor U16691 (N_16691,N_14081,N_14985);
or U16692 (N_16692,N_13219,N_13457);
nand U16693 (N_16693,N_13788,N_13869);
nand U16694 (N_16694,N_14995,N_12606);
and U16695 (N_16695,N_15729,N_15941);
and U16696 (N_16696,N_13525,N_15955);
nand U16697 (N_16697,N_14972,N_12447);
nand U16698 (N_16698,N_15953,N_12657);
nand U16699 (N_16699,N_13903,N_15170);
and U16700 (N_16700,N_15700,N_13969);
or U16701 (N_16701,N_15805,N_14020);
and U16702 (N_16702,N_13631,N_13622);
and U16703 (N_16703,N_15891,N_13153);
or U16704 (N_16704,N_14116,N_13817);
or U16705 (N_16705,N_14130,N_12425);
nor U16706 (N_16706,N_15691,N_12688);
xor U16707 (N_16707,N_15431,N_13235);
nor U16708 (N_16708,N_15476,N_15083);
nand U16709 (N_16709,N_13301,N_13314);
and U16710 (N_16710,N_13643,N_14926);
xor U16711 (N_16711,N_14411,N_14539);
or U16712 (N_16712,N_12790,N_12855);
xor U16713 (N_16713,N_12687,N_15523);
xor U16714 (N_16714,N_12883,N_14766);
and U16715 (N_16715,N_12617,N_12471);
xnor U16716 (N_16716,N_13847,N_15392);
and U16717 (N_16717,N_14414,N_14976);
and U16718 (N_16718,N_13011,N_14949);
nor U16719 (N_16719,N_14322,N_13246);
or U16720 (N_16720,N_12069,N_13501);
xnor U16721 (N_16721,N_15703,N_13095);
nor U16722 (N_16722,N_12666,N_14958);
xnor U16723 (N_16723,N_12149,N_13140);
and U16724 (N_16724,N_13504,N_15047);
nand U16725 (N_16725,N_14595,N_12561);
and U16726 (N_16726,N_14124,N_13298);
or U16727 (N_16727,N_13281,N_13997);
nand U16728 (N_16728,N_15454,N_15995);
or U16729 (N_16729,N_15566,N_14224);
xnor U16730 (N_16730,N_14099,N_14676);
nor U16731 (N_16731,N_13027,N_15650);
xor U16732 (N_16732,N_12593,N_12481);
or U16733 (N_16733,N_14978,N_15359);
nand U16734 (N_16734,N_15975,N_14956);
nor U16735 (N_16735,N_13459,N_15908);
or U16736 (N_16736,N_12060,N_13244);
and U16737 (N_16737,N_13894,N_15009);
nand U16738 (N_16738,N_14267,N_12274);
nand U16739 (N_16739,N_12827,N_15202);
xor U16740 (N_16740,N_12399,N_15903);
or U16741 (N_16741,N_13444,N_15739);
nand U16742 (N_16742,N_12405,N_13835);
nor U16743 (N_16743,N_13076,N_15243);
or U16744 (N_16744,N_12125,N_14317);
and U16745 (N_16745,N_14153,N_15917);
and U16746 (N_16746,N_14562,N_15368);
nand U16747 (N_16747,N_12567,N_14965);
nor U16748 (N_16748,N_13805,N_12062);
nand U16749 (N_16749,N_14970,N_15293);
nand U16750 (N_16750,N_15250,N_12989);
nor U16751 (N_16751,N_13764,N_14086);
or U16752 (N_16752,N_15457,N_13530);
xor U16753 (N_16753,N_12784,N_14315);
xor U16754 (N_16754,N_12661,N_14389);
nor U16755 (N_16755,N_13669,N_13337);
nor U16756 (N_16756,N_14505,N_13387);
and U16757 (N_16757,N_13772,N_14457);
xor U16758 (N_16758,N_12282,N_14866);
nand U16759 (N_16759,N_12912,N_13469);
or U16760 (N_16760,N_13977,N_13571);
xnor U16761 (N_16761,N_12680,N_15886);
or U16762 (N_16762,N_14147,N_12387);
and U16763 (N_16763,N_15376,N_12977);
nor U16764 (N_16764,N_15830,N_13085);
xnor U16765 (N_16765,N_14173,N_12092);
nor U16766 (N_16766,N_15824,N_15959);
nor U16767 (N_16767,N_14577,N_13864);
nor U16768 (N_16768,N_12783,N_12823);
nor U16769 (N_16769,N_13959,N_14090);
nand U16770 (N_16770,N_14131,N_12967);
nor U16771 (N_16771,N_13878,N_14157);
and U16772 (N_16772,N_13382,N_12836);
nand U16773 (N_16773,N_12737,N_14193);
nand U16774 (N_16774,N_14120,N_13383);
or U16775 (N_16775,N_13436,N_15984);
and U16776 (N_16776,N_14185,N_15184);
or U16777 (N_16777,N_15489,N_12168);
nor U16778 (N_16778,N_14444,N_14544);
nand U16779 (N_16779,N_13257,N_15532);
and U16780 (N_16780,N_12134,N_12150);
nand U16781 (N_16781,N_12029,N_14393);
nor U16782 (N_16782,N_13829,N_13879);
xor U16783 (N_16783,N_14599,N_12284);
or U16784 (N_16784,N_12356,N_12699);
or U16785 (N_16785,N_14062,N_14347);
or U16786 (N_16786,N_12218,N_13881);
nor U16787 (N_16787,N_13675,N_14838);
or U16788 (N_16788,N_14038,N_13616);
and U16789 (N_16789,N_13517,N_13655);
nor U16790 (N_16790,N_12540,N_13513);
nor U16791 (N_16791,N_14327,N_14757);
or U16792 (N_16792,N_12386,N_14612);
nand U16793 (N_16793,N_12146,N_14822);
nor U16794 (N_16794,N_15406,N_15636);
and U16795 (N_16795,N_15649,N_12919);
and U16796 (N_16796,N_14336,N_12368);
or U16797 (N_16797,N_13723,N_12111);
nand U16798 (N_16798,N_12299,N_12199);
and U16799 (N_16799,N_15913,N_15038);
nand U16800 (N_16800,N_14477,N_14409);
and U16801 (N_16801,N_15192,N_12649);
nor U16802 (N_16802,N_12419,N_15922);
xor U16803 (N_16803,N_12390,N_12210);
or U16804 (N_16804,N_15920,N_15945);
nand U16805 (N_16805,N_14814,N_15100);
and U16806 (N_16806,N_13164,N_15591);
nand U16807 (N_16807,N_15067,N_12288);
nor U16808 (N_16808,N_14609,N_13326);
and U16809 (N_16809,N_12660,N_14048);
nand U16810 (N_16810,N_12178,N_14381);
and U16811 (N_16811,N_13113,N_15510);
and U16812 (N_16812,N_15499,N_15329);
and U16813 (N_16813,N_14585,N_13215);
nand U16814 (N_16814,N_13422,N_15887);
and U16815 (N_16815,N_15519,N_13695);
or U16816 (N_16816,N_15089,N_15263);
xnor U16817 (N_16817,N_15114,N_12677);
nor U16818 (N_16818,N_14311,N_14089);
nand U16819 (N_16819,N_12008,N_14443);
nor U16820 (N_16820,N_14110,N_14282);
nand U16821 (N_16821,N_13756,N_13434);
nand U16822 (N_16822,N_12703,N_12499);
nand U16823 (N_16823,N_12330,N_12926);
nor U16824 (N_16824,N_13208,N_14716);
xnor U16825 (N_16825,N_15345,N_14355);
nand U16826 (N_16826,N_13472,N_15943);
nor U16827 (N_16827,N_12670,N_12483);
or U16828 (N_16828,N_12999,N_14591);
or U16829 (N_16829,N_14711,N_15331);
and U16830 (N_16830,N_13625,N_14216);
and U16831 (N_16831,N_12252,N_15665);
or U16832 (N_16832,N_13845,N_15765);
and U16833 (N_16833,N_15583,N_12151);
nand U16834 (N_16834,N_15963,N_12373);
and U16835 (N_16835,N_12577,N_12597);
nand U16836 (N_16836,N_12672,N_15546);
or U16837 (N_16837,N_13880,N_13096);
xor U16838 (N_16838,N_12935,N_13958);
and U16839 (N_16839,N_14418,N_14374);
and U16840 (N_16840,N_12081,N_14542);
and U16841 (N_16841,N_15313,N_13217);
or U16842 (N_16842,N_12009,N_13483);
nor U16843 (N_16843,N_13254,N_15827);
or U16844 (N_16844,N_15880,N_12181);
nand U16845 (N_16845,N_14528,N_14664);
or U16846 (N_16846,N_12811,N_12319);
nand U16847 (N_16847,N_13400,N_14480);
and U16848 (N_16848,N_13360,N_13603);
nor U16849 (N_16849,N_14648,N_13957);
nand U16850 (N_16850,N_13548,N_13973);
xor U16851 (N_16851,N_15153,N_15549);
xnor U16852 (N_16852,N_14287,N_14472);
and U16853 (N_16853,N_15662,N_13931);
or U16854 (N_16854,N_13359,N_12851);
xnor U16855 (N_16855,N_13460,N_13539);
nor U16856 (N_16856,N_15164,N_15373);
and U16857 (N_16857,N_15940,N_13652);
or U16858 (N_16858,N_15879,N_13156);
nor U16859 (N_16859,N_14460,N_12880);
or U16860 (N_16860,N_15442,N_12525);
xnor U16861 (N_16861,N_14773,N_12472);
nor U16862 (N_16862,N_12173,N_13888);
nand U16863 (N_16863,N_13839,N_12022);
xnor U16864 (N_16864,N_13495,N_12857);
nor U16865 (N_16865,N_14611,N_14800);
nor U16866 (N_16866,N_14525,N_12886);
and U16867 (N_16867,N_13291,N_15225);
xor U16868 (N_16868,N_15156,N_14005);
nor U16869 (N_16869,N_14937,N_12318);
nand U16870 (N_16870,N_15789,N_14470);
xor U16871 (N_16871,N_15418,N_13522);
nor U16872 (N_16872,N_12537,N_13363);
nor U16873 (N_16873,N_12986,N_14733);
nand U16874 (N_16874,N_15960,N_15020);
and U16875 (N_16875,N_12007,N_14656);
or U16876 (N_16876,N_13419,N_14990);
or U16877 (N_16877,N_14862,N_13897);
nand U16878 (N_16878,N_12119,N_14540);
and U16879 (N_16879,N_14435,N_13055);
and U16880 (N_16880,N_13081,N_12142);
xor U16881 (N_16881,N_15582,N_13478);
nand U16882 (N_16882,N_14649,N_14132);
nand U16883 (N_16883,N_14310,N_14500);
xor U16884 (N_16884,N_14077,N_14888);
or U16885 (N_16885,N_15224,N_14160);
nor U16886 (N_16886,N_14564,N_14251);
nand U16887 (N_16887,N_12532,N_14630);
or U16888 (N_16888,N_12058,N_12918);
and U16889 (N_16889,N_13370,N_15037);
xor U16890 (N_16890,N_15625,N_13560);
or U16891 (N_16891,N_14725,N_12414);
and U16892 (N_16892,N_13283,N_12716);
nand U16893 (N_16893,N_15569,N_15312);
nand U16894 (N_16894,N_13371,N_12610);
nand U16895 (N_16895,N_12908,N_12226);
xnor U16896 (N_16896,N_13236,N_15515);
nor U16897 (N_16897,N_14297,N_14183);
and U16898 (N_16898,N_13418,N_14798);
or U16899 (N_16899,N_12878,N_15607);
nor U16900 (N_16900,N_15944,N_15804);
and U16901 (N_16901,N_13157,N_13861);
xor U16902 (N_16902,N_13697,N_14922);
xnor U16903 (N_16903,N_13762,N_14572);
or U16904 (N_16904,N_15825,N_14790);
nand U16905 (N_16905,N_12991,N_12164);
nor U16906 (N_16906,N_12528,N_13405);
or U16907 (N_16907,N_13771,N_14923);
xor U16908 (N_16908,N_15587,N_13928);
nor U16909 (N_16909,N_15101,N_14424);
nor U16910 (N_16910,N_13329,N_15504);
xor U16911 (N_16911,N_14217,N_14665);
xnor U16912 (N_16912,N_15230,N_12121);
nor U16913 (N_16913,N_15685,N_13963);
xor U16914 (N_16914,N_12968,N_13229);
or U16915 (N_16915,N_15226,N_14931);
nor U16916 (N_16916,N_15852,N_13518);
or U16917 (N_16917,N_12505,N_15971);
or U16918 (N_16918,N_12618,N_13814);
nand U16919 (N_16919,N_14638,N_13125);
xor U16920 (N_16920,N_14255,N_12108);
or U16921 (N_16921,N_15484,N_13514);
xnor U16922 (N_16922,N_14452,N_15862);
or U16923 (N_16923,N_15811,N_12600);
xor U16924 (N_16924,N_13506,N_14043);
xnor U16925 (N_16925,N_14947,N_15087);
xor U16926 (N_16926,N_14478,N_14637);
or U16927 (N_16927,N_13256,N_15828);
nand U16928 (N_16928,N_15802,N_12907);
nand U16929 (N_16929,N_12627,N_13725);
or U16930 (N_16930,N_14735,N_12714);
and U16931 (N_16931,N_12201,N_12881);
or U16932 (N_16932,N_15873,N_15449);
nand U16933 (N_16933,N_12435,N_15706);
nand U16934 (N_16934,N_15005,N_15330);
or U16935 (N_16935,N_13662,N_13659);
nor U16936 (N_16936,N_12778,N_15254);
nand U16937 (N_16937,N_13391,N_15205);
nor U16938 (N_16938,N_15440,N_12161);
xnor U16939 (N_16939,N_13437,N_14220);
nand U16940 (N_16940,N_13707,N_15855);
nand U16941 (N_16941,N_12826,N_14557);
nand U16942 (N_16942,N_13035,N_13986);
and U16943 (N_16943,N_13388,N_14118);
and U16944 (N_16944,N_15275,N_15521);
xor U16945 (N_16945,N_13607,N_13013);
nand U16946 (N_16946,N_12141,N_12418);
nor U16947 (N_16947,N_14034,N_14045);
and U16948 (N_16948,N_13925,N_14677);
or U16949 (N_16949,N_15421,N_13521);
xnor U16950 (N_16950,N_15391,N_12100);
and U16951 (N_16951,N_13205,N_14328);
xnor U16952 (N_16952,N_15781,N_15834);
or U16953 (N_16953,N_15782,N_13692);
nor U16954 (N_16954,N_14953,N_15645);
nor U16955 (N_16955,N_13657,N_15950);
xor U16956 (N_16956,N_12690,N_12900);
nand U16957 (N_16957,N_13554,N_15428);
or U16958 (N_16958,N_13321,N_15938);
and U16959 (N_16959,N_15693,N_15358);
nand U16960 (N_16960,N_14345,N_12316);
xnor U16961 (N_16961,N_15899,N_13248);
xor U16962 (N_16962,N_14690,N_12705);
and U16963 (N_16963,N_15092,N_14436);
xor U16964 (N_16964,N_13990,N_12342);
xor U16965 (N_16965,N_12445,N_15750);
nor U16966 (N_16966,N_15023,N_13123);
nor U16967 (N_16967,N_13347,N_14703);
nand U16968 (N_16968,N_14640,N_15981);
or U16969 (N_16969,N_13193,N_15353);
and U16970 (N_16970,N_12715,N_13030);
or U16971 (N_16971,N_12961,N_12556);
and U16972 (N_16972,N_15161,N_13976);
nand U16973 (N_16973,N_12295,N_13150);
nor U16974 (N_16974,N_12557,N_15744);
and U16975 (N_16975,N_13552,N_12053);
or U16976 (N_16976,N_13463,N_13660);
and U16977 (N_16977,N_12787,N_14512);
and U16978 (N_16978,N_13488,N_12637);
and U16979 (N_16979,N_12939,N_15228);
and U16980 (N_16980,N_14617,N_12090);
or U16981 (N_16981,N_12979,N_15635);
nor U16982 (N_16982,N_13774,N_15674);
or U16983 (N_16983,N_15807,N_14042);
nand U16984 (N_16984,N_13553,N_14149);
xnor U16985 (N_16985,N_15840,N_12519);
nor U16986 (N_16986,N_13820,N_13080);
and U16987 (N_16987,N_14742,N_15237);
xor U16988 (N_16988,N_13747,N_12018);
xor U16989 (N_16989,N_13753,N_14222);
or U16990 (N_16990,N_14708,N_13290);
and U16991 (N_16991,N_13425,N_15116);
nor U16992 (N_16992,N_12844,N_13705);
nor U16993 (N_16993,N_12052,N_13995);
nand U16994 (N_16994,N_15355,N_14559);
or U16995 (N_16995,N_15212,N_13720);
nor U16996 (N_16996,N_14468,N_15831);
xor U16997 (N_16997,N_13541,N_15111);
nor U16998 (N_16998,N_15853,N_13674);
and U16999 (N_16999,N_15458,N_13384);
or U17000 (N_17000,N_12213,N_13187);
xor U17001 (N_17001,N_13152,N_13294);
nand U17002 (N_17002,N_12079,N_15326);
nor U17003 (N_17003,N_15093,N_15624);
nand U17004 (N_17004,N_13399,N_12854);
xor U17005 (N_17005,N_12508,N_12614);
nor U17006 (N_17006,N_15352,N_15098);
nor U17007 (N_17007,N_13075,N_14471);
xor U17008 (N_17008,N_14915,N_12945);
nand U17009 (N_17009,N_15207,N_12572);
and U17010 (N_17010,N_14758,N_15034);
nand U17011 (N_17011,N_13918,N_13121);
nand U17012 (N_17012,N_13733,N_12972);
nand U17013 (N_17013,N_14992,N_15733);
nor U17014 (N_17014,N_14176,N_12921);
nand U17015 (N_17015,N_14163,N_15925);
or U17016 (N_17016,N_12315,N_12901);
xor U17017 (N_17017,N_13516,N_12601);
nand U17018 (N_17018,N_15577,N_13367);
and U17019 (N_17019,N_12010,N_14448);
and U17020 (N_17020,N_14324,N_14605);
nor U17021 (N_17021,N_12839,N_13909);
xor U17022 (N_17022,N_12028,N_12833);
xnor U17023 (N_17023,N_12765,N_12871);
nor U17024 (N_17024,N_15520,N_12118);
xnor U17025 (N_17025,N_12285,N_13104);
xnor U17026 (N_17026,N_14545,N_13135);
nand U17027 (N_17027,N_15189,N_14809);
and U17028 (N_17028,N_14006,N_13661);
nand U17029 (N_17029,N_15004,N_15961);
nor U17030 (N_17030,N_14453,N_14463);
nor U17031 (N_17031,N_13619,N_15193);
and U17032 (N_17032,N_14806,N_14983);
nand U17033 (N_17033,N_13040,N_13738);
nor U17034 (N_17034,N_13250,N_13752);
or U17035 (N_17035,N_14485,N_13724);
nand U17036 (N_17036,N_12895,N_13018);
or U17037 (N_17037,N_12943,N_13214);
or U17038 (N_17038,N_14964,N_14706);
xnor U17039 (N_17039,N_15481,N_12452);
and U17040 (N_17040,N_12397,N_12971);
nand U17041 (N_17041,N_12693,N_13188);
nand U17042 (N_17042,N_14138,N_13389);
or U17043 (N_17043,N_13440,N_13323);
and U17044 (N_17044,N_13531,N_15122);
and U17045 (N_17045,N_12602,N_15024);
nor U17046 (N_17046,N_12303,N_14182);
or U17047 (N_17047,N_12463,N_12305);
xnor U17048 (N_17048,N_15901,N_14919);
nand U17049 (N_17049,N_14041,N_14386);
and U17050 (N_17050,N_12464,N_12581);
nand U17051 (N_17051,N_13189,N_15682);
or U17052 (N_17052,N_15654,N_13280);
nand U17053 (N_17053,N_15169,N_14624);
nand U17054 (N_17054,N_15066,N_13589);
nor U17055 (N_17055,N_14181,N_13482);
xnor U17056 (N_17056,N_15821,N_13485);
or U17057 (N_17057,N_15140,N_12937);
nor U17058 (N_17058,N_14271,N_15416);
and U17059 (N_17059,N_14817,N_12970);
or U17060 (N_17060,N_15633,N_13807);
nor U17061 (N_17061,N_14510,N_14732);
nor U17062 (N_17062,N_12437,N_15874);
and U17063 (N_17063,N_13799,N_13234);
or U17064 (N_17064,N_14977,N_13961);
or U17065 (N_17065,N_15629,N_12981);
or U17066 (N_17066,N_15154,N_12310);
nand U17067 (N_17067,N_14159,N_15120);
and U17068 (N_17068,N_13608,N_14865);
xor U17069 (N_17069,N_13266,N_12286);
or U17070 (N_17070,N_15135,N_14854);
and U17071 (N_17071,N_15160,N_13293);
xor U17072 (N_17072,N_13131,N_15895);
xor U17073 (N_17073,N_13915,N_12138);
nor U17074 (N_17074,N_14569,N_13781);
and U17075 (N_17075,N_12909,N_15456);
nor U17076 (N_17076,N_15280,N_15930);
xor U17077 (N_17077,N_14912,N_12554);
and U17078 (N_17078,N_12929,N_15639);
xor U17079 (N_17079,N_14644,N_13653);
nand U17080 (N_17080,N_14820,N_12552);
nand U17081 (N_17081,N_15262,N_12997);
and U17082 (N_17082,N_15051,N_13206);
and U17083 (N_17083,N_13685,N_13455);
nor U17084 (N_17084,N_12297,N_13806);
and U17085 (N_17085,N_15145,N_14364);
nor U17086 (N_17086,N_13004,N_15753);
or U17087 (N_17087,N_12186,N_15516);
or U17088 (N_17088,N_13380,N_15348);
nand U17089 (N_17089,N_12535,N_14392);
nand U17090 (N_17090,N_14680,N_12262);
nor U17091 (N_17091,N_15690,N_15718);
and U17092 (N_17092,N_13492,N_15932);
nor U17093 (N_17093,N_15305,N_12104);
xor U17094 (N_17094,N_12495,N_15664);
nand U17095 (N_17095,N_15282,N_14009);
nand U17096 (N_17096,N_15783,N_15919);
nor U17097 (N_17097,N_15675,N_15528);
nand U17098 (N_17098,N_14784,N_13837);
nor U17099 (N_17099,N_12650,N_14123);
nor U17100 (N_17100,N_13218,N_15375);
and U17101 (N_17101,N_13467,N_14701);
nand U17102 (N_17102,N_13320,N_14948);
and U17103 (N_17103,N_12017,N_14104);
xor U17104 (N_17104,N_13999,N_15594);
or U17105 (N_17105,N_15012,N_15535);
nand U17106 (N_17106,N_15195,N_13271);
and U17107 (N_17107,N_14370,N_15551);
and U17108 (N_17108,N_14218,N_14223);
nand U17109 (N_17109,N_12729,N_14916);
nor U17110 (N_17110,N_15541,N_13310);
or U17111 (N_17111,N_13198,N_15374);
xnor U17112 (N_17112,N_14845,N_13285);
xor U17113 (N_17113,N_14508,N_13109);
nor U17114 (N_17114,N_12539,N_12730);
or U17115 (N_17115,N_12116,N_12185);
or U17116 (N_17116,N_14553,N_13872);
xor U17117 (N_17117,N_15494,N_15091);
nor U17118 (N_17118,N_14761,N_14391);
nand U17119 (N_17119,N_14242,N_14667);
xor U17120 (N_17120,N_12786,N_13126);
nand U17121 (N_17121,N_15472,N_13843);
and U17122 (N_17122,N_14234,N_12433);
or U17123 (N_17123,N_12382,N_15780);
and U17124 (N_17124,N_15081,N_15797);
or U17125 (N_17125,N_15902,N_14008);
xnor U17126 (N_17126,N_14461,N_12165);
nand U17127 (N_17127,N_12513,N_15035);
xnor U17128 (N_17128,N_14523,N_12596);
nor U17129 (N_17129,N_12248,N_15605);
nand U17130 (N_17130,N_15994,N_14350);
or U17131 (N_17131,N_12665,N_12353);
xnor U17132 (N_17132,N_14900,N_12476);
and U17133 (N_17133,N_14633,N_12555);
xnor U17134 (N_17134,N_15396,N_13595);
nand U17135 (N_17135,N_15785,N_12003);
xor U17136 (N_17136,N_14075,N_12272);
or U17137 (N_17137,N_12188,N_14847);
or U17138 (N_17138,N_12254,N_12372);
nor U17139 (N_17139,N_13580,N_14580);
or U17140 (N_17140,N_14258,N_13439);
and U17141 (N_17141,N_15138,N_14920);
xnor U17142 (N_17142,N_15385,N_14944);
or U17143 (N_17143,N_15432,N_14314);
nand U17144 (N_17144,N_14993,N_15084);
nand U17145 (N_17145,N_13644,N_15399);
and U17146 (N_17146,N_14748,N_13711);
nor U17147 (N_17147,N_13563,N_15307);
nand U17148 (N_17148,N_13706,N_13021);
or U17149 (N_17149,N_12189,N_12037);
nand U17150 (N_17150,N_15477,N_12761);
or U17151 (N_17151,N_15016,N_14904);
xor U17152 (N_17152,N_13106,N_14537);
nor U17153 (N_17153,N_15018,N_13905);
or U17154 (N_17154,N_14950,N_15298);
xnor U17155 (N_17155,N_13162,N_14375);
xor U17156 (N_17156,N_14024,N_12169);
and U17157 (N_17157,N_15253,N_12431);
xnor U17158 (N_17158,N_13377,N_13866);
and U17159 (N_17159,N_13721,N_15656);
xnor U17160 (N_17160,N_14467,N_12671);
xnor U17161 (N_17161,N_12298,N_13955);
xnor U17162 (N_17162,N_15657,N_15609);
or U17163 (N_17163,N_15695,N_15036);
or U17164 (N_17164,N_14549,N_13613);
nand U17165 (N_17165,N_12074,N_13366);
nand U17166 (N_17166,N_14080,N_12536);
or U17167 (N_17167,N_12487,N_12669);
or U17168 (N_17168,N_13486,N_13971);
nand U17169 (N_17169,N_14365,N_12948);
nor U17170 (N_17170,N_15788,N_15561);
nand U17171 (N_17171,N_13858,N_14241);
xor U17172 (N_17172,N_15658,N_12340);
or U17173 (N_17173,N_14437,N_13374);
nand U17174 (N_17174,N_12225,N_13636);
nor U17175 (N_17175,N_12713,N_14264);
xnor U17176 (N_17176,N_12320,N_14815);
xor U17177 (N_17177,N_14481,N_12753);
or U17178 (N_17178,N_14056,N_12940);
and U17179 (N_17179,N_13841,N_15620);
nor U17180 (N_17180,N_15670,N_15102);
and U17181 (N_17181,N_12027,N_13704);
or U17182 (N_17182,N_15071,N_15812);
xnor U17183 (N_17183,N_13555,N_15220);
nand U17184 (N_17184,N_13282,N_15383);
nor U17185 (N_17185,N_13268,N_14682);
and U17186 (N_17186,N_12012,N_13648);
or U17187 (N_17187,N_15918,N_15646);
nor U17188 (N_17188,N_15040,N_14079);
nand U17189 (N_17189,N_14362,N_15796);
and U17190 (N_17190,N_12428,N_14907);
nor U17191 (N_17191,N_14669,N_13934);
nor U17192 (N_17192,N_15586,N_12204);
nand U17193 (N_17193,N_14629,N_12757);
xor U17194 (N_17194,N_15856,N_15445);
xor U17195 (N_17195,N_15201,N_14289);
nor U17196 (N_17196,N_13962,N_14312);
nand U17197 (N_17197,N_14825,N_14383);
xor U17198 (N_17198,N_15829,N_13304);
or U17199 (N_17199,N_12966,N_14551);
nor U17200 (N_17200,N_13340,N_15219);
or U17201 (N_17201,N_12592,N_13017);
or U17202 (N_17202,N_14663,N_13031);
nand U17203 (N_17203,N_13677,N_14012);
nor U17204 (N_17204,N_13342,N_13604);
nand U17205 (N_17205,N_15000,N_14823);
xor U17206 (N_17206,N_13074,N_14849);
and U17207 (N_17207,N_13892,N_13251);
or U17208 (N_17208,N_15112,N_14960);
xnor U17209 (N_17209,N_15191,N_14519);
or U17210 (N_17210,N_12879,N_13988);
xor U17211 (N_17211,N_13621,N_13222);
xor U17212 (N_17212,N_12545,N_15165);
or U17213 (N_17213,N_14743,N_13920);
or U17214 (N_17214,N_14872,N_12308);
nor U17215 (N_17215,N_14127,N_12247);
xnor U17216 (N_17216,N_13520,N_14864);
xor U17217 (N_17217,N_12478,N_13974);
and U17218 (N_17218,N_12293,N_15621);
xnor U17219 (N_17219,N_12659,N_12143);
nor U17220 (N_17220,N_12466,N_14013);
and U17221 (N_17221,N_13170,N_12875);
and U17222 (N_17222,N_13441,N_13054);
or U17223 (N_17223,N_14771,N_15793);
nand U17224 (N_17224,N_13932,N_14498);
nand U17225 (N_17225,N_12172,N_12726);
nor U17226 (N_17226,N_12934,N_13786);
nand U17227 (N_17227,N_15405,N_13225);
nor U17228 (N_17228,N_15001,N_15475);
nor U17229 (N_17229,N_14791,N_12766);
nand U17230 (N_17230,N_12475,N_14371);
or U17231 (N_17231,N_13741,N_12242);
and U17232 (N_17232,N_13717,N_13558);
or U17233 (N_17233,N_12802,N_15309);
nor U17234 (N_17234,N_12423,N_14226);
nor U17235 (N_17235,N_13299,N_15090);
or U17236 (N_17236,N_13951,N_13312);
and U17237 (N_17237,N_14177,N_14746);
nand U17238 (N_17238,N_14494,N_13335);
nand U17239 (N_17239,N_14245,N_12369);
or U17240 (N_17240,N_12624,N_13496);
nor U17241 (N_17241,N_15032,N_12153);
xor U17242 (N_17242,N_13046,N_15641);
nand U17243 (N_17243,N_13828,N_12963);
and U17244 (N_17244,N_15709,N_13242);
nor U17245 (N_17245,N_12840,N_14834);
or U17246 (N_17246,N_14534,N_14100);
or U17247 (N_17247,N_15710,N_12322);
xor U17248 (N_17248,N_14060,N_14164);
and U17249 (N_17249,N_14563,N_13186);
xnor U17250 (N_17250,N_15565,N_14119);
nand U17251 (N_17251,N_15369,N_14091);
or U17252 (N_17252,N_13420,N_12086);
xor U17253 (N_17253,N_15492,N_12439);
xor U17254 (N_17254,N_13309,N_12750);
and U17255 (N_17255,N_15760,N_14991);
and U17256 (N_17256,N_14464,N_15393);
nor U17257 (N_17257,N_15584,N_15563);
nor U17258 (N_17258,N_15300,N_12559);
nand U17259 (N_17259,N_14205,N_15545);
nand U17260 (N_17260,N_15741,N_14909);
nand U17261 (N_17261,N_15213,N_15757);
xnor U17262 (N_17262,N_14699,N_13069);
and U17263 (N_17263,N_15148,N_14065);
xnor U17264 (N_17264,N_15167,N_15726);
nand U17265 (N_17265,N_15512,N_12355);
nand U17266 (N_17266,N_14476,N_12568);
or U17267 (N_17267,N_15870,N_13577);
nand U17268 (N_17268,N_13154,N_15175);
nor U17269 (N_17269,N_15273,N_15323);
or U17270 (N_17270,N_13307,N_15272);
and U17271 (N_17271,N_14700,N_14626);
xnor U17272 (N_17272,N_12709,N_14447);
nor U17273 (N_17273,N_15697,N_13993);
or U17274 (N_17274,N_13870,N_15407);
and U17275 (N_17275,N_13564,N_14507);
and U17276 (N_17276,N_13936,N_13410);
and U17277 (N_17277,N_12697,N_13171);
xor U17278 (N_17278,N_14513,N_14652);
nor U17279 (N_17279,N_15728,N_14727);
or U17280 (N_17280,N_14842,N_15185);
xor U17281 (N_17281,N_12400,N_13333);
or U17282 (N_17282,N_12171,N_13708);
xnor U17283 (N_17283,N_13023,N_14496);
nor U17284 (N_17284,N_13003,N_14687);
xor U17285 (N_17285,N_15096,N_15465);
nand U17286 (N_17286,N_13163,N_15839);
and U17287 (N_17287,N_15806,N_13006);
and U17288 (N_17288,N_15088,N_13815);
xnor U17289 (N_17289,N_15190,N_14619);
xnor U17290 (N_17290,N_15888,N_12531);
xor U17291 (N_17291,N_13556,N_14174);
xnor U17292 (N_17292,N_14209,N_15669);
nor U17293 (N_17293,N_13230,N_12611);
nor U17294 (N_17294,N_15436,N_13423);
nor U17295 (N_17295,N_14905,N_15762);
nand U17296 (N_17296,N_13679,N_15758);
or U17297 (N_17297,N_13895,N_14092);
and U17298 (N_17298,N_13497,N_15395);
nor U17299 (N_17299,N_12430,N_14606);
and U17300 (N_17300,N_12219,N_12641);
or U17301 (N_17301,N_12917,N_12990);
xnor U17302 (N_17302,N_12167,N_14996);
xnor U17303 (N_17303,N_14273,N_14704);
or U17304 (N_17304,N_14333,N_13221);
and U17305 (N_17305,N_13343,N_14998);
and U17306 (N_17306,N_12742,N_12268);
xor U17307 (N_17307,N_14340,N_14821);
and U17308 (N_17308,N_13712,N_13407);
xnor U17309 (N_17309,N_15324,N_13305);
xor U17310 (N_17310,N_14316,N_15730);
nand U17311 (N_17311,N_14689,N_15146);
xnor U17312 (N_17312,N_13979,N_12976);
and U17313 (N_17313,N_12867,N_13025);
nand U17314 (N_17314,N_14529,N_12527);
xnor U17315 (N_17315,N_13699,N_15820);
nor U17316 (N_17316,N_14425,N_12088);
nor U17317 (N_17317,N_13789,N_13111);
and U17318 (N_17318,N_14446,N_14833);
and U17319 (N_17319,N_15965,N_14818);
or U17320 (N_17320,N_14935,N_14952);
xnor U17321 (N_17321,N_12136,N_14803);
and U17322 (N_17322,N_12388,N_14303);
nor U17323 (N_17323,N_15738,N_13836);
or U17324 (N_17324,N_15208,N_15030);
or U17325 (N_17325,N_14782,N_15248);
xor U17326 (N_17326,N_14839,N_13369);
nand U17327 (N_17327,N_12407,N_15746);
or U17328 (N_17328,N_13612,N_15079);
nand U17329 (N_17329,N_14546,N_14794);
or U17330 (N_17330,N_12916,N_13057);
xor U17331 (N_17331,N_15063,N_12885);
and U17332 (N_17332,N_14072,N_13346);
nor U17333 (N_17333,N_14608,N_12391);
and U17334 (N_17334,N_12651,N_12953);
nor U17335 (N_17335,N_14713,N_12663);
xor U17336 (N_17336,N_12462,N_12902);
or U17337 (N_17337,N_13165,N_12370);
nand U17338 (N_17338,N_15266,N_14535);
nand U17339 (N_17339,N_15719,N_15387);
or U17340 (N_17340,N_13092,N_15598);
nor U17341 (N_17341,N_14846,N_15157);
nor U17342 (N_17342,N_12751,N_15297);
xor U17343 (N_17343,N_12653,N_14527);
nand U17344 (N_17344,N_14107,N_12965);
nor U17345 (N_17345,N_12723,N_12506);
xor U17346 (N_17346,N_13043,N_15723);
and U17347 (N_17347,N_13351,N_14168);
nor U17348 (N_17348,N_13587,N_15234);
nor U17349 (N_17349,N_14899,N_15631);
nand U17350 (N_17350,N_13068,N_12270);
and U17351 (N_17351,N_14321,N_12776);
xnor U17352 (N_17352,N_14681,N_15951);
and U17353 (N_17353,N_14898,N_15045);
nor U17354 (N_17354,N_13498,N_12745);
or U17355 (N_17355,N_14702,N_15181);
or U17356 (N_17356,N_15725,N_13446);
or U17357 (N_17357,N_12117,N_13838);
nand U17358 (N_17358,N_14445,N_14228);
xor U17359 (N_17359,N_12244,N_14109);
and U17360 (N_17360,N_14334,N_12273);
nand U17361 (N_17361,N_12346,N_15689);
xor U17362 (N_17362,N_12240,N_12825);
and U17363 (N_17363,N_12793,N_15341);
nor U17364 (N_17364,N_12504,N_12038);
nand U17365 (N_17365,N_15987,N_14738);
xor U17366 (N_17366,N_14789,N_12354);
xor U17367 (N_17367,N_13240,N_15231);
and U17368 (N_17368,N_13617,N_14852);
and U17369 (N_17369,N_15600,N_15227);
nor U17370 (N_17370,N_14011,N_15052);
or U17371 (N_17371,N_13077,N_13508);
and U17372 (N_17372,N_13611,N_14869);
or U17373 (N_17373,N_15304,N_15136);
nor U17374 (N_17374,N_15106,N_12345);
and U17375 (N_17375,N_15267,N_14515);
xor U17376 (N_17376,N_13117,N_12170);
nor U17377 (N_17377,N_15284,N_13952);
or U17378 (N_17378,N_12558,N_14139);
or U17379 (N_17379,N_14777,N_12465);
xor U17380 (N_17380,N_12950,N_15483);
nand U17381 (N_17381,N_13261,N_15132);
or U17382 (N_17382,N_12080,N_13176);
nand U17383 (N_17383,N_15158,N_14429);
nor U17384 (N_17384,N_15814,N_14169);
or U17385 (N_17385,N_14180,N_13759);
nor U17386 (N_17386,N_13646,N_14087);
xor U17387 (N_17387,N_12993,N_14836);
nand U17388 (N_17388,N_12763,N_14348);
nand U17389 (N_17389,N_15271,N_13865);
and U17390 (N_17390,N_13802,N_14653);
and U17391 (N_17391,N_15011,N_15552);
xor U17392 (N_17392,N_14857,N_14335);
or U17393 (N_17393,N_15151,N_14017);
or U17394 (N_17394,N_12526,N_15119);
nor U17395 (N_17395,N_13783,N_13566);
xnor U17396 (N_17396,N_15349,N_12856);
and U17397 (N_17397,N_14567,N_15278);
xnor U17398 (N_17398,N_13512,N_12078);
nand U17399 (N_17399,N_15452,N_13179);
nor U17400 (N_17400,N_13792,N_14555);
or U17401 (N_17401,N_12511,N_12160);
or U17402 (N_17402,N_14039,N_12773);
nand U17403 (N_17403,N_14301,N_13048);
nor U17404 (N_17404,N_14252,N_13127);
nor U17405 (N_17405,N_12429,N_13593);
xor U17406 (N_17406,N_12212,N_12350);
nor U17407 (N_17407,N_13800,N_15141);
or U17408 (N_17408,N_12453,N_12949);
nor U17409 (N_17409,N_15260,N_14342);
or U17410 (N_17410,N_13020,N_13500);
xor U17411 (N_17411,N_13102,N_13448);
or U17412 (N_17412,N_12180,N_13949);
nor U17413 (N_17413,N_13549,N_13045);
nand U17414 (N_17414,N_15508,N_15573);
or U17415 (N_17415,N_13557,N_14278);
xnor U17416 (N_17416,N_14263,N_12277);
nor U17417 (N_17417,N_13204,N_14049);
nor U17418 (N_17418,N_15423,N_12214);
and U17419 (N_17419,N_14415,N_13378);
and U17420 (N_17420,N_12441,N_14747);
nand U17421 (N_17421,N_12756,N_14856);
nor U17422 (N_17422,N_13270,N_15123);
xor U17423 (N_17423,N_13041,N_15529);
nand U17424 (N_17424,N_14913,N_15777);
or U17425 (N_17425,N_12470,N_12259);
or U17426 (N_17426,N_15328,N_13908);
or U17427 (N_17427,N_14999,N_12313);
and U17428 (N_17428,N_13624,N_12542);
xnor U17429 (N_17429,N_15245,N_15702);
or U17430 (N_17430,N_12923,N_13810);
nor U17431 (N_17431,N_13145,N_12048);
nand U17432 (N_17432,N_15427,N_12727);
nand U17433 (N_17433,N_15615,N_13664);
nand U17434 (N_17434,N_14432,N_14880);
nor U17435 (N_17435,N_15701,N_12006);
nor U17436 (N_17436,N_13247,N_14647);
or U17437 (N_17437,N_14940,N_15642);
nand U17438 (N_17438,N_15363,N_12144);
nand U17439 (N_17439,N_12501,N_12517);
xor U17440 (N_17440,N_14145,N_14788);
xor U17441 (N_17441,N_15630,N_12944);
xnor U17442 (N_17442,N_13093,N_13610);
and U17443 (N_17443,N_15592,N_12183);
and U17444 (N_17444,N_15784,N_14320);
xor U17445 (N_17445,N_12762,N_12014);
nor U17446 (N_17446,N_15771,N_12590);
nand U17447 (N_17447,N_14373,N_13484);
xor U17448 (N_17448,N_14401,N_13588);
and U17449 (N_17449,N_13105,N_15044);
or U17450 (N_17450,N_15384,N_14558);
nand U17451 (N_17451,N_13777,N_12411);
nor U17452 (N_17452,N_12893,N_14492);
nor U17453 (N_17453,N_15558,N_14959);
and U17454 (N_17454,N_12585,N_15849);
nor U17455 (N_17455,N_15655,N_15134);
and U17456 (N_17456,N_12417,N_13654);
nor U17457 (N_17457,N_12998,N_12674);
xnor U17458 (N_17458,N_12550,N_14126);
nor U17459 (N_17459,N_12654,N_14053);
or U17460 (N_17460,N_12942,N_13458);
nor U17461 (N_17461,N_12523,N_14625);
nand U17462 (N_17462,N_15915,N_12489);
nor U17463 (N_17463,N_14671,N_13406);
xor U17464 (N_17464,N_12806,N_14262);
nor U17465 (N_17465,N_12711,N_13130);
or U17466 (N_17466,N_15790,N_15506);
and U17467 (N_17467,N_15127,N_13091);
and U17468 (N_17468,N_15933,N_12184);
xnor U17469 (N_17469,N_13998,N_12873);
nor U17470 (N_17470,N_12707,N_15513);
nand U17471 (N_17471,N_13812,N_15708);
xor U17472 (N_17472,N_12830,N_14341);
and U17473 (N_17473,N_13213,N_13542);
or U17474 (N_17474,N_12633,N_14243);
and U17475 (N_17475,N_13680,N_13134);
and U17476 (N_17476,N_13686,N_15188);
or U17477 (N_17477,N_13173,N_12530);
or U17478 (N_17478,N_14816,N_13220);
and U17479 (N_17479,N_15912,N_12267);
or U17480 (N_17480,N_12819,N_12522);
and U17481 (N_17481,N_14135,N_15094);
xor U17482 (N_17482,N_12675,N_14059);
nor U17483 (N_17483,N_12280,N_14069);
nand U17484 (N_17484,N_13059,N_14932);
xor U17485 (N_17485,N_15716,N_14548);
or U17486 (N_17486,N_12775,N_12706);
and U17487 (N_17487,N_13972,N_13012);
nand U17488 (N_17488,N_15916,N_15931);
and U17489 (N_17489,N_15319,N_12507);
nand U17490 (N_17490,N_12202,N_15954);
or U17491 (N_17491,N_14554,N_13014);
nand U17492 (N_17492,N_12866,N_15817);
or U17493 (N_17493,N_15335,N_12584);
xor U17494 (N_17494,N_13985,N_14003);
and U17495 (N_17495,N_13141,N_12636);
and U17496 (N_17496,N_14422,N_12749);
xor U17497 (N_17497,N_15779,N_13317);
xor U17498 (N_17498,N_14047,N_15936);
nand U17499 (N_17499,N_15264,N_14475);
nand U17500 (N_17500,N_14731,N_13524);
nor U17501 (N_17501,N_12057,N_14230);
and U17502 (N_17502,N_12874,N_14338);
or U17503 (N_17503,N_14326,N_13750);
and U17504 (N_17504,N_12311,N_15731);
or U17505 (N_17505,N_12396,N_12992);
nor U17506 (N_17506,N_15818,N_14305);
and U17507 (N_17507,N_14812,N_14627);
nand U17508 (N_17508,N_15696,N_12936);
and U17509 (N_17509,N_14103,N_12314);
xor U17510 (N_17510,N_15289,N_14421);
xnor U17511 (N_17511,N_14190,N_14155);
nand U17512 (N_17512,N_12640,N_12514);
xor U17513 (N_17513,N_14486,N_13211);
and U17514 (N_17514,N_12089,N_14221);
nor U17515 (N_17515,N_13965,N_15952);
xor U17516 (N_17516,N_14951,N_12234);
xnor U17517 (N_17517,N_14651,N_14189);
xnor U17518 (N_17518,N_13975,N_12911);
or U17519 (N_17519,N_12162,N_12915);
and U17520 (N_17520,N_14851,N_15007);
nor U17521 (N_17521,N_14497,N_13007);
xor U17522 (N_17522,N_14683,N_15398);
or U17523 (N_17523,N_14691,N_15595);
or U17524 (N_17524,N_13565,N_15740);
or U17525 (N_17525,N_13714,N_12594);
and U17526 (N_17526,N_13534,N_12678);
nor U17527 (N_17527,N_15522,N_14574);
nand U17528 (N_17528,N_12335,N_12106);
and U17529 (N_17529,N_14455,N_15791);
nor U17530 (N_17530,N_13730,N_14509);
nor U17531 (N_17531,N_14902,N_15754);
and U17532 (N_17532,N_15676,N_13421);
nand U17533 (N_17533,N_15077,N_14430);
nand U17534 (N_17534,N_14499,N_13306);
xor U17535 (N_17535,N_13923,N_13442);
and U17536 (N_17536,N_12200,N_13203);
nor U17537 (N_17537,N_12357,N_15144);
and U17538 (N_17538,N_13010,N_12938);
xor U17539 (N_17539,N_15177,N_15909);
or U17540 (N_17540,N_15325,N_13902);
and U17541 (N_17541,N_13502,N_13334);
xnor U17542 (N_17542,N_13352,N_14692);
xor U17543 (N_17543,N_12444,N_12235);
or U17544 (N_17544,N_14405,N_14938);
and U17545 (N_17545,N_12174,N_14614);
or U17546 (N_17546,N_15883,N_13700);
nand U17547 (N_17547,N_13473,N_14586);
nor U17548 (N_17548,N_15006,N_12264);
nand U17549 (N_17549,N_13529,N_13821);
nand U17550 (N_17550,N_12668,N_14369);
xnor U17551 (N_17551,N_12389,N_14368);
xnor U17552 (N_17552,N_15988,N_14093);
and U17553 (N_17553,N_12442,N_15196);
nand U17554 (N_17554,N_14440,N_13339);
nand U17555 (N_17555,N_13431,N_15438);
and U17556 (N_17556,N_14379,N_14248);
and U17557 (N_17557,N_15269,N_12269);
nand U17558 (N_17558,N_14982,N_12084);
xnor U17559 (N_17559,N_14504,N_13906);
nor U17560 (N_17560,N_13968,N_15021);
nor U17561 (N_17561,N_12740,N_14876);
xor U17562 (N_17562,N_14167,N_15002);
and U17563 (N_17563,N_12630,N_14934);
or U17564 (N_17564,N_12824,N_13196);
and U17565 (N_17565,N_13118,N_14973);
nand U17566 (N_17566,N_13456,N_15525);
nand U17567 (N_17567,N_14867,N_12110);
nor U17568 (N_17568,N_13258,N_12843);
nor U17569 (N_17569,N_12095,N_15889);
xnor U17570 (N_17570,N_14602,N_15350);
and U17571 (N_17571,N_13948,N_13731);
xor U17572 (N_17572,N_12367,N_15469);
or U17573 (N_17573,N_13623,N_13791);
xnor U17574 (N_17574,N_13470,N_12920);
nor U17575 (N_17575,N_12817,N_13394);
nand U17576 (N_17576,N_13016,N_14388);
xnor U17577 (N_17577,N_12451,N_13641);
xnor U17578 (N_17578,N_15876,N_12236);
nor U17579 (N_17579,N_12980,N_15316);
nor U17580 (N_17580,N_14592,N_14319);
nor U17581 (N_17581,N_14166,N_12194);
and U17582 (N_17582,N_15942,N_12652);
xnor U17583 (N_17583,N_13896,N_15147);
nor U17584 (N_17584,N_14442,N_13970);
nand U17585 (N_17585,N_13311,N_12574);
nand U17586 (N_17586,N_15531,N_12384);
nor U17587 (N_17587,N_13585,N_14779);
or U17588 (N_17588,N_13029,N_13146);
nand U17589 (N_17589,N_13133,N_13409);
nand U17590 (N_17590,N_13649,N_14831);
and U17591 (N_17591,N_14352,N_13698);
xnor U17592 (N_17592,N_15073,N_13178);
or U17593 (N_17593,N_12816,N_15306);
and U17594 (N_17594,N_13107,N_15530);
and U17595 (N_17595,N_13953,N_13005);
or U17596 (N_17596,N_12454,N_13787);
and U17597 (N_17597,N_15979,N_13822);
xor U17598 (N_17598,N_13392,N_12249);
and U17599 (N_17599,N_14739,N_12794);
nand U17600 (N_17600,N_14783,N_13049);
xnor U17601 (N_17601,N_14892,N_13578);
xnor U17602 (N_17602,N_13569,N_15759);
xnor U17603 (N_17603,N_15867,N_15441);
nand U17604 (N_17604,N_15604,N_13754);
and U17605 (N_17605,N_13033,N_14302);
nand U17606 (N_17606,N_13927,N_12694);
nand U17607 (N_17607,N_12695,N_12292);
xnor U17608 (N_17608,N_14967,N_12764);
and U17609 (N_17609,N_13882,N_12094);
xor U17610 (N_17610,N_15113,N_13197);
and U17611 (N_17611,N_14621,N_15288);
xnor U17612 (N_17612,N_13372,N_15302);
or U17613 (N_17613,N_14051,N_14473);
nor U17614 (N_17614,N_15668,N_14659);
and U17615 (N_17615,N_12352,N_12845);
or U17616 (N_17616,N_14122,N_12243);
nand U17617 (N_17617,N_12964,N_12974);
and U17618 (N_17618,N_13194,N_15015);
or U17619 (N_17619,N_12955,N_15638);
and U17620 (N_17620,N_14603,N_14469);
and U17621 (N_17621,N_14837,N_15028);
and U17622 (N_17622,N_13064,N_13051);
or U17623 (N_17623,N_12432,N_15937);
or U17624 (N_17624,N_14097,N_14863);
xor U17625 (N_17625,N_15732,N_15229);
nand U17626 (N_17626,N_12604,N_13262);
nand U17627 (N_17627,N_14565,N_12689);
xnor U17628 (N_17628,N_15622,N_15617);
nor U17629 (N_17629,N_14754,N_12846);
and U17630 (N_17630,N_12145,N_13922);
and U17631 (N_17631,N_15310,N_12416);
nor U17632 (N_17632,N_13594,N_14584);
nor U17633 (N_17633,N_14694,N_15435);
xor U17634 (N_17634,N_13989,N_14843);
nand U17635 (N_17635,N_14547,N_12485);
nand U17636 (N_17636,N_14309,N_14750);
and U17637 (N_17637,N_13078,N_12323);
nand U17638 (N_17638,N_12158,N_14269);
xnor U17639 (N_17639,N_13937,N_13899);
xor U17640 (N_17640,N_14354,N_13114);
nand U17641 (N_17641,N_12177,N_12769);
xor U17642 (N_17642,N_15763,N_14085);
nand U17643 (N_17643,N_12889,N_14257);
nand U17644 (N_17644,N_13065,N_14082);
and U17645 (N_17645,N_15747,N_13886);
xor U17646 (N_17646,N_12809,N_13002);
xnor U17647 (N_17647,N_14984,N_13427);
or U17648 (N_17648,N_15978,N_12549);
or U17649 (N_17649,N_14451,N_13823);
xor U17650 (N_17650,N_12798,N_12924);
and U17651 (N_17651,N_12877,N_13857);
or U17652 (N_17652,N_12691,N_15766);
and U17653 (N_17653,N_15613,N_14431);
and U17654 (N_17654,N_12101,N_12023);
nor U17655 (N_17655,N_15043,N_14074);
and U17656 (N_17656,N_15085,N_12044);
nand U17657 (N_17657,N_14767,N_14063);
nand U17658 (N_17658,N_15417,N_13574);
nor U17659 (N_17659,N_14295,N_14491);
xnor U17660 (N_17660,N_15911,N_14792);
nand U17661 (N_17661,N_12289,N_13100);
nand U17662 (N_17662,N_14795,N_15724);
xnor U17663 (N_17663,N_12366,N_13609);
and U17664 (N_17664,N_14057,N_12903);
nand U17665 (N_17665,N_12785,N_14718);
xnor U17666 (N_17666,N_15905,N_14399);
and U17667 (N_17667,N_14588,N_13830);
nor U17668 (N_17668,N_12166,N_15130);
nand U17669 (N_17669,N_13253,N_15681);
nor U17670 (N_17670,N_15279,N_14136);
nand U17671 (N_17671,N_12488,N_12814);
nor U17672 (N_17672,N_12796,N_14636);
xor U17673 (N_17673,N_13824,N_14918);
or U17674 (N_17674,N_15705,N_13729);
and U17675 (N_17675,N_13846,N_13224);
nor U17676 (N_17676,N_15606,N_12985);
and U17677 (N_17677,N_15321,N_12205);
nand U17678 (N_17678,N_12484,N_15162);
or U17679 (N_17679,N_12051,N_15553);
xor U17680 (N_17680,N_12913,N_13891);
nand U17681 (N_17681,N_14536,N_13583);
xnor U17682 (N_17682,N_13149,N_13108);
nand U17683 (N_17683,N_15795,N_12521);
and U17684 (N_17684,N_14720,N_12518);
nor U17685 (N_17685,N_15715,N_14587);
and U17686 (N_17686,N_12190,N_13233);
or U17687 (N_17687,N_12066,N_14693);
xor U17688 (N_17688,N_13718,N_12562);
or U17689 (N_17689,N_14670,N_13330);
and U17690 (N_17690,N_14054,N_12863);
nand U17691 (N_17691,N_13630,N_15159);
and U17692 (N_17692,N_13600,N_12808);
xor U17693 (N_17693,N_15764,N_13322);
nand U17694 (N_17694,N_15470,N_14140);
and U17695 (N_17695,N_12896,N_13527);
nor U17696 (N_17696,N_12375,N_14142);
xnor U17697 (N_17697,N_15997,N_13185);
and U17698 (N_17698,N_12512,N_15017);
xnor U17699 (N_17699,N_14874,N_13606);
nand U17700 (N_17700,N_14387,N_15013);
xnor U17701 (N_17701,N_12409,N_14875);
xnor U17702 (N_17702,N_15769,N_14955);
nand U17703 (N_17703,N_15679,N_14406);
or U17704 (N_17704,N_15049,N_12931);
and U17705 (N_17705,N_13489,N_14171);
nor U17706 (N_17706,N_12619,N_13072);
nand U17707 (N_17707,N_15064,N_14613);
xnor U17708 (N_17708,N_14835,N_14813);
and U17709 (N_17709,N_13432,N_12623);
xor U17710 (N_17710,N_14590,N_12434);
and U17711 (N_17711,N_15446,N_15033);
xor U17712 (N_17712,N_13924,N_12586);
xnor U17713 (N_17713,N_13365,N_14495);
nor U17714 (N_17714,N_15362,N_13094);
nand U17715 (N_17715,N_12658,N_14520);
nand U17716 (N_17716,N_14187,N_12283);
xor U17717 (N_17717,N_12380,N_14942);
or U17718 (N_17718,N_13101,N_14407);
nand U17719 (N_17719,N_15892,N_12891);
xnor U17720 (N_17720,N_13710,N_14921);
nor U17721 (N_17721,N_12497,N_14115);
nor U17722 (N_17722,N_15845,N_13736);
nor U17723 (N_17723,N_14987,N_13088);
and U17724 (N_17724,N_14870,N_15517);
or U17725 (N_17725,N_13620,N_15107);
nand U17726 (N_17726,N_12363,N_13568);
xnor U17727 (N_17727,N_15967,N_15924);
nand U17728 (N_17728,N_12664,N_14106);
or U17729 (N_17729,N_14579,N_14256);
or U17730 (N_17730,N_15634,N_15437);
or U17731 (N_17731,N_13701,N_13581);
and U17732 (N_17732,N_13295,N_13665);
and U17733 (N_17733,N_12700,N_14827);
xor U17734 (N_17734,N_14939,N_13375);
or U17735 (N_17735,N_12102,N_15171);
xor U17736 (N_17736,N_12634,N_15808);
or U17737 (N_17737,N_12994,N_14088);
nor U17738 (N_17738,N_15986,N_13202);
nor U17739 (N_17739,N_15118,N_13263);
nor U17740 (N_17740,N_14886,N_13795);
or U17741 (N_17741,N_12042,N_12266);
xor U17742 (N_17742,N_13275,N_12736);
nand U17743 (N_17743,N_12951,N_14318);
nor U17744 (N_17744,N_14946,N_13042);
nand U17745 (N_17745,N_14709,N_13813);
nand U17746 (N_17746,N_15426,N_15287);
nor U17747 (N_17747,N_12858,N_12013);
and U17748 (N_17748,N_15082,N_15126);
or U17749 (N_17749,N_14895,N_13586);
nor U17750 (N_17750,N_12091,N_12324);
nor U17751 (N_17751,N_12376,N_14128);
and U17752 (N_17752,N_13851,N_15221);
xor U17753 (N_17753,N_12821,N_13991);
or U17754 (N_17754,N_13284,N_15743);
nor U17755 (N_17755,N_15415,N_14832);
or U17756 (N_17756,N_15907,N_14254);
xor U17757 (N_17757,N_13116,N_12135);
or U17758 (N_17758,N_15893,N_12098);
and U17759 (N_17759,N_13871,N_12643);
and U17760 (N_17760,N_13614,N_13168);
xnor U17761 (N_17761,N_13148,N_14860);
nor U17762 (N_17762,N_12612,N_12779);
xor U17763 (N_17763,N_13856,N_15861);
or U17764 (N_17764,N_13978,N_15314);
nand U17765 (N_17765,N_14027,N_13634);
xor U17766 (N_17766,N_12241,N_13067);
nand U17767 (N_17767,N_14759,N_12187);
or U17768 (N_17768,N_14114,N_12576);
or U17769 (N_17769,N_15841,N_12782);
and U17770 (N_17770,N_12097,N_12587);
and U17771 (N_17771,N_14277,N_13672);
and U17772 (N_17772,N_12588,N_12605);
and U17773 (N_17773,N_14229,N_14420);
or U17774 (N_17774,N_12130,N_13277);
xnor U17775 (N_17775,N_13832,N_14198);
or U17776 (N_17776,N_15480,N_13688);
nand U17777 (N_17777,N_13452,N_12331);
nand U17778 (N_17778,N_13877,N_13702);
nor U17779 (N_17779,N_13465,N_15455);
xnor U17780 (N_17780,N_15360,N_15022);
and U17781 (N_17781,N_12719,N_15072);
xnor U17782 (N_17782,N_15099,N_15842);
xnor U17783 (N_17783,N_15194,N_13397);
nor U17784 (N_17784,N_15075,N_12834);
and U17785 (N_17785,N_14662,N_12182);
nand U17786 (N_17786,N_13480,N_15466);
or U17787 (N_17787,N_12741,N_14963);
and U17788 (N_17788,N_15857,N_15663);
xnor U17789 (N_17789,N_12982,N_12925);
and U17790 (N_17790,N_14046,N_13401);
nor U17791 (N_17791,N_15768,N_14660);
nor U17792 (N_17792,N_13765,N_12797);
nor U17793 (N_17793,N_13996,N_14848);
nor U17794 (N_17794,N_15139,N_14989);
and U17795 (N_17795,N_14206,N_15129);
xnor U17796 (N_17796,N_13272,N_15424);
or U17797 (N_17797,N_12127,N_15562);
and U17798 (N_17798,N_14906,N_14994);
nor U17799 (N_17799,N_15524,N_12734);
nor U17800 (N_17800,N_14380,N_12406);
xor U17801 (N_17801,N_13279,N_14753);
nand U17802 (N_17802,N_15648,N_13195);
or U17803 (N_17803,N_13658,N_15031);
nor U17804 (N_17804,N_14274,N_12864);
xor U17805 (N_17805,N_14356,N_15580);
xnor U17806 (N_17806,N_14506,N_13433);
nand U17807 (N_17807,N_15488,N_15276);
and U17808 (N_17808,N_14376,N_13505);
nor U17809 (N_17809,N_14917,N_14236);
and U17810 (N_17810,N_13833,N_13690);
nor U17811 (N_17811,N_14582,N_15291);
xnor U17812 (N_17812,N_15966,N_13946);
or U17813 (N_17813,N_14067,N_13916);
nor U17814 (N_17814,N_14975,N_14583);
nor U17815 (N_17815,N_15068,N_15707);
or U17816 (N_17816,N_14201,N_12020);
xor U17817 (N_17817,N_12498,N_13356);
nor U17818 (N_17818,N_14001,N_13097);
or U17819 (N_17819,N_12546,N_15214);
xor U17820 (N_17820,N_12720,N_15187);
xor U17821 (N_17821,N_13110,N_12932);
or U17822 (N_17822,N_13670,N_14184);
nand U17823 (N_17823,N_14170,N_13264);
xor U17824 (N_17824,N_12635,N_14962);
nand U17825 (N_17825,N_13344,N_15644);
and U17826 (N_17826,N_14134,N_12206);
xor U17827 (N_17827,N_14929,N_15425);
nand U17828 (N_17828,N_13477,N_12455);
nor U17829 (N_17829,N_12056,N_15692);
nand U17830 (N_17830,N_12482,N_12743);
nand U17831 (N_17831,N_12351,N_15500);
xnor U17832 (N_17832,N_14698,N_14828);
nor U17833 (N_17833,N_15211,N_14634);
xnor U17834 (N_17834,N_12721,N_13098);
xnor U17835 (N_17835,N_12379,N_14578);
or U17836 (N_17836,N_15661,N_12656);
or U17837 (N_17837,N_12702,N_15491);
xor U17838 (N_17838,N_13954,N_15868);
nor U17839 (N_17839,N_14715,N_14741);
xor U17840 (N_17840,N_14517,N_15885);
and U17841 (N_17841,N_12616,N_13570);
nor U17842 (N_17842,N_12317,N_13276);
nand U17843 (N_17843,N_14378,N_13635);
xnor U17844 (N_17844,N_12309,N_12872);
and U17845 (N_17845,N_13760,N_14058);
nor U17846 (N_17846,N_13547,N_12112);
nor U17847 (N_17847,N_12404,N_15509);
nand U17848 (N_17848,N_12789,N_12890);
nand U17849 (N_17849,N_13642,N_15653);
nor U17850 (N_17850,N_12910,N_12347);
nand U17851 (N_17851,N_14395,N_12973);
nor U17852 (N_17852,N_12801,N_12520);
and U17853 (N_17853,N_12031,N_12995);
nor U17854 (N_17854,N_14550,N_14353);
nor U17855 (N_17855,N_14729,N_14040);
or U17856 (N_17856,N_15443,N_13615);
or U17857 (N_17857,N_13128,N_14214);
or U17858 (N_17858,N_13987,N_14151);
nand U17859 (N_17859,N_13199,N_12413);
xor U17860 (N_17860,N_14329,N_14493);
and U17861 (N_17861,N_12831,N_13292);
nand U17862 (N_17862,N_15343,N_12374);
nor U17863 (N_17863,N_15666,N_15871);
or U17864 (N_17864,N_13913,N_13132);
nor U17865 (N_17865,N_14474,N_12838);
or U17866 (N_17866,N_14029,N_14893);
or U17867 (N_17867,N_12203,N_14144);
nand U17868 (N_17868,N_14503,N_12645);
xor U17869 (N_17869,N_13819,N_15736);
nand U17870 (N_17870,N_13066,N_12772);
xor U17871 (N_17871,N_13183,N_13390);
nand U17872 (N_17872,N_13237,N_12099);
nor U17873 (N_17873,N_15168,N_14730);
nor U17874 (N_17874,N_15678,N_12746);
nand U17875 (N_17875,N_13803,N_14541);
nor U17876 (N_17876,N_13103,N_15247);
xor U17877 (N_17877,N_13945,N_15946);
nor U17878 (N_17878,N_15133,N_15397);
nand U17879 (N_17879,N_14501,N_14686);
nand U17880 (N_17880,N_15241,N_12393);
xor U17881 (N_17881,N_12631,N_12002);
nand U17882 (N_17882,N_12041,N_13885);
nor U17883 (N_17883,N_14211,N_13873);
xor U17884 (N_17884,N_12946,N_12139);
and U17885 (N_17885,N_14755,N_15414);
and U17886 (N_17886,N_13709,N_13398);
and U17887 (N_17887,N_14125,N_15614);
xnor U17888 (N_17888,N_13758,N_13844);
or U17889 (N_17889,N_15854,N_15593);
or U17890 (N_17890,N_13414,N_12344);
nor U17891 (N_17891,N_12717,N_14661);
or U17892 (N_17892,N_14238,N_14928);
xnor U17893 (N_17893,N_15463,N_15555);
and U17894 (N_17894,N_13274,N_14530);
or U17895 (N_17895,N_14339,N_12073);
and U17896 (N_17896,N_14868,N_15439);
xnor U17897 (N_17897,N_12107,N_14673);
nor U17898 (N_17898,N_15256,N_15217);
or U17899 (N_17899,N_13302,N_14290);
nand U17900 (N_17900,N_15244,N_13082);
nand U17901 (N_17901,N_13767,N_14250);
nor U17902 (N_17902,N_15010,N_14268);
nand U17903 (N_17903,N_12983,N_12302);
or U17904 (N_17904,N_15070,N_12034);
or U17905 (N_17905,N_14969,N_13744);
and U17906 (N_17906,N_12253,N_13715);
nand U17907 (N_17907,N_15843,N_14359);
xnor U17908 (N_17908,N_12957,N_12246);
or U17909 (N_17909,N_13368,N_13874);
nand U17910 (N_17910,N_12547,N_15547);
and U17911 (N_17911,N_14397,N_13947);
nor U17912 (N_17912,N_12822,N_13967);
nor U17913 (N_17913,N_12120,N_12281);
nor U17914 (N_17914,N_12338,N_14385);
or U17915 (N_17915,N_15048,N_12103);
or U17916 (N_17916,N_13691,N_15203);
and U17917 (N_17917,N_15947,N_12085);
xor U17918 (N_17918,N_15388,N_13546);
or U17919 (N_17919,N_14162,N_14412);
or U17920 (N_17920,N_13647,N_12524);
nand U17921 (N_17921,N_14396,N_15773);
nand U17922 (N_17922,N_12329,N_14571);
nand U17923 (N_17923,N_12257,N_12718);
nand U17924 (N_17924,N_15686,N_12032);
xor U17925 (N_17925,N_13567,N_15389);
or U17926 (N_17926,N_13532,N_14298);
nand U17927 (N_17927,N_15956,N_15053);
or U17928 (N_17928,N_15810,N_15632);
or U17929 (N_17929,N_14786,N_15058);
nor U17930 (N_17930,N_14419,N_13001);
or U17931 (N_17931,N_12493,N_15787);
or U17932 (N_17932,N_15074,N_13602);
or U17933 (N_17933,N_14988,N_15514);
nand U17934 (N_17934,N_12123,N_14986);
xor U17935 (N_17935,N_15518,N_13561);
or U17936 (N_17936,N_15926,N_13912);
or U17937 (N_17937,N_13073,N_14306);
and U17938 (N_17938,N_14199,N_15377);
or U17939 (N_17939,N_15412,N_12326);
xor U17940 (N_17940,N_15178,N_14927);
and U17941 (N_17941,N_14696,N_12781);
nor U17942 (N_17942,N_12927,N_13395);
nand U17943 (N_17943,N_15367,N_12364);
or U17944 (N_17944,N_13559,N_12747);
xor U17945 (N_17945,N_15969,N_14102);
nand U17946 (N_17946,N_14785,N_13601);
and U17947 (N_17947,N_14215,N_12841);
or U17948 (N_17948,N_12061,N_15218);
and U17949 (N_17949,N_13739,N_13633);
or U17950 (N_17950,N_15459,N_13260);
xor U17951 (N_17951,N_12551,N_12365);
nand U17952 (N_17952,N_12175,N_13062);
nor U17953 (N_17953,N_14685,N_13180);
and U17954 (N_17954,N_14819,N_15559);
xor U17955 (N_17955,N_15400,N_13308);
xor U17956 (N_17956,N_12812,N_14787);
xnor U17957 (N_17957,N_14576,N_12378);
nor U17958 (N_17958,N_13129,N_15311);
and U17959 (N_17959,N_15332,N_12894);
or U17960 (N_17960,N_14805,N_12456);
nor U17961 (N_17961,N_12571,N_12515);
nand U17962 (N_17962,N_12290,N_14533);
nand U17963 (N_17963,N_14531,N_14377);
nand U17964 (N_17964,N_12933,N_13693);
or U17965 (N_17965,N_12467,N_15246);
nor U17966 (N_17966,N_14344,N_15939);
xor U17967 (N_17967,N_12140,N_14679);
nand U17968 (N_17968,N_14240,N_12701);
nand U17969 (N_17969,N_13893,N_15381);
nand U17970 (N_17970,N_13509,N_14098);
xnor U17971 (N_17971,N_12328,N_12569);
xor U17972 (N_17972,N_13868,N_12256);
nor U17973 (N_17973,N_14195,N_13050);
or U17974 (N_17974,N_13656,N_15720);
xor U17975 (N_17975,N_14840,N_13550);
nor U17976 (N_17976,N_12030,N_12457);
and U17977 (N_17977,N_15197,N_14033);
and U17978 (N_17978,N_12035,N_15238);
xor U17979 (N_17979,N_14450,N_15356);
and U17980 (N_17980,N_12402,N_14675);
xnor U17981 (N_17981,N_12221,N_15792);
nor U17982 (N_17982,N_12884,N_12227);
nand U17983 (N_17983,N_15968,N_15863);
xor U17984 (N_17984,N_14178,N_15651);
nor U17985 (N_17985,N_15507,N_13191);
or U17986 (N_17986,N_12047,N_14207);
or U17987 (N_17987,N_13402,N_15180);
or U17988 (N_17988,N_12477,N_15596);
nand U17989 (N_17989,N_15299,N_14620);
nand U17990 (N_17990,N_13287,N_15095);
nand U17991 (N_17991,N_13782,N_15536);
or U17992 (N_17992,N_13994,N_14071);
nand U17993 (N_17993,N_12420,N_15900);
nand U17994 (N_17994,N_13919,N_15974);
or U17995 (N_17995,N_12033,N_15471);
nor U17996 (N_17996,N_14331,N_14622);
xnor U17997 (N_17997,N_15832,N_14456);
nor U17998 (N_17998,N_14914,N_15844);
or U17999 (N_17999,N_15914,N_14632);
or U18000 (N_18000,N_14228,N_15656);
and U18001 (N_18001,N_15171,N_14952);
xor U18002 (N_18002,N_14652,N_15777);
nand U18003 (N_18003,N_13226,N_14967);
xnor U18004 (N_18004,N_14034,N_12457);
or U18005 (N_18005,N_12410,N_13056);
or U18006 (N_18006,N_13105,N_15219);
nand U18007 (N_18007,N_13258,N_14980);
or U18008 (N_18008,N_13737,N_13532);
nand U18009 (N_18009,N_13774,N_14329);
nand U18010 (N_18010,N_12152,N_13115);
nor U18011 (N_18011,N_13071,N_12764);
or U18012 (N_18012,N_14613,N_15902);
or U18013 (N_18013,N_15325,N_14748);
nor U18014 (N_18014,N_14848,N_12332);
or U18015 (N_18015,N_14845,N_14116);
xor U18016 (N_18016,N_15815,N_15402);
or U18017 (N_18017,N_13285,N_15598);
and U18018 (N_18018,N_14581,N_13239);
nor U18019 (N_18019,N_15586,N_13590);
nor U18020 (N_18020,N_14469,N_14026);
or U18021 (N_18021,N_15929,N_13098);
nor U18022 (N_18022,N_15385,N_13338);
nand U18023 (N_18023,N_15750,N_13697);
nor U18024 (N_18024,N_13366,N_13191);
xnor U18025 (N_18025,N_13058,N_12896);
or U18026 (N_18026,N_13193,N_14774);
or U18027 (N_18027,N_14823,N_13766);
nor U18028 (N_18028,N_13871,N_14758);
nand U18029 (N_18029,N_13269,N_12034);
nand U18030 (N_18030,N_15531,N_14292);
nand U18031 (N_18031,N_14019,N_13636);
nand U18032 (N_18032,N_12062,N_12072);
xor U18033 (N_18033,N_15697,N_12638);
nor U18034 (N_18034,N_15424,N_12862);
or U18035 (N_18035,N_13077,N_13012);
and U18036 (N_18036,N_14545,N_13919);
xor U18037 (N_18037,N_13459,N_15126);
xor U18038 (N_18038,N_15428,N_15550);
xor U18039 (N_18039,N_12179,N_12444);
xnor U18040 (N_18040,N_12510,N_12213);
nor U18041 (N_18041,N_14820,N_15595);
and U18042 (N_18042,N_13854,N_12059);
nand U18043 (N_18043,N_12685,N_14086);
nand U18044 (N_18044,N_12275,N_15190);
nor U18045 (N_18045,N_13402,N_14174);
nand U18046 (N_18046,N_14555,N_15700);
and U18047 (N_18047,N_12634,N_12456);
nand U18048 (N_18048,N_13908,N_14551);
or U18049 (N_18049,N_14258,N_13523);
or U18050 (N_18050,N_13528,N_15503);
or U18051 (N_18051,N_12407,N_15048);
and U18052 (N_18052,N_12893,N_15344);
or U18053 (N_18053,N_12359,N_14251);
and U18054 (N_18054,N_15524,N_13103);
and U18055 (N_18055,N_15766,N_15786);
nor U18056 (N_18056,N_13659,N_13329);
nor U18057 (N_18057,N_15028,N_13496);
xnor U18058 (N_18058,N_12798,N_14337);
and U18059 (N_18059,N_15096,N_13317);
or U18060 (N_18060,N_12085,N_13932);
or U18061 (N_18061,N_14647,N_12548);
nand U18062 (N_18062,N_14837,N_13802);
nor U18063 (N_18063,N_15316,N_14617);
nor U18064 (N_18064,N_12399,N_14195);
nand U18065 (N_18065,N_14724,N_13599);
and U18066 (N_18066,N_13133,N_12527);
nand U18067 (N_18067,N_13593,N_15038);
nand U18068 (N_18068,N_14406,N_12429);
nand U18069 (N_18069,N_13078,N_15855);
nand U18070 (N_18070,N_14161,N_12917);
xor U18071 (N_18071,N_14885,N_15004);
xnor U18072 (N_18072,N_14367,N_12381);
nor U18073 (N_18073,N_12453,N_14881);
or U18074 (N_18074,N_12094,N_15221);
nor U18075 (N_18075,N_15584,N_12036);
and U18076 (N_18076,N_13506,N_14185);
and U18077 (N_18077,N_14859,N_14159);
nand U18078 (N_18078,N_14508,N_15036);
or U18079 (N_18079,N_13852,N_13865);
nand U18080 (N_18080,N_15023,N_15701);
or U18081 (N_18081,N_12721,N_13680);
and U18082 (N_18082,N_15727,N_13191);
nand U18083 (N_18083,N_13810,N_12197);
nand U18084 (N_18084,N_13019,N_15554);
or U18085 (N_18085,N_15869,N_14586);
nor U18086 (N_18086,N_12809,N_12065);
or U18087 (N_18087,N_15495,N_14685);
xnor U18088 (N_18088,N_12862,N_12154);
or U18089 (N_18089,N_13051,N_13445);
or U18090 (N_18090,N_14027,N_12018);
nor U18091 (N_18091,N_13816,N_14883);
and U18092 (N_18092,N_15387,N_15704);
xnor U18093 (N_18093,N_15724,N_14628);
xnor U18094 (N_18094,N_13902,N_14638);
and U18095 (N_18095,N_15676,N_15254);
or U18096 (N_18096,N_12701,N_15941);
or U18097 (N_18097,N_13482,N_13380);
or U18098 (N_18098,N_14471,N_15542);
or U18099 (N_18099,N_13337,N_12900);
xnor U18100 (N_18100,N_12611,N_15944);
and U18101 (N_18101,N_15165,N_12114);
and U18102 (N_18102,N_13933,N_14256);
or U18103 (N_18103,N_14990,N_12405);
or U18104 (N_18104,N_12858,N_13879);
xnor U18105 (N_18105,N_13239,N_15799);
nand U18106 (N_18106,N_12960,N_12346);
nand U18107 (N_18107,N_13012,N_13254);
nor U18108 (N_18108,N_15278,N_13777);
nand U18109 (N_18109,N_13224,N_15401);
nor U18110 (N_18110,N_15596,N_15833);
or U18111 (N_18111,N_15011,N_13719);
nor U18112 (N_18112,N_15175,N_12009);
and U18113 (N_18113,N_13362,N_15951);
and U18114 (N_18114,N_12642,N_12717);
or U18115 (N_18115,N_15989,N_13080);
or U18116 (N_18116,N_14603,N_15154);
xor U18117 (N_18117,N_13489,N_12436);
and U18118 (N_18118,N_15496,N_15321);
and U18119 (N_18119,N_13163,N_14246);
and U18120 (N_18120,N_13080,N_15260);
and U18121 (N_18121,N_12608,N_13038);
or U18122 (N_18122,N_13766,N_14536);
and U18123 (N_18123,N_15851,N_13625);
nand U18124 (N_18124,N_12331,N_14008);
nor U18125 (N_18125,N_14981,N_13626);
nor U18126 (N_18126,N_12289,N_14624);
xnor U18127 (N_18127,N_12343,N_14976);
and U18128 (N_18128,N_12059,N_12864);
nor U18129 (N_18129,N_12921,N_12664);
nand U18130 (N_18130,N_12481,N_15496);
nand U18131 (N_18131,N_15064,N_13808);
nor U18132 (N_18132,N_15425,N_15624);
nor U18133 (N_18133,N_14802,N_12428);
nor U18134 (N_18134,N_12494,N_13235);
nand U18135 (N_18135,N_13541,N_14327);
and U18136 (N_18136,N_12353,N_14056);
xor U18137 (N_18137,N_13724,N_12504);
nor U18138 (N_18138,N_15323,N_12180);
and U18139 (N_18139,N_13889,N_15905);
nand U18140 (N_18140,N_13983,N_12321);
nand U18141 (N_18141,N_13096,N_12271);
xnor U18142 (N_18142,N_15107,N_15587);
or U18143 (N_18143,N_13177,N_12556);
nor U18144 (N_18144,N_14932,N_14256);
and U18145 (N_18145,N_12947,N_14817);
and U18146 (N_18146,N_14341,N_12686);
nand U18147 (N_18147,N_15358,N_15429);
nor U18148 (N_18148,N_15968,N_13378);
nand U18149 (N_18149,N_12473,N_14055);
or U18150 (N_18150,N_15468,N_14870);
and U18151 (N_18151,N_12033,N_14542);
or U18152 (N_18152,N_15338,N_14494);
and U18153 (N_18153,N_15056,N_12894);
and U18154 (N_18154,N_13430,N_15609);
or U18155 (N_18155,N_13712,N_15506);
nor U18156 (N_18156,N_13899,N_15352);
xor U18157 (N_18157,N_15350,N_14518);
and U18158 (N_18158,N_14108,N_12583);
xnor U18159 (N_18159,N_13028,N_15260);
xor U18160 (N_18160,N_13173,N_15377);
and U18161 (N_18161,N_14591,N_14464);
or U18162 (N_18162,N_14883,N_13894);
nor U18163 (N_18163,N_13666,N_14365);
nor U18164 (N_18164,N_15297,N_14450);
nor U18165 (N_18165,N_12754,N_12735);
and U18166 (N_18166,N_13636,N_15377);
xnor U18167 (N_18167,N_12811,N_14448);
xnor U18168 (N_18168,N_14773,N_12404);
nand U18169 (N_18169,N_13966,N_12253);
nor U18170 (N_18170,N_15799,N_15649);
or U18171 (N_18171,N_12407,N_14143);
nor U18172 (N_18172,N_15639,N_15630);
or U18173 (N_18173,N_14047,N_13821);
nor U18174 (N_18174,N_12610,N_14459);
nor U18175 (N_18175,N_13728,N_12656);
xnor U18176 (N_18176,N_15845,N_14552);
nor U18177 (N_18177,N_15085,N_12261);
and U18178 (N_18178,N_15643,N_13686);
nor U18179 (N_18179,N_15507,N_14744);
nand U18180 (N_18180,N_14334,N_14252);
nor U18181 (N_18181,N_14509,N_14188);
and U18182 (N_18182,N_14335,N_15443);
or U18183 (N_18183,N_12310,N_13522);
nand U18184 (N_18184,N_12571,N_13590);
xor U18185 (N_18185,N_12833,N_12211);
nor U18186 (N_18186,N_15538,N_15211);
or U18187 (N_18187,N_12228,N_13884);
or U18188 (N_18188,N_15194,N_14465);
and U18189 (N_18189,N_15715,N_12406);
nor U18190 (N_18190,N_15433,N_15662);
and U18191 (N_18191,N_13343,N_12482);
or U18192 (N_18192,N_13795,N_15634);
xnor U18193 (N_18193,N_15186,N_15116);
or U18194 (N_18194,N_15976,N_14951);
nor U18195 (N_18195,N_12704,N_12730);
and U18196 (N_18196,N_15641,N_12149);
nor U18197 (N_18197,N_15359,N_14431);
xor U18198 (N_18198,N_13364,N_15793);
xor U18199 (N_18199,N_12928,N_15120);
xor U18200 (N_18200,N_15541,N_12472);
and U18201 (N_18201,N_12857,N_12572);
and U18202 (N_18202,N_15810,N_13979);
and U18203 (N_18203,N_15675,N_13539);
nor U18204 (N_18204,N_15375,N_15547);
nor U18205 (N_18205,N_12814,N_13785);
and U18206 (N_18206,N_13398,N_12847);
nand U18207 (N_18207,N_12764,N_12241);
nor U18208 (N_18208,N_15477,N_12100);
nor U18209 (N_18209,N_15785,N_12397);
or U18210 (N_18210,N_13019,N_13970);
and U18211 (N_18211,N_13178,N_15581);
and U18212 (N_18212,N_13186,N_12105);
and U18213 (N_18213,N_15614,N_12704);
nor U18214 (N_18214,N_13543,N_13092);
nor U18215 (N_18215,N_13111,N_13662);
nor U18216 (N_18216,N_15351,N_13471);
xnor U18217 (N_18217,N_13196,N_12911);
nor U18218 (N_18218,N_12030,N_15673);
nor U18219 (N_18219,N_12545,N_13723);
and U18220 (N_18220,N_14407,N_12558);
xnor U18221 (N_18221,N_13212,N_14741);
and U18222 (N_18222,N_15695,N_12258);
nand U18223 (N_18223,N_12615,N_13558);
xor U18224 (N_18224,N_12166,N_13270);
xnor U18225 (N_18225,N_13110,N_13321);
and U18226 (N_18226,N_13561,N_12454);
nand U18227 (N_18227,N_13332,N_15036);
nor U18228 (N_18228,N_13995,N_12556);
nor U18229 (N_18229,N_14176,N_12830);
or U18230 (N_18230,N_15873,N_12871);
nor U18231 (N_18231,N_14459,N_12664);
nand U18232 (N_18232,N_13051,N_12642);
xor U18233 (N_18233,N_14120,N_14778);
nor U18234 (N_18234,N_15612,N_13663);
or U18235 (N_18235,N_15823,N_13128);
nor U18236 (N_18236,N_14386,N_12729);
and U18237 (N_18237,N_12447,N_12651);
or U18238 (N_18238,N_15324,N_12561);
and U18239 (N_18239,N_13492,N_12806);
and U18240 (N_18240,N_15421,N_14131);
nor U18241 (N_18241,N_13792,N_15296);
and U18242 (N_18242,N_15711,N_14429);
and U18243 (N_18243,N_15842,N_13254);
xor U18244 (N_18244,N_13644,N_14320);
or U18245 (N_18245,N_14460,N_14834);
nand U18246 (N_18246,N_15916,N_13767);
nor U18247 (N_18247,N_13706,N_12942);
or U18248 (N_18248,N_12913,N_14314);
and U18249 (N_18249,N_15976,N_15982);
and U18250 (N_18250,N_14905,N_13729);
nand U18251 (N_18251,N_13971,N_14033);
nand U18252 (N_18252,N_14116,N_14554);
xor U18253 (N_18253,N_12275,N_14486);
and U18254 (N_18254,N_13202,N_14983);
or U18255 (N_18255,N_13320,N_13774);
xnor U18256 (N_18256,N_14183,N_13644);
or U18257 (N_18257,N_13569,N_15058);
and U18258 (N_18258,N_13607,N_14283);
xor U18259 (N_18259,N_12807,N_13739);
and U18260 (N_18260,N_14292,N_14742);
nand U18261 (N_18261,N_15165,N_13961);
xor U18262 (N_18262,N_13503,N_12926);
nand U18263 (N_18263,N_15883,N_14596);
and U18264 (N_18264,N_13626,N_13547);
nor U18265 (N_18265,N_13616,N_14346);
nor U18266 (N_18266,N_13313,N_12201);
and U18267 (N_18267,N_12950,N_14735);
and U18268 (N_18268,N_15736,N_15515);
or U18269 (N_18269,N_14310,N_14690);
xnor U18270 (N_18270,N_12214,N_12055);
or U18271 (N_18271,N_13704,N_14676);
nand U18272 (N_18272,N_14655,N_14457);
or U18273 (N_18273,N_13752,N_13563);
nor U18274 (N_18274,N_12823,N_12347);
or U18275 (N_18275,N_14775,N_12266);
nand U18276 (N_18276,N_12242,N_12523);
nor U18277 (N_18277,N_13100,N_15584);
nand U18278 (N_18278,N_14599,N_15306);
xnor U18279 (N_18279,N_14237,N_14217);
or U18280 (N_18280,N_12582,N_15390);
xnor U18281 (N_18281,N_14412,N_15117);
nor U18282 (N_18282,N_14098,N_13862);
or U18283 (N_18283,N_12314,N_13470);
or U18284 (N_18284,N_12239,N_12929);
and U18285 (N_18285,N_13426,N_15964);
and U18286 (N_18286,N_13425,N_12702);
xnor U18287 (N_18287,N_13543,N_15766);
or U18288 (N_18288,N_15336,N_15052);
xnor U18289 (N_18289,N_12835,N_15108);
or U18290 (N_18290,N_13001,N_13807);
and U18291 (N_18291,N_12677,N_15320);
nor U18292 (N_18292,N_12986,N_12837);
or U18293 (N_18293,N_14426,N_12417);
nand U18294 (N_18294,N_13252,N_14694);
xnor U18295 (N_18295,N_15870,N_12821);
xnor U18296 (N_18296,N_13933,N_15844);
or U18297 (N_18297,N_14283,N_13152);
xnor U18298 (N_18298,N_15047,N_12787);
xnor U18299 (N_18299,N_15371,N_15798);
or U18300 (N_18300,N_14249,N_15236);
xnor U18301 (N_18301,N_12412,N_13861);
and U18302 (N_18302,N_15365,N_13650);
nor U18303 (N_18303,N_12616,N_13394);
and U18304 (N_18304,N_13663,N_14324);
or U18305 (N_18305,N_12530,N_15570);
nand U18306 (N_18306,N_15229,N_14534);
xnor U18307 (N_18307,N_13497,N_14406);
or U18308 (N_18308,N_15182,N_13086);
and U18309 (N_18309,N_14601,N_14286);
nor U18310 (N_18310,N_13984,N_12322);
or U18311 (N_18311,N_15208,N_15882);
xor U18312 (N_18312,N_13827,N_13790);
nor U18313 (N_18313,N_15669,N_15329);
and U18314 (N_18314,N_14041,N_12119);
nand U18315 (N_18315,N_14045,N_14742);
or U18316 (N_18316,N_14688,N_14355);
nand U18317 (N_18317,N_13326,N_14475);
nand U18318 (N_18318,N_15225,N_15728);
nor U18319 (N_18319,N_15654,N_13410);
or U18320 (N_18320,N_14946,N_13741);
and U18321 (N_18321,N_15208,N_14561);
nand U18322 (N_18322,N_12076,N_15514);
xnor U18323 (N_18323,N_14943,N_14814);
nor U18324 (N_18324,N_14871,N_15661);
and U18325 (N_18325,N_14964,N_13684);
and U18326 (N_18326,N_12208,N_15897);
xnor U18327 (N_18327,N_14850,N_15971);
xnor U18328 (N_18328,N_14623,N_15097);
and U18329 (N_18329,N_13807,N_12235);
and U18330 (N_18330,N_13046,N_14221);
or U18331 (N_18331,N_13875,N_15678);
or U18332 (N_18332,N_12865,N_12937);
and U18333 (N_18333,N_15673,N_14629);
and U18334 (N_18334,N_14934,N_15590);
or U18335 (N_18335,N_12391,N_13167);
and U18336 (N_18336,N_12403,N_12515);
nand U18337 (N_18337,N_15239,N_12085);
and U18338 (N_18338,N_13742,N_12064);
xnor U18339 (N_18339,N_14271,N_13866);
nor U18340 (N_18340,N_15857,N_13696);
or U18341 (N_18341,N_12189,N_12554);
xnor U18342 (N_18342,N_12652,N_15041);
xor U18343 (N_18343,N_13257,N_14909);
nand U18344 (N_18344,N_15528,N_13628);
or U18345 (N_18345,N_12826,N_14224);
nand U18346 (N_18346,N_14390,N_13192);
nor U18347 (N_18347,N_15140,N_12822);
nor U18348 (N_18348,N_12934,N_15434);
nor U18349 (N_18349,N_12140,N_14966);
xor U18350 (N_18350,N_12389,N_15904);
xnor U18351 (N_18351,N_15681,N_15908);
nand U18352 (N_18352,N_14555,N_15141);
nor U18353 (N_18353,N_12334,N_12614);
nand U18354 (N_18354,N_14195,N_14898);
and U18355 (N_18355,N_14061,N_14947);
nor U18356 (N_18356,N_12006,N_15537);
nor U18357 (N_18357,N_12935,N_15297);
and U18358 (N_18358,N_13994,N_12905);
xnor U18359 (N_18359,N_14169,N_15975);
nand U18360 (N_18360,N_14041,N_14143);
nand U18361 (N_18361,N_14000,N_12516);
nand U18362 (N_18362,N_14314,N_15572);
nand U18363 (N_18363,N_13393,N_14197);
nor U18364 (N_18364,N_12041,N_13031);
nand U18365 (N_18365,N_14415,N_12564);
nor U18366 (N_18366,N_14861,N_14645);
xor U18367 (N_18367,N_12626,N_14335);
or U18368 (N_18368,N_14515,N_15720);
xor U18369 (N_18369,N_13463,N_14113);
or U18370 (N_18370,N_14924,N_14466);
or U18371 (N_18371,N_12056,N_15526);
or U18372 (N_18372,N_14941,N_12838);
nand U18373 (N_18373,N_12123,N_13644);
or U18374 (N_18374,N_14502,N_13157);
nor U18375 (N_18375,N_15934,N_14948);
and U18376 (N_18376,N_12987,N_13151);
or U18377 (N_18377,N_15874,N_12890);
and U18378 (N_18378,N_14684,N_14747);
nor U18379 (N_18379,N_15527,N_15492);
and U18380 (N_18380,N_14473,N_15126);
nand U18381 (N_18381,N_12371,N_13371);
or U18382 (N_18382,N_13766,N_13858);
or U18383 (N_18383,N_14733,N_14337);
or U18384 (N_18384,N_15899,N_14199);
nor U18385 (N_18385,N_12470,N_14890);
nand U18386 (N_18386,N_14610,N_13261);
nor U18387 (N_18387,N_14029,N_13531);
nand U18388 (N_18388,N_13769,N_14531);
nor U18389 (N_18389,N_14342,N_15582);
and U18390 (N_18390,N_14513,N_14046);
xnor U18391 (N_18391,N_14005,N_12251);
nand U18392 (N_18392,N_15893,N_14770);
or U18393 (N_18393,N_15787,N_13769);
xnor U18394 (N_18394,N_15389,N_14437);
and U18395 (N_18395,N_12661,N_13194);
nor U18396 (N_18396,N_12595,N_13733);
nand U18397 (N_18397,N_14685,N_14232);
nor U18398 (N_18398,N_14177,N_12951);
and U18399 (N_18399,N_15294,N_15284);
nor U18400 (N_18400,N_14876,N_14974);
nor U18401 (N_18401,N_14323,N_14596);
nor U18402 (N_18402,N_14953,N_12938);
and U18403 (N_18403,N_15316,N_14971);
or U18404 (N_18404,N_14788,N_12686);
xor U18405 (N_18405,N_13335,N_12250);
or U18406 (N_18406,N_14306,N_13996);
nor U18407 (N_18407,N_14508,N_12398);
xnor U18408 (N_18408,N_13684,N_12437);
or U18409 (N_18409,N_13778,N_12600);
and U18410 (N_18410,N_13301,N_13337);
nand U18411 (N_18411,N_13140,N_13248);
or U18412 (N_18412,N_14292,N_13739);
or U18413 (N_18413,N_13726,N_12605);
and U18414 (N_18414,N_14195,N_13826);
nand U18415 (N_18415,N_15592,N_14435);
xor U18416 (N_18416,N_15585,N_14447);
and U18417 (N_18417,N_15116,N_12616);
nor U18418 (N_18418,N_13582,N_15609);
and U18419 (N_18419,N_12704,N_15809);
or U18420 (N_18420,N_15708,N_12129);
and U18421 (N_18421,N_15376,N_14052);
nand U18422 (N_18422,N_15203,N_15975);
nand U18423 (N_18423,N_15231,N_13860);
xnor U18424 (N_18424,N_12613,N_15720);
and U18425 (N_18425,N_12873,N_13299);
xor U18426 (N_18426,N_13696,N_12544);
and U18427 (N_18427,N_12190,N_13615);
xor U18428 (N_18428,N_13701,N_13772);
nor U18429 (N_18429,N_15133,N_14113);
nor U18430 (N_18430,N_14634,N_15235);
xor U18431 (N_18431,N_14900,N_14400);
or U18432 (N_18432,N_12130,N_14781);
or U18433 (N_18433,N_12061,N_12073);
nor U18434 (N_18434,N_12649,N_14201);
and U18435 (N_18435,N_14221,N_14701);
or U18436 (N_18436,N_15236,N_12671);
or U18437 (N_18437,N_14813,N_15976);
and U18438 (N_18438,N_14374,N_12867);
or U18439 (N_18439,N_15823,N_13924);
nor U18440 (N_18440,N_12877,N_12327);
nand U18441 (N_18441,N_12960,N_12696);
or U18442 (N_18442,N_15148,N_14785);
or U18443 (N_18443,N_12742,N_15654);
or U18444 (N_18444,N_15681,N_14025);
and U18445 (N_18445,N_13496,N_13565);
nand U18446 (N_18446,N_13927,N_12864);
or U18447 (N_18447,N_13641,N_12830);
xor U18448 (N_18448,N_14927,N_12527);
xor U18449 (N_18449,N_13345,N_14439);
and U18450 (N_18450,N_14268,N_13941);
xnor U18451 (N_18451,N_12876,N_12749);
and U18452 (N_18452,N_15239,N_12650);
xor U18453 (N_18453,N_14188,N_15755);
nor U18454 (N_18454,N_14197,N_12418);
and U18455 (N_18455,N_12388,N_12500);
nand U18456 (N_18456,N_14601,N_14586);
xnor U18457 (N_18457,N_12451,N_15282);
and U18458 (N_18458,N_14957,N_14318);
and U18459 (N_18459,N_15893,N_13405);
nand U18460 (N_18460,N_15220,N_13484);
nor U18461 (N_18461,N_12948,N_12083);
xor U18462 (N_18462,N_12667,N_14760);
nor U18463 (N_18463,N_13974,N_13780);
and U18464 (N_18464,N_13982,N_12454);
xnor U18465 (N_18465,N_14395,N_13997);
nor U18466 (N_18466,N_13086,N_13253);
or U18467 (N_18467,N_14735,N_15272);
xnor U18468 (N_18468,N_15039,N_12575);
and U18469 (N_18469,N_14128,N_14355);
nor U18470 (N_18470,N_15234,N_15051);
and U18471 (N_18471,N_15711,N_15827);
xnor U18472 (N_18472,N_13297,N_15615);
and U18473 (N_18473,N_13934,N_14755);
nor U18474 (N_18474,N_15470,N_15209);
xor U18475 (N_18475,N_12616,N_15879);
and U18476 (N_18476,N_12480,N_13773);
nand U18477 (N_18477,N_13772,N_14531);
or U18478 (N_18478,N_14917,N_14798);
and U18479 (N_18479,N_12599,N_15903);
xnor U18480 (N_18480,N_12772,N_14005);
and U18481 (N_18481,N_14438,N_13292);
or U18482 (N_18482,N_12790,N_14854);
or U18483 (N_18483,N_14341,N_13776);
and U18484 (N_18484,N_15957,N_15174);
xnor U18485 (N_18485,N_15125,N_13043);
xnor U18486 (N_18486,N_14220,N_12435);
or U18487 (N_18487,N_13397,N_12333);
nor U18488 (N_18488,N_15566,N_14752);
nor U18489 (N_18489,N_12069,N_15869);
nor U18490 (N_18490,N_15736,N_12281);
xnor U18491 (N_18491,N_12703,N_12395);
or U18492 (N_18492,N_12141,N_15910);
and U18493 (N_18493,N_14250,N_12296);
and U18494 (N_18494,N_15690,N_15276);
and U18495 (N_18495,N_14834,N_12736);
xor U18496 (N_18496,N_15427,N_15511);
nor U18497 (N_18497,N_14896,N_14179);
and U18498 (N_18498,N_12731,N_15527);
nor U18499 (N_18499,N_15291,N_13582);
or U18500 (N_18500,N_15616,N_14249);
xnor U18501 (N_18501,N_13267,N_14030);
and U18502 (N_18502,N_14262,N_12252);
xnor U18503 (N_18503,N_13350,N_15027);
nand U18504 (N_18504,N_13812,N_13914);
xnor U18505 (N_18505,N_12232,N_12353);
nand U18506 (N_18506,N_13938,N_12172);
or U18507 (N_18507,N_15560,N_14426);
nand U18508 (N_18508,N_14344,N_14566);
nor U18509 (N_18509,N_13747,N_15009);
and U18510 (N_18510,N_12356,N_12221);
nand U18511 (N_18511,N_15236,N_13181);
or U18512 (N_18512,N_14189,N_15185);
nor U18513 (N_18513,N_14799,N_12011);
and U18514 (N_18514,N_14650,N_13761);
or U18515 (N_18515,N_13825,N_12934);
nand U18516 (N_18516,N_12215,N_14729);
xor U18517 (N_18517,N_15080,N_15093);
nand U18518 (N_18518,N_13148,N_14690);
or U18519 (N_18519,N_14675,N_12713);
xor U18520 (N_18520,N_12920,N_12928);
and U18521 (N_18521,N_13961,N_15011);
and U18522 (N_18522,N_13730,N_12507);
nand U18523 (N_18523,N_13857,N_14696);
and U18524 (N_18524,N_12916,N_12768);
nor U18525 (N_18525,N_13654,N_15507);
and U18526 (N_18526,N_12913,N_14864);
xor U18527 (N_18527,N_12846,N_12936);
or U18528 (N_18528,N_12440,N_14336);
and U18529 (N_18529,N_13458,N_14861);
nand U18530 (N_18530,N_13559,N_13454);
xor U18531 (N_18531,N_14766,N_12380);
xor U18532 (N_18532,N_13082,N_12249);
and U18533 (N_18533,N_15478,N_15516);
nor U18534 (N_18534,N_13170,N_15676);
and U18535 (N_18535,N_13226,N_15290);
or U18536 (N_18536,N_15029,N_14197);
nand U18537 (N_18537,N_13914,N_12700);
and U18538 (N_18538,N_14730,N_14006);
nor U18539 (N_18539,N_15249,N_13823);
nor U18540 (N_18540,N_13750,N_12412);
nand U18541 (N_18541,N_12936,N_12828);
or U18542 (N_18542,N_12694,N_14042);
nor U18543 (N_18543,N_13737,N_14541);
nor U18544 (N_18544,N_12288,N_12941);
nand U18545 (N_18545,N_14740,N_15352);
nor U18546 (N_18546,N_13387,N_12272);
xor U18547 (N_18547,N_13957,N_13153);
xnor U18548 (N_18548,N_14364,N_12609);
nor U18549 (N_18549,N_15998,N_15401);
xnor U18550 (N_18550,N_12329,N_14306);
xnor U18551 (N_18551,N_12701,N_14253);
nor U18552 (N_18552,N_15690,N_13439);
and U18553 (N_18553,N_13580,N_14189);
and U18554 (N_18554,N_13408,N_14455);
and U18555 (N_18555,N_12915,N_13393);
nand U18556 (N_18556,N_12911,N_13331);
nand U18557 (N_18557,N_13909,N_14800);
nor U18558 (N_18558,N_13174,N_12161);
and U18559 (N_18559,N_14847,N_14084);
or U18560 (N_18560,N_14011,N_13161);
or U18561 (N_18561,N_15260,N_12566);
xor U18562 (N_18562,N_12258,N_13853);
xor U18563 (N_18563,N_15657,N_12563);
nand U18564 (N_18564,N_15620,N_14560);
xnor U18565 (N_18565,N_13043,N_12260);
nand U18566 (N_18566,N_13482,N_12721);
xor U18567 (N_18567,N_12888,N_13226);
and U18568 (N_18568,N_12702,N_12624);
or U18569 (N_18569,N_12765,N_15488);
or U18570 (N_18570,N_14238,N_14541);
nor U18571 (N_18571,N_14406,N_13788);
xor U18572 (N_18572,N_15560,N_15646);
xnor U18573 (N_18573,N_15963,N_15120);
and U18574 (N_18574,N_15159,N_12207);
nand U18575 (N_18575,N_13002,N_12695);
xnor U18576 (N_18576,N_14898,N_15539);
xor U18577 (N_18577,N_13830,N_15069);
or U18578 (N_18578,N_13140,N_14831);
nor U18579 (N_18579,N_15142,N_14948);
xor U18580 (N_18580,N_13802,N_12856);
xnor U18581 (N_18581,N_12024,N_15289);
nand U18582 (N_18582,N_12940,N_13725);
nand U18583 (N_18583,N_12402,N_13002);
or U18584 (N_18584,N_13872,N_15363);
xor U18585 (N_18585,N_14535,N_14084);
and U18586 (N_18586,N_15304,N_15825);
nand U18587 (N_18587,N_14908,N_12038);
xor U18588 (N_18588,N_12436,N_13021);
nand U18589 (N_18589,N_15250,N_13210);
xor U18590 (N_18590,N_14805,N_14068);
nor U18591 (N_18591,N_14179,N_15453);
xor U18592 (N_18592,N_14120,N_14122);
and U18593 (N_18593,N_12455,N_13435);
nand U18594 (N_18594,N_12041,N_13728);
nand U18595 (N_18595,N_12971,N_12978);
or U18596 (N_18596,N_13039,N_13755);
xnor U18597 (N_18597,N_13414,N_13870);
or U18598 (N_18598,N_15384,N_15661);
or U18599 (N_18599,N_12555,N_14715);
xnor U18600 (N_18600,N_13690,N_12632);
nor U18601 (N_18601,N_14899,N_15825);
xnor U18602 (N_18602,N_13133,N_14702);
nand U18603 (N_18603,N_14643,N_13468);
xnor U18604 (N_18604,N_13877,N_13040);
and U18605 (N_18605,N_14473,N_13398);
xnor U18606 (N_18606,N_14307,N_15739);
nor U18607 (N_18607,N_15083,N_14589);
and U18608 (N_18608,N_12802,N_15385);
nand U18609 (N_18609,N_14668,N_14647);
or U18610 (N_18610,N_15317,N_14039);
and U18611 (N_18611,N_13824,N_13357);
nor U18612 (N_18612,N_13086,N_15144);
and U18613 (N_18613,N_12741,N_13577);
and U18614 (N_18614,N_12994,N_15190);
xor U18615 (N_18615,N_15544,N_15372);
nor U18616 (N_18616,N_13915,N_12698);
nor U18617 (N_18617,N_15511,N_15269);
xnor U18618 (N_18618,N_13539,N_13383);
or U18619 (N_18619,N_15821,N_14326);
nor U18620 (N_18620,N_15191,N_15279);
nand U18621 (N_18621,N_14062,N_13664);
xor U18622 (N_18622,N_12367,N_15145);
nand U18623 (N_18623,N_12921,N_14838);
and U18624 (N_18624,N_14366,N_15927);
nand U18625 (N_18625,N_12205,N_12312);
nand U18626 (N_18626,N_14141,N_13958);
nor U18627 (N_18627,N_15510,N_15338);
or U18628 (N_18628,N_12667,N_12656);
nor U18629 (N_18629,N_12402,N_13110);
nand U18630 (N_18630,N_13858,N_15008);
nand U18631 (N_18631,N_12310,N_15372);
or U18632 (N_18632,N_13611,N_12000);
nand U18633 (N_18633,N_15063,N_15819);
and U18634 (N_18634,N_15981,N_12070);
and U18635 (N_18635,N_13480,N_12355);
nand U18636 (N_18636,N_12272,N_14431);
nand U18637 (N_18637,N_14051,N_13376);
nor U18638 (N_18638,N_13353,N_12114);
or U18639 (N_18639,N_14337,N_14355);
xnor U18640 (N_18640,N_15816,N_13184);
nand U18641 (N_18641,N_14698,N_14597);
nor U18642 (N_18642,N_12560,N_12020);
nor U18643 (N_18643,N_12665,N_12269);
and U18644 (N_18644,N_15120,N_14922);
xnor U18645 (N_18645,N_13246,N_15228);
xnor U18646 (N_18646,N_14678,N_15536);
or U18647 (N_18647,N_15934,N_14650);
or U18648 (N_18648,N_14240,N_14194);
and U18649 (N_18649,N_12975,N_13777);
xor U18650 (N_18650,N_13496,N_12603);
nand U18651 (N_18651,N_14230,N_15453);
nor U18652 (N_18652,N_13592,N_13665);
nand U18653 (N_18653,N_12820,N_14087);
or U18654 (N_18654,N_15717,N_15554);
nand U18655 (N_18655,N_14355,N_13326);
or U18656 (N_18656,N_13683,N_12347);
nand U18657 (N_18657,N_14270,N_14394);
or U18658 (N_18658,N_15672,N_15579);
nand U18659 (N_18659,N_15037,N_13576);
nand U18660 (N_18660,N_15783,N_13034);
or U18661 (N_18661,N_15585,N_15685);
nand U18662 (N_18662,N_15031,N_14199);
nor U18663 (N_18663,N_13318,N_15268);
and U18664 (N_18664,N_15696,N_15290);
xnor U18665 (N_18665,N_12393,N_15068);
nand U18666 (N_18666,N_13889,N_14208);
or U18667 (N_18667,N_14517,N_12625);
xnor U18668 (N_18668,N_13502,N_12715);
nor U18669 (N_18669,N_12115,N_15075);
nand U18670 (N_18670,N_12753,N_13471);
nand U18671 (N_18671,N_13346,N_14635);
or U18672 (N_18672,N_15767,N_14172);
nor U18673 (N_18673,N_13947,N_14345);
nor U18674 (N_18674,N_13894,N_13317);
and U18675 (N_18675,N_14090,N_12596);
or U18676 (N_18676,N_13992,N_12504);
and U18677 (N_18677,N_15213,N_12763);
nand U18678 (N_18678,N_13213,N_12335);
and U18679 (N_18679,N_15312,N_12244);
nor U18680 (N_18680,N_14880,N_14909);
and U18681 (N_18681,N_12610,N_12823);
nor U18682 (N_18682,N_12748,N_14931);
nor U18683 (N_18683,N_14549,N_14594);
or U18684 (N_18684,N_12906,N_14748);
nand U18685 (N_18685,N_15983,N_15188);
xnor U18686 (N_18686,N_13401,N_13399);
xnor U18687 (N_18687,N_14553,N_12160);
nor U18688 (N_18688,N_15753,N_15197);
nor U18689 (N_18689,N_15663,N_13533);
or U18690 (N_18690,N_14528,N_14143);
or U18691 (N_18691,N_14547,N_12974);
and U18692 (N_18692,N_15116,N_14056);
or U18693 (N_18693,N_14890,N_12232);
and U18694 (N_18694,N_14938,N_14740);
or U18695 (N_18695,N_15303,N_12401);
and U18696 (N_18696,N_12966,N_15994);
nor U18697 (N_18697,N_15048,N_12430);
xnor U18698 (N_18698,N_14801,N_15136);
nor U18699 (N_18699,N_12095,N_14029);
or U18700 (N_18700,N_15315,N_13570);
nand U18701 (N_18701,N_14345,N_13937);
nor U18702 (N_18702,N_14482,N_13315);
and U18703 (N_18703,N_15068,N_15368);
nand U18704 (N_18704,N_15620,N_14903);
nand U18705 (N_18705,N_13596,N_12680);
or U18706 (N_18706,N_13168,N_13645);
nand U18707 (N_18707,N_13346,N_14851);
and U18708 (N_18708,N_13193,N_15401);
or U18709 (N_18709,N_15106,N_15518);
xnor U18710 (N_18710,N_12006,N_12351);
or U18711 (N_18711,N_15741,N_12633);
and U18712 (N_18712,N_15195,N_12721);
nand U18713 (N_18713,N_12627,N_14112);
or U18714 (N_18714,N_12928,N_14564);
or U18715 (N_18715,N_15080,N_14086);
or U18716 (N_18716,N_13137,N_12148);
and U18717 (N_18717,N_12750,N_15559);
nand U18718 (N_18718,N_13000,N_12264);
xnor U18719 (N_18719,N_15208,N_14788);
nor U18720 (N_18720,N_14867,N_12357);
xor U18721 (N_18721,N_15694,N_14455);
and U18722 (N_18722,N_12897,N_12104);
and U18723 (N_18723,N_15277,N_13241);
nand U18724 (N_18724,N_13428,N_13666);
and U18725 (N_18725,N_14277,N_12163);
nand U18726 (N_18726,N_13985,N_12162);
and U18727 (N_18727,N_14172,N_15979);
or U18728 (N_18728,N_15383,N_15883);
xnor U18729 (N_18729,N_15801,N_14540);
xnor U18730 (N_18730,N_12842,N_12366);
or U18731 (N_18731,N_13864,N_13827);
or U18732 (N_18732,N_14671,N_13775);
nand U18733 (N_18733,N_12930,N_13164);
or U18734 (N_18734,N_12094,N_15514);
nand U18735 (N_18735,N_15939,N_14152);
or U18736 (N_18736,N_14861,N_12087);
xnor U18737 (N_18737,N_14687,N_15011);
nand U18738 (N_18738,N_15427,N_14627);
nor U18739 (N_18739,N_15049,N_13262);
and U18740 (N_18740,N_14256,N_15241);
xor U18741 (N_18741,N_15965,N_15261);
and U18742 (N_18742,N_15257,N_15786);
nand U18743 (N_18743,N_13166,N_13835);
or U18744 (N_18744,N_13198,N_15037);
nand U18745 (N_18745,N_15309,N_12522);
xnor U18746 (N_18746,N_13273,N_12675);
nand U18747 (N_18747,N_13789,N_15853);
nor U18748 (N_18748,N_15077,N_15383);
xor U18749 (N_18749,N_12256,N_12027);
nor U18750 (N_18750,N_14519,N_13321);
nand U18751 (N_18751,N_12229,N_13338);
or U18752 (N_18752,N_12120,N_15123);
and U18753 (N_18753,N_13348,N_15654);
nand U18754 (N_18754,N_13561,N_15125);
nand U18755 (N_18755,N_12305,N_13329);
or U18756 (N_18756,N_13597,N_15216);
nand U18757 (N_18757,N_14405,N_13661);
nor U18758 (N_18758,N_13359,N_12756);
or U18759 (N_18759,N_14438,N_13056);
and U18760 (N_18760,N_12964,N_14755);
and U18761 (N_18761,N_14567,N_12169);
and U18762 (N_18762,N_12831,N_13289);
nand U18763 (N_18763,N_13768,N_14260);
nand U18764 (N_18764,N_14592,N_15723);
nand U18765 (N_18765,N_14450,N_12045);
and U18766 (N_18766,N_12882,N_14686);
nor U18767 (N_18767,N_12748,N_12783);
nor U18768 (N_18768,N_14644,N_15589);
xnor U18769 (N_18769,N_13960,N_14451);
and U18770 (N_18770,N_13461,N_15003);
or U18771 (N_18771,N_14924,N_13658);
nor U18772 (N_18772,N_12426,N_15225);
xnor U18773 (N_18773,N_13084,N_12837);
nor U18774 (N_18774,N_15599,N_15023);
and U18775 (N_18775,N_14384,N_13775);
or U18776 (N_18776,N_15155,N_12417);
nor U18777 (N_18777,N_15637,N_12871);
or U18778 (N_18778,N_15393,N_15503);
nand U18779 (N_18779,N_15056,N_13819);
xnor U18780 (N_18780,N_15906,N_15880);
or U18781 (N_18781,N_15467,N_14061);
or U18782 (N_18782,N_12325,N_13682);
and U18783 (N_18783,N_13443,N_12229);
nand U18784 (N_18784,N_13827,N_15091);
nor U18785 (N_18785,N_14888,N_13836);
and U18786 (N_18786,N_12455,N_14779);
nand U18787 (N_18787,N_14769,N_14009);
xor U18788 (N_18788,N_14657,N_13962);
and U18789 (N_18789,N_15117,N_12180);
and U18790 (N_18790,N_12952,N_15814);
xor U18791 (N_18791,N_12011,N_14834);
or U18792 (N_18792,N_15642,N_12722);
xor U18793 (N_18793,N_15246,N_13120);
nand U18794 (N_18794,N_15823,N_14624);
and U18795 (N_18795,N_12785,N_15986);
nand U18796 (N_18796,N_14520,N_12834);
nor U18797 (N_18797,N_13987,N_12077);
nor U18798 (N_18798,N_15226,N_14258);
and U18799 (N_18799,N_14521,N_14081);
and U18800 (N_18800,N_15949,N_14903);
or U18801 (N_18801,N_14966,N_13980);
and U18802 (N_18802,N_14057,N_12779);
xnor U18803 (N_18803,N_13167,N_12509);
nand U18804 (N_18804,N_15470,N_14043);
nand U18805 (N_18805,N_13047,N_14509);
and U18806 (N_18806,N_15736,N_12909);
xor U18807 (N_18807,N_14080,N_14058);
xnor U18808 (N_18808,N_13961,N_14585);
nand U18809 (N_18809,N_15226,N_12510);
nor U18810 (N_18810,N_15080,N_15957);
or U18811 (N_18811,N_14721,N_12288);
nand U18812 (N_18812,N_15582,N_14766);
nor U18813 (N_18813,N_13210,N_14352);
nor U18814 (N_18814,N_12070,N_13277);
and U18815 (N_18815,N_12120,N_15605);
and U18816 (N_18816,N_12940,N_15685);
xnor U18817 (N_18817,N_13910,N_15198);
or U18818 (N_18818,N_13397,N_13469);
nor U18819 (N_18819,N_15283,N_15572);
nand U18820 (N_18820,N_15012,N_13433);
and U18821 (N_18821,N_12799,N_12090);
nand U18822 (N_18822,N_14789,N_15286);
nor U18823 (N_18823,N_14037,N_14708);
or U18824 (N_18824,N_13517,N_15469);
nor U18825 (N_18825,N_12784,N_13840);
nor U18826 (N_18826,N_12830,N_13867);
xnor U18827 (N_18827,N_15532,N_12668);
or U18828 (N_18828,N_13474,N_13846);
or U18829 (N_18829,N_15810,N_12625);
or U18830 (N_18830,N_14279,N_14394);
nor U18831 (N_18831,N_14049,N_14219);
or U18832 (N_18832,N_14595,N_13097);
and U18833 (N_18833,N_15107,N_12948);
or U18834 (N_18834,N_12150,N_14331);
xor U18835 (N_18835,N_12612,N_13642);
and U18836 (N_18836,N_12111,N_13387);
nor U18837 (N_18837,N_12168,N_12274);
nor U18838 (N_18838,N_12140,N_14852);
xnor U18839 (N_18839,N_12746,N_15658);
or U18840 (N_18840,N_14778,N_15067);
xor U18841 (N_18841,N_13959,N_12386);
nand U18842 (N_18842,N_13125,N_15949);
or U18843 (N_18843,N_13850,N_15809);
or U18844 (N_18844,N_13926,N_13908);
nand U18845 (N_18845,N_12008,N_12940);
xnor U18846 (N_18846,N_13524,N_12703);
nor U18847 (N_18847,N_15806,N_13549);
and U18848 (N_18848,N_14572,N_13353);
or U18849 (N_18849,N_13621,N_13007);
nand U18850 (N_18850,N_14392,N_13126);
or U18851 (N_18851,N_14243,N_13393);
nand U18852 (N_18852,N_14682,N_13222);
nand U18853 (N_18853,N_14206,N_14122);
and U18854 (N_18854,N_14743,N_13515);
xor U18855 (N_18855,N_15783,N_12912);
or U18856 (N_18856,N_15858,N_13533);
nand U18857 (N_18857,N_13307,N_13446);
and U18858 (N_18858,N_13622,N_12332);
nand U18859 (N_18859,N_14315,N_12876);
nor U18860 (N_18860,N_14383,N_14168);
nand U18861 (N_18861,N_15919,N_13577);
xnor U18862 (N_18862,N_15621,N_14147);
xor U18863 (N_18863,N_14197,N_13254);
and U18864 (N_18864,N_15630,N_15581);
xnor U18865 (N_18865,N_12737,N_14881);
or U18866 (N_18866,N_12216,N_12044);
and U18867 (N_18867,N_13522,N_15498);
or U18868 (N_18868,N_13034,N_12346);
nor U18869 (N_18869,N_12328,N_12422);
or U18870 (N_18870,N_13921,N_14837);
xor U18871 (N_18871,N_14966,N_13742);
or U18872 (N_18872,N_13665,N_12562);
or U18873 (N_18873,N_13300,N_15813);
or U18874 (N_18874,N_14346,N_13693);
nor U18875 (N_18875,N_15422,N_14318);
nor U18876 (N_18876,N_14955,N_14244);
and U18877 (N_18877,N_15862,N_15880);
nor U18878 (N_18878,N_12604,N_15213);
nor U18879 (N_18879,N_12644,N_15596);
nand U18880 (N_18880,N_15693,N_14265);
nor U18881 (N_18881,N_13427,N_14916);
nor U18882 (N_18882,N_12053,N_12436);
xor U18883 (N_18883,N_15059,N_12679);
or U18884 (N_18884,N_12803,N_15128);
nor U18885 (N_18885,N_12432,N_12001);
nor U18886 (N_18886,N_12168,N_15527);
nand U18887 (N_18887,N_13960,N_12604);
and U18888 (N_18888,N_13368,N_13279);
nand U18889 (N_18889,N_14926,N_13451);
nor U18890 (N_18890,N_15463,N_13751);
nand U18891 (N_18891,N_12296,N_12132);
and U18892 (N_18892,N_15141,N_13734);
xnor U18893 (N_18893,N_14296,N_13004);
xnor U18894 (N_18894,N_15836,N_15165);
nor U18895 (N_18895,N_15582,N_14937);
and U18896 (N_18896,N_13342,N_14290);
or U18897 (N_18897,N_14619,N_12782);
or U18898 (N_18898,N_14509,N_13857);
or U18899 (N_18899,N_13871,N_13321);
or U18900 (N_18900,N_12889,N_15834);
and U18901 (N_18901,N_12486,N_14780);
or U18902 (N_18902,N_14678,N_13890);
and U18903 (N_18903,N_13962,N_12465);
nand U18904 (N_18904,N_12016,N_12926);
or U18905 (N_18905,N_12655,N_13814);
nor U18906 (N_18906,N_12682,N_13273);
nand U18907 (N_18907,N_13551,N_12407);
nand U18908 (N_18908,N_12014,N_14111);
nor U18909 (N_18909,N_12358,N_13693);
nand U18910 (N_18910,N_12522,N_13564);
or U18911 (N_18911,N_13139,N_14047);
nand U18912 (N_18912,N_13515,N_12127);
and U18913 (N_18913,N_15673,N_14728);
nor U18914 (N_18914,N_13811,N_12589);
nor U18915 (N_18915,N_15415,N_12059);
nand U18916 (N_18916,N_13091,N_12378);
nand U18917 (N_18917,N_14384,N_14151);
xnor U18918 (N_18918,N_15689,N_15145);
nand U18919 (N_18919,N_13076,N_15155);
and U18920 (N_18920,N_15819,N_14856);
nand U18921 (N_18921,N_14123,N_13614);
or U18922 (N_18922,N_12107,N_14637);
nor U18923 (N_18923,N_15721,N_15848);
nor U18924 (N_18924,N_15538,N_15508);
and U18925 (N_18925,N_15968,N_13298);
and U18926 (N_18926,N_14988,N_15722);
nand U18927 (N_18927,N_14779,N_15247);
or U18928 (N_18928,N_15839,N_15579);
nor U18929 (N_18929,N_13351,N_15185);
or U18930 (N_18930,N_15107,N_12694);
nand U18931 (N_18931,N_15358,N_15105);
nand U18932 (N_18932,N_12988,N_13740);
or U18933 (N_18933,N_13582,N_13645);
or U18934 (N_18934,N_14110,N_12781);
and U18935 (N_18935,N_15949,N_13764);
nand U18936 (N_18936,N_14499,N_12613);
and U18937 (N_18937,N_13422,N_15298);
nand U18938 (N_18938,N_12914,N_12702);
and U18939 (N_18939,N_12628,N_12697);
and U18940 (N_18940,N_12320,N_13951);
xor U18941 (N_18941,N_13841,N_15228);
nand U18942 (N_18942,N_14913,N_13911);
nor U18943 (N_18943,N_12020,N_14660);
nand U18944 (N_18944,N_14723,N_13939);
and U18945 (N_18945,N_13422,N_14113);
and U18946 (N_18946,N_15327,N_13785);
and U18947 (N_18947,N_14247,N_15597);
nor U18948 (N_18948,N_13290,N_12344);
nor U18949 (N_18949,N_12834,N_13056);
xor U18950 (N_18950,N_13792,N_13870);
nor U18951 (N_18951,N_14346,N_12760);
or U18952 (N_18952,N_14354,N_12710);
nand U18953 (N_18953,N_14618,N_12982);
and U18954 (N_18954,N_15629,N_15566);
nor U18955 (N_18955,N_12754,N_15050);
xor U18956 (N_18956,N_13196,N_14507);
or U18957 (N_18957,N_14134,N_13688);
xor U18958 (N_18958,N_14772,N_14292);
or U18959 (N_18959,N_12423,N_13919);
xor U18960 (N_18960,N_12000,N_15619);
nand U18961 (N_18961,N_15451,N_12839);
and U18962 (N_18962,N_14357,N_15524);
nor U18963 (N_18963,N_13347,N_13309);
and U18964 (N_18964,N_14739,N_15773);
nor U18965 (N_18965,N_13208,N_15262);
and U18966 (N_18966,N_14842,N_15143);
and U18967 (N_18967,N_12665,N_15482);
nor U18968 (N_18968,N_13114,N_13286);
nand U18969 (N_18969,N_15286,N_14619);
or U18970 (N_18970,N_12382,N_15823);
nor U18971 (N_18971,N_13263,N_14989);
xnor U18972 (N_18972,N_14364,N_15022);
nor U18973 (N_18973,N_15272,N_14348);
or U18974 (N_18974,N_14515,N_15768);
xor U18975 (N_18975,N_12047,N_15780);
xor U18976 (N_18976,N_15304,N_13070);
nor U18977 (N_18977,N_13096,N_14336);
or U18978 (N_18978,N_12258,N_14684);
or U18979 (N_18979,N_13107,N_12162);
nor U18980 (N_18980,N_13240,N_14257);
nor U18981 (N_18981,N_14519,N_15526);
and U18982 (N_18982,N_14220,N_13797);
nand U18983 (N_18983,N_15381,N_13516);
xnor U18984 (N_18984,N_14891,N_13274);
xor U18985 (N_18985,N_15495,N_13149);
or U18986 (N_18986,N_14287,N_12301);
nor U18987 (N_18987,N_15590,N_15602);
nand U18988 (N_18988,N_13924,N_13833);
and U18989 (N_18989,N_14804,N_12839);
or U18990 (N_18990,N_15754,N_15215);
nand U18991 (N_18991,N_13974,N_15986);
nand U18992 (N_18992,N_15898,N_14144);
nand U18993 (N_18993,N_13421,N_13878);
and U18994 (N_18994,N_13371,N_12269);
xnor U18995 (N_18995,N_12852,N_15344);
nor U18996 (N_18996,N_14374,N_15753);
or U18997 (N_18997,N_15697,N_12328);
nor U18998 (N_18998,N_13074,N_13574);
xnor U18999 (N_18999,N_15967,N_14710);
xnor U19000 (N_19000,N_12704,N_15017);
xnor U19001 (N_19001,N_14716,N_14208);
nor U19002 (N_19002,N_13070,N_15430);
xor U19003 (N_19003,N_15709,N_13631);
and U19004 (N_19004,N_12654,N_13873);
nor U19005 (N_19005,N_12890,N_12576);
and U19006 (N_19006,N_12457,N_12703);
nand U19007 (N_19007,N_14780,N_14503);
nand U19008 (N_19008,N_13482,N_13063);
xor U19009 (N_19009,N_13220,N_12781);
nand U19010 (N_19010,N_13509,N_12945);
or U19011 (N_19011,N_13798,N_13677);
nand U19012 (N_19012,N_12195,N_13403);
or U19013 (N_19013,N_12376,N_14974);
and U19014 (N_19014,N_14551,N_13790);
or U19015 (N_19015,N_12016,N_12410);
nor U19016 (N_19016,N_13095,N_12799);
or U19017 (N_19017,N_15023,N_14151);
and U19018 (N_19018,N_13299,N_14537);
xor U19019 (N_19019,N_13405,N_13519);
nor U19020 (N_19020,N_12974,N_12721);
or U19021 (N_19021,N_12793,N_12588);
nand U19022 (N_19022,N_15863,N_15259);
or U19023 (N_19023,N_15684,N_14914);
nor U19024 (N_19024,N_15331,N_12273);
xnor U19025 (N_19025,N_12768,N_13466);
or U19026 (N_19026,N_12155,N_13342);
nor U19027 (N_19027,N_15664,N_12613);
xnor U19028 (N_19028,N_15323,N_15356);
and U19029 (N_19029,N_12368,N_12788);
or U19030 (N_19030,N_12419,N_12423);
or U19031 (N_19031,N_15125,N_15592);
nor U19032 (N_19032,N_15574,N_14547);
xnor U19033 (N_19033,N_12194,N_14786);
or U19034 (N_19034,N_13819,N_15259);
and U19035 (N_19035,N_14173,N_13886);
or U19036 (N_19036,N_13525,N_14950);
xnor U19037 (N_19037,N_13153,N_13777);
or U19038 (N_19038,N_13471,N_12999);
nand U19039 (N_19039,N_15556,N_12333);
and U19040 (N_19040,N_12084,N_15071);
xor U19041 (N_19041,N_13209,N_15714);
xnor U19042 (N_19042,N_14284,N_14847);
or U19043 (N_19043,N_14164,N_13790);
xnor U19044 (N_19044,N_15399,N_15122);
xor U19045 (N_19045,N_15074,N_15209);
nand U19046 (N_19046,N_13636,N_14924);
and U19047 (N_19047,N_12447,N_13032);
nand U19048 (N_19048,N_12200,N_14675);
nand U19049 (N_19049,N_13888,N_12638);
and U19050 (N_19050,N_13418,N_14706);
and U19051 (N_19051,N_14205,N_12898);
or U19052 (N_19052,N_12845,N_14701);
and U19053 (N_19053,N_12127,N_13129);
and U19054 (N_19054,N_12200,N_13672);
and U19055 (N_19055,N_14045,N_14801);
or U19056 (N_19056,N_15242,N_13108);
nor U19057 (N_19057,N_15986,N_15592);
and U19058 (N_19058,N_13886,N_12493);
xor U19059 (N_19059,N_15548,N_14875);
nand U19060 (N_19060,N_15061,N_15283);
nand U19061 (N_19061,N_13482,N_14749);
xnor U19062 (N_19062,N_13811,N_13440);
nand U19063 (N_19063,N_12764,N_13536);
xnor U19064 (N_19064,N_13494,N_15428);
nand U19065 (N_19065,N_15388,N_13124);
nor U19066 (N_19066,N_13234,N_12560);
nor U19067 (N_19067,N_14128,N_13606);
or U19068 (N_19068,N_15340,N_13958);
nand U19069 (N_19069,N_12907,N_14473);
and U19070 (N_19070,N_14968,N_15529);
nand U19071 (N_19071,N_12089,N_15912);
nand U19072 (N_19072,N_13549,N_14544);
and U19073 (N_19073,N_13586,N_13298);
and U19074 (N_19074,N_14210,N_13543);
nand U19075 (N_19075,N_15950,N_13216);
and U19076 (N_19076,N_15631,N_12215);
nor U19077 (N_19077,N_15673,N_15054);
xor U19078 (N_19078,N_13070,N_12573);
or U19079 (N_19079,N_13973,N_12589);
nor U19080 (N_19080,N_14119,N_13649);
nand U19081 (N_19081,N_13835,N_15248);
and U19082 (N_19082,N_12030,N_15836);
and U19083 (N_19083,N_13166,N_14465);
nand U19084 (N_19084,N_13548,N_15611);
nor U19085 (N_19085,N_13977,N_12255);
or U19086 (N_19086,N_15571,N_14036);
nor U19087 (N_19087,N_15452,N_14821);
nor U19088 (N_19088,N_14935,N_14121);
nor U19089 (N_19089,N_14706,N_12071);
or U19090 (N_19090,N_12926,N_13597);
xor U19091 (N_19091,N_15781,N_12579);
nor U19092 (N_19092,N_12103,N_14312);
nor U19093 (N_19093,N_12223,N_15512);
nand U19094 (N_19094,N_13268,N_15103);
nand U19095 (N_19095,N_14363,N_15412);
and U19096 (N_19096,N_14400,N_13231);
xnor U19097 (N_19097,N_12733,N_12205);
nand U19098 (N_19098,N_14074,N_15610);
and U19099 (N_19099,N_15377,N_13639);
or U19100 (N_19100,N_15002,N_15192);
xnor U19101 (N_19101,N_12026,N_14740);
or U19102 (N_19102,N_12856,N_14751);
and U19103 (N_19103,N_15836,N_13410);
or U19104 (N_19104,N_15600,N_12822);
or U19105 (N_19105,N_13315,N_15942);
and U19106 (N_19106,N_14935,N_14122);
nor U19107 (N_19107,N_15719,N_13713);
nand U19108 (N_19108,N_12921,N_15363);
or U19109 (N_19109,N_15344,N_12408);
and U19110 (N_19110,N_15943,N_14136);
or U19111 (N_19111,N_14259,N_12918);
and U19112 (N_19112,N_14910,N_15489);
and U19113 (N_19113,N_15848,N_15433);
and U19114 (N_19114,N_13623,N_12593);
nor U19115 (N_19115,N_15623,N_14245);
xor U19116 (N_19116,N_12805,N_14026);
nor U19117 (N_19117,N_12004,N_14611);
and U19118 (N_19118,N_13370,N_15088);
nor U19119 (N_19119,N_15906,N_13634);
and U19120 (N_19120,N_14305,N_14487);
or U19121 (N_19121,N_15596,N_15394);
or U19122 (N_19122,N_15009,N_14003);
and U19123 (N_19123,N_13807,N_13214);
xnor U19124 (N_19124,N_12120,N_14963);
nand U19125 (N_19125,N_14024,N_12750);
or U19126 (N_19126,N_15544,N_13235);
and U19127 (N_19127,N_13912,N_15579);
or U19128 (N_19128,N_13869,N_12171);
xor U19129 (N_19129,N_14856,N_15513);
nand U19130 (N_19130,N_12614,N_14107);
nand U19131 (N_19131,N_12184,N_14767);
xor U19132 (N_19132,N_12828,N_13887);
and U19133 (N_19133,N_14477,N_14953);
and U19134 (N_19134,N_13336,N_13553);
or U19135 (N_19135,N_14364,N_12172);
nand U19136 (N_19136,N_15819,N_14032);
or U19137 (N_19137,N_15317,N_13231);
nor U19138 (N_19138,N_14216,N_15509);
xor U19139 (N_19139,N_15650,N_15328);
and U19140 (N_19140,N_15963,N_13497);
and U19141 (N_19141,N_12018,N_12734);
nand U19142 (N_19142,N_14519,N_13694);
or U19143 (N_19143,N_15921,N_13757);
or U19144 (N_19144,N_15907,N_14095);
xnor U19145 (N_19145,N_14703,N_12462);
nor U19146 (N_19146,N_14357,N_14552);
xor U19147 (N_19147,N_15597,N_12183);
or U19148 (N_19148,N_12640,N_15424);
nand U19149 (N_19149,N_12696,N_12536);
or U19150 (N_19150,N_15732,N_13751);
xnor U19151 (N_19151,N_12818,N_13714);
nor U19152 (N_19152,N_14220,N_14837);
and U19153 (N_19153,N_12768,N_12804);
or U19154 (N_19154,N_14572,N_12809);
nand U19155 (N_19155,N_13152,N_13351);
nand U19156 (N_19156,N_13739,N_14901);
nand U19157 (N_19157,N_15917,N_15196);
xnor U19158 (N_19158,N_13111,N_13176);
nand U19159 (N_19159,N_14150,N_13274);
xnor U19160 (N_19160,N_13728,N_14661);
nor U19161 (N_19161,N_15042,N_15517);
nor U19162 (N_19162,N_12588,N_12113);
and U19163 (N_19163,N_12080,N_14068);
nor U19164 (N_19164,N_14311,N_14985);
or U19165 (N_19165,N_13052,N_12280);
xor U19166 (N_19166,N_13017,N_12637);
nand U19167 (N_19167,N_13644,N_13784);
nor U19168 (N_19168,N_14082,N_15797);
xnor U19169 (N_19169,N_15417,N_14488);
and U19170 (N_19170,N_13171,N_14058);
nor U19171 (N_19171,N_14814,N_14534);
nand U19172 (N_19172,N_13051,N_15307);
nand U19173 (N_19173,N_13722,N_13117);
nor U19174 (N_19174,N_12610,N_15465);
or U19175 (N_19175,N_15491,N_13197);
nor U19176 (N_19176,N_13025,N_14162);
or U19177 (N_19177,N_12883,N_13314);
xor U19178 (N_19178,N_13252,N_12172);
and U19179 (N_19179,N_12011,N_15306);
or U19180 (N_19180,N_13460,N_15356);
nand U19181 (N_19181,N_15985,N_14937);
and U19182 (N_19182,N_14377,N_15445);
and U19183 (N_19183,N_15378,N_15404);
nor U19184 (N_19184,N_15966,N_13194);
nand U19185 (N_19185,N_14283,N_15911);
xor U19186 (N_19186,N_12217,N_14756);
and U19187 (N_19187,N_15355,N_15633);
nand U19188 (N_19188,N_12570,N_12501);
xnor U19189 (N_19189,N_13227,N_13165);
nand U19190 (N_19190,N_15966,N_13034);
nor U19191 (N_19191,N_13075,N_15709);
and U19192 (N_19192,N_15042,N_13944);
or U19193 (N_19193,N_14222,N_15577);
or U19194 (N_19194,N_12658,N_13966);
xnor U19195 (N_19195,N_14630,N_13527);
and U19196 (N_19196,N_12782,N_12131);
or U19197 (N_19197,N_15833,N_15920);
or U19198 (N_19198,N_13948,N_13224);
nand U19199 (N_19199,N_13043,N_12146);
or U19200 (N_19200,N_13679,N_13209);
or U19201 (N_19201,N_13393,N_13853);
and U19202 (N_19202,N_12680,N_14547);
xnor U19203 (N_19203,N_14435,N_15864);
nor U19204 (N_19204,N_12501,N_12514);
nor U19205 (N_19205,N_15398,N_15357);
or U19206 (N_19206,N_14392,N_15568);
or U19207 (N_19207,N_12595,N_14559);
and U19208 (N_19208,N_15331,N_12918);
xnor U19209 (N_19209,N_13726,N_12353);
nor U19210 (N_19210,N_15355,N_14949);
nor U19211 (N_19211,N_12868,N_15986);
xor U19212 (N_19212,N_14683,N_15467);
nor U19213 (N_19213,N_14893,N_15637);
or U19214 (N_19214,N_12256,N_12185);
and U19215 (N_19215,N_12758,N_15442);
xnor U19216 (N_19216,N_14274,N_12313);
and U19217 (N_19217,N_15305,N_12731);
and U19218 (N_19218,N_12332,N_12165);
nand U19219 (N_19219,N_12124,N_15341);
nand U19220 (N_19220,N_13436,N_14014);
and U19221 (N_19221,N_15858,N_13790);
or U19222 (N_19222,N_13538,N_14304);
xor U19223 (N_19223,N_12478,N_14895);
xor U19224 (N_19224,N_15876,N_15358);
or U19225 (N_19225,N_15367,N_13763);
nand U19226 (N_19226,N_13786,N_12317);
and U19227 (N_19227,N_14911,N_15663);
nor U19228 (N_19228,N_15987,N_14100);
xor U19229 (N_19229,N_13453,N_12048);
xnor U19230 (N_19230,N_15232,N_14487);
nor U19231 (N_19231,N_12283,N_14869);
or U19232 (N_19232,N_14587,N_15265);
nor U19233 (N_19233,N_15922,N_14632);
nor U19234 (N_19234,N_14238,N_14337);
nor U19235 (N_19235,N_14240,N_14184);
and U19236 (N_19236,N_12098,N_14777);
nor U19237 (N_19237,N_13718,N_14324);
or U19238 (N_19238,N_13356,N_13652);
and U19239 (N_19239,N_12212,N_14691);
nand U19240 (N_19240,N_13833,N_13418);
and U19241 (N_19241,N_13664,N_12557);
or U19242 (N_19242,N_13178,N_12093);
nand U19243 (N_19243,N_13472,N_13622);
nor U19244 (N_19244,N_12552,N_15949);
nor U19245 (N_19245,N_15367,N_15113);
or U19246 (N_19246,N_13473,N_15719);
and U19247 (N_19247,N_15107,N_15537);
and U19248 (N_19248,N_13470,N_14116);
nor U19249 (N_19249,N_12538,N_13796);
and U19250 (N_19250,N_13850,N_15796);
or U19251 (N_19251,N_15133,N_15287);
nand U19252 (N_19252,N_13693,N_14476);
and U19253 (N_19253,N_14250,N_15206);
or U19254 (N_19254,N_15990,N_14677);
nor U19255 (N_19255,N_15519,N_13657);
or U19256 (N_19256,N_13722,N_14009);
and U19257 (N_19257,N_15742,N_15154);
nor U19258 (N_19258,N_13440,N_14142);
xnor U19259 (N_19259,N_13671,N_13793);
xor U19260 (N_19260,N_15432,N_15238);
and U19261 (N_19261,N_13922,N_15839);
or U19262 (N_19262,N_14894,N_14164);
nor U19263 (N_19263,N_14814,N_15572);
and U19264 (N_19264,N_13756,N_15940);
xnor U19265 (N_19265,N_15932,N_15469);
or U19266 (N_19266,N_14208,N_12138);
xnor U19267 (N_19267,N_13739,N_12275);
xor U19268 (N_19268,N_13209,N_14796);
and U19269 (N_19269,N_14681,N_14410);
nand U19270 (N_19270,N_14906,N_14028);
xnor U19271 (N_19271,N_14522,N_15700);
and U19272 (N_19272,N_12297,N_15641);
xnor U19273 (N_19273,N_13076,N_12112);
nand U19274 (N_19274,N_12360,N_12674);
nor U19275 (N_19275,N_13344,N_15994);
or U19276 (N_19276,N_15703,N_13097);
and U19277 (N_19277,N_13764,N_15581);
xor U19278 (N_19278,N_12680,N_12805);
or U19279 (N_19279,N_14760,N_15871);
xnor U19280 (N_19280,N_12700,N_12818);
nand U19281 (N_19281,N_14128,N_13318);
and U19282 (N_19282,N_14892,N_12210);
and U19283 (N_19283,N_13126,N_12887);
nand U19284 (N_19284,N_15991,N_15140);
xor U19285 (N_19285,N_14850,N_13514);
or U19286 (N_19286,N_14469,N_14336);
nand U19287 (N_19287,N_15430,N_15530);
nand U19288 (N_19288,N_12394,N_12787);
nor U19289 (N_19289,N_13030,N_15738);
xnor U19290 (N_19290,N_13283,N_12439);
nor U19291 (N_19291,N_12935,N_15099);
nor U19292 (N_19292,N_12715,N_14988);
and U19293 (N_19293,N_14575,N_14462);
nand U19294 (N_19294,N_12176,N_12177);
nand U19295 (N_19295,N_12549,N_14840);
and U19296 (N_19296,N_12449,N_13968);
xnor U19297 (N_19297,N_14205,N_15595);
or U19298 (N_19298,N_15766,N_12595);
or U19299 (N_19299,N_15877,N_13989);
and U19300 (N_19300,N_15631,N_12909);
xor U19301 (N_19301,N_15495,N_14570);
or U19302 (N_19302,N_12961,N_13547);
nand U19303 (N_19303,N_12180,N_13173);
xnor U19304 (N_19304,N_13465,N_15900);
or U19305 (N_19305,N_14002,N_12756);
nor U19306 (N_19306,N_13614,N_13693);
and U19307 (N_19307,N_13987,N_14870);
xor U19308 (N_19308,N_14649,N_15797);
nor U19309 (N_19309,N_15988,N_15876);
and U19310 (N_19310,N_13115,N_13863);
xor U19311 (N_19311,N_13593,N_15961);
nand U19312 (N_19312,N_13676,N_15142);
xnor U19313 (N_19313,N_14648,N_15310);
nand U19314 (N_19314,N_14841,N_14128);
and U19315 (N_19315,N_12044,N_14987);
and U19316 (N_19316,N_15323,N_12463);
xnor U19317 (N_19317,N_12145,N_14343);
nor U19318 (N_19318,N_13133,N_13159);
nand U19319 (N_19319,N_14262,N_12479);
xnor U19320 (N_19320,N_12750,N_15977);
and U19321 (N_19321,N_12806,N_15523);
and U19322 (N_19322,N_13373,N_12003);
nand U19323 (N_19323,N_14993,N_15073);
nor U19324 (N_19324,N_15556,N_15953);
and U19325 (N_19325,N_15867,N_13219);
nand U19326 (N_19326,N_13576,N_13289);
or U19327 (N_19327,N_14605,N_15454);
and U19328 (N_19328,N_14184,N_12547);
nor U19329 (N_19329,N_15394,N_12758);
nor U19330 (N_19330,N_14045,N_12992);
or U19331 (N_19331,N_14280,N_13059);
xor U19332 (N_19332,N_15398,N_13692);
nand U19333 (N_19333,N_15991,N_14911);
nor U19334 (N_19334,N_12323,N_12827);
or U19335 (N_19335,N_12504,N_12128);
nor U19336 (N_19336,N_12201,N_15685);
or U19337 (N_19337,N_13054,N_12460);
nand U19338 (N_19338,N_13449,N_13695);
xnor U19339 (N_19339,N_14154,N_15932);
xnor U19340 (N_19340,N_14593,N_14807);
xor U19341 (N_19341,N_14761,N_15583);
xnor U19342 (N_19342,N_13285,N_12404);
or U19343 (N_19343,N_15270,N_15810);
nand U19344 (N_19344,N_15064,N_13403);
xor U19345 (N_19345,N_12994,N_12779);
and U19346 (N_19346,N_12605,N_15465);
nor U19347 (N_19347,N_12865,N_14305);
nor U19348 (N_19348,N_15431,N_13331);
and U19349 (N_19349,N_12678,N_15882);
or U19350 (N_19350,N_13228,N_14259);
nor U19351 (N_19351,N_15403,N_13549);
xnor U19352 (N_19352,N_15775,N_15415);
or U19353 (N_19353,N_14088,N_12715);
nor U19354 (N_19354,N_15283,N_13036);
or U19355 (N_19355,N_15414,N_12658);
or U19356 (N_19356,N_15773,N_12294);
and U19357 (N_19357,N_15308,N_13342);
and U19358 (N_19358,N_13559,N_12286);
xor U19359 (N_19359,N_15747,N_15030);
xnor U19360 (N_19360,N_15748,N_13039);
and U19361 (N_19361,N_12589,N_12471);
nor U19362 (N_19362,N_14363,N_12142);
xnor U19363 (N_19363,N_14884,N_15013);
xor U19364 (N_19364,N_12176,N_15496);
or U19365 (N_19365,N_13065,N_14729);
and U19366 (N_19366,N_12223,N_14485);
and U19367 (N_19367,N_13771,N_14010);
nand U19368 (N_19368,N_14714,N_12798);
xnor U19369 (N_19369,N_15227,N_12133);
nand U19370 (N_19370,N_13579,N_12102);
nand U19371 (N_19371,N_13172,N_13642);
xnor U19372 (N_19372,N_12074,N_14853);
xor U19373 (N_19373,N_15666,N_15220);
nand U19374 (N_19374,N_14286,N_15933);
and U19375 (N_19375,N_12086,N_14515);
nor U19376 (N_19376,N_14518,N_13350);
or U19377 (N_19377,N_12612,N_12633);
nand U19378 (N_19378,N_14317,N_15726);
and U19379 (N_19379,N_12074,N_13256);
and U19380 (N_19380,N_14197,N_13856);
xnor U19381 (N_19381,N_14911,N_13476);
and U19382 (N_19382,N_14128,N_15337);
or U19383 (N_19383,N_12378,N_12053);
xor U19384 (N_19384,N_14815,N_15415);
xnor U19385 (N_19385,N_15692,N_14800);
xnor U19386 (N_19386,N_13081,N_12544);
and U19387 (N_19387,N_15691,N_12564);
nor U19388 (N_19388,N_14186,N_15881);
or U19389 (N_19389,N_14986,N_15490);
xor U19390 (N_19390,N_14530,N_15052);
and U19391 (N_19391,N_14183,N_14751);
nor U19392 (N_19392,N_12285,N_14212);
or U19393 (N_19393,N_12472,N_15876);
nor U19394 (N_19394,N_14611,N_15477);
nor U19395 (N_19395,N_13295,N_14678);
and U19396 (N_19396,N_13484,N_13725);
or U19397 (N_19397,N_13292,N_14969);
or U19398 (N_19398,N_13803,N_12278);
nand U19399 (N_19399,N_13839,N_14419);
and U19400 (N_19400,N_12165,N_13058);
and U19401 (N_19401,N_13658,N_14499);
nand U19402 (N_19402,N_15129,N_13531);
and U19403 (N_19403,N_12338,N_15031);
or U19404 (N_19404,N_13764,N_13347);
nor U19405 (N_19405,N_12938,N_15816);
nand U19406 (N_19406,N_14993,N_14699);
nor U19407 (N_19407,N_15757,N_13261);
and U19408 (N_19408,N_13021,N_15205);
nand U19409 (N_19409,N_13510,N_12512);
nor U19410 (N_19410,N_13574,N_12922);
xor U19411 (N_19411,N_14476,N_13048);
nand U19412 (N_19412,N_13703,N_12453);
xor U19413 (N_19413,N_15216,N_15281);
and U19414 (N_19414,N_14191,N_14174);
or U19415 (N_19415,N_12190,N_13506);
xnor U19416 (N_19416,N_12805,N_13672);
or U19417 (N_19417,N_12901,N_12214);
or U19418 (N_19418,N_12197,N_14191);
nand U19419 (N_19419,N_15749,N_12579);
nor U19420 (N_19420,N_12259,N_12570);
xor U19421 (N_19421,N_14027,N_12248);
and U19422 (N_19422,N_13722,N_14461);
or U19423 (N_19423,N_13806,N_14714);
or U19424 (N_19424,N_15873,N_12816);
nand U19425 (N_19425,N_13425,N_15451);
and U19426 (N_19426,N_13368,N_15661);
or U19427 (N_19427,N_14213,N_15245);
and U19428 (N_19428,N_14876,N_12792);
xor U19429 (N_19429,N_15446,N_13375);
or U19430 (N_19430,N_12449,N_14412);
nand U19431 (N_19431,N_13446,N_13879);
nor U19432 (N_19432,N_14805,N_12340);
nand U19433 (N_19433,N_15456,N_13619);
nand U19434 (N_19434,N_14644,N_12257);
or U19435 (N_19435,N_14179,N_14041);
xnor U19436 (N_19436,N_12533,N_14039);
and U19437 (N_19437,N_15388,N_15082);
nor U19438 (N_19438,N_14382,N_13879);
nand U19439 (N_19439,N_12474,N_12688);
and U19440 (N_19440,N_13267,N_13569);
xnor U19441 (N_19441,N_12052,N_14752);
nand U19442 (N_19442,N_13068,N_12355);
nor U19443 (N_19443,N_12372,N_15646);
nand U19444 (N_19444,N_12379,N_12929);
nand U19445 (N_19445,N_14859,N_15380);
nor U19446 (N_19446,N_12965,N_12373);
nor U19447 (N_19447,N_15434,N_12541);
xnor U19448 (N_19448,N_15375,N_13663);
nand U19449 (N_19449,N_13497,N_14691);
xor U19450 (N_19450,N_13064,N_12591);
nand U19451 (N_19451,N_13200,N_13089);
xnor U19452 (N_19452,N_15259,N_13274);
nor U19453 (N_19453,N_14811,N_13415);
and U19454 (N_19454,N_12202,N_15088);
nor U19455 (N_19455,N_12835,N_14216);
nand U19456 (N_19456,N_12715,N_12435);
nand U19457 (N_19457,N_15605,N_15841);
xor U19458 (N_19458,N_14974,N_15893);
nor U19459 (N_19459,N_15508,N_12128);
and U19460 (N_19460,N_12075,N_12238);
and U19461 (N_19461,N_14469,N_12244);
nand U19462 (N_19462,N_15669,N_13161);
or U19463 (N_19463,N_15924,N_14702);
and U19464 (N_19464,N_15076,N_12908);
xnor U19465 (N_19465,N_13881,N_15325);
or U19466 (N_19466,N_13112,N_14716);
nand U19467 (N_19467,N_15136,N_13973);
xor U19468 (N_19468,N_13826,N_13687);
nand U19469 (N_19469,N_13635,N_14833);
nand U19470 (N_19470,N_13521,N_14874);
and U19471 (N_19471,N_12169,N_14467);
xor U19472 (N_19472,N_14878,N_14980);
and U19473 (N_19473,N_14013,N_15152);
xor U19474 (N_19474,N_15910,N_15992);
or U19475 (N_19475,N_12835,N_12710);
nor U19476 (N_19476,N_12419,N_13976);
nand U19477 (N_19477,N_14535,N_14438);
and U19478 (N_19478,N_12091,N_15881);
and U19479 (N_19479,N_15579,N_12085);
or U19480 (N_19480,N_15764,N_15807);
nor U19481 (N_19481,N_15765,N_12286);
or U19482 (N_19482,N_14641,N_14413);
xor U19483 (N_19483,N_15027,N_15032);
nor U19484 (N_19484,N_14880,N_13009);
nand U19485 (N_19485,N_15525,N_15069);
nand U19486 (N_19486,N_15519,N_14771);
xnor U19487 (N_19487,N_15171,N_15162);
and U19488 (N_19488,N_13958,N_12203);
xor U19489 (N_19489,N_13183,N_13217);
nor U19490 (N_19490,N_13821,N_13759);
or U19491 (N_19491,N_14330,N_14218);
and U19492 (N_19492,N_12977,N_15430);
and U19493 (N_19493,N_14455,N_13971);
or U19494 (N_19494,N_14124,N_14454);
nand U19495 (N_19495,N_13667,N_12635);
nand U19496 (N_19496,N_14952,N_14430);
xnor U19497 (N_19497,N_15156,N_15038);
or U19498 (N_19498,N_13951,N_15712);
xnor U19499 (N_19499,N_12569,N_14596);
or U19500 (N_19500,N_14636,N_15671);
nor U19501 (N_19501,N_13287,N_12489);
nand U19502 (N_19502,N_15922,N_15641);
nor U19503 (N_19503,N_14778,N_13845);
or U19504 (N_19504,N_12148,N_12574);
nor U19505 (N_19505,N_15679,N_15161);
and U19506 (N_19506,N_15223,N_14485);
xor U19507 (N_19507,N_13883,N_14096);
xor U19508 (N_19508,N_15078,N_15329);
xnor U19509 (N_19509,N_14898,N_14285);
nor U19510 (N_19510,N_15538,N_14320);
or U19511 (N_19511,N_14019,N_13060);
or U19512 (N_19512,N_15709,N_12149);
and U19513 (N_19513,N_12918,N_12722);
nor U19514 (N_19514,N_14063,N_12841);
nand U19515 (N_19515,N_15985,N_12388);
xor U19516 (N_19516,N_15288,N_14184);
nand U19517 (N_19517,N_12156,N_12648);
and U19518 (N_19518,N_13697,N_14423);
nor U19519 (N_19519,N_14941,N_13508);
nand U19520 (N_19520,N_14258,N_13557);
and U19521 (N_19521,N_13639,N_13832);
nand U19522 (N_19522,N_14289,N_13815);
nand U19523 (N_19523,N_12446,N_12542);
xnor U19524 (N_19524,N_13829,N_12742);
and U19525 (N_19525,N_14137,N_13614);
nor U19526 (N_19526,N_15286,N_14821);
or U19527 (N_19527,N_12027,N_14952);
nand U19528 (N_19528,N_13618,N_13248);
and U19529 (N_19529,N_12329,N_14168);
nor U19530 (N_19530,N_13647,N_15464);
nor U19531 (N_19531,N_14960,N_12570);
nand U19532 (N_19532,N_14038,N_14158);
xnor U19533 (N_19533,N_14591,N_13828);
nor U19534 (N_19534,N_12719,N_12587);
nand U19535 (N_19535,N_12229,N_12011);
xor U19536 (N_19536,N_12825,N_12278);
nand U19537 (N_19537,N_12643,N_12605);
nor U19538 (N_19538,N_14724,N_12489);
xor U19539 (N_19539,N_14791,N_12666);
or U19540 (N_19540,N_13016,N_12572);
or U19541 (N_19541,N_15458,N_13793);
xor U19542 (N_19542,N_14166,N_14802);
nand U19543 (N_19543,N_12968,N_15673);
xnor U19544 (N_19544,N_15804,N_14700);
or U19545 (N_19545,N_13887,N_12736);
xnor U19546 (N_19546,N_12522,N_15369);
or U19547 (N_19547,N_13163,N_14406);
and U19548 (N_19548,N_12973,N_15300);
nor U19549 (N_19549,N_14977,N_13246);
nand U19550 (N_19550,N_14664,N_15722);
xnor U19551 (N_19551,N_12232,N_12252);
nand U19552 (N_19552,N_14641,N_14507);
or U19553 (N_19553,N_15906,N_15570);
and U19554 (N_19554,N_14340,N_12853);
xor U19555 (N_19555,N_12972,N_13721);
nand U19556 (N_19556,N_12025,N_14927);
xnor U19557 (N_19557,N_15879,N_15908);
xnor U19558 (N_19558,N_12759,N_14336);
and U19559 (N_19559,N_14008,N_15011);
nand U19560 (N_19560,N_13941,N_12463);
xnor U19561 (N_19561,N_14038,N_13221);
or U19562 (N_19562,N_15229,N_15415);
xor U19563 (N_19563,N_15069,N_12852);
nor U19564 (N_19564,N_14974,N_15011);
and U19565 (N_19565,N_14789,N_15525);
xnor U19566 (N_19566,N_12802,N_12219);
xor U19567 (N_19567,N_14137,N_15669);
and U19568 (N_19568,N_12173,N_14877);
and U19569 (N_19569,N_14626,N_14911);
or U19570 (N_19570,N_14778,N_14676);
or U19571 (N_19571,N_13728,N_13167);
xor U19572 (N_19572,N_12197,N_15600);
nand U19573 (N_19573,N_15852,N_15411);
nand U19574 (N_19574,N_12198,N_14065);
nand U19575 (N_19575,N_15809,N_13534);
and U19576 (N_19576,N_12719,N_15888);
xnor U19577 (N_19577,N_13724,N_13227);
xnor U19578 (N_19578,N_13024,N_15192);
and U19579 (N_19579,N_15489,N_15751);
nor U19580 (N_19580,N_14709,N_13773);
nor U19581 (N_19581,N_15450,N_13352);
and U19582 (N_19582,N_13398,N_14429);
or U19583 (N_19583,N_14502,N_12079);
xnor U19584 (N_19584,N_13629,N_15312);
nand U19585 (N_19585,N_15600,N_15479);
nor U19586 (N_19586,N_12577,N_12370);
nand U19587 (N_19587,N_13835,N_12911);
nor U19588 (N_19588,N_15936,N_15799);
nand U19589 (N_19589,N_12108,N_12426);
nand U19590 (N_19590,N_13811,N_12358);
nand U19591 (N_19591,N_14354,N_15971);
or U19592 (N_19592,N_12777,N_15899);
xnor U19593 (N_19593,N_13982,N_13522);
xor U19594 (N_19594,N_14969,N_13934);
or U19595 (N_19595,N_12267,N_13233);
xnor U19596 (N_19596,N_12206,N_12085);
or U19597 (N_19597,N_14319,N_15006);
nand U19598 (N_19598,N_13742,N_15852);
and U19599 (N_19599,N_14945,N_12685);
nor U19600 (N_19600,N_15803,N_13295);
nand U19601 (N_19601,N_14506,N_13586);
and U19602 (N_19602,N_15467,N_14199);
xnor U19603 (N_19603,N_15769,N_12545);
nand U19604 (N_19604,N_12614,N_12877);
and U19605 (N_19605,N_14768,N_12806);
or U19606 (N_19606,N_13614,N_15113);
or U19607 (N_19607,N_14445,N_13310);
nor U19608 (N_19608,N_15262,N_14229);
or U19609 (N_19609,N_13960,N_15637);
xor U19610 (N_19610,N_13610,N_15136);
or U19611 (N_19611,N_13903,N_15426);
and U19612 (N_19612,N_15937,N_12569);
xnor U19613 (N_19613,N_12374,N_15488);
nor U19614 (N_19614,N_13603,N_12553);
nor U19615 (N_19615,N_14173,N_14388);
nor U19616 (N_19616,N_14245,N_12353);
xnor U19617 (N_19617,N_14346,N_15368);
and U19618 (N_19618,N_13505,N_13694);
or U19619 (N_19619,N_13556,N_15074);
and U19620 (N_19620,N_12564,N_13043);
and U19621 (N_19621,N_12736,N_12149);
xnor U19622 (N_19622,N_12815,N_15586);
nor U19623 (N_19623,N_15152,N_13039);
and U19624 (N_19624,N_15275,N_14421);
nand U19625 (N_19625,N_13179,N_15926);
or U19626 (N_19626,N_12604,N_12409);
or U19627 (N_19627,N_14251,N_15870);
and U19628 (N_19628,N_15853,N_15108);
and U19629 (N_19629,N_15068,N_14834);
xor U19630 (N_19630,N_13099,N_13556);
nand U19631 (N_19631,N_14615,N_12624);
and U19632 (N_19632,N_12940,N_15999);
xor U19633 (N_19633,N_13067,N_13080);
nor U19634 (N_19634,N_14864,N_14180);
xor U19635 (N_19635,N_12655,N_14959);
nor U19636 (N_19636,N_12470,N_13527);
or U19637 (N_19637,N_14236,N_15856);
and U19638 (N_19638,N_13150,N_13625);
xnor U19639 (N_19639,N_12175,N_14444);
nand U19640 (N_19640,N_14960,N_14174);
nand U19641 (N_19641,N_14913,N_13864);
xnor U19642 (N_19642,N_14684,N_14941);
xor U19643 (N_19643,N_15505,N_13577);
xor U19644 (N_19644,N_13021,N_14858);
nand U19645 (N_19645,N_12657,N_12531);
or U19646 (N_19646,N_15736,N_14684);
or U19647 (N_19647,N_15511,N_13350);
nand U19648 (N_19648,N_12388,N_14324);
nand U19649 (N_19649,N_15332,N_14801);
xnor U19650 (N_19650,N_13324,N_15956);
nand U19651 (N_19651,N_14618,N_14501);
and U19652 (N_19652,N_12386,N_13010);
or U19653 (N_19653,N_15396,N_14438);
xnor U19654 (N_19654,N_13577,N_12463);
nor U19655 (N_19655,N_15701,N_15146);
xor U19656 (N_19656,N_15900,N_12507);
and U19657 (N_19657,N_13522,N_14957);
nand U19658 (N_19658,N_13079,N_12998);
and U19659 (N_19659,N_15264,N_15779);
nor U19660 (N_19660,N_13235,N_12071);
nor U19661 (N_19661,N_12735,N_15816);
xor U19662 (N_19662,N_12690,N_12675);
or U19663 (N_19663,N_13633,N_13030);
nor U19664 (N_19664,N_14134,N_12393);
xor U19665 (N_19665,N_14359,N_13029);
nand U19666 (N_19666,N_12815,N_12730);
nor U19667 (N_19667,N_14763,N_12721);
nor U19668 (N_19668,N_14934,N_14785);
and U19669 (N_19669,N_15174,N_12718);
or U19670 (N_19670,N_13976,N_15010);
xor U19671 (N_19671,N_14446,N_14038);
and U19672 (N_19672,N_14263,N_12109);
nand U19673 (N_19673,N_13736,N_13617);
and U19674 (N_19674,N_12144,N_14713);
xor U19675 (N_19675,N_15450,N_14690);
nand U19676 (N_19676,N_15932,N_15333);
nand U19677 (N_19677,N_13196,N_12209);
and U19678 (N_19678,N_14814,N_14268);
and U19679 (N_19679,N_12466,N_15540);
and U19680 (N_19680,N_12259,N_13385);
or U19681 (N_19681,N_13584,N_14309);
xor U19682 (N_19682,N_14975,N_15124);
xnor U19683 (N_19683,N_15173,N_15375);
nor U19684 (N_19684,N_12083,N_14586);
nor U19685 (N_19685,N_12153,N_14879);
xor U19686 (N_19686,N_15949,N_14444);
xnor U19687 (N_19687,N_14842,N_13069);
nor U19688 (N_19688,N_13494,N_14538);
and U19689 (N_19689,N_12775,N_15576);
nor U19690 (N_19690,N_13917,N_14209);
or U19691 (N_19691,N_13866,N_15246);
or U19692 (N_19692,N_12688,N_12162);
and U19693 (N_19693,N_12853,N_15635);
or U19694 (N_19694,N_13091,N_14469);
nor U19695 (N_19695,N_14632,N_12648);
and U19696 (N_19696,N_13458,N_15627);
or U19697 (N_19697,N_15959,N_14438);
and U19698 (N_19698,N_15783,N_13654);
xor U19699 (N_19699,N_15663,N_13289);
xor U19700 (N_19700,N_12710,N_13241);
or U19701 (N_19701,N_14960,N_14474);
xor U19702 (N_19702,N_13035,N_12195);
and U19703 (N_19703,N_13188,N_15810);
nand U19704 (N_19704,N_12274,N_12244);
and U19705 (N_19705,N_14189,N_12874);
and U19706 (N_19706,N_12540,N_14625);
and U19707 (N_19707,N_15958,N_13269);
xnor U19708 (N_19708,N_15624,N_14203);
xnor U19709 (N_19709,N_12613,N_12077);
or U19710 (N_19710,N_14163,N_14715);
or U19711 (N_19711,N_15939,N_15518);
or U19712 (N_19712,N_12032,N_13881);
or U19713 (N_19713,N_13310,N_14842);
xor U19714 (N_19714,N_13411,N_12012);
nand U19715 (N_19715,N_15446,N_12208);
xor U19716 (N_19716,N_15892,N_15891);
or U19717 (N_19717,N_14544,N_15880);
and U19718 (N_19718,N_13894,N_14441);
and U19719 (N_19719,N_13992,N_12401);
nand U19720 (N_19720,N_15970,N_13479);
nor U19721 (N_19721,N_12901,N_13049);
and U19722 (N_19722,N_12101,N_15621);
nand U19723 (N_19723,N_14897,N_15215);
nor U19724 (N_19724,N_13149,N_13643);
nor U19725 (N_19725,N_15624,N_14856);
and U19726 (N_19726,N_14962,N_12001);
xnor U19727 (N_19727,N_12208,N_14777);
nand U19728 (N_19728,N_14772,N_12301);
xor U19729 (N_19729,N_13882,N_13765);
nand U19730 (N_19730,N_13663,N_12788);
xnor U19731 (N_19731,N_12902,N_15380);
xnor U19732 (N_19732,N_14640,N_15175);
and U19733 (N_19733,N_15066,N_13821);
nand U19734 (N_19734,N_14477,N_13383);
and U19735 (N_19735,N_12056,N_14302);
or U19736 (N_19736,N_14429,N_13798);
nor U19737 (N_19737,N_15003,N_13705);
or U19738 (N_19738,N_14022,N_13809);
nor U19739 (N_19739,N_14289,N_14382);
or U19740 (N_19740,N_12497,N_13821);
and U19741 (N_19741,N_12170,N_12704);
xor U19742 (N_19742,N_15064,N_14515);
xor U19743 (N_19743,N_12943,N_13099);
and U19744 (N_19744,N_13103,N_14313);
and U19745 (N_19745,N_12674,N_13201);
xor U19746 (N_19746,N_15961,N_13107);
nor U19747 (N_19747,N_12517,N_14793);
nand U19748 (N_19748,N_12951,N_15351);
nor U19749 (N_19749,N_12237,N_13475);
and U19750 (N_19750,N_15657,N_13593);
nand U19751 (N_19751,N_12809,N_15327);
nand U19752 (N_19752,N_15413,N_13330);
xor U19753 (N_19753,N_14881,N_15051);
or U19754 (N_19754,N_15195,N_12466);
and U19755 (N_19755,N_15578,N_14181);
xnor U19756 (N_19756,N_15837,N_13055);
and U19757 (N_19757,N_12786,N_14202);
xor U19758 (N_19758,N_15197,N_13984);
nor U19759 (N_19759,N_14453,N_12820);
nor U19760 (N_19760,N_13415,N_14722);
nor U19761 (N_19761,N_13649,N_15997);
nand U19762 (N_19762,N_13217,N_15929);
and U19763 (N_19763,N_12364,N_14707);
nand U19764 (N_19764,N_13460,N_15078);
xor U19765 (N_19765,N_15726,N_12180);
nand U19766 (N_19766,N_12450,N_14182);
and U19767 (N_19767,N_12830,N_15078);
and U19768 (N_19768,N_12692,N_15395);
xnor U19769 (N_19769,N_13095,N_13710);
or U19770 (N_19770,N_14174,N_15776);
xor U19771 (N_19771,N_14118,N_15724);
and U19772 (N_19772,N_15616,N_13905);
nor U19773 (N_19773,N_15293,N_15565);
or U19774 (N_19774,N_12630,N_12844);
xnor U19775 (N_19775,N_15866,N_12636);
xor U19776 (N_19776,N_13484,N_14914);
nor U19777 (N_19777,N_13661,N_15546);
xor U19778 (N_19778,N_14776,N_13644);
xnor U19779 (N_19779,N_12526,N_12605);
nand U19780 (N_19780,N_14493,N_12703);
or U19781 (N_19781,N_13139,N_12190);
nand U19782 (N_19782,N_12413,N_12933);
xnor U19783 (N_19783,N_12519,N_15815);
or U19784 (N_19784,N_12773,N_13786);
nand U19785 (N_19785,N_13741,N_12126);
nand U19786 (N_19786,N_12489,N_13918);
or U19787 (N_19787,N_12924,N_15725);
or U19788 (N_19788,N_13375,N_12770);
or U19789 (N_19789,N_12232,N_12091);
and U19790 (N_19790,N_13503,N_12117);
nor U19791 (N_19791,N_14139,N_15227);
xnor U19792 (N_19792,N_13831,N_13422);
or U19793 (N_19793,N_15627,N_14952);
xnor U19794 (N_19794,N_13400,N_12937);
xor U19795 (N_19795,N_13446,N_12586);
xnor U19796 (N_19796,N_14779,N_12642);
xnor U19797 (N_19797,N_12897,N_13763);
xor U19798 (N_19798,N_12799,N_15965);
nor U19799 (N_19799,N_15674,N_12524);
nand U19800 (N_19800,N_13236,N_15562);
and U19801 (N_19801,N_13634,N_15963);
nand U19802 (N_19802,N_14511,N_14186);
nor U19803 (N_19803,N_15065,N_13382);
or U19804 (N_19804,N_13952,N_15170);
and U19805 (N_19805,N_13835,N_15289);
xor U19806 (N_19806,N_15480,N_13550);
xnor U19807 (N_19807,N_15056,N_15945);
nand U19808 (N_19808,N_15820,N_15203);
nand U19809 (N_19809,N_15598,N_12564);
and U19810 (N_19810,N_13674,N_12861);
or U19811 (N_19811,N_13828,N_15564);
or U19812 (N_19812,N_12633,N_14312);
nor U19813 (N_19813,N_15083,N_12777);
or U19814 (N_19814,N_12949,N_14072);
or U19815 (N_19815,N_14504,N_14379);
nand U19816 (N_19816,N_13263,N_15601);
and U19817 (N_19817,N_14350,N_15343);
nor U19818 (N_19818,N_13075,N_13522);
or U19819 (N_19819,N_15204,N_12160);
nand U19820 (N_19820,N_12424,N_13961);
nor U19821 (N_19821,N_12115,N_13508);
and U19822 (N_19822,N_12767,N_12839);
or U19823 (N_19823,N_14771,N_12719);
nand U19824 (N_19824,N_15370,N_14190);
nor U19825 (N_19825,N_12778,N_14863);
xor U19826 (N_19826,N_12466,N_14890);
nand U19827 (N_19827,N_13918,N_14820);
or U19828 (N_19828,N_15250,N_12393);
or U19829 (N_19829,N_15471,N_12901);
xor U19830 (N_19830,N_13585,N_15739);
and U19831 (N_19831,N_12876,N_12022);
xor U19832 (N_19832,N_12387,N_12226);
nand U19833 (N_19833,N_14815,N_15860);
nor U19834 (N_19834,N_15079,N_14001);
or U19835 (N_19835,N_13564,N_15407);
nand U19836 (N_19836,N_15355,N_15008);
and U19837 (N_19837,N_12868,N_13925);
nor U19838 (N_19838,N_14320,N_12297);
xnor U19839 (N_19839,N_14877,N_14978);
nor U19840 (N_19840,N_14976,N_12474);
nand U19841 (N_19841,N_12191,N_12352);
nor U19842 (N_19842,N_13675,N_15129);
xnor U19843 (N_19843,N_13550,N_15804);
or U19844 (N_19844,N_14921,N_14699);
nand U19845 (N_19845,N_13835,N_14591);
nor U19846 (N_19846,N_14560,N_15573);
xnor U19847 (N_19847,N_13669,N_12420);
nor U19848 (N_19848,N_15728,N_12026);
or U19849 (N_19849,N_15103,N_12654);
nor U19850 (N_19850,N_12143,N_14966);
xor U19851 (N_19851,N_13849,N_13311);
xnor U19852 (N_19852,N_12102,N_13898);
nand U19853 (N_19853,N_13962,N_15884);
or U19854 (N_19854,N_13585,N_15850);
nand U19855 (N_19855,N_15140,N_12333);
and U19856 (N_19856,N_12841,N_12964);
xnor U19857 (N_19857,N_14252,N_15471);
and U19858 (N_19858,N_13017,N_12609);
xnor U19859 (N_19859,N_12315,N_15881);
and U19860 (N_19860,N_15374,N_14216);
or U19861 (N_19861,N_12343,N_13231);
or U19862 (N_19862,N_13638,N_15574);
or U19863 (N_19863,N_13506,N_14516);
nand U19864 (N_19864,N_15394,N_15375);
and U19865 (N_19865,N_12298,N_13770);
xor U19866 (N_19866,N_14386,N_13527);
nor U19867 (N_19867,N_15845,N_13244);
or U19868 (N_19868,N_12660,N_15194);
nor U19869 (N_19869,N_13621,N_14183);
and U19870 (N_19870,N_12297,N_15314);
nand U19871 (N_19871,N_15340,N_13757);
xnor U19872 (N_19872,N_12795,N_14051);
nor U19873 (N_19873,N_12141,N_12440);
nor U19874 (N_19874,N_12386,N_13343);
xor U19875 (N_19875,N_13867,N_13015);
and U19876 (N_19876,N_12918,N_14233);
or U19877 (N_19877,N_14850,N_13477);
nor U19878 (N_19878,N_14117,N_14731);
or U19879 (N_19879,N_15403,N_15798);
xnor U19880 (N_19880,N_14833,N_13469);
xnor U19881 (N_19881,N_15700,N_13499);
xnor U19882 (N_19882,N_13284,N_12811);
nand U19883 (N_19883,N_13424,N_15860);
and U19884 (N_19884,N_13217,N_13887);
xor U19885 (N_19885,N_12024,N_14028);
nor U19886 (N_19886,N_14293,N_15443);
nor U19887 (N_19887,N_15534,N_14086);
nand U19888 (N_19888,N_14561,N_14580);
xor U19889 (N_19889,N_13168,N_13298);
and U19890 (N_19890,N_14602,N_12448);
and U19891 (N_19891,N_15710,N_15036);
xor U19892 (N_19892,N_13421,N_12507);
nor U19893 (N_19893,N_14216,N_12558);
and U19894 (N_19894,N_13251,N_13967);
or U19895 (N_19895,N_14741,N_14435);
and U19896 (N_19896,N_14142,N_12005);
nor U19897 (N_19897,N_12882,N_12359);
xor U19898 (N_19898,N_13717,N_13847);
nor U19899 (N_19899,N_13067,N_13268);
xor U19900 (N_19900,N_15811,N_14975);
or U19901 (N_19901,N_14166,N_14740);
and U19902 (N_19902,N_13103,N_13745);
nor U19903 (N_19903,N_14919,N_13149);
xor U19904 (N_19904,N_15458,N_14918);
nand U19905 (N_19905,N_14807,N_13040);
nand U19906 (N_19906,N_15386,N_13176);
xor U19907 (N_19907,N_12492,N_13265);
nand U19908 (N_19908,N_12951,N_15393);
xnor U19909 (N_19909,N_15738,N_14481);
xor U19910 (N_19910,N_15987,N_14383);
nand U19911 (N_19911,N_14177,N_13707);
xor U19912 (N_19912,N_15150,N_12156);
xor U19913 (N_19913,N_13633,N_13820);
xnor U19914 (N_19914,N_14713,N_12431);
xnor U19915 (N_19915,N_13868,N_12467);
xor U19916 (N_19916,N_14832,N_13939);
nor U19917 (N_19917,N_15312,N_12679);
and U19918 (N_19918,N_12351,N_14978);
xor U19919 (N_19919,N_14226,N_14580);
nor U19920 (N_19920,N_12920,N_12966);
nand U19921 (N_19921,N_15261,N_13103);
or U19922 (N_19922,N_14216,N_14641);
nand U19923 (N_19923,N_14667,N_15594);
nand U19924 (N_19924,N_14499,N_12397);
or U19925 (N_19925,N_14618,N_14435);
xor U19926 (N_19926,N_14887,N_14967);
xor U19927 (N_19927,N_15153,N_14307);
and U19928 (N_19928,N_13671,N_12506);
xor U19929 (N_19929,N_14090,N_13380);
and U19930 (N_19930,N_14487,N_12096);
and U19931 (N_19931,N_13428,N_15782);
nor U19932 (N_19932,N_15195,N_14664);
and U19933 (N_19933,N_13462,N_15170);
and U19934 (N_19934,N_15924,N_15516);
nand U19935 (N_19935,N_14257,N_13914);
nor U19936 (N_19936,N_12619,N_12955);
xor U19937 (N_19937,N_14727,N_12705);
and U19938 (N_19938,N_15551,N_12188);
xor U19939 (N_19939,N_12132,N_14605);
nand U19940 (N_19940,N_12492,N_14682);
xnor U19941 (N_19941,N_15574,N_12932);
or U19942 (N_19942,N_14211,N_13451);
nand U19943 (N_19943,N_14271,N_12209);
nor U19944 (N_19944,N_13138,N_14943);
xnor U19945 (N_19945,N_12391,N_12804);
nand U19946 (N_19946,N_15870,N_14935);
xnor U19947 (N_19947,N_15217,N_15550);
or U19948 (N_19948,N_13194,N_13898);
and U19949 (N_19949,N_14875,N_13449);
xnor U19950 (N_19950,N_12490,N_15067);
xor U19951 (N_19951,N_14576,N_14897);
xor U19952 (N_19952,N_12565,N_15851);
nor U19953 (N_19953,N_15124,N_13145);
nor U19954 (N_19954,N_12353,N_13670);
nor U19955 (N_19955,N_13670,N_14687);
xor U19956 (N_19956,N_12983,N_12811);
nor U19957 (N_19957,N_15591,N_15017);
xor U19958 (N_19958,N_12885,N_14528);
xnor U19959 (N_19959,N_13507,N_13640);
and U19960 (N_19960,N_14989,N_12012);
and U19961 (N_19961,N_12703,N_14596);
or U19962 (N_19962,N_12694,N_14364);
xor U19963 (N_19963,N_15538,N_14647);
nand U19964 (N_19964,N_14303,N_15274);
nor U19965 (N_19965,N_13363,N_14068);
nand U19966 (N_19966,N_14168,N_14368);
or U19967 (N_19967,N_12352,N_12376);
and U19968 (N_19968,N_15502,N_15501);
and U19969 (N_19969,N_13876,N_15101);
nor U19970 (N_19970,N_15513,N_15082);
xor U19971 (N_19971,N_13968,N_13925);
or U19972 (N_19972,N_13184,N_14668);
or U19973 (N_19973,N_12072,N_14460);
or U19974 (N_19974,N_14883,N_15297);
or U19975 (N_19975,N_14020,N_13230);
or U19976 (N_19976,N_12999,N_15492);
nor U19977 (N_19977,N_12924,N_13372);
nor U19978 (N_19978,N_15956,N_13365);
or U19979 (N_19979,N_14802,N_15921);
xor U19980 (N_19980,N_12178,N_15905);
xor U19981 (N_19981,N_15127,N_15699);
nor U19982 (N_19982,N_13763,N_15560);
nand U19983 (N_19983,N_15637,N_13550);
or U19984 (N_19984,N_13217,N_13007);
or U19985 (N_19985,N_13460,N_14134);
or U19986 (N_19986,N_13388,N_15407);
nand U19987 (N_19987,N_15956,N_15568);
xnor U19988 (N_19988,N_14275,N_15194);
nor U19989 (N_19989,N_15404,N_13916);
or U19990 (N_19990,N_15831,N_12512);
or U19991 (N_19991,N_15221,N_13831);
and U19992 (N_19992,N_15357,N_12289);
nor U19993 (N_19993,N_12668,N_12888);
xor U19994 (N_19994,N_13946,N_14669);
or U19995 (N_19995,N_12898,N_12753);
and U19996 (N_19996,N_14596,N_15252);
or U19997 (N_19997,N_13328,N_12138);
and U19998 (N_19998,N_14646,N_13982);
nor U19999 (N_19999,N_14321,N_14344);
xnor UO_0 (O_0,N_17805,N_17922);
nand UO_1 (O_1,N_18139,N_17095);
nand UO_2 (O_2,N_18239,N_17296);
and UO_3 (O_3,N_17357,N_17262);
nor UO_4 (O_4,N_18732,N_16020);
or UO_5 (O_5,N_17625,N_16895);
xnor UO_6 (O_6,N_17438,N_16313);
xnor UO_7 (O_7,N_19903,N_16413);
and UO_8 (O_8,N_17132,N_18831);
or UO_9 (O_9,N_16355,N_18520);
nand UO_10 (O_10,N_19690,N_16595);
nand UO_11 (O_11,N_19694,N_18272);
or UO_12 (O_12,N_18430,N_17499);
nand UO_13 (O_13,N_18173,N_16078);
and UO_14 (O_14,N_18772,N_16878);
or UO_15 (O_15,N_17003,N_16821);
and UO_16 (O_16,N_19034,N_18331);
and UO_17 (O_17,N_18653,N_19471);
nor UO_18 (O_18,N_18363,N_16926);
xnor UO_19 (O_19,N_17611,N_19066);
and UO_20 (O_20,N_19072,N_16281);
xor UO_21 (O_21,N_17530,N_18290);
or UO_22 (O_22,N_19865,N_18746);
or UO_23 (O_23,N_19809,N_16223);
nor UO_24 (O_24,N_16094,N_18843);
and UO_25 (O_25,N_16669,N_17066);
and UO_26 (O_26,N_19122,N_18518);
nor UO_27 (O_27,N_16412,N_16470);
xor UO_28 (O_28,N_16684,N_18055);
xor UO_29 (O_29,N_16351,N_17400);
nor UO_30 (O_30,N_19074,N_16051);
or UO_31 (O_31,N_18972,N_16408);
xor UO_32 (O_32,N_16201,N_17565);
or UO_33 (O_33,N_16916,N_17350);
and UO_34 (O_34,N_18293,N_18465);
or UO_35 (O_35,N_18914,N_17954);
and UO_36 (O_36,N_16573,N_16786);
nand UO_37 (O_37,N_18416,N_17420);
nor UO_38 (O_38,N_17079,N_19245);
nor UO_39 (O_39,N_18115,N_17012);
or UO_40 (O_40,N_17483,N_17308);
xor UO_41 (O_41,N_17090,N_16808);
xor UO_42 (O_42,N_17681,N_19312);
xnor UO_43 (O_43,N_18069,N_19933);
and UO_44 (O_44,N_17541,N_18533);
nand UO_45 (O_45,N_19500,N_18714);
xnor UO_46 (O_46,N_19255,N_19431);
nand UO_47 (O_47,N_19923,N_19898);
xor UO_48 (O_48,N_18094,N_17471);
nor UO_49 (O_49,N_19545,N_19221);
nand UO_50 (O_50,N_19730,N_16559);
or UO_51 (O_51,N_17594,N_18191);
xnor UO_52 (O_52,N_19417,N_17705);
or UO_53 (O_53,N_16672,N_16479);
and UO_54 (O_54,N_16892,N_16268);
nand UO_55 (O_55,N_16175,N_16165);
or UO_56 (O_56,N_18026,N_16317);
xnor UO_57 (O_57,N_19563,N_16161);
nand UO_58 (O_58,N_17761,N_17288);
nand UO_59 (O_59,N_16650,N_19727);
xnor UO_60 (O_60,N_16241,N_18281);
nor UO_61 (O_61,N_16059,N_19383);
or UO_62 (O_62,N_16577,N_19733);
nor UO_63 (O_63,N_16485,N_16216);
xor UO_64 (O_64,N_18954,N_18707);
or UO_65 (O_65,N_17547,N_16400);
nor UO_66 (O_66,N_17494,N_17279);
or UO_67 (O_67,N_18809,N_17539);
xor UO_68 (O_68,N_17669,N_17026);
or UO_69 (O_69,N_17719,N_16171);
xnor UO_70 (O_70,N_19190,N_17127);
xor UO_71 (O_71,N_17800,N_19883);
nor UO_72 (O_72,N_17624,N_18436);
xor UO_73 (O_73,N_19736,N_19161);
or UO_74 (O_74,N_17024,N_16659);
nand UO_75 (O_75,N_19956,N_19979);
and UO_76 (O_76,N_18901,N_18612);
nor UO_77 (O_77,N_18717,N_19673);
xnor UO_78 (O_78,N_19065,N_17071);
nand UO_79 (O_79,N_17216,N_18559);
nor UO_80 (O_80,N_16364,N_19951);
or UO_81 (O_81,N_19099,N_18644);
or UO_82 (O_82,N_17419,N_16826);
xor UO_83 (O_83,N_16536,N_19705);
nor UO_84 (O_84,N_16472,N_18317);
nor UO_85 (O_85,N_19095,N_17403);
nor UO_86 (O_86,N_16658,N_19256);
or UO_87 (O_87,N_16076,N_19360);
nand UO_88 (O_88,N_17889,N_19076);
nand UO_89 (O_89,N_18903,N_17323);
nand UO_90 (O_90,N_17425,N_17882);
xor UO_91 (O_91,N_18154,N_16347);
or UO_92 (O_92,N_18813,N_16637);
or UO_93 (O_93,N_17641,N_19588);
nand UO_94 (O_94,N_19743,N_16745);
nor UO_95 (O_95,N_16299,N_18542);
and UO_96 (O_96,N_18641,N_16862);
nand UO_97 (O_97,N_16775,N_16972);
xnor UO_98 (O_98,N_18906,N_17157);
nand UO_99 (O_99,N_19087,N_16079);
or UO_100 (O_100,N_17162,N_18788);
nor UO_101 (O_101,N_16064,N_17407);
and UO_102 (O_102,N_19139,N_18712);
xnor UO_103 (O_103,N_19414,N_19701);
and UO_104 (O_104,N_17172,N_17204);
or UO_105 (O_105,N_18636,N_16032);
and UO_106 (O_106,N_16893,N_16083);
or UO_107 (O_107,N_19262,N_18184);
or UO_108 (O_108,N_17595,N_16876);
nand UO_109 (O_109,N_19362,N_16462);
nor UO_110 (O_110,N_18091,N_19040);
or UO_111 (O_111,N_19550,N_16609);
nor UO_112 (O_112,N_19141,N_18930);
xor UO_113 (O_113,N_17390,N_19842);
and UO_114 (O_114,N_16785,N_19128);
and UO_115 (O_115,N_16710,N_18213);
nand UO_116 (O_116,N_17199,N_16690);
or UO_117 (O_117,N_18498,N_16586);
nand UO_118 (O_118,N_18517,N_17433);
nand UO_119 (O_119,N_17999,N_18877);
or UO_120 (O_120,N_17383,N_19918);
nand UO_121 (O_121,N_17802,N_19806);
nand UO_122 (O_122,N_16236,N_16113);
nor UO_123 (O_123,N_19821,N_16954);
xor UO_124 (O_124,N_18098,N_17015);
nand UO_125 (O_125,N_19791,N_16763);
xor UO_126 (O_126,N_16771,N_17418);
or UO_127 (O_127,N_16789,N_18480);
and UO_128 (O_128,N_16084,N_16978);
nand UO_129 (O_129,N_17720,N_17630);
nor UO_130 (O_130,N_16434,N_19257);
nand UO_131 (O_131,N_17063,N_17974);
xor UO_132 (O_132,N_19780,N_16626);
nor UO_133 (O_133,N_17727,N_17311);
or UO_134 (O_134,N_19039,N_19697);
or UO_135 (O_135,N_16103,N_18525);
xor UO_136 (O_136,N_16698,N_17502);
or UO_137 (O_137,N_19592,N_18087);
nand UO_138 (O_138,N_19770,N_18850);
nor UO_139 (O_139,N_19032,N_19014);
nand UO_140 (O_140,N_18616,N_19186);
or UO_141 (O_141,N_17074,N_19651);
nand UO_142 (O_142,N_19031,N_17245);
nand UO_143 (O_143,N_17227,N_19146);
xnor UO_144 (O_144,N_17010,N_19748);
xnor UO_145 (O_145,N_17891,N_16404);
xor UO_146 (O_146,N_16425,N_16327);
nor UO_147 (O_147,N_16029,N_18793);
or UO_148 (O_148,N_19523,N_16508);
nand UO_149 (O_149,N_19521,N_17154);
and UO_150 (O_150,N_18401,N_17743);
xor UO_151 (O_151,N_17602,N_17560);
nor UO_152 (O_152,N_17573,N_19797);
nand UO_153 (O_153,N_19193,N_16143);
xor UO_154 (O_154,N_19882,N_17214);
or UO_155 (O_155,N_19910,N_16579);
nor UO_156 (O_156,N_16499,N_16787);
and UO_157 (O_157,N_18546,N_18387);
xor UO_158 (O_158,N_18198,N_19543);
nor UO_159 (O_159,N_19771,N_19115);
or UO_160 (O_160,N_16604,N_18169);
xor UO_161 (O_161,N_18068,N_18875);
nor UO_162 (O_162,N_19790,N_16623);
xor UO_163 (O_163,N_18507,N_17294);
xor UO_164 (O_164,N_19136,N_17117);
nand UO_165 (O_165,N_17533,N_19375);
and UO_166 (O_166,N_18691,N_18593);
and UO_167 (O_167,N_19213,N_18421);
nor UO_168 (O_168,N_18816,N_17778);
or UO_169 (O_169,N_17623,N_19202);
xor UO_170 (O_170,N_18602,N_18880);
nand UO_171 (O_171,N_18858,N_18755);
or UO_172 (O_172,N_16861,N_18832);
xor UO_173 (O_173,N_17459,N_17796);
nand UO_174 (O_174,N_18164,N_18805);
nand UO_175 (O_175,N_18766,N_19063);
nor UO_176 (O_176,N_17924,N_19599);
and UO_177 (O_177,N_18127,N_18841);
and UO_178 (O_178,N_16209,N_18722);
nand UO_179 (O_179,N_16294,N_19472);
nand UO_180 (O_180,N_19699,N_19426);
or UO_181 (O_181,N_16885,N_19096);
or UO_182 (O_182,N_19579,N_18837);
and UO_183 (O_183,N_19005,N_18979);
and UO_184 (O_184,N_19456,N_17029);
nor UO_185 (O_185,N_19269,N_17041);
or UO_186 (O_186,N_19795,N_19449);
nor UO_187 (O_187,N_18202,N_16418);
xor UO_188 (O_188,N_18754,N_19985);
xnor UO_189 (O_189,N_16320,N_16751);
or UO_190 (O_190,N_19966,N_18973);
or UO_191 (O_191,N_16894,N_16133);
or UO_192 (O_192,N_16431,N_17442);
nor UO_193 (O_193,N_19636,N_18771);
and UO_194 (O_194,N_19843,N_16122);
or UO_195 (O_195,N_16461,N_18409);
xnor UO_196 (O_196,N_18427,N_18125);
and UO_197 (O_197,N_18051,N_18188);
or UO_198 (O_198,N_18304,N_17316);
or UO_199 (O_199,N_18016,N_17488);
nand UO_200 (O_200,N_16114,N_18523);
nor UO_201 (O_201,N_17057,N_18611);
or UO_202 (O_202,N_16965,N_17808);
or UO_203 (O_203,N_18578,N_16065);
xor UO_204 (O_204,N_17904,N_17476);
nor UO_205 (O_205,N_18099,N_19053);
nor UO_206 (O_206,N_16187,N_19899);
or UO_207 (O_207,N_17998,N_18340);
nor UO_208 (O_208,N_16244,N_19715);
xor UO_209 (O_209,N_16551,N_19676);
and UO_210 (O_210,N_19451,N_16641);
nand UO_211 (O_211,N_18565,N_16318);
or UO_212 (O_212,N_17171,N_17161);
and UO_213 (O_213,N_18506,N_19007);
or UO_214 (O_214,N_17485,N_17464);
nor UO_215 (O_215,N_16362,N_18660);
nor UO_216 (O_216,N_18513,N_16052);
xor UO_217 (O_217,N_19098,N_17265);
xnor UO_218 (O_218,N_18615,N_17572);
nor UO_219 (O_219,N_17859,N_17503);
and UO_220 (O_220,N_17359,N_17803);
and UO_221 (O_221,N_16359,N_17426);
or UO_222 (O_222,N_16055,N_17763);
xnor UO_223 (O_223,N_16386,N_19420);
nand UO_224 (O_224,N_19316,N_19288);
nor UO_225 (O_225,N_18854,N_19153);
or UO_226 (O_226,N_16600,N_19744);
nor UO_227 (O_227,N_16913,N_16396);
nand UO_228 (O_228,N_19050,N_18940);
nand UO_229 (O_229,N_16645,N_18534);
xnor UO_230 (O_230,N_17562,N_19224);
xor UO_231 (O_231,N_18379,N_18134);
xnor UO_232 (O_232,N_18635,N_17376);
xnor UO_233 (O_233,N_19038,N_16923);
nand UO_234 (O_234,N_18695,N_18167);
and UO_235 (O_235,N_19261,N_16360);
nand UO_236 (O_236,N_18121,N_18275);
nor UO_237 (O_237,N_16014,N_18784);
or UO_238 (O_238,N_19688,N_18935);
xnor UO_239 (O_239,N_18680,N_16633);
nor UO_240 (O_240,N_16330,N_19560);
and UO_241 (O_241,N_16819,N_19574);
nand UO_242 (O_242,N_19815,N_18742);
nor UO_243 (O_243,N_19160,N_17457);
nor UO_244 (O_244,N_18630,N_16211);
and UO_245 (O_245,N_16802,N_17021);
and UO_246 (O_246,N_17082,N_19530);
nand UO_247 (O_247,N_18392,N_19212);
xnor UO_248 (O_248,N_16679,N_17233);
nand UO_249 (O_249,N_16603,N_16120);
nand UO_250 (O_250,N_17860,N_16621);
nor UO_251 (O_251,N_19984,N_17596);
or UO_252 (O_252,N_18162,N_17759);
and UO_253 (O_253,N_18958,N_16872);
or UO_254 (O_254,N_19057,N_19369);
xor UO_255 (O_255,N_18758,N_16963);
xnor UO_256 (O_256,N_19081,N_19615);
nor UO_257 (O_257,N_16562,N_18848);
nor UO_258 (O_258,N_17421,N_19779);
xnor UO_259 (O_259,N_19011,N_18027);
nor UO_260 (O_260,N_16995,N_19515);
or UO_261 (O_261,N_16915,N_19080);
nand UO_262 (O_262,N_17219,N_17581);
and UO_263 (O_263,N_17374,N_19646);
nand UO_264 (O_264,N_17513,N_18295);
and UO_265 (O_265,N_17023,N_16448);
and UO_266 (O_266,N_16357,N_18760);
or UO_267 (O_267,N_19285,N_16410);
or UO_268 (O_268,N_16944,N_18529);
and UO_269 (O_269,N_18731,N_17121);
and UO_270 (O_270,N_17575,N_19764);
xnor UO_271 (O_271,N_17109,N_16903);
xor UO_272 (O_272,N_19195,N_17823);
nor UO_273 (O_273,N_19739,N_19091);
nand UO_274 (O_274,N_16740,N_19405);
nor UO_275 (O_275,N_16339,N_19975);
or UO_276 (O_276,N_17788,N_16050);
and UO_277 (O_277,N_16532,N_16516);
nand UO_278 (O_278,N_17437,N_16304);
nand UO_279 (O_279,N_17222,N_16261);
nor UO_280 (O_280,N_17051,N_18763);
and UO_281 (O_281,N_18528,N_18647);
xor UO_282 (O_282,N_19496,N_18283);
and UO_283 (O_283,N_18195,N_17837);
and UO_284 (O_284,N_18526,N_18938);
nor UO_285 (O_285,N_17470,N_17568);
xor UO_286 (O_286,N_17138,N_18800);
nand UO_287 (O_287,N_16452,N_17058);
xor UO_288 (O_288,N_19149,N_19816);
xor UO_289 (O_289,N_17806,N_18751);
nand UO_290 (O_290,N_17155,N_19168);
and UO_291 (O_291,N_16530,N_18962);
and UO_292 (O_292,N_17001,N_16912);
nor UO_293 (O_293,N_18496,N_16942);
or UO_294 (O_294,N_17116,N_18738);
and UO_295 (O_295,N_19434,N_19798);
and UO_296 (O_296,N_19206,N_19183);
or UO_297 (O_297,N_19029,N_17203);
or UO_298 (O_298,N_16728,N_16292);
and UO_299 (O_299,N_16678,N_17632);
or UO_300 (O_300,N_17713,N_16908);
nand UO_301 (O_301,N_17535,N_18866);
nand UO_302 (O_302,N_16146,N_17552);
nor UO_303 (O_303,N_16089,N_19859);
nor UO_304 (O_304,N_19838,N_17968);
nor UO_305 (O_305,N_19504,N_16484);
nand UO_306 (O_306,N_19056,N_16964);
xnor UO_307 (O_307,N_17570,N_19246);
xor UO_308 (O_308,N_17527,N_16665);
and UO_309 (O_309,N_16384,N_19633);
nor UO_310 (O_310,N_18560,N_18224);
and UO_311 (O_311,N_19772,N_19858);
and UO_312 (O_312,N_18050,N_17797);
or UO_313 (O_313,N_18160,N_17181);
or UO_314 (O_314,N_17258,N_18662);
nand UO_315 (O_315,N_16013,N_16156);
nor UO_316 (O_316,N_16831,N_17926);
xor UO_317 (O_317,N_16153,N_16361);
xor UO_318 (O_318,N_16858,N_17319);
or UO_319 (O_319,N_16619,N_18199);
nor UO_320 (O_320,N_18483,N_19223);
and UO_321 (O_321,N_18827,N_16909);
or UO_322 (O_322,N_19318,N_16765);
nand UO_323 (O_323,N_17887,N_18589);
nand UO_324 (O_324,N_17297,N_16841);
or UO_325 (O_325,N_16905,N_19959);
and UO_326 (O_326,N_19915,N_16128);
xnor UO_327 (O_327,N_16818,N_17179);
xnor UO_328 (O_328,N_16402,N_18092);
xor UO_329 (O_329,N_17659,N_16277);
and UO_330 (O_330,N_17923,N_17615);
nand UO_331 (O_331,N_18384,N_17396);
nor UO_332 (O_332,N_19696,N_19265);
xnor UO_333 (O_333,N_18745,N_17008);
nand UO_334 (O_334,N_16662,N_18613);
or UO_335 (O_335,N_18209,N_17993);
xnor UO_336 (O_336,N_17025,N_18690);
and UO_337 (O_337,N_16928,N_19216);
and UO_338 (O_338,N_18472,N_19308);
xor UO_339 (O_339,N_19203,N_17380);
nand UO_340 (O_340,N_18113,N_18952);
nor UO_341 (O_341,N_16697,N_17660);
or UO_342 (O_342,N_16300,N_19019);
and UO_343 (O_343,N_16343,N_16742);
and UO_344 (O_344,N_18795,N_19766);
xor UO_345 (O_345,N_18670,N_16950);
xnor UO_346 (O_346,N_19864,N_19848);
or UO_347 (O_347,N_18485,N_19547);
nor UO_348 (O_348,N_18874,N_19231);
and UO_349 (O_349,N_17062,N_18884);
nand UO_350 (O_350,N_16298,N_18457);
nor UO_351 (O_351,N_17620,N_18112);
nor UO_352 (O_352,N_17367,N_19682);
nand UO_353 (O_353,N_16139,N_16220);
or UO_354 (O_354,N_18334,N_17545);
nand UO_355 (O_355,N_19896,N_18073);
nand UO_356 (O_356,N_19296,N_19823);
xnor UO_357 (O_357,N_17783,N_16420);
nand UO_358 (O_358,N_17128,N_17080);
xnor UO_359 (O_359,N_16403,N_16456);
nand UO_360 (O_360,N_16132,N_17820);
and UO_361 (O_361,N_19954,N_16951);
nor UO_362 (O_362,N_17756,N_16254);
or UO_363 (O_363,N_19327,N_19556);
nor UO_364 (O_364,N_17139,N_17643);
or UO_365 (O_365,N_19526,N_16068);
nor UO_366 (O_366,N_16239,N_18364);
nand UO_367 (O_367,N_18614,N_18661);
nor UO_368 (O_368,N_18425,N_19897);
nor UO_369 (O_369,N_17857,N_17431);
and UO_370 (O_370,N_17867,N_16968);
or UO_371 (O_371,N_18646,N_16938);
xnor UO_372 (O_372,N_17178,N_18428);
and UO_373 (O_373,N_16323,N_16778);
xor UO_374 (O_374,N_18415,N_19716);
xor UO_375 (O_375,N_19608,N_18872);
xnor UO_376 (O_376,N_19097,N_18219);
xor UO_377 (O_377,N_18651,N_19343);
xor UO_378 (O_378,N_19884,N_16801);
nand UO_379 (O_379,N_19799,N_18978);
nand UO_380 (O_380,N_19124,N_17406);
nand UO_381 (O_381,N_17828,N_18140);
nand UO_382 (O_382,N_16038,N_16154);
nor UO_383 (O_383,N_17208,N_19323);
or UO_384 (O_384,N_16714,N_19570);
nand UO_385 (O_385,N_16019,N_18251);
nand UO_386 (O_386,N_18684,N_19960);
xor UO_387 (O_387,N_17014,N_19225);
xnor UO_388 (O_388,N_17105,N_16467);
and UO_389 (O_389,N_16601,N_17584);
or UO_390 (O_390,N_17957,N_19048);
xor UO_391 (O_391,N_18607,N_16011);
xnor UO_392 (O_392,N_18103,N_18277);
nand UO_393 (O_393,N_19501,N_16002);
and UO_394 (O_394,N_17355,N_18390);
or UO_395 (O_395,N_18354,N_19169);
nand UO_396 (O_396,N_18012,N_18944);
xnor UO_397 (O_397,N_19622,N_16733);
or UO_398 (O_398,N_16870,N_16830);
nor UO_399 (O_399,N_18204,N_19970);
nor UO_400 (O_400,N_16054,N_18532);
and UO_401 (O_401,N_18942,N_18061);
xor UO_402 (O_402,N_18945,N_17666);
or UO_403 (O_403,N_16387,N_17861);
nand UO_404 (O_404,N_16764,N_18551);
and UO_405 (O_405,N_16656,N_18564);
nand UO_406 (O_406,N_17656,N_18497);
nand UO_407 (O_407,N_18900,N_17671);
xnor UO_408 (O_408,N_16016,N_17031);
and UO_409 (O_409,N_18727,N_18923);
nor UO_410 (O_410,N_18200,N_18348);
and UO_411 (O_411,N_19925,N_19906);
nand UO_412 (O_412,N_17410,N_17149);
nand UO_413 (O_413,N_19295,N_17416);
and UO_414 (O_414,N_17781,N_16943);
nand UO_415 (O_415,N_17606,N_19601);
nand UO_416 (O_416,N_17772,N_16984);
nor UO_417 (O_417,N_16664,N_16449);
nand UO_418 (O_418,N_16811,N_16611);
nor UO_419 (O_419,N_16231,N_17475);
and UO_420 (O_420,N_17614,N_18159);
or UO_421 (O_421,N_16095,N_19656);
nand UO_422 (O_422,N_17716,N_17566);
and UO_423 (O_423,N_18461,N_19176);
or UO_424 (O_424,N_16533,N_16193);
xor UO_425 (O_425,N_17280,N_16711);
and UO_426 (O_426,N_18932,N_18448);
and UO_427 (O_427,N_17220,N_16554);
nor UO_428 (O_428,N_16702,N_19937);
nand UO_429 (O_429,N_19765,N_16306);
xnor UO_430 (O_430,N_18396,N_18654);
nor UO_431 (O_431,N_17236,N_19981);
and UO_432 (O_432,N_19982,N_16582);
nor UO_433 (O_433,N_17393,N_18381);
xnor UO_434 (O_434,N_17571,N_18860);
and UO_435 (O_435,N_18176,N_16373);
nand UO_436 (O_436,N_18898,N_16824);
nand UO_437 (O_437,N_16825,N_17901);
xnor UO_438 (O_438,N_18309,N_17622);
or UO_439 (O_439,N_19429,N_19752);
nor UO_440 (O_440,N_18752,N_16260);
nor UO_441 (O_441,N_17833,N_17723);
nor UO_442 (O_442,N_19909,N_17942);
and UO_443 (O_443,N_18132,N_19393);
nor UO_444 (O_444,N_18502,N_17588);
xor UO_445 (O_445,N_18696,N_19827);
nand UO_446 (O_446,N_17776,N_18734);
nor UO_447 (O_447,N_16377,N_19055);
nor UO_448 (O_448,N_18212,N_18385);
nor UO_449 (O_449,N_19365,N_17304);
xnor UO_450 (O_450,N_18965,N_17246);
nor UO_451 (O_451,N_17834,N_18861);
and UO_452 (O_452,N_18320,N_17771);
or UO_453 (O_453,N_16009,N_19381);
nand UO_454 (O_454,N_18287,N_18035);
or UO_455 (O_455,N_18966,N_18798);
and UO_456 (O_456,N_16585,N_18242);
or UO_457 (O_457,N_17388,N_16097);
nand UO_458 (O_458,N_16827,N_17972);
nor UO_459 (O_459,N_19814,N_17945);
nor UO_460 (O_460,N_16866,N_16003);
nand UO_461 (O_461,N_17436,N_17381);
xnor UO_462 (O_462,N_19746,N_19445);
nand UO_463 (O_463,N_18253,N_18301);
nor UO_464 (O_464,N_17697,N_18405);
or UO_465 (O_465,N_17831,N_16379);
nor UO_466 (O_466,N_16197,N_16196);
nor UO_467 (O_467,N_19747,N_18422);
and UO_468 (O_468,N_19349,N_17338);
nor UO_469 (O_469,N_18685,N_18522);
or UO_470 (O_470,N_17491,N_19654);
and UO_471 (O_471,N_18263,N_17125);
nor UO_472 (O_472,N_17306,N_16864);
or UO_473 (O_473,N_16838,N_16624);
or UO_474 (O_474,N_19969,N_19470);
and UO_475 (O_475,N_19968,N_18325);
or UO_476 (O_476,N_18270,N_18913);
and UO_477 (O_477,N_17988,N_17613);
nand UO_478 (O_478,N_18362,N_19760);
xor UO_479 (O_479,N_19667,N_19582);
nor UO_480 (O_480,N_16071,N_19494);
xor UO_481 (O_481,N_19287,N_19590);
nor UO_482 (O_482,N_16266,N_17192);
nand UO_483 (O_483,N_19524,N_18886);
nand UO_484 (O_484,N_16502,N_18006);
and UO_485 (O_485,N_19914,N_17967);
or UO_486 (O_486,N_17962,N_18137);
nor UO_487 (O_487,N_16353,N_19152);
xor UO_488 (O_488,N_19242,N_19930);
nor UO_489 (O_489,N_19596,N_17300);
nor UO_490 (O_490,N_18141,N_17890);
and UO_491 (O_491,N_16018,N_19532);
and UO_492 (O_492,N_18530,N_17352);
or UO_493 (O_493,N_18737,N_16301);
nand UO_494 (O_494,N_18241,N_19461);
xnor UO_495 (O_495,N_16026,N_17708);
nand UO_496 (O_496,N_17682,N_18245);
and UO_497 (O_497,N_16776,N_19077);
and UO_498 (O_498,N_18101,N_19527);
nor UO_499 (O_499,N_17473,N_18700);
or UO_500 (O_500,N_17270,N_17629);
nand UO_501 (O_501,N_16494,N_18269);
nor UO_502 (O_502,N_19140,N_18896);
nor UO_503 (O_503,N_17439,N_18531);
or UO_504 (O_504,N_19416,N_19713);
xor UO_505 (O_505,N_18208,N_17856);
and UO_506 (O_506,N_19710,N_19067);
xor UO_507 (O_507,N_18215,N_18868);
and UO_508 (O_508,N_19535,N_19569);
and UO_509 (O_509,N_19782,N_16227);
nand UO_510 (O_510,N_19967,N_17638);
and UO_511 (O_511,N_19692,N_19600);
xnor UO_512 (O_512,N_17740,N_19133);
and UO_513 (O_513,N_16726,N_18211);
or UO_514 (O_514,N_18587,N_18779);
nand UO_515 (O_515,N_17838,N_17042);
nor UO_516 (O_516,N_18077,N_16411);
xor UO_517 (O_517,N_16008,N_19380);
nand UO_518 (O_518,N_17460,N_18033);
nand UO_519 (O_519,N_18739,N_17885);
nand UO_520 (O_520,N_19384,N_16590);
or UO_521 (O_521,N_19228,N_16245);
or UO_522 (O_522,N_17081,N_17409);
nand UO_523 (O_523,N_18487,N_19093);
nor UO_524 (O_524,N_18135,N_19276);
and UO_525 (O_525,N_17534,N_17531);
nor UO_526 (O_526,N_17863,N_19252);
nor UO_527 (O_527,N_17709,N_16321);
nor UO_528 (O_528,N_18072,N_17871);
nand UO_529 (O_529,N_19613,N_16203);
nand UO_530 (O_530,N_17905,N_18210);
nand UO_531 (O_531,N_18667,N_16924);
or UO_532 (O_532,N_17906,N_19222);
xnor UO_533 (O_533,N_17469,N_16644);
xor UO_534 (O_534,N_16720,N_16657);
or UO_535 (O_535,N_16031,N_17553);
and UO_536 (O_536,N_19554,N_19513);
or UO_537 (O_537,N_19333,N_17718);
nand UO_538 (O_538,N_19536,N_19480);
xor UO_539 (O_539,N_18484,N_16986);
and UO_540 (O_540,N_18538,N_16112);
nand UO_541 (O_541,N_17432,N_16072);
nand UO_542 (O_542,N_17980,N_17982);
or UO_543 (O_543,N_19366,N_19507);
nand UO_544 (O_544,N_19758,N_17295);
and UO_545 (O_545,N_17362,N_17005);
or UO_546 (O_546,N_18096,N_18246);
nand UO_547 (O_547,N_16087,N_17268);
nand UO_548 (O_548,N_17549,N_17052);
and UO_549 (O_549,N_16988,N_18553);
xor UO_550 (O_550,N_16162,N_19240);
and UO_551 (O_551,N_17649,N_16759);
and UO_552 (O_552,N_17035,N_18575);
and UO_553 (O_553,N_16289,N_18781);
or UO_554 (O_554,N_17101,N_18663);
or UO_555 (O_555,N_18192,N_19350);
or UO_556 (O_556,N_19476,N_18820);
or UO_557 (O_557,N_17053,N_18438);
xor UO_558 (O_558,N_19232,N_17913);
or UO_559 (O_559,N_16842,N_19759);
xor UO_560 (O_560,N_16110,N_19244);
nand UO_561 (O_561,N_19753,N_17391);
nor UO_562 (O_562,N_16166,N_17250);
and UO_563 (O_563,N_19943,N_18366);
or UO_564 (O_564,N_16389,N_16845);
and UO_565 (O_565,N_17564,N_17912);
or UO_566 (O_566,N_16476,N_19237);
nand UO_567 (O_567,N_17399,N_17599);
nand UO_568 (O_568,N_19348,N_18687);
xor UO_569 (O_569,N_16832,N_17446);
nand UO_570 (O_570,N_16541,N_16232);
or UO_571 (O_571,N_17548,N_18312);
nand UO_572 (O_572,N_16605,N_17687);
nand UO_573 (O_573,N_16980,N_18378);
or UO_574 (O_574,N_19266,N_19948);
or UO_575 (O_575,N_16440,N_17382);
nand UO_576 (O_576,N_19593,N_18839);
nand UO_577 (O_577,N_19992,N_18961);
xor UO_578 (O_578,N_18509,N_18501);
nor UO_579 (O_579,N_17559,N_17729);
nor UO_580 (O_580,N_19172,N_16552);
nor UO_581 (O_581,N_16174,N_17508);
nand UO_582 (O_582,N_19197,N_17970);
or UO_583 (O_583,N_19397,N_18493);
or UO_584 (O_584,N_19553,N_17969);
or UO_585 (O_585,N_19044,N_17722);
or UO_586 (O_586,N_19844,N_18711);
nand UO_587 (O_587,N_16136,N_18922);
or UO_588 (O_588,N_19181,N_19155);
nand UO_589 (O_589,N_16933,N_16427);
nor UO_590 (O_590,N_19549,N_18144);
nor UO_591 (O_591,N_18371,N_16741);
or UO_592 (O_592,N_16617,N_16836);
nand UO_593 (O_593,N_18720,N_18203);
xnor UO_594 (O_594,N_19300,N_16085);
and UO_595 (O_595,N_17546,N_17160);
nor UO_596 (O_596,N_18170,N_16865);
nor UO_597 (O_597,N_17255,N_16628);
and UO_598 (O_598,N_19273,N_16075);
nand UO_599 (O_599,N_19486,N_16725);
nand UO_600 (O_600,N_19455,N_19630);
xnor UO_601 (O_601,N_17757,N_18997);
nor UO_602 (O_602,N_18036,N_18057);
nand UO_603 (O_603,N_19386,N_19990);
and UO_604 (O_604,N_16137,N_18273);
and UO_605 (O_605,N_19459,N_18910);
xor UO_606 (O_606,N_16115,N_16446);
nor UO_607 (O_607,N_18770,N_19046);
or UO_608 (O_608,N_19834,N_18076);
nor UO_609 (O_609,N_19901,N_19218);
or UO_610 (O_610,N_19407,N_16473);
and UO_611 (O_611,N_18454,N_18572);
nor UO_612 (O_612,N_19111,N_16464);
or UO_613 (O_613,N_18468,N_19317);
nand UO_614 (O_614,N_17816,N_18413);
xor UO_615 (O_615,N_18310,N_17115);
nor UO_616 (O_616,N_18492,N_19423);
or UO_617 (O_617,N_18086,N_18231);
nand UO_618 (O_618,N_19489,N_19488);
nand UO_619 (O_619,N_17443,N_16850);
or UO_620 (O_620,N_18873,N_16246);
xnor UO_621 (O_621,N_19619,N_19114);
nand UO_622 (O_622,N_19732,N_19977);
and UO_623 (O_623,N_16519,N_17617);
xor UO_624 (O_624,N_17845,N_18562);
nor UO_625 (O_625,N_16037,N_17618);
nor UO_626 (O_626,N_16217,N_17777);
and UO_627 (O_627,N_18693,N_17811);
nor UO_628 (O_628,N_16701,N_18840);
or UO_629 (O_629,N_19170,N_17879);
nor UO_630 (O_630,N_16506,N_16757);
or UO_631 (O_631,N_17894,N_16708);
nand UO_632 (O_632,N_18618,N_17018);
nor UO_633 (O_633,N_19890,N_18315);
xnor UO_634 (O_634,N_19717,N_17389);
and UO_635 (O_635,N_16800,N_18114);
or UO_636 (O_636,N_16738,N_19936);
nor UO_637 (O_637,N_17411,N_16767);
and UO_638 (O_638,N_19495,N_19587);
xor UO_639 (O_639,N_18443,N_16560);
nor UO_640 (O_640,N_17704,N_19640);
and UO_641 (O_641,N_18426,N_19525);
nand UO_642 (O_642,N_18234,N_19413);
and UO_643 (O_643,N_16340,N_18059);
nor UO_644 (O_644,N_16381,N_18014);
or UO_645 (O_645,N_16372,N_18814);
and UO_646 (O_646,N_18605,N_18929);
nor UO_647 (O_647,N_16610,N_17987);
or UO_648 (O_648,N_17078,N_16067);
nor UO_649 (O_649,N_17450,N_16371);
xnor UO_650 (O_650,N_17169,N_17324);
nor UO_651 (O_651,N_16990,N_16345);
nor UO_652 (O_652,N_18108,N_17070);
nand UO_653 (O_653,N_16206,N_18959);
or UO_654 (O_654,N_16178,N_18339);
or UO_655 (O_655,N_19670,N_16415);
nand UO_656 (O_656,N_17123,N_16392);
nand UO_657 (O_657,N_19179,N_18808);
nor UO_658 (O_658,N_18220,N_16971);
xor UO_659 (O_659,N_16048,N_16471);
nand UO_660 (O_660,N_18306,N_19757);
or UO_661 (O_661,N_19877,N_19132);
nand UO_662 (O_662,N_18626,N_19649);
and UO_663 (O_663,N_17166,N_18721);
or UO_664 (O_664,N_18276,N_16495);
xnor UO_665 (O_665,N_19347,N_16302);
nand UO_666 (O_666,N_16282,N_17337);
or UO_667 (O_667,N_18183,N_18318);
nor UO_668 (O_668,N_16293,N_17205);
xor UO_669 (O_669,N_18931,N_16525);
or UO_670 (O_670,N_19824,N_16914);
nand UO_671 (O_671,N_16730,N_16760);
nor UO_672 (O_672,N_17509,N_19928);
or UO_673 (O_673,N_16660,N_19541);
xor UO_674 (O_674,N_17846,N_16949);
or UO_675 (O_675,N_18600,N_19687);
and UO_676 (O_676,N_17445,N_16442);
xnor UO_677 (O_677,N_16140,N_19306);
nor UO_678 (O_678,N_16843,N_19478);
xor UO_679 (O_679,N_19562,N_19329);
xor UO_680 (O_680,N_17835,N_17554);
xnor UO_681 (O_681,N_19326,N_19483);
or UO_682 (O_682,N_19638,N_19851);
and UO_683 (O_683,N_19807,N_18918);
nand UO_684 (O_684,N_16338,N_19719);
and UO_685 (O_685,N_18155,N_18994);
nand UO_686 (O_686,N_18021,N_18028);
xor UO_687 (O_687,N_17981,N_18743);
xor UO_688 (O_688,N_17985,N_17586);
nor UO_689 (O_689,N_18812,N_16627);
and UO_690 (O_690,N_19102,N_16540);
nor UO_691 (O_691,N_17375,N_19891);
xor UO_692 (O_692,N_17747,N_18372);
or UO_693 (O_693,N_17069,N_16689);
xnor UO_694 (O_694,N_18597,N_18622);
nor UO_695 (O_695,N_16695,N_18268);
or UO_696 (O_696,N_16225,N_18744);
and UO_697 (O_697,N_18729,N_17020);
nand UO_698 (O_698,N_18129,N_18672);
nand UO_699 (O_699,N_18566,N_18953);
nor UO_700 (O_700,N_16940,N_19900);
nand UO_701 (O_701,N_18280,N_17866);
and UO_702 (O_702,N_18664,N_16642);
nand UO_703 (O_703,N_16534,N_16107);
xnor UO_704 (O_704,N_16931,N_18568);
nor UO_705 (O_705,N_17185,N_17461);
nand UO_706 (O_706,N_16388,N_18503);
or UO_707 (O_707,N_19411,N_16511);
nor UO_708 (O_708,N_17692,N_18311);
nand UO_709 (O_709,N_16957,N_17975);
xnor UO_710 (O_710,N_18897,N_17663);
nor UO_711 (O_711,N_19201,N_17320);
or UO_712 (O_712,N_16123,N_17850);
xor UO_713 (O_713,N_17810,N_16233);
or UO_714 (O_714,N_18638,N_17369);
xnor UO_715 (O_715,N_16907,N_16398);
and UO_716 (O_716,N_18193,N_17516);
or UO_717 (O_717,N_17271,N_18045);
and UO_718 (O_718,N_19776,N_19430);
or UO_719 (O_719,N_18040,N_16817);
or UO_720 (O_720,N_17458,N_18267);
or UO_721 (O_721,N_16074,N_16691);
and UO_722 (O_722,N_19204,N_16385);
nor UO_723 (O_723,N_18074,N_17793);
xnor UO_724 (O_724,N_17048,N_18093);
xnor UO_725 (O_725,N_18571,N_19741);
and UO_726 (O_726,N_16699,N_17273);
and UO_727 (O_727,N_17392,N_16921);
and UO_728 (O_728,N_16999,N_17263);
or UO_729 (O_729,N_19991,N_18089);
or UO_730 (O_730,N_18990,N_17394);
and UO_731 (O_731,N_18826,N_16739);
nand UO_732 (O_732,N_18624,N_17480);
xor UO_733 (O_733,N_18237,N_17941);
nor UO_734 (O_734,N_18852,N_18083);
and UO_735 (O_735,N_17318,N_17211);
and UO_736 (O_736,N_17496,N_18056);
and UO_737 (O_737,N_17868,N_17452);
xor UO_738 (O_738,N_17751,N_16257);
or UO_739 (O_739,N_19506,N_16612);
and UO_740 (O_740,N_17415,N_18955);
xor UO_741 (O_741,N_19761,N_16267);
nor UO_742 (O_742,N_17345,N_19808);
and UO_743 (O_743,N_17683,N_18004);
xor UO_744 (O_744,N_17523,N_16394);
or UO_745 (O_745,N_18512,N_19374);
nand UO_746 (O_746,N_18064,N_19085);
nand UO_747 (O_747,N_19505,N_17848);
and UO_748 (O_748,N_18674,N_16976);
nor UO_749 (O_749,N_18388,N_16010);
xnor UO_750 (O_750,N_16737,N_16788);
nor UO_751 (O_751,N_18504,N_17328);
xnor UO_752 (O_752,N_17699,N_17501);
nand UO_753 (O_753,N_17537,N_18265);
or UO_754 (O_754,N_18984,N_17137);
nor UO_755 (O_755,N_16030,N_16028);
nor UO_756 (O_756,N_16395,N_19534);
and UO_757 (O_757,N_17817,N_18123);
nor UO_758 (O_758,N_16513,N_17886);
xnor UO_759 (O_759,N_16129,N_18969);
nand UO_760 (O_760,N_18608,N_17610);
nor UO_761 (O_761,N_16955,N_16027);
or UO_762 (O_762,N_19006,N_16130);
xor UO_763 (O_763,N_17744,N_16189);
nor UO_764 (O_764,N_17385,N_16992);
nor UO_765 (O_765,N_19293,N_19177);
nand UO_766 (O_766,N_18893,N_19784);
nor UO_767 (O_767,N_17874,N_19607);
nor UO_768 (O_768,N_19718,N_16614);
nand UO_769 (O_769,N_16149,N_16109);
and UO_770 (O_770,N_18547,N_18029);
and UO_771 (O_771,N_17786,N_18833);
and UO_772 (O_772,N_18153,N_16015);
xor UO_773 (O_773,N_16295,N_17884);
nor UO_774 (O_774,N_18818,N_19831);
xor UO_775 (O_775,N_19946,N_19629);
nand UO_776 (O_776,N_16458,N_18227);
nor UO_777 (O_777,N_18133,N_16994);
nand UO_778 (O_778,N_19491,N_16514);
or UO_779 (O_779,N_17898,N_16447);
and UO_780 (O_780,N_18937,N_17767);
nor UO_781 (O_781,N_19993,N_17423);
xnor UO_782 (O_782,N_17291,N_17707);
or UO_783 (O_783,N_18181,N_18494);
nor UO_784 (O_784,N_19934,N_17574);
or UO_785 (O_785,N_17468,N_17038);
nand UO_786 (O_786,N_17500,N_17033);
nor UO_787 (O_787,N_19330,N_19291);
xnor UO_788 (O_788,N_19196,N_17978);
and UO_789 (O_789,N_19778,N_19902);
nor UO_790 (O_790,N_19116,N_16316);
and UO_791 (O_791,N_17717,N_16597);
nand UO_792 (O_792,N_17131,N_19026);
nand UO_793 (O_793,N_17881,N_19150);
and UO_794 (O_794,N_16046,N_18197);
nand UO_795 (O_795,N_19631,N_18186);
nor UO_796 (O_796,N_18975,N_18338);
and UO_797 (O_797,N_16004,N_16953);
xor UO_798 (O_798,N_17919,N_18609);
and UO_799 (O_799,N_16033,N_16521);
nor UO_800 (O_800,N_17056,N_16922);
nor UO_801 (O_801,N_19517,N_19873);
nand UO_802 (O_802,N_19371,N_17290);
nor UO_803 (O_803,N_16041,N_16546);
and UO_804 (O_804,N_18150,N_18182);
or UO_805 (O_805,N_17274,N_18569);
nand UO_806 (O_806,N_16583,N_17334);
or UO_807 (O_807,N_17193,N_16378);
nor UO_808 (O_808,N_16273,N_18190);
or UO_809 (O_809,N_18681,N_19043);
and UO_810 (O_810,N_18750,N_19822);
nand UO_811 (O_811,N_19028,N_17691);
and UO_812 (O_812,N_17854,N_19792);
nor UO_813 (O_813,N_17030,N_16224);
nand UO_814 (O_814,N_19643,N_16539);
nand UO_815 (O_815,N_19389,N_19283);
nand UO_816 (O_816,N_18920,N_19709);
xor UO_817 (O_817,N_16734,N_18095);
nand UO_818 (O_818,N_18682,N_16335);
xnor UO_819 (O_819,N_16365,N_19278);
and UO_820 (O_820,N_17472,N_17198);
and UO_821 (O_821,N_16683,N_19740);
and UO_822 (O_822,N_16564,N_17226);
or UO_823 (O_823,N_16488,N_17735);
nand UO_824 (O_824,N_19134,N_16319);
or UO_825 (O_825,N_19100,N_16671);
xnor UO_826 (O_826,N_17813,N_16797);
and UO_827 (O_827,N_19301,N_19737);
nand UO_828 (O_828,N_17909,N_16263);
or UO_829 (O_829,N_18053,N_19083);
nor UO_830 (O_830,N_19837,N_19749);
nand UO_831 (O_831,N_19767,N_16791);
nor UO_832 (O_832,N_16177,N_17801);
nor UO_833 (O_833,N_16962,N_19775);
or UO_834 (O_834,N_17944,N_19463);
nor UO_835 (O_835,N_19684,N_19800);
xnor UO_836 (O_836,N_18765,N_16634);
nand UO_837 (O_837,N_17899,N_19774);
nand UO_838 (O_838,N_19439,N_19609);
nand UO_839 (O_839,N_16444,N_19135);
and UO_840 (O_840,N_18165,N_19567);
and UO_841 (O_841,N_17165,N_16503);
and UO_842 (O_842,N_18459,N_17339);
nand UO_843 (O_843,N_18100,N_19325);
xnor UO_844 (O_844,N_19872,N_16682);
xor UO_845 (O_845,N_17332,N_17822);
and UO_846 (O_846,N_19805,N_18450);
nor UO_847 (O_847,N_19290,N_18999);
nand UO_848 (O_848,N_17371,N_16237);
nand UO_849 (O_849,N_17313,N_19401);
xnor UO_850 (O_850,N_16712,N_19514);
xor UO_851 (O_851,N_16873,N_19723);
nor UO_852 (O_852,N_19700,N_16017);
and UO_853 (O_853,N_17156,N_17603);
or UO_854 (O_854,N_18577,N_18736);
nand UO_855 (O_855,N_17135,N_18177);
nand UO_856 (O_856,N_17658,N_17243);
nor UO_857 (O_857,N_16661,N_18917);
nor UO_858 (O_858,N_16346,N_18032);
xnor UO_859 (O_859,N_16898,N_18157);
nor UO_860 (O_860,N_17883,N_19691);
nand UO_861 (O_861,N_17739,N_17929);
and UO_862 (O_862,N_17825,N_17124);
xnor UO_863 (O_863,N_17685,N_16837);
or UO_864 (O_864,N_19625,N_18617);
nor UO_865 (O_865,N_19650,N_19427);
and UO_866 (O_866,N_16520,N_17260);
nor UO_867 (O_867,N_18658,N_16341);
nand UO_868 (O_868,N_19103,N_19385);
nor UO_869 (O_869,N_19400,N_19129);
or UO_870 (O_870,N_16553,N_16407);
xnor UO_871 (O_871,N_17447,N_16615);
nand UO_872 (O_872,N_19118,N_16249);
or UO_873 (O_873,N_16192,N_19591);
xnor UO_874 (O_874,N_19829,N_19437);
nor UO_875 (O_875,N_16587,N_19487);
and UO_876 (O_876,N_17348,N_17932);
nor UO_877 (O_877,N_17915,N_16598);
and UO_878 (O_878,N_19158,N_16550);
or UO_879 (O_879,N_16145,N_18710);
or UO_880 (O_880,N_18803,N_18424);
or UO_881 (O_881,N_18998,N_19832);
nor UO_882 (O_882,N_18688,N_18490);
nand UO_883 (O_883,N_17827,N_19839);
nor UO_884 (O_884,N_18701,N_18453);
and UO_885 (O_885,N_18588,N_18289);
nand UO_886 (O_886,N_17465,N_17679);
nand UO_887 (O_887,N_16592,N_17766);
nand UO_888 (O_888,N_18733,N_18715);
nor UO_889 (O_889,N_17103,N_16429);
nor UO_890 (O_890,N_17217,N_18995);
xor UO_891 (O_891,N_19345,N_18474);
or UO_892 (O_892,N_16758,N_18433);
or UO_893 (O_893,N_19689,N_16840);
and UO_894 (O_894,N_19905,N_17307);
or UO_895 (O_895,N_16815,N_18499);
xor UO_896 (O_896,N_17888,N_18048);
nand UO_897 (O_897,N_16483,N_18407);
nand UO_898 (O_898,N_16173,N_19363);
nand UO_899 (O_899,N_16001,N_16498);
nand UO_900 (O_900,N_17147,N_18313);
or UO_901 (O_901,N_16045,N_16352);
or UO_902 (O_902,N_19572,N_17215);
nand UO_903 (O_903,N_19382,N_19332);
nor UO_904 (O_904,N_18895,N_16331);
nor UO_905 (O_905,N_17664,N_19904);
nor UO_906 (O_906,N_17853,N_19616);
xor UO_907 (O_907,N_18957,N_19321);
and UO_908 (O_908,N_18365,N_19109);
or UO_909 (O_909,N_16518,N_17202);
and UO_910 (O_910,N_18374,N_19162);
or UO_911 (O_911,N_18561,N_16368);
nand UO_912 (O_912,N_18307,N_18206);
nand UO_913 (O_913,N_19557,N_19352);
xor UO_914 (O_914,N_19756,N_17737);
or UO_915 (O_915,N_18261,N_17873);
and UO_916 (O_916,N_16329,N_19302);
nor UO_917 (O_917,N_16575,N_18777);
or UO_918 (O_918,N_16799,N_18382);
nor UO_919 (O_919,N_17164,N_18326);
nor UO_920 (O_920,N_16493,N_16896);
xor UO_921 (O_921,N_16348,N_19919);
xnor UO_922 (O_922,N_19107,N_17186);
xnor UO_923 (O_923,N_16308,N_18435);
nor UO_924 (O_924,N_17959,N_16556);
and UO_925 (O_925,N_17336,N_17481);
and UO_926 (O_926,N_18023,N_17113);
nor UO_927 (O_927,N_17938,N_19751);
nor UO_928 (O_928,N_18677,N_17449);
nand UO_929 (O_929,N_19292,N_17544);
or UO_930 (O_930,N_18604,N_19679);
nand UO_931 (O_931,N_18105,N_17301);
nand UO_932 (O_932,N_17864,N_18869);
nand UO_933 (O_933,N_18558,N_17591);
nor UO_934 (O_934,N_17206,N_19519);
nand UO_935 (O_935,N_17983,N_18226);
nor UO_936 (O_936,N_18797,N_18394);
and UO_937 (O_937,N_18718,N_19578);
nor UO_938 (O_938,N_16163,N_16234);
and UO_939 (O_939,N_16901,N_19368);
and UO_940 (O_940,N_18065,N_19922);
or UO_941 (O_941,N_17106,N_16088);
nand UO_942 (O_942,N_17903,N_18757);
xor UO_943 (O_943,N_19516,N_17765);
xnor UO_944 (O_944,N_18266,N_19452);
nand UO_945 (O_945,N_19704,N_17150);
xnor UO_946 (O_946,N_17314,N_17143);
xor UO_947 (O_947,N_17684,N_18119);
and UO_948 (O_948,N_17555,N_17519);
nand UO_949 (O_949,N_19313,N_19618);
nor UO_950 (O_950,N_19920,N_16142);
xnor UO_951 (O_951,N_18104,N_19886);
nor UO_952 (O_952,N_18031,N_18500);
and UO_953 (O_953,N_16375,N_16491);
xnor UO_954 (O_954,N_16252,N_17770);
nand UO_955 (O_955,N_16925,N_17764);
xor UO_956 (O_956,N_17726,N_18904);
or UO_957 (O_957,N_16736,N_19185);
xor UO_958 (O_958,N_18970,N_19171);
nand UO_959 (O_959,N_19324,N_17605);
or UO_960 (O_960,N_18775,N_19275);
nand UO_961 (O_961,N_17668,N_18963);
nand UO_962 (O_962,N_19681,N_18521);
nand UO_963 (O_963,N_17855,N_17696);
xnor UO_964 (O_964,N_17167,N_19319);
and UO_965 (O_965,N_19617,N_18883);
or UO_966 (O_966,N_16311,N_17830);
nand UO_967 (O_967,N_16680,N_18991);
nand UO_968 (O_968,N_19441,N_19750);
or UO_969 (O_969,N_19577,N_19395);
nor UO_970 (O_970,N_18549,N_18864);
xnor UO_971 (O_971,N_17908,N_18001);
nor UO_972 (O_972,N_16124,N_16782);
xnor UO_973 (O_973,N_18899,N_19214);
nor UO_974 (O_974,N_19184,N_19680);
xnor UO_975 (O_975,N_19840,N_19215);
nor UO_976 (O_976,N_17824,N_19000);
or UO_977 (O_977,N_19208,N_16401);
xor UO_978 (O_978,N_18038,N_19230);
xnor UO_979 (O_979,N_16127,N_17870);
or UO_980 (O_980,N_17402,N_19175);
and UO_981 (O_981,N_18330,N_19853);
or UO_982 (O_982,N_19341,N_16945);
xnor UO_983 (O_983,N_18619,N_19166);
nand UO_984 (O_984,N_16073,N_18620);
nand UO_985 (O_985,N_16445,N_16947);
xnor UO_986 (O_986,N_18637,N_17804);
nor UO_987 (O_987,N_18919,N_19314);
or UO_988 (O_988,N_17637,N_16570);
nor UO_989 (O_989,N_17344,N_17712);
or UO_990 (O_990,N_16285,N_19127);
xnor UO_991 (O_991,N_16803,N_19274);
or UO_992 (O_992,N_18025,N_19191);
and UO_993 (O_993,N_17950,N_17734);
nor UO_994 (O_994,N_19008,N_16996);
xnor UO_995 (O_995,N_19151,N_16426);
or UO_996 (O_996,N_19399,N_17928);
xnor UO_997 (O_997,N_16622,N_19089);
or UO_998 (O_998,N_17329,N_16279);
xnor UO_999 (O_999,N_17939,N_18570);
or UO_1000 (O_1000,N_17773,N_17940);
xnor UO_1001 (O_1001,N_17997,N_17521);
nor UO_1002 (O_1002,N_18423,N_17577);
or UO_1003 (O_1003,N_18563,N_17467);
and UO_1004 (O_1004,N_16526,N_19078);
nand UO_1005 (O_1005,N_17677,N_17807);
xnor UO_1006 (O_1006,N_16283,N_18058);
nand UO_1007 (O_1007,N_19916,N_19131);
nand UO_1008 (O_1008,N_16709,N_18748);
xor UO_1009 (O_1009,N_19503,N_17207);
or UO_1010 (O_1010,N_18319,N_19509);
and UO_1011 (O_1011,N_17522,N_18704);
nand UO_1012 (O_1012,N_16212,N_19086);
xnor UO_1013 (O_1013,N_18228,N_18264);
nor UO_1014 (O_1014,N_19061,N_18294);
and UO_1015 (O_1015,N_17096,N_16489);
and UO_1016 (O_1016,N_16463,N_16121);
xor UO_1017 (O_1017,N_18085,N_16258);
nand UO_1018 (O_1018,N_16416,N_18369);
and UO_1019 (O_1019,N_18846,N_16846);
nand UO_1020 (O_1020,N_19512,N_19893);
nor UO_1021 (O_1021,N_17264,N_16970);
or UO_1022 (O_1022,N_18406,N_17358);
nor UO_1023 (O_1023,N_19762,N_18708);
nor UO_1024 (O_1024,N_16205,N_18951);
nand UO_1025 (O_1025,N_17512,N_19199);
nand UO_1026 (O_1026,N_19479,N_17815);
or UO_1027 (O_1027,N_18921,N_17673);
nand UO_1028 (O_1028,N_17518,N_19989);
xor UO_1029 (O_1029,N_16569,N_16118);
or UO_1030 (O_1030,N_16250,N_16053);
nand UO_1031 (O_1031,N_16430,N_18097);
and UO_1032 (O_1032,N_18475,N_19789);
nand UO_1033 (O_1033,N_18482,N_19672);
and UO_1034 (O_1034,N_17711,N_18713);
or UO_1035 (O_1035,N_18080,N_16284);
or UO_1036 (O_1036,N_17576,N_19403);
nand UO_1037 (O_1037,N_17176,N_19342);
and UO_1038 (O_1038,N_16287,N_17067);
xnor UO_1039 (O_1039,N_16198,N_19425);
xnor UO_1040 (O_1040,N_18462,N_16989);
or UO_1041 (O_1041,N_16852,N_18432);
and UO_1042 (O_1042,N_18019,N_16510);
xor UO_1043 (O_1043,N_19745,N_18753);
and UO_1044 (O_1044,N_19391,N_17745);
nand UO_1045 (O_1045,N_18466,N_16290);
xor UO_1046 (O_1046,N_19529,N_16666);
nand UO_1047 (O_1047,N_16638,N_19714);
xnor UO_1048 (O_1048,N_17395,N_17372);
nand UO_1049 (O_1049,N_17044,N_17130);
or UO_1050 (O_1050,N_16305,N_18802);
and UO_1051 (O_1051,N_19540,N_17934);
and UO_1052 (O_1052,N_18335,N_17902);
and UO_1053 (O_1053,N_16269,N_17742);
or UO_1054 (O_1054,N_17466,N_16935);
and UO_1055 (O_1055,N_17184,N_16007);
or UO_1056 (O_1056,N_18926,N_18885);
nand UO_1057 (O_1057,N_17829,N_16883);
or UO_1058 (O_1058,N_18665,N_18907);
nor UO_1059 (O_1059,N_18557,N_17897);
xor UO_1060 (O_1060,N_17240,N_19668);
and UO_1061 (O_1061,N_16889,N_18018);
or UO_1062 (O_1062,N_19997,N_18316);
and UO_1063 (O_1063,N_18633,N_19049);
xnor UO_1064 (O_1064,N_16823,N_19473);
xnor UO_1065 (O_1065,N_18151,N_16475);
nand UO_1066 (O_1066,N_17780,N_16807);
and UO_1067 (O_1067,N_19678,N_16578);
xnor UO_1068 (O_1068,N_18207,N_17843);
and UO_1069 (O_1069,N_18889,N_18550);
nand UO_1070 (O_1070,N_19887,N_18376);
nor UO_1071 (O_1071,N_16006,N_16369);
nand UO_1072 (O_1072,N_19857,N_19156);
and UO_1073 (O_1073,N_17286,N_16497);
and UO_1074 (O_1074,N_18156,N_18686);
or UO_1075 (O_1075,N_16750,N_18789);
nor UO_1076 (O_1076,N_17036,N_18214);
nand UO_1077 (O_1077,N_19999,N_16828);
nor UO_1078 (O_1078,N_16676,N_18987);
nand UO_1079 (O_1079,N_18222,N_18463);
or UO_1080 (O_1080,N_19464,N_16397);
and UO_1081 (O_1081,N_17598,N_17118);
nand UO_1082 (O_1082,N_17910,N_16435);
nor UO_1083 (O_1083,N_17107,N_18260);
nand UO_1084 (O_1084,N_16542,N_19648);
or UO_1085 (O_1085,N_17225,N_16936);
nand UO_1086 (O_1086,N_19379,N_17784);
or UO_1087 (O_1087,N_19238,N_16576);
or UO_1088 (O_1088,N_19339,N_16956);
nand UO_1089 (O_1089,N_17492,N_16204);
nor UO_1090 (O_1090,N_19677,N_17792);
xnor UO_1091 (O_1091,N_18801,N_19159);
or UO_1092 (O_1092,N_17059,N_18735);
xnor UO_1093 (O_1093,N_19602,N_18106);
nor UO_1094 (O_1094,N_17730,N_17049);
xnor UO_1095 (O_1095,N_16024,N_18767);
and UO_1096 (O_1096,N_17917,N_16370);
nand UO_1097 (O_1097,N_19801,N_17343);
nand UO_1098 (O_1098,N_19305,N_18741);
nor UO_1099 (O_1099,N_17412,N_16755);
nand UO_1100 (O_1100,N_19833,N_16186);
or UO_1101 (O_1101,N_16286,N_17511);
nand UO_1102 (O_1102,N_19810,N_18163);
nand UO_1103 (O_1103,N_17189,N_18252);
or UO_1104 (O_1104,N_17633,N_17634);
xor UO_1105 (O_1105,N_17093,N_17931);
xor UO_1106 (O_1106,N_19950,N_19852);
xnor UO_1107 (O_1107,N_17277,N_17563);
and UO_1108 (O_1108,N_16460,N_18782);
nor UO_1109 (O_1109,N_18705,N_18337);
and UO_1110 (O_1110,N_17256,N_19973);
nand UO_1111 (O_1111,N_17144,N_17238);
and UO_1112 (O_1112,N_18440,N_17930);
or UO_1113 (O_1113,N_16276,N_16322);
xor UO_1114 (O_1114,N_17842,N_16061);
xor UO_1115 (O_1115,N_17040,N_18403);
nor UO_1116 (O_1116,N_17645,N_17746);
or UO_1117 (O_1117,N_17317,N_19537);
nand UO_1118 (O_1118,N_18044,N_17953);
nand UO_1119 (O_1119,N_19498,N_16466);
nor UO_1120 (O_1120,N_18419,N_17342);
or UO_1121 (O_1121,N_16793,N_17790);
and UO_1122 (O_1122,N_19538,N_17141);
xor UO_1123 (O_1123,N_17153,N_19598);
nand UO_1124 (O_1124,N_19239,N_19337);
or UO_1125 (O_1125,N_18540,N_19294);
and UO_1126 (O_1126,N_18567,N_16310);
or UO_1127 (O_1127,N_16930,N_17272);
and UO_1128 (O_1128,N_18650,N_16230);
or UO_1129 (O_1129,N_19856,N_19793);
nor UO_1130 (O_1130,N_17017,N_17714);
and UO_1131 (O_1131,N_18329,N_18481);
or UO_1132 (O_1132,N_17194,N_19268);
nand UO_1133 (O_1133,N_18908,N_19738);
and UO_1134 (O_1134,N_17686,N_18343);
xnor UO_1135 (O_1135,N_18473,N_16548);
or UO_1136 (O_1136,N_18358,N_18892);
and UO_1137 (O_1137,N_16366,N_18989);
xor UO_1138 (O_1138,N_19024,N_19013);
or UO_1139 (O_1139,N_16565,N_18305);
or UO_1140 (O_1140,N_17335,N_18391);
nand UO_1141 (O_1141,N_17774,N_16766);
xnor UO_1142 (O_1142,N_18460,N_16982);
nand UO_1143 (O_1143,N_19361,N_19448);
xor UO_1144 (O_1144,N_19804,N_19531);
or UO_1145 (O_1145,N_19344,N_16303);
or UO_1146 (O_1146,N_16784,N_16781);
nand UO_1147 (O_1147,N_17989,N_17787);
or UO_1148 (O_1148,N_19041,N_19861);
nor UO_1149 (O_1149,N_16099,N_16333);
or UO_1150 (O_1150,N_17333,N_19580);
nand UO_1151 (O_1151,N_18017,N_17920);
and UO_1152 (O_1152,N_19889,N_17949);
and UO_1153 (O_1153,N_17769,N_17960);
nand UO_1154 (O_1154,N_18015,N_16747);
nor UO_1155 (O_1155,N_19163,N_16307);
xor UO_1156 (O_1156,N_16653,N_17267);
nor UO_1157 (O_1157,N_16164,N_18323);
xnor UO_1158 (O_1158,N_19398,N_17210);
nor UO_1159 (O_1159,N_16455,N_18389);
and UO_1160 (O_1160,N_19335,N_18879);
xnor UO_1161 (O_1161,N_17180,N_18933);
nor UO_1162 (O_1162,N_19854,N_18314);
and UO_1163 (O_1163,N_19112,N_18467);
or UO_1164 (O_1164,N_16969,N_17111);
nor UO_1165 (O_1165,N_17505,N_19555);
nand UO_1166 (O_1166,N_18126,N_19182);
xor UO_1167 (O_1167,N_18902,N_19895);
nand UO_1168 (O_1168,N_19663,N_19036);
xnor UO_1169 (O_1169,N_18916,N_18934);
or UO_1170 (O_1170,N_18218,N_16391);
xnor UO_1171 (O_1171,N_17782,N_17626);
nand UO_1172 (O_1172,N_17609,N_16772);
xor UO_1173 (O_1173,N_19907,N_16779);
nor UO_1174 (O_1174,N_16704,N_16135);
xnor UO_1175 (O_1175,N_19863,N_19009);
nor UO_1176 (O_1176,N_16356,N_17612);
or UO_1177 (O_1177,N_17799,N_18259);
and UO_1178 (O_1178,N_17768,N_16875);
nand UO_1179 (O_1179,N_19944,N_17520);
or UO_1180 (O_1180,N_18668,N_16229);
and UO_1181 (O_1181,N_19945,N_19867);
or UO_1182 (O_1182,N_17373,N_16918);
nor UO_1183 (O_1183,N_17955,N_19236);
and UO_1184 (O_1184,N_16686,N_18442);
nand UO_1185 (O_1185,N_19045,N_16571);
nand UO_1186 (O_1186,N_19198,N_17247);
xnor UO_1187 (O_1187,N_16834,N_16794);
or UO_1188 (O_1188,N_17758,N_16428);
nand UO_1189 (O_1189,N_18943,N_16131);
or UO_1190 (O_1190,N_19062,N_18300);
or UO_1191 (O_1191,N_17055,N_18102);
or UO_1192 (O_1192,N_16919,N_19396);
nand UO_1193 (O_1193,N_19052,N_18845);
nor UO_1194 (O_1194,N_17514,N_16670);
xor UO_1195 (O_1195,N_16749,N_19189);
and UO_1196 (O_1196,N_18773,N_19082);
nand UO_1197 (O_1197,N_18187,N_16549);
nand UO_1198 (O_1198,N_19286,N_19387);
nor UO_1199 (O_1199,N_16066,N_18062);
nor UO_1200 (O_1200,N_18847,N_16315);
xor UO_1201 (O_1201,N_18429,N_16188);
or UO_1202 (O_1202,N_16792,N_19027);
nor UO_1203 (O_1203,N_19603,N_19641);
nand UO_1204 (O_1204,N_17878,N_18118);
nand UO_1205 (O_1205,N_17585,N_19174);
and UO_1206 (O_1206,N_18699,N_17738);
nor UO_1207 (O_1207,N_16342,N_19147);
or UO_1208 (O_1208,N_17099,N_18996);
or UO_1209 (O_1209,N_16451,N_16256);
nand UO_1210 (O_1210,N_19015,N_16185);
xnor UO_1211 (O_1211,N_19020,N_18147);
or UO_1212 (O_1212,N_17911,N_17689);
and UO_1213 (O_1213,N_18324,N_18111);
nand UO_1214 (O_1214,N_16545,N_17809);
nor UO_1215 (O_1215,N_19518,N_18747);
nand UO_1216 (O_1216,N_16649,N_16703);
nor UO_1217 (O_1217,N_16328,N_16039);
and UO_1218 (O_1218,N_16780,N_16443);
xor UO_1219 (O_1219,N_18070,N_17578);
xnor UO_1220 (O_1220,N_16034,N_19359);
and UO_1221 (O_1221,N_16242,N_18723);
nand UO_1222 (O_1222,N_17557,N_18678);
and UO_1223 (O_1223,N_18941,N_19972);
nor UO_1224 (O_1224,N_17754,N_17852);
and UO_1225 (O_1225,N_16899,N_19390);
and UO_1226 (O_1226,N_18175,N_18726);
and UO_1227 (O_1227,N_19552,N_19546);
and UO_1228 (O_1228,N_16868,N_16863);
and UO_1229 (O_1229,N_18982,N_17914);
xnor UO_1230 (O_1230,N_16959,N_17429);
xnor UO_1231 (O_1231,N_18806,N_16000);
xor UO_1232 (O_1232,N_16681,N_18201);
nor UO_1233 (O_1233,N_17858,N_19025);
and UO_1234 (O_1234,N_16867,N_18887);
nor UO_1235 (O_1235,N_16182,N_17146);
or UO_1236 (O_1236,N_19334,N_19734);
xnor UO_1237 (O_1237,N_19706,N_18631);
and UO_1238 (O_1238,N_16155,N_18645);
and UO_1239 (O_1239,N_16106,N_16414);
nand UO_1240 (O_1240,N_18464,N_18081);
nor UO_1241 (O_1241,N_18471,N_18915);
nor UO_1242 (O_1242,N_16974,N_18341);
or UO_1243 (O_1243,N_17405,N_17463);
xnor UO_1244 (O_1244,N_17340,N_19624);
nor UO_1245 (O_1245,N_17068,N_17259);
or UO_1246 (O_1246,N_17401,N_16620);
xnor UO_1247 (O_1247,N_17986,N_16069);
or UO_1248 (O_1248,N_17724,N_16639);
nand UO_1249 (O_1249,N_19662,N_19284);
or UO_1250 (O_1250,N_16454,N_18764);
nor UO_1251 (O_1251,N_19825,N_18881);
or UO_1252 (O_1252,N_17456,N_16474);
nand UO_1253 (O_1253,N_19270,N_19217);
nor UO_1254 (O_1254,N_17435,N_18888);
nand UO_1255 (O_1255,N_19377,N_16987);
nor UO_1256 (O_1256,N_18333,N_19939);
and UO_1257 (O_1257,N_18810,N_19628);
xor UO_1258 (O_1258,N_17916,N_18282);
nand UO_1259 (O_1259,N_17579,N_18447);
and UO_1260 (O_1260,N_17151,N_17009);
nor UO_1261 (O_1261,N_19440,N_19932);
nand UO_1262 (O_1262,N_18949,N_17200);
and UO_1263 (O_1263,N_17601,N_17195);
or UO_1264 (O_1264,N_17839,N_19113);
nand UO_1265 (O_1265,N_17022,N_18357);
nand UO_1266 (O_1266,N_18724,N_18456);
xor UO_1267 (O_1267,N_17701,N_19742);
xor UO_1268 (O_1268,N_16958,N_16480);
nand UO_1269 (O_1269,N_18434,N_19685);
nor UO_1270 (O_1270,N_18360,N_17693);
nor UO_1271 (O_1271,N_16693,N_19485);
nor UO_1272 (O_1272,N_16507,N_18152);
or UO_1273 (O_1273,N_17976,N_17540);
nor UO_1274 (O_1274,N_16851,N_17152);
nor UO_1275 (O_1275,N_16423,N_18939);
nand UO_1276 (O_1276,N_17364,N_17821);
xor UO_1277 (O_1277,N_18233,N_16380);
nand UO_1278 (O_1278,N_16278,N_16692);
nor UO_1279 (O_1279,N_17736,N_19584);
and UO_1280 (O_1280,N_18063,N_17148);
or UO_1281 (O_1281,N_16505,N_19438);
xor UO_1282 (O_1282,N_16477,N_19340);
or UO_1283 (O_1283,N_17175,N_16555);
or UO_1284 (O_1284,N_17646,N_18037);
nor UO_1285 (O_1285,N_17963,N_18470);
xnor UO_1286 (O_1286,N_19958,N_19355);
nand UO_1287 (O_1287,N_17750,N_17604);
nor UO_1288 (O_1288,N_16732,N_16879);
nand UO_1289 (O_1289,N_16208,N_16890);
nor UO_1290 (O_1290,N_18327,N_18205);
nor UO_1291 (O_1291,N_16181,N_18000);
nand UO_1292 (O_1292,N_19874,N_16183);
nor UO_1293 (O_1293,N_19264,N_18347);
or UO_1294 (O_1294,N_16116,N_16468);
nor UO_1295 (O_1295,N_18621,N_18034);
nand UO_1296 (O_1296,N_19322,N_18543);
nor UO_1297 (O_1297,N_19632,N_19983);
xor UO_1298 (O_1298,N_17083,N_17441);
and UO_1299 (O_1299,N_18544,N_17209);
xor UO_1300 (O_1300,N_16096,N_18948);
nand UO_1301 (O_1301,N_19787,N_18656);
and UO_1302 (O_1302,N_19754,N_16218);
or UO_1303 (O_1303,N_17876,N_17397);
xor UO_1304 (O_1304,N_18655,N_19627);
nand UO_1305 (O_1305,N_19373,N_16902);
xnor UO_1306 (O_1306,N_18332,N_16228);
nand UO_1307 (O_1307,N_19227,N_16663);
and UO_1308 (O_1308,N_18249,N_16544);
or UO_1309 (O_1309,N_17600,N_16752);
or UO_1310 (O_1310,N_16332,N_16528);
and UO_1311 (O_1311,N_18248,N_19702);
nand UO_1312 (O_1312,N_19145,N_16805);
or UO_1313 (O_1313,N_17346,N_17497);
nand UO_1314 (O_1314,N_17991,N_17430);
and UO_1315 (O_1315,N_19443,N_17054);
xnor UO_1316 (O_1316,N_18545,N_16882);
and UO_1317 (O_1317,N_16856,N_18185);
nand UO_1318 (O_1318,N_17748,N_17064);
or UO_1319 (O_1319,N_17417,N_18976);
xor UO_1320 (O_1320,N_18274,N_18003);
or UO_1321 (O_1321,N_19279,N_16607);
nand UO_1322 (O_1322,N_17650,N_17387);
xor UO_1323 (O_1323,N_17506,N_17102);
nor UO_1324 (O_1324,N_19477,N_17569);
and UO_1325 (O_1325,N_18643,N_19017);
or UO_1326 (O_1326,N_16296,N_17814);
xnor UO_1327 (O_1327,N_19406,N_18519);
xor UO_1328 (O_1328,N_16631,N_16441);
or UO_1329 (O_1329,N_17170,N_19465);
and UO_1330 (O_1330,N_18247,N_19998);
nand UO_1331 (O_1331,N_19054,N_19875);
and UO_1332 (O_1332,N_18759,N_16062);
xor UO_1333 (O_1333,N_16770,N_17925);
nor UO_1334 (O_1334,N_16151,N_19721);
or UO_1335 (O_1335,N_19576,N_19660);
nor UO_1336 (O_1336,N_16522,N_19871);
nand UO_1337 (O_1337,N_18640,N_16647);
xnor UO_1338 (O_1338,N_16904,N_18437);
or UO_1339 (O_1339,N_18495,N_19653);
or UO_1340 (O_1340,N_18988,N_19432);
nor UO_1341 (O_1341,N_17943,N_16602);
xnor UO_1342 (O_1342,N_18925,N_16023);
nor UO_1343 (O_1343,N_17635,N_16210);
or UO_1344 (O_1344,N_16376,N_18967);
and UO_1345 (O_1345,N_19468,N_18352);
nor UO_1346 (O_1346,N_19788,N_18174);
nor UO_1347 (O_1347,N_18876,N_16700);
and UO_1348 (O_1348,N_17826,N_19482);
and UO_1349 (O_1349,N_17619,N_17112);
nor UO_1350 (O_1350,N_18859,N_18375);
nand UO_1351 (O_1351,N_17731,N_17840);
or UO_1352 (O_1352,N_16147,N_18629);
nor UO_1353 (O_1353,N_18591,N_16309);
and UO_1354 (O_1354,N_17795,N_17034);
or UO_1355 (O_1355,N_19575,N_18299);
nor UO_1356 (O_1356,N_17229,N_18478);
nor UO_1357 (O_1357,N_16629,N_17662);
nor UO_1358 (O_1358,N_18556,N_19880);
and UO_1359 (O_1359,N_18993,N_18346);
nand UO_1360 (O_1360,N_19621,N_19454);
nand UO_1361 (O_1361,N_17379,N_19652);
xnor UO_1362 (O_1362,N_17341,N_19119);
and UO_1363 (O_1363,N_17958,N_19929);
nor UO_1364 (O_1364,N_18355,N_17670);
xor UO_1365 (O_1365,N_16713,N_19620);
xnor UO_1366 (O_1366,N_17948,N_16580);
nand UO_1367 (O_1367,N_16668,N_19961);
or UO_1368 (O_1368,N_18756,N_17174);
nand UO_1369 (O_1369,N_16717,N_16724);
and UO_1370 (O_1370,N_17741,N_19725);
xnor UO_1371 (O_1371,N_17104,N_18821);
nand UO_1372 (O_1372,N_17278,N_18595);
or UO_1373 (O_1373,N_18666,N_17961);
nand UO_1374 (O_1374,N_18510,N_19304);
nor UO_1375 (O_1375,N_19539,N_17728);
and UO_1376 (O_1376,N_16409,N_17524);
nand UO_1377 (O_1377,N_19209,N_17120);
xor UO_1378 (O_1378,N_17515,N_18774);
xnor UO_1379 (O_1379,N_18288,N_17100);
nand UO_1380 (O_1380,N_18377,N_19481);
nand UO_1381 (O_1381,N_16314,N_16465);
or UO_1382 (O_1382,N_18870,N_19544);
xnor UO_1383 (O_1383,N_19818,N_19247);
xnor UO_1384 (O_1384,N_17479,N_18977);
xor UO_1385 (O_1385,N_18652,N_18728);
xor UO_1386 (O_1386,N_19912,N_16795);
nor UO_1387 (O_1387,N_16326,N_18171);
xor UO_1388 (O_1388,N_18030,N_18709);
and UO_1389 (O_1389,N_17119,N_17039);
or UO_1390 (O_1390,N_18117,N_18488);
and UO_1391 (O_1391,N_18393,N_18703);
and UO_1392 (O_1392,N_19059,N_19965);
nand UO_1393 (O_1393,N_17657,N_19611);
nand UO_1394 (O_1394,N_19931,N_17413);
xor UO_1395 (O_1395,N_16929,N_18420);
nand UO_1396 (O_1396,N_17002,N_16675);
and UO_1397 (O_1397,N_19565,N_17676);
nor UO_1398 (O_1398,N_17517,N_18968);
or UO_1399 (O_1399,N_19794,N_18149);
xnor UO_1400 (O_1400,N_19402,N_18842);
nand UO_1401 (O_1401,N_17453,N_16527);
nor UO_1402 (O_1402,N_16635,N_16961);
or UO_1403 (O_1403,N_16117,N_17937);
xor UO_1404 (O_1404,N_19033,N_19769);
xnor UO_1405 (O_1405,N_18020,N_19346);
nand UO_1406 (O_1406,N_17896,N_16172);
nor UO_1407 (O_1407,N_17289,N_19735);
or UO_1408 (O_1408,N_17187,N_16561);
and UO_1409 (O_1409,N_18255,N_16297);
or UO_1410 (O_1410,N_17098,N_17498);
xor UO_1411 (O_1411,N_19802,N_16568);
nor UO_1412 (O_1412,N_18361,N_19462);
xnor UO_1413 (O_1413,N_19303,N_16158);
nand UO_1414 (O_1414,N_18344,N_19253);
nor UO_1415 (O_1415,N_16291,N_19994);
nor UO_1416 (O_1416,N_18829,N_16453);
nand UO_1417 (O_1417,N_16822,N_19693);
and UO_1418 (O_1418,N_17642,N_19561);
or UO_1419 (O_1419,N_16860,N_17298);
xor UO_1420 (O_1420,N_19051,N_18956);
and UO_1421 (O_1421,N_18791,N_16082);
nor UO_1422 (O_1422,N_17789,N_18236);
nand UO_1423 (O_1423,N_19866,N_16848);
and UO_1424 (O_1424,N_19378,N_19315);
nand UO_1425 (O_1425,N_19828,N_19233);
or UO_1426 (O_1426,N_17849,N_16920);
nor UO_1427 (O_1427,N_16854,N_18552);
and UO_1428 (O_1428,N_16529,N_16450);
xor UO_1429 (O_1429,N_17028,N_17644);
and UO_1430 (O_1430,N_16729,N_19388);
xor UO_1431 (O_1431,N_19297,N_19207);
nand UO_1432 (O_1432,N_18168,N_16457);
or UO_1433 (O_1433,N_17007,N_18657);
and UO_1434 (O_1434,N_18830,N_16200);
nor UO_1435 (O_1435,N_17349,N_19282);
nor UO_1436 (O_1436,N_18455,N_17665);
nor UO_1437 (O_1437,N_18469,N_16207);
nor UO_1438 (O_1438,N_17951,N_19942);
xnor UO_1439 (O_1439,N_19499,N_18166);
nand UO_1440 (O_1440,N_19299,N_16235);
nand UO_1441 (O_1441,N_18238,N_17283);
nor UO_1442 (O_1442,N_16180,N_19415);
xnor UO_1443 (O_1443,N_18581,N_19938);
and UO_1444 (O_1444,N_18778,N_17356);
or UO_1445 (O_1445,N_19356,N_17794);
xnor UO_1446 (O_1446,N_19073,N_17086);
or UO_1447 (O_1447,N_16572,N_16213);
and UO_1448 (O_1448,N_19328,N_16424);
nor UO_1449 (O_1449,N_19845,N_18986);
and UO_1450 (O_1450,N_16835,N_19605);
or UO_1451 (O_1451,N_16855,N_17221);
nor UO_1452 (O_1452,N_16673,N_16880);
or UO_1453 (O_1453,N_18194,N_19962);
xnor UO_1454 (O_1454,N_16796,N_17322);
or UO_1455 (O_1455,N_18225,N_18863);
and UO_1456 (O_1456,N_17482,N_18090);
nor UO_1457 (O_1457,N_17841,N_16618);
nor UO_1458 (O_1458,N_17652,N_17292);
xor UO_1459 (O_1459,N_18909,N_18350);
or UO_1460 (O_1460,N_16481,N_19595);
or UO_1461 (O_1461,N_16652,N_17462);
and UO_1462 (O_1462,N_17129,N_17234);
xor UO_1463 (O_1463,N_16934,N_19796);
nor UO_1464 (O_1464,N_16091,N_16715);
or UO_1465 (O_1465,N_17434,N_18749);
or UO_1466 (O_1466,N_16981,N_19655);
nand UO_1467 (O_1467,N_19589,N_18142);
or UO_1468 (O_1468,N_19876,N_19855);
and UO_1469 (O_1469,N_18476,N_18278);
and UO_1470 (O_1470,N_18370,N_17072);
nand UO_1471 (O_1471,N_17414,N_19148);
nand UO_1472 (O_1472,N_18853,N_19908);
nand UO_1473 (O_1473,N_19811,N_17995);
or UO_1474 (O_1474,N_18516,N_17016);
or UO_1475 (O_1475,N_18109,N_17145);
and UO_1476 (O_1476,N_16280,N_19018);
or UO_1477 (O_1477,N_19783,N_19850);
xnor UO_1478 (O_1478,N_19558,N_17061);
and UO_1479 (O_1479,N_17188,N_18912);
nand UO_1480 (O_1480,N_17936,N_18862);
nand UO_1481 (O_1481,N_19187,N_17237);
nor UO_1482 (O_1482,N_16176,N_17640);
nand UO_1483 (O_1483,N_19583,N_19243);
or UO_1484 (O_1484,N_19458,N_17556);
and UO_1485 (O_1485,N_18297,N_17110);
or UO_1486 (O_1486,N_16419,N_18116);
and UO_1487 (O_1487,N_18719,N_17363);
and UO_1488 (O_1488,N_17386,N_19004);
or UO_1489 (O_1489,N_19533,N_17851);
or UO_1490 (O_1490,N_16170,N_19594);
nand UO_1491 (O_1491,N_18971,N_18511);
and UO_1492 (O_1492,N_17760,N_16221);
and UO_1493 (O_1493,N_19862,N_16086);
xor UO_1494 (O_1494,N_16985,N_18303);
and UO_1495 (O_1495,N_17495,N_17085);
xor UO_1496 (O_1496,N_18254,N_17654);
or UO_1497 (O_1497,N_16354,N_16643);
or UO_1498 (O_1498,N_17084,N_17580);
and UO_1499 (O_1499,N_16044,N_19508);
and UO_1500 (O_1500,N_16492,N_19351);
nand UO_1501 (O_1501,N_19178,N_17688);
nand UO_1502 (O_1502,N_16058,N_16104);
xnor UO_1503 (O_1503,N_16723,N_17651);
nor UO_1504 (O_1504,N_17918,N_16591);
nand UO_1505 (O_1505,N_17303,N_18284);
nand UO_1506 (O_1506,N_19484,N_18128);
nor UO_1507 (O_1507,N_16952,N_17275);
xor UO_1508 (O_1508,N_16159,N_17880);
and UO_1509 (O_1509,N_18807,N_18675);
xnor UO_1510 (O_1510,N_16501,N_18894);
or UO_1511 (O_1511,N_17330,N_16625);
xnor UO_1512 (O_1512,N_16667,N_19917);
and UO_1513 (O_1513,N_19404,N_16998);
and UO_1514 (O_1514,N_19921,N_19320);
nor UO_1515 (O_1515,N_17558,N_17608);
or UO_1516 (O_1516,N_18669,N_19722);
nand UO_1517 (O_1517,N_17242,N_16654);
nand UO_1518 (O_1518,N_19606,N_18683);
and UO_1519 (O_1519,N_17354,N_18342);
or UO_1520 (O_1520,N_19957,N_18400);
or UO_1521 (O_1521,N_19211,N_17353);
or UO_1522 (O_1522,N_17710,N_19205);
nor UO_1523 (O_1523,N_19935,N_19070);
xnor UO_1524 (O_1524,N_18223,N_18642);
and UO_1525 (O_1525,N_19661,N_16255);
nor UO_1526 (O_1526,N_18013,N_16336);
or UO_1527 (O_1527,N_19671,N_19104);
nor UO_1528 (O_1528,N_19947,N_18229);
xnor UO_1529 (O_1529,N_19030,N_16581);
nor UO_1530 (O_1530,N_17197,N_17361);
or UO_1531 (O_1531,N_19941,N_18232);
xor UO_1532 (O_1532,N_19192,N_17996);
nand UO_1533 (O_1533,N_16312,N_18580);
or UO_1534 (O_1534,N_17700,N_19002);
xnor UO_1535 (O_1535,N_19436,N_17935);
or UO_1536 (O_1536,N_16160,N_17196);
nand UO_1537 (O_1537,N_16975,N_19435);
nor UO_1538 (O_1538,N_19258,N_16190);
nor UO_1539 (O_1539,N_16705,N_17907);
xor UO_1540 (O_1540,N_17674,N_19071);
and UO_1541 (O_1541,N_18368,N_16144);
xor UO_1542 (O_1542,N_18823,N_17567);
nand UO_1543 (O_1543,N_18790,N_16081);
and UO_1544 (O_1544,N_19878,N_19781);
nor UO_1545 (O_1545,N_16215,N_18794);
nor UO_1546 (O_1546,N_19474,N_16438);
or UO_1547 (O_1547,N_17755,N_17752);
nor UO_1548 (O_1548,N_16515,N_16469);
nand UO_1549 (O_1549,N_18671,N_17076);
xor UO_1550 (O_1550,N_16270,N_19272);
xor UO_1551 (O_1551,N_17990,N_19101);
nor UO_1552 (O_1552,N_19870,N_19110);
or UO_1553 (O_1553,N_16363,N_17370);
or UO_1554 (O_1554,N_17698,N_17404);
and UO_1555 (O_1555,N_16983,N_16537);
or UO_1556 (O_1556,N_17134,N_19894);
nand UO_1557 (O_1557,N_18787,N_19248);
or UO_1558 (O_1558,N_19064,N_17984);
xnor UO_1559 (O_1559,N_17092,N_17971);
nor UO_1560 (O_1560,N_19639,N_16844);
or UO_1561 (O_1561,N_16721,N_19974);
xnor UO_1562 (O_1562,N_18189,N_18271);
nand UO_1563 (O_1563,N_16496,N_16262);
nand UO_1564 (O_1564,N_19137,N_17097);
nor UO_1565 (O_1565,N_19035,N_17847);
or UO_1566 (O_1566,N_18010,N_18445);
and UO_1567 (O_1567,N_18983,N_17032);
nand UO_1568 (O_1568,N_19971,N_18002);
nor UO_1569 (O_1569,N_19235,N_18216);
and UO_1570 (O_1570,N_16405,N_18537);
nand UO_1571 (O_1571,N_16422,N_19986);
and UO_1572 (O_1572,N_17680,N_16043);
nand UO_1573 (O_1573,N_16253,N_16119);
and UO_1574 (O_1574,N_19298,N_16874);
or UO_1575 (O_1575,N_18698,N_17478);
nand UO_1576 (O_1576,N_16967,N_19010);
or UO_1577 (O_1577,N_19428,N_19502);
nand UO_1578 (O_1578,N_16393,N_18950);
or UO_1579 (O_1579,N_17293,N_18819);
or UO_1580 (O_1580,N_18291,N_16324);
or UO_1581 (O_1581,N_16383,N_16040);
and UO_1582 (O_1582,N_16243,N_16169);
nand UO_1583 (O_1583,N_18449,N_17347);
nand UO_1584 (O_1584,N_19447,N_17140);
xnor UO_1585 (O_1585,N_16849,N_19669);
nand UO_1586 (O_1586,N_19707,N_19785);
or UO_1587 (O_1587,N_18536,N_19708);
xnor UO_1588 (O_1588,N_17444,N_19566);
nand UO_1589 (O_1589,N_19370,N_16523);
or UO_1590 (O_1590,N_17933,N_17212);
and UO_1591 (O_1591,N_16344,N_18761);
or UO_1592 (O_1592,N_16753,N_17428);
or UO_1593 (O_1593,N_16487,N_18452);
nand UO_1594 (O_1594,N_18648,N_16829);
nor UO_1595 (O_1595,N_17733,N_19869);
nand UO_1596 (O_1596,N_19309,N_18410);
nor UO_1597 (O_1597,N_17715,N_18479);
nor UO_1598 (O_1598,N_19571,N_19995);
nor UO_1599 (O_1599,N_18582,N_18441);
nor UO_1600 (O_1600,N_17966,N_18196);
nand UO_1601 (O_1601,N_19892,N_19460);
xor UO_1602 (O_1602,N_19418,N_19419);
xor UO_1603 (O_1603,N_17422,N_17892);
or UO_1604 (O_1604,N_17702,N_18024);
nor UO_1605 (O_1605,N_17947,N_19281);
nand UO_1606 (O_1606,N_18799,N_18849);
and UO_1607 (O_1607,N_16271,N_17360);
nand UO_1608 (O_1608,N_18046,N_17325);
nor UO_1609 (O_1609,N_18865,N_18009);
nor UO_1610 (O_1610,N_19820,N_18279);
nor UO_1611 (O_1611,N_18835,N_19364);
and UO_1612 (O_1612,N_19642,N_16251);
or UO_1613 (O_1613,N_18404,N_17490);
and UO_1614 (O_1614,N_16134,N_18768);
nand UO_1615 (O_1615,N_16727,N_16790);
nand UO_1616 (O_1616,N_19658,N_16259);
and UO_1617 (O_1617,N_18120,N_18180);
and UO_1618 (O_1618,N_16264,N_19069);
or UO_1619 (O_1619,N_19755,N_18047);
or UO_1620 (O_1620,N_18725,N_18878);
xnor UO_1621 (O_1621,N_17869,N_18444);
or UO_1622 (O_1622,N_16886,N_17703);
or UO_1623 (O_1623,N_17013,N_19836);
or UO_1624 (O_1624,N_18411,N_16202);
nor UO_1625 (O_1625,N_19157,N_18397);
nor UO_1626 (O_1626,N_18584,N_17077);
xnor UO_1627 (O_1627,N_18412,N_16716);
nand UO_1628 (O_1628,N_18359,N_16524);
nor UO_1629 (O_1629,N_16694,N_19585);
and UO_1630 (O_1630,N_16272,N_18417);
xor UO_1631 (O_1631,N_18054,N_16588);
or UO_1632 (O_1632,N_16288,N_16148);
nor UO_1633 (O_1633,N_16813,N_19422);
xor UO_1634 (O_1634,N_18786,N_19647);
nand UO_1635 (O_1635,N_17087,N_19976);
nand UO_1636 (O_1636,N_19949,N_17142);
nor UO_1637 (O_1637,N_19126,N_19559);
or UO_1638 (O_1638,N_19092,N_17973);
nand UO_1639 (O_1639,N_17173,N_19826);
nand UO_1640 (O_1640,N_17536,N_17695);
and UO_1641 (O_1641,N_18610,N_18947);
nor UO_1642 (O_1642,N_18178,N_19924);
or UO_1643 (O_1643,N_16869,N_18179);
or UO_1644 (O_1644,N_16478,N_18395);
xor UO_1645 (O_1645,N_19497,N_19090);
and UO_1646 (O_1646,N_17921,N_16960);
xor UO_1647 (O_1647,N_19581,N_17487);
nor UO_1648 (O_1648,N_19683,N_18505);
xor UO_1649 (O_1649,N_17252,N_19444);
or UO_1650 (O_1650,N_19469,N_19331);
and UO_1651 (O_1651,N_19637,N_16157);
nand UO_1652 (O_1652,N_17281,N_19913);
nor UO_1653 (O_1653,N_18590,N_19259);
xnor UO_1654 (O_1654,N_17900,N_19354);
and UO_1655 (O_1655,N_19450,N_18573);
nor UO_1656 (O_1656,N_16077,N_16910);
nor UO_1657 (O_1657,N_18515,N_19675);
and UO_1658 (O_1658,N_18946,N_17253);
and UO_1659 (O_1659,N_17875,N_16535);
or UO_1660 (O_1660,N_19597,N_17019);
or UO_1661 (O_1661,N_16022,N_19786);
or UO_1662 (O_1662,N_18964,N_19421);
nand UO_1663 (O_1663,N_19927,N_19564);
nand UO_1664 (O_1664,N_17525,N_18598);
and UO_1665 (O_1665,N_19830,N_17182);
nand UO_1666 (O_1666,N_18980,N_18005);
nor UO_1667 (O_1667,N_16881,N_16439);
or UO_1668 (O_1668,N_19835,N_17694);
nor UO_1669 (O_1669,N_18052,N_16812);
xnor UO_1670 (O_1670,N_16238,N_17653);
xnor UO_1671 (O_1671,N_19442,N_19120);
or UO_1672 (O_1672,N_19042,N_16941);
and UO_1673 (O_1673,N_16859,N_18541);
xor UO_1674 (O_1674,N_19079,N_16543);
nand UO_1675 (O_1675,N_19138,N_19254);
or UO_1676 (O_1676,N_18408,N_17351);
nor UO_1677 (O_1677,N_19586,N_16406);
nand UO_1678 (O_1678,N_18351,N_16195);
nand UO_1679 (O_1679,N_16482,N_17302);
nor UO_1680 (O_1680,N_18308,N_18836);
or UO_1681 (O_1681,N_18130,N_18049);
xnor UO_1682 (O_1682,N_18579,N_19075);
nor UO_1683 (O_1683,N_16012,N_19277);
xor UO_1684 (O_1684,N_18322,N_17529);
xor UO_1685 (O_1685,N_17060,N_19358);
or UO_1686 (O_1686,N_17477,N_16735);
xnor UO_1687 (O_1687,N_16382,N_17628);
or UO_1688 (O_1688,N_16433,N_17779);
nand UO_1689 (O_1689,N_19955,N_18599);
and UO_1690 (O_1690,N_17592,N_19409);
xor UO_1691 (O_1691,N_18486,N_19105);
nor UO_1692 (O_1692,N_17384,N_16138);
xnor UO_1693 (O_1693,N_17424,N_18292);
nand UO_1694 (O_1694,N_17377,N_16150);
nor UO_1695 (O_1695,N_16589,N_19173);
nand UO_1696 (O_1696,N_16275,N_17590);
and UO_1697 (O_1697,N_18785,N_17607);
or UO_1698 (O_1698,N_16098,N_18974);
xor UO_1699 (O_1699,N_16646,N_19475);
nand UO_1700 (O_1700,N_17956,N_19664);
nand UO_1701 (O_1701,N_19644,N_18353);
or UO_1702 (O_1702,N_16437,N_18356);
and UO_1703 (O_1703,N_18060,N_16754);
xor UO_1704 (O_1704,N_18349,N_18871);
or UO_1705 (O_1705,N_17587,N_18689);
nand UO_1706 (O_1706,N_19988,N_16655);
and UO_1707 (O_1707,N_17844,N_16798);
or UO_1708 (O_1708,N_16613,N_17532);
nor UO_1709 (O_1709,N_19446,N_16100);
xnor UO_1710 (O_1710,N_18172,N_18082);
xnor UO_1711 (O_1711,N_16056,N_18321);
nand UO_1712 (O_1712,N_19610,N_16558);
nand UO_1713 (O_1713,N_19068,N_17589);
or UO_1714 (O_1714,N_18345,N_19144);
nand UO_1715 (O_1715,N_16141,N_18258);
and UO_1716 (O_1716,N_17365,N_18380);
nand UO_1717 (O_1717,N_19803,N_17621);
or UO_1718 (O_1718,N_17126,N_17309);
or UO_1719 (O_1719,N_18240,N_19963);
nor UO_1720 (O_1720,N_18084,N_18514);
or UO_1721 (O_1721,N_17133,N_18792);
nand UO_1722 (O_1722,N_17276,N_17927);
nand UO_1723 (O_1723,N_16191,N_17593);
or UO_1724 (O_1724,N_19164,N_17979);
xor UO_1725 (O_1725,N_17261,N_19686);
nand UO_1726 (O_1726,N_18583,N_18627);
xor UO_1727 (O_1727,N_17675,N_17510);
nand UO_1728 (O_1728,N_17177,N_18890);
nor UO_1729 (O_1729,N_19879,N_16167);
nand UO_1730 (O_1730,N_17448,N_17315);
or UO_1731 (O_1731,N_16774,N_17454);
nand UO_1732 (O_1732,N_19037,N_19645);
and UO_1733 (O_1733,N_16566,N_16325);
nand UO_1734 (O_1734,N_16247,N_17994);
nor UO_1735 (O_1735,N_16334,N_19307);
or UO_1736 (O_1736,N_16888,N_19490);
or UO_1737 (O_1737,N_19634,N_19987);
nand UO_1738 (O_1738,N_18161,N_18697);
xor UO_1739 (O_1739,N_17647,N_18985);
nor UO_1740 (O_1740,N_16105,N_16584);
and UO_1741 (O_1741,N_17706,N_19311);
or UO_1742 (O_1742,N_17287,N_18527);
and UO_1743 (O_1743,N_16512,N_16630);
xnor UO_1744 (O_1744,N_16417,N_19433);
and UO_1745 (O_1745,N_16021,N_18256);
or UO_1746 (O_1746,N_16762,N_19726);
or UO_1747 (O_1747,N_16677,N_17241);
or UO_1748 (O_1748,N_19047,N_17721);
or UO_1749 (O_1749,N_16707,N_17305);
xor UO_1750 (O_1750,N_16718,N_19022);
nand UO_1751 (O_1751,N_18491,N_16891);
nor UO_1752 (O_1752,N_19453,N_18535);
and UO_1753 (O_1753,N_19674,N_17493);
nor UO_1754 (O_1754,N_19888,N_18508);
and UO_1755 (O_1755,N_18992,N_18659);
nand UO_1756 (O_1756,N_19467,N_16399);
nand UO_1757 (O_1757,N_18131,N_19868);
nor UO_1758 (O_1758,N_18431,N_18882);
and UO_1759 (O_1759,N_18762,N_18244);
or UO_1760 (O_1760,N_17285,N_17977);
nor UO_1761 (O_1761,N_18911,N_16979);
xnor UO_1762 (O_1762,N_17368,N_16946);
xnor UO_1763 (O_1763,N_19229,N_16731);
nand UO_1764 (O_1764,N_17667,N_19280);
xor UO_1765 (O_1765,N_17331,N_16640);
nor UO_1766 (O_1766,N_19763,N_18439);
and UO_1767 (O_1767,N_16102,N_18302);
nand UO_1768 (O_1768,N_17284,N_18548);
nor UO_1769 (O_1769,N_18007,N_18706);
xnor UO_1770 (O_1770,N_19310,N_16199);
xnor UO_1771 (O_1771,N_17321,N_18676);
xor UO_1772 (O_1772,N_16993,N_17616);
nand UO_1773 (O_1773,N_17224,N_19626);
and UO_1774 (O_1774,N_17819,N_18451);
nand UO_1775 (O_1775,N_18022,N_19720);
nand UO_1776 (O_1776,N_17168,N_19376);
and UO_1777 (O_1777,N_16814,N_18822);
or UO_1778 (O_1778,N_18336,N_19121);
nand UO_1779 (O_1779,N_18373,N_19130);
xor UO_1780 (O_1780,N_17639,N_19094);
nor UO_1781 (O_1781,N_19980,N_19817);
nand UO_1782 (O_1782,N_16421,N_17254);
xor UO_1783 (O_1783,N_18328,N_16804);
xnor UO_1784 (O_1784,N_19952,N_16820);
nand UO_1785 (O_1785,N_17378,N_18414);
nand UO_1786 (O_1786,N_16092,N_18217);
and UO_1787 (O_1787,N_18649,N_18539);
and UO_1788 (O_1788,N_17798,N_17818);
or UO_1789 (O_1789,N_18524,N_18928);
and UO_1790 (O_1790,N_18143,N_16047);
or UO_1791 (O_1791,N_18838,N_19978);
xor UO_1792 (O_1792,N_18574,N_17791);
or UO_1793 (O_1793,N_17690,N_18066);
and UO_1794 (O_1794,N_17489,N_17655);
and UO_1795 (O_1795,N_16432,N_16005);
nand UO_1796 (O_1796,N_19847,N_17239);
or UO_1797 (O_1797,N_17269,N_18594);
xor UO_1798 (O_1798,N_18716,N_18110);
xor UO_1799 (O_1799,N_19542,N_19940);
or UO_1800 (O_1800,N_16743,N_16687);
nor UO_1801 (O_1801,N_16906,N_19635);
or UO_1802 (O_1802,N_17832,N_19226);
or UO_1803 (O_1803,N_16504,N_18867);
nand UO_1804 (O_1804,N_16884,N_19528);
nand UO_1805 (O_1805,N_17257,N_18694);
xor UO_1806 (O_1806,N_17045,N_19154);
nand UO_1807 (O_1807,N_19728,N_17248);
and UO_1808 (O_1808,N_16853,N_19372);
xor UO_1809 (O_1809,N_19060,N_17282);
xor UO_1810 (O_1810,N_16035,N_19125);
nor UO_1811 (O_1811,N_17408,N_16636);
nor UO_1812 (O_1812,N_16080,N_17504);
and UO_1813 (O_1813,N_18042,N_18008);
xor UO_1814 (O_1814,N_19250,N_16126);
xor UO_1815 (O_1815,N_17000,N_18398);
nor UO_1816 (O_1816,N_18138,N_17526);
nor UO_1817 (O_1817,N_17094,N_16060);
or UO_1818 (O_1818,N_19165,N_16593);
nand UO_1819 (O_1819,N_17895,N_16337);
nand UO_1820 (O_1820,N_17163,N_16696);
nor UO_1821 (O_1821,N_16226,N_18891);
and UO_1822 (O_1822,N_19773,N_19510);
and UO_1823 (O_1823,N_16632,N_16773);
xnor UO_1824 (O_1824,N_17636,N_19210);
nor UO_1825 (O_1825,N_17451,N_16374);
xor UO_1826 (O_1826,N_16274,N_17136);
nor UO_1827 (O_1827,N_18576,N_19012);
nor UO_1828 (O_1828,N_19143,N_19001);
nand UO_1829 (O_1829,N_18780,N_16184);
or UO_1830 (O_1830,N_17046,N_18458);
and UO_1831 (O_1831,N_17004,N_16685);
nand UO_1832 (O_1832,N_16390,N_19466);
and UO_1833 (O_1833,N_19841,N_19271);
and UO_1834 (O_1834,N_16036,N_16746);
nor UO_1835 (O_1835,N_19964,N_16877);
nor UO_1836 (O_1836,N_18804,N_18122);
nand UO_1837 (O_1837,N_17543,N_19106);
or UO_1838 (O_1838,N_19777,N_19003);
nand UO_1839 (O_1839,N_17775,N_19234);
and UO_1840 (O_1840,N_17678,N_19357);
and UO_1841 (O_1841,N_17965,N_17213);
xnor UO_1842 (O_1842,N_18078,N_16563);
nand UO_1843 (O_1843,N_19424,N_16857);
nand UO_1844 (O_1844,N_17872,N_16932);
nor UO_1845 (O_1845,N_18828,N_16596);
nor UO_1846 (O_1846,N_19084,N_16688);
nor UO_1847 (O_1847,N_17244,N_19819);
nand UO_1848 (O_1848,N_19860,N_17648);
xor UO_1849 (O_1849,N_16101,N_18257);
nand UO_1850 (O_1850,N_16517,N_19289);
nor UO_1851 (O_1851,N_16557,N_19698);
nand UO_1852 (O_1852,N_19711,N_17050);
nor UO_1853 (O_1853,N_16917,N_19604);
and UO_1854 (O_1854,N_18606,N_16911);
nand UO_1855 (O_1855,N_19263,N_19522);
nand UO_1856 (O_1856,N_19511,N_19695);
nor UO_1857 (O_1857,N_18796,N_17753);
and UO_1858 (O_1858,N_19729,N_16722);
nor UO_1859 (O_1859,N_18834,N_19573);
and UO_1860 (O_1860,N_16265,N_18402);
and UO_1861 (O_1861,N_17672,N_19392);
nor UO_1862 (O_1862,N_19180,N_16049);
or UO_1863 (O_1863,N_16997,N_17812);
nand UO_1864 (O_1864,N_19367,N_16179);
and UO_1865 (O_1865,N_16547,N_16927);
nand UO_1866 (O_1866,N_18811,N_18625);
nand UO_1867 (O_1867,N_18844,N_18555);
nand UO_1868 (O_1868,N_19336,N_16783);
nand UO_1869 (O_1869,N_16608,N_17065);
and UO_1870 (O_1870,N_19659,N_16214);
or UO_1871 (O_1871,N_16222,N_18298);
and UO_1872 (O_1872,N_17108,N_16349);
nor UO_1873 (O_1873,N_18554,N_17232);
and UO_1874 (O_1874,N_18079,N_17011);
nor UO_1875 (O_1875,N_16973,N_16937);
xnor UO_1876 (O_1876,N_18067,N_16219);
nor UO_1877 (O_1877,N_18039,N_19016);
nor UO_1878 (O_1878,N_16436,N_19614);
xor UO_1879 (O_1879,N_19167,N_17725);
xor UO_1880 (O_1880,N_19665,N_19724);
or UO_1881 (O_1881,N_17231,N_16509);
and UO_1882 (O_1882,N_19813,N_18634);
or UO_1883 (O_1883,N_17661,N_16809);
or UO_1884 (O_1884,N_17027,N_17047);
or UO_1885 (O_1885,N_16531,N_16025);
or UO_1886 (O_1886,N_16240,N_19712);
xnor UO_1887 (O_1887,N_18817,N_16500);
and UO_1888 (O_1888,N_19249,N_18146);
and UO_1889 (O_1889,N_19551,N_17223);
and UO_1890 (O_1890,N_18740,N_17583);
xor UO_1891 (O_1891,N_19123,N_18235);
xnor UO_1892 (O_1892,N_18477,N_18815);
or UO_1893 (O_1893,N_19623,N_16616);
nor UO_1894 (O_1894,N_19219,N_17631);
xnor UO_1895 (O_1895,N_19353,N_17992);
or UO_1896 (O_1896,N_17597,N_16887);
xnor UO_1897 (O_1897,N_19953,N_17582);
or UO_1898 (O_1898,N_19260,N_16769);
xor UO_1899 (O_1899,N_18586,N_19703);
nand UO_1900 (O_1900,N_18043,N_19058);
or UO_1901 (O_1901,N_18107,N_18960);
nand UO_1902 (O_1902,N_17561,N_16063);
or UO_1903 (O_1903,N_16350,N_16648);
and UO_1904 (O_1904,N_18489,N_18418);
nor UO_1905 (O_1905,N_17946,N_19666);
xnor UO_1906 (O_1906,N_18632,N_16108);
and UO_1907 (O_1907,N_18075,N_16367);
and UO_1908 (O_1908,N_17550,N_16816);
xnor UO_1909 (O_1909,N_17037,N_17266);
nor UO_1910 (O_1910,N_17427,N_17893);
nand UO_1911 (O_1911,N_17785,N_19410);
nor UO_1912 (O_1912,N_19846,N_16538);
and UO_1913 (O_1913,N_17542,N_19088);
nor UO_1914 (O_1914,N_17191,N_17326);
xnor UO_1915 (O_1915,N_16459,N_17190);
and UO_1916 (O_1916,N_19911,N_17122);
nand UO_1917 (O_1917,N_17732,N_17228);
nand UO_1918 (O_1918,N_17528,N_16777);
xor UO_1919 (O_1919,N_16490,N_17312);
or UO_1920 (O_1920,N_17073,N_19267);
nand UO_1921 (O_1921,N_18286,N_18088);
or UO_1922 (O_1922,N_19200,N_18148);
xor UO_1923 (O_1923,N_18679,N_18905);
and UO_1924 (O_1924,N_19188,N_16111);
xnor UO_1925 (O_1925,N_16152,N_18673);
nor UO_1926 (O_1926,N_18221,N_19548);
xnor UO_1927 (O_1927,N_19731,N_18011);
nor UO_1928 (O_1928,N_18367,N_18855);
or UO_1929 (O_1929,N_17310,N_16768);
and UO_1930 (O_1930,N_19520,N_17507);
and UO_1931 (O_1931,N_16358,N_18383);
nand UO_1932 (O_1932,N_18639,N_19412);
xnor UO_1933 (O_1933,N_17089,N_17091);
or UO_1934 (O_1934,N_18769,N_18592);
or UO_1935 (O_1935,N_17862,N_16839);
and UO_1936 (O_1936,N_16674,N_18936);
xor UO_1937 (O_1937,N_18124,N_19812);
nand UO_1938 (O_1938,N_19926,N_17159);
or UO_1939 (O_1939,N_16871,N_19457);
or UO_1940 (O_1940,N_16070,N_17484);
nand UO_1941 (O_1941,N_17964,N_17455);
xnor UO_1942 (O_1942,N_19241,N_16042);
or UO_1943 (O_1943,N_19885,N_17235);
nand UO_1944 (O_1944,N_19768,N_18230);
nand UO_1945 (O_1945,N_19568,N_18071);
or UO_1946 (O_1946,N_16748,N_18296);
or UO_1947 (O_1947,N_16093,N_17865);
xor UO_1948 (O_1948,N_18136,N_19849);
xor UO_1949 (O_1949,N_16567,N_18243);
xnor UO_1950 (O_1950,N_18596,N_17249);
and UO_1951 (O_1951,N_18857,N_17006);
nor UO_1952 (O_1952,N_18145,N_18603);
xor UO_1953 (O_1953,N_18927,N_18981);
xnor UO_1954 (O_1954,N_19881,N_16833);
nor UO_1955 (O_1955,N_17366,N_16651);
and UO_1956 (O_1956,N_18730,N_18856);
and UO_1957 (O_1957,N_16594,N_19117);
or UO_1958 (O_1958,N_16599,N_18702);
nand UO_1959 (O_1959,N_16806,N_18158);
or UO_1960 (O_1960,N_17952,N_19108);
and UO_1961 (O_1961,N_17877,N_17627);
or UO_1962 (O_1962,N_16125,N_16090);
or UO_1963 (O_1963,N_18041,N_18824);
xnor UO_1964 (O_1964,N_16486,N_16574);
and UO_1965 (O_1965,N_19493,N_17486);
and UO_1966 (O_1966,N_19021,N_16977);
nand UO_1967 (O_1967,N_17299,N_19220);
nor UO_1968 (O_1968,N_18446,N_17075);
and UO_1969 (O_1969,N_16756,N_19408);
or UO_1970 (O_1970,N_17183,N_17088);
and UO_1971 (O_1971,N_19394,N_18851);
or UO_1972 (O_1972,N_17836,N_17230);
and UO_1973 (O_1973,N_16194,N_17201);
xnor UO_1974 (O_1974,N_18285,N_18825);
nand UO_1975 (O_1975,N_17218,N_18262);
xor UO_1976 (O_1976,N_17043,N_19996);
nor UO_1977 (O_1977,N_17398,N_18783);
and UO_1978 (O_1978,N_18399,N_16966);
and UO_1979 (O_1979,N_16810,N_16706);
and UO_1980 (O_1980,N_17158,N_18692);
nor UO_1981 (O_1981,N_17538,N_16847);
xor UO_1982 (O_1982,N_18386,N_18776);
and UO_1983 (O_1983,N_17749,N_16900);
xor UO_1984 (O_1984,N_16948,N_17114);
nand UO_1985 (O_1985,N_19142,N_16991);
xor UO_1986 (O_1986,N_17551,N_19612);
xor UO_1987 (O_1987,N_18628,N_19194);
xor UO_1988 (O_1988,N_19338,N_18924);
xnor UO_1989 (O_1989,N_16168,N_17440);
nor UO_1990 (O_1990,N_16897,N_19657);
nor UO_1991 (O_1991,N_16761,N_17762);
xor UO_1992 (O_1992,N_19251,N_16719);
or UO_1993 (O_1993,N_16939,N_18601);
or UO_1994 (O_1994,N_18623,N_17251);
and UO_1995 (O_1995,N_16744,N_16248);
nand UO_1996 (O_1996,N_19492,N_18585);
and UO_1997 (O_1997,N_16606,N_19023);
nor UO_1998 (O_1998,N_17474,N_18250);
xor UO_1999 (O_1999,N_16057,N_17327);
and UO_2000 (O_2000,N_16104,N_19974);
or UO_2001 (O_2001,N_18994,N_18337);
and UO_2002 (O_2002,N_17301,N_19142);
nor UO_2003 (O_2003,N_18476,N_18879);
nand UO_2004 (O_2004,N_16605,N_18251);
and UO_2005 (O_2005,N_17001,N_18213);
nor UO_2006 (O_2006,N_17472,N_17800);
and UO_2007 (O_2007,N_17213,N_16260);
nor UO_2008 (O_2008,N_17120,N_17636);
and UO_2009 (O_2009,N_16078,N_16125);
and UO_2010 (O_2010,N_19034,N_16219);
nor UO_2011 (O_2011,N_18059,N_19754);
nor UO_2012 (O_2012,N_18571,N_16646);
nand UO_2013 (O_2013,N_18627,N_16429);
nand UO_2014 (O_2014,N_16529,N_19045);
and UO_2015 (O_2015,N_19112,N_19156);
nor UO_2016 (O_2016,N_17467,N_16736);
nor UO_2017 (O_2017,N_17466,N_17703);
or UO_2018 (O_2018,N_19905,N_17082);
nor UO_2019 (O_2019,N_19532,N_18365);
xor UO_2020 (O_2020,N_18964,N_19347);
nand UO_2021 (O_2021,N_16561,N_16966);
or UO_2022 (O_2022,N_16345,N_16523);
nand UO_2023 (O_2023,N_18441,N_16487);
nand UO_2024 (O_2024,N_16147,N_17331);
nand UO_2025 (O_2025,N_17033,N_19323);
xnor UO_2026 (O_2026,N_19331,N_17642);
and UO_2027 (O_2027,N_17633,N_17610);
and UO_2028 (O_2028,N_18130,N_18859);
nand UO_2029 (O_2029,N_17079,N_18539);
or UO_2030 (O_2030,N_16678,N_17269);
and UO_2031 (O_2031,N_16341,N_16261);
xor UO_2032 (O_2032,N_16167,N_19375);
and UO_2033 (O_2033,N_17832,N_18643);
nand UO_2034 (O_2034,N_17745,N_19982);
nor UO_2035 (O_2035,N_19224,N_18194);
or UO_2036 (O_2036,N_17680,N_17985);
and UO_2037 (O_2037,N_16323,N_16976);
nor UO_2038 (O_2038,N_19223,N_17888);
or UO_2039 (O_2039,N_18935,N_19308);
or UO_2040 (O_2040,N_19202,N_19985);
nand UO_2041 (O_2041,N_19317,N_16581);
nand UO_2042 (O_2042,N_19384,N_17839);
or UO_2043 (O_2043,N_16043,N_18733);
nand UO_2044 (O_2044,N_16273,N_19496);
nor UO_2045 (O_2045,N_18692,N_19277);
nand UO_2046 (O_2046,N_17939,N_17078);
and UO_2047 (O_2047,N_17373,N_16507);
xnor UO_2048 (O_2048,N_16523,N_16508);
nor UO_2049 (O_2049,N_16425,N_19613);
nor UO_2050 (O_2050,N_18804,N_17583);
or UO_2051 (O_2051,N_16891,N_17629);
xor UO_2052 (O_2052,N_18962,N_18461);
xnor UO_2053 (O_2053,N_19306,N_18704);
nor UO_2054 (O_2054,N_18257,N_18223);
nor UO_2055 (O_2055,N_19692,N_16007);
nor UO_2056 (O_2056,N_17176,N_17393);
nand UO_2057 (O_2057,N_16628,N_16050);
nand UO_2058 (O_2058,N_17720,N_19336);
nor UO_2059 (O_2059,N_19472,N_18503);
xor UO_2060 (O_2060,N_16036,N_16303);
nor UO_2061 (O_2061,N_18877,N_17356);
nor UO_2062 (O_2062,N_16974,N_17306);
xor UO_2063 (O_2063,N_19108,N_16011);
xnor UO_2064 (O_2064,N_17369,N_17432);
or UO_2065 (O_2065,N_18362,N_19316);
nand UO_2066 (O_2066,N_16087,N_16831);
or UO_2067 (O_2067,N_17818,N_18645);
nor UO_2068 (O_2068,N_18836,N_17759);
and UO_2069 (O_2069,N_16611,N_16512);
nand UO_2070 (O_2070,N_18108,N_17733);
xor UO_2071 (O_2071,N_18093,N_16570);
and UO_2072 (O_2072,N_16538,N_18556);
xor UO_2073 (O_2073,N_19763,N_17624);
and UO_2074 (O_2074,N_19561,N_19173);
or UO_2075 (O_2075,N_17790,N_19533);
xor UO_2076 (O_2076,N_18437,N_19904);
or UO_2077 (O_2077,N_17620,N_16116);
nand UO_2078 (O_2078,N_17911,N_17001);
or UO_2079 (O_2079,N_16793,N_18127);
xor UO_2080 (O_2080,N_16083,N_19032);
and UO_2081 (O_2081,N_18305,N_18393);
and UO_2082 (O_2082,N_17755,N_19238);
nand UO_2083 (O_2083,N_16847,N_17057);
or UO_2084 (O_2084,N_18927,N_16384);
xnor UO_2085 (O_2085,N_17861,N_18895);
and UO_2086 (O_2086,N_18622,N_18435);
nand UO_2087 (O_2087,N_17450,N_16261);
nor UO_2088 (O_2088,N_17435,N_16869);
and UO_2089 (O_2089,N_16094,N_18188);
xor UO_2090 (O_2090,N_19933,N_16630);
xor UO_2091 (O_2091,N_16831,N_17309);
nand UO_2092 (O_2092,N_17308,N_17143);
nand UO_2093 (O_2093,N_16915,N_18562);
nand UO_2094 (O_2094,N_16054,N_16590);
nor UO_2095 (O_2095,N_17614,N_18277);
nor UO_2096 (O_2096,N_19865,N_18211);
or UO_2097 (O_2097,N_16261,N_17354);
nand UO_2098 (O_2098,N_18528,N_19578);
nand UO_2099 (O_2099,N_18359,N_18899);
and UO_2100 (O_2100,N_19850,N_18822);
and UO_2101 (O_2101,N_18462,N_16450);
nand UO_2102 (O_2102,N_16890,N_16604);
and UO_2103 (O_2103,N_19587,N_17279);
nand UO_2104 (O_2104,N_16728,N_18939);
and UO_2105 (O_2105,N_18941,N_17062);
xnor UO_2106 (O_2106,N_17978,N_18569);
and UO_2107 (O_2107,N_16216,N_19120);
xnor UO_2108 (O_2108,N_17333,N_16994);
nand UO_2109 (O_2109,N_18982,N_16659);
and UO_2110 (O_2110,N_16455,N_16887);
nand UO_2111 (O_2111,N_16796,N_16121);
and UO_2112 (O_2112,N_19626,N_19289);
and UO_2113 (O_2113,N_19341,N_16947);
nand UO_2114 (O_2114,N_16662,N_17218);
nor UO_2115 (O_2115,N_16895,N_17509);
nand UO_2116 (O_2116,N_17761,N_16761);
nor UO_2117 (O_2117,N_18630,N_19642);
nand UO_2118 (O_2118,N_17666,N_18901);
xnor UO_2119 (O_2119,N_17288,N_17599);
or UO_2120 (O_2120,N_19459,N_17660);
or UO_2121 (O_2121,N_18643,N_19154);
xor UO_2122 (O_2122,N_16951,N_18074);
xor UO_2123 (O_2123,N_17520,N_18493);
nor UO_2124 (O_2124,N_16192,N_18143);
or UO_2125 (O_2125,N_18465,N_17932);
nand UO_2126 (O_2126,N_16492,N_18429);
xor UO_2127 (O_2127,N_18961,N_17898);
nand UO_2128 (O_2128,N_18339,N_17571);
and UO_2129 (O_2129,N_16839,N_16458);
nor UO_2130 (O_2130,N_18969,N_16353);
or UO_2131 (O_2131,N_18271,N_19012);
or UO_2132 (O_2132,N_17061,N_17885);
and UO_2133 (O_2133,N_17984,N_17530);
xnor UO_2134 (O_2134,N_18160,N_16380);
nand UO_2135 (O_2135,N_19867,N_17735);
or UO_2136 (O_2136,N_18419,N_18085);
and UO_2137 (O_2137,N_19280,N_18354);
nor UO_2138 (O_2138,N_16294,N_17334);
nand UO_2139 (O_2139,N_18997,N_16960);
xnor UO_2140 (O_2140,N_16051,N_17645);
nor UO_2141 (O_2141,N_18575,N_16199);
and UO_2142 (O_2142,N_17246,N_16437);
and UO_2143 (O_2143,N_17931,N_18361);
and UO_2144 (O_2144,N_17688,N_18042);
and UO_2145 (O_2145,N_19359,N_17799);
nand UO_2146 (O_2146,N_16518,N_19789);
or UO_2147 (O_2147,N_19759,N_18220);
nor UO_2148 (O_2148,N_17751,N_16643);
and UO_2149 (O_2149,N_19921,N_16756);
xor UO_2150 (O_2150,N_16860,N_16132);
nand UO_2151 (O_2151,N_19238,N_16807);
nor UO_2152 (O_2152,N_18898,N_19399);
nand UO_2153 (O_2153,N_17610,N_18170);
nor UO_2154 (O_2154,N_17309,N_19256);
xor UO_2155 (O_2155,N_17819,N_19859);
nor UO_2156 (O_2156,N_19072,N_17879);
or UO_2157 (O_2157,N_16744,N_16152);
or UO_2158 (O_2158,N_18615,N_17433);
nor UO_2159 (O_2159,N_17129,N_19464);
xor UO_2160 (O_2160,N_19434,N_18863);
or UO_2161 (O_2161,N_17569,N_16785);
nand UO_2162 (O_2162,N_17621,N_18583);
and UO_2163 (O_2163,N_17870,N_19118);
and UO_2164 (O_2164,N_16894,N_19708);
xnor UO_2165 (O_2165,N_18585,N_17638);
xor UO_2166 (O_2166,N_17111,N_18427);
nor UO_2167 (O_2167,N_19842,N_18554);
xnor UO_2168 (O_2168,N_17736,N_18990);
nand UO_2169 (O_2169,N_17779,N_16274);
or UO_2170 (O_2170,N_18225,N_18667);
and UO_2171 (O_2171,N_19095,N_17694);
xor UO_2172 (O_2172,N_17060,N_19595);
or UO_2173 (O_2173,N_17729,N_18418);
or UO_2174 (O_2174,N_18570,N_19764);
nor UO_2175 (O_2175,N_18190,N_16299);
nand UO_2176 (O_2176,N_19968,N_17542);
xor UO_2177 (O_2177,N_17793,N_16800);
or UO_2178 (O_2178,N_19120,N_17861);
nand UO_2179 (O_2179,N_17716,N_18541);
xor UO_2180 (O_2180,N_18285,N_19719);
nand UO_2181 (O_2181,N_16110,N_18950);
xor UO_2182 (O_2182,N_17144,N_17520);
and UO_2183 (O_2183,N_16781,N_19888);
nand UO_2184 (O_2184,N_16171,N_18982);
nand UO_2185 (O_2185,N_17526,N_18180);
and UO_2186 (O_2186,N_16464,N_19742);
or UO_2187 (O_2187,N_17932,N_17949);
nor UO_2188 (O_2188,N_18823,N_17757);
nand UO_2189 (O_2189,N_17821,N_16751);
nor UO_2190 (O_2190,N_16120,N_19130);
nand UO_2191 (O_2191,N_16661,N_17841);
and UO_2192 (O_2192,N_17292,N_16501);
or UO_2193 (O_2193,N_18877,N_17206);
and UO_2194 (O_2194,N_19953,N_17732);
or UO_2195 (O_2195,N_19185,N_16751);
or UO_2196 (O_2196,N_17019,N_16349);
and UO_2197 (O_2197,N_16006,N_18373);
and UO_2198 (O_2198,N_16246,N_17709);
or UO_2199 (O_2199,N_18900,N_19349);
nor UO_2200 (O_2200,N_18826,N_18112);
nand UO_2201 (O_2201,N_18289,N_17774);
and UO_2202 (O_2202,N_16241,N_17843);
and UO_2203 (O_2203,N_16102,N_17139);
or UO_2204 (O_2204,N_17648,N_16745);
or UO_2205 (O_2205,N_17769,N_17440);
xnor UO_2206 (O_2206,N_19294,N_17840);
nor UO_2207 (O_2207,N_19590,N_17125);
and UO_2208 (O_2208,N_19585,N_18116);
or UO_2209 (O_2209,N_17603,N_18727);
or UO_2210 (O_2210,N_19120,N_19063);
nor UO_2211 (O_2211,N_18643,N_18376);
nor UO_2212 (O_2212,N_17524,N_19806);
or UO_2213 (O_2213,N_19087,N_19178);
and UO_2214 (O_2214,N_19445,N_18147);
or UO_2215 (O_2215,N_16657,N_19174);
and UO_2216 (O_2216,N_18601,N_19926);
xnor UO_2217 (O_2217,N_19633,N_16155);
or UO_2218 (O_2218,N_17877,N_19891);
nor UO_2219 (O_2219,N_17956,N_17036);
and UO_2220 (O_2220,N_17902,N_18233);
xor UO_2221 (O_2221,N_18586,N_16047);
and UO_2222 (O_2222,N_17640,N_18866);
nor UO_2223 (O_2223,N_17300,N_19480);
xnor UO_2224 (O_2224,N_19626,N_17319);
or UO_2225 (O_2225,N_19682,N_17865);
nand UO_2226 (O_2226,N_18165,N_19146);
or UO_2227 (O_2227,N_17191,N_19676);
xnor UO_2228 (O_2228,N_18111,N_17387);
or UO_2229 (O_2229,N_18337,N_19429);
or UO_2230 (O_2230,N_19150,N_19938);
and UO_2231 (O_2231,N_16067,N_19198);
and UO_2232 (O_2232,N_17040,N_18908);
nor UO_2233 (O_2233,N_18201,N_19096);
or UO_2234 (O_2234,N_17395,N_17596);
and UO_2235 (O_2235,N_19579,N_19602);
nand UO_2236 (O_2236,N_17954,N_19247);
or UO_2237 (O_2237,N_17416,N_16589);
nor UO_2238 (O_2238,N_17102,N_18058);
or UO_2239 (O_2239,N_18570,N_17008);
xnor UO_2240 (O_2240,N_17993,N_18577);
nand UO_2241 (O_2241,N_18092,N_18174);
xor UO_2242 (O_2242,N_17195,N_17679);
and UO_2243 (O_2243,N_16966,N_17811);
nand UO_2244 (O_2244,N_18572,N_16224);
nor UO_2245 (O_2245,N_16113,N_17078);
and UO_2246 (O_2246,N_18459,N_16187);
nor UO_2247 (O_2247,N_17389,N_17471);
xnor UO_2248 (O_2248,N_19138,N_18149);
and UO_2249 (O_2249,N_16708,N_18851);
xor UO_2250 (O_2250,N_16279,N_17998);
and UO_2251 (O_2251,N_17981,N_17662);
or UO_2252 (O_2252,N_19209,N_16406);
or UO_2253 (O_2253,N_18667,N_18538);
nor UO_2254 (O_2254,N_19221,N_17574);
and UO_2255 (O_2255,N_18279,N_18799);
nand UO_2256 (O_2256,N_16266,N_18333);
xnor UO_2257 (O_2257,N_19634,N_17149);
nor UO_2258 (O_2258,N_17160,N_16113);
nor UO_2259 (O_2259,N_17160,N_19367);
and UO_2260 (O_2260,N_18580,N_17657);
and UO_2261 (O_2261,N_19498,N_16509);
nor UO_2262 (O_2262,N_18618,N_17713);
xor UO_2263 (O_2263,N_16483,N_17403);
nand UO_2264 (O_2264,N_16676,N_16840);
or UO_2265 (O_2265,N_16195,N_16883);
nand UO_2266 (O_2266,N_19784,N_17981);
or UO_2267 (O_2267,N_16742,N_16012);
and UO_2268 (O_2268,N_19986,N_18041);
or UO_2269 (O_2269,N_18756,N_16264);
nor UO_2270 (O_2270,N_16521,N_19012);
and UO_2271 (O_2271,N_16964,N_17455);
or UO_2272 (O_2272,N_17945,N_18731);
xor UO_2273 (O_2273,N_17879,N_17347);
nand UO_2274 (O_2274,N_19663,N_17346);
or UO_2275 (O_2275,N_19474,N_16082);
and UO_2276 (O_2276,N_16565,N_16771);
or UO_2277 (O_2277,N_18148,N_18775);
nand UO_2278 (O_2278,N_17053,N_19127);
or UO_2279 (O_2279,N_16293,N_18905);
xnor UO_2280 (O_2280,N_16718,N_17898);
or UO_2281 (O_2281,N_19965,N_17719);
nor UO_2282 (O_2282,N_17612,N_19090);
and UO_2283 (O_2283,N_18503,N_16710);
and UO_2284 (O_2284,N_19028,N_19537);
nand UO_2285 (O_2285,N_17433,N_16882);
and UO_2286 (O_2286,N_19251,N_17581);
and UO_2287 (O_2287,N_18461,N_19191);
or UO_2288 (O_2288,N_19203,N_19409);
xnor UO_2289 (O_2289,N_19043,N_16676);
and UO_2290 (O_2290,N_16265,N_16490);
or UO_2291 (O_2291,N_19188,N_18307);
nand UO_2292 (O_2292,N_16640,N_19303);
and UO_2293 (O_2293,N_19828,N_17129);
nor UO_2294 (O_2294,N_19825,N_19002);
xor UO_2295 (O_2295,N_19469,N_18523);
nand UO_2296 (O_2296,N_19313,N_17261);
xnor UO_2297 (O_2297,N_19702,N_19796);
and UO_2298 (O_2298,N_18064,N_17850);
xor UO_2299 (O_2299,N_18972,N_19927);
or UO_2300 (O_2300,N_18447,N_17370);
xnor UO_2301 (O_2301,N_18848,N_18761);
nand UO_2302 (O_2302,N_19020,N_18144);
nand UO_2303 (O_2303,N_19241,N_19154);
or UO_2304 (O_2304,N_18091,N_18706);
xnor UO_2305 (O_2305,N_18991,N_19698);
and UO_2306 (O_2306,N_16951,N_16536);
or UO_2307 (O_2307,N_17462,N_19481);
xnor UO_2308 (O_2308,N_16626,N_16180);
xor UO_2309 (O_2309,N_18204,N_16359);
or UO_2310 (O_2310,N_16383,N_18658);
or UO_2311 (O_2311,N_18879,N_16433);
xor UO_2312 (O_2312,N_18900,N_18568);
nand UO_2313 (O_2313,N_18816,N_16861);
and UO_2314 (O_2314,N_16465,N_18308);
and UO_2315 (O_2315,N_19135,N_17762);
xnor UO_2316 (O_2316,N_17896,N_17431);
nand UO_2317 (O_2317,N_17823,N_16009);
xor UO_2318 (O_2318,N_19391,N_17755);
nand UO_2319 (O_2319,N_17320,N_17129);
nand UO_2320 (O_2320,N_16540,N_17096);
nor UO_2321 (O_2321,N_18889,N_16792);
nand UO_2322 (O_2322,N_16682,N_16100);
xnor UO_2323 (O_2323,N_17450,N_16056);
nand UO_2324 (O_2324,N_16365,N_17030);
nand UO_2325 (O_2325,N_18804,N_18839);
nand UO_2326 (O_2326,N_18987,N_17701);
nand UO_2327 (O_2327,N_19512,N_19611);
or UO_2328 (O_2328,N_16628,N_18927);
and UO_2329 (O_2329,N_19405,N_17251);
xor UO_2330 (O_2330,N_16026,N_16480);
nor UO_2331 (O_2331,N_19549,N_19214);
nor UO_2332 (O_2332,N_17970,N_18129);
nand UO_2333 (O_2333,N_18307,N_18148);
or UO_2334 (O_2334,N_18488,N_16805);
or UO_2335 (O_2335,N_18730,N_16496);
xor UO_2336 (O_2336,N_19953,N_19275);
and UO_2337 (O_2337,N_18998,N_18537);
and UO_2338 (O_2338,N_18612,N_18324);
nor UO_2339 (O_2339,N_19982,N_17632);
xor UO_2340 (O_2340,N_19058,N_18049);
xor UO_2341 (O_2341,N_17848,N_19145);
nand UO_2342 (O_2342,N_19217,N_19857);
nand UO_2343 (O_2343,N_17697,N_16591);
xor UO_2344 (O_2344,N_18909,N_17814);
or UO_2345 (O_2345,N_18668,N_17946);
nand UO_2346 (O_2346,N_17116,N_17461);
and UO_2347 (O_2347,N_16140,N_19393);
nor UO_2348 (O_2348,N_16207,N_18096);
or UO_2349 (O_2349,N_17357,N_17328);
nand UO_2350 (O_2350,N_19046,N_19163);
or UO_2351 (O_2351,N_16103,N_18621);
or UO_2352 (O_2352,N_17497,N_17601);
and UO_2353 (O_2353,N_17301,N_17694);
xnor UO_2354 (O_2354,N_16202,N_18502);
nor UO_2355 (O_2355,N_16419,N_18181);
nor UO_2356 (O_2356,N_19144,N_19049);
xor UO_2357 (O_2357,N_18203,N_19486);
or UO_2358 (O_2358,N_16749,N_17963);
nand UO_2359 (O_2359,N_19319,N_16757);
xnor UO_2360 (O_2360,N_17563,N_16386);
and UO_2361 (O_2361,N_17471,N_19904);
and UO_2362 (O_2362,N_16301,N_17120);
and UO_2363 (O_2363,N_19388,N_16749);
nand UO_2364 (O_2364,N_19284,N_16958);
nand UO_2365 (O_2365,N_19464,N_19863);
xnor UO_2366 (O_2366,N_16177,N_17135);
xor UO_2367 (O_2367,N_19691,N_17221);
nor UO_2368 (O_2368,N_17638,N_19960);
nand UO_2369 (O_2369,N_18093,N_18379);
nand UO_2370 (O_2370,N_18063,N_16857);
nand UO_2371 (O_2371,N_17782,N_17131);
or UO_2372 (O_2372,N_17078,N_17291);
xor UO_2373 (O_2373,N_19997,N_18895);
nor UO_2374 (O_2374,N_18656,N_16044);
nand UO_2375 (O_2375,N_16230,N_18320);
or UO_2376 (O_2376,N_19081,N_16233);
and UO_2377 (O_2377,N_19309,N_19331);
or UO_2378 (O_2378,N_16440,N_19936);
xor UO_2379 (O_2379,N_18113,N_19768);
nor UO_2380 (O_2380,N_19577,N_16125);
nand UO_2381 (O_2381,N_18327,N_17800);
nand UO_2382 (O_2382,N_18335,N_19200);
nand UO_2383 (O_2383,N_19113,N_16701);
nor UO_2384 (O_2384,N_18971,N_18246);
xor UO_2385 (O_2385,N_17382,N_19193);
nor UO_2386 (O_2386,N_16084,N_19704);
nand UO_2387 (O_2387,N_19569,N_19790);
xnor UO_2388 (O_2388,N_17390,N_19796);
and UO_2389 (O_2389,N_18817,N_19966);
nor UO_2390 (O_2390,N_16996,N_18999);
and UO_2391 (O_2391,N_19281,N_19923);
xor UO_2392 (O_2392,N_19614,N_17094);
xnor UO_2393 (O_2393,N_17712,N_19091);
or UO_2394 (O_2394,N_19166,N_18413);
and UO_2395 (O_2395,N_16854,N_17601);
and UO_2396 (O_2396,N_17121,N_19254);
or UO_2397 (O_2397,N_18943,N_16770);
or UO_2398 (O_2398,N_19860,N_17295);
xor UO_2399 (O_2399,N_18563,N_17239);
nor UO_2400 (O_2400,N_19610,N_17345);
and UO_2401 (O_2401,N_17674,N_16678);
xor UO_2402 (O_2402,N_19246,N_18812);
xnor UO_2403 (O_2403,N_18366,N_19302);
and UO_2404 (O_2404,N_19387,N_18581);
nand UO_2405 (O_2405,N_19542,N_16020);
or UO_2406 (O_2406,N_19739,N_16083);
and UO_2407 (O_2407,N_16829,N_17724);
nor UO_2408 (O_2408,N_17896,N_17973);
xnor UO_2409 (O_2409,N_19727,N_18449);
or UO_2410 (O_2410,N_17415,N_17273);
and UO_2411 (O_2411,N_18934,N_18236);
nor UO_2412 (O_2412,N_19292,N_17159);
and UO_2413 (O_2413,N_17493,N_18000);
or UO_2414 (O_2414,N_19861,N_18068);
or UO_2415 (O_2415,N_16390,N_18020);
and UO_2416 (O_2416,N_17803,N_19899);
nand UO_2417 (O_2417,N_17378,N_18296);
nor UO_2418 (O_2418,N_16706,N_18454);
nor UO_2419 (O_2419,N_17279,N_18743);
and UO_2420 (O_2420,N_16263,N_19433);
and UO_2421 (O_2421,N_19983,N_17122);
xor UO_2422 (O_2422,N_18867,N_19011);
nand UO_2423 (O_2423,N_18007,N_16171);
xnor UO_2424 (O_2424,N_19389,N_19897);
nor UO_2425 (O_2425,N_19882,N_18125);
or UO_2426 (O_2426,N_16608,N_16691);
nand UO_2427 (O_2427,N_19620,N_17786);
and UO_2428 (O_2428,N_17670,N_17800);
xnor UO_2429 (O_2429,N_18268,N_19299);
and UO_2430 (O_2430,N_19408,N_17502);
xor UO_2431 (O_2431,N_19827,N_17381);
or UO_2432 (O_2432,N_19549,N_17526);
xnor UO_2433 (O_2433,N_18221,N_18317);
nand UO_2434 (O_2434,N_16775,N_18759);
nand UO_2435 (O_2435,N_16988,N_18397);
and UO_2436 (O_2436,N_19535,N_19768);
nor UO_2437 (O_2437,N_18950,N_17979);
or UO_2438 (O_2438,N_17625,N_18014);
xnor UO_2439 (O_2439,N_19921,N_18652);
and UO_2440 (O_2440,N_16836,N_16180);
and UO_2441 (O_2441,N_17443,N_18118);
xnor UO_2442 (O_2442,N_16574,N_18612);
or UO_2443 (O_2443,N_18948,N_18770);
xor UO_2444 (O_2444,N_17104,N_18119);
and UO_2445 (O_2445,N_19980,N_17801);
or UO_2446 (O_2446,N_16453,N_16870);
and UO_2447 (O_2447,N_17663,N_18340);
and UO_2448 (O_2448,N_19256,N_19531);
xnor UO_2449 (O_2449,N_17966,N_18339);
xnor UO_2450 (O_2450,N_17515,N_16423);
nor UO_2451 (O_2451,N_18928,N_17331);
nor UO_2452 (O_2452,N_16048,N_19211);
or UO_2453 (O_2453,N_16500,N_19231);
xnor UO_2454 (O_2454,N_19246,N_18632);
or UO_2455 (O_2455,N_17963,N_17931);
or UO_2456 (O_2456,N_19238,N_17898);
xnor UO_2457 (O_2457,N_19017,N_17054);
nand UO_2458 (O_2458,N_18784,N_16836);
nand UO_2459 (O_2459,N_17380,N_17130);
or UO_2460 (O_2460,N_18862,N_18234);
or UO_2461 (O_2461,N_19590,N_17840);
xnor UO_2462 (O_2462,N_19923,N_19199);
and UO_2463 (O_2463,N_19365,N_17070);
xnor UO_2464 (O_2464,N_19564,N_19149);
nor UO_2465 (O_2465,N_18398,N_16816);
or UO_2466 (O_2466,N_17989,N_16522);
and UO_2467 (O_2467,N_16833,N_16754);
nor UO_2468 (O_2468,N_16127,N_16604);
xnor UO_2469 (O_2469,N_16062,N_17804);
xnor UO_2470 (O_2470,N_17339,N_16618);
and UO_2471 (O_2471,N_16175,N_17878);
nor UO_2472 (O_2472,N_17535,N_17364);
nand UO_2473 (O_2473,N_17801,N_19197);
nor UO_2474 (O_2474,N_17756,N_17516);
or UO_2475 (O_2475,N_16636,N_17776);
and UO_2476 (O_2476,N_17737,N_17262);
nand UO_2477 (O_2477,N_18065,N_18290);
or UO_2478 (O_2478,N_18423,N_18127);
nor UO_2479 (O_2479,N_16022,N_17147);
and UO_2480 (O_2480,N_17517,N_19873);
and UO_2481 (O_2481,N_18254,N_18828);
and UO_2482 (O_2482,N_18850,N_19356);
nand UO_2483 (O_2483,N_18263,N_16892);
and UO_2484 (O_2484,N_19658,N_16606);
xor UO_2485 (O_2485,N_19129,N_17284);
and UO_2486 (O_2486,N_18161,N_19336);
xor UO_2487 (O_2487,N_17997,N_19828);
nand UO_2488 (O_2488,N_18226,N_17337);
nand UO_2489 (O_2489,N_17815,N_16395);
nor UO_2490 (O_2490,N_19116,N_17452);
nand UO_2491 (O_2491,N_18754,N_17214);
nor UO_2492 (O_2492,N_19471,N_19718);
or UO_2493 (O_2493,N_19209,N_19618);
nor UO_2494 (O_2494,N_19898,N_18109);
xor UO_2495 (O_2495,N_19100,N_17904);
nor UO_2496 (O_2496,N_19054,N_17305);
and UO_2497 (O_2497,N_16665,N_17174);
nand UO_2498 (O_2498,N_19407,N_17575);
nor UO_2499 (O_2499,N_18129,N_16523);
endmodule